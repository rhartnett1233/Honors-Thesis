module AND2_X1( A1, A2, ZN );
  input A1;
  input A2;
  //input_done

  output ZN;
  //output_done

  //wire_done

  assign ZN = A1 & A2;
endmodule


module OR2_X1( A1, A2, ZN );
  input A1;
  input A2;
  //input_done

  output ZN;
  //output_done

  //wire_done

  assign ZN = A1 | A2;
endmodule

module INV_X1( A, ZN );
  input A;
  //input_done

  output ZN;
  //output_done

  //wire_done
  
  assign ZN = ~A;
endmodule

module scale2_0 ( in, inbar, out, outbar );

  input wire [7:0] in;
  input wire [7:0] inbar;
//input_done

  output wire [7:0] out;
  output wire [7:0] outbar;
//output_done

  wire in_0;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_1;
  wire in_7;
  wire n11;
  wire n12;
  wire n13;
  wire n14;
  wire n15;
  wire n16;
  wire n17;
  wire n18;
  wire n19;
  wire n20;
  wire in_0bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_1bar;
  wire in_7bar;
  wire n11bar;
  wire n12bar;
  wire n13bar;
  wire n14bar;
  wire n15bar;
  wire n16bar;
  wire n17bar;
  wire n18bar;
  wire n19bar;
  wire n20bar;
//wire_done

  assign in_0 = in[0];
  assign out[7] = in_6;
  assign in_6  = in[6];
  assign out[6] = in_5;
  assign in_5  = in[5];
  assign out[5] = in_4;
  assign in_4  = in[4];
  assign out[2] = in_1;
  assign in_1  = in[1];
  assign out[0] = in_7;
  assign in_7  = in[7];
  assign in_0bar = inbar[0];
  assign outbar[7] = in_6bar;
  assign in_6bar = inbar[6];
  assign outbar[6] = in_5bar;
  assign in_5bar = inbar[5];
  assign outbar[5] = in_4bar;
  assign in_4bar = inbar[4];
  assign outbar[2] = in_1bar;
  assign in_1bar = inbar[1];
  assign outbar[0] = in_7bar;
  assign in_7bar = inbar[7];
//assign_done

  assign n20bar = in_7;
  assign n20 = in_7bar;
  assign n19bar = in[3];
  assign n19 = inbar[3];
  assign n18bar = in[2];
  assign n18 = inbar[2];
  assign n17bar = in_0;
  assign n17 = in_0bar;
  OR2_X1 U5 ( .A1(n16), .A2(n15), .ZN(out[4]) );
  AND2_X1 U5bar ( .A1(n16bar), .A2(n15bar), .ZN(outbar[4]) );
  AND2_X1 U6 ( .A1(in[3]), .A2(n20), .ZN(n15) );
  OR2_X1 U6bar ( .A1(inbar[3]), .A2(n20bar), .ZN(n15bar) );
  AND2_X1 U7 ( .A1(in_7), .A2(n19), .ZN(n16) );
  OR2_X1 U7bar ( .A1(in_7bar), .A2(n19bar), .ZN(n16bar) );
  OR2_X1 U8 ( .A1(n14), .A2(n13), .ZN(out[3]) );
  AND2_X1 U8bar ( .A1(n14bar), .A2(n13bar), .ZN(outbar[3]) );
  AND2_X1 U9 ( .A1(in[2]), .A2(n20), .ZN(n13) );
  OR2_X1 U9bar ( .A1(inbar[2]), .A2(n20bar), .ZN(n13bar) );
  AND2_X1 U10 ( .A1(in_7), .A2(n18), .ZN(n14) );
  OR2_X1 U10bar ( .A1(in_7bar), .A2(n18bar), .ZN(n14bar) );
  OR2_X1 U11 ( .A1(n12), .A2(n11), .ZN(out[1]) );
  AND2_X1 U11bar ( .A1(n12bar), .A2(n11bar), .ZN(outbar[1]) );
  AND2_X1 U12 ( .A1(in_0), .A2(n20), .ZN(n11) );
  OR2_X1 U12bar ( .A1(in_0bar), .A2(n20bar), .ZN(n11bar) );
  AND2_X1 U13 ( .A1(in_7), .A2(n17), .ZN(n12) );
  OR2_X1 U13bar ( .A1(in_7bar), .A2(n17bar), .ZN(n12bar) );
endmodule

module byteXor_0 ( a, abar, b, bbar, y, ybar );

  input wire [7:0] a;
  input wire [7:0] b;
  input wire [7:0] abar;
  input wire [7:0] bbar;
//input_done

  output wire [7:0] y;
  output wire [7:0] ybar;
//output_done

  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n33bar;
  wire n34bar;
  wire n35bar;
  wire n36bar;
  wire n37bar;
  wire n38bar;
  wire n39bar;
  wire n40bar;
  wire n41bar;
  wire n42bar;
  wire n43bar;
  wire n44bar;
  wire n45bar;
  wire n46bar;
  wire n47bar;
  wire n48bar;
  wire n49bar;
  wire n50bar;
  wire n51bar;
  wire n52bar;
  wire n53bar;
  wire n54bar;
  wire n55bar;
  wire n56bar;
  wire n57bar;
  wire n58bar;
  wire n59bar;
  wire n60bar;
  wire n61bar;
  wire n62bar;
  wire n63bar;
  wire n64bar;
//wire_done

 //assign_done

  assign n64bar = n47;
  assign n64 = n47bar;
  assign n63bar = a[7];
  assign n63 = abar[7];
  assign n62bar = n45;
  assign n62 = n45bar;
  assign n61bar = a[6];
  assign n61 = abar[6];
  assign n60bar = n43;
  assign n60 = n43bar;
  assign n59bar = a[5];
  assign n59 = abar[5];
  assign n58bar = n41;
  assign n58 = n41bar;
  assign n57bar = a[4];
  assign n57 = abar[4];
  assign n56bar = n39;
  assign n56 = n39bar;
  assign n55bar = a[3];
  assign n55 = abar[3];
  assign n54bar = n37;
  assign n54 = n37bar;
  assign n53bar = a[2];
  assign n53 = abar[2];
  assign n52bar = n35;
  assign n52 = n35bar;
  assign n51bar = a[1];
  assign n51 = abar[1];
  assign n50bar = n33;
  assign n50 = n33bar;
  assign n49bar = a[0];
  assign n49 = abar[0];
  OR2_X1 U17 ( .A1(n48), .A2(n64), .ZN(y[7]) );
  AND2_X1 U17bar ( .A1(n48bar), .A2(n64bar), .ZN(ybar[7]) );
  OR2_X1 U18 ( .A1(n63), .A2(b[7]), .ZN(n47) );
  AND2_X1 U18bar ( .A1(n63bar), .A2(bbar[7]), .ZN(n47bar) );
  AND2_X1 U19 ( .A1(b[7]), .A2(n63), .ZN(n48) );
  OR2_X1 U19bar ( .A1(bbar[7]), .A2(n63bar), .ZN(n48bar) );
  OR2_X1 U20 ( .A1(n46), .A2(n62), .ZN(y[6]) );
  AND2_X1 U20bar ( .A1(n46bar), .A2(n62bar), .ZN(ybar[6]) );
  OR2_X1 U21 ( .A1(n61), .A2(b[6]), .ZN(n45) );
  AND2_X1 U21bar ( .A1(n61bar), .A2(bbar[6]), .ZN(n45bar) );
  AND2_X1 U22 ( .A1(b[6]), .A2(n61), .ZN(n46) );
  OR2_X1 U22bar ( .A1(bbar[6]), .A2(n61bar), .ZN(n46bar) );
  OR2_X1 U23 ( .A1(n44), .A2(n60), .ZN(y[5]) );
  AND2_X1 U23bar ( .A1(n44bar), .A2(n60bar), .ZN(ybar[5]) );
  OR2_X1 U24 ( .A1(n59), .A2(b[5]), .ZN(n43) );
  AND2_X1 U24bar ( .A1(n59bar), .A2(bbar[5]), .ZN(n43bar) );
  AND2_X1 U25 ( .A1(b[5]), .A2(n59), .ZN(n44) );
  OR2_X1 U25bar ( .A1(bbar[5]), .A2(n59bar), .ZN(n44bar) );
  OR2_X1 U26 ( .A1(n42), .A2(n58), .ZN(y[4]) );
  AND2_X1 U26bar ( .A1(n42bar), .A2(n58bar), .ZN(ybar[4]) );
  OR2_X1 U27 ( .A1(n57), .A2(b[4]), .ZN(n41) );
  AND2_X1 U27bar ( .A1(n57bar), .A2(bbar[4]), .ZN(n41bar) );
  AND2_X1 U28 ( .A1(b[4]), .A2(n57), .ZN(n42) );
  OR2_X1 U28bar ( .A1(bbar[4]), .A2(n57bar), .ZN(n42bar) );
  OR2_X1 U29 ( .A1(n40), .A2(n56), .ZN(y[3]) );
  AND2_X1 U29bar ( .A1(n40bar), .A2(n56bar), .ZN(ybar[3]) );
  OR2_X1 U30 ( .A1(n55), .A2(b[3]), .ZN(n39) );
  AND2_X1 U30bar ( .A1(n55bar), .A2(bbar[3]), .ZN(n39bar) );
  AND2_X1 U31 ( .A1(b[3]), .A2(n55), .ZN(n40) );
  OR2_X1 U31bar ( .A1(bbar[3]), .A2(n55bar), .ZN(n40bar) );
  OR2_X1 U32 ( .A1(n38), .A2(n54), .ZN(y[2]) );
  AND2_X1 U32bar ( .A1(n38bar), .A2(n54bar), .ZN(ybar[2]) );
  OR2_X1 U33 ( .A1(n53), .A2(b[2]), .ZN(n37) );
  AND2_X1 U33bar ( .A1(n53bar), .A2(bbar[2]), .ZN(n37bar) );
  AND2_X1 U34 ( .A1(b[2]), .A2(n53), .ZN(n38) );
  OR2_X1 U34bar ( .A1(bbar[2]), .A2(n53bar), .ZN(n38bar) );
  OR2_X1 U35 ( .A1(n36), .A2(n52), .ZN(y[1]) );
  AND2_X1 U35bar ( .A1(n36bar), .A2(n52bar), .ZN(ybar[1]) );
  OR2_X1 U36 ( .A1(n51), .A2(b[1]), .ZN(n35) );
  AND2_X1 U36bar ( .A1(n51bar), .A2(bbar[1]), .ZN(n35bar) );
  AND2_X1 U37 ( .A1(b[1]), .A2(n51), .ZN(n36) );
  OR2_X1 U37bar ( .A1(bbar[1]), .A2(n51bar), .ZN(n36bar) );
  OR2_X1 U38 ( .A1(n34), .A2(n50), .ZN(y[0]) );
  AND2_X1 U38bar ( .A1(n34bar), .A2(n50bar), .ZN(ybar[0]) );
  OR2_X1 U39 ( .A1(n49), .A2(b[0]), .ZN(n33) );
  AND2_X1 U39bar ( .A1(n49bar), .A2(bbar[0]), .ZN(n33bar) );
  AND2_X1 U40 ( .A1(b[0]), .A2(n49), .ZN(n34) );
  OR2_X1 U40bar ( .A1(bbar[0]), .A2(n49bar), .ZN(n34bar) );
endmodule

module byteXor4_0 ( a, abar, b, bbar, c, cbar, d, dbar, y, ybar );

  input wire [7:0] a;
  input wire [7:0] b;
  input wire [7:0] c;
  input wire [7:0] d;
  input wire [7:0] abar;
  input wire [7:0] bbar;
  input wire [7:0] cbar;
  input wire [7:0] dbar;
//input_done

  output wire [7:0] y;
  output wire [7:0] ybar;
//output_done

  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n113bar;
  wire n114bar;
  wire n115bar;
  wire n116bar;
  wire n117bar;
  wire n118bar;
  wire n119bar;
  wire n120bar;
  wire n121bar;
  wire n122bar;
  wire n123bar;
  wire n124bar;
  wire n125bar;
  wire n126bar;
  wire n127bar;
  wire n128bar;
  wire n129bar;
  wire n130bar;
  wire n131bar;
  wire n132bar;
  wire n133bar;
  wire n134bar;
  wire n135bar;
  wire n136bar;
  wire n137bar;
  wire n138bar;
  wire n139bar;
  wire n140bar;
  wire n141bar;
  wire n142bar;
  wire n143bar;
  wire n144bar;
  wire n145bar;
  wire n146bar;
  wire n147bar;
  wire n148bar;
  wire n149bar;
  wire n150bar;
  wire n151bar;
  wire n152bar;
  wire n153bar;
  wire n154bar;
  wire n155bar;
  wire n156bar;
  wire n157bar;
  wire n158bar;
  wire n159bar;
  wire n160bar;
  wire n161bar;
  wire n162bar;
  wire n163bar;
  wire n164bar;
  wire n165bar;
  wire n166bar;
  wire n167bar;
  wire n168bar;
  wire n169bar;
  wire n170bar;
  wire n171bar;
  wire n172bar;
  wire n173bar;
  wire n174bar;
  wire n175bar;
  wire n176bar;
  wire n177bar;
  wire n178bar;
  wire n179bar;
  wire n180bar;
  wire n181bar;
  wire n182bar;
  wire n183bar;
  wire n184bar;
  wire n185bar;
  wire n186bar;
  wire n187bar;
  wire n188bar;
  wire n189bar;
  wire n190bar;
  wire n191bar;
  wire n192bar;
  wire n193bar;
  wire n194bar;
  wire n195bar;
  wire n196bar;
  wire n197bar;
  wire n198bar;
  wire n199bar;
  wire n200bar;
  wire n201bar;
  wire n202bar;
  wire n203bar;
  wire n204bar;
  wire n205bar;
  wire n206bar;
  wire n207bar;
  wire n208bar;
  wire n209bar;
  wire n210bar;
  wire n211bar;
  wire n212bar;
  wire n213bar;
  wire n214bar;
  wire n215bar;
  wire n216bar;
  wire n217bar;
  wire n218bar;
  wire n219bar;
  wire n220bar;
  wire n221bar;
  wire n222bar;
  wire n223bar;
  wire n224bar;
//wire_done

 //assign_done

  assign n224bar = n175;
  assign n224 = n175bar;
  assign n223bar = a[7];
  assign n223 = abar[7];
  assign n222bar = n167;
  assign n222 = n167bar;
  assign n221bar = a[6];
  assign n221 = abar[6];
  assign n220bar = n159;
  assign n220 = n159bar;
  assign n219bar = a[5];
  assign n219 = abar[5];
  assign n218bar = n151;
  assign n218 = n151bar;
  assign n217bar = a[4];
  assign n217 = abar[4];
  assign n216bar = n143;
  assign n216 = n143bar;
  assign n215bar = a[3];
  assign n215 = abar[3];
  assign n214bar = n135;
  assign n214 = n135bar;
  assign n213bar = a[2];
  assign n213 = abar[2];
  assign n212bar = n127;
  assign n212 = n127bar;
  assign n211bar = a[1];
  assign n211 = abar[1];
  assign n210bar = n119;
  assign n210 = n119bar;
  assign n209bar = a[0];
  assign n209 = abar[0];
  assign n208bar = b[7];
  assign n208 = bbar[7];
  assign n207bar = b[6];
  assign n207 = bbar[6];
  assign n206bar = b[5];
  assign n206 = bbar[5];
  assign n205bar = b[4];
  assign n205 = bbar[4];
  assign n204bar = b[3];
  assign n204 = bbar[3];
  assign n203bar = b[2];
  assign n203 = bbar[2];
  assign n202bar = b[1];
  assign n202 = bbar[1];
  assign n201bar = b[0];
  assign n201 = bbar[0];
  assign n200bar = n171;
  assign n200 = n171bar;
  assign n199bar = c[7];
  assign n199 = cbar[7];
  assign n198bar = n163;
  assign n198 = n163bar;
  assign n197bar = c[6];
  assign n197 = cbar[6];
  assign n196bar = n155;
  assign n196 = n155bar;
  assign n195bar = c[5];
  assign n195 = cbar[5];
  assign n194bar = n147;
  assign n194 = n147bar;
  assign n193bar = c[4];
  assign n193 = cbar[4];
  assign n192bar = n139;
  assign n192 = n139bar;
  assign n191bar = c[3];
  assign n191 = cbar[3];
  assign n190bar = n131;
  assign n190 = n131bar;
  assign n189bar = c[2];
  assign n189 = cbar[2];
  assign n188bar = n123;
  assign n188 = n123bar;
  assign n187bar = c[1];
  assign n187 = cbar[1];
  assign n186bar = n115;
  assign n186 = n115bar;
  assign n185bar = c[0];
  assign n185 = cbar[0];
  assign n184bar = d[7];
  assign n184 = dbar[7];
  assign n183bar = d[6];
  assign n183 = dbar[6];
  assign n182bar = d[5];
  assign n182 = dbar[5];
  assign n181bar = d[4];
  assign n181 = dbar[4];
  assign n180bar = d[3];
  assign n180 = dbar[3];
  assign n179bar = d[2];
  assign n179 = dbar[2];
  assign n178bar = d[1];
  assign n178 = dbar[1];
  assign n177bar = d[0];
  assign n177 = dbar[0];
  OR2_X1 U49 ( .A1(n176), .A2(n224), .ZN(y[7]) );
  AND2_X1 U49bar ( .A1(n176bar), .A2(n224bar), .ZN(ybar[7]) );
  OR2_X1 U50 ( .A1(n174), .A2(n200), .ZN(n175) );
  AND2_X1 U50bar ( .A1(n174bar), .A2(n200bar), .ZN(n175bar) );
  AND2_X1 U51 ( .A1(n200), .A2(n174), .ZN(n176) );
  OR2_X1 U51bar ( .A1(n200bar), .A2(n174bar), .ZN(n176bar) );
  AND2_X1 U52 ( .A1(n173), .A2(n172), .ZN(n174) );
  OR2_X1 U52bar ( .A1(n173bar), .A2(n172bar), .ZN(n174bar) );
  OR2_X1 U53 ( .A1(n223), .A2(b[7]), .ZN(n172) );
  AND2_X1 U53bar ( .A1(n223bar), .A2(bbar[7]), .ZN(n172bar) );
  OR2_X1 U54 ( .A1(n208), .A2(a[7]), .ZN(n173) );
  AND2_X1 U54bar ( .A1(n208bar), .A2(abar[7]), .ZN(n173bar) );
  AND2_X1 U55 ( .A1(n170), .A2(n169), .ZN(n171) );
  OR2_X1 U55bar ( .A1(n170bar), .A2(n169bar), .ZN(n171bar) );
  OR2_X1 U56 ( .A1(n199), .A2(d[7]), .ZN(n169) );
  AND2_X1 U56bar ( .A1(n199bar), .A2(dbar[7]), .ZN(n169bar) );
  OR2_X1 U57 ( .A1(n184), .A2(c[7]), .ZN(n170) );
  AND2_X1 U57bar ( .A1(n184bar), .A2(cbar[7]), .ZN(n170bar) );
  OR2_X1 U58 ( .A1(n168), .A2(n222), .ZN(y[6]) );
  AND2_X1 U58bar ( .A1(n168bar), .A2(n222bar), .ZN(ybar[6]) );
  OR2_X1 U59 ( .A1(n166), .A2(n198), .ZN(n167) );
  AND2_X1 U59bar ( .A1(n166bar), .A2(n198bar), .ZN(n167bar) );
  AND2_X1 U60 ( .A1(n198), .A2(n166), .ZN(n168) );
  OR2_X1 U60bar ( .A1(n198bar), .A2(n166bar), .ZN(n168bar) );
  AND2_X1 U61 ( .A1(n165), .A2(n164), .ZN(n166) );
  OR2_X1 U61bar ( .A1(n165bar), .A2(n164bar), .ZN(n166bar) );
  OR2_X1 U62 ( .A1(n221), .A2(b[6]), .ZN(n164) );
  AND2_X1 U62bar ( .A1(n221bar), .A2(bbar[6]), .ZN(n164bar) );
  OR2_X1 U63 ( .A1(n207), .A2(a[6]), .ZN(n165) );
  AND2_X1 U63bar ( .A1(n207bar), .A2(abar[6]), .ZN(n165bar) );
  AND2_X1 U64 ( .A1(n162), .A2(n161), .ZN(n163) );
  OR2_X1 U64bar ( .A1(n162bar), .A2(n161bar), .ZN(n163bar) );
  OR2_X1 U65 ( .A1(n197), .A2(d[6]), .ZN(n161) );
  AND2_X1 U65bar ( .A1(n197bar), .A2(dbar[6]), .ZN(n161bar) );
  OR2_X1 U66 ( .A1(n183), .A2(c[6]), .ZN(n162) );
  AND2_X1 U66bar ( .A1(n183bar), .A2(cbar[6]), .ZN(n162bar) );
  OR2_X1 U67 ( .A1(n160), .A2(n220), .ZN(y[5]) );
  AND2_X1 U67bar ( .A1(n160bar), .A2(n220bar), .ZN(ybar[5]) );
  OR2_X1 U68 ( .A1(n158), .A2(n196), .ZN(n159) );
  AND2_X1 U68bar ( .A1(n158bar), .A2(n196bar), .ZN(n159bar) );
  AND2_X1 U69 ( .A1(n196), .A2(n158), .ZN(n160) );
  OR2_X1 U69bar ( .A1(n196bar), .A2(n158bar), .ZN(n160bar) );
  AND2_X1 U70 ( .A1(n157), .A2(n156), .ZN(n158) );
  OR2_X1 U70bar ( .A1(n157bar), .A2(n156bar), .ZN(n158bar) );
  OR2_X1 U71 ( .A1(n219), .A2(b[5]), .ZN(n156) );
  AND2_X1 U71bar ( .A1(n219bar), .A2(bbar[5]), .ZN(n156bar) );
  OR2_X1 U72 ( .A1(n206), .A2(a[5]), .ZN(n157) );
  AND2_X1 U72bar ( .A1(n206bar), .A2(abar[5]), .ZN(n157bar) );
  AND2_X1 U73 ( .A1(n154), .A2(n153), .ZN(n155) );
  OR2_X1 U73bar ( .A1(n154bar), .A2(n153bar), .ZN(n155bar) );
  OR2_X1 U74 ( .A1(n195), .A2(d[5]), .ZN(n153) );
  AND2_X1 U74bar ( .A1(n195bar), .A2(dbar[5]), .ZN(n153bar) );
  OR2_X1 U75 ( .A1(n182), .A2(c[5]), .ZN(n154) );
  AND2_X1 U75bar ( .A1(n182bar), .A2(cbar[5]), .ZN(n154bar) );
  OR2_X1 U76 ( .A1(n152), .A2(n218), .ZN(y[4]) );
  AND2_X1 U76bar ( .A1(n152bar), .A2(n218bar), .ZN(ybar[4]) );
  OR2_X1 U77 ( .A1(n150), .A2(n194), .ZN(n151) );
  AND2_X1 U77bar ( .A1(n150bar), .A2(n194bar), .ZN(n151bar) );
  AND2_X1 U78 ( .A1(n194), .A2(n150), .ZN(n152) );
  OR2_X1 U78bar ( .A1(n194bar), .A2(n150bar), .ZN(n152bar) );
  AND2_X1 U79 ( .A1(n149), .A2(n148), .ZN(n150) );
  OR2_X1 U79bar ( .A1(n149bar), .A2(n148bar), .ZN(n150bar) );
  OR2_X1 U80 ( .A1(n217), .A2(b[4]), .ZN(n148) );
  AND2_X1 U80bar ( .A1(n217bar), .A2(bbar[4]), .ZN(n148bar) );
  OR2_X1 U81 ( .A1(n205), .A2(a[4]), .ZN(n149) );
  AND2_X1 U81bar ( .A1(n205bar), .A2(abar[4]), .ZN(n149bar) );
  AND2_X1 U82 ( .A1(n146), .A2(n145), .ZN(n147) );
  OR2_X1 U82bar ( .A1(n146bar), .A2(n145bar), .ZN(n147bar) );
  OR2_X1 U83 ( .A1(n193), .A2(d[4]), .ZN(n145) );
  AND2_X1 U83bar ( .A1(n193bar), .A2(dbar[4]), .ZN(n145bar) );
  OR2_X1 U84 ( .A1(n181), .A2(c[4]), .ZN(n146) );
  AND2_X1 U84bar ( .A1(n181bar), .A2(cbar[4]), .ZN(n146bar) );
  OR2_X1 U85 ( .A1(n144), .A2(n216), .ZN(y[3]) );
  AND2_X1 U85bar ( .A1(n144bar), .A2(n216bar), .ZN(ybar[3]) );
  OR2_X1 U86 ( .A1(n142), .A2(n192), .ZN(n143) );
  AND2_X1 U86bar ( .A1(n142bar), .A2(n192bar), .ZN(n143bar) );
  AND2_X1 U87 ( .A1(n192), .A2(n142), .ZN(n144) );
  OR2_X1 U87bar ( .A1(n192bar), .A2(n142bar), .ZN(n144bar) );
  AND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(n142) );
  OR2_X1 U88bar ( .A1(n141bar), .A2(n140bar), .ZN(n142bar) );
  OR2_X1 U89 ( .A1(n215), .A2(b[3]), .ZN(n140) );
  AND2_X1 U89bar ( .A1(n215bar), .A2(bbar[3]), .ZN(n140bar) );
  OR2_X1 U90 ( .A1(n204), .A2(a[3]), .ZN(n141) );
  AND2_X1 U90bar ( .A1(n204bar), .A2(abar[3]), .ZN(n141bar) );
  AND2_X1 U91 ( .A1(n138), .A2(n137), .ZN(n139) );
  OR2_X1 U91bar ( .A1(n138bar), .A2(n137bar), .ZN(n139bar) );
  OR2_X1 U92 ( .A1(n191), .A2(d[3]), .ZN(n137) );
  AND2_X1 U92bar ( .A1(n191bar), .A2(dbar[3]), .ZN(n137bar) );
  OR2_X1 U93 ( .A1(n180), .A2(c[3]), .ZN(n138) );
  AND2_X1 U93bar ( .A1(n180bar), .A2(cbar[3]), .ZN(n138bar) );
  OR2_X1 U94 ( .A1(n136), .A2(n214), .ZN(y[2]) );
  AND2_X1 U94bar ( .A1(n136bar), .A2(n214bar), .ZN(ybar[2]) );
  OR2_X1 U95 ( .A1(n134), .A2(n190), .ZN(n135) );
  AND2_X1 U95bar ( .A1(n134bar), .A2(n190bar), .ZN(n135bar) );
  AND2_X1 U96 ( .A1(n190), .A2(n134), .ZN(n136) );
  OR2_X1 U96bar ( .A1(n190bar), .A2(n134bar), .ZN(n136bar) );
  AND2_X1 U97 ( .A1(n133), .A2(n132), .ZN(n134) );
  OR2_X1 U97bar ( .A1(n133bar), .A2(n132bar), .ZN(n134bar) );
  OR2_X1 U98 ( .A1(n213), .A2(b[2]), .ZN(n132) );
  AND2_X1 U98bar ( .A1(n213bar), .A2(bbar[2]), .ZN(n132bar) );
  OR2_X1 U99 ( .A1(n203), .A2(a[2]), .ZN(n133) );
  AND2_X1 U99bar ( .A1(n203bar), .A2(abar[2]), .ZN(n133bar) );
  AND2_X1 U100 ( .A1(n130), .A2(n129), .ZN(n131) );
  OR2_X1 U100bar ( .A1(n130bar), .A2(n129bar), .ZN(n131bar) );
  OR2_X1 U101 ( .A1(n189), .A2(d[2]), .ZN(n129) );
  AND2_X1 U101bar ( .A1(n189bar), .A2(dbar[2]), .ZN(n129bar) );
  OR2_X1 U102 ( .A1(n179), .A2(c[2]), .ZN(n130) );
  AND2_X1 U102bar ( .A1(n179bar), .A2(cbar[2]), .ZN(n130bar) );
  OR2_X1 U103 ( .A1(n128), .A2(n212), .ZN(y[1]) );
  AND2_X1 U103bar ( .A1(n128bar), .A2(n212bar), .ZN(ybar[1]) );
  OR2_X1 U104 ( .A1(n126), .A2(n188), .ZN(n127) );
  AND2_X1 U104bar ( .A1(n126bar), .A2(n188bar), .ZN(n127bar) );
  AND2_X1 U105 ( .A1(n188), .A2(n126), .ZN(n128) );
  OR2_X1 U105bar ( .A1(n188bar), .A2(n126bar), .ZN(n128bar) );
  AND2_X1 U106 ( .A1(n125), .A2(n124), .ZN(n126) );
  OR2_X1 U106bar ( .A1(n125bar), .A2(n124bar), .ZN(n126bar) );
  OR2_X1 U107 ( .A1(n211), .A2(b[1]), .ZN(n124) );
  AND2_X1 U107bar ( .A1(n211bar), .A2(bbar[1]), .ZN(n124bar) );
  OR2_X1 U108 ( .A1(n202), .A2(a[1]), .ZN(n125) );
  AND2_X1 U108bar ( .A1(n202bar), .A2(abar[1]), .ZN(n125bar) );
  AND2_X1 U109 ( .A1(n122), .A2(n121), .ZN(n123) );
  OR2_X1 U109bar ( .A1(n122bar), .A2(n121bar), .ZN(n123bar) );
  OR2_X1 U110 ( .A1(n187), .A2(d[1]), .ZN(n121) );
  AND2_X1 U110bar ( .A1(n187bar), .A2(dbar[1]), .ZN(n121bar) );
  OR2_X1 U111 ( .A1(n178), .A2(c[1]), .ZN(n122) );
  AND2_X1 U111bar ( .A1(n178bar), .A2(cbar[1]), .ZN(n122bar) );
  OR2_X1 U112 ( .A1(n120), .A2(n210), .ZN(y[0]) );
  AND2_X1 U112bar ( .A1(n120bar), .A2(n210bar), .ZN(ybar[0]) );
  OR2_X1 U113 ( .A1(n118), .A2(n186), .ZN(n119) );
  AND2_X1 U113bar ( .A1(n118bar), .A2(n186bar), .ZN(n119bar) );
  AND2_X1 U114 ( .A1(n186), .A2(n118), .ZN(n120) );
  OR2_X1 U114bar ( .A1(n186bar), .A2(n118bar), .ZN(n120bar) );
  AND2_X1 U115 ( .A1(n117), .A2(n116), .ZN(n118) );
  OR2_X1 U115bar ( .A1(n117bar), .A2(n116bar), .ZN(n118bar) );
  OR2_X1 U116 ( .A1(n209), .A2(b[0]), .ZN(n116) );
  AND2_X1 U116bar ( .A1(n209bar), .A2(bbar[0]), .ZN(n116bar) );
  OR2_X1 U117 ( .A1(n201), .A2(a[0]), .ZN(n117) );
  AND2_X1 U117bar ( .A1(n201bar), .A2(abar[0]), .ZN(n117bar) );
  AND2_X1 U118 ( .A1(n114), .A2(n113), .ZN(n115) );
  OR2_X1 U118bar ( .A1(n114bar), .A2(n113bar), .ZN(n115bar) );
  OR2_X1 U119 ( .A1(n185), .A2(d[0]), .ZN(n113) );
  AND2_X1 U119bar ( .A1(n185bar), .A2(dbar[0]), .ZN(n113bar) );
  OR2_X1 U120 ( .A1(n177), .A2(c[0]), .ZN(n114) );
  AND2_X1 U120bar ( .A1(n177bar), .A2(cbar[0]), .ZN(n114bar) );
endmodule

module scale2_13 ( in, inbar, out, outbar );

  input wire [7:0] in;
  input wire [7:0] inbar;
//input_done

  output wire [7:0] out;
  output wire [7:0] outbar;
//output_done

  wire in_0;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_1;
  wire in_7;
  wire n11;
  wire n12;
  wire n13;
  wire n14;
  wire n15;
  wire n16;
  wire n17;
  wire n18;
  wire n19;
  wire n20;
  wire in_0bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_1bar;
  wire in_7bar;
  wire n11bar;
  wire n12bar;
  wire n13bar;
  wire n14bar;
  wire n15bar;
  wire n16bar;
  wire n17bar;
  wire n18bar;
  wire n19bar;
  wire n20bar;
//wire_done

  assign in_0 = in[0];
  assign out[7] = in_6;
  assign in_6  = in[6];
  assign out[6] = in_5;
  assign in_5  = in[5];
  assign out[5] = in_4;
  assign in_4  = in[4];
  assign out[2] = in_1;
  assign in_1  = in[1];
  assign out[0] = in_7;
  assign in_7  = in[7];
  assign in_0bar = inbar[0];
  assign outbar[7] = in_6bar;
  assign in_6bar = inbar[6];
  assign outbar[6] = in_5bar;
  assign in_5bar = inbar[5];
  assign outbar[5] = in_4bar;
  assign in_4bar = inbar[4];
  assign outbar[2] = in_1bar;
  assign in_1bar = inbar[1];
  assign outbar[0] = in_7bar;
  assign in_7bar = inbar[7];
//assign_done

  assign n20bar = in_7;
  assign n20 = in_7bar;
  assign n19bar = in[3];
  assign n19 = inbar[3];
  assign n18bar = in[2];
  assign n18 = inbar[2];
  assign n17bar = in_0;
  assign n17 = in_0bar;
  OR2_X1 U5 ( .A1(n16), .A2(n15), .ZN(out[4]) );
  AND2_X1 U5bar ( .A1(n16bar), .A2(n15bar), .ZN(outbar[4]) );
  AND2_X1 U6 ( .A1(in[3]), .A2(n20), .ZN(n15) );
  OR2_X1 U6bar ( .A1(inbar[3]), .A2(n20bar), .ZN(n15bar) );
  AND2_X1 U7 ( .A1(in_7), .A2(n19), .ZN(n16) );
  OR2_X1 U7bar ( .A1(in_7bar), .A2(n19bar), .ZN(n16bar) );
  OR2_X1 U8 ( .A1(n14), .A2(n13), .ZN(out[3]) );
  AND2_X1 U8bar ( .A1(n14bar), .A2(n13bar), .ZN(outbar[3]) );
  AND2_X1 U9 ( .A1(in[2]), .A2(n20), .ZN(n13) );
  OR2_X1 U9bar ( .A1(inbar[2]), .A2(n20bar), .ZN(n13bar) );
  AND2_X1 U10 ( .A1(in_7), .A2(n18), .ZN(n14) );
  OR2_X1 U10bar ( .A1(in_7bar), .A2(n18bar), .ZN(n14bar) );
  OR2_X1 U11 ( .A1(n12), .A2(n11), .ZN(out[1]) );
  AND2_X1 U11bar ( .A1(n12bar), .A2(n11bar), .ZN(outbar[1]) );
  AND2_X1 U12 ( .A1(in_0), .A2(n20), .ZN(n11) );
  OR2_X1 U12bar ( .A1(in_0bar), .A2(n20bar), .ZN(n11bar) );
  AND2_X1 U13 ( .A1(in_7), .A2(n17), .ZN(n12) );
  OR2_X1 U13bar ( .A1(in_7bar), .A2(n17bar), .ZN(n12bar) );
endmodule

module scale2_14 ( in, inbar, out, outbar );

  input wire [7:0] in;
  input wire [7:0] inbar;
//input_done

  output wire [7:0] out;
  output wire [7:0] outbar;
//output_done

  wire in_0;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_1;
  wire in_7;
  wire n11;
  wire n12;
  wire n13;
  wire n14;
  wire n15;
  wire n16;
  wire n17;
  wire n18;
  wire n19;
  wire n20;
  wire in_0bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_1bar;
  wire in_7bar;
  wire n11bar;
  wire n12bar;
  wire n13bar;
  wire n14bar;
  wire n15bar;
  wire n16bar;
  wire n17bar;
  wire n18bar;
  wire n19bar;
  wire n20bar;
//wire_done

  assign in_0 = in[0];
  assign out[7] = in_6;
  assign in_6  = in[6];
  assign out[6] = in_5;
  assign in_5  = in[5];
  assign out[5] = in_4;
  assign in_4  = in[4];
  assign out[2] = in_1;
  assign in_1  = in[1];
  assign out[0] = in_7;
  assign in_7  = in[7];
  assign in_0bar = inbar[0];
  assign outbar[7] = in_6bar;
  assign in_6bar = inbar[6];
  assign outbar[6] = in_5bar;
  assign in_5bar = inbar[5];
  assign outbar[5] = in_4bar;
  assign in_4bar = inbar[4];
  assign outbar[2] = in_1bar;
  assign in_1bar = inbar[1];
  assign outbar[0] = in_7bar;
  assign in_7bar = inbar[7];
//assign_done

  assign n20bar = in_7;
  assign n20 = in_7bar;
  assign n19bar = in[3];
  assign n19 = inbar[3];
  assign n18bar = in[2];
  assign n18 = inbar[2];
  assign n17bar = in_0;
  assign n17 = in_0bar;
  OR2_X1 U5 ( .A1(n16), .A2(n15), .ZN(out[4]) );
  AND2_X1 U5bar ( .A1(n16bar), .A2(n15bar), .ZN(outbar[4]) );
  AND2_X1 U6 ( .A1(in[3]), .A2(n20), .ZN(n15) );
  OR2_X1 U6bar ( .A1(inbar[3]), .A2(n20bar), .ZN(n15bar) );
  AND2_X1 U7 ( .A1(in_7), .A2(n19), .ZN(n16) );
  OR2_X1 U7bar ( .A1(in_7bar), .A2(n19bar), .ZN(n16bar) );
  OR2_X1 U8 ( .A1(n14), .A2(n13), .ZN(out[3]) );
  AND2_X1 U8bar ( .A1(n14bar), .A2(n13bar), .ZN(outbar[3]) );
  AND2_X1 U9 ( .A1(in[2]), .A2(n20), .ZN(n13) );
  OR2_X1 U9bar ( .A1(inbar[2]), .A2(n20bar), .ZN(n13bar) );
  AND2_X1 U10 ( .A1(in_7), .A2(n18), .ZN(n14) );
  OR2_X1 U10bar ( .A1(in_7bar), .A2(n18bar), .ZN(n14bar) );
  OR2_X1 U11 ( .A1(n12), .A2(n11), .ZN(out[1]) );
  AND2_X1 U11bar ( .A1(n12bar), .A2(n11bar), .ZN(outbar[1]) );
  AND2_X1 U12 ( .A1(in_0), .A2(n20), .ZN(n11) );
  OR2_X1 U12bar ( .A1(in_0bar), .A2(n20bar), .ZN(n11bar) );
  AND2_X1 U13 ( .A1(in_7), .A2(n17), .ZN(n12) );
  OR2_X1 U13bar ( .A1(in_7bar), .A2(n17bar), .ZN(n12bar) );
endmodule

module scale2_15 ( in, inbar, out, outbar );

  input wire [7:0] in;
  input wire [7:0] inbar;
//input_done

  output wire [7:0] out;
  output wire [7:0] outbar;
//output_done

  wire in_0;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_1;
  wire in_7;
  wire n11;
  wire n12;
  wire n13;
  wire n14;
  wire n15;
  wire n16;
  wire n17;
  wire n18;
  wire n19;
  wire n20;
  wire in_0bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_1bar;
  wire in_7bar;
  wire n11bar;
  wire n12bar;
  wire n13bar;
  wire n14bar;
  wire n15bar;
  wire n16bar;
  wire n17bar;
  wire n18bar;
  wire n19bar;
  wire n20bar;
//wire_done

  assign in_0 = in[0];
  assign out[7] = in_6;
  assign in_6  = in[6];
  assign out[6] = in_5;
  assign in_5  = in[5];
  assign out[5] = in_4;
  assign in_4  = in[4];
  assign out[2] = in_1;
  assign in_1  = in[1];
  assign out[0] = in_7;
  assign in_7  = in[7];
  assign in_0bar = inbar[0];
  assign outbar[7] = in_6bar;
  assign in_6bar = inbar[6];
  assign outbar[6] = in_5bar;
  assign in_5bar = inbar[5];
  assign outbar[5] = in_4bar;
  assign in_4bar = inbar[4];
  assign outbar[2] = in_1bar;
  assign in_1bar = inbar[1];
  assign outbar[0] = in_7bar;
  assign in_7bar = inbar[7];
//assign_done

  assign n20bar = in_7;
  assign n20 = in_7bar;
  assign n19bar = in[3];
  assign n19 = inbar[3];
  assign n18bar = in[2];
  assign n18 = inbar[2];
  assign n17bar = in_0;
  assign n17 = in_0bar;
  OR2_X1 U5 ( .A1(n16), .A2(n15), .ZN(out[4]) );
  AND2_X1 U5bar ( .A1(n16bar), .A2(n15bar), .ZN(outbar[4]) );
  AND2_X1 U6 ( .A1(in[3]), .A2(n20), .ZN(n15) );
  OR2_X1 U6bar ( .A1(inbar[3]), .A2(n20bar), .ZN(n15bar) );
  AND2_X1 U7 ( .A1(in_7), .A2(n19), .ZN(n16) );
  OR2_X1 U7bar ( .A1(in_7bar), .A2(n19bar), .ZN(n16bar) );
  OR2_X1 U8 ( .A1(n14), .A2(n13), .ZN(out[3]) );
  AND2_X1 U8bar ( .A1(n14bar), .A2(n13bar), .ZN(outbar[3]) );
  AND2_X1 U9 ( .A1(in[2]), .A2(n20), .ZN(n13) );
  OR2_X1 U9bar ( .A1(inbar[2]), .A2(n20bar), .ZN(n13bar) );
  AND2_X1 U10 ( .A1(in_7), .A2(n18), .ZN(n14) );
  OR2_X1 U10bar ( .A1(in_7bar), .A2(n18bar), .ZN(n14bar) );
  OR2_X1 U11 ( .A1(n12), .A2(n11), .ZN(out[1]) );
  AND2_X1 U11bar ( .A1(n12bar), .A2(n11bar), .ZN(outbar[1]) );
  AND2_X1 U12 ( .A1(in_0), .A2(n20), .ZN(n11) );
  OR2_X1 U12bar ( .A1(in_0bar), .A2(n20bar), .ZN(n11bar) );
  AND2_X1 U13 ( .A1(in_7), .A2(n17), .ZN(n12) );
  OR2_X1 U13bar ( .A1(in_7bar), .A2(n17bar), .ZN(n12bar) );
endmodule

module byteXor_14 ( a, abar, b, bbar, y, ybar );

  input wire [7:0] a;
  input wire [7:0] b;
  input wire [7:0] abar;
  input wire [7:0] bbar;
//input_done

  output wire [7:0] y;
  output wire [7:0] ybar;
//output_done

  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n33bar;
  wire n34bar;
  wire n35bar;
  wire n36bar;
  wire n37bar;
  wire n38bar;
  wire n39bar;
  wire n40bar;
  wire n41bar;
  wire n42bar;
  wire n43bar;
  wire n44bar;
  wire n45bar;
  wire n46bar;
  wire n47bar;
  wire n48bar;
  wire n49bar;
  wire n50bar;
  wire n51bar;
  wire n52bar;
  wire n53bar;
  wire n54bar;
  wire n55bar;
  wire n56bar;
  wire n57bar;
  wire n58bar;
  wire n59bar;
  wire n60bar;
  wire n61bar;
  wire n62bar;
  wire n63bar;
  wire n64bar;
//wire_done

 //assign_done

  assign n64bar = n47;
  assign n64 = n47bar;
  assign n63bar = a[7];
  assign n63 = abar[7];
  assign n62bar = n45;
  assign n62 = n45bar;
  assign n61bar = a[6];
  assign n61 = abar[6];
  assign n60bar = n43;
  assign n60 = n43bar;
  assign n59bar = a[5];
  assign n59 = abar[5];
  assign n58bar = n41;
  assign n58 = n41bar;
  assign n57bar = a[4];
  assign n57 = abar[4];
  assign n56bar = n39;
  assign n56 = n39bar;
  assign n55bar = a[3];
  assign n55 = abar[3];
  assign n54bar = n37;
  assign n54 = n37bar;
  assign n53bar = a[2];
  assign n53 = abar[2];
  assign n52bar = n35;
  assign n52 = n35bar;
  assign n51bar = a[1];
  assign n51 = abar[1];
  assign n50bar = n33;
  assign n50 = n33bar;
  assign n49bar = a[0];
  assign n49 = abar[0];
  OR2_X1 U17 ( .A1(n48), .A2(n64), .ZN(y[7]) );
  AND2_X1 U17bar ( .A1(n48bar), .A2(n64bar), .ZN(ybar[7]) );
  OR2_X1 U18 ( .A1(n63), .A2(b[7]), .ZN(n47) );
  AND2_X1 U18bar ( .A1(n63bar), .A2(bbar[7]), .ZN(n47bar) );
  AND2_X1 U19 ( .A1(b[7]), .A2(n63), .ZN(n48) );
  OR2_X1 U19bar ( .A1(bbar[7]), .A2(n63bar), .ZN(n48bar) );
  OR2_X1 U20 ( .A1(n46), .A2(n62), .ZN(y[6]) );
  AND2_X1 U20bar ( .A1(n46bar), .A2(n62bar), .ZN(ybar[6]) );
  OR2_X1 U21 ( .A1(n61), .A2(b[6]), .ZN(n45) );
  AND2_X1 U21bar ( .A1(n61bar), .A2(bbar[6]), .ZN(n45bar) );
  AND2_X1 U22 ( .A1(b[6]), .A2(n61), .ZN(n46) );
  OR2_X1 U22bar ( .A1(bbar[6]), .A2(n61bar), .ZN(n46bar) );
  OR2_X1 U23 ( .A1(n44), .A2(n60), .ZN(y[5]) );
  AND2_X1 U23bar ( .A1(n44bar), .A2(n60bar), .ZN(ybar[5]) );
  OR2_X1 U24 ( .A1(n59), .A2(b[5]), .ZN(n43) );
  AND2_X1 U24bar ( .A1(n59bar), .A2(bbar[5]), .ZN(n43bar) );
  AND2_X1 U25 ( .A1(b[5]), .A2(n59), .ZN(n44) );
  OR2_X1 U25bar ( .A1(bbar[5]), .A2(n59bar), .ZN(n44bar) );
  OR2_X1 U26 ( .A1(n42), .A2(n58), .ZN(y[4]) );
  AND2_X1 U26bar ( .A1(n42bar), .A2(n58bar), .ZN(ybar[4]) );
  OR2_X1 U27 ( .A1(n57), .A2(b[4]), .ZN(n41) );
  AND2_X1 U27bar ( .A1(n57bar), .A2(bbar[4]), .ZN(n41bar) );
  AND2_X1 U28 ( .A1(b[4]), .A2(n57), .ZN(n42) );
  OR2_X1 U28bar ( .A1(bbar[4]), .A2(n57bar), .ZN(n42bar) );
  OR2_X1 U29 ( .A1(n40), .A2(n56), .ZN(y[3]) );
  AND2_X1 U29bar ( .A1(n40bar), .A2(n56bar), .ZN(ybar[3]) );
  OR2_X1 U30 ( .A1(n55), .A2(b[3]), .ZN(n39) );
  AND2_X1 U30bar ( .A1(n55bar), .A2(bbar[3]), .ZN(n39bar) );
  AND2_X1 U31 ( .A1(b[3]), .A2(n55), .ZN(n40) );
  OR2_X1 U31bar ( .A1(bbar[3]), .A2(n55bar), .ZN(n40bar) );
  OR2_X1 U32 ( .A1(n38), .A2(n54), .ZN(y[2]) );
  AND2_X1 U32bar ( .A1(n38bar), .A2(n54bar), .ZN(ybar[2]) );
  OR2_X1 U33 ( .A1(n53), .A2(b[2]), .ZN(n37) );
  AND2_X1 U33bar ( .A1(n53bar), .A2(bbar[2]), .ZN(n37bar) );
  AND2_X1 U34 ( .A1(b[2]), .A2(n53), .ZN(n38) );
  OR2_X1 U34bar ( .A1(bbar[2]), .A2(n53bar), .ZN(n38bar) );
  OR2_X1 U35 ( .A1(n36), .A2(n52), .ZN(y[1]) );
  AND2_X1 U35bar ( .A1(n36bar), .A2(n52bar), .ZN(ybar[1]) );
  OR2_X1 U36 ( .A1(n51), .A2(b[1]), .ZN(n35) );
  AND2_X1 U36bar ( .A1(n51bar), .A2(bbar[1]), .ZN(n35bar) );
  AND2_X1 U37 ( .A1(b[1]), .A2(n51), .ZN(n36) );
  OR2_X1 U37bar ( .A1(bbar[1]), .A2(n51bar), .ZN(n36bar) );
  OR2_X1 U38 ( .A1(n34), .A2(n50), .ZN(y[0]) );
  AND2_X1 U38bar ( .A1(n34bar), .A2(n50bar), .ZN(ybar[0]) );
  OR2_X1 U39 ( .A1(n49), .A2(b[0]), .ZN(n33) );
  AND2_X1 U39bar ( .A1(n49bar), .A2(bbar[0]), .ZN(n33bar) );
  AND2_X1 U40 ( .A1(b[0]), .A2(n49), .ZN(n34) );
  OR2_X1 U40bar ( .A1(bbar[0]), .A2(n49bar), .ZN(n34bar) );
endmodule

module byteXor_15 ( a, abar, b, bbar, y, ybar );

  input wire [7:0] a;
  input wire [7:0] b;
  input wire [7:0] abar;
  input wire [7:0] bbar;
//input_done

  output wire [7:0] y;
  output wire [7:0] ybar;
//output_done

  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n33bar;
  wire n34bar;
  wire n35bar;
  wire n36bar;
  wire n37bar;
  wire n38bar;
  wire n39bar;
  wire n40bar;
  wire n41bar;
  wire n42bar;
  wire n43bar;
  wire n44bar;
  wire n45bar;
  wire n46bar;
  wire n47bar;
  wire n48bar;
  wire n49bar;
  wire n50bar;
  wire n51bar;
  wire n52bar;
  wire n53bar;
  wire n54bar;
  wire n55bar;
  wire n56bar;
  wire n57bar;
  wire n58bar;
  wire n59bar;
  wire n60bar;
  wire n61bar;
  wire n62bar;
  wire n63bar;
  wire n64bar;
//wire_done

 //assign_done

  assign n64bar = n47;
  assign n64 = n47bar;
  assign n63bar = a[7];
  assign n63 = abar[7];
  assign n62bar = n45;
  assign n62 = n45bar;
  assign n61bar = a[6];
  assign n61 = abar[6];
  assign n60bar = n43;
  assign n60 = n43bar;
  assign n59bar = a[5];
  assign n59 = abar[5];
  assign n58bar = n41;
  assign n58 = n41bar;
  assign n57bar = a[4];
  assign n57 = abar[4];
  assign n56bar = n39;
  assign n56 = n39bar;
  assign n55bar = a[3];
  assign n55 = abar[3];
  assign n54bar = n37;
  assign n54 = n37bar;
  assign n53bar = a[2];
  assign n53 = abar[2];
  assign n52bar = n35;
  assign n52 = n35bar;
  assign n51bar = a[1];
  assign n51 = abar[1];
  assign n50bar = n33;
  assign n50 = n33bar;
  assign n49bar = a[0];
  assign n49 = abar[0];
  OR2_X1 U17 ( .A1(n48), .A2(n64), .ZN(y[7]) );
  AND2_X1 U17bar ( .A1(n48bar), .A2(n64bar), .ZN(ybar[7]) );
  OR2_X1 U18 ( .A1(n63), .A2(b[7]), .ZN(n47) );
  AND2_X1 U18bar ( .A1(n63bar), .A2(bbar[7]), .ZN(n47bar) );
  AND2_X1 U19 ( .A1(b[7]), .A2(n63), .ZN(n48) );
  OR2_X1 U19bar ( .A1(bbar[7]), .A2(n63bar), .ZN(n48bar) );
  OR2_X1 U20 ( .A1(n46), .A2(n62), .ZN(y[6]) );
  AND2_X1 U20bar ( .A1(n46bar), .A2(n62bar), .ZN(ybar[6]) );
  OR2_X1 U21 ( .A1(n61), .A2(b[6]), .ZN(n45) );
  AND2_X1 U21bar ( .A1(n61bar), .A2(bbar[6]), .ZN(n45bar) );
  AND2_X1 U22 ( .A1(b[6]), .A2(n61), .ZN(n46) );
  OR2_X1 U22bar ( .A1(bbar[6]), .A2(n61bar), .ZN(n46bar) );
  OR2_X1 U23 ( .A1(n44), .A2(n60), .ZN(y[5]) );
  AND2_X1 U23bar ( .A1(n44bar), .A2(n60bar), .ZN(ybar[5]) );
  OR2_X1 U24 ( .A1(n59), .A2(b[5]), .ZN(n43) );
  AND2_X1 U24bar ( .A1(n59bar), .A2(bbar[5]), .ZN(n43bar) );
  AND2_X1 U25 ( .A1(b[5]), .A2(n59), .ZN(n44) );
  OR2_X1 U25bar ( .A1(bbar[5]), .A2(n59bar), .ZN(n44bar) );
  OR2_X1 U26 ( .A1(n42), .A2(n58), .ZN(y[4]) );
  AND2_X1 U26bar ( .A1(n42bar), .A2(n58bar), .ZN(ybar[4]) );
  OR2_X1 U27 ( .A1(n57), .A2(b[4]), .ZN(n41) );
  AND2_X1 U27bar ( .A1(n57bar), .A2(bbar[4]), .ZN(n41bar) );
  AND2_X1 U28 ( .A1(b[4]), .A2(n57), .ZN(n42) );
  OR2_X1 U28bar ( .A1(bbar[4]), .A2(n57bar), .ZN(n42bar) );
  OR2_X1 U29 ( .A1(n40), .A2(n56), .ZN(y[3]) );
  AND2_X1 U29bar ( .A1(n40bar), .A2(n56bar), .ZN(ybar[3]) );
  OR2_X1 U30 ( .A1(n55), .A2(b[3]), .ZN(n39) );
  AND2_X1 U30bar ( .A1(n55bar), .A2(bbar[3]), .ZN(n39bar) );
  AND2_X1 U31 ( .A1(b[3]), .A2(n55), .ZN(n40) );
  OR2_X1 U31bar ( .A1(bbar[3]), .A2(n55bar), .ZN(n40bar) );
  OR2_X1 U32 ( .A1(n38), .A2(n54), .ZN(y[2]) );
  AND2_X1 U32bar ( .A1(n38bar), .A2(n54bar), .ZN(ybar[2]) );
  OR2_X1 U33 ( .A1(n53), .A2(b[2]), .ZN(n37) );
  AND2_X1 U33bar ( .A1(n53bar), .A2(bbar[2]), .ZN(n37bar) );
  AND2_X1 U34 ( .A1(b[2]), .A2(n53), .ZN(n38) );
  OR2_X1 U34bar ( .A1(bbar[2]), .A2(n53bar), .ZN(n38bar) );
  OR2_X1 U35 ( .A1(n36), .A2(n52), .ZN(y[1]) );
  AND2_X1 U35bar ( .A1(n36bar), .A2(n52bar), .ZN(ybar[1]) );
  OR2_X1 U36 ( .A1(n51), .A2(b[1]), .ZN(n35) );
  AND2_X1 U36bar ( .A1(n51bar), .A2(bbar[1]), .ZN(n35bar) );
  AND2_X1 U37 ( .A1(b[1]), .A2(n51), .ZN(n36) );
  OR2_X1 U37bar ( .A1(bbar[1]), .A2(n51bar), .ZN(n36bar) );
  OR2_X1 U38 ( .A1(n34), .A2(n50), .ZN(y[0]) );
  AND2_X1 U38bar ( .A1(n34bar), .A2(n50bar), .ZN(ybar[0]) );
  OR2_X1 U39 ( .A1(n49), .A2(b[0]), .ZN(n33) );
  AND2_X1 U39bar ( .A1(n49bar), .A2(bbar[0]), .ZN(n33bar) );
  AND2_X1 U40 ( .A1(b[0]), .A2(n49), .ZN(n34) );
  OR2_X1 U40bar ( .A1(bbar[0]), .A2(n49bar), .ZN(n34bar) );
endmodule

module byteXor_16 ( a, abar, b, bbar, y, ybar );

  input wire [7:0] a;
  input wire [7:0] b;
  input wire [7:0] abar;
  input wire [7:0] bbar;
//input_done

  output wire [7:0] y;
  output wire [7:0] ybar;
//output_done

  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n33bar;
  wire n34bar;
  wire n35bar;
  wire n36bar;
  wire n37bar;
  wire n38bar;
  wire n39bar;
  wire n40bar;
  wire n41bar;
  wire n42bar;
  wire n43bar;
  wire n44bar;
  wire n45bar;
  wire n46bar;
  wire n47bar;
  wire n48bar;
  wire n49bar;
  wire n50bar;
  wire n51bar;
  wire n52bar;
  wire n53bar;
  wire n54bar;
  wire n55bar;
  wire n56bar;
  wire n57bar;
  wire n58bar;
  wire n59bar;
  wire n60bar;
  wire n61bar;
  wire n62bar;
  wire n63bar;
  wire n64bar;
//wire_done

 //assign_done

  assign n64bar = n47;
  assign n64 = n47bar;
  assign n63bar = a[7];
  assign n63 = abar[7];
  assign n62bar = n45;
  assign n62 = n45bar;
  assign n61bar = a[6];
  assign n61 = abar[6];
  assign n60bar = n43;
  assign n60 = n43bar;
  assign n59bar = a[5];
  assign n59 = abar[5];
  assign n58bar = n41;
  assign n58 = n41bar;
  assign n57bar = a[4];
  assign n57 = abar[4];
  assign n56bar = n39;
  assign n56 = n39bar;
  assign n55bar = a[3];
  assign n55 = abar[3];
  assign n54bar = n37;
  assign n54 = n37bar;
  assign n53bar = a[2];
  assign n53 = abar[2];
  assign n52bar = n35;
  assign n52 = n35bar;
  assign n51bar = a[1];
  assign n51 = abar[1];
  assign n50bar = n33;
  assign n50 = n33bar;
  assign n49bar = a[0];
  assign n49 = abar[0];
  OR2_X1 U17 ( .A1(n48), .A2(n64), .ZN(y[7]) );
  AND2_X1 U17bar ( .A1(n48bar), .A2(n64bar), .ZN(ybar[7]) );
  OR2_X1 U18 ( .A1(n63), .A2(b[7]), .ZN(n47) );
  AND2_X1 U18bar ( .A1(n63bar), .A2(bbar[7]), .ZN(n47bar) );
  AND2_X1 U19 ( .A1(b[7]), .A2(n63), .ZN(n48) );
  OR2_X1 U19bar ( .A1(bbar[7]), .A2(n63bar), .ZN(n48bar) );
  OR2_X1 U20 ( .A1(n46), .A2(n62), .ZN(y[6]) );
  AND2_X1 U20bar ( .A1(n46bar), .A2(n62bar), .ZN(ybar[6]) );
  OR2_X1 U21 ( .A1(n61), .A2(b[6]), .ZN(n45) );
  AND2_X1 U21bar ( .A1(n61bar), .A2(bbar[6]), .ZN(n45bar) );
  AND2_X1 U22 ( .A1(b[6]), .A2(n61), .ZN(n46) );
  OR2_X1 U22bar ( .A1(bbar[6]), .A2(n61bar), .ZN(n46bar) );
  OR2_X1 U23 ( .A1(n44), .A2(n60), .ZN(y[5]) );
  AND2_X1 U23bar ( .A1(n44bar), .A2(n60bar), .ZN(ybar[5]) );
  OR2_X1 U24 ( .A1(n59), .A2(b[5]), .ZN(n43) );
  AND2_X1 U24bar ( .A1(n59bar), .A2(bbar[5]), .ZN(n43bar) );
  AND2_X1 U25 ( .A1(b[5]), .A2(n59), .ZN(n44) );
  OR2_X1 U25bar ( .A1(bbar[5]), .A2(n59bar), .ZN(n44bar) );
  OR2_X1 U26 ( .A1(n42), .A2(n58), .ZN(y[4]) );
  AND2_X1 U26bar ( .A1(n42bar), .A2(n58bar), .ZN(ybar[4]) );
  OR2_X1 U27 ( .A1(n57), .A2(b[4]), .ZN(n41) );
  AND2_X1 U27bar ( .A1(n57bar), .A2(bbar[4]), .ZN(n41bar) );
  AND2_X1 U28 ( .A1(b[4]), .A2(n57), .ZN(n42) );
  OR2_X1 U28bar ( .A1(bbar[4]), .A2(n57bar), .ZN(n42bar) );
  OR2_X1 U29 ( .A1(n40), .A2(n56), .ZN(y[3]) );
  AND2_X1 U29bar ( .A1(n40bar), .A2(n56bar), .ZN(ybar[3]) );
  OR2_X1 U30 ( .A1(n55), .A2(b[3]), .ZN(n39) );
  AND2_X1 U30bar ( .A1(n55bar), .A2(bbar[3]), .ZN(n39bar) );
  AND2_X1 U31 ( .A1(b[3]), .A2(n55), .ZN(n40) );
  OR2_X1 U31bar ( .A1(bbar[3]), .A2(n55bar), .ZN(n40bar) );
  OR2_X1 U32 ( .A1(n38), .A2(n54), .ZN(y[2]) );
  AND2_X1 U32bar ( .A1(n38bar), .A2(n54bar), .ZN(ybar[2]) );
  OR2_X1 U33 ( .A1(n53), .A2(b[2]), .ZN(n37) );
  AND2_X1 U33bar ( .A1(n53bar), .A2(bbar[2]), .ZN(n37bar) );
  AND2_X1 U34 ( .A1(b[2]), .A2(n53), .ZN(n38) );
  OR2_X1 U34bar ( .A1(bbar[2]), .A2(n53bar), .ZN(n38bar) );
  OR2_X1 U35 ( .A1(n36), .A2(n52), .ZN(y[1]) );
  AND2_X1 U35bar ( .A1(n36bar), .A2(n52bar), .ZN(ybar[1]) );
  OR2_X1 U36 ( .A1(n51), .A2(b[1]), .ZN(n35) );
  AND2_X1 U36bar ( .A1(n51bar), .A2(bbar[1]), .ZN(n35bar) );
  AND2_X1 U37 ( .A1(b[1]), .A2(n51), .ZN(n36) );
  OR2_X1 U37bar ( .A1(bbar[1]), .A2(n51bar), .ZN(n36bar) );
  OR2_X1 U38 ( .A1(n34), .A2(n50), .ZN(y[0]) );
  AND2_X1 U38bar ( .A1(n34bar), .A2(n50bar), .ZN(ybar[0]) );
  OR2_X1 U39 ( .A1(n49), .A2(b[0]), .ZN(n33) );
  AND2_X1 U39bar ( .A1(n49bar), .A2(bbar[0]), .ZN(n33bar) );
  AND2_X1 U40 ( .A1(b[0]), .A2(n49), .ZN(n34) );
  OR2_X1 U40bar ( .A1(bbar[0]), .A2(n49bar), .ZN(n34bar) );
endmodule

module byteXor4_13 ( a, abar, b, bbar, c, cbar, d, dbar, y, ybar );

  input wire [7:0] a;
  input wire [7:0] b;
  input wire [7:0] c;
  input wire [7:0] d;
  input wire [7:0] abar;
  input wire [7:0] bbar;
  input wire [7:0] cbar;
  input wire [7:0] dbar;
//input_done

  output wire [7:0] y;
  output wire [7:0] ybar;
//output_done

  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n113bar;
  wire n114bar;
  wire n115bar;
  wire n116bar;
  wire n117bar;
  wire n118bar;
  wire n119bar;
  wire n120bar;
  wire n121bar;
  wire n122bar;
  wire n123bar;
  wire n124bar;
  wire n125bar;
  wire n126bar;
  wire n127bar;
  wire n128bar;
  wire n129bar;
  wire n130bar;
  wire n131bar;
  wire n132bar;
  wire n133bar;
  wire n134bar;
  wire n135bar;
  wire n136bar;
  wire n137bar;
  wire n138bar;
  wire n139bar;
  wire n140bar;
  wire n141bar;
  wire n142bar;
  wire n143bar;
  wire n144bar;
  wire n145bar;
  wire n146bar;
  wire n147bar;
  wire n148bar;
  wire n149bar;
  wire n150bar;
  wire n151bar;
  wire n152bar;
  wire n153bar;
  wire n154bar;
  wire n155bar;
  wire n156bar;
  wire n157bar;
  wire n158bar;
  wire n159bar;
  wire n160bar;
  wire n161bar;
  wire n162bar;
  wire n163bar;
  wire n164bar;
  wire n165bar;
  wire n166bar;
  wire n167bar;
  wire n168bar;
  wire n169bar;
  wire n170bar;
  wire n171bar;
  wire n172bar;
  wire n173bar;
  wire n174bar;
  wire n175bar;
  wire n176bar;
  wire n177bar;
  wire n178bar;
  wire n179bar;
  wire n180bar;
  wire n181bar;
  wire n182bar;
  wire n183bar;
  wire n184bar;
  wire n185bar;
  wire n186bar;
  wire n187bar;
  wire n188bar;
  wire n189bar;
  wire n190bar;
  wire n191bar;
  wire n192bar;
  wire n193bar;
  wire n194bar;
  wire n195bar;
  wire n196bar;
  wire n197bar;
  wire n198bar;
  wire n199bar;
  wire n200bar;
  wire n201bar;
  wire n202bar;
  wire n203bar;
  wire n204bar;
  wire n205bar;
  wire n206bar;
  wire n207bar;
  wire n208bar;
  wire n209bar;
  wire n210bar;
  wire n211bar;
  wire n212bar;
  wire n213bar;
  wire n214bar;
  wire n215bar;
  wire n216bar;
  wire n217bar;
  wire n218bar;
  wire n219bar;
  wire n220bar;
  wire n221bar;
  wire n222bar;
  wire n223bar;
  wire n224bar;
//wire_done

 //assign_done

  assign n224bar = n175;
  assign n224 = n175bar;
  assign n223bar = a[7];
  assign n223 = abar[7];
  assign n222bar = n167;
  assign n222 = n167bar;
  assign n221bar = a[6];
  assign n221 = abar[6];
  assign n220bar = n159;
  assign n220 = n159bar;
  assign n219bar = a[5];
  assign n219 = abar[5];
  assign n218bar = n151;
  assign n218 = n151bar;
  assign n217bar = a[4];
  assign n217 = abar[4];
  assign n216bar = n143;
  assign n216 = n143bar;
  assign n215bar = a[3];
  assign n215 = abar[3];
  assign n214bar = n135;
  assign n214 = n135bar;
  assign n213bar = a[2];
  assign n213 = abar[2];
  assign n212bar = n127;
  assign n212 = n127bar;
  assign n211bar = a[1];
  assign n211 = abar[1];
  assign n210bar = n119;
  assign n210 = n119bar;
  assign n209bar = a[0];
  assign n209 = abar[0];
  assign n208bar = b[7];
  assign n208 = bbar[7];
  assign n207bar = b[6];
  assign n207 = bbar[6];
  assign n206bar = b[5];
  assign n206 = bbar[5];
  assign n205bar = b[4];
  assign n205 = bbar[4];
  assign n204bar = b[3];
  assign n204 = bbar[3];
  assign n203bar = b[2];
  assign n203 = bbar[2];
  assign n202bar = b[1];
  assign n202 = bbar[1];
  assign n201bar = b[0];
  assign n201 = bbar[0];
  assign n200bar = n171;
  assign n200 = n171bar;
  assign n199bar = c[7];
  assign n199 = cbar[7];
  assign n198bar = n163;
  assign n198 = n163bar;
  assign n197bar = c[6];
  assign n197 = cbar[6];
  assign n196bar = n155;
  assign n196 = n155bar;
  assign n195bar = c[5];
  assign n195 = cbar[5];
  assign n194bar = n147;
  assign n194 = n147bar;
  assign n193bar = c[4];
  assign n193 = cbar[4];
  assign n192bar = n139;
  assign n192 = n139bar;
  assign n191bar = c[3];
  assign n191 = cbar[3];
  assign n190bar = n131;
  assign n190 = n131bar;
  assign n189bar = c[2];
  assign n189 = cbar[2];
  assign n188bar = n123;
  assign n188 = n123bar;
  assign n187bar = c[1];
  assign n187 = cbar[1];
  assign n186bar = n115;
  assign n186 = n115bar;
  assign n185bar = c[0];
  assign n185 = cbar[0];
  assign n184bar = d[7];
  assign n184 = dbar[7];
  assign n183bar = d[6];
  assign n183 = dbar[6];
  assign n182bar = d[5];
  assign n182 = dbar[5];
  assign n181bar = d[4];
  assign n181 = dbar[4];
  assign n180bar = d[3];
  assign n180 = dbar[3];
  assign n179bar = d[2];
  assign n179 = dbar[2];
  assign n178bar = d[1];
  assign n178 = dbar[1];
  assign n177bar = d[0];
  assign n177 = dbar[0];
  OR2_X1 U49 ( .A1(n176), .A2(n224), .ZN(y[7]) );
  AND2_X1 U49bar ( .A1(n176bar), .A2(n224bar), .ZN(ybar[7]) );
  OR2_X1 U50 ( .A1(n174), .A2(n200), .ZN(n175) );
  AND2_X1 U50bar ( .A1(n174bar), .A2(n200bar), .ZN(n175bar) );
  AND2_X1 U51 ( .A1(n200), .A2(n174), .ZN(n176) );
  OR2_X1 U51bar ( .A1(n200bar), .A2(n174bar), .ZN(n176bar) );
  AND2_X1 U52 ( .A1(n173), .A2(n172), .ZN(n174) );
  OR2_X1 U52bar ( .A1(n173bar), .A2(n172bar), .ZN(n174bar) );
  OR2_X1 U53 ( .A1(n223), .A2(b[7]), .ZN(n172) );
  AND2_X1 U53bar ( .A1(n223bar), .A2(bbar[7]), .ZN(n172bar) );
  OR2_X1 U54 ( .A1(n208), .A2(a[7]), .ZN(n173) );
  AND2_X1 U54bar ( .A1(n208bar), .A2(abar[7]), .ZN(n173bar) );
  AND2_X1 U55 ( .A1(n170), .A2(n169), .ZN(n171) );
  OR2_X1 U55bar ( .A1(n170bar), .A2(n169bar), .ZN(n171bar) );
  OR2_X1 U56 ( .A1(n199), .A2(d[7]), .ZN(n169) );
  AND2_X1 U56bar ( .A1(n199bar), .A2(dbar[7]), .ZN(n169bar) );
  OR2_X1 U57 ( .A1(n184), .A2(c[7]), .ZN(n170) );
  AND2_X1 U57bar ( .A1(n184bar), .A2(cbar[7]), .ZN(n170bar) );
  OR2_X1 U58 ( .A1(n168), .A2(n222), .ZN(y[6]) );
  AND2_X1 U58bar ( .A1(n168bar), .A2(n222bar), .ZN(ybar[6]) );
  OR2_X1 U59 ( .A1(n166), .A2(n198), .ZN(n167) );
  AND2_X1 U59bar ( .A1(n166bar), .A2(n198bar), .ZN(n167bar) );
  AND2_X1 U60 ( .A1(n198), .A2(n166), .ZN(n168) );
  OR2_X1 U60bar ( .A1(n198bar), .A2(n166bar), .ZN(n168bar) );
  AND2_X1 U61 ( .A1(n165), .A2(n164), .ZN(n166) );
  OR2_X1 U61bar ( .A1(n165bar), .A2(n164bar), .ZN(n166bar) );
  OR2_X1 U62 ( .A1(n221), .A2(b[6]), .ZN(n164) );
  AND2_X1 U62bar ( .A1(n221bar), .A2(bbar[6]), .ZN(n164bar) );
  OR2_X1 U63 ( .A1(n207), .A2(a[6]), .ZN(n165) );
  AND2_X1 U63bar ( .A1(n207bar), .A2(abar[6]), .ZN(n165bar) );
  AND2_X1 U64 ( .A1(n162), .A2(n161), .ZN(n163) );
  OR2_X1 U64bar ( .A1(n162bar), .A2(n161bar), .ZN(n163bar) );
  OR2_X1 U65 ( .A1(n197), .A2(d[6]), .ZN(n161) );
  AND2_X1 U65bar ( .A1(n197bar), .A2(dbar[6]), .ZN(n161bar) );
  OR2_X1 U66 ( .A1(n183), .A2(c[6]), .ZN(n162) );
  AND2_X1 U66bar ( .A1(n183bar), .A2(cbar[6]), .ZN(n162bar) );
  OR2_X1 U67 ( .A1(n160), .A2(n220), .ZN(y[5]) );
  AND2_X1 U67bar ( .A1(n160bar), .A2(n220bar), .ZN(ybar[5]) );
  OR2_X1 U68 ( .A1(n158), .A2(n196), .ZN(n159) );
  AND2_X1 U68bar ( .A1(n158bar), .A2(n196bar), .ZN(n159bar) );
  AND2_X1 U69 ( .A1(n196), .A2(n158), .ZN(n160) );
  OR2_X1 U69bar ( .A1(n196bar), .A2(n158bar), .ZN(n160bar) );
  AND2_X1 U70 ( .A1(n157), .A2(n156), .ZN(n158) );
  OR2_X1 U70bar ( .A1(n157bar), .A2(n156bar), .ZN(n158bar) );
  OR2_X1 U71 ( .A1(n219), .A2(b[5]), .ZN(n156) );
  AND2_X1 U71bar ( .A1(n219bar), .A2(bbar[5]), .ZN(n156bar) );
  OR2_X1 U72 ( .A1(n206), .A2(a[5]), .ZN(n157) );
  AND2_X1 U72bar ( .A1(n206bar), .A2(abar[5]), .ZN(n157bar) );
  AND2_X1 U73 ( .A1(n154), .A2(n153), .ZN(n155) );
  OR2_X1 U73bar ( .A1(n154bar), .A2(n153bar), .ZN(n155bar) );
  OR2_X1 U74 ( .A1(n195), .A2(d[5]), .ZN(n153) );
  AND2_X1 U74bar ( .A1(n195bar), .A2(dbar[5]), .ZN(n153bar) );
  OR2_X1 U75 ( .A1(n182), .A2(c[5]), .ZN(n154) );
  AND2_X1 U75bar ( .A1(n182bar), .A2(cbar[5]), .ZN(n154bar) );
  OR2_X1 U76 ( .A1(n152), .A2(n218), .ZN(y[4]) );
  AND2_X1 U76bar ( .A1(n152bar), .A2(n218bar), .ZN(ybar[4]) );
  OR2_X1 U77 ( .A1(n150), .A2(n194), .ZN(n151) );
  AND2_X1 U77bar ( .A1(n150bar), .A2(n194bar), .ZN(n151bar) );
  AND2_X1 U78 ( .A1(n194), .A2(n150), .ZN(n152) );
  OR2_X1 U78bar ( .A1(n194bar), .A2(n150bar), .ZN(n152bar) );
  AND2_X1 U79 ( .A1(n149), .A2(n148), .ZN(n150) );
  OR2_X1 U79bar ( .A1(n149bar), .A2(n148bar), .ZN(n150bar) );
  OR2_X1 U80 ( .A1(n217), .A2(b[4]), .ZN(n148) );
  AND2_X1 U80bar ( .A1(n217bar), .A2(bbar[4]), .ZN(n148bar) );
  OR2_X1 U81 ( .A1(n205), .A2(a[4]), .ZN(n149) );
  AND2_X1 U81bar ( .A1(n205bar), .A2(abar[4]), .ZN(n149bar) );
  AND2_X1 U82 ( .A1(n146), .A2(n145), .ZN(n147) );
  OR2_X1 U82bar ( .A1(n146bar), .A2(n145bar), .ZN(n147bar) );
  OR2_X1 U83 ( .A1(n193), .A2(d[4]), .ZN(n145) );
  AND2_X1 U83bar ( .A1(n193bar), .A2(dbar[4]), .ZN(n145bar) );
  OR2_X1 U84 ( .A1(n181), .A2(c[4]), .ZN(n146) );
  AND2_X1 U84bar ( .A1(n181bar), .A2(cbar[4]), .ZN(n146bar) );
  OR2_X1 U85 ( .A1(n144), .A2(n216), .ZN(y[3]) );
  AND2_X1 U85bar ( .A1(n144bar), .A2(n216bar), .ZN(ybar[3]) );
  OR2_X1 U86 ( .A1(n142), .A2(n192), .ZN(n143) );
  AND2_X1 U86bar ( .A1(n142bar), .A2(n192bar), .ZN(n143bar) );
  AND2_X1 U87 ( .A1(n192), .A2(n142), .ZN(n144) );
  OR2_X1 U87bar ( .A1(n192bar), .A2(n142bar), .ZN(n144bar) );
  AND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(n142) );
  OR2_X1 U88bar ( .A1(n141bar), .A2(n140bar), .ZN(n142bar) );
  OR2_X1 U89 ( .A1(n215), .A2(b[3]), .ZN(n140) );
  AND2_X1 U89bar ( .A1(n215bar), .A2(bbar[3]), .ZN(n140bar) );
  OR2_X1 U90 ( .A1(n204), .A2(a[3]), .ZN(n141) );
  AND2_X1 U90bar ( .A1(n204bar), .A2(abar[3]), .ZN(n141bar) );
  AND2_X1 U91 ( .A1(n138), .A2(n137), .ZN(n139) );
  OR2_X1 U91bar ( .A1(n138bar), .A2(n137bar), .ZN(n139bar) );
  OR2_X1 U92 ( .A1(n191), .A2(d[3]), .ZN(n137) );
  AND2_X1 U92bar ( .A1(n191bar), .A2(dbar[3]), .ZN(n137bar) );
  OR2_X1 U93 ( .A1(n180), .A2(c[3]), .ZN(n138) );
  AND2_X1 U93bar ( .A1(n180bar), .A2(cbar[3]), .ZN(n138bar) );
  OR2_X1 U94 ( .A1(n136), .A2(n214), .ZN(y[2]) );
  AND2_X1 U94bar ( .A1(n136bar), .A2(n214bar), .ZN(ybar[2]) );
  OR2_X1 U95 ( .A1(n134), .A2(n190), .ZN(n135) );
  AND2_X1 U95bar ( .A1(n134bar), .A2(n190bar), .ZN(n135bar) );
  AND2_X1 U96 ( .A1(n190), .A2(n134), .ZN(n136) );
  OR2_X1 U96bar ( .A1(n190bar), .A2(n134bar), .ZN(n136bar) );
  AND2_X1 U97 ( .A1(n133), .A2(n132), .ZN(n134) );
  OR2_X1 U97bar ( .A1(n133bar), .A2(n132bar), .ZN(n134bar) );
  OR2_X1 U98 ( .A1(n213), .A2(b[2]), .ZN(n132) );
  AND2_X1 U98bar ( .A1(n213bar), .A2(bbar[2]), .ZN(n132bar) );
  OR2_X1 U99 ( .A1(n203), .A2(a[2]), .ZN(n133) );
  AND2_X1 U99bar ( .A1(n203bar), .A2(abar[2]), .ZN(n133bar) );
  AND2_X1 U100 ( .A1(n130), .A2(n129), .ZN(n131) );
  OR2_X1 U100bar ( .A1(n130bar), .A2(n129bar), .ZN(n131bar) );
  OR2_X1 U101 ( .A1(n189), .A2(d[2]), .ZN(n129) );
  AND2_X1 U101bar ( .A1(n189bar), .A2(dbar[2]), .ZN(n129bar) );
  OR2_X1 U102 ( .A1(n179), .A2(c[2]), .ZN(n130) );
  AND2_X1 U102bar ( .A1(n179bar), .A2(cbar[2]), .ZN(n130bar) );
  OR2_X1 U103 ( .A1(n128), .A2(n212), .ZN(y[1]) );
  AND2_X1 U103bar ( .A1(n128bar), .A2(n212bar), .ZN(ybar[1]) );
  OR2_X1 U104 ( .A1(n126), .A2(n188), .ZN(n127) );
  AND2_X1 U104bar ( .A1(n126bar), .A2(n188bar), .ZN(n127bar) );
  AND2_X1 U105 ( .A1(n188), .A2(n126), .ZN(n128) );
  OR2_X1 U105bar ( .A1(n188bar), .A2(n126bar), .ZN(n128bar) );
  AND2_X1 U106 ( .A1(n125), .A2(n124), .ZN(n126) );
  OR2_X1 U106bar ( .A1(n125bar), .A2(n124bar), .ZN(n126bar) );
  OR2_X1 U107 ( .A1(n211), .A2(b[1]), .ZN(n124) );
  AND2_X1 U107bar ( .A1(n211bar), .A2(bbar[1]), .ZN(n124bar) );
  OR2_X1 U108 ( .A1(n202), .A2(a[1]), .ZN(n125) );
  AND2_X1 U108bar ( .A1(n202bar), .A2(abar[1]), .ZN(n125bar) );
  AND2_X1 U109 ( .A1(n122), .A2(n121), .ZN(n123) );
  OR2_X1 U109bar ( .A1(n122bar), .A2(n121bar), .ZN(n123bar) );
  OR2_X1 U110 ( .A1(n187), .A2(d[1]), .ZN(n121) );
  AND2_X1 U110bar ( .A1(n187bar), .A2(dbar[1]), .ZN(n121bar) );
  OR2_X1 U111 ( .A1(n178), .A2(c[1]), .ZN(n122) );
  AND2_X1 U111bar ( .A1(n178bar), .A2(cbar[1]), .ZN(n122bar) );
  OR2_X1 U112 ( .A1(n120), .A2(n210), .ZN(y[0]) );
  AND2_X1 U112bar ( .A1(n120bar), .A2(n210bar), .ZN(ybar[0]) );
  OR2_X1 U113 ( .A1(n118), .A2(n186), .ZN(n119) );
  AND2_X1 U113bar ( .A1(n118bar), .A2(n186bar), .ZN(n119bar) );
  AND2_X1 U114 ( .A1(n186), .A2(n118), .ZN(n120) );
  OR2_X1 U114bar ( .A1(n186bar), .A2(n118bar), .ZN(n120bar) );
  AND2_X1 U115 ( .A1(n117), .A2(n116), .ZN(n118) );
  OR2_X1 U115bar ( .A1(n117bar), .A2(n116bar), .ZN(n118bar) );
  OR2_X1 U116 ( .A1(n209), .A2(b[0]), .ZN(n116) );
  AND2_X1 U116bar ( .A1(n209bar), .A2(bbar[0]), .ZN(n116bar) );
  OR2_X1 U117 ( .A1(n201), .A2(a[0]), .ZN(n117) );
  AND2_X1 U117bar ( .A1(n201bar), .A2(abar[0]), .ZN(n117bar) );
  AND2_X1 U118 ( .A1(n114), .A2(n113), .ZN(n115) );
  OR2_X1 U118bar ( .A1(n114bar), .A2(n113bar), .ZN(n115bar) );
  OR2_X1 U119 ( .A1(n185), .A2(d[0]), .ZN(n113) );
  AND2_X1 U119bar ( .A1(n185bar), .A2(dbar[0]), .ZN(n113bar) );
  OR2_X1 U120 ( .A1(n177), .A2(c[0]), .ZN(n114) );
  AND2_X1 U120bar ( .A1(n177bar), .A2(cbar[0]), .ZN(n114bar) );
endmodule

module byteXor4_14 ( a, abar, b, bbar, c, cbar, d, dbar, y, ybar );

  input wire [7:0] a;
  input wire [7:0] b;
  input wire [7:0] c;
  input wire [7:0] d;
  input wire [7:0] abar;
  input wire [7:0] bbar;
  input wire [7:0] cbar;
  input wire [7:0] dbar;
//input_done

  output wire [7:0] y;
  output wire [7:0] ybar;
//output_done

  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n113bar;
  wire n114bar;
  wire n115bar;
  wire n116bar;
  wire n117bar;
  wire n118bar;
  wire n119bar;
  wire n120bar;
  wire n121bar;
  wire n122bar;
  wire n123bar;
  wire n124bar;
  wire n125bar;
  wire n126bar;
  wire n127bar;
  wire n128bar;
  wire n129bar;
  wire n130bar;
  wire n131bar;
  wire n132bar;
  wire n133bar;
  wire n134bar;
  wire n135bar;
  wire n136bar;
  wire n137bar;
  wire n138bar;
  wire n139bar;
  wire n140bar;
  wire n141bar;
  wire n142bar;
  wire n143bar;
  wire n144bar;
  wire n145bar;
  wire n146bar;
  wire n147bar;
  wire n148bar;
  wire n149bar;
  wire n150bar;
  wire n151bar;
  wire n152bar;
  wire n153bar;
  wire n154bar;
  wire n155bar;
  wire n156bar;
  wire n157bar;
  wire n158bar;
  wire n159bar;
  wire n160bar;
  wire n161bar;
  wire n162bar;
  wire n163bar;
  wire n164bar;
  wire n165bar;
  wire n166bar;
  wire n167bar;
  wire n168bar;
  wire n169bar;
  wire n170bar;
  wire n171bar;
  wire n172bar;
  wire n173bar;
  wire n174bar;
  wire n175bar;
  wire n176bar;
  wire n177bar;
  wire n178bar;
  wire n179bar;
  wire n180bar;
  wire n181bar;
  wire n182bar;
  wire n183bar;
  wire n184bar;
  wire n185bar;
  wire n186bar;
  wire n187bar;
  wire n188bar;
  wire n189bar;
  wire n190bar;
  wire n191bar;
  wire n192bar;
  wire n193bar;
  wire n194bar;
  wire n195bar;
  wire n196bar;
  wire n197bar;
  wire n198bar;
  wire n199bar;
  wire n200bar;
  wire n201bar;
  wire n202bar;
  wire n203bar;
  wire n204bar;
  wire n205bar;
  wire n206bar;
  wire n207bar;
  wire n208bar;
  wire n209bar;
  wire n210bar;
  wire n211bar;
  wire n212bar;
  wire n213bar;
  wire n214bar;
  wire n215bar;
  wire n216bar;
  wire n217bar;
  wire n218bar;
  wire n219bar;
  wire n220bar;
  wire n221bar;
  wire n222bar;
  wire n223bar;
  wire n224bar;
//wire_done

 //assign_done

  assign n224bar = n175;
  assign n224 = n175bar;
  assign n223bar = a[7];
  assign n223 = abar[7];
  assign n222bar = n167;
  assign n222 = n167bar;
  assign n221bar = a[6];
  assign n221 = abar[6];
  assign n220bar = n159;
  assign n220 = n159bar;
  assign n219bar = a[5];
  assign n219 = abar[5];
  assign n218bar = n151;
  assign n218 = n151bar;
  assign n217bar = a[4];
  assign n217 = abar[4];
  assign n216bar = n143;
  assign n216 = n143bar;
  assign n215bar = a[3];
  assign n215 = abar[3];
  assign n214bar = n135;
  assign n214 = n135bar;
  assign n213bar = a[2];
  assign n213 = abar[2];
  assign n212bar = n127;
  assign n212 = n127bar;
  assign n211bar = a[1];
  assign n211 = abar[1];
  assign n210bar = n119;
  assign n210 = n119bar;
  assign n209bar = a[0];
  assign n209 = abar[0];
  assign n208bar = b[7];
  assign n208 = bbar[7];
  assign n207bar = b[6];
  assign n207 = bbar[6];
  assign n206bar = b[5];
  assign n206 = bbar[5];
  assign n205bar = b[4];
  assign n205 = bbar[4];
  assign n204bar = b[3];
  assign n204 = bbar[3];
  assign n203bar = b[2];
  assign n203 = bbar[2];
  assign n202bar = b[1];
  assign n202 = bbar[1];
  assign n201bar = b[0];
  assign n201 = bbar[0];
  assign n200bar = n171;
  assign n200 = n171bar;
  assign n199bar = c[7];
  assign n199 = cbar[7];
  assign n198bar = n163;
  assign n198 = n163bar;
  assign n197bar = c[6];
  assign n197 = cbar[6];
  assign n196bar = n155;
  assign n196 = n155bar;
  assign n195bar = c[5];
  assign n195 = cbar[5];
  assign n194bar = n147;
  assign n194 = n147bar;
  assign n193bar = c[4];
  assign n193 = cbar[4];
  assign n192bar = n139;
  assign n192 = n139bar;
  assign n191bar = c[3];
  assign n191 = cbar[3];
  assign n190bar = n131;
  assign n190 = n131bar;
  assign n189bar = c[2];
  assign n189 = cbar[2];
  assign n188bar = n123;
  assign n188 = n123bar;
  assign n187bar = c[1];
  assign n187 = cbar[1];
  assign n186bar = n115;
  assign n186 = n115bar;
  assign n185bar = c[0];
  assign n185 = cbar[0];
  assign n184bar = d[7];
  assign n184 = dbar[7];
  assign n183bar = d[6];
  assign n183 = dbar[6];
  assign n182bar = d[5];
  assign n182 = dbar[5];
  assign n181bar = d[4];
  assign n181 = dbar[4];
  assign n180bar = d[3];
  assign n180 = dbar[3];
  assign n179bar = d[2];
  assign n179 = dbar[2];
  assign n178bar = d[1];
  assign n178 = dbar[1];
  assign n177bar = d[0];
  assign n177 = dbar[0];
  OR2_X1 U49 ( .A1(n176), .A2(n224), .ZN(y[7]) );
  AND2_X1 U49bar ( .A1(n176bar), .A2(n224bar), .ZN(ybar[7]) );
  OR2_X1 U50 ( .A1(n174), .A2(n200), .ZN(n175) );
  AND2_X1 U50bar ( .A1(n174bar), .A2(n200bar), .ZN(n175bar) );
  AND2_X1 U51 ( .A1(n200), .A2(n174), .ZN(n176) );
  OR2_X1 U51bar ( .A1(n200bar), .A2(n174bar), .ZN(n176bar) );
  AND2_X1 U52 ( .A1(n173), .A2(n172), .ZN(n174) );
  OR2_X1 U52bar ( .A1(n173bar), .A2(n172bar), .ZN(n174bar) );
  OR2_X1 U53 ( .A1(n223), .A2(b[7]), .ZN(n172) );
  AND2_X1 U53bar ( .A1(n223bar), .A2(bbar[7]), .ZN(n172bar) );
  OR2_X1 U54 ( .A1(n208), .A2(a[7]), .ZN(n173) );
  AND2_X1 U54bar ( .A1(n208bar), .A2(abar[7]), .ZN(n173bar) );
  AND2_X1 U55 ( .A1(n170), .A2(n169), .ZN(n171) );
  OR2_X1 U55bar ( .A1(n170bar), .A2(n169bar), .ZN(n171bar) );
  OR2_X1 U56 ( .A1(n199), .A2(d[7]), .ZN(n169) );
  AND2_X1 U56bar ( .A1(n199bar), .A2(dbar[7]), .ZN(n169bar) );
  OR2_X1 U57 ( .A1(n184), .A2(c[7]), .ZN(n170) );
  AND2_X1 U57bar ( .A1(n184bar), .A2(cbar[7]), .ZN(n170bar) );
  OR2_X1 U58 ( .A1(n168), .A2(n222), .ZN(y[6]) );
  AND2_X1 U58bar ( .A1(n168bar), .A2(n222bar), .ZN(ybar[6]) );
  OR2_X1 U59 ( .A1(n166), .A2(n198), .ZN(n167) );
  AND2_X1 U59bar ( .A1(n166bar), .A2(n198bar), .ZN(n167bar) );
  AND2_X1 U60 ( .A1(n198), .A2(n166), .ZN(n168) );
  OR2_X1 U60bar ( .A1(n198bar), .A2(n166bar), .ZN(n168bar) );
  AND2_X1 U61 ( .A1(n165), .A2(n164), .ZN(n166) );
  OR2_X1 U61bar ( .A1(n165bar), .A2(n164bar), .ZN(n166bar) );
  OR2_X1 U62 ( .A1(n221), .A2(b[6]), .ZN(n164) );
  AND2_X1 U62bar ( .A1(n221bar), .A2(bbar[6]), .ZN(n164bar) );
  OR2_X1 U63 ( .A1(n207), .A2(a[6]), .ZN(n165) );
  AND2_X1 U63bar ( .A1(n207bar), .A2(abar[6]), .ZN(n165bar) );
  AND2_X1 U64 ( .A1(n162), .A2(n161), .ZN(n163) );
  OR2_X1 U64bar ( .A1(n162bar), .A2(n161bar), .ZN(n163bar) );
  OR2_X1 U65 ( .A1(n197), .A2(d[6]), .ZN(n161) );
  AND2_X1 U65bar ( .A1(n197bar), .A2(dbar[6]), .ZN(n161bar) );
  OR2_X1 U66 ( .A1(n183), .A2(c[6]), .ZN(n162) );
  AND2_X1 U66bar ( .A1(n183bar), .A2(cbar[6]), .ZN(n162bar) );
  OR2_X1 U67 ( .A1(n160), .A2(n220), .ZN(y[5]) );
  AND2_X1 U67bar ( .A1(n160bar), .A2(n220bar), .ZN(ybar[5]) );
  OR2_X1 U68 ( .A1(n158), .A2(n196), .ZN(n159) );
  AND2_X1 U68bar ( .A1(n158bar), .A2(n196bar), .ZN(n159bar) );
  AND2_X1 U69 ( .A1(n196), .A2(n158), .ZN(n160) );
  OR2_X1 U69bar ( .A1(n196bar), .A2(n158bar), .ZN(n160bar) );
  AND2_X1 U70 ( .A1(n157), .A2(n156), .ZN(n158) );
  OR2_X1 U70bar ( .A1(n157bar), .A2(n156bar), .ZN(n158bar) );
  OR2_X1 U71 ( .A1(n219), .A2(b[5]), .ZN(n156) );
  AND2_X1 U71bar ( .A1(n219bar), .A2(bbar[5]), .ZN(n156bar) );
  OR2_X1 U72 ( .A1(n206), .A2(a[5]), .ZN(n157) );
  AND2_X1 U72bar ( .A1(n206bar), .A2(abar[5]), .ZN(n157bar) );
  AND2_X1 U73 ( .A1(n154), .A2(n153), .ZN(n155) );
  OR2_X1 U73bar ( .A1(n154bar), .A2(n153bar), .ZN(n155bar) );
  OR2_X1 U74 ( .A1(n195), .A2(d[5]), .ZN(n153) );
  AND2_X1 U74bar ( .A1(n195bar), .A2(dbar[5]), .ZN(n153bar) );
  OR2_X1 U75 ( .A1(n182), .A2(c[5]), .ZN(n154) );
  AND2_X1 U75bar ( .A1(n182bar), .A2(cbar[5]), .ZN(n154bar) );
  OR2_X1 U76 ( .A1(n152), .A2(n218), .ZN(y[4]) );
  AND2_X1 U76bar ( .A1(n152bar), .A2(n218bar), .ZN(ybar[4]) );
  OR2_X1 U77 ( .A1(n150), .A2(n194), .ZN(n151) );
  AND2_X1 U77bar ( .A1(n150bar), .A2(n194bar), .ZN(n151bar) );
  AND2_X1 U78 ( .A1(n194), .A2(n150), .ZN(n152) );
  OR2_X1 U78bar ( .A1(n194bar), .A2(n150bar), .ZN(n152bar) );
  AND2_X1 U79 ( .A1(n149), .A2(n148), .ZN(n150) );
  OR2_X1 U79bar ( .A1(n149bar), .A2(n148bar), .ZN(n150bar) );
  OR2_X1 U80 ( .A1(n217), .A2(b[4]), .ZN(n148) );
  AND2_X1 U80bar ( .A1(n217bar), .A2(bbar[4]), .ZN(n148bar) );
  OR2_X1 U81 ( .A1(n205), .A2(a[4]), .ZN(n149) );
  AND2_X1 U81bar ( .A1(n205bar), .A2(abar[4]), .ZN(n149bar) );
  AND2_X1 U82 ( .A1(n146), .A2(n145), .ZN(n147) );
  OR2_X1 U82bar ( .A1(n146bar), .A2(n145bar), .ZN(n147bar) );
  OR2_X1 U83 ( .A1(n193), .A2(d[4]), .ZN(n145) );
  AND2_X1 U83bar ( .A1(n193bar), .A2(dbar[4]), .ZN(n145bar) );
  OR2_X1 U84 ( .A1(n181), .A2(c[4]), .ZN(n146) );
  AND2_X1 U84bar ( .A1(n181bar), .A2(cbar[4]), .ZN(n146bar) );
  OR2_X1 U85 ( .A1(n144), .A2(n216), .ZN(y[3]) );
  AND2_X1 U85bar ( .A1(n144bar), .A2(n216bar), .ZN(ybar[3]) );
  OR2_X1 U86 ( .A1(n142), .A2(n192), .ZN(n143) );
  AND2_X1 U86bar ( .A1(n142bar), .A2(n192bar), .ZN(n143bar) );
  AND2_X1 U87 ( .A1(n192), .A2(n142), .ZN(n144) );
  OR2_X1 U87bar ( .A1(n192bar), .A2(n142bar), .ZN(n144bar) );
  AND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(n142) );
  OR2_X1 U88bar ( .A1(n141bar), .A2(n140bar), .ZN(n142bar) );
  OR2_X1 U89 ( .A1(n215), .A2(b[3]), .ZN(n140) );
  AND2_X1 U89bar ( .A1(n215bar), .A2(bbar[3]), .ZN(n140bar) );
  OR2_X1 U90 ( .A1(n204), .A2(a[3]), .ZN(n141) );
  AND2_X1 U90bar ( .A1(n204bar), .A2(abar[3]), .ZN(n141bar) );
  AND2_X1 U91 ( .A1(n138), .A2(n137), .ZN(n139) );
  OR2_X1 U91bar ( .A1(n138bar), .A2(n137bar), .ZN(n139bar) );
  OR2_X1 U92 ( .A1(n191), .A2(d[3]), .ZN(n137) );
  AND2_X1 U92bar ( .A1(n191bar), .A2(dbar[3]), .ZN(n137bar) );
  OR2_X1 U93 ( .A1(n180), .A2(c[3]), .ZN(n138) );
  AND2_X1 U93bar ( .A1(n180bar), .A2(cbar[3]), .ZN(n138bar) );
  OR2_X1 U94 ( .A1(n136), .A2(n214), .ZN(y[2]) );
  AND2_X1 U94bar ( .A1(n136bar), .A2(n214bar), .ZN(ybar[2]) );
  OR2_X1 U95 ( .A1(n134), .A2(n190), .ZN(n135) );
  AND2_X1 U95bar ( .A1(n134bar), .A2(n190bar), .ZN(n135bar) );
  AND2_X1 U96 ( .A1(n190), .A2(n134), .ZN(n136) );
  OR2_X1 U96bar ( .A1(n190bar), .A2(n134bar), .ZN(n136bar) );
  AND2_X1 U97 ( .A1(n133), .A2(n132), .ZN(n134) );
  OR2_X1 U97bar ( .A1(n133bar), .A2(n132bar), .ZN(n134bar) );
  OR2_X1 U98 ( .A1(n213), .A2(b[2]), .ZN(n132) );
  AND2_X1 U98bar ( .A1(n213bar), .A2(bbar[2]), .ZN(n132bar) );
  OR2_X1 U99 ( .A1(n203), .A2(a[2]), .ZN(n133) );
  AND2_X1 U99bar ( .A1(n203bar), .A2(abar[2]), .ZN(n133bar) );
  AND2_X1 U100 ( .A1(n130), .A2(n129), .ZN(n131) );
  OR2_X1 U100bar ( .A1(n130bar), .A2(n129bar), .ZN(n131bar) );
  OR2_X1 U101 ( .A1(n189), .A2(d[2]), .ZN(n129) );
  AND2_X1 U101bar ( .A1(n189bar), .A2(dbar[2]), .ZN(n129bar) );
  OR2_X1 U102 ( .A1(n179), .A2(c[2]), .ZN(n130) );
  AND2_X1 U102bar ( .A1(n179bar), .A2(cbar[2]), .ZN(n130bar) );
  OR2_X1 U103 ( .A1(n128), .A2(n212), .ZN(y[1]) );
  AND2_X1 U103bar ( .A1(n128bar), .A2(n212bar), .ZN(ybar[1]) );
  OR2_X1 U104 ( .A1(n126), .A2(n188), .ZN(n127) );
  AND2_X1 U104bar ( .A1(n126bar), .A2(n188bar), .ZN(n127bar) );
  AND2_X1 U105 ( .A1(n188), .A2(n126), .ZN(n128) );
  OR2_X1 U105bar ( .A1(n188bar), .A2(n126bar), .ZN(n128bar) );
  AND2_X1 U106 ( .A1(n125), .A2(n124), .ZN(n126) );
  OR2_X1 U106bar ( .A1(n125bar), .A2(n124bar), .ZN(n126bar) );
  OR2_X1 U107 ( .A1(n211), .A2(b[1]), .ZN(n124) );
  AND2_X1 U107bar ( .A1(n211bar), .A2(bbar[1]), .ZN(n124bar) );
  OR2_X1 U108 ( .A1(n202), .A2(a[1]), .ZN(n125) );
  AND2_X1 U108bar ( .A1(n202bar), .A2(abar[1]), .ZN(n125bar) );
  AND2_X1 U109 ( .A1(n122), .A2(n121), .ZN(n123) );
  OR2_X1 U109bar ( .A1(n122bar), .A2(n121bar), .ZN(n123bar) );
  OR2_X1 U110 ( .A1(n187), .A2(d[1]), .ZN(n121) );
  AND2_X1 U110bar ( .A1(n187bar), .A2(dbar[1]), .ZN(n121bar) );
  OR2_X1 U111 ( .A1(n178), .A2(c[1]), .ZN(n122) );
  AND2_X1 U111bar ( .A1(n178bar), .A2(cbar[1]), .ZN(n122bar) );
  OR2_X1 U112 ( .A1(n120), .A2(n210), .ZN(y[0]) );
  AND2_X1 U112bar ( .A1(n120bar), .A2(n210bar), .ZN(ybar[0]) );
  OR2_X1 U113 ( .A1(n118), .A2(n186), .ZN(n119) );
  AND2_X1 U113bar ( .A1(n118bar), .A2(n186bar), .ZN(n119bar) );
  AND2_X1 U114 ( .A1(n186), .A2(n118), .ZN(n120) );
  OR2_X1 U114bar ( .A1(n186bar), .A2(n118bar), .ZN(n120bar) );
  AND2_X1 U115 ( .A1(n117), .A2(n116), .ZN(n118) );
  OR2_X1 U115bar ( .A1(n117bar), .A2(n116bar), .ZN(n118bar) );
  OR2_X1 U116 ( .A1(n209), .A2(b[0]), .ZN(n116) );
  AND2_X1 U116bar ( .A1(n209bar), .A2(bbar[0]), .ZN(n116bar) );
  OR2_X1 U117 ( .A1(n201), .A2(a[0]), .ZN(n117) );
  AND2_X1 U117bar ( .A1(n201bar), .A2(abar[0]), .ZN(n117bar) );
  AND2_X1 U118 ( .A1(n114), .A2(n113), .ZN(n115) );
  OR2_X1 U118bar ( .A1(n114bar), .A2(n113bar), .ZN(n115bar) );
  OR2_X1 U119 ( .A1(n185), .A2(d[0]), .ZN(n113) );
  AND2_X1 U119bar ( .A1(n185bar), .A2(dbar[0]), .ZN(n113bar) );
  OR2_X1 U120 ( .A1(n177), .A2(c[0]), .ZN(n114) );
  AND2_X1 U120bar ( .A1(n177bar), .A2(cbar[0]), .ZN(n114bar) );
endmodule

module byteXor4_15 ( a, abar, b, bbar, c, cbar, d, dbar, y, ybar );

  input wire [7:0] a;
  input wire [7:0] b;
  input wire [7:0] c;
  input wire [7:0] d;
  input wire [7:0] abar;
  input wire [7:0] bbar;
  input wire [7:0] cbar;
  input wire [7:0] dbar;
//input_done

  output wire [7:0] y;
  output wire [7:0] ybar;
//output_done

  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n113bar;
  wire n114bar;
  wire n115bar;
  wire n116bar;
  wire n117bar;
  wire n118bar;
  wire n119bar;
  wire n120bar;
  wire n121bar;
  wire n122bar;
  wire n123bar;
  wire n124bar;
  wire n125bar;
  wire n126bar;
  wire n127bar;
  wire n128bar;
  wire n129bar;
  wire n130bar;
  wire n131bar;
  wire n132bar;
  wire n133bar;
  wire n134bar;
  wire n135bar;
  wire n136bar;
  wire n137bar;
  wire n138bar;
  wire n139bar;
  wire n140bar;
  wire n141bar;
  wire n142bar;
  wire n143bar;
  wire n144bar;
  wire n145bar;
  wire n146bar;
  wire n147bar;
  wire n148bar;
  wire n149bar;
  wire n150bar;
  wire n151bar;
  wire n152bar;
  wire n153bar;
  wire n154bar;
  wire n155bar;
  wire n156bar;
  wire n157bar;
  wire n158bar;
  wire n159bar;
  wire n160bar;
  wire n161bar;
  wire n162bar;
  wire n163bar;
  wire n164bar;
  wire n165bar;
  wire n166bar;
  wire n167bar;
  wire n168bar;
  wire n169bar;
  wire n170bar;
  wire n171bar;
  wire n172bar;
  wire n173bar;
  wire n174bar;
  wire n175bar;
  wire n176bar;
  wire n177bar;
  wire n178bar;
  wire n179bar;
  wire n180bar;
  wire n181bar;
  wire n182bar;
  wire n183bar;
  wire n184bar;
  wire n185bar;
  wire n186bar;
  wire n187bar;
  wire n188bar;
  wire n189bar;
  wire n190bar;
  wire n191bar;
  wire n192bar;
  wire n193bar;
  wire n194bar;
  wire n195bar;
  wire n196bar;
  wire n197bar;
  wire n198bar;
  wire n199bar;
  wire n200bar;
  wire n201bar;
  wire n202bar;
  wire n203bar;
  wire n204bar;
  wire n205bar;
  wire n206bar;
  wire n207bar;
  wire n208bar;
  wire n209bar;
  wire n210bar;
  wire n211bar;
  wire n212bar;
  wire n213bar;
  wire n214bar;
  wire n215bar;
  wire n216bar;
  wire n217bar;
  wire n218bar;
  wire n219bar;
  wire n220bar;
  wire n221bar;
  wire n222bar;
  wire n223bar;
  wire n224bar;
//wire_done

 //assign_done

  assign n224bar = n175;
  assign n224 = n175bar;
  assign n223bar = a[7];
  assign n223 = abar[7];
  assign n222bar = n167;
  assign n222 = n167bar;
  assign n221bar = a[6];
  assign n221 = abar[6];
  assign n220bar = n159;
  assign n220 = n159bar;
  assign n219bar = a[5];
  assign n219 = abar[5];
  assign n218bar = n151;
  assign n218 = n151bar;
  assign n217bar = a[4];
  assign n217 = abar[4];
  assign n216bar = n143;
  assign n216 = n143bar;
  assign n215bar = a[3];
  assign n215 = abar[3];
  assign n214bar = n135;
  assign n214 = n135bar;
  assign n213bar = a[2];
  assign n213 = abar[2];
  assign n212bar = n127;
  assign n212 = n127bar;
  assign n211bar = a[1];
  assign n211 = abar[1];
  assign n210bar = n119;
  assign n210 = n119bar;
  assign n209bar = a[0];
  assign n209 = abar[0];
  assign n208bar = b[7];
  assign n208 = bbar[7];
  assign n207bar = b[6];
  assign n207 = bbar[6];
  assign n206bar = b[5];
  assign n206 = bbar[5];
  assign n205bar = b[4];
  assign n205 = bbar[4];
  assign n204bar = b[3];
  assign n204 = bbar[3];
  assign n203bar = b[2];
  assign n203 = bbar[2];
  assign n202bar = b[1];
  assign n202 = bbar[1];
  assign n201bar = b[0];
  assign n201 = bbar[0];
  assign n200bar = n171;
  assign n200 = n171bar;
  assign n199bar = c[7];
  assign n199 = cbar[7];
  assign n198bar = n163;
  assign n198 = n163bar;
  assign n197bar = c[6];
  assign n197 = cbar[6];
  assign n196bar = n155;
  assign n196 = n155bar;
  assign n195bar = c[5];
  assign n195 = cbar[5];
  assign n194bar = n147;
  assign n194 = n147bar;
  assign n193bar = c[4];
  assign n193 = cbar[4];
  assign n192bar = n139;
  assign n192 = n139bar;
  assign n191bar = c[3];
  assign n191 = cbar[3];
  assign n190bar = n131;
  assign n190 = n131bar;
  assign n189bar = c[2];
  assign n189 = cbar[2];
  assign n188bar = n123;
  assign n188 = n123bar;
  assign n187bar = c[1];
  assign n187 = cbar[1];
  assign n186bar = n115;
  assign n186 = n115bar;
  assign n185bar = c[0];
  assign n185 = cbar[0];
  assign n184bar = d[7];
  assign n184 = dbar[7];
  assign n183bar = d[6];
  assign n183 = dbar[6];
  assign n182bar = d[5];
  assign n182 = dbar[5];
  assign n181bar = d[4];
  assign n181 = dbar[4];
  assign n180bar = d[3];
  assign n180 = dbar[3];
  assign n179bar = d[2];
  assign n179 = dbar[2];
  assign n178bar = d[1];
  assign n178 = dbar[1];
  assign n177bar = d[0];
  assign n177 = dbar[0];
  OR2_X1 U49 ( .A1(n176), .A2(n224), .ZN(y[7]) );
  AND2_X1 U49bar ( .A1(n176bar), .A2(n224bar), .ZN(ybar[7]) );
  OR2_X1 U50 ( .A1(n174), .A2(n200), .ZN(n175) );
  AND2_X1 U50bar ( .A1(n174bar), .A2(n200bar), .ZN(n175bar) );
  AND2_X1 U51 ( .A1(n200), .A2(n174), .ZN(n176) );
  OR2_X1 U51bar ( .A1(n200bar), .A2(n174bar), .ZN(n176bar) );
  AND2_X1 U52 ( .A1(n173), .A2(n172), .ZN(n174) );
  OR2_X1 U52bar ( .A1(n173bar), .A2(n172bar), .ZN(n174bar) );
  OR2_X1 U53 ( .A1(n223), .A2(b[7]), .ZN(n172) );
  AND2_X1 U53bar ( .A1(n223bar), .A2(bbar[7]), .ZN(n172bar) );
  OR2_X1 U54 ( .A1(n208), .A2(a[7]), .ZN(n173) );
  AND2_X1 U54bar ( .A1(n208bar), .A2(abar[7]), .ZN(n173bar) );
  AND2_X1 U55 ( .A1(n170), .A2(n169), .ZN(n171) );
  OR2_X1 U55bar ( .A1(n170bar), .A2(n169bar), .ZN(n171bar) );
  OR2_X1 U56 ( .A1(n199), .A2(d[7]), .ZN(n169) );
  AND2_X1 U56bar ( .A1(n199bar), .A2(dbar[7]), .ZN(n169bar) );
  OR2_X1 U57 ( .A1(n184), .A2(c[7]), .ZN(n170) );
  AND2_X1 U57bar ( .A1(n184bar), .A2(cbar[7]), .ZN(n170bar) );
  OR2_X1 U58 ( .A1(n168), .A2(n222), .ZN(y[6]) );
  AND2_X1 U58bar ( .A1(n168bar), .A2(n222bar), .ZN(ybar[6]) );
  OR2_X1 U59 ( .A1(n166), .A2(n198), .ZN(n167) );
  AND2_X1 U59bar ( .A1(n166bar), .A2(n198bar), .ZN(n167bar) );
  AND2_X1 U60 ( .A1(n198), .A2(n166), .ZN(n168) );
  OR2_X1 U60bar ( .A1(n198bar), .A2(n166bar), .ZN(n168bar) );
  AND2_X1 U61 ( .A1(n165), .A2(n164), .ZN(n166) );
  OR2_X1 U61bar ( .A1(n165bar), .A2(n164bar), .ZN(n166bar) );
  OR2_X1 U62 ( .A1(n221), .A2(b[6]), .ZN(n164) );
  AND2_X1 U62bar ( .A1(n221bar), .A2(bbar[6]), .ZN(n164bar) );
  OR2_X1 U63 ( .A1(n207), .A2(a[6]), .ZN(n165) );
  AND2_X1 U63bar ( .A1(n207bar), .A2(abar[6]), .ZN(n165bar) );
  AND2_X1 U64 ( .A1(n162), .A2(n161), .ZN(n163) );
  OR2_X1 U64bar ( .A1(n162bar), .A2(n161bar), .ZN(n163bar) );
  OR2_X1 U65 ( .A1(n197), .A2(d[6]), .ZN(n161) );
  AND2_X1 U65bar ( .A1(n197bar), .A2(dbar[6]), .ZN(n161bar) );
  OR2_X1 U66 ( .A1(n183), .A2(c[6]), .ZN(n162) );
  AND2_X1 U66bar ( .A1(n183bar), .A2(cbar[6]), .ZN(n162bar) );
  OR2_X1 U67 ( .A1(n160), .A2(n220), .ZN(y[5]) );
  AND2_X1 U67bar ( .A1(n160bar), .A2(n220bar), .ZN(ybar[5]) );
  OR2_X1 U68 ( .A1(n158), .A2(n196), .ZN(n159) );
  AND2_X1 U68bar ( .A1(n158bar), .A2(n196bar), .ZN(n159bar) );
  AND2_X1 U69 ( .A1(n196), .A2(n158), .ZN(n160) );
  OR2_X1 U69bar ( .A1(n196bar), .A2(n158bar), .ZN(n160bar) );
  AND2_X1 U70 ( .A1(n157), .A2(n156), .ZN(n158) );
  OR2_X1 U70bar ( .A1(n157bar), .A2(n156bar), .ZN(n158bar) );
  OR2_X1 U71 ( .A1(n219), .A2(b[5]), .ZN(n156) );
  AND2_X1 U71bar ( .A1(n219bar), .A2(bbar[5]), .ZN(n156bar) );
  OR2_X1 U72 ( .A1(n206), .A2(a[5]), .ZN(n157) );
  AND2_X1 U72bar ( .A1(n206bar), .A2(abar[5]), .ZN(n157bar) );
  AND2_X1 U73 ( .A1(n154), .A2(n153), .ZN(n155) );
  OR2_X1 U73bar ( .A1(n154bar), .A2(n153bar), .ZN(n155bar) );
  OR2_X1 U74 ( .A1(n195), .A2(d[5]), .ZN(n153) );
  AND2_X1 U74bar ( .A1(n195bar), .A2(dbar[5]), .ZN(n153bar) );
  OR2_X1 U75 ( .A1(n182), .A2(c[5]), .ZN(n154) );
  AND2_X1 U75bar ( .A1(n182bar), .A2(cbar[5]), .ZN(n154bar) );
  OR2_X1 U76 ( .A1(n152), .A2(n218), .ZN(y[4]) );
  AND2_X1 U76bar ( .A1(n152bar), .A2(n218bar), .ZN(ybar[4]) );
  OR2_X1 U77 ( .A1(n150), .A2(n194), .ZN(n151) );
  AND2_X1 U77bar ( .A1(n150bar), .A2(n194bar), .ZN(n151bar) );
  AND2_X1 U78 ( .A1(n194), .A2(n150), .ZN(n152) );
  OR2_X1 U78bar ( .A1(n194bar), .A2(n150bar), .ZN(n152bar) );
  AND2_X1 U79 ( .A1(n149), .A2(n148), .ZN(n150) );
  OR2_X1 U79bar ( .A1(n149bar), .A2(n148bar), .ZN(n150bar) );
  OR2_X1 U80 ( .A1(n217), .A2(b[4]), .ZN(n148) );
  AND2_X1 U80bar ( .A1(n217bar), .A2(bbar[4]), .ZN(n148bar) );
  OR2_X1 U81 ( .A1(n205), .A2(a[4]), .ZN(n149) );
  AND2_X1 U81bar ( .A1(n205bar), .A2(abar[4]), .ZN(n149bar) );
  AND2_X1 U82 ( .A1(n146), .A2(n145), .ZN(n147) );
  OR2_X1 U82bar ( .A1(n146bar), .A2(n145bar), .ZN(n147bar) );
  OR2_X1 U83 ( .A1(n193), .A2(d[4]), .ZN(n145) );
  AND2_X1 U83bar ( .A1(n193bar), .A2(dbar[4]), .ZN(n145bar) );
  OR2_X1 U84 ( .A1(n181), .A2(c[4]), .ZN(n146) );
  AND2_X1 U84bar ( .A1(n181bar), .A2(cbar[4]), .ZN(n146bar) );
  OR2_X1 U85 ( .A1(n144), .A2(n216), .ZN(y[3]) );
  AND2_X1 U85bar ( .A1(n144bar), .A2(n216bar), .ZN(ybar[3]) );
  OR2_X1 U86 ( .A1(n142), .A2(n192), .ZN(n143) );
  AND2_X1 U86bar ( .A1(n142bar), .A2(n192bar), .ZN(n143bar) );
  AND2_X1 U87 ( .A1(n192), .A2(n142), .ZN(n144) );
  OR2_X1 U87bar ( .A1(n192bar), .A2(n142bar), .ZN(n144bar) );
  AND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(n142) );
  OR2_X1 U88bar ( .A1(n141bar), .A2(n140bar), .ZN(n142bar) );
  OR2_X1 U89 ( .A1(n215), .A2(b[3]), .ZN(n140) );
  AND2_X1 U89bar ( .A1(n215bar), .A2(bbar[3]), .ZN(n140bar) );
  OR2_X1 U90 ( .A1(n204), .A2(a[3]), .ZN(n141) );
  AND2_X1 U90bar ( .A1(n204bar), .A2(abar[3]), .ZN(n141bar) );
  AND2_X1 U91 ( .A1(n138), .A2(n137), .ZN(n139) );
  OR2_X1 U91bar ( .A1(n138bar), .A2(n137bar), .ZN(n139bar) );
  OR2_X1 U92 ( .A1(n191), .A2(d[3]), .ZN(n137) );
  AND2_X1 U92bar ( .A1(n191bar), .A2(dbar[3]), .ZN(n137bar) );
  OR2_X1 U93 ( .A1(n180), .A2(c[3]), .ZN(n138) );
  AND2_X1 U93bar ( .A1(n180bar), .A2(cbar[3]), .ZN(n138bar) );
  OR2_X1 U94 ( .A1(n136), .A2(n214), .ZN(y[2]) );
  AND2_X1 U94bar ( .A1(n136bar), .A2(n214bar), .ZN(ybar[2]) );
  OR2_X1 U95 ( .A1(n134), .A2(n190), .ZN(n135) );
  AND2_X1 U95bar ( .A1(n134bar), .A2(n190bar), .ZN(n135bar) );
  AND2_X1 U96 ( .A1(n190), .A2(n134), .ZN(n136) );
  OR2_X1 U96bar ( .A1(n190bar), .A2(n134bar), .ZN(n136bar) );
  AND2_X1 U97 ( .A1(n133), .A2(n132), .ZN(n134) );
  OR2_X1 U97bar ( .A1(n133bar), .A2(n132bar), .ZN(n134bar) );
  OR2_X1 U98 ( .A1(n213), .A2(b[2]), .ZN(n132) );
  AND2_X1 U98bar ( .A1(n213bar), .A2(bbar[2]), .ZN(n132bar) );
  OR2_X1 U99 ( .A1(n203), .A2(a[2]), .ZN(n133) );
  AND2_X1 U99bar ( .A1(n203bar), .A2(abar[2]), .ZN(n133bar) );
  AND2_X1 U100 ( .A1(n130), .A2(n129), .ZN(n131) );
  OR2_X1 U100bar ( .A1(n130bar), .A2(n129bar), .ZN(n131bar) );
  OR2_X1 U101 ( .A1(n189), .A2(d[2]), .ZN(n129) );
  AND2_X1 U101bar ( .A1(n189bar), .A2(dbar[2]), .ZN(n129bar) );
  OR2_X1 U102 ( .A1(n179), .A2(c[2]), .ZN(n130) );
  AND2_X1 U102bar ( .A1(n179bar), .A2(cbar[2]), .ZN(n130bar) );
  OR2_X1 U103 ( .A1(n128), .A2(n212), .ZN(y[1]) );
  AND2_X1 U103bar ( .A1(n128bar), .A2(n212bar), .ZN(ybar[1]) );
  OR2_X1 U104 ( .A1(n126), .A2(n188), .ZN(n127) );
  AND2_X1 U104bar ( .A1(n126bar), .A2(n188bar), .ZN(n127bar) );
  AND2_X1 U105 ( .A1(n188), .A2(n126), .ZN(n128) );
  OR2_X1 U105bar ( .A1(n188bar), .A2(n126bar), .ZN(n128bar) );
  AND2_X1 U106 ( .A1(n125), .A2(n124), .ZN(n126) );
  OR2_X1 U106bar ( .A1(n125bar), .A2(n124bar), .ZN(n126bar) );
  OR2_X1 U107 ( .A1(n211), .A2(b[1]), .ZN(n124) );
  AND2_X1 U107bar ( .A1(n211bar), .A2(bbar[1]), .ZN(n124bar) );
  OR2_X1 U108 ( .A1(n202), .A2(a[1]), .ZN(n125) );
  AND2_X1 U108bar ( .A1(n202bar), .A2(abar[1]), .ZN(n125bar) );
  AND2_X1 U109 ( .A1(n122), .A2(n121), .ZN(n123) );
  OR2_X1 U109bar ( .A1(n122bar), .A2(n121bar), .ZN(n123bar) );
  OR2_X1 U110 ( .A1(n187), .A2(d[1]), .ZN(n121) );
  AND2_X1 U110bar ( .A1(n187bar), .A2(dbar[1]), .ZN(n121bar) );
  OR2_X1 U111 ( .A1(n178), .A2(c[1]), .ZN(n122) );
  AND2_X1 U111bar ( .A1(n178bar), .A2(cbar[1]), .ZN(n122bar) );
  OR2_X1 U112 ( .A1(n120), .A2(n210), .ZN(y[0]) );
  AND2_X1 U112bar ( .A1(n120bar), .A2(n210bar), .ZN(ybar[0]) );
  OR2_X1 U113 ( .A1(n118), .A2(n186), .ZN(n119) );
  AND2_X1 U113bar ( .A1(n118bar), .A2(n186bar), .ZN(n119bar) );
  AND2_X1 U114 ( .A1(n186), .A2(n118), .ZN(n120) );
  OR2_X1 U114bar ( .A1(n186bar), .A2(n118bar), .ZN(n120bar) );
  AND2_X1 U115 ( .A1(n117), .A2(n116), .ZN(n118) );
  OR2_X1 U115bar ( .A1(n117bar), .A2(n116bar), .ZN(n118bar) );
  OR2_X1 U116 ( .A1(n209), .A2(b[0]), .ZN(n116) );
  AND2_X1 U116bar ( .A1(n209bar), .A2(bbar[0]), .ZN(n116bar) );
  OR2_X1 U117 ( .A1(n201), .A2(a[0]), .ZN(n117) );
  AND2_X1 U117bar ( .A1(n201bar), .A2(abar[0]), .ZN(n117bar) );
  AND2_X1 U118 ( .A1(n114), .A2(n113), .ZN(n115) );
  OR2_X1 U118bar ( .A1(n114bar), .A2(n113bar), .ZN(n115bar) );
  OR2_X1 U119 ( .A1(n185), .A2(d[0]), .ZN(n113) );
  AND2_X1 U119bar ( .A1(n185bar), .A2(dbar[0]), .ZN(n113bar) );
  OR2_X1 U120 ( .A1(n177), .A2(c[0]), .ZN(n114) );
  AND2_X1 U120bar ( .A1(n177bar), .A2(cbar[0]), .ZN(n114bar) );
endmodule

module mixCol_0 ( in, inbar, out, outbar );


  input wire [31:0] in;
  input wire [31:0] inbar;
//input_done

  output wire [31:0] out;
  output wire [31:0] outbar;
//output_done

  wire [7:0] b0_s2;
  wire [7:0] b1_s2;
  wire [7:0] b2_s2;
  wire [7:0] b3_s2;
  wire [7:0] b0_s3;
  wire [7:0] b1_s3;
  wire [7:0] b2_s3;
  wire [7:0] b3_s3;

  wire [7:0] b0_s2bar;
  wire [7:0] b1_s2bar;
  wire [7:0] b2_s2bar;
  wire [7:0] b3_s2bar;
  wire [7:0] b0_s3bar;
  wire [7:0] b1_s3bar;
  wire [7:0] b2_s3bar;
  wire [7:0] b3_s3bar;
//wire_done

 //assign_done

  scale2_0 b0_scale2 ( .in(in[31:24]), .inbar(inbar[31:24]), .out(b0_s2), .outbar(b0_s2bar) );
  scale2_15 b1_scale2 ( .in(in[23:16]), .inbar(inbar[23:16]), .out(b1_s2), .outbar(b1_s2bar) );
  scale2_14 b2_scale2 ( .in(in[15:8]), .inbar(inbar[15:8]), .out(b2_s2), .outbar(b2_s2bar) );
  scale2_13 b3_scale2 ( .in(in[7:0]), .inbar(inbar[7:0]), .out(b3_s2), .outbar(b3_s2bar) );

  byteXor_0 b0_scale3 ( .a(in[31:24]), .abar(inbar[31:24]), .b(b0_s2), .bbar(b0_s2bar), .y(b0_s3), .ybar(b0_s3bar) );
  byteXor_16 b1_scale3 ( .a(in[23:16]), .abar(inbar[23:16]), .b(b1_s2), .bbar(b1_s2bar), .y(b1_s3), .ybar(b1_s3bar) );
  byteXor_15 b2_scale3 ( .a(in[15:8]), .abar(inbar[15:8]), .b(b2_s2), .bbar(b2_s2bar), .y(b2_s3), .ybar(b2_s3bar) );
  byteXor_14 b3_scale3 ( .a(in[7:0]), .abar(inbar[7:0]), .b(b3_s2), .bbar(b3_s2bar), .y(b3_s3), .ybar(b3_s3bar) );

  byteXor4_0 out0 ( .a(b0_s2), .abar(b0_s2bar), .b(b1_s3), .bbar(b1_s3bar), .c(in[15:8]), .cbar(inbar[15:8]),
       .d(in[7:0]), .dbar(inbar[7:0]), .y(out[31:24]), .ybar(outbar[31:24]) );
  byteXor4_15 out1 ( .a(in[31:24]), .abar(inbar[31:24]), .b(b1_s2), .bbar(b1_s2bar), .c(b2_s3), .cbar(b2_s3bar),
       .d(in[7:0]), .dbar(inbar[7:0]), .y(out[23:16]), .ybar(outbar[23:16]) );
  byteXor4_14 out2 ( .a(in[31:24]), .abar(inbar[31:24]), .b(in[23:16]), .bbar(inbar[23:16]), .c(b2_s2), .cbar(b2_s2bar),
       .d(b3_s3), .dbar(b3_s3bar), .y(out[15:8]), .ybar(outbar[15:8]) );
  byteXor4_13 out3 ( .a(b0_s3), .abar(b0_s3bar), .b(in[23:16]), .bbar(inbar[23:16]), .c(in[15:8]), .cbar(inbar[15:8]),
       .d(b3_s2), .dbar(b3_s2bar), .y(out[7:0]), .ybar(outbar[7:0]) );
endmodule

module scale2_1 ( in, inbar, out, outbar );

  input wire [7:0] in;
  input wire [7:0] inbar;
//input_done

  output wire [7:0] out;
  output wire [7:0] outbar;
//output_done

  wire in_0;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_1;
  wire in_7;
  wire n11;
  wire n12;
  wire n13;
  wire n14;
  wire n15;
  wire n16;
  wire n17;
  wire n18;
  wire n19;
  wire n20;
  wire in_0bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_1bar;
  wire in_7bar;
  wire n11bar;
  wire n12bar;
  wire n13bar;
  wire n14bar;
  wire n15bar;
  wire n16bar;
  wire n17bar;
  wire n18bar;
  wire n19bar;
  wire n20bar;
//wire_done

  assign in_0 = in[0];
  assign out[7] = in_6;
  assign in_6  = in[6];
  assign out[6] = in_5;
  assign in_5  = in[5];
  assign out[5] = in_4;
  assign in_4  = in[4];
  assign out[2] = in_1;
  assign in_1  = in[1];
  assign out[0] = in_7;
  assign in_7  = in[7];
  assign in_0bar = inbar[0];
  assign outbar[7] = in_6bar;
  assign in_6bar = inbar[6];
  assign outbar[6] = in_5bar;
  assign in_5bar = inbar[5];
  assign outbar[5] = in_4bar;
  assign in_4bar = inbar[4];
  assign outbar[2] = in_1bar;
  assign in_1bar = inbar[1];
  assign outbar[0] = in_7bar;
  assign in_7bar = inbar[7];
//assign_done

  assign n20bar = in_7;
  assign n20 = in_7bar;
  assign n19bar = in[3];
  assign n19 = inbar[3];
  assign n18bar = in[2];
  assign n18 = inbar[2];
  assign n17bar = in_0;
  assign n17 = in_0bar;
  OR2_X1 U5 ( .A1(n16), .A2(n15), .ZN(out[4]) );
  AND2_X1 U5bar ( .A1(n16bar), .A2(n15bar), .ZN(outbar[4]) );
  AND2_X1 U6 ( .A1(in[3]), .A2(n20), .ZN(n15) );
  OR2_X1 U6bar ( .A1(inbar[3]), .A2(n20bar), .ZN(n15bar) );
  AND2_X1 U7 ( .A1(in_7), .A2(n19), .ZN(n16) );
  OR2_X1 U7bar ( .A1(in_7bar), .A2(n19bar), .ZN(n16bar) );
  OR2_X1 U8 ( .A1(n14), .A2(n13), .ZN(out[3]) );
  AND2_X1 U8bar ( .A1(n14bar), .A2(n13bar), .ZN(outbar[3]) );
  AND2_X1 U9 ( .A1(in[2]), .A2(n20), .ZN(n13) );
  OR2_X1 U9bar ( .A1(inbar[2]), .A2(n20bar), .ZN(n13bar) );
  AND2_X1 U10 ( .A1(in_7), .A2(n18), .ZN(n14) );
  OR2_X1 U10bar ( .A1(in_7bar), .A2(n18bar), .ZN(n14bar) );
  OR2_X1 U11 ( .A1(n12), .A2(n11), .ZN(out[1]) );
  AND2_X1 U11bar ( .A1(n12bar), .A2(n11bar), .ZN(outbar[1]) );
  AND2_X1 U12 ( .A1(in_0), .A2(n20), .ZN(n11) );
  OR2_X1 U12bar ( .A1(in_0bar), .A2(n20bar), .ZN(n11bar) );
  AND2_X1 U13 ( .A1(in_7), .A2(n17), .ZN(n12) );
  OR2_X1 U13bar ( .A1(in_7bar), .A2(n17bar), .ZN(n12bar) );
endmodule

module scale2_2 ( in, inbar, out, outbar );

  input wire [7:0] in;
  input wire [7:0] inbar;
//input_done

  output wire [7:0] out;
  output wire [7:0] outbar;
//output_done

  wire in_0;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_1;
  wire in_7;
  wire n11;
  wire n12;
  wire n13;
  wire n14;
  wire n15;
  wire n16;
  wire n17;
  wire n18;
  wire n19;
  wire n20;
  wire in_0bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_1bar;
  wire in_7bar;
  wire n11bar;
  wire n12bar;
  wire n13bar;
  wire n14bar;
  wire n15bar;
  wire n16bar;
  wire n17bar;
  wire n18bar;
  wire n19bar;
  wire n20bar;
//wire_done

  assign in_0 = in[0];
  assign out[7] = in_6;
  assign in_6  = in[6];
  assign out[6] = in_5;
  assign in_5  = in[5];
  assign out[5] = in_4;
  assign in_4  = in[4];
  assign out[2] = in_1;
  assign in_1  = in[1];
  assign out[0] = in_7;
  assign in_7  = in[7];
  assign in_0bar = inbar[0];
  assign outbar[7] = in_6bar;
  assign in_6bar = inbar[6];
  assign outbar[6] = in_5bar;
  assign in_5bar = inbar[5];
  assign outbar[5] = in_4bar;
  assign in_4bar = inbar[4];
  assign outbar[2] = in_1bar;
  assign in_1bar = inbar[1];
  assign outbar[0] = in_7bar;
  assign in_7bar = inbar[7];
//assign_done

  assign n20bar = in_7;
  assign n20 = in_7bar;
  assign n19bar = in[3];
  assign n19 = inbar[3];
  assign n18bar = in[2];
  assign n18 = inbar[2];
  assign n17bar = in_0;
  assign n17 = in_0bar;
  OR2_X1 U5 ( .A1(n16), .A2(n15), .ZN(out[4]) );
  AND2_X1 U5bar ( .A1(n16bar), .A2(n15bar), .ZN(outbar[4]) );
  AND2_X1 U6 ( .A1(in[3]), .A2(n20), .ZN(n15) );
  OR2_X1 U6bar ( .A1(inbar[3]), .A2(n20bar), .ZN(n15bar) );
  AND2_X1 U7 ( .A1(in_7), .A2(n19), .ZN(n16) );
  OR2_X1 U7bar ( .A1(in_7bar), .A2(n19bar), .ZN(n16bar) );
  OR2_X1 U8 ( .A1(n14), .A2(n13), .ZN(out[3]) );
  AND2_X1 U8bar ( .A1(n14bar), .A2(n13bar), .ZN(outbar[3]) );
  AND2_X1 U9 ( .A1(in[2]), .A2(n20), .ZN(n13) );
  OR2_X1 U9bar ( .A1(inbar[2]), .A2(n20bar), .ZN(n13bar) );
  AND2_X1 U10 ( .A1(in_7), .A2(n18), .ZN(n14) );
  OR2_X1 U10bar ( .A1(in_7bar), .A2(n18bar), .ZN(n14bar) );
  OR2_X1 U11 ( .A1(n12), .A2(n11), .ZN(out[1]) );
  AND2_X1 U11bar ( .A1(n12bar), .A2(n11bar), .ZN(outbar[1]) );
  AND2_X1 U12 ( .A1(in_0), .A2(n20), .ZN(n11) );
  OR2_X1 U12bar ( .A1(in_0bar), .A2(n20bar), .ZN(n11bar) );
  AND2_X1 U13 ( .A1(in_7), .A2(n17), .ZN(n12) );
  OR2_X1 U13bar ( .A1(in_7bar), .A2(n17bar), .ZN(n12bar) );
endmodule

module scale2_3 ( in, inbar, out, outbar );

  input wire [7:0] in;
  input wire [7:0] inbar;
//input_done

  output wire [7:0] out;
  output wire [7:0] outbar;
//output_done

  wire in_0;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_1;
  wire in_7;
  wire n11;
  wire n12;
  wire n13;
  wire n14;
  wire n15;
  wire n16;
  wire n17;
  wire n18;
  wire n19;
  wire n20;
  wire in_0bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_1bar;
  wire in_7bar;
  wire n11bar;
  wire n12bar;
  wire n13bar;
  wire n14bar;
  wire n15bar;
  wire n16bar;
  wire n17bar;
  wire n18bar;
  wire n19bar;
  wire n20bar;
//wire_done

  assign in_0 = in[0];
  assign out[7] = in_6;
  assign in_6  = in[6];
  assign out[6] = in_5;
  assign in_5  = in[5];
  assign out[5] = in_4;
  assign in_4  = in[4];
  assign out[2] = in_1;
  assign in_1  = in[1];
  assign out[0] = in_7;
  assign in_7  = in[7];
  assign in_0bar = inbar[0];
  assign outbar[7] = in_6bar;
  assign in_6bar = inbar[6];
  assign outbar[6] = in_5bar;
  assign in_5bar = inbar[5];
  assign outbar[5] = in_4bar;
  assign in_4bar = inbar[4];
  assign outbar[2] = in_1bar;
  assign in_1bar = inbar[1];
  assign outbar[0] = in_7bar;
  assign in_7bar = inbar[7];
//assign_done

  assign n20bar = in_7;
  assign n20 = in_7bar;
  assign n19bar = in[3];
  assign n19 = inbar[3];
  assign n18bar = in[2];
  assign n18 = inbar[2];
  assign n17bar = in_0;
  assign n17 = in_0bar;
  OR2_X1 U5 ( .A1(n16), .A2(n15), .ZN(out[4]) );
  AND2_X1 U5bar ( .A1(n16bar), .A2(n15bar), .ZN(outbar[4]) );
  AND2_X1 U6 ( .A1(in[3]), .A2(n20), .ZN(n15) );
  OR2_X1 U6bar ( .A1(inbar[3]), .A2(n20bar), .ZN(n15bar) );
  AND2_X1 U7 ( .A1(in_7), .A2(n19), .ZN(n16) );
  OR2_X1 U7bar ( .A1(in_7bar), .A2(n19bar), .ZN(n16bar) );
  OR2_X1 U8 ( .A1(n14), .A2(n13), .ZN(out[3]) );
  AND2_X1 U8bar ( .A1(n14bar), .A2(n13bar), .ZN(outbar[3]) );
  AND2_X1 U9 ( .A1(in[2]), .A2(n20), .ZN(n13) );
  OR2_X1 U9bar ( .A1(inbar[2]), .A2(n20bar), .ZN(n13bar) );
  AND2_X1 U10 ( .A1(in_7), .A2(n18), .ZN(n14) );
  OR2_X1 U10bar ( .A1(in_7bar), .A2(n18bar), .ZN(n14bar) );
  OR2_X1 U11 ( .A1(n12), .A2(n11), .ZN(out[1]) );
  AND2_X1 U11bar ( .A1(n12bar), .A2(n11bar), .ZN(outbar[1]) );
  AND2_X1 U12 ( .A1(in_0), .A2(n20), .ZN(n11) );
  OR2_X1 U12bar ( .A1(in_0bar), .A2(n20bar), .ZN(n11bar) );
  AND2_X1 U13 ( .A1(in_7), .A2(n17), .ZN(n12) );
  OR2_X1 U13bar ( .A1(in_7bar), .A2(n17bar), .ZN(n12bar) );
endmodule

module scale2_4 ( in, inbar, out, outbar );

  input wire [7:0] in;
  input wire [7:0] inbar;
//input_done

  output wire [7:0] out;
  output wire [7:0] outbar;
//output_done

  wire in_0;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_1;
  wire in_7;
  wire n11;
  wire n12;
  wire n13;
  wire n14;
  wire n15;
  wire n16;
  wire n17;
  wire n18;
  wire n19;
  wire n20;
  wire in_0bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_1bar;
  wire in_7bar;
  wire n11bar;
  wire n12bar;
  wire n13bar;
  wire n14bar;
  wire n15bar;
  wire n16bar;
  wire n17bar;
  wire n18bar;
  wire n19bar;
  wire n20bar;
//wire_done

  assign in_0 = in[0];
  assign out[7] = in_6;
  assign in_6  = in[6];
  assign out[6] = in_5;
  assign in_5  = in[5];
  assign out[5] = in_4;
  assign in_4  = in[4];
  assign out[2] = in_1;
  assign in_1  = in[1];
  assign out[0] = in_7;
  assign in_7  = in[7];
  assign in_0bar = inbar[0];
  assign outbar[7] = in_6bar;
  assign in_6bar = inbar[6];
  assign outbar[6] = in_5bar;
  assign in_5bar = inbar[5];
  assign outbar[5] = in_4bar;
  assign in_4bar = inbar[4];
  assign outbar[2] = in_1bar;
  assign in_1bar = inbar[1];
  assign outbar[0] = in_7bar;
  assign in_7bar = inbar[7];
//assign_done

  assign n20bar = in_7;
  assign n20 = in_7bar;
  assign n19bar = in[3];
  assign n19 = inbar[3];
  assign n18bar = in[2];
  assign n18 = inbar[2];
  assign n17bar = in_0;
  assign n17 = in_0bar;
  OR2_X1 U5 ( .A1(n16), .A2(n15), .ZN(out[4]) );
  AND2_X1 U5bar ( .A1(n16bar), .A2(n15bar), .ZN(outbar[4]) );
  AND2_X1 U6 ( .A1(in[3]), .A2(n20), .ZN(n15) );
  OR2_X1 U6bar ( .A1(inbar[3]), .A2(n20bar), .ZN(n15bar) );
  AND2_X1 U7 ( .A1(in_7), .A2(n19), .ZN(n16) );
  OR2_X1 U7bar ( .A1(in_7bar), .A2(n19bar), .ZN(n16bar) );
  OR2_X1 U8 ( .A1(n14), .A2(n13), .ZN(out[3]) );
  AND2_X1 U8bar ( .A1(n14bar), .A2(n13bar), .ZN(outbar[3]) );
  AND2_X1 U9 ( .A1(in[2]), .A2(n20), .ZN(n13) );
  OR2_X1 U9bar ( .A1(inbar[2]), .A2(n20bar), .ZN(n13bar) );
  AND2_X1 U10 ( .A1(in_7), .A2(n18), .ZN(n14) );
  OR2_X1 U10bar ( .A1(in_7bar), .A2(n18bar), .ZN(n14bar) );
  OR2_X1 U11 ( .A1(n12), .A2(n11), .ZN(out[1]) );
  AND2_X1 U11bar ( .A1(n12bar), .A2(n11bar), .ZN(outbar[1]) );
  AND2_X1 U12 ( .A1(in_0), .A2(n20), .ZN(n11) );
  OR2_X1 U12bar ( .A1(in_0bar), .A2(n20bar), .ZN(n11bar) );
  AND2_X1 U13 ( .A1(in_7), .A2(n17), .ZN(n12) );
  OR2_X1 U13bar ( .A1(in_7bar), .A2(n17bar), .ZN(n12bar) );
endmodule

module byteXor_2 ( a, abar, b, bbar, y, ybar );

  input wire [7:0] a;
  input wire [7:0] b;
  input wire [7:0] abar;
  input wire [7:0] bbar;
//input_done

  output wire [7:0] y;
  output wire [7:0] ybar;
//output_done

  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n33bar;
  wire n34bar;
  wire n35bar;
  wire n36bar;
  wire n37bar;
  wire n38bar;
  wire n39bar;
  wire n40bar;
  wire n41bar;
  wire n42bar;
  wire n43bar;
  wire n44bar;
  wire n45bar;
  wire n46bar;
  wire n47bar;
  wire n48bar;
  wire n49bar;
  wire n50bar;
  wire n51bar;
  wire n52bar;
  wire n53bar;
  wire n54bar;
  wire n55bar;
  wire n56bar;
  wire n57bar;
  wire n58bar;
  wire n59bar;
  wire n60bar;
  wire n61bar;
  wire n62bar;
  wire n63bar;
  wire n64bar;
//wire_done

 //assign_done

  assign n64bar = n47;
  assign n64 = n47bar;
  assign n63bar = a[7];
  assign n63 = abar[7];
  assign n62bar = n45;
  assign n62 = n45bar;
  assign n61bar = a[6];
  assign n61 = abar[6];
  assign n60bar = n43;
  assign n60 = n43bar;
  assign n59bar = a[5];
  assign n59 = abar[5];
  assign n58bar = n41;
  assign n58 = n41bar;
  assign n57bar = a[4];
  assign n57 = abar[4];
  assign n56bar = n39;
  assign n56 = n39bar;
  assign n55bar = a[3];
  assign n55 = abar[3];
  assign n54bar = n37;
  assign n54 = n37bar;
  assign n53bar = a[2];
  assign n53 = abar[2];
  assign n52bar = n35;
  assign n52 = n35bar;
  assign n51bar = a[1];
  assign n51 = abar[1];
  assign n50bar = n33;
  assign n50 = n33bar;
  assign n49bar = a[0];
  assign n49 = abar[0];
  OR2_X1 U17 ( .A1(n48), .A2(n64), .ZN(y[7]) );
  AND2_X1 U17bar ( .A1(n48bar), .A2(n64bar), .ZN(ybar[7]) );
  OR2_X1 U18 ( .A1(n63), .A2(b[7]), .ZN(n47) );
  AND2_X1 U18bar ( .A1(n63bar), .A2(bbar[7]), .ZN(n47bar) );
  AND2_X1 U19 ( .A1(b[7]), .A2(n63), .ZN(n48) );
  OR2_X1 U19bar ( .A1(bbar[7]), .A2(n63bar), .ZN(n48bar) );
  OR2_X1 U20 ( .A1(n46), .A2(n62), .ZN(y[6]) );
  AND2_X1 U20bar ( .A1(n46bar), .A2(n62bar), .ZN(ybar[6]) );
  OR2_X1 U21 ( .A1(n61), .A2(b[6]), .ZN(n45) );
  AND2_X1 U21bar ( .A1(n61bar), .A2(bbar[6]), .ZN(n45bar) );
  AND2_X1 U22 ( .A1(b[6]), .A2(n61), .ZN(n46) );
  OR2_X1 U22bar ( .A1(bbar[6]), .A2(n61bar), .ZN(n46bar) );
  OR2_X1 U23 ( .A1(n44), .A2(n60), .ZN(y[5]) );
  AND2_X1 U23bar ( .A1(n44bar), .A2(n60bar), .ZN(ybar[5]) );
  OR2_X1 U24 ( .A1(n59), .A2(b[5]), .ZN(n43) );
  AND2_X1 U24bar ( .A1(n59bar), .A2(bbar[5]), .ZN(n43bar) );
  AND2_X1 U25 ( .A1(b[5]), .A2(n59), .ZN(n44) );
  OR2_X1 U25bar ( .A1(bbar[5]), .A2(n59bar), .ZN(n44bar) );
  OR2_X1 U26 ( .A1(n42), .A2(n58), .ZN(y[4]) );
  AND2_X1 U26bar ( .A1(n42bar), .A2(n58bar), .ZN(ybar[4]) );
  OR2_X1 U27 ( .A1(n57), .A2(b[4]), .ZN(n41) );
  AND2_X1 U27bar ( .A1(n57bar), .A2(bbar[4]), .ZN(n41bar) );
  AND2_X1 U28 ( .A1(b[4]), .A2(n57), .ZN(n42) );
  OR2_X1 U28bar ( .A1(bbar[4]), .A2(n57bar), .ZN(n42bar) );
  OR2_X1 U29 ( .A1(n40), .A2(n56), .ZN(y[3]) );
  AND2_X1 U29bar ( .A1(n40bar), .A2(n56bar), .ZN(ybar[3]) );
  OR2_X1 U30 ( .A1(n55), .A2(b[3]), .ZN(n39) );
  AND2_X1 U30bar ( .A1(n55bar), .A2(bbar[3]), .ZN(n39bar) );
  AND2_X1 U31 ( .A1(b[3]), .A2(n55), .ZN(n40) );
  OR2_X1 U31bar ( .A1(bbar[3]), .A2(n55bar), .ZN(n40bar) );
  OR2_X1 U32 ( .A1(n38), .A2(n54), .ZN(y[2]) );
  AND2_X1 U32bar ( .A1(n38bar), .A2(n54bar), .ZN(ybar[2]) );
  OR2_X1 U33 ( .A1(n53), .A2(b[2]), .ZN(n37) );
  AND2_X1 U33bar ( .A1(n53bar), .A2(bbar[2]), .ZN(n37bar) );
  AND2_X1 U34 ( .A1(b[2]), .A2(n53), .ZN(n38) );
  OR2_X1 U34bar ( .A1(bbar[2]), .A2(n53bar), .ZN(n38bar) );
  OR2_X1 U35 ( .A1(n36), .A2(n52), .ZN(y[1]) );
  AND2_X1 U35bar ( .A1(n36bar), .A2(n52bar), .ZN(ybar[1]) );
  OR2_X1 U36 ( .A1(n51), .A2(b[1]), .ZN(n35) );
  AND2_X1 U36bar ( .A1(n51bar), .A2(bbar[1]), .ZN(n35bar) );
  AND2_X1 U37 ( .A1(b[1]), .A2(n51), .ZN(n36) );
  OR2_X1 U37bar ( .A1(bbar[1]), .A2(n51bar), .ZN(n36bar) );
  OR2_X1 U38 ( .A1(n34), .A2(n50), .ZN(y[0]) );
  AND2_X1 U38bar ( .A1(n34bar), .A2(n50bar), .ZN(ybar[0]) );
  OR2_X1 U39 ( .A1(n49), .A2(b[0]), .ZN(n33) );
  AND2_X1 U39bar ( .A1(n49bar), .A2(bbar[0]), .ZN(n33bar) );
  AND2_X1 U40 ( .A1(b[0]), .A2(n49), .ZN(n34) );
  OR2_X1 U40bar ( .A1(bbar[0]), .A2(n49bar), .ZN(n34bar) );
endmodule

module byteXor_3 ( a, abar, b, bbar, y, ybar );

  input wire [7:0] a;
  input wire [7:0] b;
  input wire [7:0] abar;
  input wire [7:0] bbar;
//input_done

  output wire [7:0] y;
  output wire [7:0] ybar;
//output_done

  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n33bar;
  wire n34bar;
  wire n35bar;
  wire n36bar;
  wire n37bar;
  wire n38bar;
  wire n39bar;
  wire n40bar;
  wire n41bar;
  wire n42bar;
  wire n43bar;
  wire n44bar;
  wire n45bar;
  wire n46bar;
  wire n47bar;
  wire n48bar;
  wire n49bar;
  wire n50bar;
  wire n51bar;
  wire n52bar;
  wire n53bar;
  wire n54bar;
  wire n55bar;
  wire n56bar;
  wire n57bar;
  wire n58bar;
  wire n59bar;
  wire n60bar;
  wire n61bar;
  wire n62bar;
  wire n63bar;
  wire n64bar;
//wire_done

 //assign_done

  assign n64bar = n47;
  assign n64 = n47bar;
  assign n63bar = a[7];
  assign n63 = abar[7];
  assign n62bar = n45;
  assign n62 = n45bar;
  assign n61bar = a[6];
  assign n61 = abar[6];
  assign n60bar = n43;
  assign n60 = n43bar;
  assign n59bar = a[5];
  assign n59 = abar[5];
  assign n58bar = n41;
  assign n58 = n41bar;
  assign n57bar = a[4];
  assign n57 = abar[4];
  assign n56bar = n39;
  assign n56 = n39bar;
  assign n55bar = a[3];
  assign n55 = abar[3];
  assign n54bar = n37;
  assign n54 = n37bar;
  assign n53bar = a[2];
  assign n53 = abar[2];
  assign n52bar = n35;
  assign n52 = n35bar;
  assign n51bar = a[1];
  assign n51 = abar[1];
  assign n50bar = n33;
  assign n50 = n33bar;
  assign n49bar = a[0];
  assign n49 = abar[0];
  OR2_X1 U17 ( .A1(n48), .A2(n64), .ZN(y[7]) );
  AND2_X1 U17bar ( .A1(n48bar), .A2(n64bar), .ZN(ybar[7]) );
  OR2_X1 U18 ( .A1(n63), .A2(b[7]), .ZN(n47) );
  AND2_X1 U18bar ( .A1(n63bar), .A2(bbar[7]), .ZN(n47bar) );
  AND2_X1 U19 ( .A1(b[7]), .A2(n63), .ZN(n48) );
  OR2_X1 U19bar ( .A1(bbar[7]), .A2(n63bar), .ZN(n48bar) );
  OR2_X1 U20 ( .A1(n46), .A2(n62), .ZN(y[6]) );
  AND2_X1 U20bar ( .A1(n46bar), .A2(n62bar), .ZN(ybar[6]) );
  OR2_X1 U21 ( .A1(n61), .A2(b[6]), .ZN(n45) );
  AND2_X1 U21bar ( .A1(n61bar), .A2(bbar[6]), .ZN(n45bar) );
  AND2_X1 U22 ( .A1(b[6]), .A2(n61), .ZN(n46) );
  OR2_X1 U22bar ( .A1(bbar[6]), .A2(n61bar), .ZN(n46bar) );
  OR2_X1 U23 ( .A1(n44), .A2(n60), .ZN(y[5]) );
  AND2_X1 U23bar ( .A1(n44bar), .A2(n60bar), .ZN(ybar[5]) );
  OR2_X1 U24 ( .A1(n59), .A2(b[5]), .ZN(n43) );
  AND2_X1 U24bar ( .A1(n59bar), .A2(bbar[5]), .ZN(n43bar) );
  AND2_X1 U25 ( .A1(b[5]), .A2(n59), .ZN(n44) );
  OR2_X1 U25bar ( .A1(bbar[5]), .A2(n59bar), .ZN(n44bar) );
  OR2_X1 U26 ( .A1(n42), .A2(n58), .ZN(y[4]) );
  AND2_X1 U26bar ( .A1(n42bar), .A2(n58bar), .ZN(ybar[4]) );
  OR2_X1 U27 ( .A1(n57), .A2(b[4]), .ZN(n41) );
  AND2_X1 U27bar ( .A1(n57bar), .A2(bbar[4]), .ZN(n41bar) );
  AND2_X1 U28 ( .A1(b[4]), .A2(n57), .ZN(n42) );
  OR2_X1 U28bar ( .A1(bbar[4]), .A2(n57bar), .ZN(n42bar) );
  OR2_X1 U29 ( .A1(n40), .A2(n56), .ZN(y[3]) );
  AND2_X1 U29bar ( .A1(n40bar), .A2(n56bar), .ZN(ybar[3]) );
  OR2_X1 U30 ( .A1(n55), .A2(b[3]), .ZN(n39) );
  AND2_X1 U30bar ( .A1(n55bar), .A2(bbar[3]), .ZN(n39bar) );
  AND2_X1 U31 ( .A1(b[3]), .A2(n55), .ZN(n40) );
  OR2_X1 U31bar ( .A1(bbar[3]), .A2(n55bar), .ZN(n40bar) );
  OR2_X1 U32 ( .A1(n38), .A2(n54), .ZN(y[2]) );
  AND2_X1 U32bar ( .A1(n38bar), .A2(n54bar), .ZN(ybar[2]) );
  OR2_X1 U33 ( .A1(n53), .A2(b[2]), .ZN(n37) );
  AND2_X1 U33bar ( .A1(n53bar), .A2(bbar[2]), .ZN(n37bar) );
  AND2_X1 U34 ( .A1(b[2]), .A2(n53), .ZN(n38) );
  OR2_X1 U34bar ( .A1(bbar[2]), .A2(n53bar), .ZN(n38bar) );
  OR2_X1 U35 ( .A1(n36), .A2(n52), .ZN(y[1]) );
  AND2_X1 U35bar ( .A1(n36bar), .A2(n52bar), .ZN(ybar[1]) );
  OR2_X1 U36 ( .A1(n51), .A2(b[1]), .ZN(n35) );
  AND2_X1 U36bar ( .A1(n51bar), .A2(bbar[1]), .ZN(n35bar) );
  AND2_X1 U37 ( .A1(b[1]), .A2(n51), .ZN(n36) );
  OR2_X1 U37bar ( .A1(bbar[1]), .A2(n51bar), .ZN(n36bar) );
  OR2_X1 U38 ( .A1(n34), .A2(n50), .ZN(y[0]) );
  AND2_X1 U38bar ( .A1(n34bar), .A2(n50bar), .ZN(ybar[0]) );
  OR2_X1 U39 ( .A1(n49), .A2(b[0]), .ZN(n33) );
  AND2_X1 U39bar ( .A1(n49bar), .A2(bbar[0]), .ZN(n33bar) );
  AND2_X1 U40 ( .A1(b[0]), .A2(n49), .ZN(n34) );
  OR2_X1 U40bar ( .A1(bbar[0]), .A2(n49bar), .ZN(n34bar) );
endmodule

module byteXor_4 ( a, abar, b, bbar, y, ybar );

  input wire [7:0] a;
  input wire [7:0] b;
  input wire [7:0] abar;
  input wire [7:0] bbar;
//input_done

  output wire [7:0] y;
  output wire [7:0] ybar;
//output_done

  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n33bar;
  wire n34bar;
  wire n35bar;
  wire n36bar;
  wire n37bar;
  wire n38bar;
  wire n39bar;
  wire n40bar;
  wire n41bar;
  wire n42bar;
  wire n43bar;
  wire n44bar;
  wire n45bar;
  wire n46bar;
  wire n47bar;
  wire n48bar;
  wire n49bar;
  wire n50bar;
  wire n51bar;
  wire n52bar;
  wire n53bar;
  wire n54bar;
  wire n55bar;
  wire n56bar;
  wire n57bar;
  wire n58bar;
  wire n59bar;
  wire n60bar;
  wire n61bar;
  wire n62bar;
  wire n63bar;
  wire n64bar;
//wire_done

 //assign_done

  assign n64bar = n47;
  assign n64 = n47bar;
  assign n63bar = a[7];
  assign n63 = abar[7];
  assign n62bar = n45;
  assign n62 = n45bar;
  assign n61bar = a[6];
  assign n61 = abar[6];
  assign n60bar = n43;
  assign n60 = n43bar;
  assign n59bar = a[5];
  assign n59 = abar[5];
  assign n58bar = n41;
  assign n58 = n41bar;
  assign n57bar = a[4];
  assign n57 = abar[4];
  assign n56bar = n39;
  assign n56 = n39bar;
  assign n55bar = a[3];
  assign n55 = abar[3];
  assign n54bar = n37;
  assign n54 = n37bar;
  assign n53bar = a[2];
  assign n53 = abar[2];
  assign n52bar = n35;
  assign n52 = n35bar;
  assign n51bar = a[1];
  assign n51 = abar[1];
  assign n50bar = n33;
  assign n50 = n33bar;
  assign n49bar = a[0];
  assign n49 = abar[0];
  OR2_X1 U17 ( .A1(n48), .A2(n64), .ZN(y[7]) );
  AND2_X1 U17bar ( .A1(n48bar), .A2(n64bar), .ZN(ybar[7]) );
  OR2_X1 U18 ( .A1(n63), .A2(b[7]), .ZN(n47) );
  AND2_X1 U18bar ( .A1(n63bar), .A2(bbar[7]), .ZN(n47bar) );
  AND2_X1 U19 ( .A1(b[7]), .A2(n63), .ZN(n48) );
  OR2_X1 U19bar ( .A1(bbar[7]), .A2(n63bar), .ZN(n48bar) );
  OR2_X1 U20 ( .A1(n46), .A2(n62), .ZN(y[6]) );
  AND2_X1 U20bar ( .A1(n46bar), .A2(n62bar), .ZN(ybar[6]) );
  OR2_X1 U21 ( .A1(n61), .A2(b[6]), .ZN(n45) );
  AND2_X1 U21bar ( .A1(n61bar), .A2(bbar[6]), .ZN(n45bar) );
  AND2_X1 U22 ( .A1(b[6]), .A2(n61), .ZN(n46) );
  OR2_X1 U22bar ( .A1(bbar[6]), .A2(n61bar), .ZN(n46bar) );
  OR2_X1 U23 ( .A1(n44), .A2(n60), .ZN(y[5]) );
  AND2_X1 U23bar ( .A1(n44bar), .A2(n60bar), .ZN(ybar[5]) );
  OR2_X1 U24 ( .A1(n59), .A2(b[5]), .ZN(n43) );
  AND2_X1 U24bar ( .A1(n59bar), .A2(bbar[5]), .ZN(n43bar) );
  AND2_X1 U25 ( .A1(b[5]), .A2(n59), .ZN(n44) );
  OR2_X1 U25bar ( .A1(bbar[5]), .A2(n59bar), .ZN(n44bar) );
  OR2_X1 U26 ( .A1(n42), .A2(n58), .ZN(y[4]) );
  AND2_X1 U26bar ( .A1(n42bar), .A2(n58bar), .ZN(ybar[4]) );
  OR2_X1 U27 ( .A1(n57), .A2(b[4]), .ZN(n41) );
  AND2_X1 U27bar ( .A1(n57bar), .A2(bbar[4]), .ZN(n41bar) );
  AND2_X1 U28 ( .A1(b[4]), .A2(n57), .ZN(n42) );
  OR2_X1 U28bar ( .A1(bbar[4]), .A2(n57bar), .ZN(n42bar) );
  OR2_X1 U29 ( .A1(n40), .A2(n56), .ZN(y[3]) );
  AND2_X1 U29bar ( .A1(n40bar), .A2(n56bar), .ZN(ybar[3]) );
  OR2_X1 U30 ( .A1(n55), .A2(b[3]), .ZN(n39) );
  AND2_X1 U30bar ( .A1(n55bar), .A2(bbar[3]), .ZN(n39bar) );
  AND2_X1 U31 ( .A1(b[3]), .A2(n55), .ZN(n40) );
  OR2_X1 U31bar ( .A1(bbar[3]), .A2(n55bar), .ZN(n40bar) );
  OR2_X1 U32 ( .A1(n38), .A2(n54), .ZN(y[2]) );
  AND2_X1 U32bar ( .A1(n38bar), .A2(n54bar), .ZN(ybar[2]) );
  OR2_X1 U33 ( .A1(n53), .A2(b[2]), .ZN(n37) );
  AND2_X1 U33bar ( .A1(n53bar), .A2(bbar[2]), .ZN(n37bar) );
  AND2_X1 U34 ( .A1(b[2]), .A2(n53), .ZN(n38) );
  OR2_X1 U34bar ( .A1(bbar[2]), .A2(n53bar), .ZN(n38bar) );
  OR2_X1 U35 ( .A1(n36), .A2(n52), .ZN(y[1]) );
  AND2_X1 U35bar ( .A1(n36bar), .A2(n52bar), .ZN(ybar[1]) );
  OR2_X1 U36 ( .A1(n51), .A2(b[1]), .ZN(n35) );
  AND2_X1 U36bar ( .A1(n51bar), .A2(bbar[1]), .ZN(n35bar) );
  AND2_X1 U37 ( .A1(b[1]), .A2(n51), .ZN(n36) );
  OR2_X1 U37bar ( .A1(bbar[1]), .A2(n51bar), .ZN(n36bar) );
  OR2_X1 U38 ( .A1(n34), .A2(n50), .ZN(y[0]) );
  AND2_X1 U38bar ( .A1(n34bar), .A2(n50bar), .ZN(ybar[0]) );
  OR2_X1 U39 ( .A1(n49), .A2(b[0]), .ZN(n33) );
  AND2_X1 U39bar ( .A1(n49bar), .A2(bbar[0]), .ZN(n33bar) );
  AND2_X1 U40 ( .A1(b[0]), .A2(n49), .ZN(n34) );
  OR2_X1 U40bar ( .A1(bbar[0]), .A2(n49bar), .ZN(n34bar) );
endmodule

module byteXor_5 ( a, abar, b, bbar, y, ybar );

  input wire [7:0] a;
  input wire [7:0] b;
  input wire [7:0] abar;
  input wire [7:0] bbar;
//input_done

  output wire [7:0] y;
  output wire [7:0] ybar;
//output_done

  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n33bar;
  wire n34bar;
  wire n35bar;
  wire n36bar;
  wire n37bar;
  wire n38bar;
  wire n39bar;
  wire n40bar;
  wire n41bar;
  wire n42bar;
  wire n43bar;
  wire n44bar;
  wire n45bar;
  wire n46bar;
  wire n47bar;
  wire n48bar;
  wire n49bar;
  wire n50bar;
  wire n51bar;
  wire n52bar;
  wire n53bar;
  wire n54bar;
  wire n55bar;
  wire n56bar;
  wire n57bar;
  wire n58bar;
  wire n59bar;
  wire n60bar;
  wire n61bar;
  wire n62bar;
  wire n63bar;
  wire n64bar;
//wire_done

 //assign_done

  assign n64bar = n47;
  assign n64 = n47bar;
  assign n63bar = a[7];
  assign n63 = abar[7];
  assign n62bar = n45;
  assign n62 = n45bar;
  assign n61bar = a[6];
  assign n61 = abar[6];
  assign n60bar = n43;
  assign n60 = n43bar;
  assign n59bar = a[5];
  assign n59 = abar[5];
  assign n58bar = n41;
  assign n58 = n41bar;
  assign n57bar = a[4];
  assign n57 = abar[4];
  assign n56bar = n39;
  assign n56 = n39bar;
  assign n55bar = a[3];
  assign n55 = abar[3];
  assign n54bar = n37;
  assign n54 = n37bar;
  assign n53bar = a[2];
  assign n53 = abar[2];
  assign n52bar = n35;
  assign n52 = n35bar;
  assign n51bar = a[1];
  assign n51 = abar[1];
  assign n50bar = n33;
  assign n50 = n33bar;
  assign n49bar = a[0];
  assign n49 = abar[0];
  OR2_X1 U17 ( .A1(n48), .A2(n64), .ZN(y[7]) );
  AND2_X1 U17bar ( .A1(n48bar), .A2(n64bar), .ZN(ybar[7]) );
  OR2_X1 U18 ( .A1(n63), .A2(b[7]), .ZN(n47) );
  AND2_X1 U18bar ( .A1(n63bar), .A2(bbar[7]), .ZN(n47bar) );
  AND2_X1 U19 ( .A1(b[7]), .A2(n63), .ZN(n48) );
  OR2_X1 U19bar ( .A1(bbar[7]), .A2(n63bar), .ZN(n48bar) );
  OR2_X1 U20 ( .A1(n46), .A2(n62), .ZN(y[6]) );
  AND2_X1 U20bar ( .A1(n46bar), .A2(n62bar), .ZN(ybar[6]) );
  OR2_X1 U21 ( .A1(n61), .A2(b[6]), .ZN(n45) );
  AND2_X1 U21bar ( .A1(n61bar), .A2(bbar[6]), .ZN(n45bar) );
  AND2_X1 U22 ( .A1(b[6]), .A2(n61), .ZN(n46) );
  OR2_X1 U22bar ( .A1(bbar[6]), .A2(n61bar), .ZN(n46bar) );
  OR2_X1 U23 ( .A1(n44), .A2(n60), .ZN(y[5]) );
  AND2_X1 U23bar ( .A1(n44bar), .A2(n60bar), .ZN(ybar[5]) );
  OR2_X1 U24 ( .A1(n59), .A2(b[5]), .ZN(n43) );
  AND2_X1 U24bar ( .A1(n59bar), .A2(bbar[5]), .ZN(n43bar) );
  AND2_X1 U25 ( .A1(b[5]), .A2(n59), .ZN(n44) );
  OR2_X1 U25bar ( .A1(bbar[5]), .A2(n59bar), .ZN(n44bar) );
  OR2_X1 U26 ( .A1(n42), .A2(n58), .ZN(y[4]) );
  AND2_X1 U26bar ( .A1(n42bar), .A2(n58bar), .ZN(ybar[4]) );
  OR2_X1 U27 ( .A1(n57), .A2(b[4]), .ZN(n41) );
  AND2_X1 U27bar ( .A1(n57bar), .A2(bbar[4]), .ZN(n41bar) );
  AND2_X1 U28 ( .A1(b[4]), .A2(n57), .ZN(n42) );
  OR2_X1 U28bar ( .A1(bbar[4]), .A2(n57bar), .ZN(n42bar) );
  OR2_X1 U29 ( .A1(n40), .A2(n56), .ZN(y[3]) );
  AND2_X1 U29bar ( .A1(n40bar), .A2(n56bar), .ZN(ybar[3]) );
  OR2_X1 U30 ( .A1(n55), .A2(b[3]), .ZN(n39) );
  AND2_X1 U30bar ( .A1(n55bar), .A2(bbar[3]), .ZN(n39bar) );
  AND2_X1 U31 ( .A1(b[3]), .A2(n55), .ZN(n40) );
  OR2_X1 U31bar ( .A1(bbar[3]), .A2(n55bar), .ZN(n40bar) );
  OR2_X1 U32 ( .A1(n38), .A2(n54), .ZN(y[2]) );
  AND2_X1 U32bar ( .A1(n38bar), .A2(n54bar), .ZN(ybar[2]) );
  OR2_X1 U33 ( .A1(n53), .A2(b[2]), .ZN(n37) );
  AND2_X1 U33bar ( .A1(n53bar), .A2(bbar[2]), .ZN(n37bar) );
  AND2_X1 U34 ( .A1(b[2]), .A2(n53), .ZN(n38) );
  OR2_X1 U34bar ( .A1(bbar[2]), .A2(n53bar), .ZN(n38bar) );
  OR2_X1 U35 ( .A1(n36), .A2(n52), .ZN(y[1]) );
  AND2_X1 U35bar ( .A1(n36bar), .A2(n52bar), .ZN(ybar[1]) );
  OR2_X1 U36 ( .A1(n51), .A2(b[1]), .ZN(n35) );
  AND2_X1 U36bar ( .A1(n51bar), .A2(bbar[1]), .ZN(n35bar) );
  AND2_X1 U37 ( .A1(b[1]), .A2(n51), .ZN(n36) );
  OR2_X1 U37bar ( .A1(bbar[1]), .A2(n51bar), .ZN(n36bar) );
  OR2_X1 U38 ( .A1(n34), .A2(n50), .ZN(y[0]) );
  AND2_X1 U38bar ( .A1(n34bar), .A2(n50bar), .ZN(ybar[0]) );
  OR2_X1 U39 ( .A1(n49), .A2(b[0]), .ZN(n33) );
  AND2_X1 U39bar ( .A1(n49bar), .A2(bbar[0]), .ZN(n33bar) );
  AND2_X1 U40 ( .A1(b[0]), .A2(n49), .ZN(n34) );
  OR2_X1 U40bar ( .A1(bbar[0]), .A2(n49bar), .ZN(n34bar) );
endmodule

module byteXor4_1 ( a, abar, b, bbar, c, cbar, d, dbar, y, ybar );

  input wire [7:0] a;
  input wire [7:0] b;
  input wire [7:0] c;
  input wire [7:0] d;
  input wire [7:0] abar;
  input wire [7:0] bbar;
  input wire [7:0] cbar;
  input wire [7:0] dbar;
//input_done

  output wire [7:0] y;
  output wire [7:0] ybar;
//output_done

  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n113bar;
  wire n114bar;
  wire n115bar;
  wire n116bar;
  wire n117bar;
  wire n118bar;
  wire n119bar;
  wire n120bar;
  wire n121bar;
  wire n122bar;
  wire n123bar;
  wire n124bar;
  wire n125bar;
  wire n126bar;
  wire n127bar;
  wire n128bar;
  wire n129bar;
  wire n130bar;
  wire n131bar;
  wire n132bar;
  wire n133bar;
  wire n134bar;
  wire n135bar;
  wire n136bar;
  wire n137bar;
  wire n138bar;
  wire n139bar;
  wire n140bar;
  wire n141bar;
  wire n142bar;
  wire n143bar;
  wire n144bar;
  wire n145bar;
  wire n146bar;
  wire n147bar;
  wire n148bar;
  wire n149bar;
  wire n150bar;
  wire n151bar;
  wire n152bar;
  wire n153bar;
  wire n154bar;
  wire n155bar;
  wire n156bar;
  wire n157bar;
  wire n158bar;
  wire n159bar;
  wire n160bar;
  wire n161bar;
  wire n162bar;
  wire n163bar;
  wire n164bar;
  wire n165bar;
  wire n166bar;
  wire n167bar;
  wire n168bar;
  wire n169bar;
  wire n170bar;
  wire n171bar;
  wire n172bar;
  wire n173bar;
  wire n174bar;
  wire n175bar;
  wire n176bar;
  wire n177bar;
  wire n178bar;
  wire n179bar;
  wire n180bar;
  wire n181bar;
  wire n182bar;
  wire n183bar;
  wire n184bar;
  wire n185bar;
  wire n186bar;
  wire n187bar;
  wire n188bar;
  wire n189bar;
  wire n190bar;
  wire n191bar;
  wire n192bar;
  wire n193bar;
  wire n194bar;
  wire n195bar;
  wire n196bar;
  wire n197bar;
  wire n198bar;
  wire n199bar;
  wire n200bar;
  wire n201bar;
  wire n202bar;
  wire n203bar;
  wire n204bar;
  wire n205bar;
  wire n206bar;
  wire n207bar;
  wire n208bar;
  wire n209bar;
  wire n210bar;
  wire n211bar;
  wire n212bar;
  wire n213bar;
  wire n214bar;
  wire n215bar;
  wire n216bar;
  wire n217bar;
  wire n218bar;
  wire n219bar;
  wire n220bar;
  wire n221bar;
  wire n222bar;
  wire n223bar;
  wire n224bar;
//wire_done

 //assign_done

  assign n224bar = n175;
  assign n224 = n175bar;
  assign n223bar = a[7];
  assign n223 = abar[7];
  assign n222bar = n167;
  assign n222 = n167bar;
  assign n221bar = a[6];
  assign n221 = abar[6];
  assign n220bar = n159;
  assign n220 = n159bar;
  assign n219bar = a[5];
  assign n219 = abar[5];
  assign n218bar = n151;
  assign n218 = n151bar;
  assign n217bar = a[4];
  assign n217 = abar[4];
  assign n216bar = n143;
  assign n216 = n143bar;
  assign n215bar = a[3];
  assign n215 = abar[3];
  assign n214bar = n135;
  assign n214 = n135bar;
  assign n213bar = a[2];
  assign n213 = abar[2];
  assign n212bar = n127;
  assign n212 = n127bar;
  assign n211bar = a[1];
  assign n211 = abar[1];
  assign n210bar = n119;
  assign n210 = n119bar;
  assign n209bar = a[0];
  assign n209 = abar[0];
  assign n208bar = b[7];
  assign n208 = bbar[7];
  assign n207bar = b[6];
  assign n207 = bbar[6];
  assign n206bar = b[5];
  assign n206 = bbar[5];
  assign n205bar = b[4];
  assign n205 = bbar[4];
  assign n204bar = b[3];
  assign n204 = bbar[3];
  assign n203bar = b[2];
  assign n203 = bbar[2];
  assign n202bar = b[1];
  assign n202 = bbar[1];
  assign n201bar = b[0];
  assign n201 = bbar[0];
  assign n200bar = n171;
  assign n200 = n171bar;
  assign n199bar = c[7];
  assign n199 = cbar[7];
  assign n198bar = n163;
  assign n198 = n163bar;
  assign n197bar = c[6];
  assign n197 = cbar[6];
  assign n196bar = n155;
  assign n196 = n155bar;
  assign n195bar = c[5];
  assign n195 = cbar[5];
  assign n194bar = n147;
  assign n194 = n147bar;
  assign n193bar = c[4];
  assign n193 = cbar[4];
  assign n192bar = n139;
  assign n192 = n139bar;
  assign n191bar = c[3];
  assign n191 = cbar[3];
  assign n190bar = n131;
  assign n190 = n131bar;
  assign n189bar = c[2];
  assign n189 = cbar[2];
  assign n188bar = n123;
  assign n188 = n123bar;
  assign n187bar = c[1];
  assign n187 = cbar[1];
  assign n186bar = n115;
  assign n186 = n115bar;
  assign n185bar = c[0];
  assign n185 = cbar[0];
  assign n184bar = d[7];
  assign n184 = dbar[7];
  assign n183bar = d[6];
  assign n183 = dbar[6];
  assign n182bar = d[5];
  assign n182 = dbar[5];
  assign n181bar = d[4];
  assign n181 = dbar[4];
  assign n180bar = d[3];
  assign n180 = dbar[3];
  assign n179bar = d[2];
  assign n179 = dbar[2];
  assign n178bar = d[1];
  assign n178 = dbar[1];
  assign n177bar = d[0];
  assign n177 = dbar[0];
  OR2_X1 U49 ( .A1(n176), .A2(n224), .ZN(y[7]) );
  AND2_X1 U49bar ( .A1(n176bar), .A2(n224bar), .ZN(ybar[7]) );
  OR2_X1 U50 ( .A1(n174), .A2(n200), .ZN(n175) );
  AND2_X1 U50bar ( .A1(n174bar), .A2(n200bar), .ZN(n175bar) );
  AND2_X1 U51 ( .A1(n200), .A2(n174), .ZN(n176) );
  OR2_X1 U51bar ( .A1(n200bar), .A2(n174bar), .ZN(n176bar) );
  AND2_X1 U52 ( .A1(n173), .A2(n172), .ZN(n174) );
  OR2_X1 U52bar ( .A1(n173bar), .A2(n172bar), .ZN(n174bar) );
  OR2_X1 U53 ( .A1(n223), .A2(b[7]), .ZN(n172) );
  AND2_X1 U53bar ( .A1(n223bar), .A2(bbar[7]), .ZN(n172bar) );
  OR2_X1 U54 ( .A1(n208), .A2(a[7]), .ZN(n173) );
  AND2_X1 U54bar ( .A1(n208bar), .A2(abar[7]), .ZN(n173bar) );
  AND2_X1 U55 ( .A1(n170), .A2(n169), .ZN(n171) );
  OR2_X1 U55bar ( .A1(n170bar), .A2(n169bar), .ZN(n171bar) );
  OR2_X1 U56 ( .A1(n199), .A2(d[7]), .ZN(n169) );
  AND2_X1 U56bar ( .A1(n199bar), .A2(dbar[7]), .ZN(n169bar) );
  OR2_X1 U57 ( .A1(n184), .A2(c[7]), .ZN(n170) );
  AND2_X1 U57bar ( .A1(n184bar), .A2(cbar[7]), .ZN(n170bar) );
  OR2_X1 U58 ( .A1(n168), .A2(n222), .ZN(y[6]) );
  AND2_X1 U58bar ( .A1(n168bar), .A2(n222bar), .ZN(ybar[6]) );
  OR2_X1 U59 ( .A1(n166), .A2(n198), .ZN(n167) );
  AND2_X1 U59bar ( .A1(n166bar), .A2(n198bar), .ZN(n167bar) );
  AND2_X1 U60 ( .A1(n198), .A2(n166), .ZN(n168) );
  OR2_X1 U60bar ( .A1(n198bar), .A2(n166bar), .ZN(n168bar) );
  AND2_X1 U61 ( .A1(n165), .A2(n164), .ZN(n166) );
  OR2_X1 U61bar ( .A1(n165bar), .A2(n164bar), .ZN(n166bar) );
  OR2_X1 U62 ( .A1(n221), .A2(b[6]), .ZN(n164) );
  AND2_X1 U62bar ( .A1(n221bar), .A2(bbar[6]), .ZN(n164bar) );
  OR2_X1 U63 ( .A1(n207), .A2(a[6]), .ZN(n165) );
  AND2_X1 U63bar ( .A1(n207bar), .A2(abar[6]), .ZN(n165bar) );
  AND2_X1 U64 ( .A1(n162), .A2(n161), .ZN(n163) );
  OR2_X1 U64bar ( .A1(n162bar), .A2(n161bar), .ZN(n163bar) );
  OR2_X1 U65 ( .A1(n197), .A2(d[6]), .ZN(n161) );
  AND2_X1 U65bar ( .A1(n197bar), .A2(dbar[6]), .ZN(n161bar) );
  OR2_X1 U66 ( .A1(n183), .A2(c[6]), .ZN(n162) );
  AND2_X1 U66bar ( .A1(n183bar), .A2(cbar[6]), .ZN(n162bar) );
  OR2_X1 U67 ( .A1(n160), .A2(n220), .ZN(y[5]) );
  AND2_X1 U67bar ( .A1(n160bar), .A2(n220bar), .ZN(ybar[5]) );
  OR2_X1 U68 ( .A1(n158), .A2(n196), .ZN(n159) );
  AND2_X1 U68bar ( .A1(n158bar), .A2(n196bar), .ZN(n159bar) );
  AND2_X1 U69 ( .A1(n196), .A2(n158), .ZN(n160) );
  OR2_X1 U69bar ( .A1(n196bar), .A2(n158bar), .ZN(n160bar) );
  AND2_X1 U70 ( .A1(n157), .A2(n156), .ZN(n158) );
  OR2_X1 U70bar ( .A1(n157bar), .A2(n156bar), .ZN(n158bar) );
  OR2_X1 U71 ( .A1(n219), .A2(b[5]), .ZN(n156) );
  AND2_X1 U71bar ( .A1(n219bar), .A2(bbar[5]), .ZN(n156bar) );
  OR2_X1 U72 ( .A1(n206), .A2(a[5]), .ZN(n157) );
  AND2_X1 U72bar ( .A1(n206bar), .A2(abar[5]), .ZN(n157bar) );
  AND2_X1 U73 ( .A1(n154), .A2(n153), .ZN(n155) );
  OR2_X1 U73bar ( .A1(n154bar), .A2(n153bar), .ZN(n155bar) );
  OR2_X1 U74 ( .A1(n195), .A2(d[5]), .ZN(n153) );
  AND2_X1 U74bar ( .A1(n195bar), .A2(dbar[5]), .ZN(n153bar) );
  OR2_X1 U75 ( .A1(n182), .A2(c[5]), .ZN(n154) );
  AND2_X1 U75bar ( .A1(n182bar), .A2(cbar[5]), .ZN(n154bar) );
  OR2_X1 U76 ( .A1(n152), .A2(n218), .ZN(y[4]) );
  AND2_X1 U76bar ( .A1(n152bar), .A2(n218bar), .ZN(ybar[4]) );
  OR2_X1 U77 ( .A1(n150), .A2(n194), .ZN(n151) );
  AND2_X1 U77bar ( .A1(n150bar), .A2(n194bar), .ZN(n151bar) );
  AND2_X1 U78 ( .A1(n194), .A2(n150), .ZN(n152) );
  OR2_X1 U78bar ( .A1(n194bar), .A2(n150bar), .ZN(n152bar) );
  AND2_X1 U79 ( .A1(n149), .A2(n148), .ZN(n150) );
  OR2_X1 U79bar ( .A1(n149bar), .A2(n148bar), .ZN(n150bar) );
  OR2_X1 U80 ( .A1(n217), .A2(b[4]), .ZN(n148) );
  AND2_X1 U80bar ( .A1(n217bar), .A2(bbar[4]), .ZN(n148bar) );
  OR2_X1 U81 ( .A1(n205), .A2(a[4]), .ZN(n149) );
  AND2_X1 U81bar ( .A1(n205bar), .A2(abar[4]), .ZN(n149bar) );
  AND2_X1 U82 ( .A1(n146), .A2(n145), .ZN(n147) );
  OR2_X1 U82bar ( .A1(n146bar), .A2(n145bar), .ZN(n147bar) );
  OR2_X1 U83 ( .A1(n193), .A2(d[4]), .ZN(n145) );
  AND2_X1 U83bar ( .A1(n193bar), .A2(dbar[4]), .ZN(n145bar) );
  OR2_X1 U84 ( .A1(n181), .A2(c[4]), .ZN(n146) );
  AND2_X1 U84bar ( .A1(n181bar), .A2(cbar[4]), .ZN(n146bar) );
  OR2_X1 U85 ( .A1(n144), .A2(n216), .ZN(y[3]) );
  AND2_X1 U85bar ( .A1(n144bar), .A2(n216bar), .ZN(ybar[3]) );
  OR2_X1 U86 ( .A1(n142), .A2(n192), .ZN(n143) );
  AND2_X1 U86bar ( .A1(n142bar), .A2(n192bar), .ZN(n143bar) );
  AND2_X1 U87 ( .A1(n192), .A2(n142), .ZN(n144) );
  OR2_X1 U87bar ( .A1(n192bar), .A2(n142bar), .ZN(n144bar) );
  AND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(n142) );
  OR2_X1 U88bar ( .A1(n141bar), .A2(n140bar), .ZN(n142bar) );
  OR2_X1 U89 ( .A1(n215), .A2(b[3]), .ZN(n140) );
  AND2_X1 U89bar ( .A1(n215bar), .A2(bbar[3]), .ZN(n140bar) );
  OR2_X1 U90 ( .A1(n204), .A2(a[3]), .ZN(n141) );
  AND2_X1 U90bar ( .A1(n204bar), .A2(abar[3]), .ZN(n141bar) );
  AND2_X1 U91 ( .A1(n138), .A2(n137), .ZN(n139) );
  OR2_X1 U91bar ( .A1(n138bar), .A2(n137bar), .ZN(n139bar) );
  OR2_X1 U92 ( .A1(n191), .A2(d[3]), .ZN(n137) );
  AND2_X1 U92bar ( .A1(n191bar), .A2(dbar[3]), .ZN(n137bar) );
  OR2_X1 U93 ( .A1(n180), .A2(c[3]), .ZN(n138) );
  AND2_X1 U93bar ( .A1(n180bar), .A2(cbar[3]), .ZN(n138bar) );
  OR2_X1 U94 ( .A1(n136), .A2(n214), .ZN(y[2]) );
  AND2_X1 U94bar ( .A1(n136bar), .A2(n214bar), .ZN(ybar[2]) );
  OR2_X1 U95 ( .A1(n134), .A2(n190), .ZN(n135) );
  AND2_X1 U95bar ( .A1(n134bar), .A2(n190bar), .ZN(n135bar) );
  AND2_X1 U96 ( .A1(n190), .A2(n134), .ZN(n136) );
  OR2_X1 U96bar ( .A1(n190bar), .A2(n134bar), .ZN(n136bar) );
  AND2_X1 U97 ( .A1(n133), .A2(n132), .ZN(n134) );
  OR2_X1 U97bar ( .A1(n133bar), .A2(n132bar), .ZN(n134bar) );
  OR2_X1 U98 ( .A1(n213), .A2(b[2]), .ZN(n132) );
  AND2_X1 U98bar ( .A1(n213bar), .A2(bbar[2]), .ZN(n132bar) );
  OR2_X1 U99 ( .A1(n203), .A2(a[2]), .ZN(n133) );
  AND2_X1 U99bar ( .A1(n203bar), .A2(abar[2]), .ZN(n133bar) );
  AND2_X1 U100 ( .A1(n130), .A2(n129), .ZN(n131) );
  OR2_X1 U100bar ( .A1(n130bar), .A2(n129bar), .ZN(n131bar) );
  OR2_X1 U101 ( .A1(n189), .A2(d[2]), .ZN(n129) );
  AND2_X1 U101bar ( .A1(n189bar), .A2(dbar[2]), .ZN(n129bar) );
  OR2_X1 U102 ( .A1(n179), .A2(c[2]), .ZN(n130) );
  AND2_X1 U102bar ( .A1(n179bar), .A2(cbar[2]), .ZN(n130bar) );
  OR2_X1 U103 ( .A1(n128), .A2(n212), .ZN(y[1]) );
  AND2_X1 U103bar ( .A1(n128bar), .A2(n212bar), .ZN(ybar[1]) );
  OR2_X1 U104 ( .A1(n126), .A2(n188), .ZN(n127) );
  AND2_X1 U104bar ( .A1(n126bar), .A2(n188bar), .ZN(n127bar) );
  AND2_X1 U105 ( .A1(n188), .A2(n126), .ZN(n128) );
  OR2_X1 U105bar ( .A1(n188bar), .A2(n126bar), .ZN(n128bar) );
  AND2_X1 U106 ( .A1(n125), .A2(n124), .ZN(n126) );
  OR2_X1 U106bar ( .A1(n125bar), .A2(n124bar), .ZN(n126bar) );
  OR2_X1 U107 ( .A1(n211), .A2(b[1]), .ZN(n124) );
  AND2_X1 U107bar ( .A1(n211bar), .A2(bbar[1]), .ZN(n124bar) );
  OR2_X1 U108 ( .A1(n202), .A2(a[1]), .ZN(n125) );
  AND2_X1 U108bar ( .A1(n202bar), .A2(abar[1]), .ZN(n125bar) );
  AND2_X1 U109 ( .A1(n122), .A2(n121), .ZN(n123) );
  OR2_X1 U109bar ( .A1(n122bar), .A2(n121bar), .ZN(n123bar) );
  OR2_X1 U110 ( .A1(n187), .A2(d[1]), .ZN(n121) );
  AND2_X1 U110bar ( .A1(n187bar), .A2(dbar[1]), .ZN(n121bar) );
  OR2_X1 U111 ( .A1(n178), .A2(c[1]), .ZN(n122) );
  AND2_X1 U111bar ( .A1(n178bar), .A2(cbar[1]), .ZN(n122bar) );
  OR2_X1 U112 ( .A1(n120), .A2(n210), .ZN(y[0]) );
  AND2_X1 U112bar ( .A1(n120bar), .A2(n210bar), .ZN(ybar[0]) );
  OR2_X1 U113 ( .A1(n118), .A2(n186), .ZN(n119) );
  AND2_X1 U113bar ( .A1(n118bar), .A2(n186bar), .ZN(n119bar) );
  AND2_X1 U114 ( .A1(n186), .A2(n118), .ZN(n120) );
  OR2_X1 U114bar ( .A1(n186bar), .A2(n118bar), .ZN(n120bar) );
  AND2_X1 U115 ( .A1(n117), .A2(n116), .ZN(n118) );
  OR2_X1 U115bar ( .A1(n117bar), .A2(n116bar), .ZN(n118bar) );
  OR2_X1 U116 ( .A1(n209), .A2(b[0]), .ZN(n116) );
  AND2_X1 U116bar ( .A1(n209bar), .A2(bbar[0]), .ZN(n116bar) );
  OR2_X1 U117 ( .A1(n201), .A2(a[0]), .ZN(n117) );
  AND2_X1 U117bar ( .A1(n201bar), .A2(abar[0]), .ZN(n117bar) );
  AND2_X1 U118 ( .A1(n114), .A2(n113), .ZN(n115) );
  OR2_X1 U118bar ( .A1(n114bar), .A2(n113bar), .ZN(n115bar) );
  OR2_X1 U119 ( .A1(n185), .A2(d[0]), .ZN(n113) );
  AND2_X1 U119bar ( .A1(n185bar), .A2(dbar[0]), .ZN(n113bar) );
  OR2_X1 U120 ( .A1(n177), .A2(c[0]), .ZN(n114) );
  AND2_X1 U120bar ( .A1(n177bar), .A2(cbar[0]), .ZN(n114bar) );
endmodule

module byteXor4_2 ( a, abar, b, bbar, c, cbar, d, dbar, y, ybar );

  input wire [7:0] a;
  input wire [7:0] b;
  input wire [7:0] c;
  input wire [7:0] d;
  input wire [7:0] abar;
  input wire [7:0] bbar;
  input wire [7:0] cbar;
  input wire [7:0] dbar;
//input_done

  output wire [7:0] y;
  output wire [7:0] ybar;
//output_done

  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n113bar;
  wire n114bar;
  wire n115bar;
  wire n116bar;
  wire n117bar;
  wire n118bar;
  wire n119bar;
  wire n120bar;
  wire n121bar;
  wire n122bar;
  wire n123bar;
  wire n124bar;
  wire n125bar;
  wire n126bar;
  wire n127bar;
  wire n128bar;
  wire n129bar;
  wire n130bar;
  wire n131bar;
  wire n132bar;
  wire n133bar;
  wire n134bar;
  wire n135bar;
  wire n136bar;
  wire n137bar;
  wire n138bar;
  wire n139bar;
  wire n140bar;
  wire n141bar;
  wire n142bar;
  wire n143bar;
  wire n144bar;
  wire n145bar;
  wire n146bar;
  wire n147bar;
  wire n148bar;
  wire n149bar;
  wire n150bar;
  wire n151bar;
  wire n152bar;
  wire n153bar;
  wire n154bar;
  wire n155bar;
  wire n156bar;
  wire n157bar;
  wire n158bar;
  wire n159bar;
  wire n160bar;
  wire n161bar;
  wire n162bar;
  wire n163bar;
  wire n164bar;
  wire n165bar;
  wire n166bar;
  wire n167bar;
  wire n168bar;
  wire n169bar;
  wire n170bar;
  wire n171bar;
  wire n172bar;
  wire n173bar;
  wire n174bar;
  wire n175bar;
  wire n176bar;
  wire n177bar;
  wire n178bar;
  wire n179bar;
  wire n180bar;
  wire n181bar;
  wire n182bar;
  wire n183bar;
  wire n184bar;
  wire n185bar;
  wire n186bar;
  wire n187bar;
  wire n188bar;
  wire n189bar;
  wire n190bar;
  wire n191bar;
  wire n192bar;
  wire n193bar;
  wire n194bar;
  wire n195bar;
  wire n196bar;
  wire n197bar;
  wire n198bar;
  wire n199bar;
  wire n200bar;
  wire n201bar;
  wire n202bar;
  wire n203bar;
  wire n204bar;
  wire n205bar;
  wire n206bar;
  wire n207bar;
  wire n208bar;
  wire n209bar;
  wire n210bar;
  wire n211bar;
  wire n212bar;
  wire n213bar;
  wire n214bar;
  wire n215bar;
  wire n216bar;
  wire n217bar;
  wire n218bar;
  wire n219bar;
  wire n220bar;
  wire n221bar;
  wire n222bar;
  wire n223bar;
  wire n224bar;
//wire_done

 //assign_done

  assign n224bar = n175;
  assign n224 = n175bar;
  assign n223bar = a[7];
  assign n223 = abar[7];
  assign n222bar = n167;
  assign n222 = n167bar;
  assign n221bar = a[6];
  assign n221 = abar[6];
  assign n220bar = n159;
  assign n220 = n159bar;
  assign n219bar = a[5];
  assign n219 = abar[5];
  assign n218bar = n151;
  assign n218 = n151bar;
  assign n217bar = a[4];
  assign n217 = abar[4];
  assign n216bar = n143;
  assign n216 = n143bar;
  assign n215bar = a[3];
  assign n215 = abar[3];
  assign n214bar = n135;
  assign n214 = n135bar;
  assign n213bar = a[2];
  assign n213 = abar[2];
  assign n212bar = n127;
  assign n212 = n127bar;
  assign n211bar = a[1];
  assign n211 = abar[1];
  assign n210bar = n119;
  assign n210 = n119bar;
  assign n209bar = a[0];
  assign n209 = abar[0];
  assign n208bar = b[7];
  assign n208 = bbar[7];
  assign n207bar = b[6];
  assign n207 = bbar[6];
  assign n206bar = b[5];
  assign n206 = bbar[5];
  assign n205bar = b[4];
  assign n205 = bbar[4];
  assign n204bar = b[3];
  assign n204 = bbar[3];
  assign n203bar = b[2];
  assign n203 = bbar[2];
  assign n202bar = b[1];
  assign n202 = bbar[1];
  assign n201bar = b[0];
  assign n201 = bbar[0];
  assign n200bar = n171;
  assign n200 = n171bar;
  assign n199bar = c[7];
  assign n199 = cbar[7];
  assign n198bar = n163;
  assign n198 = n163bar;
  assign n197bar = c[6];
  assign n197 = cbar[6];
  assign n196bar = n155;
  assign n196 = n155bar;
  assign n195bar = c[5];
  assign n195 = cbar[5];
  assign n194bar = n147;
  assign n194 = n147bar;
  assign n193bar = c[4];
  assign n193 = cbar[4];
  assign n192bar = n139;
  assign n192 = n139bar;
  assign n191bar = c[3];
  assign n191 = cbar[3];
  assign n190bar = n131;
  assign n190 = n131bar;
  assign n189bar = c[2];
  assign n189 = cbar[2];
  assign n188bar = n123;
  assign n188 = n123bar;
  assign n187bar = c[1];
  assign n187 = cbar[1];
  assign n186bar = n115;
  assign n186 = n115bar;
  assign n185bar = c[0];
  assign n185 = cbar[0];
  assign n184bar = d[7];
  assign n184 = dbar[7];
  assign n183bar = d[6];
  assign n183 = dbar[6];
  assign n182bar = d[5];
  assign n182 = dbar[5];
  assign n181bar = d[4];
  assign n181 = dbar[4];
  assign n180bar = d[3];
  assign n180 = dbar[3];
  assign n179bar = d[2];
  assign n179 = dbar[2];
  assign n178bar = d[1];
  assign n178 = dbar[1];
  assign n177bar = d[0];
  assign n177 = dbar[0];
  OR2_X1 U49 ( .A1(n176), .A2(n224), .ZN(y[7]) );
  AND2_X1 U49bar ( .A1(n176bar), .A2(n224bar), .ZN(ybar[7]) );
  OR2_X1 U50 ( .A1(n174), .A2(n200), .ZN(n175) );
  AND2_X1 U50bar ( .A1(n174bar), .A2(n200bar), .ZN(n175bar) );
  AND2_X1 U51 ( .A1(n200), .A2(n174), .ZN(n176) );
  OR2_X1 U51bar ( .A1(n200bar), .A2(n174bar), .ZN(n176bar) );
  AND2_X1 U52 ( .A1(n173), .A2(n172), .ZN(n174) );
  OR2_X1 U52bar ( .A1(n173bar), .A2(n172bar), .ZN(n174bar) );
  OR2_X1 U53 ( .A1(n223), .A2(b[7]), .ZN(n172) );
  AND2_X1 U53bar ( .A1(n223bar), .A2(bbar[7]), .ZN(n172bar) );
  OR2_X1 U54 ( .A1(n208), .A2(a[7]), .ZN(n173) );
  AND2_X1 U54bar ( .A1(n208bar), .A2(abar[7]), .ZN(n173bar) );
  AND2_X1 U55 ( .A1(n170), .A2(n169), .ZN(n171) );
  OR2_X1 U55bar ( .A1(n170bar), .A2(n169bar), .ZN(n171bar) );
  OR2_X1 U56 ( .A1(n199), .A2(d[7]), .ZN(n169) );
  AND2_X1 U56bar ( .A1(n199bar), .A2(dbar[7]), .ZN(n169bar) );
  OR2_X1 U57 ( .A1(n184), .A2(c[7]), .ZN(n170) );
  AND2_X1 U57bar ( .A1(n184bar), .A2(cbar[7]), .ZN(n170bar) );
  OR2_X1 U58 ( .A1(n168), .A2(n222), .ZN(y[6]) );
  AND2_X1 U58bar ( .A1(n168bar), .A2(n222bar), .ZN(ybar[6]) );
  OR2_X1 U59 ( .A1(n166), .A2(n198), .ZN(n167) );
  AND2_X1 U59bar ( .A1(n166bar), .A2(n198bar), .ZN(n167bar) );
  AND2_X1 U60 ( .A1(n198), .A2(n166), .ZN(n168) );
  OR2_X1 U60bar ( .A1(n198bar), .A2(n166bar), .ZN(n168bar) );
  AND2_X1 U61 ( .A1(n165), .A2(n164), .ZN(n166) );
  OR2_X1 U61bar ( .A1(n165bar), .A2(n164bar), .ZN(n166bar) );
  OR2_X1 U62 ( .A1(n221), .A2(b[6]), .ZN(n164) );
  AND2_X1 U62bar ( .A1(n221bar), .A2(bbar[6]), .ZN(n164bar) );
  OR2_X1 U63 ( .A1(n207), .A2(a[6]), .ZN(n165) );
  AND2_X1 U63bar ( .A1(n207bar), .A2(abar[6]), .ZN(n165bar) );
  AND2_X1 U64 ( .A1(n162), .A2(n161), .ZN(n163) );
  OR2_X1 U64bar ( .A1(n162bar), .A2(n161bar), .ZN(n163bar) );
  OR2_X1 U65 ( .A1(n197), .A2(d[6]), .ZN(n161) );
  AND2_X1 U65bar ( .A1(n197bar), .A2(dbar[6]), .ZN(n161bar) );
  OR2_X1 U66 ( .A1(n183), .A2(c[6]), .ZN(n162) );
  AND2_X1 U66bar ( .A1(n183bar), .A2(cbar[6]), .ZN(n162bar) );
  OR2_X1 U67 ( .A1(n160), .A2(n220), .ZN(y[5]) );
  AND2_X1 U67bar ( .A1(n160bar), .A2(n220bar), .ZN(ybar[5]) );
  OR2_X1 U68 ( .A1(n158), .A2(n196), .ZN(n159) );
  AND2_X1 U68bar ( .A1(n158bar), .A2(n196bar), .ZN(n159bar) );
  AND2_X1 U69 ( .A1(n196), .A2(n158), .ZN(n160) );
  OR2_X1 U69bar ( .A1(n196bar), .A2(n158bar), .ZN(n160bar) );
  AND2_X1 U70 ( .A1(n157), .A2(n156), .ZN(n158) );
  OR2_X1 U70bar ( .A1(n157bar), .A2(n156bar), .ZN(n158bar) );
  OR2_X1 U71 ( .A1(n219), .A2(b[5]), .ZN(n156) );
  AND2_X1 U71bar ( .A1(n219bar), .A2(bbar[5]), .ZN(n156bar) );
  OR2_X1 U72 ( .A1(n206), .A2(a[5]), .ZN(n157) );
  AND2_X1 U72bar ( .A1(n206bar), .A2(abar[5]), .ZN(n157bar) );
  AND2_X1 U73 ( .A1(n154), .A2(n153), .ZN(n155) );
  OR2_X1 U73bar ( .A1(n154bar), .A2(n153bar), .ZN(n155bar) );
  OR2_X1 U74 ( .A1(n195), .A2(d[5]), .ZN(n153) );
  AND2_X1 U74bar ( .A1(n195bar), .A2(dbar[5]), .ZN(n153bar) );
  OR2_X1 U75 ( .A1(n182), .A2(c[5]), .ZN(n154) );
  AND2_X1 U75bar ( .A1(n182bar), .A2(cbar[5]), .ZN(n154bar) );
  OR2_X1 U76 ( .A1(n152), .A2(n218), .ZN(y[4]) );
  AND2_X1 U76bar ( .A1(n152bar), .A2(n218bar), .ZN(ybar[4]) );
  OR2_X1 U77 ( .A1(n150), .A2(n194), .ZN(n151) );
  AND2_X1 U77bar ( .A1(n150bar), .A2(n194bar), .ZN(n151bar) );
  AND2_X1 U78 ( .A1(n194), .A2(n150), .ZN(n152) );
  OR2_X1 U78bar ( .A1(n194bar), .A2(n150bar), .ZN(n152bar) );
  AND2_X1 U79 ( .A1(n149), .A2(n148), .ZN(n150) );
  OR2_X1 U79bar ( .A1(n149bar), .A2(n148bar), .ZN(n150bar) );
  OR2_X1 U80 ( .A1(n217), .A2(b[4]), .ZN(n148) );
  AND2_X1 U80bar ( .A1(n217bar), .A2(bbar[4]), .ZN(n148bar) );
  OR2_X1 U81 ( .A1(n205), .A2(a[4]), .ZN(n149) );
  AND2_X1 U81bar ( .A1(n205bar), .A2(abar[4]), .ZN(n149bar) );
  AND2_X1 U82 ( .A1(n146), .A2(n145), .ZN(n147) );
  OR2_X1 U82bar ( .A1(n146bar), .A2(n145bar), .ZN(n147bar) );
  OR2_X1 U83 ( .A1(n193), .A2(d[4]), .ZN(n145) );
  AND2_X1 U83bar ( .A1(n193bar), .A2(dbar[4]), .ZN(n145bar) );
  OR2_X1 U84 ( .A1(n181), .A2(c[4]), .ZN(n146) );
  AND2_X1 U84bar ( .A1(n181bar), .A2(cbar[4]), .ZN(n146bar) );
  OR2_X1 U85 ( .A1(n144), .A2(n216), .ZN(y[3]) );
  AND2_X1 U85bar ( .A1(n144bar), .A2(n216bar), .ZN(ybar[3]) );
  OR2_X1 U86 ( .A1(n142), .A2(n192), .ZN(n143) );
  AND2_X1 U86bar ( .A1(n142bar), .A2(n192bar), .ZN(n143bar) );
  AND2_X1 U87 ( .A1(n192), .A2(n142), .ZN(n144) );
  OR2_X1 U87bar ( .A1(n192bar), .A2(n142bar), .ZN(n144bar) );
  AND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(n142) );
  OR2_X1 U88bar ( .A1(n141bar), .A2(n140bar), .ZN(n142bar) );
  OR2_X1 U89 ( .A1(n215), .A2(b[3]), .ZN(n140) );
  AND2_X1 U89bar ( .A1(n215bar), .A2(bbar[3]), .ZN(n140bar) );
  OR2_X1 U90 ( .A1(n204), .A2(a[3]), .ZN(n141) );
  AND2_X1 U90bar ( .A1(n204bar), .A2(abar[3]), .ZN(n141bar) );
  AND2_X1 U91 ( .A1(n138), .A2(n137), .ZN(n139) );
  OR2_X1 U91bar ( .A1(n138bar), .A2(n137bar), .ZN(n139bar) );
  OR2_X1 U92 ( .A1(n191), .A2(d[3]), .ZN(n137) );
  AND2_X1 U92bar ( .A1(n191bar), .A2(dbar[3]), .ZN(n137bar) );
  OR2_X1 U93 ( .A1(n180), .A2(c[3]), .ZN(n138) );
  AND2_X1 U93bar ( .A1(n180bar), .A2(cbar[3]), .ZN(n138bar) );
  OR2_X1 U94 ( .A1(n136), .A2(n214), .ZN(y[2]) );
  AND2_X1 U94bar ( .A1(n136bar), .A2(n214bar), .ZN(ybar[2]) );
  OR2_X1 U95 ( .A1(n134), .A2(n190), .ZN(n135) );
  AND2_X1 U95bar ( .A1(n134bar), .A2(n190bar), .ZN(n135bar) );
  AND2_X1 U96 ( .A1(n190), .A2(n134), .ZN(n136) );
  OR2_X1 U96bar ( .A1(n190bar), .A2(n134bar), .ZN(n136bar) );
  AND2_X1 U97 ( .A1(n133), .A2(n132), .ZN(n134) );
  OR2_X1 U97bar ( .A1(n133bar), .A2(n132bar), .ZN(n134bar) );
  OR2_X1 U98 ( .A1(n213), .A2(b[2]), .ZN(n132) );
  AND2_X1 U98bar ( .A1(n213bar), .A2(bbar[2]), .ZN(n132bar) );
  OR2_X1 U99 ( .A1(n203), .A2(a[2]), .ZN(n133) );
  AND2_X1 U99bar ( .A1(n203bar), .A2(abar[2]), .ZN(n133bar) );
  AND2_X1 U100 ( .A1(n130), .A2(n129), .ZN(n131) );
  OR2_X1 U100bar ( .A1(n130bar), .A2(n129bar), .ZN(n131bar) );
  OR2_X1 U101 ( .A1(n189), .A2(d[2]), .ZN(n129) );
  AND2_X1 U101bar ( .A1(n189bar), .A2(dbar[2]), .ZN(n129bar) );
  OR2_X1 U102 ( .A1(n179), .A2(c[2]), .ZN(n130) );
  AND2_X1 U102bar ( .A1(n179bar), .A2(cbar[2]), .ZN(n130bar) );
  OR2_X1 U103 ( .A1(n128), .A2(n212), .ZN(y[1]) );
  AND2_X1 U103bar ( .A1(n128bar), .A2(n212bar), .ZN(ybar[1]) );
  OR2_X1 U104 ( .A1(n126), .A2(n188), .ZN(n127) );
  AND2_X1 U104bar ( .A1(n126bar), .A2(n188bar), .ZN(n127bar) );
  AND2_X1 U105 ( .A1(n188), .A2(n126), .ZN(n128) );
  OR2_X1 U105bar ( .A1(n188bar), .A2(n126bar), .ZN(n128bar) );
  AND2_X1 U106 ( .A1(n125), .A2(n124), .ZN(n126) );
  OR2_X1 U106bar ( .A1(n125bar), .A2(n124bar), .ZN(n126bar) );
  OR2_X1 U107 ( .A1(n211), .A2(b[1]), .ZN(n124) );
  AND2_X1 U107bar ( .A1(n211bar), .A2(bbar[1]), .ZN(n124bar) );
  OR2_X1 U108 ( .A1(n202), .A2(a[1]), .ZN(n125) );
  AND2_X1 U108bar ( .A1(n202bar), .A2(abar[1]), .ZN(n125bar) );
  AND2_X1 U109 ( .A1(n122), .A2(n121), .ZN(n123) );
  OR2_X1 U109bar ( .A1(n122bar), .A2(n121bar), .ZN(n123bar) );
  OR2_X1 U110 ( .A1(n187), .A2(d[1]), .ZN(n121) );
  AND2_X1 U110bar ( .A1(n187bar), .A2(dbar[1]), .ZN(n121bar) );
  OR2_X1 U111 ( .A1(n178), .A2(c[1]), .ZN(n122) );
  AND2_X1 U111bar ( .A1(n178bar), .A2(cbar[1]), .ZN(n122bar) );
  OR2_X1 U112 ( .A1(n120), .A2(n210), .ZN(y[0]) );
  AND2_X1 U112bar ( .A1(n120bar), .A2(n210bar), .ZN(ybar[0]) );
  OR2_X1 U113 ( .A1(n118), .A2(n186), .ZN(n119) );
  AND2_X1 U113bar ( .A1(n118bar), .A2(n186bar), .ZN(n119bar) );
  AND2_X1 U114 ( .A1(n186), .A2(n118), .ZN(n120) );
  OR2_X1 U114bar ( .A1(n186bar), .A2(n118bar), .ZN(n120bar) );
  AND2_X1 U115 ( .A1(n117), .A2(n116), .ZN(n118) );
  OR2_X1 U115bar ( .A1(n117bar), .A2(n116bar), .ZN(n118bar) );
  OR2_X1 U116 ( .A1(n209), .A2(b[0]), .ZN(n116) );
  AND2_X1 U116bar ( .A1(n209bar), .A2(bbar[0]), .ZN(n116bar) );
  OR2_X1 U117 ( .A1(n201), .A2(a[0]), .ZN(n117) );
  AND2_X1 U117bar ( .A1(n201bar), .A2(abar[0]), .ZN(n117bar) );
  AND2_X1 U118 ( .A1(n114), .A2(n113), .ZN(n115) );
  OR2_X1 U118bar ( .A1(n114bar), .A2(n113bar), .ZN(n115bar) );
  OR2_X1 U119 ( .A1(n185), .A2(d[0]), .ZN(n113) );
  AND2_X1 U119bar ( .A1(n185bar), .A2(dbar[0]), .ZN(n113bar) );
  OR2_X1 U120 ( .A1(n177), .A2(c[0]), .ZN(n114) );
  AND2_X1 U120bar ( .A1(n177bar), .A2(cbar[0]), .ZN(n114bar) );
endmodule

module byteXor4_3 ( a, abar, b, bbar, c, cbar, d, dbar, y, ybar );

  input wire [7:0] a;
  input wire [7:0] b;
  input wire [7:0] c;
  input wire [7:0] d;
  input wire [7:0] abar;
  input wire [7:0] bbar;
  input wire [7:0] cbar;
  input wire [7:0] dbar;
//input_done

  output wire [7:0] y;
  output wire [7:0] ybar;
//output_done

  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n113bar;
  wire n114bar;
  wire n115bar;
  wire n116bar;
  wire n117bar;
  wire n118bar;
  wire n119bar;
  wire n120bar;
  wire n121bar;
  wire n122bar;
  wire n123bar;
  wire n124bar;
  wire n125bar;
  wire n126bar;
  wire n127bar;
  wire n128bar;
  wire n129bar;
  wire n130bar;
  wire n131bar;
  wire n132bar;
  wire n133bar;
  wire n134bar;
  wire n135bar;
  wire n136bar;
  wire n137bar;
  wire n138bar;
  wire n139bar;
  wire n140bar;
  wire n141bar;
  wire n142bar;
  wire n143bar;
  wire n144bar;
  wire n145bar;
  wire n146bar;
  wire n147bar;
  wire n148bar;
  wire n149bar;
  wire n150bar;
  wire n151bar;
  wire n152bar;
  wire n153bar;
  wire n154bar;
  wire n155bar;
  wire n156bar;
  wire n157bar;
  wire n158bar;
  wire n159bar;
  wire n160bar;
  wire n161bar;
  wire n162bar;
  wire n163bar;
  wire n164bar;
  wire n165bar;
  wire n166bar;
  wire n167bar;
  wire n168bar;
  wire n169bar;
  wire n170bar;
  wire n171bar;
  wire n172bar;
  wire n173bar;
  wire n174bar;
  wire n175bar;
  wire n176bar;
  wire n177bar;
  wire n178bar;
  wire n179bar;
  wire n180bar;
  wire n181bar;
  wire n182bar;
  wire n183bar;
  wire n184bar;
  wire n185bar;
  wire n186bar;
  wire n187bar;
  wire n188bar;
  wire n189bar;
  wire n190bar;
  wire n191bar;
  wire n192bar;
  wire n193bar;
  wire n194bar;
  wire n195bar;
  wire n196bar;
  wire n197bar;
  wire n198bar;
  wire n199bar;
  wire n200bar;
  wire n201bar;
  wire n202bar;
  wire n203bar;
  wire n204bar;
  wire n205bar;
  wire n206bar;
  wire n207bar;
  wire n208bar;
  wire n209bar;
  wire n210bar;
  wire n211bar;
  wire n212bar;
  wire n213bar;
  wire n214bar;
  wire n215bar;
  wire n216bar;
  wire n217bar;
  wire n218bar;
  wire n219bar;
  wire n220bar;
  wire n221bar;
  wire n222bar;
  wire n223bar;
  wire n224bar;
//wire_done

 //assign_done

  assign n224bar = n175;
  assign n224 = n175bar;
  assign n223bar = a[7];
  assign n223 = abar[7];
  assign n222bar = n167;
  assign n222 = n167bar;
  assign n221bar = a[6];
  assign n221 = abar[6];
  assign n220bar = n159;
  assign n220 = n159bar;
  assign n219bar = a[5];
  assign n219 = abar[5];
  assign n218bar = n151;
  assign n218 = n151bar;
  assign n217bar = a[4];
  assign n217 = abar[4];
  assign n216bar = n143;
  assign n216 = n143bar;
  assign n215bar = a[3];
  assign n215 = abar[3];
  assign n214bar = n135;
  assign n214 = n135bar;
  assign n213bar = a[2];
  assign n213 = abar[2];
  assign n212bar = n127;
  assign n212 = n127bar;
  assign n211bar = a[1];
  assign n211 = abar[1];
  assign n210bar = n119;
  assign n210 = n119bar;
  assign n209bar = a[0];
  assign n209 = abar[0];
  assign n208bar = b[7];
  assign n208 = bbar[7];
  assign n207bar = b[6];
  assign n207 = bbar[6];
  assign n206bar = b[5];
  assign n206 = bbar[5];
  assign n205bar = b[4];
  assign n205 = bbar[4];
  assign n204bar = b[3];
  assign n204 = bbar[3];
  assign n203bar = b[2];
  assign n203 = bbar[2];
  assign n202bar = b[1];
  assign n202 = bbar[1];
  assign n201bar = b[0];
  assign n201 = bbar[0];
  assign n200bar = n171;
  assign n200 = n171bar;
  assign n199bar = c[7];
  assign n199 = cbar[7];
  assign n198bar = n163;
  assign n198 = n163bar;
  assign n197bar = c[6];
  assign n197 = cbar[6];
  assign n196bar = n155;
  assign n196 = n155bar;
  assign n195bar = c[5];
  assign n195 = cbar[5];
  assign n194bar = n147;
  assign n194 = n147bar;
  assign n193bar = c[4];
  assign n193 = cbar[4];
  assign n192bar = n139;
  assign n192 = n139bar;
  assign n191bar = c[3];
  assign n191 = cbar[3];
  assign n190bar = n131;
  assign n190 = n131bar;
  assign n189bar = c[2];
  assign n189 = cbar[2];
  assign n188bar = n123;
  assign n188 = n123bar;
  assign n187bar = c[1];
  assign n187 = cbar[1];
  assign n186bar = n115;
  assign n186 = n115bar;
  assign n185bar = c[0];
  assign n185 = cbar[0];
  assign n184bar = d[7];
  assign n184 = dbar[7];
  assign n183bar = d[6];
  assign n183 = dbar[6];
  assign n182bar = d[5];
  assign n182 = dbar[5];
  assign n181bar = d[4];
  assign n181 = dbar[4];
  assign n180bar = d[3];
  assign n180 = dbar[3];
  assign n179bar = d[2];
  assign n179 = dbar[2];
  assign n178bar = d[1];
  assign n178 = dbar[1];
  assign n177bar = d[0];
  assign n177 = dbar[0];
  OR2_X1 U49 ( .A1(n176), .A2(n224), .ZN(y[7]) );
  AND2_X1 U49bar ( .A1(n176bar), .A2(n224bar), .ZN(ybar[7]) );
  OR2_X1 U50 ( .A1(n174), .A2(n200), .ZN(n175) );
  AND2_X1 U50bar ( .A1(n174bar), .A2(n200bar), .ZN(n175bar) );
  AND2_X1 U51 ( .A1(n200), .A2(n174), .ZN(n176) );
  OR2_X1 U51bar ( .A1(n200bar), .A2(n174bar), .ZN(n176bar) );
  AND2_X1 U52 ( .A1(n173), .A2(n172), .ZN(n174) );
  OR2_X1 U52bar ( .A1(n173bar), .A2(n172bar), .ZN(n174bar) );
  OR2_X1 U53 ( .A1(n223), .A2(b[7]), .ZN(n172) );
  AND2_X1 U53bar ( .A1(n223bar), .A2(bbar[7]), .ZN(n172bar) );
  OR2_X1 U54 ( .A1(n208), .A2(a[7]), .ZN(n173) );
  AND2_X1 U54bar ( .A1(n208bar), .A2(abar[7]), .ZN(n173bar) );
  AND2_X1 U55 ( .A1(n170), .A2(n169), .ZN(n171) );
  OR2_X1 U55bar ( .A1(n170bar), .A2(n169bar), .ZN(n171bar) );
  OR2_X1 U56 ( .A1(n199), .A2(d[7]), .ZN(n169) );
  AND2_X1 U56bar ( .A1(n199bar), .A2(dbar[7]), .ZN(n169bar) );
  OR2_X1 U57 ( .A1(n184), .A2(c[7]), .ZN(n170) );
  AND2_X1 U57bar ( .A1(n184bar), .A2(cbar[7]), .ZN(n170bar) );
  OR2_X1 U58 ( .A1(n168), .A2(n222), .ZN(y[6]) );
  AND2_X1 U58bar ( .A1(n168bar), .A2(n222bar), .ZN(ybar[6]) );
  OR2_X1 U59 ( .A1(n166), .A2(n198), .ZN(n167) );
  AND2_X1 U59bar ( .A1(n166bar), .A2(n198bar), .ZN(n167bar) );
  AND2_X1 U60 ( .A1(n198), .A2(n166), .ZN(n168) );
  OR2_X1 U60bar ( .A1(n198bar), .A2(n166bar), .ZN(n168bar) );
  AND2_X1 U61 ( .A1(n165), .A2(n164), .ZN(n166) );
  OR2_X1 U61bar ( .A1(n165bar), .A2(n164bar), .ZN(n166bar) );
  OR2_X1 U62 ( .A1(n221), .A2(b[6]), .ZN(n164) );
  AND2_X1 U62bar ( .A1(n221bar), .A2(bbar[6]), .ZN(n164bar) );
  OR2_X1 U63 ( .A1(n207), .A2(a[6]), .ZN(n165) );
  AND2_X1 U63bar ( .A1(n207bar), .A2(abar[6]), .ZN(n165bar) );
  AND2_X1 U64 ( .A1(n162), .A2(n161), .ZN(n163) );
  OR2_X1 U64bar ( .A1(n162bar), .A2(n161bar), .ZN(n163bar) );
  OR2_X1 U65 ( .A1(n197), .A2(d[6]), .ZN(n161) );
  AND2_X1 U65bar ( .A1(n197bar), .A2(dbar[6]), .ZN(n161bar) );
  OR2_X1 U66 ( .A1(n183), .A2(c[6]), .ZN(n162) );
  AND2_X1 U66bar ( .A1(n183bar), .A2(cbar[6]), .ZN(n162bar) );
  OR2_X1 U67 ( .A1(n160), .A2(n220), .ZN(y[5]) );
  AND2_X1 U67bar ( .A1(n160bar), .A2(n220bar), .ZN(ybar[5]) );
  OR2_X1 U68 ( .A1(n158), .A2(n196), .ZN(n159) );
  AND2_X1 U68bar ( .A1(n158bar), .A2(n196bar), .ZN(n159bar) );
  AND2_X1 U69 ( .A1(n196), .A2(n158), .ZN(n160) );
  OR2_X1 U69bar ( .A1(n196bar), .A2(n158bar), .ZN(n160bar) );
  AND2_X1 U70 ( .A1(n157), .A2(n156), .ZN(n158) );
  OR2_X1 U70bar ( .A1(n157bar), .A2(n156bar), .ZN(n158bar) );
  OR2_X1 U71 ( .A1(n219), .A2(b[5]), .ZN(n156) );
  AND2_X1 U71bar ( .A1(n219bar), .A2(bbar[5]), .ZN(n156bar) );
  OR2_X1 U72 ( .A1(n206), .A2(a[5]), .ZN(n157) );
  AND2_X1 U72bar ( .A1(n206bar), .A2(abar[5]), .ZN(n157bar) );
  AND2_X1 U73 ( .A1(n154), .A2(n153), .ZN(n155) );
  OR2_X1 U73bar ( .A1(n154bar), .A2(n153bar), .ZN(n155bar) );
  OR2_X1 U74 ( .A1(n195), .A2(d[5]), .ZN(n153) );
  AND2_X1 U74bar ( .A1(n195bar), .A2(dbar[5]), .ZN(n153bar) );
  OR2_X1 U75 ( .A1(n182), .A2(c[5]), .ZN(n154) );
  AND2_X1 U75bar ( .A1(n182bar), .A2(cbar[5]), .ZN(n154bar) );
  OR2_X1 U76 ( .A1(n152), .A2(n218), .ZN(y[4]) );
  AND2_X1 U76bar ( .A1(n152bar), .A2(n218bar), .ZN(ybar[4]) );
  OR2_X1 U77 ( .A1(n150), .A2(n194), .ZN(n151) );
  AND2_X1 U77bar ( .A1(n150bar), .A2(n194bar), .ZN(n151bar) );
  AND2_X1 U78 ( .A1(n194), .A2(n150), .ZN(n152) );
  OR2_X1 U78bar ( .A1(n194bar), .A2(n150bar), .ZN(n152bar) );
  AND2_X1 U79 ( .A1(n149), .A2(n148), .ZN(n150) );
  OR2_X1 U79bar ( .A1(n149bar), .A2(n148bar), .ZN(n150bar) );
  OR2_X1 U80 ( .A1(n217), .A2(b[4]), .ZN(n148) );
  AND2_X1 U80bar ( .A1(n217bar), .A2(bbar[4]), .ZN(n148bar) );
  OR2_X1 U81 ( .A1(n205), .A2(a[4]), .ZN(n149) );
  AND2_X1 U81bar ( .A1(n205bar), .A2(abar[4]), .ZN(n149bar) );
  AND2_X1 U82 ( .A1(n146), .A2(n145), .ZN(n147) );
  OR2_X1 U82bar ( .A1(n146bar), .A2(n145bar), .ZN(n147bar) );
  OR2_X1 U83 ( .A1(n193), .A2(d[4]), .ZN(n145) );
  AND2_X1 U83bar ( .A1(n193bar), .A2(dbar[4]), .ZN(n145bar) );
  OR2_X1 U84 ( .A1(n181), .A2(c[4]), .ZN(n146) );
  AND2_X1 U84bar ( .A1(n181bar), .A2(cbar[4]), .ZN(n146bar) );
  OR2_X1 U85 ( .A1(n144), .A2(n216), .ZN(y[3]) );
  AND2_X1 U85bar ( .A1(n144bar), .A2(n216bar), .ZN(ybar[3]) );
  OR2_X1 U86 ( .A1(n142), .A2(n192), .ZN(n143) );
  AND2_X1 U86bar ( .A1(n142bar), .A2(n192bar), .ZN(n143bar) );
  AND2_X1 U87 ( .A1(n192), .A2(n142), .ZN(n144) );
  OR2_X1 U87bar ( .A1(n192bar), .A2(n142bar), .ZN(n144bar) );
  AND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(n142) );
  OR2_X1 U88bar ( .A1(n141bar), .A2(n140bar), .ZN(n142bar) );
  OR2_X1 U89 ( .A1(n215), .A2(b[3]), .ZN(n140) );
  AND2_X1 U89bar ( .A1(n215bar), .A2(bbar[3]), .ZN(n140bar) );
  OR2_X1 U90 ( .A1(n204), .A2(a[3]), .ZN(n141) );
  AND2_X1 U90bar ( .A1(n204bar), .A2(abar[3]), .ZN(n141bar) );
  AND2_X1 U91 ( .A1(n138), .A2(n137), .ZN(n139) );
  OR2_X1 U91bar ( .A1(n138bar), .A2(n137bar), .ZN(n139bar) );
  OR2_X1 U92 ( .A1(n191), .A2(d[3]), .ZN(n137) );
  AND2_X1 U92bar ( .A1(n191bar), .A2(dbar[3]), .ZN(n137bar) );
  OR2_X1 U93 ( .A1(n180), .A2(c[3]), .ZN(n138) );
  AND2_X1 U93bar ( .A1(n180bar), .A2(cbar[3]), .ZN(n138bar) );
  OR2_X1 U94 ( .A1(n136), .A2(n214), .ZN(y[2]) );
  AND2_X1 U94bar ( .A1(n136bar), .A2(n214bar), .ZN(ybar[2]) );
  OR2_X1 U95 ( .A1(n134), .A2(n190), .ZN(n135) );
  AND2_X1 U95bar ( .A1(n134bar), .A2(n190bar), .ZN(n135bar) );
  AND2_X1 U96 ( .A1(n190), .A2(n134), .ZN(n136) );
  OR2_X1 U96bar ( .A1(n190bar), .A2(n134bar), .ZN(n136bar) );
  AND2_X1 U97 ( .A1(n133), .A2(n132), .ZN(n134) );
  OR2_X1 U97bar ( .A1(n133bar), .A2(n132bar), .ZN(n134bar) );
  OR2_X1 U98 ( .A1(n213), .A2(b[2]), .ZN(n132) );
  AND2_X1 U98bar ( .A1(n213bar), .A2(bbar[2]), .ZN(n132bar) );
  OR2_X1 U99 ( .A1(n203), .A2(a[2]), .ZN(n133) );
  AND2_X1 U99bar ( .A1(n203bar), .A2(abar[2]), .ZN(n133bar) );
  AND2_X1 U100 ( .A1(n130), .A2(n129), .ZN(n131) );
  OR2_X1 U100bar ( .A1(n130bar), .A2(n129bar), .ZN(n131bar) );
  OR2_X1 U101 ( .A1(n189), .A2(d[2]), .ZN(n129) );
  AND2_X1 U101bar ( .A1(n189bar), .A2(dbar[2]), .ZN(n129bar) );
  OR2_X1 U102 ( .A1(n179), .A2(c[2]), .ZN(n130) );
  AND2_X1 U102bar ( .A1(n179bar), .A2(cbar[2]), .ZN(n130bar) );
  OR2_X1 U103 ( .A1(n128), .A2(n212), .ZN(y[1]) );
  AND2_X1 U103bar ( .A1(n128bar), .A2(n212bar), .ZN(ybar[1]) );
  OR2_X1 U104 ( .A1(n126), .A2(n188), .ZN(n127) );
  AND2_X1 U104bar ( .A1(n126bar), .A2(n188bar), .ZN(n127bar) );
  AND2_X1 U105 ( .A1(n188), .A2(n126), .ZN(n128) );
  OR2_X1 U105bar ( .A1(n188bar), .A2(n126bar), .ZN(n128bar) );
  AND2_X1 U106 ( .A1(n125), .A2(n124), .ZN(n126) );
  OR2_X1 U106bar ( .A1(n125bar), .A2(n124bar), .ZN(n126bar) );
  OR2_X1 U107 ( .A1(n211), .A2(b[1]), .ZN(n124) );
  AND2_X1 U107bar ( .A1(n211bar), .A2(bbar[1]), .ZN(n124bar) );
  OR2_X1 U108 ( .A1(n202), .A2(a[1]), .ZN(n125) );
  AND2_X1 U108bar ( .A1(n202bar), .A2(abar[1]), .ZN(n125bar) );
  AND2_X1 U109 ( .A1(n122), .A2(n121), .ZN(n123) );
  OR2_X1 U109bar ( .A1(n122bar), .A2(n121bar), .ZN(n123bar) );
  OR2_X1 U110 ( .A1(n187), .A2(d[1]), .ZN(n121) );
  AND2_X1 U110bar ( .A1(n187bar), .A2(dbar[1]), .ZN(n121bar) );
  OR2_X1 U111 ( .A1(n178), .A2(c[1]), .ZN(n122) );
  AND2_X1 U111bar ( .A1(n178bar), .A2(cbar[1]), .ZN(n122bar) );
  OR2_X1 U112 ( .A1(n120), .A2(n210), .ZN(y[0]) );
  AND2_X1 U112bar ( .A1(n120bar), .A2(n210bar), .ZN(ybar[0]) );
  OR2_X1 U113 ( .A1(n118), .A2(n186), .ZN(n119) );
  AND2_X1 U113bar ( .A1(n118bar), .A2(n186bar), .ZN(n119bar) );
  AND2_X1 U114 ( .A1(n186), .A2(n118), .ZN(n120) );
  OR2_X1 U114bar ( .A1(n186bar), .A2(n118bar), .ZN(n120bar) );
  AND2_X1 U115 ( .A1(n117), .A2(n116), .ZN(n118) );
  OR2_X1 U115bar ( .A1(n117bar), .A2(n116bar), .ZN(n118bar) );
  OR2_X1 U116 ( .A1(n209), .A2(b[0]), .ZN(n116) );
  AND2_X1 U116bar ( .A1(n209bar), .A2(bbar[0]), .ZN(n116bar) );
  OR2_X1 U117 ( .A1(n201), .A2(a[0]), .ZN(n117) );
  AND2_X1 U117bar ( .A1(n201bar), .A2(abar[0]), .ZN(n117bar) );
  AND2_X1 U118 ( .A1(n114), .A2(n113), .ZN(n115) );
  OR2_X1 U118bar ( .A1(n114bar), .A2(n113bar), .ZN(n115bar) );
  OR2_X1 U119 ( .A1(n185), .A2(d[0]), .ZN(n113) );
  AND2_X1 U119bar ( .A1(n185bar), .A2(dbar[0]), .ZN(n113bar) );
  OR2_X1 U120 ( .A1(n177), .A2(c[0]), .ZN(n114) );
  AND2_X1 U120bar ( .A1(n177bar), .A2(cbar[0]), .ZN(n114bar) );
endmodule

module byteXor4_4 ( a, abar, b, bbar, c, cbar, d, dbar, y, ybar );

  input wire [7:0] a;
  input wire [7:0] b;
  input wire [7:0] c;
  input wire [7:0] d;
  input wire [7:0] abar;
  input wire [7:0] bbar;
  input wire [7:0] cbar;
  input wire [7:0] dbar;
//input_done

  output wire [7:0] y;
  output wire [7:0] ybar;
//output_done

  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n113bar;
  wire n114bar;
  wire n115bar;
  wire n116bar;
  wire n117bar;
  wire n118bar;
  wire n119bar;
  wire n120bar;
  wire n121bar;
  wire n122bar;
  wire n123bar;
  wire n124bar;
  wire n125bar;
  wire n126bar;
  wire n127bar;
  wire n128bar;
  wire n129bar;
  wire n130bar;
  wire n131bar;
  wire n132bar;
  wire n133bar;
  wire n134bar;
  wire n135bar;
  wire n136bar;
  wire n137bar;
  wire n138bar;
  wire n139bar;
  wire n140bar;
  wire n141bar;
  wire n142bar;
  wire n143bar;
  wire n144bar;
  wire n145bar;
  wire n146bar;
  wire n147bar;
  wire n148bar;
  wire n149bar;
  wire n150bar;
  wire n151bar;
  wire n152bar;
  wire n153bar;
  wire n154bar;
  wire n155bar;
  wire n156bar;
  wire n157bar;
  wire n158bar;
  wire n159bar;
  wire n160bar;
  wire n161bar;
  wire n162bar;
  wire n163bar;
  wire n164bar;
  wire n165bar;
  wire n166bar;
  wire n167bar;
  wire n168bar;
  wire n169bar;
  wire n170bar;
  wire n171bar;
  wire n172bar;
  wire n173bar;
  wire n174bar;
  wire n175bar;
  wire n176bar;
  wire n177bar;
  wire n178bar;
  wire n179bar;
  wire n180bar;
  wire n181bar;
  wire n182bar;
  wire n183bar;
  wire n184bar;
  wire n185bar;
  wire n186bar;
  wire n187bar;
  wire n188bar;
  wire n189bar;
  wire n190bar;
  wire n191bar;
  wire n192bar;
  wire n193bar;
  wire n194bar;
  wire n195bar;
  wire n196bar;
  wire n197bar;
  wire n198bar;
  wire n199bar;
  wire n200bar;
  wire n201bar;
  wire n202bar;
  wire n203bar;
  wire n204bar;
  wire n205bar;
  wire n206bar;
  wire n207bar;
  wire n208bar;
  wire n209bar;
  wire n210bar;
  wire n211bar;
  wire n212bar;
  wire n213bar;
  wire n214bar;
  wire n215bar;
  wire n216bar;
  wire n217bar;
  wire n218bar;
  wire n219bar;
  wire n220bar;
  wire n221bar;
  wire n222bar;
  wire n223bar;
  wire n224bar;
//wire_done

 //assign_done

  assign n224bar = n175;
  assign n224 = n175bar;
  assign n223bar = a[7];
  assign n223 = abar[7];
  assign n222bar = n167;
  assign n222 = n167bar;
  assign n221bar = a[6];
  assign n221 = abar[6];
  assign n220bar = n159;
  assign n220 = n159bar;
  assign n219bar = a[5];
  assign n219 = abar[5];
  assign n218bar = n151;
  assign n218 = n151bar;
  assign n217bar = a[4];
  assign n217 = abar[4];
  assign n216bar = n143;
  assign n216 = n143bar;
  assign n215bar = a[3];
  assign n215 = abar[3];
  assign n214bar = n135;
  assign n214 = n135bar;
  assign n213bar = a[2];
  assign n213 = abar[2];
  assign n212bar = n127;
  assign n212 = n127bar;
  assign n211bar = a[1];
  assign n211 = abar[1];
  assign n210bar = n119;
  assign n210 = n119bar;
  assign n209bar = a[0];
  assign n209 = abar[0];
  assign n208bar = b[7];
  assign n208 = bbar[7];
  assign n207bar = b[6];
  assign n207 = bbar[6];
  assign n206bar = b[5];
  assign n206 = bbar[5];
  assign n205bar = b[4];
  assign n205 = bbar[4];
  assign n204bar = b[3];
  assign n204 = bbar[3];
  assign n203bar = b[2];
  assign n203 = bbar[2];
  assign n202bar = b[1];
  assign n202 = bbar[1];
  assign n201bar = b[0];
  assign n201 = bbar[0];
  assign n200bar = n171;
  assign n200 = n171bar;
  assign n199bar = c[7];
  assign n199 = cbar[7];
  assign n198bar = n163;
  assign n198 = n163bar;
  assign n197bar = c[6];
  assign n197 = cbar[6];
  assign n196bar = n155;
  assign n196 = n155bar;
  assign n195bar = c[5];
  assign n195 = cbar[5];
  assign n194bar = n147;
  assign n194 = n147bar;
  assign n193bar = c[4];
  assign n193 = cbar[4];
  assign n192bar = n139;
  assign n192 = n139bar;
  assign n191bar = c[3];
  assign n191 = cbar[3];
  assign n190bar = n131;
  assign n190 = n131bar;
  assign n189bar = c[2];
  assign n189 = cbar[2];
  assign n188bar = n123;
  assign n188 = n123bar;
  assign n187bar = c[1];
  assign n187 = cbar[1];
  assign n186bar = n115;
  assign n186 = n115bar;
  assign n185bar = c[0];
  assign n185 = cbar[0];
  assign n184bar = d[7];
  assign n184 = dbar[7];
  assign n183bar = d[6];
  assign n183 = dbar[6];
  assign n182bar = d[5];
  assign n182 = dbar[5];
  assign n181bar = d[4];
  assign n181 = dbar[4];
  assign n180bar = d[3];
  assign n180 = dbar[3];
  assign n179bar = d[2];
  assign n179 = dbar[2];
  assign n178bar = d[1];
  assign n178 = dbar[1];
  assign n177bar = d[0];
  assign n177 = dbar[0];
  OR2_X1 U49 ( .A1(n176), .A2(n224), .ZN(y[7]) );
  AND2_X1 U49bar ( .A1(n176bar), .A2(n224bar), .ZN(ybar[7]) );
  OR2_X1 U50 ( .A1(n174), .A2(n200), .ZN(n175) );
  AND2_X1 U50bar ( .A1(n174bar), .A2(n200bar), .ZN(n175bar) );
  AND2_X1 U51 ( .A1(n200), .A2(n174), .ZN(n176) );
  OR2_X1 U51bar ( .A1(n200bar), .A2(n174bar), .ZN(n176bar) );
  AND2_X1 U52 ( .A1(n173), .A2(n172), .ZN(n174) );
  OR2_X1 U52bar ( .A1(n173bar), .A2(n172bar), .ZN(n174bar) );
  OR2_X1 U53 ( .A1(n223), .A2(b[7]), .ZN(n172) );
  AND2_X1 U53bar ( .A1(n223bar), .A2(bbar[7]), .ZN(n172bar) );
  OR2_X1 U54 ( .A1(n208), .A2(a[7]), .ZN(n173) );
  AND2_X1 U54bar ( .A1(n208bar), .A2(abar[7]), .ZN(n173bar) );
  AND2_X1 U55 ( .A1(n170), .A2(n169), .ZN(n171) );
  OR2_X1 U55bar ( .A1(n170bar), .A2(n169bar), .ZN(n171bar) );
  OR2_X1 U56 ( .A1(n199), .A2(d[7]), .ZN(n169) );
  AND2_X1 U56bar ( .A1(n199bar), .A2(dbar[7]), .ZN(n169bar) );
  OR2_X1 U57 ( .A1(n184), .A2(c[7]), .ZN(n170) );
  AND2_X1 U57bar ( .A1(n184bar), .A2(cbar[7]), .ZN(n170bar) );
  OR2_X1 U58 ( .A1(n168), .A2(n222), .ZN(y[6]) );
  AND2_X1 U58bar ( .A1(n168bar), .A2(n222bar), .ZN(ybar[6]) );
  OR2_X1 U59 ( .A1(n166), .A2(n198), .ZN(n167) );
  AND2_X1 U59bar ( .A1(n166bar), .A2(n198bar), .ZN(n167bar) );
  AND2_X1 U60 ( .A1(n198), .A2(n166), .ZN(n168) );
  OR2_X1 U60bar ( .A1(n198bar), .A2(n166bar), .ZN(n168bar) );
  AND2_X1 U61 ( .A1(n165), .A2(n164), .ZN(n166) );
  OR2_X1 U61bar ( .A1(n165bar), .A2(n164bar), .ZN(n166bar) );
  OR2_X1 U62 ( .A1(n221), .A2(b[6]), .ZN(n164) );
  AND2_X1 U62bar ( .A1(n221bar), .A2(bbar[6]), .ZN(n164bar) );
  OR2_X1 U63 ( .A1(n207), .A2(a[6]), .ZN(n165) );
  AND2_X1 U63bar ( .A1(n207bar), .A2(abar[6]), .ZN(n165bar) );
  AND2_X1 U64 ( .A1(n162), .A2(n161), .ZN(n163) );
  OR2_X1 U64bar ( .A1(n162bar), .A2(n161bar), .ZN(n163bar) );
  OR2_X1 U65 ( .A1(n197), .A2(d[6]), .ZN(n161) );
  AND2_X1 U65bar ( .A1(n197bar), .A2(dbar[6]), .ZN(n161bar) );
  OR2_X1 U66 ( .A1(n183), .A2(c[6]), .ZN(n162) );
  AND2_X1 U66bar ( .A1(n183bar), .A2(cbar[6]), .ZN(n162bar) );
  OR2_X1 U67 ( .A1(n160), .A2(n220), .ZN(y[5]) );
  AND2_X1 U67bar ( .A1(n160bar), .A2(n220bar), .ZN(ybar[5]) );
  OR2_X1 U68 ( .A1(n158), .A2(n196), .ZN(n159) );
  AND2_X1 U68bar ( .A1(n158bar), .A2(n196bar), .ZN(n159bar) );
  AND2_X1 U69 ( .A1(n196), .A2(n158), .ZN(n160) );
  OR2_X1 U69bar ( .A1(n196bar), .A2(n158bar), .ZN(n160bar) );
  AND2_X1 U70 ( .A1(n157), .A2(n156), .ZN(n158) );
  OR2_X1 U70bar ( .A1(n157bar), .A2(n156bar), .ZN(n158bar) );
  OR2_X1 U71 ( .A1(n219), .A2(b[5]), .ZN(n156) );
  AND2_X1 U71bar ( .A1(n219bar), .A2(bbar[5]), .ZN(n156bar) );
  OR2_X1 U72 ( .A1(n206), .A2(a[5]), .ZN(n157) );
  AND2_X1 U72bar ( .A1(n206bar), .A2(abar[5]), .ZN(n157bar) );
  AND2_X1 U73 ( .A1(n154), .A2(n153), .ZN(n155) );
  OR2_X1 U73bar ( .A1(n154bar), .A2(n153bar), .ZN(n155bar) );
  OR2_X1 U74 ( .A1(n195), .A2(d[5]), .ZN(n153) );
  AND2_X1 U74bar ( .A1(n195bar), .A2(dbar[5]), .ZN(n153bar) );
  OR2_X1 U75 ( .A1(n182), .A2(c[5]), .ZN(n154) );
  AND2_X1 U75bar ( .A1(n182bar), .A2(cbar[5]), .ZN(n154bar) );
  OR2_X1 U76 ( .A1(n152), .A2(n218), .ZN(y[4]) );
  AND2_X1 U76bar ( .A1(n152bar), .A2(n218bar), .ZN(ybar[4]) );
  OR2_X1 U77 ( .A1(n150), .A2(n194), .ZN(n151) );
  AND2_X1 U77bar ( .A1(n150bar), .A2(n194bar), .ZN(n151bar) );
  AND2_X1 U78 ( .A1(n194), .A2(n150), .ZN(n152) );
  OR2_X1 U78bar ( .A1(n194bar), .A2(n150bar), .ZN(n152bar) );
  AND2_X1 U79 ( .A1(n149), .A2(n148), .ZN(n150) );
  OR2_X1 U79bar ( .A1(n149bar), .A2(n148bar), .ZN(n150bar) );
  OR2_X1 U80 ( .A1(n217), .A2(b[4]), .ZN(n148) );
  AND2_X1 U80bar ( .A1(n217bar), .A2(bbar[4]), .ZN(n148bar) );
  OR2_X1 U81 ( .A1(n205), .A2(a[4]), .ZN(n149) );
  AND2_X1 U81bar ( .A1(n205bar), .A2(abar[4]), .ZN(n149bar) );
  AND2_X1 U82 ( .A1(n146), .A2(n145), .ZN(n147) );
  OR2_X1 U82bar ( .A1(n146bar), .A2(n145bar), .ZN(n147bar) );
  OR2_X1 U83 ( .A1(n193), .A2(d[4]), .ZN(n145) );
  AND2_X1 U83bar ( .A1(n193bar), .A2(dbar[4]), .ZN(n145bar) );
  OR2_X1 U84 ( .A1(n181), .A2(c[4]), .ZN(n146) );
  AND2_X1 U84bar ( .A1(n181bar), .A2(cbar[4]), .ZN(n146bar) );
  OR2_X1 U85 ( .A1(n144), .A2(n216), .ZN(y[3]) );
  AND2_X1 U85bar ( .A1(n144bar), .A2(n216bar), .ZN(ybar[3]) );
  OR2_X1 U86 ( .A1(n142), .A2(n192), .ZN(n143) );
  AND2_X1 U86bar ( .A1(n142bar), .A2(n192bar), .ZN(n143bar) );
  AND2_X1 U87 ( .A1(n192), .A2(n142), .ZN(n144) );
  OR2_X1 U87bar ( .A1(n192bar), .A2(n142bar), .ZN(n144bar) );
  AND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(n142) );
  OR2_X1 U88bar ( .A1(n141bar), .A2(n140bar), .ZN(n142bar) );
  OR2_X1 U89 ( .A1(n215), .A2(b[3]), .ZN(n140) );
  AND2_X1 U89bar ( .A1(n215bar), .A2(bbar[3]), .ZN(n140bar) );
  OR2_X1 U90 ( .A1(n204), .A2(a[3]), .ZN(n141) );
  AND2_X1 U90bar ( .A1(n204bar), .A2(abar[3]), .ZN(n141bar) );
  AND2_X1 U91 ( .A1(n138), .A2(n137), .ZN(n139) );
  OR2_X1 U91bar ( .A1(n138bar), .A2(n137bar), .ZN(n139bar) );
  OR2_X1 U92 ( .A1(n191), .A2(d[3]), .ZN(n137) );
  AND2_X1 U92bar ( .A1(n191bar), .A2(dbar[3]), .ZN(n137bar) );
  OR2_X1 U93 ( .A1(n180), .A2(c[3]), .ZN(n138) );
  AND2_X1 U93bar ( .A1(n180bar), .A2(cbar[3]), .ZN(n138bar) );
  OR2_X1 U94 ( .A1(n136), .A2(n214), .ZN(y[2]) );
  AND2_X1 U94bar ( .A1(n136bar), .A2(n214bar), .ZN(ybar[2]) );
  OR2_X1 U95 ( .A1(n134), .A2(n190), .ZN(n135) );
  AND2_X1 U95bar ( .A1(n134bar), .A2(n190bar), .ZN(n135bar) );
  AND2_X1 U96 ( .A1(n190), .A2(n134), .ZN(n136) );
  OR2_X1 U96bar ( .A1(n190bar), .A2(n134bar), .ZN(n136bar) );
  AND2_X1 U97 ( .A1(n133), .A2(n132), .ZN(n134) );
  OR2_X1 U97bar ( .A1(n133bar), .A2(n132bar), .ZN(n134bar) );
  OR2_X1 U98 ( .A1(n213), .A2(b[2]), .ZN(n132) );
  AND2_X1 U98bar ( .A1(n213bar), .A2(bbar[2]), .ZN(n132bar) );
  OR2_X1 U99 ( .A1(n203), .A2(a[2]), .ZN(n133) );
  AND2_X1 U99bar ( .A1(n203bar), .A2(abar[2]), .ZN(n133bar) );
  AND2_X1 U100 ( .A1(n130), .A2(n129), .ZN(n131) );
  OR2_X1 U100bar ( .A1(n130bar), .A2(n129bar), .ZN(n131bar) );
  OR2_X1 U101 ( .A1(n189), .A2(d[2]), .ZN(n129) );
  AND2_X1 U101bar ( .A1(n189bar), .A2(dbar[2]), .ZN(n129bar) );
  OR2_X1 U102 ( .A1(n179), .A2(c[2]), .ZN(n130) );
  AND2_X1 U102bar ( .A1(n179bar), .A2(cbar[2]), .ZN(n130bar) );
  OR2_X1 U103 ( .A1(n128), .A2(n212), .ZN(y[1]) );
  AND2_X1 U103bar ( .A1(n128bar), .A2(n212bar), .ZN(ybar[1]) );
  OR2_X1 U104 ( .A1(n126), .A2(n188), .ZN(n127) );
  AND2_X1 U104bar ( .A1(n126bar), .A2(n188bar), .ZN(n127bar) );
  AND2_X1 U105 ( .A1(n188), .A2(n126), .ZN(n128) );
  OR2_X1 U105bar ( .A1(n188bar), .A2(n126bar), .ZN(n128bar) );
  AND2_X1 U106 ( .A1(n125), .A2(n124), .ZN(n126) );
  OR2_X1 U106bar ( .A1(n125bar), .A2(n124bar), .ZN(n126bar) );
  OR2_X1 U107 ( .A1(n211), .A2(b[1]), .ZN(n124) );
  AND2_X1 U107bar ( .A1(n211bar), .A2(bbar[1]), .ZN(n124bar) );
  OR2_X1 U108 ( .A1(n202), .A2(a[1]), .ZN(n125) );
  AND2_X1 U108bar ( .A1(n202bar), .A2(abar[1]), .ZN(n125bar) );
  AND2_X1 U109 ( .A1(n122), .A2(n121), .ZN(n123) );
  OR2_X1 U109bar ( .A1(n122bar), .A2(n121bar), .ZN(n123bar) );
  OR2_X1 U110 ( .A1(n187), .A2(d[1]), .ZN(n121) );
  AND2_X1 U110bar ( .A1(n187bar), .A2(dbar[1]), .ZN(n121bar) );
  OR2_X1 U111 ( .A1(n178), .A2(c[1]), .ZN(n122) );
  AND2_X1 U111bar ( .A1(n178bar), .A2(cbar[1]), .ZN(n122bar) );
  OR2_X1 U112 ( .A1(n120), .A2(n210), .ZN(y[0]) );
  AND2_X1 U112bar ( .A1(n120bar), .A2(n210bar), .ZN(ybar[0]) );
  OR2_X1 U113 ( .A1(n118), .A2(n186), .ZN(n119) );
  AND2_X1 U113bar ( .A1(n118bar), .A2(n186bar), .ZN(n119bar) );
  AND2_X1 U114 ( .A1(n186), .A2(n118), .ZN(n120) );
  OR2_X1 U114bar ( .A1(n186bar), .A2(n118bar), .ZN(n120bar) );
  AND2_X1 U115 ( .A1(n117), .A2(n116), .ZN(n118) );
  OR2_X1 U115bar ( .A1(n117bar), .A2(n116bar), .ZN(n118bar) );
  OR2_X1 U116 ( .A1(n209), .A2(b[0]), .ZN(n116) );
  AND2_X1 U116bar ( .A1(n209bar), .A2(bbar[0]), .ZN(n116bar) );
  OR2_X1 U117 ( .A1(n201), .A2(a[0]), .ZN(n117) );
  AND2_X1 U117bar ( .A1(n201bar), .A2(abar[0]), .ZN(n117bar) );
  AND2_X1 U118 ( .A1(n114), .A2(n113), .ZN(n115) );
  OR2_X1 U118bar ( .A1(n114bar), .A2(n113bar), .ZN(n115bar) );
  OR2_X1 U119 ( .A1(n185), .A2(d[0]), .ZN(n113) );
  AND2_X1 U119bar ( .A1(n185bar), .A2(dbar[0]), .ZN(n113bar) );
  OR2_X1 U120 ( .A1(n177), .A2(c[0]), .ZN(n114) );
  AND2_X1 U120bar ( .A1(n177bar), .A2(cbar[0]), .ZN(n114bar) );
endmodule

module mixCol_1 ( in, inbar, out, outbar );

  input wire [31:0] in;
  input wire [31:0] inbar;
//input_done

  output wire [31:0] out;
  output wire [31:0] outbar;
//output_done

  wire [7:0] b0_s2;
  wire [7:0] b1_s2;
  wire [7:0] b2_s2;
  wire [7:0] b3_s2;
  wire [7:0] b0_s3;
  wire [7:0] b1_s3;
  wire [7:0] b2_s3;
  wire [7:0] b3_s3;

  wire [7:0] b0_s2bar;
  wire [7:0] b1_s2bar;
  wire [7:0] b2_s2bar;
  wire [7:0] b3_s2bar;
  wire [7:0] b0_s3bar;
  wire [7:0] b1_s3bar;
  wire [7:0] b2_s3bar;
  wire [7:0] b3_s3bar;
//wire_done

 //assign_done

  scale2_4 b0_scale2 ( .in(in[31:24]), .inbar(inbar[31:24]), .out(b0_s2), .outbar(b0_s2bar) );
  scale2_3 b1_scale2 ( .in(in[23:16]), .inbar(inbar[23:16]), .out(b1_s2), .outbar(b1_s2bar) );
  scale2_2 b2_scale2 ( .in(in[15:8]), .inbar(inbar[15:8]), .out(b2_s2), .outbar(b2_s2bar) );
  scale2_1 b3_scale2 ( .in(in[7:0]), .inbar(inbar[7:0]), .out(b3_s2), .outbar(b3_s2bar) );

  byteXor_5 b0_scale3 ( .a(in[31:24]), .abar(inbar[31:24]), .b(b0_s2), .bbar(b0_s2bar), .y(b0_s3), .ybar(b0_s3bar) );
  byteXor_4 b1_scale3 ( .a(in[23:16]), .abar(inbar[23:16]), .b(b1_s2), .bbar(b1_s2bar), .y(b1_s3), .ybar(b1_s3bar) );
  byteXor_3 b2_scale3 ( .a(in[15:8]), .abar(inbar[15:8]), .b(b2_s2), .bbar(b2_s2bar), .y(b2_s3), .ybar(b2_s3bar) );
  byteXor_2 b3_scale3 ( .a(in[7:0]), .abar(inbar[7:0]), .b(b3_s2), .bbar(b3_s2bar), .y(b3_s3), .ybar(b3_s3bar) );

  byteXor4_4 out0 ( .a(b0_s2), .abar(b0_s2bar), .b(b1_s3), .bbar(b1_s3bar), .c(in[15:8]), .cbar(inbar[15:8]),
       .d(in[7:0]), .dbar(inbar[7:0]), .y(out[31:24]), .ybar(outbar[31:24]) );
  byteXor4_3 out1 ( .a(in[31:24]), .abar(inbar[31:24]), .b(b1_s2), .bbar(b1_s2bar), .c(b2_s3), .cbar(b2_s3bar),
       .d(in[7:0]), .dbar(inbar[7:0]), .y(out[23:16]), .ybar(outbar[23:16]) );
  byteXor4_2 out2 ( .a(in[31:24]), .abar(inbar[31:24]), .b(in[23:16]), .bbar(inbar[23:16]), .c(b2_s2), .cbar(b2_s2bar),
       .d(b3_s3), .dbar(b3_s3bar), .y(out[15:8]), .ybar(outbar[15:8]) );
  byteXor4_1 out3 ( .a(b0_s3), .abar(b0_s3bar), .b(in[23:16]), .bbar(inbar[23:16]), .c(in[15:8]), .cbar(inbar[15:8]),
       .d(b3_s2), .dbar(b3_s2bar), .y(out[7:0]), .ybar(outbar[7:0]) );
endmodule

module scale2_5 ( in, inbar, out, outbar );

  input wire [7:0] in;
  input wire [7:0] inbar;
//input_done

  output wire [7:0] out;
  output wire [7:0] outbar;
//output_done

  wire in_0;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_1;
  wire in_7;
  wire n11;
  wire n12;
  wire n13;
  wire n14;
  wire n15;
  wire n16;
  wire n17;
  wire n18;
  wire n19;
  wire n20;
  wire in_0bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_1bar;
  wire in_7bar;
  wire n11bar;
  wire n12bar;
  wire n13bar;
  wire n14bar;
  wire n15bar;
  wire n16bar;
  wire n17bar;
  wire n18bar;
  wire n19bar;
  wire n20bar;
//wire_done

  assign in_0 = in[0];
  assign out[7] = in_6;
  assign in_6  = in[6];
  assign out[6] = in_5;
  assign in_5  = in[5];
  assign out[5] = in_4;
  assign in_4  = in[4];
  assign out[2] = in_1;
  assign in_1  = in[1];
  assign out[0] = in_7;
  assign in_7  = in[7];
  assign in_0bar = inbar[0];
  assign outbar[7] = in_6bar;
  assign in_6bar = inbar[6];
  assign outbar[6] = in_5bar;
  assign in_5bar = inbar[5];
  assign outbar[5] = in_4bar;
  assign in_4bar = inbar[4];
  assign outbar[2] = in_1bar;
  assign in_1bar = inbar[1];
  assign outbar[0] = in_7bar;
  assign in_7bar = inbar[7];
//assign_done

  assign n20bar = in_7;
  assign n20 = in_7bar;
  assign n19bar = in[3];
  assign n19 = inbar[3];
  assign n18bar = in[2];
  assign n18 = inbar[2];
  assign n17bar = in_0;
  assign n17 = in_0bar;
  OR2_X1 U5 ( .A1(n16), .A2(n15), .ZN(out[4]) );
  AND2_X1 U5bar ( .A1(n16bar), .A2(n15bar), .ZN(outbar[4]) );
  AND2_X1 U6 ( .A1(in[3]), .A2(n20), .ZN(n15) );
  OR2_X1 U6bar ( .A1(inbar[3]), .A2(n20bar), .ZN(n15bar) );
  AND2_X1 U7 ( .A1(in_7), .A2(n19), .ZN(n16) );
  OR2_X1 U7bar ( .A1(in_7bar), .A2(n19bar), .ZN(n16bar) );
  OR2_X1 U8 ( .A1(n14), .A2(n13), .ZN(out[3]) );
  AND2_X1 U8bar ( .A1(n14bar), .A2(n13bar), .ZN(outbar[3]) );
  AND2_X1 U9 ( .A1(in[2]), .A2(n20), .ZN(n13) );
  OR2_X1 U9bar ( .A1(inbar[2]), .A2(n20bar), .ZN(n13bar) );
  AND2_X1 U10 ( .A1(in_7), .A2(n18), .ZN(n14) );
  OR2_X1 U10bar ( .A1(in_7bar), .A2(n18bar), .ZN(n14bar) );
  OR2_X1 U11 ( .A1(n12), .A2(n11), .ZN(out[1]) );
  AND2_X1 U11bar ( .A1(n12bar), .A2(n11bar), .ZN(outbar[1]) );
  AND2_X1 U12 ( .A1(in_0), .A2(n20), .ZN(n11) );
  OR2_X1 U12bar ( .A1(in_0bar), .A2(n20bar), .ZN(n11bar) );
  AND2_X1 U13 ( .A1(in_7), .A2(n17), .ZN(n12) );
  OR2_X1 U13bar ( .A1(in_7bar), .A2(n17bar), .ZN(n12bar) );
endmodule

module scale2_6 ( in, inbar, out, outbar );

  input wire [7:0] in;
  input wire [7:0] inbar;
//input_done

  output wire [7:0] out;
  output wire [7:0] outbar;
//output_done

  wire in_0;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_1;
  wire in_7;
  wire n11;
  wire n12;
  wire n13;
  wire n14;
  wire n15;
  wire n16;
  wire n17;
  wire n18;
  wire n19;
  wire n20;
  wire in_0bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_1bar;
  wire in_7bar;
  wire n11bar;
  wire n12bar;
  wire n13bar;
  wire n14bar;
  wire n15bar;
  wire n16bar;
  wire n17bar;
  wire n18bar;
  wire n19bar;
  wire n20bar;
//wire_done

  assign in_0 = in[0];
  assign out[7] = in_6;
  assign in_6  = in[6];
  assign out[6] = in_5;
  assign in_5  = in[5];
  assign out[5] = in_4;
  assign in_4  = in[4];
  assign out[2] = in_1;
  assign in_1  = in[1];
  assign out[0] = in_7;
  assign in_7  = in[7];
  assign in_0bar = inbar[0];
  assign outbar[7] = in_6bar;
  assign in_6bar = inbar[6];
  assign outbar[6] = in_5bar;
  assign in_5bar = inbar[5];
  assign outbar[5] = in_4bar;
  assign in_4bar = inbar[4];
  assign outbar[2] = in_1bar;
  assign in_1bar = inbar[1];
  assign outbar[0] = in_7bar;
  assign in_7bar = inbar[7];
//assign_done

  assign n20bar = in_7;
  assign n20 = in_7bar;
  assign n19bar = in[3];
  assign n19 = inbar[3];
  assign n18bar = in[2];
  assign n18 = inbar[2];
  assign n17bar = in_0;
  assign n17 = in_0bar;
  OR2_X1 U5 ( .A1(n16), .A2(n15), .ZN(out[4]) );
  AND2_X1 U5bar ( .A1(n16bar), .A2(n15bar), .ZN(outbar[4]) );
  AND2_X1 U6 ( .A1(in[3]), .A2(n20), .ZN(n15) );
  OR2_X1 U6bar ( .A1(inbar[3]), .A2(n20bar), .ZN(n15bar) );
  AND2_X1 U7 ( .A1(in_7), .A2(n19), .ZN(n16) );
  OR2_X1 U7bar ( .A1(in_7bar), .A2(n19bar), .ZN(n16bar) );
  OR2_X1 U8 ( .A1(n14), .A2(n13), .ZN(out[3]) );
  AND2_X1 U8bar ( .A1(n14bar), .A2(n13bar), .ZN(outbar[3]) );
  AND2_X1 U9 ( .A1(in[2]), .A2(n20), .ZN(n13) );
  OR2_X1 U9bar ( .A1(inbar[2]), .A2(n20bar), .ZN(n13bar) );
  AND2_X1 U10 ( .A1(in_7), .A2(n18), .ZN(n14) );
  OR2_X1 U10bar ( .A1(in_7bar), .A2(n18bar), .ZN(n14bar) );
  OR2_X1 U11 ( .A1(n12), .A2(n11), .ZN(out[1]) );
  AND2_X1 U11bar ( .A1(n12bar), .A2(n11bar), .ZN(outbar[1]) );
  AND2_X1 U12 ( .A1(in_0), .A2(n20), .ZN(n11) );
  OR2_X1 U12bar ( .A1(in_0bar), .A2(n20bar), .ZN(n11bar) );
  AND2_X1 U13 ( .A1(in_7), .A2(n17), .ZN(n12) );
  OR2_X1 U13bar ( .A1(in_7bar), .A2(n17bar), .ZN(n12bar) );
endmodule

module scale2_7 ( in, inbar, out, outbar );

  input wire [7:0] in;
  input wire [7:0] inbar;
//input_done

  output wire [7:0] out;
  output wire [7:0] outbar;
//output_done

  wire in_0;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_1;
  wire in_7;
  wire n11;
  wire n12;
  wire n13;
  wire n14;
  wire n15;
  wire n16;
  wire n17;
  wire n18;
  wire n19;
  wire n20;
  wire in_0bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_1bar;
  wire in_7bar;
  wire n11bar;
  wire n12bar;
  wire n13bar;
  wire n14bar;
  wire n15bar;
  wire n16bar;
  wire n17bar;
  wire n18bar;
  wire n19bar;
  wire n20bar;
//wire_done

  assign in_0 = in[0];
  assign out[7] = in_6;
  assign in_6  = in[6];
  assign out[6] = in_5;
  assign in_5  = in[5];
  assign out[5] = in_4;
  assign in_4  = in[4];
  assign out[2] = in_1;
  assign in_1  = in[1];
  assign out[0] = in_7;
  assign in_7  = in[7];
  assign in_0bar = inbar[0];
  assign outbar[7] = in_6bar;
  assign in_6bar = inbar[6];
  assign outbar[6] = in_5bar;
  assign in_5bar = inbar[5];
  assign outbar[5] = in_4bar;
  assign in_4bar = inbar[4];
  assign outbar[2] = in_1bar;
  assign in_1bar = inbar[1];
  assign outbar[0] = in_7bar;
  assign in_7bar = inbar[7];
//assign_done

  assign n20bar = in_7;
  assign n20 = in_7bar;
  assign n19bar = in[3];
  assign n19 = inbar[3];
  assign n18bar = in[2];
  assign n18 = inbar[2];
  assign n17bar = in_0;
  assign n17 = in_0bar;
  OR2_X1 U5 ( .A1(n16), .A2(n15), .ZN(out[4]) );
  AND2_X1 U5bar ( .A1(n16bar), .A2(n15bar), .ZN(outbar[4]) );
  AND2_X1 U6 ( .A1(in[3]), .A2(n20), .ZN(n15) );
  OR2_X1 U6bar ( .A1(inbar[3]), .A2(n20bar), .ZN(n15bar) );
  AND2_X1 U7 ( .A1(in_7), .A2(n19), .ZN(n16) );
  OR2_X1 U7bar ( .A1(in_7bar), .A2(n19bar), .ZN(n16bar) );
  OR2_X1 U8 ( .A1(n14), .A2(n13), .ZN(out[3]) );
  AND2_X1 U8bar ( .A1(n14bar), .A2(n13bar), .ZN(outbar[3]) );
  AND2_X1 U9 ( .A1(in[2]), .A2(n20), .ZN(n13) );
  OR2_X1 U9bar ( .A1(inbar[2]), .A2(n20bar), .ZN(n13bar) );
  AND2_X1 U10 ( .A1(in_7), .A2(n18), .ZN(n14) );
  OR2_X1 U10bar ( .A1(in_7bar), .A2(n18bar), .ZN(n14bar) );
  OR2_X1 U11 ( .A1(n12), .A2(n11), .ZN(out[1]) );
  AND2_X1 U11bar ( .A1(n12bar), .A2(n11bar), .ZN(outbar[1]) );
  AND2_X1 U12 ( .A1(in_0), .A2(n20), .ZN(n11) );
  OR2_X1 U12bar ( .A1(in_0bar), .A2(n20bar), .ZN(n11bar) );
  AND2_X1 U13 ( .A1(in_7), .A2(n17), .ZN(n12) );
  OR2_X1 U13bar ( .A1(in_7bar), .A2(n17bar), .ZN(n12bar) );
endmodule

module scale2_8 ( in, inbar, out, outbar );

  input wire [7:0] in;
  input wire [7:0] inbar;
//input_done

  output wire [7:0] out;
  output wire [7:0] outbar;
//output_done

  wire in_0;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_1;
  wire in_7;
  wire n11;
  wire n12;
  wire n13;
  wire n14;
  wire n15;
  wire n16;
  wire n17;
  wire n18;
  wire n19;
  wire n20;
  wire in_0bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_1bar;
  wire in_7bar;
  wire n11bar;
  wire n12bar;
  wire n13bar;
  wire n14bar;
  wire n15bar;
  wire n16bar;
  wire n17bar;
  wire n18bar;
  wire n19bar;
  wire n20bar;
//wire_done

  assign in_0 = in[0];
  assign out[7] = in_6;
  assign in_6  = in[6];
  assign out[6] = in_5;
  assign in_5  = in[5];
  assign out[5] = in_4;
  assign in_4  = in[4];
  assign out[2] = in_1;
  assign in_1  = in[1];
  assign out[0] = in_7;
  assign in_7  = in[7];
  assign in_0bar = inbar[0];
  assign outbar[7] = in_6bar;
  assign in_6bar = inbar[6];
  assign outbar[6] = in_5bar;
  assign in_5bar = inbar[5];
  assign outbar[5] = in_4bar;
  assign in_4bar = inbar[4];
  assign outbar[2] = in_1bar;
  assign in_1bar = inbar[1];
  assign outbar[0] = in_7bar;
  assign in_7bar = inbar[7];
//assign_done

  assign n20bar = in_7;
  assign n20 = in_7bar;
  assign n19bar = in[3];
  assign n19 = inbar[3];
  assign n18bar = in[2];
  assign n18 = inbar[2];
  assign n17bar = in_0;
  assign n17 = in_0bar;
  OR2_X1 U5 ( .A1(n16), .A2(n15), .ZN(out[4]) );
  AND2_X1 U5bar ( .A1(n16bar), .A2(n15bar), .ZN(outbar[4]) );
  AND2_X1 U6 ( .A1(in[3]), .A2(n20), .ZN(n15) );
  OR2_X1 U6bar ( .A1(inbar[3]), .A2(n20bar), .ZN(n15bar) );
  AND2_X1 U7 ( .A1(in_7), .A2(n19), .ZN(n16) );
  OR2_X1 U7bar ( .A1(in_7bar), .A2(n19bar), .ZN(n16bar) );
  OR2_X1 U8 ( .A1(n14), .A2(n13), .ZN(out[3]) );
  AND2_X1 U8bar ( .A1(n14bar), .A2(n13bar), .ZN(outbar[3]) );
  AND2_X1 U9 ( .A1(in[2]), .A2(n20), .ZN(n13) );
  OR2_X1 U9bar ( .A1(inbar[2]), .A2(n20bar), .ZN(n13bar) );
  AND2_X1 U10 ( .A1(in_7), .A2(n18), .ZN(n14) );
  OR2_X1 U10bar ( .A1(in_7bar), .A2(n18bar), .ZN(n14bar) );
  OR2_X1 U11 ( .A1(n12), .A2(n11), .ZN(out[1]) );
  AND2_X1 U11bar ( .A1(n12bar), .A2(n11bar), .ZN(outbar[1]) );
  AND2_X1 U12 ( .A1(in_0), .A2(n20), .ZN(n11) );
  OR2_X1 U12bar ( .A1(in_0bar), .A2(n20bar), .ZN(n11bar) );
  AND2_X1 U13 ( .A1(in_7), .A2(n17), .ZN(n12) );
  OR2_X1 U13bar ( .A1(in_7bar), .A2(n17bar), .ZN(n12bar) );
endmodule

module byteXor_6 ( a, abar, b, bbar, y, ybar );

  input wire [7:0] a;
  input wire [7:0] b;
  input wire [7:0] abar;
  input wire [7:0] bbar;
//input_done

  output wire [7:0] y;
  output wire [7:0] ybar;
//output_done

  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n33bar;
  wire n34bar;
  wire n35bar;
  wire n36bar;
  wire n37bar;
  wire n38bar;
  wire n39bar;
  wire n40bar;
  wire n41bar;
  wire n42bar;
  wire n43bar;
  wire n44bar;
  wire n45bar;
  wire n46bar;
  wire n47bar;
  wire n48bar;
  wire n49bar;
  wire n50bar;
  wire n51bar;
  wire n52bar;
  wire n53bar;
  wire n54bar;
  wire n55bar;
  wire n56bar;
  wire n57bar;
  wire n58bar;
  wire n59bar;
  wire n60bar;
  wire n61bar;
  wire n62bar;
  wire n63bar;
  wire n64bar;
//wire_done

 //assign_done

  assign n64bar = n47;
  assign n64 = n47bar;
  assign n63bar = a[7];
  assign n63 = abar[7];
  assign n62bar = n45;
  assign n62 = n45bar;
  assign n61bar = a[6];
  assign n61 = abar[6];
  assign n60bar = n43;
  assign n60 = n43bar;
  assign n59bar = a[5];
  assign n59 = abar[5];
  assign n58bar = n41;
  assign n58 = n41bar;
  assign n57bar = a[4];
  assign n57 = abar[4];
  assign n56bar = n39;
  assign n56 = n39bar;
  assign n55bar = a[3];
  assign n55 = abar[3];
  assign n54bar = n37;
  assign n54 = n37bar;
  assign n53bar = a[2];
  assign n53 = abar[2];
  assign n52bar = n35;
  assign n52 = n35bar;
  assign n51bar = a[1];
  assign n51 = abar[1];
  assign n50bar = n33;
  assign n50 = n33bar;
  assign n49bar = a[0];
  assign n49 = abar[0];
  OR2_X1 U17 ( .A1(n48), .A2(n64), .ZN(y[7]) );
  AND2_X1 U17bar ( .A1(n48bar), .A2(n64bar), .ZN(ybar[7]) );
  OR2_X1 U18 ( .A1(n63), .A2(b[7]), .ZN(n47) );
  AND2_X1 U18bar ( .A1(n63bar), .A2(bbar[7]), .ZN(n47bar) );
  AND2_X1 U19 ( .A1(b[7]), .A2(n63), .ZN(n48) );
  OR2_X1 U19bar ( .A1(bbar[7]), .A2(n63bar), .ZN(n48bar) );
  OR2_X1 U20 ( .A1(n46), .A2(n62), .ZN(y[6]) );
  AND2_X1 U20bar ( .A1(n46bar), .A2(n62bar), .ZN(ybar[6]) );
  OR2_X1 U21 ( .A1(n61), .A2(b[6]), .ZN(n45) );
  AND2_X1 U21bar ( .A1(n61bar), .A2(bbar[6]), .ZN(n45bar) );
  AND2_X1 U22 ( .A1(b[6]), .A2(n61), .ZN(n46) );
  OR2_X1 U22bar ( .A1(bbar[6]), .A2(n61bar), .ZN(n46bar) );
  OR2_X1 U23 ( .A1(n44), .A2(n60), .ZN(y[5]) );
  AND2_X1 U23bar ( .A1(n44bar), .A2(n60bar), .ZN(ybar[5]) );
  OR2_X1 U24 ( .A1(n59), .A2(b[5]), .ZN(n43) );
  AND2_X1 U24bar ( .A1(n59bar), .A2(bbar[5]), .ZN(n43bar) );
  AND2_X1 U25 ( .A1(b[5]), .A2(n59), .ZN(n44) );
  OR2_X1 U25bar ( .A1(bbar[5]), .A2(n59bar), .ZN(n44bar) );
  OR2_X1 U26 ( .A1(n42), .A2(n58), .ZN(y[4]) );
  AND2_X1 U26bar ( .A1(n42bar), .A2(n58bar), .ZN(ybar[4]) );
  OR2_X1 U27 ( .A1(n57), .A2(b[4]), .ZN(n41) );
  AND2_X1 U27bar ( .A1(n57bar), .A2(bbar[4]), .ZN(n41bar) );
  AND2_X1 U28 ( .A1(b[4]), .A2(n57), .ZN(n42) );
  OR2_X1 U28bar ( .A1(bbar[4]), .A2(n57bar), .ZN(n42bar) );
  OR2_X1 U29 ( .A1(n40), .A2(n56), .ZN(y[3]) );
  AND2_X1 U29bar ( .A1(n40bar), .A2(n56bar), .ZN(ybar[3]) );
  OR2_X1 U30 ( .A1(n55), .A2(b[3]), .ZN(n39) );
  AND2_X1 U30bar ( .A1(n55bar), .A2(bbar[3]), .ZN(n39bar) );
  AND2_X1 U31 ( .A1(b[3]), .A2(n55), .ZN(n40) );
  OR2_X1 U31bar ( .A1(bbar[3]), .A2(n55bar), .ZN(n40bar) );
  OR2_X1 U32 ( .A1(n38), .A2(n54), .ZN(y[2]) );
  AND2_X1 U32bar ( .A1(n38bar), .A2(n54bar), .ZN(ybar[2]) );
  OR2_X1 U33 ( .A1(n53), .A2(b[2]), .ZN(n37) );
  AND2_X1 U33bar ( .A1(n53bar), .A2(bbar[2]), .ZN(n37bar) );
  AND2_X1 U34 ( .A1(b[2]), .A2(n53), .ZN(n38) );
  OR2_X1 U34bar ( .A1(bbar[2]), .A2(n53bar), .ZN(n38bar) );
  OR2_X1 U35 ( .A1(n36), .A2(n52), .ZN(y[1]) );
  AND2_X1 U35bar ( .A1(n36bar), .A2(n52bar), .ZN(ybar[1]) );
  OR2_X1 U36 ( .A1(n51), .A2(b[1]), .ZN(n35) );
  AND2_X1 U36bar ( .A1(n51bar), .A2(bbar[1]), .ZN(n35bar) );
  AND2_X1 U37 ( .A1(b[1]), .A2(n51), .ZN(n36) );
  OR2_X1 U37bar ( .A1(bbar[1]), .A2(n51bar), .ZN(n36bar) );
  OR2_X1 U38 ( .A1(n34), .A2(n50), .ZN(y[0]) );
  AND2_X1 U38bar ( .A1(n34bar), .A2(n50bar), .ZN(ybar[0]) );
  OR2_X1 U39 ( .A1(n49), .A2(b[0]), .ZN(n33) );
  AND2_X1 U39bar ( .A1(n49bar), .A2(bbar[0]), .ZN(n33bar) );
  AND2_X1 U40 ( .A1(b[0]), .A2(n49), .ZN(n34) );
  OR2_X1 U40bar ( .A1(bbar[0]), .A2(n49bar), .ZN(n34bar) );
endmodule

module byteXor_7 ( a, abar, b, bbar, y, ybar );

  input wire [7:0] a;
  input wire [7:0] b;
  input wire [7:0] abar;
  input wire [7:0] bbar;
//input_done

  output wire [7:0] y;
  output wire [7:0] ybar;
//output_done

  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n33bar;
  wire n34bar;
  wire n35bar;
  wire n36bar;
  wire n37bar;
  wire n38bar;
  wire n39bar;
  wire n40bar;
  wire n41bar;
  wire n42bar;
  wire n43bar;
  wire n44bar;
  wire n45bar;
  wire n46bar;
  wire n47bar;
  wire n48bar;
  wire n49bar;
  wire n50bar;
  wire n51bar;
  wire n52bar;
  wire n53bar;
  wire n54bar;
  wire n55bar;
  wire n56bar;
  wire n57bar;
  wire n58bar;
  wire n59bar;
  wire n60bar;
  wire n61bar;
  wire n62bar;
  wire n63bar;
  wire n64bar;
//wire_done

 //assign_done

  assign n64bar = n47;
  assign n64 = n47bar;
  assign n63bar = a[7];
  assign n63 = abar[7];
  assign n62bar = n45;
  assign n62 = n45bar;
  assign n61bar = a[6];
  assign n61 = abar[6];
  assign n60bar = n43;
  assign n60 = n43bar;
  assign n59bar = a[5];
  assign n59 = abar[5];
  assign n58bar = n41;
  assign n58 = n41bar;
  assign n57bar = a[4];
  assign n57 = abar[4];
  assign n56bar = n39;
  assign n56 = n39bar;
  assign n55bar = a[3];
  assign n55 = abar[3];
  assign n54bar = n37;
  assign n54 = n37bar;
  assign n53bar = a[2];
  assign n53 = abar[2];
  assign n52bar = n35;
  assign n52 = n35bar;
  assign n51bar = a[1];
  assign n51 = abar[1];
  assign n50bar = n33;
  assign n50 = n33bar;
  assign n49bar = a[0];
  assign n49 = abar[0];
  OR2_X1 U17 ( .A1(n48), .A2(n64), .ZN(y[7]) );
  AND2_X1 U17bar ( .A1(n48bar), .A2(n64bar), .ZN(ybar[7]) );
  OR2_X1 U18 ( .A1(n63), .A2(b[7]), .ZN(n47) );
  AND2_X1 U18bar ( .A1(n63bar), .A2(bbar[7]), .ZN(n47bar) );
  AND2_X1 U19 ( .A1(b[7]), .A2(n63), .ZN(n48) );
  OR2_X1 U19bar ( .A1(bbar[7]), .A2(n63bar), .ZN(n48bar) );
  OR2_X1 U20 ( .A1(n46), .A2(n62), .ZN(y[6]) );
  AND2_X1 U20bar ( .A1(n46bar), .A2(n62bar), .ZN(ybar[6]) );
  OR2_X1 U21 ( .A1(n61), .A2(b[6]), .ZN(n45) );
  AND2_X1 U21bar ( .A1(n61bar), .A2(bbar[6]), .ZN(n45bar) );
  AND2_X1 U22 ( .A1(b[6]), .A2(n61), .ZN(n46) );
  OR2_X1 U22bar ( .A1(bbar[6]), .A2(n61bar), .ZN(n46bar) );
  OR2_X1 U23 ( .A1(n44), .A2(n60), .ZN(y[5]) );
  AND2_X1 U23bar ( .A1(n44bar), .A2(n60bar), .ZN(ybar[5]) );
  OR2_X1 U24 ( .A1(n59), .A2(b[5]), .ZN(n43) );
  AND2_X1 U24bar ( .A1(n59bar), .A2(bbar[5]), .ZN(n43bar) );
  AND2_X1 U25 ( .A1(b[5]), .A2(n59), .ZN(n44) );
  OR2_X1 U25bar ( .A1(bbar[5]), .A2(n59bar), .ZN(n44bar) );
  OR2_X1 U26 ( .A1(n42), .A2(n58), .ZN(y[4]) );
  AND2_X1 U26bar ( .A1(n42bar), .A2(n58bar), .ZN(ybar[4]) );
  OR2_X1 U27 ( .A1(n57), .A2(b[4]), .ZN(n41) );
  AND2_X1 U27bar ( .A1(n57bar), .A2(bbar[4]), .ZN(n41bar) );
  AND2_X1 U28 ( .A1(b[4]), .A2(n57), .ZN(n42) );
  OR2_X1 U28bar ( .A1(bbar[4]), .A2(n57bar), .ZN(n42bar) );
  OR2_X1 U29 ( .A1(n40), .A2(n56), .ZN(y[3]) );
  AND2_X1 U29bar ( .A1(n40bar), .A2(n56bar), .ZN(ybar[3]) );
  OR2_X1 U30 ( .A1(n55), .A2(b[3]), .ZN(n39) );
  AND2_X1 U30bar ( .A1(n55bar), .A2(bbar[3]), .ZN(n39bar) );
  AND2_X1 U31 ( .A1(b[3]), .A2(n55), .ZN(n40) );
  OR2_X1 U31bar ( .A1(bbar[3]), .A2(n55bar), .ZN(n40bar) );
  OR2_X1 U32 ( .A1(n38), .A2(n54), .ZN(y[2]) );
  AND2_X1 U32bar ( .A1(n38bar), .A2(n54bar), .ZN(ybar[2]) );
  OR2_X1 U33 ( .A1(n53), .A2(b[2]), .ZN(n37) );
  AND2_X1 U33bar ( .A1(n53bar), .A2(bbar[2]), .ZN(n37bar) );
  AND2_X1 U34 ( .A1(b[2]), .A2(n53), .ZN(n38) );
  OR2_X1 U34bar ( .A1(bbar[2]), .A2(n53bar), .ZN(n38bar) );
  OR2_X1 U35 ( .A1(n36), .A2(n52), .ZN(y[1]) );
  AND2_X1 U35bar ( .A1(n36bar), .A2(n52bar), .ZN(ybar[1]) );
  OR2_X1 U36 ( .A1(n51), .A2(b[1]), .ZN(n35) );
  AND2_X1 U36bar ( .A1(n51bar), .A2(bbar[1]), .ZN(n35bar) );
  AND2_X1 U37 ( .A1(b[1]), .A2(n51), .ZN(n36) );
  OR2_X1 U37bar ( .A1(bbar[1]), .A2(n51bar), .ZN(n36bar) );
  OR2_X1 U38 ( .A1(n34), .A2(n50), .ZN(y[0]) );
  AND2_X1 U38bar ( .A1(n34bar), .A2(n50bar), .ZN(ybar[0]) );
  OR2_X1 U39 ( .A1(n49), .A2(b[0]), .ZN(n33) );
  AND2_X1 U39bar ( .A1(n49bar), .A2(bbar[0]), .ZN(n33bar) );
  AND2_X1 U40 ( .A1(b[0]), .A2(n49), .ZN(n34) );
  OR2_X1 U40bar ( .A1(bbar[0]), .A2(n49bar), .ZN(n34bar) );
endmodule

module byteXor_8 ( a, abar, b, bbar, y, ybar );

  input wire [7:0] a;
  input wire [7:0] b;
  input wire [7:0] abar;
  input wire [7:0] bbar;
//input_done

  output wire [7:0] y;
  output wire [7:0] ybar;
//output_done

  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n33bar;
  wire n34bar;
  wire n35bar;
  wire n36bar;
  wire n37bar;
  wire n38bar;
  wire n39bar;
  wire n40bar;
  wire n41bar;
  wire n42bar;
  wire n43bar;
  wire n44bar;
  wire n45bar;
  wire n46bar;
  wire n47bar;
  wire n48bar;
  wire n49bar;
  wire n50bar;
  wire n51bar;
  wire n52bar;
  wire n53bar;
  wire n54bar;
  wire n55bar;
  wire n56bar;
  wire n57bar;
  wire n58bar;
  wire n59bar;
  wire n60bar;
  wire n61bar;
  wire n62bar;
  wire n63bar;
  wire n64bar;
//wire_done

 //assign_done

  assign n64bar = n47;
  assign n64 = n47bar;
  assign n63bar = a[7];
  assign n63 = abar[7];
  assign n62bar = n45;
  assign n62 = n45bar;
  assign n61bar = a[6];
  assign n61 = abar[6];
  assign n60bar = n43;
  assign n60 = n43bar;
  assign n59bar = a[5];
  assign n59 = abar[5];
  assign n58bar = n41;
  assign n58 = n41bar;
  assign n57bar = a[4];
  assign n57 = abar[4];
  assign n56bar = n39;
  assign n56 = n39bar;
  assign n55bar = a[3];
  assign n55 = abar[3];
  assign n54bar = n37;
  assign n54 = n37bar;
  assign n53bar = a[2];
  assign n53 = abar[2];
  assign n52bar = n35;
  assign n52 = n35bar;
  assign n51bar = a[1];
  assign n51 = abar[1];
  assign n50bar = n33;
  assign n50 = n33bar;
  assign n49bar = a[0];
  assign n49 = abar[0];
  OR2_X1 U17 ( .A1(n48), .A2(n64), .ZN(y[7]) );
  AND2_X1 U17bar ( .A1(n48bar), .A2(n64bar), .ZN(ybar[7]) );
  OR2_X1 U18 ( .A1(n63), .A2(b[7]), .ZN(n47) );
  AND2_X1 U18bar ( .A1(n63bar), .A2(bbar[7]), .ZN(n47bar) );
  AND2_X1 U19 ( .A1(b[7]), .A2(n63), .ZN(n48) );
  OR2_X1 U19bar ( .A1(bbar[7]), .A2(n63bar), .ZN(n48bar) );
  OR2_X1 U20 ( .A1(n46), .A2(n62), .ZN(y[6]) );
  AND2_X1 U20bar ( .A1(n46bar), .A2(n62bar), .ZN(ybar[6]) );
  OR2_X1 U21 ( .A1(n61), .A2(b[6]), .ZN(n45) );
  AND2_X1 U21bar ( .A1(n61bar), .A2(bbar[6]), .ZN(n45bar) );
  AND2_X1 U22 ( .A1(b[6]), .A2(n61), .ZN(n46) );
  OR2_X1 U22bar ( .A1(bbar[6]), .A2(n61bar), .ZN(n46bar) );
  OR2_X1 U23 ( .A1(n44), .A2(n60), .ZN(y[5]) );
  AND2_X1 U23bar ( .A1(n44bar), .A2(n60bar), .ZN(ybar[5]) );
  OR2_X1 U24 ( .A1(n59), .A2(b[5]), .ZN(n43) );
  AND2_X1 U24bar ( .A1(n59bar), .A2(bbar[5]), .ZN(n43bar) );
  AND2_X1 U25 ( .A1(b[5]), .A2(n59), .ZN(n44) );
  OR2_X1 U25bar ( .A1(bbar[5]), .A2(n59bar), .ZN(n44bar) );
  OR2_X1 U26 ( .A1(n42), .A2(n58), .ZN(y[4]) );
  AND2_X1 U26bar ( .A1(n42bar), .A2(n58bar), .ZN(ybar[4]) );
  OR2_X1 U27 ( .A1(n57), .A2(b[4]), .ZN(n41) );
  AND2_X1 U27bar ( .A1(n57bar), .A2(bbar[4]), .ZN(n41bar) );
  AND2_X1 U28 ( .A1(b[4]), .A2(n57), .ZN(n42) );
  OR2_X1 U28bar ( .A1(bbar[4]), .A2(n57bar), .ZN(n42bar) );
  OR2_X1 U29 ( .A1(n40), .A2(n56), .ZN(y[3]) );
  AND2_X1 U29bar ( .A1(n40bar), .A2(n56bar), .ZN(ybar[3]) );
  OR2_X1 U30 ( .A1(n55), .A2(b[3]), .ZN(n39) );
  AND2_X1 U30bar ( .A1(n55bar), .A2(bbar[3]), .ZN(n39bar) );
  AND2_X1 U31 ( .A1(b[3]), .A2(n55), .ZN(n40) );
  OR2_X1 U31bar ( .A1(bbar[3]), .A2(n55bar), .ZN(n40bar) );
  OR2_X1 U32 ( .A1(n38), .A2(n54), .ZN(y[2]) );
  AND2_X1 U32bar ( .A1(n38bar), .A2(n54bar), .ZN(ybar[2]) );
  OR2_X1 U33 ( .A1(n53), .A2(b[2]), .ZN(n37) );
  AND2_X1 U33bar ( .A1(n53bar), .A2(bbar[2]), .ZN(n37bar) );
  AND2_X1 U34 ( .A1(b[2]), .A2(n53), .ZN(n38) );
  OR2_X1 U34bar ( .A1(bbar[2]), .A2(n53bar), .ZN(n38bar) );
  OR2_X1 U35 ( .A1(n36), .A2(n52), .ZN(y[1]) );
  AND2_X1 U35bar ( .A1(n36bar), .A2(n52bar), .ZN(ybar[1]) );
  OR2_X1 U36 ( .A1(n51), .A2(b[1]), .ZN(n35) );
  AND2_X1 U36bar ( .A1(n51bar), .A2(bbar[1]), .ZN(n35bar) );
  AND2_X1 U37 ( .A1(b[1]), .A2(n51), .ZN(n36) );
  OR2_X1 U37bar ( .A1(bbar[1]), .A2(n51bar), .ZN(n36bar) );
  OR2_X1 U38 ( .A1(n34), .A2(n50), .ZN(y[0]) );
  AND2_X1 U38bar ( .A1(n34bar), .A2(n50bar), .ZN(ybar[0]) );
  OR2_X1 U39 ( .A1(n49), .A2(b[0]), .ZN(n33) );
  AND2_X1 U39bar ( .A1(n49bar), .A2(bbar[0]), .ZN(n33bar) );
  AND2_X1 U40 ( .A1(b[0]), .A2(n49), .ZN(n34) );
  OR2_X1 U40bar ( .A1(bbar[0]), .A2(n49bar), .ZN(n34bar) );
endmodule

module byteXor_9 ( a, abar, b, bbar, y, ybar );

  input wire [7:0] a;
  input wire [7:0] b;
  input wire [7:0] abar;
  input wire [7:0] bbar;
//input_done

  output wire [7:0] y;
  output wire [7:0] ybar;
//output_done

  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n33bar;
  wire n34bar;
  wire n35bar;
  wire n36bar;
  wire n37bar;
  wire n38bar;
  wire n39bar;
  wire n40bar;
  wire n41bar;
  wire n42bar;
  wire n43bar;
  wire n44bar;
  wire n45bar;
  wire n46bar;
  wire n47bar;
  wire n48bar;
  wire n49bar;
  wire n50bar;
  wire n51bar;
  wire n52bar;
  wire n53bar;
  wire n54bar;
  wire n55bar;
  wire n56bar;
  wire n57bar;
  wire n58bar;
  wire n59bar;
  wire n60bar;
  wire n61bar;
  wire n62bar;
  wire n63bar;
  wire n64bar;
//wire_done

 //assign_done

  assign n64bar = n47;
  assign n64 = n47bar;
  assign n63bar = a[7];
  assign n63 = abar[7];
  assign n62bar = n45;
  assign n62 = n45bar;
  assign n61bar = a[6];
  assign n61 = abar[6];
  assign n60bar = n43;
  assign n60 = n43bar;
  assign n59bar = a[5];
  assign n59 = abar[5];
  assign n58bar = n41;
  assign n58 = n41bar;
  assign n57bar = a[4];
  assign n57 = abar[4];
  assign n56bar = n39;
  assign n56 = n39bar;
  assign n55bar = a[3];
  assign n55 = abar[3];
  assign n54bar = n37;
  assign n54 = n37bar;
  assign n53bar = a[2];
  assign n53 = abar[2];
  assign n52bar = n35;
  assign n52 = n35bar;
  assign n51bar = a[1];
  assign n51 = abar[1];
  assign n50bar = n33;
  assign n50 = n33bar;
  assign n49bar = a[0];
  assign n49 = abar[0];
  OR2_X1 U17 ( .A1(n48), .A2(n64), .ZN(y[7]) );
  AND2_X1 U17bar ( .A1(n48bar), .A2(n64bar), .ZN(ybar[7]) );
  OR2_X1 U18 ( .A1(n63), .A2(b[7]), .ZN(n47) );
  AND2_X1 U18bar ( .A1(n63bar), .A2(bbar[7]), .ZN(n47bar) );
  AND2_X1 U19 ( .A1(b[7]), .A2(n63), .ZN(n48) );
  OR2_X1 U19bar ( .A1(bbar[7]), .A2(n63bar), .ZN(n48bar) );
  OR2_X1 U20 ( .A1(n46), .A2(n62), .ZN(y[6]) );
  AND2_X1 U20bar ( .A1(n46bar), .A2(n62bar), .ZN(ybar[6]) );
  OR2_X1 U21 ( .A1(n61), .A2(b[6]), .ZN(n45) );
  AND2_X1 U21bar ( .A1(n61bar), .A2(bbar[6]), .ZN(n45bar) );
  AND2_X1 U22 ( .A1(b[6]), .A2(n61), .ZN(n46) );
  OR2_X1 U22bar ( .A1(bbar[6]), .A2(n61bar), .ZN(n46bar) );
  OR2_X1 U23 ( .A1(n44), .A2(n60), .ZN(y[5]) );
  AND2_X1 U23bar ( .A1(n44bar), .A2(n60bar), .ZN(ybar[5]) );
  OR2_X1 U24 ( .A1(n59), .A2(b[5]), .ZN(n43) );
  AND2_X1 U24bar ( .A1(n59bar), .A2(bbar[5]), .ZN(n43bar) );
  AND2_X1 U25 ( .A1(b[5]), .A2(n59), .ZN(n44) );
  OR2_X1 U25bar ( .A1(bbar[5]), .A2(n59bar), .ZN(n44bar) );
  OR2_X1 U26 ( .A1(n42), .A2(n58), .ZN(y[4]) );
  AND2_X1 U26bar ( .A1(n42bar), .A2(n58bar), .ZN(ybar[4]) );
  OR2_X1 U27 ( .A1(n57), .A2(b[4]), .ZN(n41) );
  AND2_X1 U27bar ( .A1(n57bar), .A2(bbar[4]), .ZN(n41bar) );
  AND2_X1 U28 ( .A1(b[4]), .A2(n57), .ZN(n42) );
  OR2_X1 U28bar ( .A1(bbar[4]), .A2(n57bar), .ZN(n42bar) );
  OR2_X1 U29 ( .A1(n40), .A2(n56), .ZN(y[3]) );
  AND2_X1 U29bar ( .A1(n40bar), .A2(n56bar), .ZN(ybar[3]) );
  OR2_X1 U30 ( .A1(n55), .A2(b[3]), .ZN(n39) );
  AND2_X1 U30bar ( .A1(n55bar), .A2(bbar[3]), .ZN(n39bar) );
  AND2_X1 U31 ( .A1(b[3]), .A2(n55), .ZN(n40) );
  OR2_X1 U31bar ( .A1(bbar[3]), .A2(n55bar), .ZN(n40bar) );
  OR2_X1 U32 ( .A1(n38), .A2(n54), .ZN(y[2]) );
  AND2_X1 U32bar ( .A1(n38bar), .A2(n54bar), .ZN(ybar[2]) );
  OR2_X1 U33 ( .A1(n53), .A2(b[2]), .ZN(n37) );
  AND2_X1 U33bar ( .A1(n53bar), .A2(bbar[2]), .ZN(n37bar) );
  AND2_X1 U34 ( .A1(b[2]), .A2(n53), .ZN(n38) );
  OR2_X1 U34bar ( .A1(bbar[2]), .A2(n53bar), .ZN(n38bar) );
  OR2_X1 U35 ( .A1(n36), .A2(n52), .ZN(y[1]) );
  AND2_X1 U35bar ( .A1(n36bar), .A2(n52bar), .ZN(ybar[1]) );
  OR2_X1 U36 ( .A1(n51), .A2(b[1]), .ZN(n35) );
  AND2_X1 U36bar ( .A1(n51bar), .A2(bbar[1]), .ZN(n35bar) );
  AND2_X1 U37 ( .A1(b[1]), .A2(n51), .ZN(n36) );
  OR2_X1 U37bar ( .A1(bbar[1]), .A2(n51bar), .ZN(n36bar) );
  OR2_X1 U38 ( .A1(n34), .A2(n50), .ZN(y[0]) );
  AND2_X1 U38bar ( .A1(n34bar), .A2(n50bar), .ZN(ybar[0]) );
  OR2_X1 U39 ( .A1(n49), .A2(b[0]), .ZN(n33) );
  AND2_X1 U39bar ( .A1(n49bar), .A2(bbar[0]), .ZN(n33bar) );
  AND2_X1 U40 ( .A1(b[0]), .A2(n49), .ZN(n34) );
  OR2_X1 U40bar ( .A1(bbar[0]), .A2(n49bar), .ZN(n34bar) );
endmodule

module byteXor4_5 ( a, abar, b, bbar, c, cbar, d, dbar, y, ybar );

  input wire [7:0] a;
  input wire [7:0] b;
  input wire [7:0] c;
  input wire [7:0] d;
  input wire [7:0] abar;
  input wire [7:0] bbar;
  input wire [7:0] cbar;
  input wire [7:0] dbar;
//input_done

  output wire [7:0] y;
  output wire [7:0] ybar;
//output_done

  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n113bar;
  wire n114bar;
  wire n115bar;
  wire n116bar;
  wire n117bar;
  wire n118bar;
  wire n119bar;
  wire n120bar;
  wire n121bar;
  wire n122bar;
  wire n123bar;
  wire n124bar;
  wire n125bar;
  wire n126bar;
  wire n127bar;
  wire n128bar;
  wire n129bar;
  wire n130bar;
  wire n131bar;
  wire n132bar;
  wire n133bar;
  wire n134bar;
  wire n135bar;
  wire n136bar;
  wire n137bar;
  wire n138bar;
  wire n139bar;
  wire n140bar;
  wire n141bar;
  wire n142bar;
  wire n143bar;
  wire n144bar;
  wire n145bar;
  wire n146bar;
  wire n147bar;
  wire n148bar;
  wire n149bar;
  wire n150bar;
  wire n151bar;
  wire n152bar;
  wire n153bar;
  wire n154bar;
  wire n155bar;
  wire n156bar;
  wire n157bar;
  wire n158bar;
  wire n159bar;
  wire n160bar;
  wire n161bar;
  wire n162bar;
  wire n163bar;
  wire n164bar;
  wire n165bar;
  wire n166bar;
  wire n167bar;
  wire n168bar;
  wire n169bar;
  wire n170bar;
  wire n171bar;
  wire n172bar;
  wire n173bar;
  wire n174bar;
  wire n175bar;
  wire n176bar;
  wire n177bar;
  wire n178bar;
  wire n179bar;
  wire n180bar;
  wire n181bar;
  wire n182bar;
  wire n183bar;
  wire n184bar;
  wire n185bar;
  wire n186bar;
  wire n187bar;
  wire n188bar;
  wire n189bar;
  wire n190bar;
  wire n191bar;
  wire n192bar;
  wire n193bar;
  wire n194bar;
  wire n195bar;
  wire n196bar;
  wire n197bar;
  wire n198bar;
  wire n199bar;
  wire n200bar;
  wire n201bar;
  wire n202bar;
  wire n203bar;
  wire n204bar;
  wire n205bar;
  wire n206bar;
  wire n207bar;
  wire n208bar;
  wire n209bar;
  wire n210bar;
  wire n211bar;
  wire n212bar;
  wire n213bar;
  wire n214bar;
  wire n215bar;
  wire n216bar;
  wire n217bar;
  wire n218bar;
  wire n219bar;
  wire n220bar;
  wire n221bar;
  wire n222bar;
  wire n223bar;
  wire n224bar;
//wire_done

 //assign_done

  assign n224bar = n175;
  assign n224 = n175bar;
  assign n223bar = a[7];
  assign n223 = abar[7];
  assign n222bar = n167;
  assign n222 = n167bar;
  assign n221bar = a[6];
  assign n221 = abar[6];
  assign n220bar = n159;
  assign n220 = n159bar;
  assign n219bar = a[5];
  assign n219 = abar[5];
  assign n218bar = n151;
  assign n218 = n151bar;
  assign n217bar = a[4];
  assign n217 = abar[4];
  assign n216bar = n143;
  assign n216 = n143bar;
  assign n215bar = a[3];
  assign n215 = abar[3];
  assign n214bar = n135;
  assign n214 = n135bar;
  assign n213bar = a[2];
  assign n213 = abar[2];
  assign n212bar = n127;
  assign n212 = n127bar;
  assign n211bar = a[1];
  assign n211 = abar[1];
  assign n210bar = n119;
  assign n210 = n119bar;
  assign n209bar = a[0];
  assign n209 = abar[0];
  assign n208bar = b[7];
  assign n208 = bbar[7];
  assign n207bar = b[6];
  assign n207 = bbar[6];
  assign n206bar = b[5];
  assign n206 = bbar[5];
  assign n205bar = b[4];
  assign n205 = bbar[4];
  assign n204bar = b[3];
  assign n204 = bbar[3];
  assign n203bar = b[2];
  assign n203 = bbar[2];
  assign n202bar = b[1];
  assign n202 = bbar[1];
  assign n201bar = b[0];
  assign n201 = bbar[0];
  assign n200bar = n171;
  assign n200 = n171bar;
  assign n199bar = c[7];
  assign n199 = cbar[7];
  assign n198bar = n163;
  assign n198 = n163bar;
  assign n197bar = c[6];
  assign n197 = cbar[6];
  assign n196bar = n155;
  assign n196 = n155bar;
  assign n195bar = c[5];
  assign n195 = cbar[5];
  assign n194bar = n147;
  assign n194 = n147bar;
  assign n193bar = c[4];
  assign n193 = cbar[4];
  assign n192bar = n139;
  assign n192 = n139bar;
  assign n191bar = c[3];
  assign n191 = cbar[3];
  assign n190bar = n131;
  assign n190 = n131bar;
  assign n189bar = c[2];
  assign n189 = cbar[2];
  assign n188bar = n123;
  assign n188 = n123bar;
  assign n187bar = c[1];
  assign n187 = cbar[1];
  assign n186bar = n115;
  assign n186 = n115bar;
  assign n185bar = c[0];
  assign n185 = cbar[0];
  assign n184bar = d[7];
  assign n184 = dbar[7];
  assign n183bar = d[6];
  assign n183 = dbar[6];
  assign n182bar = d[5];
  assign n182 = dbar[5];
  assign n181bar = d[4];
  assign n181 = dbar[4];
  assign n180bar = d[3];
  assign n180 = dbar[3];
  assign n179bar = d[2];
  assign n179 = dbar[2];
  assign n178bar = d[1];
  assign n178 = dbar[1];
  assign n177bar = d[0];
  assign n177 = dbar[0];
  OR2_X1 U49 ( .A1(n176), .A2(n224), .ZN(y[7]) );
  AND2_X1 U49bar ( .A1(n176bar), .A2(n224bar), .ZN(ybar[7]) );
  OR2_X1 U50 ( .A1(n174), .A2(n200), .ZN(n175) );
  AND2_X1 U50bar ( .A1(n174bar), .A2(n200bar), .ZN(n175bar) );
  AND2_X1 U51 ( .A1(n200), .A2(n174), .ZN(n176) );
  OR2_X1 U51bar ( .A1(n200bar), .A2(n174bar), .ZN(n176bar) );
  AND2_X1 U52 ( .A1(n173), .A2(n172), .ZN(n174) );
  OR2_X1 U52bar ( .A1(n173bar), .A2(n172bar), .ZN(n174bar) );
  OR2_X1 U53 ( .A1(n223), .A2(b[7]), .ZN(n172) );
  AND2_X1 U53bar ( .A1(n223bar), .A2(bbar[7]), .ZN(n172bar) );
  OR2_X1 U54 ( .A1(n208), .A2(a[7]), .ZN(n173) );
  AND2_X1 U54bar ( .A1(n208bar), .A2(abar[7]), .ZN(n173bar) );
  AND2_X1 U55 ( .A1(n170), .A2(n169), .ZN(n171) );
  OR2_X1 U55bar ( .A1(n170bar), .A2(n169bar), .ZN(n171bar) );
  OR2_X1 U56 ( .A1(n199), .A2(d[7]), .ZN(n169) );
  AND2_X1 U56bar ( .A1(n199bar), .A2(dbar[7]), .ZN(n169bar) );
  OR2_X1 U57 ( .A1(n184), .A2(c[7]), .ZN(n170) );
  AND2_X1 U57bar ( .A1(n184bar), .A2(cbar[7]), .ZN(n170bar) );
  OR2_X1 U58 ( .A1(n168), .A2(n222), .ZN(y[6]) );
  AND2_X1 U58bar ( .A1(n168bar), .A2(n222bar), .ZN(ybar[6]) );
  OR2_X1 U59 ( .A1(n166), .A2(n198), .ZN(n167) );
  AND2_X1 U59bar ( .A1(n166bar), .A2(n198bar), .ZN(n167bar) );
  AND2_X1 U60 ( .A1(n198), .A2(n166), .ZN(n168) );
  OR2_X1 U60bar ( .A1(n198bar), .A2(n166bar), .ZN(n168bar) );
  AND2_X1 U61 ( .A1(n165), .A2(n164), .ZN(n166) );
  OR2_X1 U61bar ( .A1(n165bar), .A2(n164bar), .ZN(n166bar) );
  OR2_X1 U62 ( .A1(n221), .A2(b[6]), .ZN(n164) );
  AND2_X1 U62bar ( .A1(n221bar), .A2(bbar[6]), .ZN(n164bar) );
  OR2_X1 U63 ( .A1(n207), .A2(a[6]), .ZN(n165) );
  AND2_X1 U63bar ( .A1(n207bar), .A2(abar[6]), .ZN(n165bar) );
  AND2_X1 U64 ( .A1(n162), .A2(n161), .ZN(n163) );
  OR2_X1 U64bar ( .A1(n162bar), .A2(n161bar), .ZN(n163bar) );
  OR2_X1 U65 ( .A1(n197), .A2(d[6]), .ZN(n161) );
  AND2_X1 U65bar ( .A1(n197bar), .A2(dbar[6]), .ZN(n161bar) );
  OR2_X1 U66 ( .A1(n183), .A2(c[6]), .ZN(n162) );
  AND2_X1 U66bar ( .A1(n183bar), .A2(cbar[6]), .ZN(n162bar) );
  OR2_X1 U67 ( .A1(n160), .A2(n220), .ZN(y[5]) );
  AND2_X1 U67bar ( .A1(n160bar), .A2(n220bar), .ZN(ybar[5]) );
  OR2_X1 U68 ( .A1(n158), .A2(n196), .ZN(n159) );
  AND2_X1 U68bar ( .A1(n158bar), .A2(n196bar), .ZN(n159bar) );
  AND2_X1 U69 ( .A1(n196), .A2(n158), .ZN(n160) );
  OR2_X1 U69bar ( .A1(n196bar), .A2(n158bar), .ZN(n160bar) );
  AND2_X1 U70 ( .A1(n157), .A2(n156), .ZN(n158) );
  OR2_X1 U70bar ( .A1(n157bar), .A2(n156bar), .ZN(n158bar) );
  OR2_X1 U71 ( .A1(n219), .A2(b[5]), .ZN(n156) );
  AND2_X1 U71bar ( .A1(n219bar), .A2(bbar[5]), .ZN(n156bar) );
  OR2_X1 U72 ( .A1(n206), .A2(a[5]), .ZN(n157) );
  AND2_X1 U72bar ( .A1(n206bar), .A2(abar[5]), .ZN(n157bar) );
  AND2_X1 U73 ( .A1(n154), .A2(n153), .ZN(n155) );
  OR2_X1 U73bar ( .A1(n154bar), .A2(n153bar), .ZN(n155bar) );
  OR2_X1 U74 ( .A1(n195), .A2(d[5]), .ZN(n153) );
  AND2_X1 U74bar ( .A1(n195bar), .A2(dbar[5]), .ZN(n153bar) );
  OR2_X1 U75 ( .A1(n182), .A2(c[5]), .ZN(n154) );
  AND2_X1 U75bar ( .A1(n182bar), .A2(cbar[5]), .ZN(n154bar) );
  OR2_X1 U76 ( .A1(n152), .A2(n218), .ZN(y[4]) );
  AND2_X1 U76bar ( .A1(n152bar), .A2(n218bar), .ZN(ybar[4]) );
  OR2_X1 U77 ( .A1(n150), .A2(n194), .ZN(n151) );
  AND2_X1 U77bar ( .A1(n150bar), .A2(n194bar), .ZN(n151bar) );
  AND2_X1 U78 ( .A1(n194), .A2(n150), .ZN(n152) );
  OR2_X1 U78bar ( .A1(n194bar), .A2(n150bar), .ZN(n152bar) );
  AND2_X1 U79 ( .A1(n149), .A2(n148), .ZN(n150) );
  OR2_X1 U79bar ( .A1(n149bar), .A2(n148bar), .ZN(n150bar) );
  OR2_X1 U80 ( .A1(n217), .A2(b[4]), .ZN(n148) );
  AND2_X1 U80bar ( .A1(n217bar), .A2(bbar[4]), .ZN(n148bar) );
  OR2_X1 U81 ( .A1(n205), .A2(a[4]), .ZN(n149) );
  AND2_X1 U81bar ( .A1(n205bar), .A2(abar[4]), .ZN(n149bar) );
  AND2_X1 U82 ( .A1(n146), .A2(n145), .ZN(n147) );
  OR2_X1 U82bar ( .A1(n146bar), .A2(n145bar), .ZN(n147bar) );
  OR2_X1 U83 ( .A1(n193), .A2(d[4]), .ZN(n145) );
  AND2_X1 U83bar ( .A1(n193bar), .A2(dbar[4]), .ZN(n145bar) );
  OR2_X1 U84 ( .A1(n181), .A2(c[4]), .ZN(n146) );
  AND2_X1 U84bar ( .A1(n181bar), .A2(cbar[4]), .ZN(n146bar) );
  OR2_X1 U85 ( .A1(n144), .A2(n216), .ZN(y[3]) );
  AND2_X1 U85bar ( .A1(n144bar), .A2(n216bar), .ZN(ybar[3]) );
  OR2_X1 U86 ( .A1(n142), .A2(n192), .ZN(n143) );
  AND2_X1 U86bar ( .A1(n142bar), .A2(n192bar), .ZN(n143bar) );
  AND2_X1 U87 ( .A1(n192), .A2(n142), .ZN(n144) );
  OR2_X1 U87bar ( .A1(n192bar), .A2(n142bar), .ZN(n144bar) );
  AND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(n142) );
  OR2_X1 U88bar ( .A1(n141bar), .A2(n140bar), .ZN(n142bar) );
  OR2_X1 U89 ( .A1(n215), .A2(b[3]), .ZN(n140) );
  AND2_X1 U89bar ( .A1(n215bar), .A2(bbar[3]), .ZN(n140bar) );
  OR2_X1 U90 ( .A1(n204), .A2(a[3]), .ZN(n141) );
  AND2_X1 U90bar ( .A1(n204bar), .A2(abar[3]), .ZN(n141bar) );
  AND2_X1 U91 ( .A1(n138), .A2(n137), .ZN(n139) );
  OR2_X1 U91bar ( .A1(n138bar), .A2(n137bar), .ZN(n139bar) );
  OR2_X1 U92 ( .A1(n191), .A2(d[3]), .ZN(n137) );
  AND2_X1 U92bar ( .A1(n191bar), .A2(dbar[3]), .ZN(n137bar) );
  OR2_X1 U93 ( .A1(n180), .A2(c[3]), .ZN(n138) );
  AND2_X1 U93bar ( .A1(n180bar), .A2(cbar[3]), .ZN(n138bar) );
  OR2_X1 U94 ( .A1(n136), .A2(n214), .ZN(y[2]) );
  AND2_X1 U94bar ( .A1(n136bar), .A2(n214bar), .ZN(ybar[2]) );
  OR2_X1 U95 ( .A1(n134), .A2(n190), .ZN(n135) );
  AND2_X1 U95bar ( .A1(n134bar), .A2(n190bar), .ZN(n135bar) );
  AND2_X1 U96 ( .A1(n190), .A2(n134), .ZN(n136) );
  OR2_X1 U96bar ( .A1(n190bar), .A2(n134bar), .ZN(n136bar) );
  AND2_X1 U97 ( .A1(n133), .A2(n132), .ZN(n134) );
  OR2_X1 U97bar ( .A1(n133bar), .A2(n132bar), .ZN(n134bar) );
  OR2_X1 U98 ( .A1(n213), .A2(b[2]), .ZN(n132) );
  AND2_X1 U98bar ( .A1(n213bar), .A2(bbar[2]), .ZN(n132bar) );
  OR2_X1 U99 ( .A1(n203), .A2(a[2]), .ZN(n133) );
  AND2_X1 U99bar ( .A1(n203bar), .A2(abar[2]), .ZN(n133bar) );
  AND2_X1 U100 ( .A1(n130), .A2(n129), .ZN(n131) );
  OR2_X1 U100bar ( .A1(n130bar), .A2(n129bar), .ZN(n131bar) );
  OR2_X1 U101 ( .A1(n189), .A2(d[2]), .ZN(n129) );
  AND2_X1 U101bar ( .A1(n189bar), .A2(dbar[2]), .ZN(n129bar) );
  OR2_X1 U102 ( .A1(n179), .A2(c[2]), .ZN(n130) );
  AND2_X1 U102bar ( .A1(n179bar), .A2(cbar[2]), .ZN(n130bar) );
  OR2_X1 U103 ( .A1(n128), .A2(n212), .ZN(y[1]) );
  AND2_X1 U103bar ( .A1(n128bar), .A2(n212bar), .ZN(ybar[1]) );
  OR2_X1 U104 ( .A1(n126), .A2(n188), .ZN(n127) );
  AND2_X1 U104bar ( .A1(n126bar), .A2(n188bar), .ZN(n127bar) );
  AND2_X1 U105 ( .A1(n188), .A2(n126), .ZN(n128) );
  OR2_X1 U105bar ( .A1(n188bar), .A2(n126bar), .ZN(n128bar) );
  AND2_X1 U106 ( .A1(n125), .A2(n124), .ZN(n126) );
  OR2_X1 U106bar ( .A1(n125bar), .A2(n124bar), .ZN(n126bar) );
  OR2_X1 U107 ( .A1(n211), .A2(b[1]), .ZN(n124) );
  AND2_X1 U107bar ( .A1(n211bar), .A2(bbar[1]), .ZN(n124bar) );
  OR2_X1 U108 ( .A1(n202), .A2(a[1]), .ZN(n125) );
  AND2_X1 U108bar ( .A1(n202bar), .A2(abar[1]), .ZN(n125bar) );
  AND2_X1 U109 ( .A1(n122), .A2(n121), .ZN(n123) );
  OR2_X1 U109bar ( .A1(n122bar), .A2(n121bar), .ZN(n123bar) );
  OR2_X1 U110 ( .A1(n187), .A2(d[1]), .ZN(n121) );
  AND2_X1 U110bar ( .A1(n187bar), .A2(dbar[1]), .ZN(n121bar) );
  OR2_X1 U111 ( .A1(n178), .A2(c[1]), .ZN(n122) );
  AND2_X1 U111bar ( .A1(n178bar), .A2(cbar[1]), .ZN(n122bar) );
  OR2_X1 U112 ( .A1(n120), .A2(n210), .ZN(y[0]) );
  AND2_X1 U112bar ( .A1(n120bar), .A2(n210bar), .ZN(ybar[0]) );
  OR2_X1 U113 ( .A1(n118), .A2(n186), .ZN(n119) );
  AND2_X1 U113bar ( .A1(n118bar), .A2(n186bar), .ZN(n119bar) );
  AND2_X1 U114 ( .A1(n186), .A2(n118), .ZN(n120) );
  OR2_X1 U114bar ( .A1(n186bar), .A2(n118bar), .ZN(n120bar) );
  AND2_X1 U115 ( .A1(n117), .A2(n116), .ZN(n118) );
  OR2_X1 U115bar ( .A1(n117bar), .A2(n116bar), .ZN(n118bar) );
  OR2_X1 U116 ( .A1(n209), .A2(b[0]), .ZN(n116) );
  AND2_X1 U116bar ( .A1(n209bar), .A2(bbar[0]), .ZN(n116bar) );
  OR2_X1 U117 ( .A1(n201), .A2(a[0]), .ZN(n117) );
  AND2_X1 U117bar ( .A1(n201bar), .A2(abar[0]), .ZN(n117bar) );
  AND2_X1 U118 ( .A1(n114), .A2(n113), .ZN(n115) );
  OR2_X1 U118bar ( .A1(n114bar), .A2(n113bar), .ZN(n115bar) );
  OR2_X1 U119 ( .A1(n185), .A2(d[0]), .ZN(n113) );
  AND2_X1 U119bar ( .A1(n185bar), .A2(dbar[0]), .ZN(n113bar) );
  OR2_X1 U120 ( .A1(n177), .A2(c[0]), .ZN(n114) );
  AND2_X1 U120bar ( .A1(n177bar), .A2(cbar[0]), .ZN(n114bar) );
endmodule

module byteXor4_6 ( a, abar, b, bbar, c, cbar, d, dbar, y, ybar );

  input wire [7:0] a;
  input wire [7:0] b;
  input wire [7:0] c;
  input wire [7:0] d;
  input wire [7:0] abar;
  input wire [7:0] bbar;
  input wire [7:0] cbar;
  input wire [7:0] dbar;
//input_done

  output wire [7:0] y;
  output wire [7:0] ybar;
//output_done

  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n113bar;
  wire n114bar;
  wire n115bar;
  wire n116bar;
  wire n117bar;
  wire n118bar;
  wire n119bar;
  wire n120bar;
  wire n121bar;
  wire n122bar;
  wire n123bar;
  wire n124bar;
  wire n125bar;
  wire n126bar;
  wire n127bar;
  wire n128bar;
  wire n129bar;
  wire n130bar;
  wire n131bar;
  wire n132bar;
  wire n133bar;
  wire n134bar;
  wire n135bar;
  wire n136bar;
  wire n137bar;
  wire n138bar;
  wire n139bar;
  wire n140bar;
  wire n141bar;
  wire n142bar;
  wire n143bar;
  wire n144bar;
  wire n145bar;
  wire n146bar;
  wire n147bar;
  wire n148bar;
  wire n149bar;
  wire n150bar;
  wire n151bar;
  wire n152bar;
  wire n153bar;
  wire n154bar;
  wire n155bar;
  wire n156bar;
  wire n157bar;
  wire n158bar;
  wire n159bar;
  wire n160bar;
  wire n161bar;
  wire n162bar;
  wire n163bar;
  wire n164bar;
  wire n165bar;
  wire n166bar;
  wire n167bar;
  wire n168bar;
  wire n169bar;
  wire n170bar;
  wire n171bar;
  wire n172bar;
  wire n173bar;
  wire n174bar;
  wire n175bar;
  wire n176bar;
  wire n177bar;
  wire n178bar;
  wire n179bar;
  wire n180bar;
  wire n181bar;
  wire n182bar;
  wire n183bar;
  wire n184bar;
  wire n185bar;
  wire n186bar;
  wire n187bar;
  wire n188bar;
  wire n189bar;
  wire n190bar;
  wire n191bar;
  wire n192bar;
  wire n193bar;
  wire n194bar;
  wire n195bar;
  wire n196bar;
  wire n197bar;
  wire n198bar;
  wire n199bar;
  wire n200bar;
  wire n201bar;
  wire n202bar;
  wire n203bar;
  wire n204bar;
  wire n205bar;
  wire n206bar;
  wire n207bar;
  wire n208bar;
  wire n209bar;
  wire n210bar;
  wire n211bar;
  wire n212bar;
  wire n213bar;
  wire n214bar;
  wire n215bar;
  wire n216bar;
  wire n217bar;
  wire n218bar;
  wire n219bar;
  wire n220bar;
  wire n221bar;
  wire n222bar;
  wire n223bar;
  wire n224bar;
//wire_done

 //assign_done

  assign n224bar = n175;
  assign n224 = n175bar;
  assign n223bar = a[7];
  assign n223 = abar[7];
  assign n222bar = n167;
  assign n222 = n167bar;
  assign n221bar = a[6];
  assign n221 = abar[6];
  assign n220bar = n159;
  assign n220 = n159bar;
  assign n219bar = a[5];
  assign n219 = abar[5];
  assign n218bar = n151;
  assign n218 = n151bar;
  assign n217bar = a[4];
  assign n217 = abar[4];
  assign n216bar = n143;
  assign n216 = n143bar;
  assign n215bar = a[3];
  assign n215 = abar[3];
  assign n214bar = n135;
  assign n214 = n135bar;
  assign n213bar = a[2];
  assign n213 = abar[2];
  assign n212bar = n127;
  assign n212 = n127bar;
  assign n211bar = a[1];
  assign n211 = abar[1];
  assign n210bar = n119;
  assign n210 = n119bar;
  assign n209bar = a[0];
  assign n209 = abar[0];
  assign n208bar = b[7];
  assign n208 = bbar[7];
  assign n207bar = b[6];
  assign n207 = bbar[6];
  assign n206bar = b[5];
  assign n206 = bbar[5];
  assign n205bar = b[4];
  assign n205 = bbar[4];
  assign n204bar = b[3];
  assign n204 = bbar[3];
  assign n203bar = b[2];
  assign n203 = bbar[2];
  assign n202bar = b[1];
  assign n202 = bbar[1];
  assign n201bar = b[0];
  assign n201 = bbar[0];
  assign n200bar = n171;
  assign n200 = n171bar;
  assign n199bar = c[7];
  assign n199 = cbar[7];
  assign n198bar = n163;
  assign n198 = n163bar;
  assign n197bar = c[6];
  assign n197 = cbar[6];
  assign n196bar = n155;
  assign n196 = n155bar;
  assign n195bar = c[5];
  assign n195 = cbar[5];
  assign n194bar = n147;
  assign n194 = n147bar;
  assign n193bar = c[4];
  assign n193 = cbar[4];
  assign n192bar = n139;
  assign n192 = n139bar;
  assign n191bar = c[3];
  assign n191 = cbar[3];
  assign n190bar = n131;
  assign n190 = n131bar;
  assign n189bar = c[2];
  assign n189 = cbar[2];
  assign n188bar = n123;
  assign n188 = n123bar;
  assign n187bar = c[1];
  assign n187 = cbar[1];
  assign n186bar = n115;
  assign n186 = n115bar;
  assign n185bar = c[0];
  assign n185 = cbar[0];
  assign n184bar = d[7];
  assign n184 = dbar[7];
  assign n183bar = d[6];
  assign n183 = dbar[6];
  assign n182bar = d[5];
  assign n182 = dbar[5];
  assign n181bar = d[4];
  assign n181 = dbar[4];
  assign n180bar = d[3];
  assign n180 = dbar[3];
  assign n179bar = d[2];
  assign n179 = dbar[2];
  assign n178bar = d[1];
  assign n178 = dbar[1];
  assign n177bar = d[0];
  assign n177 = dbar[0];
  OR2_X1 U49 ( .A1(n176), .A2(n224), .ZN(y[7]) );
  AND2_X1 U49bar ( .A1(n176bar), .A2(n224bar), .ZN(ybar[7]) );
  OR2_X1 U50 ( .A1(n174), .A2(n200), .ZN(n175) );
  AND2_X1 U50bar ( .A1(n174bar), .A2(n200bar), .ZN(n175bar) );
  AND2_X1 U51 ( .A1(n200), .A2(n174), .ZN(n176) );
  OR2_X1 U51bar ( .A1(n200bar), .A2(n174bar), .ZN(n176bar) );
  AND2_X1 U52 ( .A1(n173), .A2(n172), .ZN(n174) );
  OR2_X1 U52bar ( .A1(n173bar), .A2(n172bar), .ZN(n174bar) );
  OR2_X1 U53 ( .A1(n223), .A2(b[7]), .ZN(n172) );
  AND2_X1 U53bar ( .A1(n223bar), .A2(bbar[7]), .ZN(n172bar) );
  OR2_X1 U54 ( .A1(n208), .A2(a[7]), .ZN(n173) );
  AND2_X1 U54bar ( .A1(n208bar), .A2(abar[7]), .ZN(n173bar) );
  AND2_X1 U55 ( .A1(n170), .A2(n169), .ZN(n171) );
  OR2_X1 U55bar ( .A1(n170bar), .A2(n169bar), .ZN(n171bar) );
  OR2_X1 U56 ( .A1(n199), .A2(d[7]), .ZN(n169) );
  AND2_X1 U56bar ( .A1(n199bar), .A2(dbar[7]), .ZN(n169bar) );
  OR2_X1 U57 ( .A1(n184), .A2(c[7]), .ZN(n170) );
  AND2_X1 U57bar ( .A1(n184bar), .A2(cbar[7]), .ZN(n170bar) );
  OR2_X1 U58 ( .A1(n168), .A2(n222), .ZN(y[6]) );
  AND2_X1 U58bar ( .A1(n168bar), .A2(n222bar), .ZN(ybar[6]) );
  OR2_X1 U59 ( .A1(n166), .A2(n198), .ZN(n167) );
  AND2_X1 U59bar ( .A1(n166bar), .A2(n198bar), .ZN(n167bar) );
  AND2_X1 U60 ( .A1(n198), .A2(n166), .ZN(n168) );
  OR2_X1 U60bar ( .A1(n198bar), .A2(n166bar), .ZN(n168bar) );
  AND2_X1 U61 ( .A1(n165), .A2(n164), .ZN(n166) );
  OR2_X1 U61bar ( .A1(n165bar), .A2(n164bar), .ZN(n166bar) );
  OR2_X1 U62 ( .A1(n221), .A2(b[6]), .ZN(n164) );
  AND2_X1 U62bar ( .A1(n221bar), .A2(bbar[6]), .ZN(n164bar) );
  OR2_X1 U63 ( .A1(n207), .A2(a[6]), .ZN(n165) );
  AND2_X1 U63bar ( .A1(n207bar), .A2(abar[6]), .ZN(n165bar) );
  AND2_X1 U64 ( .A1(n162), .A2(n161), .ZN(n163) );
  OR2_X1 U64bar ( .A1(n162bar), .A2(n161bar), .ZN(n163bar) );
  OR2_X1 U65 ( .A1(n197), .A2(d[6]), .ZN(n161) );
  AND2_X1 U65bar ( .A1(n197bar), .A2(dbar[6]), .ZN(n161bar) );
  OR2_X1 U66 ( .A1(n183), .A2(c[6]), .ZN(n162) );
  AND2_X1 U66bar ( .A1(n183bar), .A2(cbar[6]), .ZN(n162bar) );
  OR2_X1 U67 ( .A1(n160), .A2(n220), .ZN(y[5]) );
  AND2_X1 U67bar ( .A1(n160bar), .A2(n220bar), .ZN(ybar[5]) );
  OR2_X1 U68 ( .A1(n158), .A2(n196), .ZN(n159) );
  AND2_X1 U68bar ( .A1(n158bar), .A2(n196bar), .ZN(n159bar) );
  AND2_X1 U69 ( .A1(n196), .A2(n158), .ZN(n160) );
  OR2_X1 U69bar ( .A1(n196bar), .A2(n158bar), .ZN(n160bar) );
  AND2_X1 U70 ( .A1(n157), .A2(n156), .ZN(n158) );
  OR2_X1 U70bar ( .A1(n157bar), .A2(n156bar), .ZN(n158bar) );
  OR2_X1 U71 ( .A1(n219), .A2(b[5]), .ZN(n156) );
  AND2_X1 U71bar ( .A1(n219bar), .A2(bbar[5]), .ZN(n156bar) );
  OR2_X1 U72 ( .A1(n206), .A2(a[5]), .ZN(n157) );
  AND2_X1 U72bar ( .A1(n206bar), .A2(abar[5]), .ZN(n157bar) );
  AND2_X1 U73 ( .A1(n154), .A2(n153), .ZN(n155) );
  OR2_X1 U73bar ( .A1(n154bar), .A2(n153bar), .ZN(n155bar) );
  OR2_X1 U74 ( .A1(n195), .A2(d[5]), .ZN(n153) );
  AND2_X1 U74bar ( .A1(n195bar), .A2(dbar[5]), .ZN(n153bar) );
  OR2_X1 U75 ( .A1(n182), .A2(c[5]), .ZN(n154) );
  AND2_X1 U75bar ( .A1(n182bar), .A2(cbar[5]), .ZN(n154bar) );
  OR2_X1 U76 ( .A1(n152), .A2(n218), .ZN(y[4]) );
  AND2_X1 U76bar ( .A1(n152bar), .A2(n218bar), .ZN(ybar[4]) );
  OR2_X1 U77 ( .A1(n150), .A2(n194), .ZN(n151) );
  AND2_X1 U77bar ( .A1(n150bar), .A2(n194bar), .ZN(n151bar) );
  AND2_X1 U78 ( .A1(n194), .A2(n150), .ZN(n152) );
  OR2_X1 U78bar ( .A1(n194bar), .A2(n150bar), .ZN(n152bar) );
  AND2_X1 U79 ( .A1(n149), .A2(n148), .ZN(n150) );
  OR2_X1 U79bar ( .A1(n149bar), .A2(n148bar), .ZN(n150bar) );
  OR2_X1 U80 ( .A1(n217), .A2(b[4]), .ZN(n148) );
  AND2_X1 U80bar ( .A1(n217bar), .A2(bbar[4]), .ZN(n148bar) );
  OR2_X1 U81 ( .A1(n205), .A2(a[4]), .ZN(n149) );
  AND2_X1 U81bar ( .A1(n205bar), .A2(abar[4]), .ZN(n149bar) );
  AND2_X1 U82 ( .A1(n146), .A2(n145), .ZN(n147) );
  OR2_X1 U82bar ( .A1(n146bar), .A2(n145bar), .ZN(n147bar) );
  OR2_X1 U83 ( .A1(n193), .A2(d[4]), .ZN(n145) );
  AND2_X1 U83bar ( .A1(n193bar), .A2(dbar[4]), .ZN(n145bar) );
  OR2_X1 U84 ( .A1(n181), .A2(c[4]), .ZN(n146) );
  AND2_X1 U84bar ( .A1(n181bar), .A2(cbar[4]), .ZN(n146bar) );
  OR2_X1 U85 ( .A1(n144), .A2(n216), .ZN(y[3]) );
  AND2_X1 U85bar ( .A1(n144bar), .A2(n216bar), .ZN(ybar[3]) );
  OR2_X1 U86 ( .A1(n142), .A2(n192), .ZN(n143) );
  AND2_X1 U86bar ( .A1(n142bar), .A2(n192bar), .ZN(n143bar) );
  AND2_X1 U87 ( .A1(n192), .A2(n142), .ZN(n144) );
  OR2_X1 U87bar ( .A1(n192bar), .A2(n142bar), .ZN(n144bar) );
  AND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(n142) );
  OR2_X1 U88bar ( .A1(n141bar), .A2(n140bar), .ZN(n142bar) );
  OR2_X1 U89 ( .A1(n215), .A2(b[3]), .ZN(n140) );
  AND2_X1 U89bar ( .A1(n215bar), .A2(bbar[3]), .ZN(n140bar) );
  OR2_X1 U90 ( .A1(n204), .A2(a[3]), .ZN(n141) );
  AND2_X1 U90bar ( .A1(n204bar), .A2(abar[3]), .ZN(n141bar) );
  AND2_X1 U91 ( .A1(n138), .A2(n137), .ZN(n139) );
  OR2_X1 U91bar ( .A1(n138bar), .A2(n137bar), .ZN(n139bar) );
  OR2_X1 U92 ( .A1(n191), .A2(d[3]), .ZN(n137) );
  AND2_X1 U92bar ( .A1(n191bar), .A2(dbar[3]), .ZN(n137bar) );
  OR2_X1 U93 ( .A1(n180), .A2(c[3]), .ZN(n138) );
  AND2_X1 U93bar ( .A1(n180bar), .A2(cbar[3]), .ZN(n138bar) );
  OR2_X1 U94 ( .A1(n136), .A2(n214), .ZN(y[2]) );
  AND2_X1 U94bar ( .A1(n136bar), .A2(n214bar), .ZN(ybar[2]) );
  OR2_X1 U95 ( .A1(n134), .A2(n190), .ZN(n135) );
  AND2_X1 U95bar ( .A1(n134bar), .A2(n190bar), .ZN(n135bar) );
  AND2_X1 U96 ( .A1(n190), .A2(n134), .ZN(n136) );
  OR2_X1 U96bar ( .A1(n190bar), .A2(n134bar), .ZN(n136bar) );
  AND2_X1 U97 ( .A1(n133), .A2(n132), .ZN(n134) );
  OR2_X1 U97bar ( .A1(n133bar), .A2(n132bar), .ZN(n134bar) );
  OR2_X1 U98 ( .A1(n213), .A2(b[2]), .ZN(n132) );
  AND2_X1 U98bar ( .A1(n213bar), .A2(bbar[2]), .ZN(n132bar) );
  OR2_X1 U99 ( .A1(n203), .A2(a[2]), .ZN(n133) );
  AND2_X1 U99bar ( .A1(n203bar), .A2(abar[2]), .ZN(n133bar) );
  AND2_X1 U100 ( .A1(n130), .A2(n129), .ZN(n131) );
  OR2_X1 U100bar ( .A1(n130bar), .A2(n129bar), .ZN(n131bar) );
  OR2_X1 U101 ( .A1(n189), .A2(d[2]), .ZN(n129) );
  AND2_X1 U101bar ( .A1(n189bar), .A2(dbar[2]), .ZN(n129bar) );
  OR2_X1 U102 ( .A1(n179), .A2(c[2]), .ZN(n130) );
  AND2_X1 U102bar ( .A1(n179bar), .A2(cbar[2]), .ZN(n130bar) );
  OR2_X1 U103 ( .A1(n128), .A2(n212), .ZN(y[1]) );
  AND2_X1 U103bar ( .A1(n128bar), .A2(n212bar), .ZN(ybar[1]) );
  OR2_X1 U104 ( .A1(n126), .A2(n188), .ZN(n127) );
  AND2_X1 U104bar ( .A1(n126bar), .A2(n188bar), .ZN(n127bar) );
  AND2_X1 U105 ( .A1(n188), .A2(n126), .ZN(n128) );
  OR2_X1 U105bar ( .A1(n188bar), .A2(n126bar), .ZN(n128bar) );
  AND2_X1 U106 ( .A1(n125), .A2(n124), .ZN(n126) );
  OR2_X1 U106bar ( .A1(n125bar), .A2(n124bar), .ZN(n126bar) );
  OR2_X1 U107 ( .A1(n211), .A2(b[1]), .ZN(n124) );
  AND2_X1 U107bar ( .A1(n211bar), .A2(bbar[1]), .ZN(n124bar) );
  OR2_X1 U108 ( .A1(n202), .A2(a[1]), .ZN(n125) );
  AND2_X1 U108bar ( .A1(n202bar), .A2(abar[1]), .ZN(n125bar) );
  AND2_X1 U109 ( .A1(n122), .A2(n121), .ZN(n123) );
  OR2_X1 U109bar ( .A1(n122bar), .A2(n121bar), .ZN(n123bar) );
  OR2_X1 U110 ( .A1(n187), .A2(d[1]), .ZN(n121) );
  AND2_X1 U110bar ( .A1(n187bar), .A2(dbar[1]), .ZN(n121bar) );
  OR2_X1 U111 ( .A1(n178), .A2(c[1]), .ZN(n122) );
  AND2_X1 U111bar ( .A1(n178bar), .A2(cbar[1]), .ZN(n122bar) );
  OR2_X1 U112 ( .A1(n120), .A2(n210), .ZN(y[0]) );
  AND2_X1 U112bar ( .A1(n120bar), .A2(n210bar), .ZN(ybar[0]) );
  OR2_X1 U113 ( .A1(n118), .A2(n186), .ZN(n119) );
  AND2_X1 U113bar ( .A1(n118bar), .A2(n186bar), .ZN(n119bar) );
  AND2_X1 U114 ( .A1(n186), .A2(n118), .ZN(n120) );
  OR2_X1 U114bar ( .A1(n186bar), .A2(n118bar), .ZN(n120bar) );
  AND2_X1 U115 ( .A1(n117), .A2(n116), .ZN(n118) );
  OR2_X1 U115bar ( .A1(n117bar), .A2(n116bar), .ZN(n118bar) );
  OR2_X1 U116 ( .A1(n209), .A2(b[0]), .ZN(n116) );
  AND2_X1 U116bar ( .A1(n209bar), .A2(bbar[0]), .ZN(n116bar) );
  OR2_X1 U117 ( .A1(n201), .A2(a[0]), .ZN(n117) );
  AND2_X1 U117bar ( .A1(n201bar), .A2(abar[0]), .ZN(n117bar) );
  AND2_X1 U118 ( .A1(n114), .A2(n113), .ZN(n115) );
  OR2_X1 U118bar ( .A1(n114bar), .A2(n113bar), .ZN(n115bar) );
  OR2_X1 U119 ( .A1(n185), .A2(d[0]), .ZN(n113) );
  AND2_X1 U119bar ( .A1(n185bar), .A2(dbar[0]), .ZN(n113bar) );
  OR2_X1 U120 ( .A1(n177), .A2(c[0]), .ZN(n114) );
  AND2_X1 U120bar ( .A1(n177bar), .A2(cbar[0]), .ZN(n114bar) );
endmodule

module byteXor4_7 ( a, abar, b, bbar, c, cbar, d, dbar, y, ybar );

  input wire [7:0] a;
  input wire [7:0] b;
  input wire [7:0] c;
  input wire [7:0] d;
  input wire [7:0] abar;
  input wire [7:0] bbar;
  input wire [7:0] cbar;
  input wire [7:0] dbar;
//input_done

  output wire [7:0] y;
  output wire [7:0] ybar;
//output_done

  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n113bar;
  wire n114bar;
  wire n115bar;
  wire n116bar;
  wire n117bar;
  wire n118bar;
  wire n119bar;
  wire n120bar;
  wire n121bar;
  wire n122bar;
  wire n123bar;
  wire n124bar;
  wire n125bar;
  wire n126bar;
  wire n127bar;
  wire n128bar;
  wire n129bar;
  wire n130bar;
  wire n131bar;
  wire n132bar;
  wire n133bar;
  wire n134bar;
  wire n135bar;
  wire n136bar;
  wire n137bar;
  wire n138bar;
  wire n139bar;
  wire n140bar;
  wire n141bar;
  wire n142bar;
  wire n143bar;
  wire n144bar;
  wire n145bar;
  wire n146bar;
  wire n147bar;
  wire n148bar;
  wire n149bar;
  wire n150bar;
  wire n151bar;
  wire n152bar;
  wire n153bar;
  wire n154bar;
  wire n155bar;
  wire n156bar;
  wire n157bar;
  wire n158bar;
  wire n159bar;
  wire n160bar;
  wire n161bar;
  wire n162bar;
  wire n163bar;
  wire n164bar;
  wire n165bar;
  wire n166bar;
  wire n167bar;
  wire n168bar;
  wire n169bar;
  wire n170bar;
  wire n171bar;
  wire n172bar;
  wire n173bar;
  wire n174bar;
  wire n175bar;
  wire n176bar;
  wire n177bar;
  wire n178bar;
  wire n179bar;
  wire n180bar;
  wire n181bar;
  wire n182bar;
  wire n183bar;
  wire n184bar;
  wire n185bar;
  wire n186bar;
  wire n187bar;
  wire n188bar;
  wire n189bar;
  wire n190bar;
  wire n191bar;
  wire n192bar;
  wire n193bar;
  wire n194bar;
  wire n195bar;
  wire n196bar;
  wire n197bar;
  wire n198bar;
  wire n199bar;
  wire n200bar;
  wire n201bar;
  wire n202bar;
  wire n203bar;
  wire n204bar;
  wire n205bar;
  wire n206bar;
  wire n207bar;
  wire n208bar;
  wire n209bar;
  wire n210bar;
  wire n211bar;
  wire n212bar;
  wire n213bar;
  wire n214bar;
  wire n215bar;
  wire n216bar;
  wire n217bar;
  wire n218bar;
  wire n219bar;
  wire n220bar;
  wire n221bar;
  wire n222bar;
  wire n223bar;
  wire n224bar;
//wire_done

 //assign_done

  assign n224bar = n175;
  assign n224 = n175bar;
  assign n223bar = a[7];
  assign n223 = abar[7];
  assign n222bar = n167;
  assign n222 = n167bar;
  assign n221bar = a[6];
  assign n221 = abar[6];
  assign n220bar = n159;
  assign n220 = n159bar;
  assign n219bar = a[5];
  assign n219 = abar[5];
  assign n218bar = n151;
  assign n218 = n151bar;
  assign n217bar = a[4];
  assign n217 = abar[4];
  assign n216bar = n143;
  assign n216 = n143bar;
  assign n215bar = a[3];
  assign n215 = abar[3];
  assign n214bar = n135;
  assign n214 = n135bar;
  assign n213bar = a[2];
  assign n213 = abar[2];
  assign n212bar = n127;
  assign n212 = n127bar;
  assign n211bar = a[1];
  assign n211 = abar[1];
  assign n210bar = n119;
  assign n210 = n119bar;
  assign n209bar = a[0];
  assign n209 = abar[0];
  assign n208bar = b[7];
  assign n208 = bbar[7];
  assign n207bar = b[6];
  assign n207 = bbar[6];
  assign n206bar = b[5];
  assign n206 = bbar[5];
  assign n205bar = b[4];
  assign n205 = bbar[4];
  assign n204bar = b[3];
  assign n204 = bbar[3];
  assign n203bar = b[2];
  assign n203 = bbar[2];
  assign n202bar = b[1];
  assign n202 = bbar[1];
  assign n201bar = b[0];
  assign n201 = bbar[0];
  assign n200bar = n171;
  assign n200 = n171bar;
  assign n199bar = c[7];
  assign n199 = cbar[7];
  assign n198bar = n163;
  assign n198 = n163bar;
  assign n197bar = c[6];
  assign n197 = cbar[6];
  assign n196bar = n155;
  assign n196 = n155bar;
  assign n195bar = c[5];
  assign n195 = cbar[5];
  assign n194bar = n147;
  assign n194 = n147bar;
  assign n193bar = c[4];
  assign n193 = cbar[4];
  assign n192bar = n139;
  assign n192 = n139bar;
  assign n191bar = c[3];
  assign n191 = cbar[3];
  assign n190bar = n131;
  assign n190 = n131bar;
  assign n189bar = c[2];
  assign n189 = cbar[2];
  assign n188bar = n123;
  assign n188 = n123bar;
  assign n187bar = c[1];
  assign n187 = cbar[1];
  assign n186bar = n115;
  assign n186 = n115bar;
  assign n185bar = c[0];
  assign n185 = cbar[0];
  assign n184bar = d[7];
  assign n184 = dbar[7];
  assign n183bar = d[6];
  assign n183 = dbar[6];
  assign n182bar = d[5];
  assign n182 = dbar[5];
  assign n181bar = d[4];
  assign n181 = dbar[4];
  assign n180bar = d[3];
  assign n180 = dbar[3];
  assign n179bar = d[2];
  assign n179 = dbar[2];
  assign n178bar = d[1];
  assign n178 = dbar[1];
  assign n177bar = d[0];
  assign n177 = dbar[0];
  OR2_X1 U49 ( .A1(n176), .A2(n224), .ZN(y[7]) );
  AND2_X1 U49bar ( .A1(n176bar), .A2(n224bar), .ZN(ybar[7]) );
  OR2_X1 U50 ( .A1(n174), .A2(n200), .ZN(n175) );
  AND2_X1 U50bar ( .A1(n174bar), .A2(n200bar), .ZN(n175bar) );
  AND2_X1 U51 ( .A1(n200), .A2(n174), .ZN(n176) );
  OR2_X1 U51bar ( .A1(n200bar), .A2(n174bar), .ZN(n176bar) );
  AND2_X1 U52 ( .A1(n173), .A2(n172), .ZN(n174) );
  OR2_X1 U52bar ( .A1(n173bar), .A2(n172bar), .ZN(n174bar) );
  OR2_X1 U53 ( .A1(n223), .A2(b[7]), .ZN(n172) );
  AND2_X1 U53bar ( .A1(n223bar), .A2(bbar[7]), .ZN(n172bar) );
  OR2_X1 U54 ( .A1(n208), .A2(a[7]), .ZN(n173) );
  AND2_X1 U54bar ( .A1(n208bar), .A2(abar[7]), .ZN(n173bar) );
  AND2_X1 U55 ( .A1(n170), .A2(n169), .ZN(n171) );
  OR2_X1 U55bar ( .A1(n170bar), .A2(n169bar), .ZN(n171bar) );
  OR2_X1 U56 ( .A1(n199), .A2(d[7]), .ZN(n169) );
  AND2_X1 U56bar ( .A1(n199bar), .A2(dbar[7]), .ZN(n169bar) );
  OR2_X1 U57 ( .A1(n184), .A2(c[7]), .ZN(n170) );
  AND2_X1 U57bar ( .A1(n184bar), .A2(cbar[7]), .ZN(n170bar) );
  OR2_X1 U58 ( .A1(n168), .A2(n222), .ZN(y[6]) );
  AND2_X1 U58bar ( .A1(n168bar), .A2(n222bar), .ZN(ybar[6]) );
  OR2_X1 U59 ( .A1(n166), .A2(n198), .ZN(n167) );
  AND2_X1 U59bar ( .A1(n166bar), .A2(n198bar), .ZN(n167bar) );
  AND2_X1 U60 ( .A1(n198), .A2(n166), .ZN(n168) );
  OR2_X1 U60bar ( .A1(n198bar), .A2(n166bar), .ZN(n168bar) );
  AND2_X1 U61 ( .A1(n165), .A2(n164), .ZN(n166) );
  OR2_X1 U61bar ( .A1(n165bar), .A2(n164bar), .ZN(n166bar) );
  OR2_X1 U62 ( .A1(n221), .A2(b[6]), .ZN(n164) );
  AND2_X1 U62bar ( .A1(n221bar), .A2(bbar[6]), .ZN(n164bar) );
  OR2_X1 U63 ( .A1(n207), .A2(a[6]), .ZN(n165) );
  AND2_X1 U63bar ( .A1(n207bar), .A2(abar[6]), .ZN(n165bar) );
  AND2_X1 U64 ( .A1(n162), .A2(n161), .ZN(n163) );
  OR2_X1 U64bar ( .A1(n162bar), .A2(n161bar), .ZN(n163bar) );
  OR2_X1 U65 ( .A1(n197), .A2(d[6]), .ZN(n161) );
  AND2_X1 U65bar ( .A1(n197bar), .A2(dbar[6]), .ZN(n161bar) );
  OR2_X1 U66 ( .A1(n183), .A2(c[6]), .ZN(n162) );
  AND2_X1 U66bar ( .A1(n183bar), .A2(cbar[6]), .ZN(n162bar) );
  OR2_X1 U67 ( .A1(n160), .A2(n220), .ZN(y[5]) );
  AND2_X1 U67bar ( .A1(n160bar), .A2(n220bar), .ZN(ybar[5]) );
  OR2_X1 U68 ( .A1(n158), .A2(n196), .ZN(n159) );
  AND2_X1 U68bar ( .A1(n158bar), .A2(n196bar), .ZN(n159bar) );
  AND2_X1 U69 ( .A1(n196), .A2(n158), .ZN(n160) );
  OR2_X1 U69bar ( .A1(n196bar), .A2(n158bar), .ZN(n160bar) );
  AND2_X1 U70 ( .A1(n157), .A2(n156), .ZN(n158) );
  OR2_X1 U70bar ( .A1(n157bar), .A2(n156bar), .ZN(n158bar) );
  OR2_X1 U71 ( .A1(n219), .A2(b[5]), .ZN(n156) );
  AND2_X1 U71bar ( .A1(n219bar), .A2(bbar[5]), .ZN(n156bar) );
  OR2_X1 U72 ( .A1(n206), .A2(a[5]), .ZN(n157) );
  AND2_X1 U72bar ( .A1(n206bar), .A2(abar[5]), .ZN(n157bar) );
  AND2_X1 U73 ( .A1(n154), .A2(n153), .ZN(n155) );
  OR2_X1 U73bar ( .A1(n154bar), .A2(n153bar), .ZN(n155bar) );
  OR2_X1 U74 ( .A1(n195), .A2(d[5]), .ZN(n153) );
  AND2_X1 U74bar ( .A1(n195bar), .A2(dbar[5]), .ZN(n153bar) );
  OR2_X1 U75 ( .A1(n182), .A2(c[5]), .ZN(n154) );
  AND2_X1 U75bar ( .A1(n182bar), .A2(cbar[5]), .ZN(n154bar) );
  OR2_X1 U76 ( .A1(n152), .A2(n218), .ZN(y[4]) );
  AND2_X1 U76bar ( .A1(n152bar), .A2(n218bar), .ZN(ybar[4]) );
  OR2_X1 U77 ( .A1(n150), .A2(n194), .ZN(n151) );
  AND2_X1 U77bar ( .A1(n150bar), .A2(n194bar), .ZN(n151bar) );
  AND2_X1 U78 ( .A1(n194), .A2(n150), .ZN(n152) );
  OR2_X1 U78bar ( .A1(n194bar), .A2(n150bar), .ZN(n152bar) );
  AND2_X1 U79 ( .A1(n149), .A2(n148), .ZN(n150) );
  OR2_X1 U79bar ( .A1(n149bar), .A2(n148bar), .ZN(n150bar) );
  OR2_X1 U80 ( .A1(n217), .A2(b[4]), .ZN(n148) );
  AND2_X1 U80bar ( .A1(n217bar), .A2(bbar[4]), .ZN(n148bar) );
  OR2_X1 U81 ( .A1(n205), .A2(a[4]), .ZN(n149) );
  AND2_X1 U81bar ( .A1(n205bar), .A2(abar[4]), .ZN(n149bar) );
  AND2_X1 U82 ( .A1(n146), .A2(n145), .ZN(n147) );
  OR2_X1 U82bar ( .A1(n146bar), .A2(n145bar), .ZN(n147bar) );
  OR2_X1 U83 ( .A1(n193), .A2(d[4]), .ZN(n145) );
  AND2_X1 U83bar ( .A1(n193bar), .A2(dbar[4]), .ZN(n145bar) );
  OR2_X1 U84 ( .A1(n181), .A2(c[4]), .ZN(n146) );
  AND2_X1 U84bar ( .A1(n181bar), .A2(cbar[4]), .ZN(n146bar) );
  OR2_X1 U85 ( .A1(n144), .A2(n216), .ZN(y[3]) );
  AND2_X1 U85bar ( .A1(n144bar), .A2(n216bar), .ZN(ybar[3]) );
  OR2_X1 U86 ( .A1(n142), .A2(n192), .ZN(n143) );
  AND2_X1 U86bar ( .A1(n142bar), .A2(n192bar), .ZN(n143bar) );
  AND2_X1 U87 ( .A1(n192), .A2(n142), .ZN(n144) );
  OR2_X1 U87bar ( .A1(n192bar), .A2(n142bar), .ZN(n144bar) );
  AND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(n142) );
  OR2_X1 U88bar ( .A1(n141bar), .A2(n140bar), .ZN(n142bar) );
  OR2_X1 U89 ( .A1(n215), .A2(b[3]), .ZN(n140) );
  AND2_X1 U89bar ( .A1(n215bar), .A2(bbar[3]), .ZN(n140bar) );
  OR2_X1 U90 ( .A1(n204), .A2(a[3]), .ZN(n141) );
  AND2_X1 U90bar ( .A1(n204bar), .A2(abar[3]), .ZN(n141bar) );
  AND2_X1 U91 ( .A1(n138), .A2(n137), .ZN(n139) );
  OR2_X1 U91bar ( .A1(n138bar), .A2(n137bar), .ZN(n139bar) );
  OR2_X1 U92 ( .A1(n191), .A2(d[3]), .ZN(n137) );
  AND2_X1 U92bar ( .A1(n191bar), .A2(dbar[3]), .ZN(n137bar) );
  OR2_X1 U93 ( .A1(n180), .A2(c[3]), .ZN(n138) );
  AND2_X1 U93bar ( .A1(n180bar), .A2(cbar[3]), .ZN(n138bar) );
  OR2_X1 U94 ( .A1(n136), .A2(n214), .ZN(y[2]) );
  AND2_X1 U94bar ( .A1(n136bar), .A2(n214bar), .ZN(ybar[2]) );
  OR2_X1 U95 ( .A1(n134), .A2(n190), .ZN(n135) );
  AND2_X1 U95bar ( .A1(n134bar), .A2(n190bar), .ZN(n135bar) );
  AND2_X1 U96 ( .A1(n190), .A2(n134), .ZN(n136) );
  OR2_X1 U96bar ( .A1(n190bar), .A2(n134bar), .ZN(n136bar) );
  AND2_X1 U97 ( .A1(n133), .A2(n132), .ZN(n134) );
  OR2_X1 U97bar ( .A1(n133bar), .A2(n132bar), .ZN(n134bar) );
  OR2_X1 U98 ( .A1(n213), .A2(b[2]), .ZN(n132) );
  AND2_X1 U98bar ( .A1(n213bar), .A2(bbar[2]), .ZN(n132bar) );
  OR2_X1 U99 ( .A1(n203), .A2(a[2]), .ZN(n133) );
  AND2_X1 U99bar ( .A1(n203bar), .A2(abar[2]), .ZN(n133bar) );
  AND2_X1 U100 ( .A1(n130), .A2(n129), .ZN(n131) );
  OR2_X1 U100bar ( .A1(n130bar), .A2(n129bar), .ZN(n131bar) );
  OR2_X1 U101 ( .A1(n189), .A2(d[2]), .ZN(n129) );
  AND2_X1 U101bar ( .A1(n189bar), .A2(dbar[2]), .ZN(n129bar) );
  OR2_X1 U102 ( .A1(n179), .A2(c[2]), .ZN(n130) );
  AND2_X1 U102bar ( .A1(n179bar), .A2(cbar[2]), .ZN(n130bar) );
  OR2_X1 U103 ( .A1(n128), .A2(n212), .ZN(y[1]) );
  AND2_X1 U103bar ( .A1(n128bar), .A2(n212bar), .ZN(ybar[1]) );
  OR2_X1 U104 ( .A1(n126), .A2(n188), .ZN(n127) );
  AND2_X1 U104bar ( .A1(n126bar), .A2(n188bar), .ZN(n127bar) );
  AND2_X1 U105 ( .A1(n188), .A2(n126), .ZN(n128) );
  OR2_X1 U105bar ( .A1(n188bar), .A2(n126bar), .ZN(n128bar) );
  AND2_X1 U106 ( .A1(n125), .A2(n124), .ZN(n126) );
  OR2_X1 U106bar ( .A1(n125bar), .A2(n124bar), .ZN(n126bar) );
  OR2_X1 U107 ( .A1(n211), .A2(b[1]), .ZN(n124) );
  AND2_X1 U107bar ( .A1(n211bar), .A2(bbar[1]), .ZN(n124bar) );
  OR2_X1 U108 ( .A1(n202), .A2(a[1]), .ZN(n125) );
  AND2_X1 U108bar ( .A1(n202bar), .A2(abar[1]), .ZN(n125bar) );
  AND2_X1 U109 ( .A1(n122), .A2(n121), .ZN(n123) );
  OR2_X1 U109bar ( .A1(n122bar), .A2(n121bar), .ZN(n123bar) );
  OR2_X1 U110 ( .A1(n187), .A2(d[1]), .ZN(n121) );
  AND2_X1 U110bar ( .A1(n187bar), .A2(dbar[1]), .ZN(n121bar) );
  OR2_X1 U111 ( .A1(n178), .A2(c[1]), .ZN(n122) );
  AND2_X1 U111bar ( .A1(n178bar), .A2(cbar[1]), .ZN(n122bar) );
  OR2_X1 U112 ( .A1(n120), .A2(n210), .ZN(y[0]) );
  AND2_X1 U112bar ( .A1(n120bar), .A2(n210bar), .ZN(ybar[0]) );
  OR2_X1 U113 ( .A1(n118), .A2(n186), .ZN(n119) );
  AND2_X1 U113bar ( .A1(n118bar), .A2(n186bar), .ZN(n119bar) );
  AND2_X1 U114 ( .A1(n186), .A2(n118), .ZN(n120) );
  OR2_X1 U114bar ( .A1(n186bar), .A2(n118bar), .ZN(n120bar) );
  AND2_X1 U115 ( .A1(n117), .A2(n116), .ZN(n118) );
  OR2_X1 U115bar ( .A1(n117bar), .A2(n116bar), .ZN(n118bar) );
  OR2_X1 U116 ( .A1(n209), .A2(b[0]), .ZN(n116) );
  AND2_X1 U116bar ( .A1(n209bar), .A2(bbar[0]), .ZN(n116bar) );
  OR2_X1 U117 ( .A1(n201), .A2(a[0]), .ZN(n117) );
  AND2_X1 U117bar ( .A1(n201bar), .A2(abar[0]), .ZN(n117bar) );
  AND2_X1 U118 ( .A1(n114), .A2(n113), .ZN(n115) );
  OR2_X1 U118bar ( .A1(n114bar), .A2(n113bar), .ZN(n115bar) );
  OR2_X1 U119 ( .A1(n185), .A2(d[0]), .ZN(n113) );
  AND2_X1 U119bar ( .A1(n185bar), .A2(dbar[0]), .ZN(n113bar) );
  OR2_X1 U120 ( .A1(n177), .A2(c[0]), .ZN(n114) );
  AND2_X1 U120bar ( .A1(n177bar), .A2(cbar[0]), .ZN(n114bar) );
endmodule

module byteXor4_8 ( a, abar, b, bbar, c, cbar, d, dbar, y, ybar );

  input wire [7:0] a;
  input wire [7:0] b;
  input wire [7:0] c;
  input wire [7:0] d;
  input wire [7:0] abar;
  input wire [7:0] bbar;
  input wire [7:0] cbar;
  input wire [7:0] dbar;
//input_done

  output wire [7:0] y;
  output wire [7:0] ybar;
//output_done

  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n113bar;
  wire n114bar;
  wire n115bar;
  wire n116bar;
  wire n117bar;
  wire n118bar;
  wire n119bar;
  wire n120bar;
  wire n121bar;
  wire n122bar;
  wire n123bar;
  wire n124bar;
  wire n125bar;
  wire n126bar;
  wire n127bar;
  wire n128bar;
  wire n129bar;
  wire n130bar;
  wire n131bar;
  wire n132bar;
  wire n133bar;
  wire n134bar;
  wire n135bar;
  wire n136bar;
  wire n137bar;
  wire n138bar;
  wire n139bar;
  wire n140bar;
  wire n141bar;
  wire n142bar;
  wire n143bar;
  wire n144bar;
  wire n145bar;
  wire n146bar;
  wire n147bar;
  wire n148bar;
  wire n149bar;
  wire n150bar;
  wire n151bar;
  wire n152bar;
  wire n153bar;
  wire n154bar;
  wire n155bar;
  wire n156bar;
  wire n157bar;
  wire n158bar;
  wire n159bar;
  wire n160bar;
  wire n161bar;
  wire n162bar;
  wire n163bar;
  wire n164bar;
  wire n165bar;
  wire n166bar;
  wire n167bar;
  wire n168bar;
  wire n169bar;
  wire n170bar;
  wire n171bar;
  wire n172bar;
  wire n173bar;
  wire n174bar;
  wire n175bar;
  wire n176bar;
  wire n177bar;
  wire n178bar;
  wire n179bar;
  wire n180bar;
  wire n181bar;
  wire n182bar;
  wire n183bar;
  wire n184bar;
  wire n185bar;
  wire n186bar;
  wire n187bar;
  wire n188bar;
  wire n189bar;
  wire n190bar;
  wire n191bar;
  wire n192bar;
  wire n193bar;
  wire n194bar;
  wire n195bar;
  wire n196bar;
  wire n197bar;
  wire n198bar;
  wire n199bar;
  wire n200bar;
  wire n201bar;
  wire n202bar;
  wire n203bar;
  wire n204bar;
  wire n205bar;
  wire n206bar;
  wire n207bar;
  wire n208bar;
  wire n209bar;
  wire n210bar;
  wire n211bar;
  wire n212bar;
  wire n213bar;
  wire n214bar;
  wire n215bar;
  wire n216bar;
  wire n217bar;
  wire n218bar;
  wire n219bar;
  wire n220bar;
  wire n221bar;
  wire n222bar;
  wire n223bar;
  wire n224bar;
//wire_done

 //assign_done

  assign n224bar = n175;
  assign n224 = n175bar;
  assign n223bar = a[7];
  assign n223 = abar[7];
  assign n222bar = n167;
  assign n222 = n167bar;
  assign n221bar = a[6];
  assign n221 = abar[6];
  assign n220bar = n159;
  assign n220 = n159bar;
  assign n219bar = a[5];
  assign n219 = abar[5];
  assign n218bar = n151;
  assign n218 = n151bar;
  assign n217bar = a[4];
  assign n217 = abar[4];
  assign n216bar = n143;
  assign n216 = n143bar;
  assign n215bar = a[3];
  assign n215 = abar[3];
  assign n214bar = n135;
  assign n214 = n135bar;
  assign n213bar = a[2];
  assign n213 = abar[2];
  assign n212bar = n127;
  assign n212 = n127bar;
  assign n211bar = a[1];
  assign n211 = abar[1];
  assign n210bar = n119;
  assign n210 = n119bar;
  assign n209bar = a[0];
  assign n209 = abar[0];
  assign n208bar = b[7];
  assign n208 = bbar[7];
  assign n207bar = b[6];
  assign n207 = bbar[6];
  assign n206bar = b[5];
  assign n206 = bbar[5];
  assign n205bar = b[4];
  assign n205 = bbar[4];
  assign n204bar = b[3];
  assign n204 = bbar[3];
  assign n203bar = b[2];
  assign n203 = bbar[2];
  assign n202bar = b[1];
  assign n202 = bbar[1];
  assign n201bar = b[0];
  assign n201 = bbar[0];
  assign n200bar = n171;
  assign n200 = n171bar;
  assign n199bar = c[7];
  assign n199 = cbar[7];
  assign n198bar = n163;
  assign n198 = n163bar;
  assign n197bar = c[6];
  assign n197 = cbar[6];
  assign n196bar = n155;
  assign n196 = n155bar;
  assign n195bar = c[5];
  assign n195 = cbar[5];
  assign n194bar = n147;
  assign n194 = n147bar;
  assign n193bar = c[4];
  assign n193 = cbar[4];
  assign n192bar = n139;
  assign n192 = n139bar;
  assign n191bar = c[3];
  assign n191 = cbar[3];
  assign n190bar = n131;
  assign n190 = n131bar;
  assign n189bar = c[2];
  assign n189 = cbar[2];
  assign n188bar = n123;
  assign n188 = n123bar;
  assign n187bar = c[1];
  assign n187 = cbar[1];
  assign n186bar = n115;
  assign n186 = n115bar;
  assign n185bar = c[0];
  assign n185 = cbar[0];
  assign n184bar = d[7];
  assign n184 = dbar[7];
  assign n183bar = d[6];
  assign n183 = dbar[6];
  assign n182bar = d[5];
  assign n182 = dbar[5];
  assign n181bar = d[4];
  assign n181 = dbar[4];
  assign n180bar = d[3];
  assign n180 = dbar[3];
  assign n179bar = d[2];
  assign n179 = dbar[2];
  assign n178bar = d[1];
  assign n178 = dbar[1];
  assign n177bar = d[0];
  assign n177 = dbar[0];
  OR2_X1 U49 ( .A1(n176), .A2(n224), .ZN(y[7]) );
  AND2_X1 U49bar ( .A1(n176bar), .A2(n224bar), .ZN(ybar[7]) );
  OR2_X1 U50 ( .A1(n174), .A2(n200), .ZN(n175) );
  AND2_X1 U50bar ( .A1(n174bar), .A2(n200bar), .ZN(n175bar) );
  AND2_X1 U51 ( .A1(n200), .A2(n174), .ZN(n176) );
  OR2_X1 U51bar ( .A1(n200bar), .A2(n174bar), .ZN(n176bar) );
  AND2_X1 U52 ( .A1(n173), .A2(n172), .ZN(n174) );
  OR2_X1 U52bar ( .A1(n173bar), .A2(n172bar), .ZN(n174bar) );
  OR2_X1 U53 ( .A1(n223), .A2(b[7]), .ZN(n172) );
  AND2_X1 U53bar ( .A1(n223bar), .A2(bbar[7]), .ZN(n172bar) );
  OR2_X1 U54 ( .A1(n208), .A2(a[7]), .ZN(n173) );
  AND2_X1 U54bar ( .A1(n208bar), .A2(abar[7]), .ZN(n173bar) );
  AND2_X1 U55 ( .A1(n170), .A2(n169), .ZN(n171) );
  OR2_X1 U55bar ( .A1(n170bar), .A2(n169bar), .ZN(n171bar) );
  OR2_X1 U56 ( .A1(n199), .A2(d[7]), .ZN(n169) );
  AND2_X1 U56bar ( .A1(n199bar), .A2(dbar[7]), .ZN(n169bar) );
  OR2_X1 U57 ( .A1(n184), .A2(c[7]), .ZN(n170) );
  AND2_X1 U57bar ( .A1(n184bar), .A2(cbar[7]), .ZN(n170bar) );
  OR2_X1 U58 ( .A1(n168), .A2(n222), .ZN(y[6]) );
  AND2_X1 U58bar ( .A1(n168bar), .A2(n222bar), .ZN(ybar[6]) );
  OR2_X1 U59 ( .A1(n166), .A2(n198), .ZN(n167) );
  AND2_X1 U59bar ( .A1(n166bar), .A2(n198bar), .ZN(n167bar) );
  AND2_X1 U60 ( .A1(n198), .A2(n166), .ZN(n168) );
  OR2_X1 U60bar ( .A1(n198bar), .A2(n166bar), .ZN(n168bar) );
  AND2_X1 U61 ( .A1(n165), .A2(n164), .ZN(n166) );
  OR2_X1 U61bar ( .A1(n165bar), .A2(n164bar), .ZN(n166bar) );
  OR2_X1 U62 ( .A1(n221), .A2(b[6]), .ZN(n164) );
  AND2_X1 U62bar ( .A1(n221bar), .A2(bbar[6]), .ZN(n164bar) );
  OR2_X1 U63 ( .A1(n207), .A2(a[6]), .ZN(n165) );
  AND2_X1 U63bar ( .A1(n207bar), .A2(abar[6]), .ZN(n165bar) );
  AND2_X1 U64 ( .A1(n162), .A2(n161), .ZN(n163) );
  OR2_X1 U64bar ( .A1(n162bar), .A2(n161bar), .ZN(n163bar) );
  OR2_X1 U65 ( .A1(n197), .A2(d[6]), .ZN(n161) );
  AND2_X1 U65bar ( .A1(n197bar), .A2(dbar[6]), .ZN(n161bar) );
  OR2_X1 U66 ( .A1(n183), .A2(c[6]), .ZN(n162) );
  AND2_X1 U66bar ( .A1(n183bar), .A2(cbar[6]), .ZN(n162bar) );
  OR2_X1 U67 ( .A1(n160), .A2(n220), .ZN(y[5]) );
  AND2_X1 U67bar ( .A1(n160bar), .A2(n220bar), .ZN(ybar[5]) );
  OR2_X1 U68 ( .A1(n158), .A2(n196), .ZN(n159) );
  AND2_X1 U68bar ( .A1(n158bar), .A2(n196bar), .ZN(n159bar) );
  AND2_X1 U69 ( .A1(n196), .A2(n158), .ZN(n160) );
  OR2_X1 U69bar ( .A1(n196bar), .A2(n158bar), .ZN(n160bar) );
  AND2_X1 U70 ( .A1(n157), .A2(n156), .ZN(n158) );
  OR2_X1 U70bar ( .A1(n157bar), .A2(n156bar), .ZN(n158bar) );
  OR2_X1 U71 ( .A1(n219), .A2(b[5]), .ZN(n156) );
  AND2_X1 U71bar ( .A1(n219bar), .A2(bbar[5]), .ZN(n156bar) );
  OR2_X1 U72 ( .A1(n206), .A2(a[5]), .ZN(n157) );
  AND2_X1 U72bar ( .A1(n206bar), .A2(abar[5]), .ZN(n157bar) );
  AND2_X1 U73 ( .A1(n154), .A2(n153), .ZN(n155) );
  OR2_X1 U73bar ( .A1(n154bar), .A2(n153bar), .ZN(n155bar) );
  OR2_X1 U74 ( .A1(n195), .A2(d[5]), .ZN(n153) );
  AND2_X1 U74bar ( .A1(n195bar), .A2(dbar[5]), .ZN(n153bar) );
  OR2_X1 U75 ( .A1(n182), .A2(c[5]), .ZN(n154) );
  AND2_X1 U75bar ( .A1(n182bar), .A2(cbar[5]), .ZN(n154bar) );
  OR2_X1 U76 ( .A1(n152), .A2(n218), .ZN(y[4]) );
  AND2_X1 U76bar ( .A1(n152bar), .A2(n218bar), .ZN(ybar[4]) );
  OR2_X1 U77 ( .A1(n150), .A2(n194), .ZN(n151) );
  AND2_X1 U77bar ( .A1(n150bar), .A2(n194bar), .ZN(n151bar) );
  AND2_X1 U78 ( .A1(n194), .A2(n150), .ZN(n152) );
  OR2_X1 U78bar ( .A1(n194bar), .A2(n150bar), .ZN(n152bar) );
  AND2_X1 U79 ( .A1(n149), .A2(n148), .ZN(n150) );
  OR2_X1 U79bar ( .A1(n149bar), .A2(n148bar), .ZN(n150bar) );
  OR2_X1 U80 ( .A1(n217), .A2(b[4]), .ZN(n148) );
  AND2_X1 U80bar ( .A1(n217bar), .A2(bbar[4]), .ZN(n148bar) );
  OR2_X1 U81 ( .A1(n205), .A2(a[4]), .ZN(n149) );
  AND2_X1 U81bar ( .A1(n205bar), .A2(abar[4]), .ZN(n149bar) );
  AND2_X1 U82 ( .A1(n146), .A2(n145), .ZN(n147) );
  OR2_X1 U82bar ( .A1(n146bar), .A2(n145bar), .ZN(n147bar) );
  OR2_X1 U83 ( .A1(n193), .A2(d[4]), .ZN(n145) );
  AND2_X1 U83bar ( .A1(n193bar), .A2(dbar[4]), .ZN(n145bar) );
  OR2_X1 U84 ( .A1(n181), .A2(c[4]), .ZN(n146) );
  AND2_X1 U84bar ( .A1(n181bar), .A2(cbar[4]), .ZN(n146bar) );
  OR2_X1 U85 ( .A1(n144), .A2(n216), .ZN(y[3]) );
  AND2_X1 U85bar ( .A1(n144bar), .A2(n216bar), .ZN(ybar[3]) );
  OR2_X1 U86 ( .A1(n142), .A2(n192), .ZN(n143) );
  AND2_X1 U86bar ( .A1(n142bar), .A2(n192bar), .ZN(n143bar) );
  AND2_X1 U87 ( .A1(n192), .A2(n142), .ZN(n144) );
  OR2_X1 U87bar ( .A1(n192bar), .A2(n142bar), .ZN(n144bar) );
  AND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(n142) );
  OR2_X1 U88bar ( .A1(n141bar), .A2(n140bar), .ZN(n142bar) );
  OR2_X1 U89 ( .A1(n215), .A2(b[3]), .ZN(n140) );
  AND2_X1 U89bar ( .A1(n215bar), .A2(bbar[3]), .ZN(n140bar) );
  OR2_X1 U90 ( .A1(n204), .A2(a[3]), .ZN(n141) );
  AND2_X1 U90bar ( .A1(n204bar), .A2(abar[3]), .ZN(n141bar) );
  AND2_X1 U91 ( .A1(n138), .A2(n137), .ZN(n139) );
  OR2_X1 U91bar ( .A1(n138bar), .A2(n137bar), .ZN(n139bar) );
  OR2_X1 U92 ( .A1(n191), .A2(d[3]), .ZN(n137) );
  AND2_X1 U92bar ( .A1(n191bar), .A2(dbar[3]), .ZN(n137bar) );
  OR2_X1 U93 ( .A1(n180), .A2(c[3]), .ZN(n138) );
  AND2_X1 U93bar ( .A1(n180bar), .A2(cbar[3]), .ZN(n138bar) );
  OR2_X1 U94 ( .A1(n136), .A2(n214), .ZN(y[2]) );
  AND2_X1 U94bar ( .A1(n136bar), .A2(n214bar), .ZN(ybar[2]) );
  OR2_X1 U95 ( .A1(n134), .A2(n190), .ZN(n135) );
  AND2_X1 U95bar ( .A1(n134bar), .A2(n190bar), .ZN(n135bar) );
  AND2_X1 U96 ( .A1(n190), .A2(n134), .ZN(n136) );
  OR2_X1 U96bar ( .A1(n190bar), .A2(n134bar), .ZN(n136bar) );
  AND2_X1 U97 ( .A1(n133), .A2(n132), .ZN(n134) );
  OR2_X1 U97bar ( .A1(n133bar), .A2(n132bar), .ZN(n134bar) );
  OR2_X1 U98 ( .A1(n213), .A2(b[2]), .ZN(n132) );
  AND2_X1 U98bar ( .A1(n213bar), .A2(bbar[2]), .ZN(n132bar) );
  OR2_X1 U99 ( .A1(n203), .A2(a[2]), .ZN(n133) );
  AND2_X1 U99bar ( .A1(n203bar), .A2(abar[2]), .ZN(n133bar) );
  AND2_X1 U100 ( .A1(n130), .A2(n129), .ZN(n131) );
  OR2_X1 U100bar ( .A1(n130bar), .A2(n129bar), .ZN(n131bar) );
  OR2_X1 U101 ( .A1(n189), .A2(d[2]), .ZN(n129) );
  AND2_X1 U101bar ( .A1(n189bar), .A2(dbar[2]), .ZN(n129bar) );
  OR2_X1 U102 ( .A1(n179), .A2(c[2]), .ZN(n130) );
  AND2_X1 U102bar ( .A1(n179bar), .A2(cbar[2]), .ZN(n130bar) );
  OR2_X1 U103 ( .A1(n128), .A2(n212), .ZN(y[1]) );
  AND2_X1 U103bar ( .A1(n128bar), .A2(n212bar), .ZN(ybar[1]) );
  OR2_X1 U104 ( .A1(n126), .A2(n188), .ZN(n127) );
  AND2_X1 U104bar ( .A1(n126bar), .A2(n188bar), .ZN(n127bar) );
  AND2_X1 U105 ( .A1(n188), .A2(n126), .ZN(n128) );
  OR2_X1 U105bar ( .A1(n188bar), .A2(n126bar), .ZN(n128bar) );
  AND2_X1 U106 ( .A1(n125), .A2(n124), .ZN(n126) );
  OR2_X1 U106bar ( .A1(n125bar), .A2(n124bar), .ZN(n126bar) );
  OR2_X1 U107 ( .A1(n211), .A2(b[1]), .ZN(n124) );
  AND2_X1 U107bar ( .A1(n211bar), .A2(bbar[1]), .ZN(n124bar) );
  OR2_X1 U108 ( .A1(n202), .A2(a[1]), .ZN(n125) );
  AND2_X1 U108bar ( .A1(n202bar), .A2(abar[1]), .ZN(n125bar) );
  AND2_X1 U109 ( .A1(n122), .A2(n121), .ZN(n123) );
  OR2_X1 U109bar ( .A1(n122bar), .A2(n121bar), .ZN(n123bar) );
  OR2_X1 U110 ( .A1(n187), .A2(d[1]), .ZN(n121) );
  AND2_X1 U110bar ( .A1(n187bar), .A2(dbar[1]), .ZN(n121bar) );
  OR2_X1 U111 ( .A1(n178), .A2(c[1]), .ZN(n122) );
  AND2_X1 U111bar ( .A1(n178bar), .A2(cbar[1]), .ZN(n122bar) );
  OR2_X1 U112 ( .A1(n120), .A2(n210), .ZN(y[0]) );
  AND2_X1 U112bar ( .A1(n120bar), .A2(n210bar), .ZN(ybar[0]) );
  OR2_X1 U113 ( .A1(n118), .A2(n186), .ZN(n119) );
  AND2_X1 U113bar ( .A1(n118bar), .A2(n186bar), .ZN(n119bar) );
  AND2_X1 U114 ( .A1(n186), .A2(n118), .ZN(n120) );
  OR2_X1 U114bar ( .A1(n186bar), .A2(n118bar), .ZN(n120bar) );
  AND2_X1 U115 ( .A1(n117), .A2(n116), .ZN(n118) );
  OR2_X1 U115bar ( .A1(n117bar), .A2(n116bar), .ZN(n118bar) );
  OR2_X1 U116 ( .A1(n209), .A2(b[0]), .ZN(n116) );
  AND2_X1 U116bar ( .A1(n209bar), .A2(bbar[0]), .ZN(n116bar) );
  OR2_X1 U117 ( .A1(n201), .A2(a[0]), .ZN(n117) );
  AND2_X1 U117bar ( .A1(n201bar), .A2(abar[0]), .ZN(n117bar) );
  AND2_X1 U118 ( .A1(n114), .A2(n113), .ZN(n115) );
  OR2_X1 U118bar ( .A1(n114bar), .A2(n113bar), .ZN(n115bar) );
  OR2_X1 U119 ( .A1(n185), .A2(d[0]), .ZN(n113) );
  AND2_X1 U119bar ( .A1(n185bar), .A2(dbar[0]), .ZN(n113bar) );
  OR2_X1 U120 ( .A1(n177), .A2(c[0]), .ZN(n114) );
  AND2_X1 U120bar ( .A1(n177bar), .A2(cbar[0]), .ZN(n114bar) );
endmodule

module mixCol_2 ( in, inbar, out, outbar );

  input wire [31:0] in;
  input wire [31:0] inbar;
//input_done

  output wire [31:0] out;
  output wire [31:0] outbar;
//output_done

  wire [7:0] b0_s2;
  wire [7:0] b1_s2;
  wire [7:0] b2_s2;
  wire [7:0] b3_s2;
  wire [7:0] b0_s3;
  wire [7:0] b1_s3;
  wire [7:0] b2_s3;
  wire [7:0] b3_s3;

  wire [7:0] b0_s2bar;
  wire [7:0] b1_s2bar;
  wire [7:0] b2_s2bar;
  wire [7:0] b3_s2bar;
  wire [7:0] b0_s3bar;
  wire [7:0] b1_s3bar;
  wire [7:0] b2_s3bar;
  wire [7:0] b3_s3bar;
//wire_done

 //assign_done

  scale2_8 b0_scale2 ( .in(in[31:24]), .inbar(inbar[31:24]), .out(b0_s2), .outbar(b0_s2bar) );
  scale2_7 b1_scale2 ( .in(in[23:16]), .inbar(inbar[23:16]), .out(b1_s2), .outbar(b1_s2bar) );
  scale2_6 b2_scale2 ( .in(in[15:8]), .inbar(inbar[15:8]), .out(b2_s2), .outbar(b2_s2bar) );
  scale2_5 b3_scale2 ( .in(in[7:0]), .inbar(inbar[7:0]), .out(b3_s2), .outbar(b3_s2bar) );

  byteXor_9 b0_scale3 ( .a(in[31:24]), .abar(inbar[31:24]), .b(b0_s2), .bbar(b0_s2bar), .y(b0_s3), .ybar(b0_s3bar) );
  byteXor_8 b1_scale3 ( .a(in[23:16]), .abar(inbar[23:16]), .b(b1_s2), .bbar(b1_s2bar), .y(b1_s3), .ybar(b1_s3bar) );
  byteXor_7 b2_scale3 ( .a(in[15:8]), .abar(inbar[15:8]), .b(b2_s2), .bbar(b2_s2bar), .y(b2_s3), .ybar(b2_s3bar) );
  byteXor_6 b3_scale3 ( .a(in[7:0]), .abar(inbar[7:0]), .b(b3_s2), .bbar(b3_s2bar), .y(b3_s3), .ybar(b3_s3bar) );

  byteXor4_8 out0 ( .a(b0_s2), .abar(b0_s2bar), .b(b1_s3), .bbar(b1_s3bar), .c(in[15:8]), .cbar(inbar[15:8]),
       .d(in[7:0]), .dbar(inbar[7:0]), .y(out[31:24]), .ybar(outbar[31:24]) );
  byteXor4_7 out1 ( .a(in[31:24]), .abar(inbar[31:24]), .b(b1_s2), .bbar(b1_s2bar), .c(b2_s3), .cbar(b2_s3bar),
       .d(in[7:0]), .dbar(inbar[7:0]), .y(out[23:16]), .ybar(outbar[23:16]) );
  byteXor4_6 out2 ( .a(in[31:24]), .abar(inbar[31:24]), .b(in[23:16]), .bbar(inbar[23:16]), .c(b2_s2), .cbar(b2_s2bar),
       .d(b3_s3), .dbar(b3_s3bar), .y(out[15:8]), .ybar(outbar[15:8]) );
  byteXor4_5 out3 ( .a(b0_s3), .abar(b0_s3bar), .b(in[23:16]), .bbar(inbar[23:16]), .c(in[15:8]), .cbar(inbar[15:8]),
       .d(b3_s2), .dbar(b3_s2bar), .y(out[7:0]), .ybar(outbar[7:0]) );
endmodule

module scale2_9 ( in, inbar, out, outbar );

  input wire [7:0] in;
  input wire [7:0] inbar;
//input_done

  output wire [7:0] out;
  output wire [7:0] outbar;
//output_done

  wire in_0;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_1;
  wire in_7;
  wire n11;
  wire n12;
  wire n13;
  wire n14;
  wire n15;
  wire n16;
  wire n17;
  wire n18;
  wire n19;
  wire n20;
  wire in_0bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_1bar;
  wire in_7bar;
  wire n11bar;
  wire n12bar;
  wire n13bar;
  wire n14bar;
  wire n15bar;
  wire n16bar;
  wire n17bar;
  wire n18bar;
  wire n19bar;
  wire n20bar;
//wire_done

  assign in_0 = in[0];
  assign out[7] = in_6;
  assign in_6  = in[6];
  assign out[6] = in_5;
  assign in_5  = in[5];
  assign out[5] = in_4;
  assign in_4  = in[4];
  assign out[2] = in_1;
  assign in_1  = in[1];
  assign out[0] = in_7;
  assign in_7  = in[7];
  assign in_0bar = inbar[0];
  assign outbar[7] = in_6bar;
  assign in_6bar = inbar[6];
  assign outbar[6] = in_5bar;
  assign in_5bar = inbar[5];
  assign outbar[5] = in_4bar;
  assign in_4bar = inbar[4];
  assign outbar[2] = in_1bar;
  assign in_1bar = inbar[1];
  assign outbar[0] = in_7bar;
  assign in_7bar = inbar[7];
//assign_done

  assign n20bar = in_7;
  assign n20 = in_7bar;
  assign n19bar = in[3];
  assign n19 = inbar[3];
  assign n18bar = in[2];
  assign n18 = inbar[2];
  assign n17bar = in_0;
  assign n17 = in_0bar;
  OR2_X1 U5 ( .A1(n16), .A2(n15), .ZN(out[4]) );
  AND2_X1 U5bar ( .A1(n16bar), .A2(n15bar), .ZN(outbar[4]) );
  AND2_X1 U6 ( .A1(in[3]), .A2(n20), .ZN(n15) );
  OR2_X1 U6bar ( .A1(inbar[3]), .A2(n20bar), .ZN(n15bar) );
  AND2_X1 U7 ( .A1(in_7), .A2(n19), .ZN(n16) );
  OR2_X1 U7bar ( .A1(in_7bar), .A2(n19bar), .ZN(n16bar) );
  OR2_X1 U8 ( .A1(n14), .A2(n13), .ZN(out[3]) );
  AND2_X1 U8bar ( .A1(n14bar), .A2(n13bar), .ZN(outbar[3]) );
  AND2_X1 U9 ( .A1(in[2]), .A2(n20), .ZN(n13) );
  OR2_X1 U9bar ( .A1(inbar[2]), .A2(n20bar), .ZN(n13bar) );
  AND2_X1 U10 ( .A1(in_7), .A2(n18), .ZN(n14) );
  OR2_X1 U10bar ( .A1(in_7bar), .A2(n18bar), .ZN(n14bar) );
  OR2_X1 U11 ( .A1(n12), .A2(n11), .ZN(out[1]) );
  AND2_X1 U11bar ( .A1(n12bar), .A2(n11bar), .ZN(outbar[1]) );
  AND2_X1 U12 ( .A1(in_0), .A2(n20), .ZN(n11) );
  OR2_X1 U12bar ( .A1(in_0bar), .A2(n20bar), .ZN(n11bar) );
  AND2_X1 U13 ( .A1(in_7), .A2(n17), .ZN(n12) );
  OR2_X1 U13bar ( .A1(in_7bar), .A2(n17bar), .ZN(n12bar) );
endmodule

module scale2_10 ( in, inbar, out, outbar );

  input wire [7:0] in;
  input wire [7:0] inbar;
//input_done

  output wire [7:0] out;
  output wire [7:0] outbar;
//output_done

  wire in_0;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_1;
  wire in_7;
  wire n11;
  wire n12;
  wire n13;
  wire n14;
  wire n15;
  wire n16;
  wire n17;
  wire n18;
  wire n19;
  wire n20;
  wire in_0bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_1bar;
  wire in_7bar;
  wire n11bar;
  wire n12bar;
  wire n13bar;
  wire n14bar;
  wire n15bar;
  wire n16bar;
  wire n17bar;
  wire n18bar;
  wire n19bar;
  wire n20bar;
//wire_done

  assign in_0 = in[0];
  assign out[7] = in_6;
  assign in_6  = in[6];
  assign out[6] = in_5;
  assign in_5  = in[5];
  assign out[5] = in_4;
  assign in_4  = in[4];
  assign out[2] = in_1;
  assign in_1  = in[1];
  assign out[0] = in_7;
  assign in_7  = in[7];
  assign in_0bar = inbar[0];
  assign outbar[7] = in_6bar;
  assign in_6bar = inbar[6];
  assign outbar[6] = in_5bar;
  assign in_5bar = inbar[5];
  assign outbar[5] = in_4bar;
  assign in_4bar = inbar[4];
  assign outbar[2] = in_1bar;
  assign in_1bar = inbar[1];
  assign outbar[0] = in_7bar;
  assign in_7bar = inbar[7];
//assign_done

  assign n20bar = in_7;
  assign n20 = in_7bar;
  assign n19bar = in[3];
  assign n19 = inbar[3];
  assign n18bar = in[2];
  assign n18 = inbar[2];
  assign n17bar = in_0;
  assign n17 = in_0bar;
  OR2_X1 U5 ( .A1(n16), .A2(n15), .ZN(out[4]) );
  AND2_X1 U5bar ( .A1(n16bar), .A2(n15bar), .ZN(outbar[4]) );
  AND2_X1 U6 ( .A1(in[3]), .A2(n20), .ZN(n15) );
  OR2_X1 U6bar ( .A1(inbar[3]), .A2(n20bar), .ZN(n15bar) );
  AND2_X1 U7 ( .A1(in_7), .A2(n19), .ZN(n16) );
  OR2_X1 U7bar ( .A1(in_7bar), .A2(n19bar), .ZN(n16bar) );
  OR2_X1 U8 ( .A1(n14), .A2(n13), .ZN(out[3]) );
  AND2_X1 U8bar ( .A1(n14bar), .A2(n13bar), .ZN(outbar[3]) );
  AND2_X1 U9 ( .A1(in[2]), .A2(n20), .ZN(n13) );
  OR2_X1 U9bar ( .A1(inbar[2]), .A2(n20bar), .ZN(n13bar) );
  AND2_X1 U10 ( .A1(in_7), .A2(n18), .ZN(n14) );
  OR2_X1 U10bar ( .A1(in_7bar), .A2(n18bar), .ZN(n14bar) );
  OR2_X1 U11 ( .A1(n12), .A2(n11), .ZN(out[1]) );
  AND2_X1 U11bar ( .A1(n12bar), .A2(n11bar), .ZN(outbar[1]) );
  AND2_X1 U12 ( .A1(in_0), .A2(n20), .ZN(n11) );
  OR2_X1 U12bar ( .A1(in_0bar), .A2(n20bar), .ZN(n11bar) );
  AND2_X1 U13 ( .A1(in_7), .A2(n17), .ZN(n12) );
  OR2_X1 U13bar ( .A1(in_7bar), .A2(n17bar), .ZN(n12bar) );
endmodule

module scale2_11 ( in, inbar, out, outbar );

  input wire [7:0] in;
  input wire [7:0] inbar;
//input_done

  output wire [7:0] out;
  output wire [7:0] outbar;
//output_done

  wire in_0;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_1;
  wire in_7;
  wire n11;
  wire n12;
  wire n13;
  wire n14;
  wire n15;
  wire n16;
  wire n17;
  wire n18;
  wire n19;
  wire n20;
  wire in_0bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_1bar;
  wire in_7bar;
  wire n11bar;
  wire n12bar;
  wire n13bar;
  wire n14bar;
  wire n15bar;
  wire n16bar;
  wire n17bar;
  wire n18bar;
  wire n19bar;
  wire n20bar;
//wire_done

  assign in_0 = in[0];
  assign out[7] = in_6;
  assign in_6  = in[6];
  assign out[6] = in_5;
  assign in_5  = in[5];
  assign out[5] = in_4;
  assign in_4  = in[4];
  assign out[2] = in_1;
  assign in_1  = in[1];
  assign out[0] = in_7;
  assign in_7  = in[7];
  assign in_0bar = inbar[0];
  assign outbar[7] = in_6bar;
  assign in_6bar = inbar[6];
  assign outbar[6] = in_5bar;
  assign in_5bar = inbar[5];
  assign outbar[5] = in_4bar;
  assign in_4bar = inbar[4];
  assign outbar[2] = in_1bar;
  assign in_1bar = inbar[1];
  assign outbar[0] = in_7bar;
  assign in_7bar = inbar[7];
//assign_done

  assign n20bar = in_7;
  assign n20 = in_7bar;
  assign n19bar = in[3];
  assign n19 = inbar[3];
  assign n18bar = in[2];
  assign n18 = inbar[2];
  assign n17bar = in_0;
  assign n17 = in_0bar;
  OR2_X1 U5 ( .A1(n16), .A2(n15), .ZN(out[4]) );
  AND2_X1 U5bar ( .A1(n16bar), .A2(n15bar), .ZN(outbar[4]) );
  AND2_X1 U6 ( .A1(in[3]), .A2(n20), .ZN(n15) );
  OR2_X1 U6bar ( .A1(inbar[3]), .A2(n20bar), .ZN(n15bar) );
  AND2_X1 U7 ( .A1(in_7), .A2(n19), .ZN(n16) );
  OR2_X1 U7bar ( .A1(in_7bar), .A2(n19bar), .ZN(n16bar) );
  OR2_X1 U8 ( .A1(n14), .A2(n13), .ZN(out[3]) );
  AND2_X1 U8bar ( .A1(n14bar), .A2(n13bar), .ZN(outbar[3]) );
  AND2_X1 U9 ( .A1(in[2]), .A2(n20), .ZN(n13) );
  OR2_X1 U9bar ( .A1(inbar[2]), .A2(n20bar), .ZN(n13bar) );
  AND2_X1 U10 ( .A1(in_7), .A2(n18), .ZN(n14) );
  OR2_X1 U10bar ( .A1(in_7bar), .A2(n18bar), .ZN(n14bar) );
  OR2_X1 U11 ( .A1(n12), .A2(n11), .ZN(out[1]) );
  AND2_X1 U11bar ( .A1(n12bar), .A2(n11bar), .ZN(outbar[1]) );
  AND2_X1 U12 ( .A1(in_0), .A2(n20), .ZN(n11) );
  OR2_X1 U12bar ( .A1(in_0bar), .A2(n20bar), .ZN(n11bar) );
  AND2_X1 U13 ( .A1(in_7), .A2(n17), .ZN(n12) );
  OR2_X1 U13bar ( .A1(in_7bar), .A2(n17bar), .ZN(n12bar) );
endmodule

module scale2_12 ( in, inbar, out, outbar );

  input wire [7:0] in;
  input wire [7:0] inbar;
//input_done

  output wire [7:0] out;
  output wire [7:0] outbar;
//output_done

  wire in_0;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_1;
  wire in_7;
  wire n11;
  wire n12;
  wire n13;
  wire n14;
  wire n15;
  wire n16;
  wire n17;
  wire n18;
  wire n19;
  wire n20;
  wire in_0bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_1bar;
  wire in_7bar;
  wire n11bar;
  wire n12bar;
  wire n13bar;
  wire n14bar;
  wire n15bar;
  wire n16bar;
  wire n17bar;
  wire n18bar;
  wire n19bar;
  wire n20bar;
//wire_done

  assign in_0 = in[0];
  assign out[7] = in_6;
  assign in_6  = in[6];
  assign out[6] = in_5;
  assign in_5  = in[5];
  assign out[5] = in_4;
  assign in_4  = in[4];
  assign out[2] = in_1;
  assign in_1  = in[1];
  assign out[0] = in_7;
  assign in_7  = in[7];
  assign in_0bar = inbar[0];
  assign outbar[7] = in_6bar;
  assign in_6bar = inbar[6];
  assign outbar[6] = in_5bar;
  assign in_5bar = inbar[5];
  assign outbar[5] = in_4bar;
  assign in_4bar = inbar[4];
  assign outbar[2] = in_1bar;
  assign in_1bar = inbar[1];
  assign outbar[0] = in_7bar;
  assign in_7bar = inbar[7];
//assign_done

  assign n20bar = in_7;
  assign n20 = in_7bar;
  assign n19bar = in[3];
  assign n19 = inbar[3];
  assign n18bar = in[2];
  assign n18 = inbar[2];
  assign n17bar = in_0;
  assign n17 = in_0bar;
  OR2_X1 U5 ( .A1(n16), .A2(n15), .ZN(out[4]) );
  AND2_X1 U5bar ( .A1(n16bar), .A2(n15bar), .ZN(outbar[4]) );
  AND2_X1 U6 ( .A1(in[3]), .A2(n20), .ZN(n15) );
  OR2_X1 U6bar ( .A1(inbar[3]), .A2(n20bar), .ZN(n15bar) );
  AND2_X1 U7 ( .A1(in_7), .A2(n19), .ZN(n16) );
  OR2_X1 U7bar ( .A1(in_7bar), .A2(n19bar), .ZN(n16bar) );
  OR2_X1 U8 ( .A1(n14), .A2(n13), .ZN(out[3]) );
  AND2_X1 U8bar ( .A1(n14bar), .A2(n13bar), .ZN(outbar[3]) );
  AND2_X1 U9 ( .A1(in[2]), .A2(n20), .ZN(n13) );
  OR2_X1 U9bar ( .A1(inbar[2]), .A2(n20bar), .ZN(n13bar) );
  AND2_X1 U10 ( .A1(in_7), .A2(n18), .ZN(n14) );
  OR2_X1 U10bar ( .A1(in_7bar), .A2(n18bar), .ZN(n14bar) );
  OR2_X1 U11 ( .A1(n12), .A2(n11), .ZN(out[1]) );
  AND2_X1 U11bar ( .A1(n12bar), .A2(n11bar), .ZN(outbar[1]) );
  AND2_X1 U12 ( .A1(in_0), .A2(n20), .ZN(n11) );
  OR2_X1 U12bar ( .A1(in_0bar), .A2(n20bar), .ZN(n11bar) );
  AND2_X1 U13 ( .A1(in_7), .A2(n17), .ZN(n12) );
  OR2_X1 U13bar ( .A1(in_7bar), .A2(n17bar), .ZN(n12bar) );
endmodule

module byteXor_10 ( a, abar, b, bbar, y, ybar );

  input wire [7:0] a;
  input wire [7:0] b;
  input wire [7:0] abar;
  input wire [7:0] bbar;
//input_done

  output wire [7:0] y;
  output wire [7:0] ybar;
//output_done

  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n33bar;
  wire n34bar;
  wire n35bar;
  wire n36bar;
  wire n37bar;
  wire n38bar;
  wire n39bar;
  wire n40bar;
  wire n41bar;
  wire n42bar;
  wire n43bar;
  wire n44bar;
  wire n45bar;
  wire n46bar;
  wire n47bar;
  wire n48bar;
  wire n49bar;
  wire n50bar;
  wire n51bar;
  wire n52bar;
  wire n53bar;
  wire n54bar;
  wire n55bar;
  wire n56bar;
  wire n57bar;
  wire n58bar;
  wire n59bar;
  wire n60bar;
  wire n61bar;
  wire n62bar;
  wire n63bar;
  wire n64bar;
//wire_done

 //assign_done

  assign n64bar = n47;
  assign n64 = n47bar;
  assign n63bar = a[7];
  assign n63 = abar[7];
  assign n62bar = n45;
  assign n62 = n45bar;
  assign n61bar = a[6];
  assign n61 = abar[6];
  assign n60bar = n43;
  assign n60 = n43bar;
  assign n59bar = a[5];
  assign n59 = abar[5];
  assign n58bar = n41;
  assign n58 = n41bar;
  assign n57bar = a[4];
  assign n57 = abar[4];
  assign n56bar = n39;
  assign n56 = n39bar;
  assign n55bar = a[3];
  assign n55 = abar[3];
  assign n54bar = n37;
  assign n54 = n37bar;
  assign n53bar = a[2];
  assign n53 = abar[2];
  assign n52bar = n35;
  assign n52 = n35bar;
  assign n51bar = a[1];
  assign n51 = abar[1];
  assign n50bar = n33;
  assign n50 = n33bar;
  assign n49bar = a[0];
  assign n49 = abar[0];
  OR2_X1 U17 ( .A1(n48), .A2(n64), .ZN(y[7]) );
  AND2_X1 U17bar ( .A1(n48bar), .A2(n64bar), .ZN(ybar[7]) );
  OR2_X1 U18 ( .A1(n63), .A2(b[7]), .ZN(n47) );
  AND2_X1 U18bar ( .A1(n63bar), .A2(bbar[7]), .ZN(n47bar) );
  AND2_X1 U19 ( .A1(b[7]), .A2(n63), .ZN(n48) );
  OR2_X1 U19bar ( .A1(bbar[7]), .A2(n63bar), .ZN(n48bar) );
  OR2_X1 U20 ( .A1(n46), .A2(n62), .ZN(y[6]) );
  AND2_X1 U20bar ( .A1(n46bar), .A2(n62bar), .ZN(ybar[6]) );
  OR2_X1 U21 ( .A1(n61), .A2(b[6]), .ZN(n45) );
  AND2_X1 U21bar ( .A1(n61bar), .A2(bbar[6]), .ZN(n45bar) );
  AND2_X1 U22 ( .A1(b[6]), .A2(n61), .ZN(n46) );
  OR2_X1 U22bar ( .A1(bbar[6]), .A2(n61bar), .ZN(n46bar) );
  OR2_X1 U23 ( .A1(n44), .A2(n60), .ZN(y[5]) );
  AND2_X1 U23bar ( .A1(n44bar), .A2(n60bar), .ZN(ybar[5]) );
  OR2_X1 U24 ( .A1(n59), .A2(b[5]), .ZN(n43) );
  AND2_X1 U24bar ( .A1(n59bar), .A2(bbar[5]), .ZN(n43bar) );
  AND2_X1 U25 ( .A1(b[5]), .A2(n59), .ZN(n44) );
  OR2_X1 U25bar ( .A1(bbar[5]), .A2(n59bar), .ZN(n44bar) );
  OR2_X1 U26 ( .A1(n42), .A2(n58), .ZN(y[4]) );
  AND2_X1 U26bar ( .A1(n42bar), .A2(n58bar), .ZN(ybar[4]) );
  OR2_X1 U27 ( .A1(n57), .A2(b[4]), .ZN(n41) );
  AND2_X1 U27bar ( .A1(n57bar), .A2(bbar[4]), .ZN(n41bar) );
  AND2_X1 U28 ( .A1(b[4]), .A2(n57), .ZN(n42) );
  OR2_X1 U28bar ( .A1(bbar[4]), .A2(n57bar), .ZN(n42bar) );
  OR2_X1 U29 ( .A1(n40), .A2(n56), .ZN(y[3]) );
  AND2_X1 U29bar ( .A1(n40bar), .A2(n56bar), .ZN(ybar[3]) );
  OR2_X1 U30 ( .A1(n55), .A2(b[3]), .ZN(n39) );
  AND2_X1 U30bar ( .A1(n55bar), .A2(bbar[3]), .ZN(n39bar) );
  AND2_X1 U31 ( .A1(b[3]), .A2(n55), .ZN(n40) );
  OR2_X1 U31bar ( .A1(bbar[3]), .A2(n55bar), .ZN(n40bar) );
  OR2_X1 U32 ( .A1(n38), .A2(n54), .ZN(y[2]) );
  AND2_X1 U32bar ( .A1(n38bar), .A2(n54bar), .ZN(ybar[2]) );
  OR2_X1 U33 ( .A1(n53), .A2(b[2]), .ZN(n37) );
  AND2_X1 U33bar ( .A1(n53bar), .A2(bbar[2]), .ZN(n37bar) );
  AND2_X1 U34 ( .A1(b[2]), .A2(n53), .ZN(n38) );
  OR2_X1 U34bar ( .A1(bbar[2]), .A2(n53bar), .ZN(n38bar) );
  OR2_X1 U35 ( .A1(n36), .A2(n52), .ZN(y[1]) );
  AND2_X1 U35bar ( .A1(n36bar), .A2(n52bar), .ZN(ybar[1]) );
  OR2_X1 U36 ( .A1(n51), .A2(b[1]), .ZN(n35) );
  AND2_X1 U36bar ( .A1(n51bar), .A2(bbar[1]), .ZN(n35bar) );
  AND2_X1 U37 ( .A1(b[1]), .A2(n51), .ZN(n36) );
  OR2_X1 U37bar ( .A1(bbar[1]), .A2(n51bar), .ZN(n36bar) );
  OR2_X1 U38 ( .A1(n34), .A2(n50), .ZN(y[0]) );
  AND2_X1 U38bar ( .A1(n34bar), .A2(n50bar), .ZN(ybar[0]) );
  OR2_X1 U39 ( .A1(n49), .A2(b[0]), .ZN(n33) );
  AND2_X1 U39bar ( .A1(n49bar), .A2(bbar[0]), .ZN(n33bar) );
  AND2_X1 U40 ( .A1(b[0]), .A2(n49), .ZN(n34) );
  OR2_X1 U40bar ( .A1(bbar[0]), .A2(n49bar), .ZN(n34bar) );
endmodule

module byteXor_11 ( a, abar, b, bbar, y, ybar );

  input wire [7:0] a;
  input wire [7:0] b;
  input wire [7:0] abar;
  input wire [7:0] bbar;
//input_done

  output wire [7:0] y;
  output wire [7:0] ybar;
//output_done

  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n33bar;
  wire n34bar;
  wire n35bar;
  wire n36bar;
  wire n37bar;
  wire n38bar;
  wire n39bar;
  wire n40bar;
  wire n41bar;
  wire n42bar;
  wire n43bar;
  wire n44bar;
  wire n45bar;
  wire n46bar;
  wire n47bar;
  wire n48bar;
  wire n49bar;
  wire n50bar;
  wire n51bar;
  wire n52bar;
  wire n53bar;
  wire n54bar;
  wire n55bar;
  wire n56bar;
  wire n57bar;
  wire n58bar;
  wire n59bar;
  wire n60bar;
  wire n61bar;
  wire n62bar;
  wire n63bar;
  wire n64bar;
//wire_done

 //assign_done

  assign n64bar = n47;
  assign n64 = n47bar;
  assign n63bar = a[7];
  assign n63 = abar[7];
  assign n62bar = n45;
  assign n62 = n45bar;
  assign n61bar = a[6];
  assign n61 = abar[6];
  assign n60bar = n43;
  assign n60 = n43bar;
  assign n59bar = a[5];
  assign n59 = abar[5];
  assign n58bar = n41;
  assign n58 = n41bar;
  assign n57bar = a[4];
  assign n57 = abar[4];
  assign n56bar = n39;
  assign n56 = n39bar;
  assign n55bar = a[3];
  assign n55 = abar[3];
  assign n54bar = n37;
  assign n54 = n37bar;
  assign n53bar = a[2];
  assign n53 = abar[2];
  assign n52bar = n35;
  assign n52 = n35bar;
  assign n51bar = a[1];
  assign n51 = abar[1];
  assign n50bar = n33;
  assign n50 = n33bar;
  assign n49bar = a[0];
  assign n49 = abar[0];
  OR2_X1 U17 ( .A1(n48), .A2(n64), .ZN(y[7]) );
  AND2_X1 U17bar ( .A1(n48bar), .A2(n64bar), .ZN(ybar[7]) );
  OR2_X1 U18 ( .A1(n63), .A2(b[7]), .ZN(n47) );
  AND2_X1 U18bar ( .A1(n63bar), .A2(bbar[7]), .ZN(n47bar) );
  AND2_X1 U19 ( .A1(b[7]), .A2(n63), .ZN(n48) );
  OR2_X1 U19bar ( .A1(bbar[7]), .A2(n63bar), .ZN(n48bar) );
  OR2_X1 U20 ( .A1(n46), .A2(n62), .ZN(y[6]) );
  AND2_X1 U20bar ( .A1(n46bar), .A2(n62bar), .ZN(ybar[6]) );
  OR2_X1 U21 ( .A1(n61), .A2(b[6]), .ZN(n45) );
  AND2_X1 U21bar ( .A1(n61bar), .A2(bbar[6]), .ZN(n45bar) );
  AND2_X1 U22 ( .A1(b[6]), .A2(n61), .ZN(n46) );
  OR2_X1 U22bar ( .A1(bbar[6]), .A2(n61bar), .ZN(n46bar) );
  OR2_X1 U23 ( .A1(n44), .A2(n60), .ZN(y[5]) );
  AND2_X1 U23bar ( .A1(n44bar), .A2(n60bar), .ZN(ybar[5]) );
  OR2_X1 U24 ( .A1(n59), .A2(b[5]), .ZN(n43) );
  AND2_X1 U24bar ( .A1(n59bar), .A2(bbar[5]), .ZN(n43bar) );
  AND2_X1 U25 ( .A1(b[5]), .A2(n59), .ZN(n44) );
  OR2_X1 U25bar ( .A1(bbar[5]), .A2(n59bar), .ZN(n44bar) );
  OR2_X1 U26 ( .A1(n42), .A2(n58), .ZN(y[4]) );
  AND2_X1 U26bar ( .A1(n42bar), .A2(n58bar), .ZN(ybar[4]) );
  OR2_X1 U27 ( .A1(n57), .A2(b[4]), .ZN(n41) );
  AND2_X1 U27bar ( .A1(n57bar), .A2(bbar[4]), .ZN(n41bar) );
  AND2_X1 U28 ( .A1(b[4]), .A2(n57), .ZN(n42) );
  OR2_X1 U28bar ( .A1(bbar[4]), .A2(n57bar), .ZN(n42bar) );
  OR2_X1 U29 ( .A1(n40), .A2(n56), .ZN(y[3]) );
  AND2_X1 U29bar ( .A1(n40bar), .A2(n56bar), .ZN(ybar[3]) );
  OR2_X1 U30 ( .A1(n55), .A2(b[3]), .ZN(n39) );
  AND2_X1 U30bar ( .A1(n55bar), .A2(bbar[3]), .ZN(n39bar) );
  AND2_X1 U31 ( .A1(b[3]), .A2(n55), .ZN(n40) );
  OR2_X1 U31bar ( .A1(bbar[3]), .A2(n55bar), .ZN(n40bar) );
  OR2_X1 U32 ( .A1(n38), .A2(n54), .ZN(y[2]) );
  AND2_X1 U32bar ( .A1(n38bar), .A2(n54bar), .ZN(ybar[2]) );
  OR2_X1 U33 ( .A1(n53), .A2(b[2]), .ZN(n37) );
  AND2_X1 U33bar ( .A1(n53bar), .A2(bbar[2]), .ZN(n37bar) );
  AND2_X1 U34 ( .A1(b[2]), .A2(n53), .ZN(n38) );
  OR2_X1 U34bar ( .A1(bbar[2]), .A2(n53bar), .ZN(n38bar) );
  OR2_X1 U35 ( .A1(n36), .A2(n52), .ZN(y[1]) );
  AND2_X1 U35bar ( .A1(n36bar), .A2(n52bar), .ZN(ybar[1]) );
  OR2_X1 U36 ( .A1(n51), .A2(b[1]), .ZN(n35) );
  AND2_X1 U36bar ( .A1(n51bar), .A2(bbar[1]), .ZN(n35bar) );
  AND2_X1 U37 ( .A1(b[1]), .A2(n51), .ZN(n36) );
  OR2_X1 U37bar ( .A1(bbar[1]), .A2(n51bar), .ZN(n36bar) );
  OR2_X1 U38 ( .A1(n34), .A2(n50), .ZN(y[0]) );
  AND2_X1 U38bar ( .A1(n34bar), .A2(n50bar), .ZN(ybar[0]) );
  OR2_X1 U39 ( .A1(n49), .A2(b[0]), .ZN(n33) );
  AND2_X1 U39bar ( .A1(n49bar), .A2(bbar[0]), .ZN(n33bar) );
  AND2_X1 U40 ( .A1(b[0]), .A2(n49), .ZN(n34) );
  OR2_X1 U40bar ( .A1(bbar[0]), .A2(n49bar), .ZN(n34bar) );
endmodule

module byteXor_12 ( a, abar, b, bbar, y, ybar );

  input wire [7:0] a;
  input wire [7:0] b;
  input wire [7:0] abar;
  input wire [7:0] bbar;
//input_done

  output wire [7:0] y;
  output wire [7:0] ybar;
//output_done

  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n33bar;
  wire n34bar;
  wire n35bar;
  wire n36bar;
  wire n37bar;
  wire n38bar;
  wire n39bar;
  wire n40bar;
  wire n41bar;
  wire n42bar;
  wire n43bar;
  wire n44bar;
  wire n45bar;
  wire n46bar;
  wire n47bar;
  wire n48bar;
  wire n49bar;
  wire n50bar;
  wire n51bar;
  wire n52bar;
  wire n53bar;
  wire n54bar;
  wire n55bar;
  wire n56bar;
  wire n57bar;
  wire n58bar;
  wire n59bar;
  wire n60bar;
  wire n61bar;
  wire n62bar;
  wire n63bar;
  wire n64bar;
//wire_done

 //assign_done

  assign n64bar = n47;
  assign n64 = n47bar;
  assign n63bar = a[7];
  assign n63 = abar[7];
  assign n62bar = n45;
  assign n62 = n45bar;
  assign n61bar = a[6];
  assign n61 = abar[6];
  assign n60bar = n43;
  assign n60 = n43bar;
  assign n59bar = a[5];
  assign n59 = abar[5];
  assign n58bar = n41;
  assign n58 = n41bar;
  assign n57bar = a[4];
  assign n57 = abar[4];
  assign n56bar = n39;
  assign n56 = n39bar;
  assign n55bar = a[3];
  assign n55 = abar[3];
  assign n54bar = n37;
  assign n54 = n37bar;
  assign n53bar = a[2];
  assign n53 = abar[2];
  assign n52bar = n35;
  assign n52 = n35bar;
  assign n51bar = a[1];
  assign n51 = abar[1];
  assign n50bar = n33;
  assign n50 = n33bar;
  assign n49bar = a[0];
  assign n49 = abar[0];
  OR2_X1 U17 ( .A1(n48), .A2(n64), .ZN(y[7]) );
  AND2_X1 U17bar ( .A1(n48bar), .A2(n64bar), .ZN(ybar[7]) );
  OR2_X1 U18 ( .A1(n63), .A2(b[7]), .ZN(n47) );
  AND2_X1 U18bar ( .A1(n63bar), .A2(bbar[7]), .ZN(n47bar) );
  AND2_X1 U19 ( .A1(b[7]), .A2(n63), .ZN(n48) );
  OR2_X1 U19bar ( .A1(bbar[7]), .A2(n63bar), .ZN(n48bar) );
  OR2_X1 U20 ( .A1(n46), .A2(n62), .ZN(y[6]) );
  AND2_X1 U20bar ( .A1(n46bar), .A2(n62bar), .ZN(ybar[6]) );
  OR2_X1 U21 ( .A1(n61), .A2(b[6]), .ZN(n45) );
  AND2_X1 U21bar ( .A1(n61bar), .A2(bbar[6]), .ZN(n45bar) );
  AND2_X1 U22 ( .A1(b[6]), .A2(n61), .ZN(n46) );
  OR2_X1 U22bar ( .A1(bbar[6]), .A2(n61bar), .ZN(n46bar) );
  OR2_X1 U23 ( .A1(n44), .A2(n60), .ZN(y[5]) );
  AND2_X1 U23bar ( .A1(n44bar), .A2(n60bar), .ZN(ybar[5]) );
  OR2_X1 U24 ( .A1(n59), .A2(b[5]), .ZN(n43) );
  AND2_X1 U24bar ( .A1(n59bar), .A2(bbar[5]), .ZN(n43bar) );
  AND2_X1 U25 ( .A1(b[5]), .A2(n59), .ZN(n44) );
  OR2_X1 U25bar ( .A1(bbar[5]), .A2(n59bar), .ZN(n44bar) );
  OR2_X1 U26 ( .A1(n42), .A2(n58), .ZN(y[4]) );
  AND2_X1 U26bar ( .A1(n42bar), .A2(n58bar), .ZN(ybar[4]) );
  OR2_X1 U27 ( .A1(n57), .A2(b[4]), .ZN(n41) );
  AND2_X1 U27bar ( .A1(n57bar), .A2(bbar[4]), .ZN(n41bar) );
  AND2_X1 U28 ( .A1(b[4]), .A2(n57), .ZN(n42) );
  OR2_X1 U28bar ( .A1(bbar[4]), .A2(n57bar), .ZN(n42bar) );
  OR2_X1 U29 ( .A1(n40), .A2(n56), .ZN(y[3]) );
  AND2_X1 U29bar ( .A1(n40bar), .A2(n56bar), .ZN(ybar[3]) );
  OR2_X1 U30 ( .A1(n55), .A2(b[3]), .ZN(n39) );
  AND2_X1 U30bar ( .A1(n55bar), .A2(bbar[3]), .ZN(n39bar) );
  AND2_X1 U31 ( .A1(b[3]), .A2(n55), .ZN(n40) );
  OR2_X1 U31bar ( .A1(bbar[3]), .A2(n55bar), .ZN(n40bar) );
  OR2_X1 U32 ( .A1(n38), .A2(n54), .ZN(y[2]) );
  AND2_X1 U32bar ( .A1(n38bar), .A2(n54bar), .ZN(ybar[2]) );
  OR2_X1 U33 ( .A1(n53), .A2(b[2]), .ZN(n37) );
  AND2_X1 U33bar ( .A1(n53bar), .A2(bbar[2]), .ZN(n37bar) );
  AND2_X1 U34 ( .A1(b[2]), .A2(n53), .ZN(n38) );
  OR2_X1 U34bar ( .A1(bbar[2]), .A2(n53bar), .ZN(n38bar) );
  OR2_X1 U35 ( .A1(n36), .A2(n52), .ZN(y[1]) );
  AND2_X1 U35bar ( .A1(n36bar), .A2(n52bar), .ZN(ybar[1]) );
  OR2_X1 U36 ( .A1(n51), .A2(b[1]), .ZN(n35) );
  AND2_X1 U36bar ( .A1(n51bar), .A2(bbar[1]), .ZN(n35bar) );
  AND2_X1 U37 ( .A1(b[1]), .A2(n51), .ZN(n36) );
  OR2_X1 U37bar ( .A1(bbar[1]), .A2(n51bar), .ZN(n36bar) );
  OR2_X1 U38 ( .A1(n34), .A2(n50), .ZN(y[0]) );
  AND2_X1 U38bar ( .A1(n34bar), .A2(n50bar), .ZN(ybar[0]) );
  OR2_X1 U39 ( .A1(n49), .A2(b[0]), .ZN(n33) );
  AND2_X1 U39bar ( .A1(n49bar), .A2(bbar[0]), .ZN(n33bar) );
  AND2_X1 U40 ( .A1(b[0]), .A2(n49), .ZN(n34) );
  OR2_X1 U40bar ( .A1(bbar[0]), .A2(n49bar), .ZN(n34bar) );
endmodule

module byteXor_13 ( a, abar, b, bbar, y, ybar );

  input wire [7:0] a;
  input wire [7:0] b;
  input wire [7:0] abar;
  input wire [7:0] bbar;
//input_done

  output wire [7:0] y;
  output wire [7:0] ybar;
//output_done

  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n33bar;
  wire n34bar;
  wire n35bar;
  wire n36bar;
  wire n37bar;
  wire n38bar;
  wire n39bar;
  wire n40bar;
  wire n41bar;
  wire n42bar;
  wire n43bar;
  wire n44bar;
  wire n45bar;
  wire n46bar;
  wire n47bar;
  wire n48bar;
  wire n49bar;
  wire n50bar;
  wire n51bar;
  wire n52bar;
  wire n53bar;
  wire n54bar;
  wire n55bar;
  wire n56bar;
  wire n57bar;
  wire n58bar;
  wire n59bar;
  wire n60bar;
  wire n61bar;
  wire n62bar;
  wire n63bar;
  wire n64bar;
//wire_done

 //assign_done

  assign n64bar = n47;
  assign n64 = n47bar;
  assign n63bar = a[7];
  assign n63 = abar[7];
  assign n62bar = n45;
  assign n62 = n45bar;
  assign n61bar = a[6];
  assign n61 = abar[6];
  assign n60bar = n43;
  assign n60 = n43bar;
  assign n59bar = a[5];
  assign n59 = abar[5];
  assign n58bar = n41;
  assign n58 = n41bar;
  assign n57bar = a[4];
  assign n57 = abar[4];
  assign n56bar = n39;
  assign n56 = n39bar;
  assign n55bar = a[3];
  assign n55 = abar[3];
  assign n54bar = n37;
  assign n54 = n37bar;
  assign n53bar = a[2];
  assign n53 = abar[2];
  assign n52bar = n35;
  assign n52 = n35bar;
  assign n51bar = a[1];
  assign n51 = abar[1];
  assign n50bar = n33;
  assign n50 = n33bar;
  assign n49bar = a[0];
  assign n49 = abar[0];
  OR2_X1 U17 ( .A1(n48), .A2(n64), .ZN(y[7]) );
  AND2_X1 U17bar ( .A1(n48bar), .A2(n64bar), .ZN(ybar[7]) );
  OR2_X1 U18 ( .A1(n63), .A2(b[7]), .ZN(n47) );
  AND2_X1 U18bar ( .A1(n63bar), .A2(bbar[7]), .ZN(n47bar) );
  AND2_X1 U19 ( .A1(b[7]), .A2(n63), .ZN(n48) );
  OR2_X1 U19bar ( .A1(bbar[7]), .A2(n63bar), .ZN(n48bar) );
  OR2_X1 U20 ( .A1(n46), .A2(n62), .ZN(y[6]) );
  AND2_X1 U20bar ( .A1(n46bar), .A2(n62bar), .ZN(ybar[6]) );
  OR2_X1 U21 ( .A1(n61), .A2(b[6]), .ZN(n45) );
  AND2_X1 U21bar ( .A1(n61bar), .A2(bbar[6]), .ZN(n45bar) );
  AND2_X1 U22 ( .A1(b[6]), .A2(n61), .ZN(n46) );
  OR2_X1 U22bar ( .A1(bbar[6]), .A2(n61bar), .ZN(n46bar) );
  OR2_X1 U23 ( .A1(n44), .A2(n60), .ZN(y[5]) );
  AND2_X1 U23bar ( .A1(n44bar), .A2(n60bar), .ZN(ybar[5]) );
  OR2_X1 U24 ( .A1(n59), .A2(b[5]), .ZN(n43) );
  AND2_X1 U24bar ( .A1(n59bar), .A2(bbar[5]), .ZN(n43bar) );
  AND2_X1 U25 ( .A1(b[5]), .A2(n59), .ZN(n44) );
  OR2_X1 U25bar ( .A1(bbar[5]), .A2(n59bar), .ZN(n44bar) );
  OR2_X1 U26 ( .A1(n42), .A2(n58), .ZN(y[4]) );
  AND2_X1 U26bar ( .A1(n42bar), .A2(n58bar), .ZN(ybar[4]) );
  OR2_X1 U27 ( .A1(n57), .A2(b[4]), .ZN(n41) );
  AND2_X1 U27bar ( .A1(n57bar), .A2(bbar[4]), .ZN(n41bar) );
  AND2_X1 U28 ( .A1(b[4]), .A2(n57), .ZN(n42) );
  OR2_X1 U28bar ( .A1(bbar[4]), .A2(n57bar), .ZN(n42bar) );
  OR2_X1 U29 ( .A1(n40), .A2(n56), .ZN(y[3]) );
  AND2_X1 U29bar ( .A1(n40bar), .A2(n56bar), .ZN(ybar[3]) );
  OR2_X1 U30 ( .A1(n55), .A2(b[3]), .ZN(n39) );
  AND2_X1 U30bar ( .A1(n55bar), .A2(bbar[3]), .ZN(n39bar) );
  AND2_X1 U31 ( .A1(b[3]), .A2(n55), .ZN(n40) );
  OR2_X1 U31bar ( .A1(bbar[3]), .A2(n55bar), .ZN(n40bar) );
  OR2_X1 U32 ( .A1(n38), .A2(n54), .ZN(y[2]) );
  AND2_X1 U32bar ( .A1(n38bar), .A2(n54bar), .ZN(ybar[2]) );
  OR2_X1 U33 ( .A1(n53), .A2(b[2]), .ZN(n37) );
  AND2_X1 U33bar ( .A1(n53bar), .A2(bbar[2]), .ZN(n37bar) );
  AND2_X1 U34 ( .A1(b[2]), .A2(n53), .ZN(n38) );
  OR2_X1 U34bar ( .A1(bbar[2]), .A2(n53bar), .ZN(n38bar) );
  OR2_X1 U35 ( .A1(n36), .A2(n52), .ZN(y[1]) );
  AND2_X1 U35bar ( .A1(n36bar), .A2(n52bar), .ZN(ybar[1]) );
  OR2_X1 U36 ( .A1(n51), .A2(b[1]), .ZN(n35) );
  AND2_X1 U36bar ( .A1(n51bar), .A2(bbar[1]), .ZN(n35bar) );
  AND2_X1 U37 ( .A1(b[1]), .A2(n51), .ZN(n36) );
  OR2_X1 U37bar ( .A1(bbar[1]), .A2(n51bar), .ZN(n36bar) );
  OR2_X1 U38 ( .A1(n34), .A2(n50), .ZN(y[0]) );
  AND2_X1 U38bar ( .A1(n34bar), .A2(n50bar), .ZN(ybar[0]) );
  OR2_X1 U39 ( .A1(n49), .A2(b[0]), .ZN(n33) );
  AND2_X1 U39bar ( .A1(n49bar), .A2(bbar[0]), .ZN(n33bar) );
  AND2_X1 U40 ( .A1(b[0]), .A2(n49), .ZN(n34) );
  OR2_X1 U40bar ( .A1(bbar[0]), .A2(n49bar), .ZN(n34bar) );
endmodule

module byteXor4_9 ( a, abar, b, bbar, c, cbar, d, dbar, y, ybar );

  input wire [7:0] a;
  input wire [7:0] b;
  input wire [7:0] c;
  input wire [7:0] d;
  input wire [7:0] abar;
  input wire [7:0] bbar;
  input wire [7:0] cbar;
  input wire [7:0] dbar;
//input_done

  output wire [7:0] y;
  output wire [7:0] ybar;
//output_done

  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n113bar;
  wire n114bar;
  wire n115bar;
  wire n116bar;
  wire n117bar;
  wire n118bar;
  wire n119bar;
  wire n120bar;
  wire n121bar;
  wire n122bar;
  wire n123bar;
  wire n124bar;
  wire n125bar;
  wire n126bar;
  wire n127bar;
  wire n128bar;
  wire n129bar;
  wire n130bar;
  wire n131bar;
  wire n132bar;
  wire n133bar;
  wire n134bar;
  wire n135bar;
  wire n136bar;
  wire n137bar;
  wire n138bar;
  wire n139bar;
  wire n140bar;
  wire n141bar;
  wire n142bar;
  wire n143bar;
  wire n144bar;
  wire n145bar;
  wire n146bar;
  wire n147bar;
  wire n148bar;
  wire n149bar;
  wire n150bar;
  wire n151bar;
  wire n152bar;
  wire n153bar;
  wire n154bar;
  wire n155bar;
  wire n156bar;
  wire n157bar;
  wire n158bar;
  wire n159bar;
  wire n160bar;
  wire n161bar;
  wire n162bar;
  wire n163bar;
  wire n164bar;
  wire n165bar;
  wire n166bar;
  wire n167bar;
  wire n168bar;
  wire n169bar;
  wire n170bar;
  wire n171bar;
  wire n172bar;
  wire n173bar;
  wire n174bar;
  wire n175bar;
  wire n176bar;
  wire n177bar;
  wire n178bar;
  wire n179bar;
  wire n180bar;
  wire n181bar;
  wire n182bar;
  wire n183bar;
  wire n184bar;
  wire n185bar;
  wire n186bar;
  wire n187bar;
  wire n188bar;
  wire n189bar;
  wire n190bar;
  wire n191bar;
  wire n192bar;
  wire n193bar;
  wire n194bar;
  wire n195bar;
  wire n196bar;
  wire n197bar;
  wire n198bar;
  wire n199bar;
  wire n200bar;
  wire n201bar;
  wire n202bar;
  wire n203bar;
  wire n204bar;
  wire n205bar;
  wire n206bar;
  wire n207bar;
  wire n208bar;
  wire n209bar;
  wire n210bar;
  wire n211bar;
  wire n212bar;
  wire n213bar;
  wire n214bar;
  wire n215bar;
  wire n216bar;
  wire n217bar;
  wire n218bar;
  wire n219bar;
  wire n220bar;
  wire n221bar;
  wire n222bar;
  wire n223bar;
  wire n224bar;
//wire_done

 //assign_done

  assign n224bar = n175;
  assign n224 = n175bar;
  assign n223bar = a[7];
  assign n223 = abar[7];
  assign n222bar = n167;
  assign n222 = n167bar;
  assign n221bar = a[6];
  assign n221 = abar[6];
  assign n220bar = n159;
  assign n220 = n159bar;
  assign n219bar = a[5];
  assign n219 = abar[5];
  assign n218bar = n151;
  assign n218 = n151bar;
  assign n217bar = a[4];
  assign n217 = abar[4];
  assign n216bar = n143;
  assign n216 = n143bar;
  assign n215bar = a[3];
  assign n215 = abar[3];
  assign n214bar = n135;
  assign n214 = n135bar;
  assign n213bar = a[2];
  assign n213 = abar[2];
  assign n212bar = n127;
  assign n212 = n127bar;
  assign n211bar = a[1];
  assign n211 = abar[1];
  assign n210bar = n119;
  assign n210 = n119bar;
  assign n209bar = a[0];
  assign n209 = abar[0];
  assign n208bar = b[7];
  assign n208 = bbar[7];
  assign n207bar = b[6];
  assign n207 = bbar[6];
  assign n206bar = b[5];
  assign n206 = bbar[5];
  assign n205bar = b[4];
  assign n205 = bbar[4];
  assign n204bar = b[3];
  assign n204 = bbar[3];
  assign n203bar = b[2];
  assign n203 = bbar[2];
  assign n202bar = b[1];
  assign n202 = bbar[1];
  assign n201bar = b[0];
  assign n201 = bbar[0];
  assign n200bar = n171;
  assign n200 = n171bar;
  assign n199bar = c[7];
  assign n199 = cbar[7];
  assign n198bar = n163;
  assign n198 = n163bar;
  assign n197bar = c[6];
  assign n197 = cbar[6];
  assign n196bar = n155;
  assign n196 = n155bar;
  assign n195bar = c[5];
  assign n195 = cbar[5];
  assign n194bar = n147;
  assign n194 = n147bar;
  assign n193bar = c[4];
  assign n193 = cbar[4];
  assign n192bar = n139;
  assign n192 = n139bar;
  assign n191bar = c[3];
  assign n191 = cbar[3];
  assign n190bar = n131;
  assign n190 = n131bar;
  assign n189bar = c[2];
  assign n189 = cbar[2];
  assign n188bar = n123;
  assign n188 = n123bar;
  assign n187bar = c[1];
  assign n187 = cbar[1];
  assign n186bar = n115;
  assign n186 = n115bar;
  assign n185bar = c[0];
  assign n185 = cbar[0];
  assign n184bar = d[7];
  assign n184 = dbar[7];
  assign n183bar = d[6];
  assign n183 = dbar[6];
  assign n182bar = d[5];
  assign n182 = dbar[5];
  assign n181bar = d[4];
  assign n181 = dbar[4];
  assign n180bar = d[3];
  assign n180 = dbar[3];
  assign n179bar = d[2];
  assign n179 = dbar[2];
  assign n178bar = d[1];
  assign n178 = dbar[1];
  assign n177bar = d[0];
  assign n177 = dbar[0];
  OR2_X1 U49 ( .A1(n176), .A2(n224), .ZN(y[7]) );
  AND2_X1 U49bar ( .A1(n176bar), .A2(n224bar), .ZN(ybar[7]) );
  OR2_X1 U50 ( .A1(n174), .A2(n200), .ZN(n175) );
  AND2_X1 U50bar ( .A1(n174bar), .A2(n200bar), .ZN(n175bar) );
  AND2_X1 U51 ( .A1(n200), .A2(n174), .ZN(n176) );
  OR2_X1 U51bar ( .A1(n200bar), .A2(n174bar), .ZN(n176bar) );
  AND2_X1 U52 ( .A1(n173), .A2(n172), .ZN(n174) );
  OR2_X1 U52bar ( .A1(n173bar), .A2(n172bar), .ZN(n174bar) );
  OR2_X1 U53 ( .A1(n223), .A2(b[7]), .ZN(n172) );
  AND2_X1 U53bar ( .A1(n223bar), .A2(bbar[7]), .ZN(n172bar) );
  OR2_X1 U54 ( .A1(n208), .A2(a[7]), .ZN(n173) );
  AND2_X1 U54bar ( .A1(n208bar), .A2(abar[7]), .ZN(n173bar) );
  AND2_X1 U55 ( .A1(n170), .A2(n169), .ZN(n171) );
  OR2_X1 U55bar ( .A1(n170bar), .A2(n169bar), .ZN(n171bar) );
  OR2_X1 U56 ( .A1(n199), .A2(d[7]), .ZN(n169) );
  AND2_X1 U56bar ( .A1(n199bar), .A2(dbar[7]), .ZN(n169bar) );
  OR2_X1 U57 ( .A1(n184), .A2(c[7]), .ZN(n170) );
  AND2_X1 U57bar ( .A1(n184bar), .A2(cbar[7]), .ZN(n170bar) );
  OR2_X1 U58 ( .A1(n168), .A2(n222), .ZN(y[6]) );
  AND2_X1 U58bar ( .A1(n168bar), .A2(n222bar), .ZN(ybar[6]) );
  OR2_X1 U59 ( .A1(n166), .A2(n198), .ZN(n167) );
  AND2_X1 U59bar ( .A1(n166bar), .A2(n198bar), .ZN(n167bar) );
  AND2_X1 U60 ( .A1(n198), .A2(n166), .ZN(n168) );
  OR2_X1 U60bar ( .A1(n198bar), .A2(n166bar), .ZN(n168bar) );
  AND2_X1 U61 ( .A1(n165), .A2(n164), .ZN(n166) );
  OR2_X1 U61bar ( .A1(n165bar), .A2(n164bar), .ZN(n166bar) );
  OR2_X1 U62 ( .A1(n221), .A2(b[6]), .ZN(n164) );
  AND2_X1 U62bar ( .A1(n221bar), .A2(bbar[6]), .ZN(n164bar) );
  OR2_X1 U63 ( .A1(n207), .A2(a[6]), .ZN(n165) );
  AND2_X1 U63bar ( .A1(n207bar), .A2(abar[6]), .ZN(n165bar) );
  AND2_X1 U64 ( .A1(n162), .A2(n161), .ZN(n163) );
  OR2_X1 U64bar ( .A1(n162bar), .A2(n161bar), .ZN(n163bar) );
  OR2_X1 U65 ( .A1(n197), .A2(d[6]), .ZN(n161) );
  AND2_X1 U65bar ( .A1(n197bar), .A2(dbar[6]), .ZN(n161bar) );
  OR2_X1 U66 ( .A1(n183), .A2(c[6]), .ZN(n162) );
  AND2_X1 U66bar ( .A1(n183bar), .A2(cbar[6]), .ZN(n162bar) );
  OR2_X1 U67 ( .A1(n160), .A2(n220), .ZN(y[5]) );
  AND2_X1 U67bar ( .A1(n160bar), .A2(n220bar), .ZN(ybar[5]) );
  OR2_X1 U68 ( .A1(n158), .A2(n196), .ZN(n159) );
  AND2_X1 U68bar ( .A1(n158bar), .A2(n196bar), .ZN(n159bar) );
  AND2_X1 U69 ( .A1(n196), .A2(n158), .ZN(n160) );
  OR2_X1 U69bar ( .A1(n196bar), .A2(n158bar), .ZN(n160bar) );
  AND2_X1 U70 ( .A1(n157), .A2(n156), .ZN(n158) );
  OR2_X1 U70bar ( .A1(n157bar), .A2(n156bar), .ZN(n158bar) );
  OR2_X1 U71 ( .A1(n219), .A2(b[5]), .ZN(n156) );
  AND2_X1 U71bar ( .A1(n219bar), .A2(bbar[5]), .ZN(n156bar) );
  OR2_X1 U72 ( .A1(n206), .A2(a[5]), .ZN(n157) );
  AND2_X1 U72bar ( .A1(n206bar), .A2(abar[5]), .ZN(n157bar) );
  AND2_X1 U73 ( .A1(n154), .A2(n153), .ZN(n155) );
  OR2_X1 U73bar ( .A1(n154bar), .A2(n153bar), .ZN(n155bar) );
  OR2_X1 U74 ( .A1(n195), .A2(d[5]), .ZN(n153) );
  AND2_X1 U74bar ( .A1(n195bar), .A2(dbar[5]), .ZN(n153bar) );
  OR2_X1 U75 ( .A1(n182), .A2(c[5]), .ZN(n154) );
  AND2_X1 U75bar ( .A1(n182bar), .A2(cbar[5]), .ZN(n154bar) );
  OR2_X1 U76 ( .A1(n152), .A2(n218), .ZN(y[4]) );
  AND2_X1 U76bar ( .A1(n152bar), .A2(n218bar), .ZN(ybar[4]) );
  OR2_X1 U77 ( .A1(n150), .A2(n194), .ZN(n151) );
  AND2_X1 U77bar ( .A1(n150bar), .A2(n194bar), .ZN(n151bar) );
  AND2_X1 U78 ( .A1(n194), .A2(n150), .ZN(n152) );
  OR2_X1 U78bar ( .A1(n194bar), .A2(n150bar), .ZN(n152bar) );
  AND2_X1 U79 ( .A1(n149), .A2(n148), .ZN(n150) );
  OR2_X1 U79bar ( .A1(n149bar), .A2(n148bar), .ZN(n150bar) );
  OR2_X1 U80 ( .A1(n217), .A2(b[4]), .ZN(n148) );
  AND2_X1 U80bar ( .A1(n217bar), .A2(bbar[4]), .ZN(n148bar) );
  OR2_X1 U81 ( .A1(n205), .A2(a[4]), .ZN(n149) );
  AND2_X1 U81bar ( .A1(n205bar), .A2(abar[4]), .ZN(n149bar) );
  AND2_X1 U82 ( .A1(n146), .A2(n145), .ZN(n147) );
  OR2_X1 U82bar ( .A1(n146bar), .A2(n145bar), .ZN(n147bar) );
  OR2_X1 U83 ( .A1(n193), .A2(d[4]), .ZN(n145) );
  AND2_X1 U83bar ( .A1(n193bar), .A2(dbar[4]), .ZN(n145bar) );
  OR2_X1 U84 ( .A1(n181), .A2(c[4]), .ZN(n146) );
  AND2_X1 U84bar ( .A1(n181bar), .A2(cbar[4]), .ZN(n146bar) );
  OR2_X1 U85 ( .A1(n144), .A2(n216), .ZN(y[3]) );
  AND2_X1 U85bar ( .A1(n144bar), .A2(n216bar), .ZN(ybar[3]) );
  OR2_X1 U86 ( .A1(n142), .A2(n192), .ZN(n143) );
  AND2_X1 U86bar ( .A1(n142bar), .A2(n192bar), .ZN(n143bar) );
  AND2_X1 U87 ( .A1(n192), .A2(n142), .ZN(n144) );
  OR2_X1 U87bar ( .A1(n192bar), .A2(n142bar), .ZN(n144bar) );
  AND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(n142) );
  OR2_X1 U88bar ( .A1(n141bar), .A2(n140bar), .ZN(n142bar) );
  OR2_X1 U89 ( .A1(n215), .A2(b[3]), .ZN(n140) );
  AND2_X1 U89bar ( .A1(n215bar), .A2(bbar[3]), .ZN(n140bar) );
  OR2_X1 U90 ( .A1(n204), .A2(a[3]), .ZN(n141) );
  AND2_X1 U90bar ( .A1(n204bar), .A2(abar[3]), .ZN(n141bar) );
  AND2_X1 U91 ( .A1(n138), .A2(n137), .ZN(n139) );
  OR2_X1 U91bar ( .A1(n138bar), .A2(n137bar), .ZN(n139bar) );
  OR2_X1 U92 ( .A1(n191), .A2(d[3]), .ZN(n137) );
  AND2_X1 U92bar ( .A1(n191bar), .A2(dbar[3]), .ZN(n137bar) );
  OR2_X1 U93 ( .A1(n180), .A2(c[3]), .ZN(n138) );
  AND2_X1 U93bar ( .A1(n180bar), .A2(cbar[3]), .ZN(n138bar) );
  OR2_X1 U94 ( .A1(n136), .A2(n214), .ZN(y[2]) );
  AND2_X1 U94bar ( .A1(n136bar), .A2(n214bar), .ZN(ybar[2]) );
  OR2_X1 U95 ( .A1(n134), .A2(n190), .ZN(n135) );
  AND2_X1 U95bar ( .A1(n134bar), .A2(n190bar), .ZN(n135bar) );
  AND2_X1 U96 ( .A1(n190), .A2(n134), .ZN(n136) );
  OR2_X1 U96bar ( .A1(n190bar), .A2(n134bar), .ZN(n136bar) );
  AND2_X1 U97 ( .A1(n133), .A2(n132), .ZN(n134) );
  OR2_X1 U97bar ( .A1(n133bar), .A2(n132bar), .ZN(n134bar) );
  OR2_X1 U98 ( .A1(n213), .A2(b[2]), .ZN(n132) );
  AND2_X1 U98bar ( .A1(n213bar), .A2(bbar[2]), .ZN(n132bar) );
  OR2_X1 U99 ( .A1(n203), .A2(a[2]), .ZN(n133) );
  AND2_X1 U99bar ( .A1(n203bar), .A2(abar[2]), .ZN(n133bar) );
  AND2_X1 U100 ( .A1(n130), .A2(n129), .ZN(n131) );
  OR2_X1 U100bar ( .A1(n130bar), .A2(n129bar), .ZN(n131bar) );
  OR2_X1 U101 ( .A1(n189), .A2(d[2]), .ZN(n129) );
  AND2_X1 U101bar ( .A1(n189bar), .A2(dbar[2]), .ZN(n129bar) );
  OR2_X1 U102 ( .A1(n179), .A2(c[2]), .ZN(n130) );
  AND2_X1 U102bar ( .A1(n179bar), .A2(cbar[2]), .ZN(n130bar) );
  OR2_X1 U103 ( .A1(n128), .A2(n212), .ZN(y[1]) );
  AND2_X1 U103bar ( .A1(n128bar), .A2(n212bar), .ZN(ybar[1]) );
  OR2_X1 U104 ( .A1(n126), .A2(n188), .ZN(n127) );
  AND2_X1 U104bar ( .A1(n126bar), .A2(n188bar), .ZN(n127bar) );
  AND2_X1 U105 ( .A1(n188), .A2(n126), .ZN(n128) );
  OR2_X1 U105bar ( .A1(n188bar), .A2(n126bar), .ZN(n128bar) );
  AND2_X1 U106 ( .A1(n125), .A2(n124), .ZN(n126) );
  OR2_X1 U106bar ( .A1(n125bar), .A2(n124bar), .ZN(n126bar) );
  OR2_X1 U107 ( .A1(n211), .A2(b[1]), .ZN(n124) );
  AND2_X1 U107bar ( .A1(n211bar), .A2(bbar[1]), .ZN(n124bar) );
  OR2_X1 U108 ( .A1(n202), .A2(a[1]), .ZN(n125) );
  AND2_X1 U108bar ( .A1(n202bar), .A2(abar[1]), .ZN(n125bar) );
  AND2_X1 U109 ( .A1(n122), .A2(n121), .ZN(n123) );
  OR2_X1 U109bar ( .A1(n122bar), .A2(n121bar), .ZN(n123bar) );
  OR2_X1 U110 ( .A1(n187), .A2(d[1]), .ZN(n121) );
  AND2_X1 U110bar ( .A1(n187bar), .A2(dbar[1]), .ZN(n121bar) );
  OR2_X1 U111 ( .A1(n178), .A2(c[1]), .ZN(n122) );
  AND2_X1 U111bar ( .A1(n178bar), .A2(cbar[1]), .ZN(n122bar) );
  OR2_X1 U112 ( .A1(n120), .A2(n210), .ZN(y[0]) );
  AND2_X1 U112bar ( .A1(n120bar), .A2(n210bar), .ZN(ybar[0]) );
  OR2_X1 U113 ( .A1(n118), .A2(n186), .ZN(n119) );
  AND2_X1 U113bar ( .A1(n118bar), .A2(n186bar), .ZN(n119bar) );
  AND2_X1 U114 ( .A1(n186), .A2(n118), .ZN(n120) );
  OR2_X1 U114bar ( .A1(n186bar), .A2(n118bar), .ZN(n120bar) );
  AND2_X1 U115 ( .A1(n117), .A2(n116), .ZN(n118) );
  OR2_X1 U115bar ( .A1(n117bar), .A2(n116bar), .ZN(n118bar) );
  OR2_X1 U116 ( .A1(n209), .A2(b[0]), .ZN(n116) );
  AND2_X1 U116bar ( .A1(n209bar), .A2(bbar[0]), .ZN(n116bar) );
  OR2_X1 U117 ( .A1(n201), .A2(a[0]), .ZN(n117) );
  AND2_X1 U117bar ( .A1(n201bar), .A2(abar[0]), .ZN(n117bar) );
  AND2_X1 U118 ( .A1(n114), .A2(n113), .ZN(n115) );
  OR2_X1 U118bar ( .A1(n114bar), .A2(n113bar), .ZN(n115bar) );
  OR2_X1 U119 ( .A1(n185), .A2(d[0]), .ZN(n113) );
  AND2_X1 U119bar ( .A1(n185bar), .A2(dbar[0]), .ZN(n113bar) );
  OR2_X1 U120 ( .A1(n177), .A2(c[0]), .ZN(n114) );
  AND2_X1 U120bar ( .A1(n177bar), .A2(cbar[0]), .ZN(n114bar) );
endmodule

module byteXor4_10 ( a, abar, b, bbar, c, cbar, d, dbar, y, ybar );

  input wire [7:0] a;
  input wire [7:0] b;
  input wire [7:0] c;
  input wire [7:0] d;
  input wire [7:0] abar;
  input wire [7:0] bbar;
  input wire [7:0] cbar;
  input wire [7:0] dbar;
//input_done

  output wire [7:0] y;
  output wire [7:0] ybar;
//output_done

  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n113bar;
  wire n114bar;
  wire n115bar;
  wire n116bar;
  wire n117bar;
  wire n118bar;
  wire n119bar;
  wire n120bar;
  wire n121bar;
  wire n122bar;
  wire n123bar;
  wire n124bar;
  wire n125bar;
  wire n126bar;
  wire n127bar;
  wire n128bar;
  wire n129bar;
  wire n130bar;
  wire n131bar;
  wire n132bar;
  wire n133bar;
  wire n134bar;
  wire n135bar;
  wire n136bar;
  wire n137bar;
  wire n138bar;
  wire n139bar;
  wire n140bar;
  wire n141bar;
  wire n142bar;
  wire n143bar;
  wire n144bar;
  wire n145bar;
  wire n146bar;
  wire n147bar;
  wire n148bar;
  wire n149bar;
  wire n150bar;
  wire n151bar;
  wire n152bar;
  wire n153bar;
  wire n154bar;
  wire n155bar;
  wire n156bar;
  wire n157bar;
  wire n158bar;
  wire n159bar;
  wire n160bar;
  wire n161bar;
  wire n162bar;
  wire n163bar;
  wire n164bar;
  wire n165bar;
  wire n166bar;
  wire n167bar;
  wire n168bar;
  wire n169bar;
  wire n170bar;
  wire n171bar;
  wire n172bar;
  wire n173bar;
  wire n174bar;
  wire n175bar;
  wire n176bar;
  wire n177bar;
  wire n178bar;
  wire n179bar;
  wire n180bar;
  wire n181bar;
  wire n182bar;
  wire n183bar;
  wire n184bar;
  wire n185bar;
  wire n186bar;
  wire n187bar;
  wire n188bar;
  wire n189bar;
  wire n190bar;
  wire n191bar;
  wire n192bar;
  wire n193bar;
  wire n194bar;
  wire n195bar;
  wire n196bar;
  wire n197bar;
  wire n198bar;
  wire n199bar;
  wire n200bar;
  wire n201bar;
  wire n202bar;
  wire n203bar;
  wire n204bar;
  wire n205bar;
  wire n206bar;
  wire n207bar;
  wire n208bar;
  wire n209bar;
  wire n210bar;
  wire n211bar;
  wire n212bar;
  wire n213bar;
  wire n214bar;
  wire n215bar;
  wire n216bar;
  wire n217bar;
  wire n218bar;
  wire n219bar;
  wire n220bar;
  wire n221bar;
  wire n222bar;
  wire n223bar;
  wire n224bar;
//wire_done

 //assign_done

  assign n224bar = n175;
  assign n224 = n175bar;
  assign n223bar = a[7];
  assign n223 = abar[7];
  assign n222bar = n167;
  assign n222 = n167bar;
  assign n221bar = a[6];
  assign n221 = abar[6];
  assign n220bar = n159;
  assign n220 = n159bar;
  assign n219bar = a[5];
  assign n219 = abar[5];
  assign n218bar = n151;
  assign n218 = n151bar;
  assign n217bar = a[4];
  assign n217 = abar[4];
  assign n216bar = n143;
  assign n216 = n143bar;
  assign n215bar = a[3];
  assign n215 = abar[3];
  assign n214bar = n135;
  assign n214 = n135bar;
  assign n213bar = a[2];
  assign n213 = abar[2];
  assign n212bar = n127;
  assign n212 = n127bar;
  assign n211bar = a[1];
  assign n211 = abar[1];
  assign n210bar = n119;
  assign n210 = n119bar;
  assign n209bar = a[0];
  assign n209 = abar[0];
  assign n208bar = b[7];
  assign n208 = bbar[7];
  assign n207bar = b[6];
  assign n207 = bbar[6];
  assign n206bar = b[5];
  assign n206 = bbar[5];
  assign n205bar = b[4];
  assign n205 = bbar[4];
  assign n204bar = b[3];
  assign n204 = bbar[3];
  assign n203bar = b[2];
  assign n203 = bbar[2];
  assign n202bar = b[1];
  assign n202 = bbar[1];
  assign n201bar = b[0];
  assign n201 = bbar[0];
  assign n200bar = n171;
  assign n200 = n171bar;
  assign n199bar = c[7];
  assign n199 = cbar[7];
  assign n198bar = n163;
  assign n198 = n163bar;
  assign n197bar = c[6];
  assign n197 = cbar[6];
  assign n196bar = n155;
  assign n196 = n155bar;
  assign n195bar = c[5];
  assign n195 = cbar[5];
  assign n194bar = n147;
  assign n194 = n147bar;
  assign n193bar = c[4];
  assign n193 = cbar[4];
  assign n192bar = n139;
  assign n192 = n139bar;
  assign n191bar = c[3];
  assign n191 = cbar[3];
  assign n190bar = n131;
  assign n190 = n131bar;
  assign n189bar = c[2];
  assign n189 = cbar[2];
  assign n188bar = n123;
  assign n188 = n123bar;
  assign n187bar = c[1];
  assign n187 = cbar[1];
  assign n186bar = n115;
  assign n186 = n115bar;
  assign n185bar = c[0];
  assign n185 = cbar[0];
  assign n184bar = d[7];
  assign n184 = dbar[7];
  assign n183bar = d[6];
  assign n183 = dbar[6];
  assign n182bar = d[5];
  assign n182 = dbar[5];
  assign n181bar = d[4];
  assign n181 = dbar[4];
  assign n180bar = d[3];
  assign n180 = dbar[3];
  assign n179bar = d[2];
  assign n179 = dbar[2];
  assign n178bar = d[1];
  assign n178 = dbar[1];
  assign n177bar = d[0];
  assign n177 = dbar[0];
  OR2_X1 U49 ( .A1(n176), .A2(n224), .ZN(y[7]) );
  AND2_X1 U49bar ( .A1(n176bar), .A2(n224bar), .ZN(ybar[7]) );
  OR2_X1 U50 ( .A1(n174), .A2(n200), .ZN(n175) );
  AND2_X1 U50bar ( .A1(n174bar), .A2(n200bar), .ZN(n175bar) );
  AND2_X1 U51 ( .A1(n200), .A2(n174), .ZN(n176) );
  OR2_X1 U51bar ( .A1(n200bar), .A2(n174bar), .ZN(n176bar) );
  AND2_X1 U52 ( .A1(n173), .A2(n172), .ZN(n174) );
  OR2_X1 U52bar ( .A1(n173bar), .A2(n172bar), .ZN(n174bar) );
  OR2_X1 U53 ( .A1(n223), .A2(b[7]), .ZN(n172) );
  AND2_X1 U53bar ( .A1(n223bar), .A2(bbar[7]), .ZN(n172bar) );
  OR2_X1 U54 ( .A1(n208), .A2(a[7]), .ZN(n173) );
  AND2_X1 U54bar ( .A1(n208bar), .A2(abar[7]), .ZN(n173bar) );
  AND2_X1 U55 ( .A1(n170), .A2(n169), .ZN(n171) );
  OR2_X1 U55bar ( .A1(n170bar), .A2(n169bar), .ZN(n171bar) );
  OR2_X1 U56 ( .A1(n199), .A2(d[7]), .ZN(n169) );
  AND2_X1 U56bar ( .A1(n199bar), .A2(dbar[7]), .ZN(n169bar) );
  OR2_X1 U57 ( .A1(n184), .A2(c[7]), .ZN(n170) );
  AND2_X1 U57bar ( .A1(n184bar), .A2(cbar[7]), .ZN(n170bar) );
  OR2_X1 U58 ( .A1(n168), .A2(n222), .ZN(y[6]) );
  AND2_X1 U58bar ( .A1(n168bar), .A2(n222bar), .ZN(ybar[6]) );
  OR2_X1 U59 ( .A1(n166), .A2(n198), .ZN(n167) );
  AND2_X1 U59bar ( .A1(n166bar), .A2(n198bar), .ZN(n167bar) );
  AND2_X1 U60 ( .A1(n198), .A2(n166), .ZN(n168) );
  OR2_X1 U60bar ( .A1(n198bar), .A2(n166bar), .ZN(n168bar) );
  AND2_X1 U61 ( .A1(n165), .A2(n164), .ZN(n166) );
  OR2_X1 U61bar ( .A1(n165bar), .A2(n164bar), .ZN(n166bar) );
  OR2_X1 U62 ( .A1(n221), .A2(b[6]), .ZN(n164) );
  AND2_X1 U62bar ( .A1(n221bar), .A2(bbar[6]), .ZN(n164bar) );
  OR2_X1 U63 ( .A1(n207), .A2(a[6]), .ZN(n165) );
  AND2_X1 U63bar ( .A1(n207bar), .A2(abar[6]), .ZN(n165bar) );
  AND2_X1 U64 ( .A1(n162), .A2(n161), .ZN(n163) );
  OR2_X1 U64bar ( .A1(n162bar), .A2(n161bar), .ZN(n163bar) );
  OR2_X1 U65 ( .A1(n197), .A2(d[6]), .ZN(n161) );
  AND2_X1 U65bar ( .A1(n197bar), .A2(dbar[6]), .ZN(n161bar) );
  OR2_X1 U66 ( .A1(n183), .A2(c[6]), .ZN(n162) );
  AND2_X1 U66bar ( .A1(n183bar), .A2(cbar[6]), .ZN(n162bar) );
  OR2_X1 U67 ( .A1(n160), .A2(n220), .ZN(y[5]) );
  AND2_X1 U67bar ( .A1(n160bar), .A2(n220bar), .ZN(ybar[5]) );
  OR2_X1 U68 ( .A1(n158), .A2(n196), .ZN(n159) );
  AND2_X1 U68bar ( .A1(n158bar), .A2(n196bar), .ZN(n159bar) );
  AND2_X1 U69 ( .A1(n196), .A2(n158), .ZN(n160) );
  OR2_X1 U69bar ( .A1(n196bar), .A2(n158bar), .ZN(n160bar) );
  AND2_X1 U70 ( .A1(n157), .A2(n156), .ZN(n158) );
  OR2_X1 U70bar ( .A1(n157bar), .A2(n156bar), .ZN(n158bar) );
  OR2_X1 U71 ( .A1(n219), .A2(b[5]), .ZN(n156) );
  AND2_X1 U71bar ( .A1(n219bar), .A2(bbar[5]), .ZN(n156bar) );
  OR2_X1 U72 ( .A1(n206), .A2(a[5]), .ZN(n157) );
  AND2_X1 U72bar ( .A1(n206bar), .A2(abar[5]), .ZN(n157bar) );
  AND2_X1 U73 ( .A1(n154), .A2(n153), .ZN(n155) );
  OR2_X1 U73bar ( .A1(n154bar), .A2(n153bar), .ZN(n155bar) );
  OR2_X1 U74 ( .A1(n195), .A2(d[5]), .ZN(n153) );
  AND2_X1 U74bar ( .A1(n195bar), .A2(dbar[5]), .ZN(n153bar) );
  OR2_X1 U75 ( .A1(n182), .A2(c[5]), .ZN(n154) );
  AND2_X1 U75bar ( .A1(n182bar), .A2(cbar[5]), .ZN(n154bar) );
  OR2_X1 U76 ( .A1(n152), .A2(n218), .ZN(y[4]) );
  AND2_X1 U76bar ( .A1(n152bar), .A2(n218bar), .ZN(ybar[4]) );
  OR2_X1 U77 ( .A1(n150), .A2(n194), .ZN(n151) );
  AND2_X1 U77bar ( .A1(n150bar), .A2(n194bar), .ZN(n151bar) );
  AND2_X1 U78 ( .A1(n194), .A2(n150), .ZN(n152) );
  OR2_X1 U78bar ( .A1(n194bar), .A2(n150bar), .ZN(n152bar) );
  AND2_X1 U79 ( .A1(n149), .A2(n148), .ZN(n150) );
  OR2_X1 U79bar ( .A1(n149bar), .A2(n148bar), .ZN(n150bar) );
  OR2_X1 U80 ( .A1(n217), .A2(b[4]), .ZN(n148) );
  AND2_X1 U80bar ( .A1(n217bar), .A2(bbar[4]), .ZN(n148bar) );
  OR2_X1 U81 ( .A1(n205), .A2(a[4]), .ZN(n149) );
  AND2_X1 U81bar ( .A1(n205bar), .A2(abar[4]), .ZN(n149bar) );
  AND2_X1 U82 ( .A1(n146), .A2(n145), .ZN(n147) );
  OR2_X1 U82bar ( .A1(n146bar), .A2(n145bar), .ZN(n147bar) );
  OR2_X1 U83 ( .A1(n193), .A2(d[4]), .ZN(n145) );
  AND2_X1 U83bar ( .A1(n193bar), .A2(dbar[4]), .ZN(n145bar) );
  OR2_X1 U84 ( .A1(n181), .A2(c[4]), .ZN(n146) );
  AND2_X1 U84bar ( .A1(n181bar), .A2(cbar[4]), .ZN(n146bar) );
  OR2_X1 U85 ( .A1(n144), .A2(n216), .ZN(y[3]) );
  AND2_X1 U85bar ( .A1(n144bar), .A2(n216bar), .ZN(ybar[3]) );
  OR2_X1 U86 ( .A1(n142), .A2(n192), .ZN(n143) );
  AND2_X1 U86bar ( .A1(n142bar), .A2(n192bar), .ZN(n143bar) );
  AND2_X1 U87 ( .A1(n192), .A2(n142), .ZN(n144) );
  OR2_X1 U87bar ( .A1(n192bar), .A2(n142bar), .ZN(n144bar) );
  AND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(n142) );
  OR2_X1 U88bar ( .A1(n141bar), .A2(n140bar), .ZN(n142bar) );
  OR2_X1 U89 ( .A1(n215), .A2(b[3]), .ZN(n140) );
  AND2_X1 U89bar ( .A1(n215bar), .A2(bbar[3]), .ZN(n140bar) );
  OR2_X1 U90 ( .A1(n204), .A2(a[3]), .ZN(n141) );
  AND2_X1 U90bar ( .A1(n204bar), .A2(abar[3]), .ZN(n141bar) );
  AND2_X1 U91 ( .A1(n138), .A2(n137), .ZN(n139) );
  OR2_X1 U91bar ( .A1(n138bar), .A2(n137bar), .ZN(n139bar) );
  OR2_X1 U92 ( .A1(n191), .A2(d[3]), .ZN(n137) );
  AND2_X1 U92bar ( .A1(n191bar), .A2(dbar[3]), .ZN(n137bar) );
  OR2_X1 U93 ( .A1(n180), .A2(c[3]), .ZN(n138) );
  AND2_X1 U93bar ( .A1(n180bar), .A2(cbar[3]), .ZN(n138bar) );
  OR2_X1 U94 ( .A1(n136), .A2(n214), .ZN(y[2]) );
  AND2_X1 U94bar ( .A1(n136bar), .A2(n214bar), .ZN(ybar[2]) );
  OR2_X1 U95 ( .A1(n134), .A2(n190), .ZN(n135) );
  AND2_X1 U95bar ( .A1(n134bar), .A2(n190bar), .ZN(n135bar) );
  AND2_X1 U96 ( .A1(n190), .A2(n134), .ZN(n136) );
  OR2_X1 U96bar ( .A1(n190bar), .A2(n134bar), .ZN(n136bar) );
  AND2_X1 U97 ( .A1(n133), .A2(n132), .ZN(n134) );
  OR2_X1 U97bar ( .A1(n133bar), .A2(n132bar), .ZN(n134bar) );
  OR2_X1 U98 ( .A1(n213), .A2(b[2]), .ZN(n132) );
  AND2_X1 U98bar ( .A1(n213bar), .A2(bbar[2]), .ZN(n132bar) );
  OR2_X1 U99 ( .A1(n203), .A2(a[2]), .ZN(n133) );
  AND2_X1 U99bar ( .A1(n203bar), .A2(abar[2]), .ZN(n133bar) );
  AND2_X1 U100 ( .A1(n130), .A2(n129), .ZN(n131) );
  OR2_X1 U100bar ( .A1(n130bar), .A2(n129bar), .ZN(n131bar) );
  OR2_X1 U101 ( .A1(n189), .A2(d[2]), .ZN(n129) );
  AND2_X1 U101bar ( .A1(n189bar), .A2(dbar[2]), .ZN(n129bar) );
  OR2_X1 U102 ( .A1(n179), .A2(c[2]), .ZN(n130) );
  AND2_X1 U102bar ( .A1(n179bar), .A2(cbar[2]), .ZN(n130bar) );
  OR2_X1 U103 ( .A1(n128), .A2(n212), .ZN(y[1]) );
  AND2_X1 U103bar ( .A1(n128bar), .A2(n212bar), .ZN(ybar[1]) );
  OR2_X1 U104 ( .A1(n126), .A2(n188), .ZN(n127) );
  AND2_X1 U104bar ( .A1(n126bar), .A2(n188bar), .ZN(n127bar) );
  AND2_X1 U105 ( .A1(n188), .A2(n126), .ZN(n128) );
  OR2_X1 U105bar ( .A1(n188bar), .A2(n126bar), .ZN(n128bar) );
  AND2_X1 U106 ( .A1(n125), .A2(n124), .ZN(n126) );
  OR2_X1 U106bar ( .A1(n125bar), .A2(n124bar), .ZN(n126bar) );
  OR2_X1 U107 ( .A1(n211), .A2(b[1]), .ZN(n124) );
  AND2_X1 U107bar ( .A1(n211bar), .A2(bbar[1]), .ZN(n124bar) );
  OR2_X1 U108 ( .A1(n202), .A2(a[1]), .ZN(n125) );
  AND2_X1 U108bar ( .A1(n202bar), .A2(abar[1]), .ZN(n125bar) );
  AND2_X1 U109 ( .A1(n122), .A2(n121), .ZN(n123) );
  OR2_X1 U109bar ( .A1(n122bar), .A2(n121bar), .ZN(n123bar) );
  OR2_X1 U110 ( .A1(n187), .A2(d[1]), .ZN(n121) );
  AND2_X1 U110bar ( .A1(n187bar), .A2(dbar[1]), .ZN(n121bar) );
  OR2_X1 U111 ( .A1(n178), .A2(c[1]), .ZN(n122) );
  AND2_X1 U111bar ( .A1(n178bar), .A2(cbar[1]), .ZN(n122bar) );
  OR2_X1 U112 ( .A1(n120), .A2(n210), .ZN(y[0]) );
  AND2_X1 U112bar ( .A1(n120bar), .A2(n210bar), .ZN(ybar[0]) );
  OR2_X1 U113 ( .A1(n118), .A2(n186), .ZN(n119) );
  AND2_X1 U113bar ( .A1(n118bar), .A2(n186bar), .ZN(n119bar) );
  AND2_X1 U114 ( .A1(n186), .A2(n118), .ZN(n120) );
  OR2_X1 U114bar ( .A1(n186bar), .A2(n118bar), .ZN(n120bar) );
  AND2_X1 U115 ( .A1(n117), .A2(n116), .ZN(n118) );
  OR2_X1 U115bar ( .A1(n117bar), .A2(n116bar), .ZN(n118bar) );
  OR2_X1 U116 ( .A1(n209), .A2(b[0]), .ZN(n116) );
  AND2_X1 U116bar ( .A1(n209bar), .A2(bbar[0]), .ZN(n116bar) );
  OR2_X1 U117 ( .A1(n201), .A2(a[0]), .ZN(n117) );
  AND2_X1 U117bar ( .A1(n201bar), .A2(abar[0]), .ZN(n117bar) );
  AND2_X1 U118 ( .A1(n114), .A2(n113), .ZN(n115) );
  OR2_X1 U118bar ( .A1(n114bar), .A2(n113bar), .ZN(n115bar) );
  OR2_X1 U119 ( .A1(n185), .A2(d[0]), .ZN(n113) );
  AND2_X1 U119bar ( .A1(n185bar), .A2(dbar[0]), .ZN(n113bar) );
  OR2_X1 U120 ( .A1(n177), .A2(c[0]), .ZN(n114) );
  AND2_X1 U120bar ( .A1(n177bar), .A2(cbar[0]), .ZN(n114bar) );
endmodule

module byteXor4_11 ( a, abar, b, bbar, c, cbar, d, dbar, y, ybar );

  input wire [7:0] a;
  input wire [7:0] b;
  input wire [7:0] c;
  input wire [7:0] d;
  input wire [7:0] abar;
  input wire [7:0] bbar;
  input wire [7:0] cbar;
  input wire [7:0] dbar;
//input_done

  output wire [7:0] y;
  output wire [7:0] ybar;
//output_done

  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n113bar;
  wire n114bar;
  wire n115bar;
  wire n116bar;
  wire n117bar;
  wire n118bar;
  wire n119bar;
  wire n120bar;
  wire n121bar;
  wire n122bar;
  wire n123bar;
  wire n124bar;
  wire n125bar;
  wire n126bar;
  wire n127bar;
  wire n128bar;
  wire n129bar;
  wire n130bar;
  wire n131bar;
  wire n132bar;
  wire n133bar;
  wire n134bar;
  wire n135bar;
  wire n136bar;
  wire n137bar;
  wire n138bar;
  wire n139bar;
  wire n140bar;
  wire n141bar;
  wire n142bar;
  wire n143bar;
  wire n144bar;
  wire n145bar;
  wire n146bar;
  wire n147bar;
  wire n148bar;
  wire n149bar;
  wire n150bar;
  wire n151bar;
  wire n152bar;
  wire n153bar;
  wire n154bar;
  wire n155bar;
  wire n156bar;
  wire n157bar;
  wire n158bar;
  wire n159bar;
  wire n160bar;
  wire n161bar;
  wire n162bar;
  wire n163bar;
  wire n164bar;
  wire n165bar;
  wire n166bar;
  wire n167bar;
  wire n168bar;
  wire n169bar;
  wire n170bar;
  wire n171bar;
  wire n172bar;
  wire n173bar;
  wire n174bar;
  wire n175bar;
  wire n176bar;
  wire n177bar;
  wire n178bar;
  wire n179bar;
  wire n180bar;
  wire n181bar;
  wire n182bar;
  wire n183bar;
  wire n184bar;
  wire n185bar;
  wire n186bar;
  wire n187bar;
  wire n188bar;
  wire n189bar;
  wire n190bar;
  wire n191bar;
  wire n192bar;
  wire n193bar;
  wire n194bar;
  wire n195bar;
  wire n196bar;
  wire n197bar;
  wire n198bar;
  wire n199bar;
  wire n200bar;
  wire n201bar;
  wire n202bar;
  wire n203bar;
  wire n204bar;
  wire n205bar;
  wire n206bar;
  wire n207bar;
  wire n208bar;
  wire n209bar;
  wire n210bar;
  wire n211bar;
  wire n212bar;
  wire n213bar;
  wire n214bar;
  wire n215bar;
  wire n216bar;
  wire n217bar;
  wire n218bar;
  wire n219bar;
  wire n220bar;
  wire n221bar;
  wire n222bar;
  wire n223bar;
  wire n224bar;
//wire_done

 //assign_done

  assign n224bar = n175;
  assign n224 = n175bar;
  assign n223bar = a[7];
  assign n223 = abar[7];
  assign n222bar = n167;
  assign n222 = n167bar;
  assign n221bar = a[6];
  assign n221 = abar[6];
  assign n220bar = n159;
  assign n220 = n159bar;
  assign n219bar = a[5];
  assign n219 = abar[5];
  assign n218bar = n151;
  assign n218 = n151bar;
  assign n217bar = a[4];
  assign n217 = abar[4];
  assign n216bar = n143;
  assign n216 = n143bar;
  assign n215bar = a[3];
  assign n215 = abar[3];
  assign n214bar = n135;
  assign n214 = n135bar;
  assign n213bar = a[2];
  assign n213 = abar[2];
  assign n212bar = n127;
  assign n212 = n127bar;
  assign n211bar = a[1];
  assign n211 = abar[1];
  assign n210bar = n119;
  assign n210 = n119bar;
  assign n209bar = a[0];
  assign n209 = abar[0];
  assign n208bar = b[7];
  assign n208 = bbar[7];
  assign n207bar = b[6];
  assign n207 = bbar[6];
  assign n206bar = b[5];
  assign n206 = bbar[5];
  assign n205bar = b[4];
  assign n205 = bbar[4];
  assign n204bar = b[3];
  assign n204 = bbar[3];
  assign n203bar = b[2];
  assign n203 = bbar[2];
  assign n202bar = b[1];
  assign n202 = bbar[1];
  assign n201bar = b[0];
  assign n201 = bbar[0];
  assign n200bar = n171;
  assign n200 = n171bar;
  assign n199bar = c[7];
  assign n199 = cbar[7];
  assign n198bar = n163;
  assign n198 = n163bar;
  assign n197bar = c[6];
  assign n197 = cbar[6];
  assign n196bar = n155;
  assign n196 = n155bar;
  assign n195bar = c[5];
  assign n195 = cbar[5];
  assign n194bar = n147;
  assign n194 = n147bar;
  assign n193bar = c[4];
  assign n193 = cbar[4];
  assign n192bar = n139;
  assign n192 = n139bar;
  assign n191bar = c[3];
  assign n191 = cbar[3];
  assign n190bar = n131;
  assign n190 = n131bar;
  assign n189bar = c[2];
  assign n189 = cbar[2];
  assign n188bar = n123;
  assign n188 = n123bar;
  assign n187bar = c[1];
  assign n187 = cbar[1];
  assign n186bar = n115;
  assign n186 = n115bar;
  assign n185bar = c[0];
  assign n185 = cbar[0];
  assign n184bar = d[7];
  assign n184 = dbar[7];
  assign n183bar = d[6];
  assign n183 = dbar[6];
  assign n182bar = d[5];
  assign n182 = dbar[5];
  assign n181bar = d[4];
  assign n181 = dbar[4];
  assign n180bar = d[3];
  assign n180 = dbar[3];
  assign n179bar = d[2];
  assign n179 = dbar[2];
  assign n178bar = d[1];
  assign n178 = dbar[1];
  assign n177bar = d[0];
  assign n177 = dbar[0];
  OR2_X1 U49 ( .A1(n176), .A2(n224), .ZN(y[7]) );
  AND2_X1 U49bar ( .A1(n176bar), .A2(n224bar), .ZN(ybar[7]) );
  OR2_X1 U50 ( .A1(n174), .A2(n200), .ZN(n175) );
  AND2_X1 U50bar ( .A1(n174bar), .A2(n200bar), .ZN(n175bar) );
  AND2_X1 U51 ( .A1(n200), .A2(n174), .ZN(n176) );
  OR2_X1 U51bar ( .A1(n200bar), .A2(n174bar), .ZN(n176bar) );
  AND2_X1 U52 ( .A1(n173), .A2(n172), .ZN(n174) );
  OR2_X1 U52bar ( .A1(n173bar), .A2(n172bar), .ZN(n174bar) );
  OR2_X1 U53 ( .A1(n223), .A2(b[7]), .ZN(n172) );
  AND2_X1 U53bar ( .A1(n223bar), .A2(bbar[7]), .ZN(n172bar) );
  OR2_X1 U54 ( .A1(n208), .A2(a[7]), .ZN(n173) );
  AND2_X1 U54bar ( .A1(n208bar), .A2(abar[7]), .ZN(n173bar) );
  AND2_X1 U55 ( .A1(n170), .A2(n169), .ZN(n171) );
  OR2_X1 U55bar ( .A1(n170bar), .A2(n169bar), .ZN(n171bar) );
  OR2_X1 U56 ( .A1(n199), .A2(d[7]), .ZN(n169) );
  AND2_X1 U56bar ( .A1(n199bar), .A2(dbar[7]), .ZN(n169bar) );
  OR2_X1 U57 ( .A1(n184), .A2(c[7]), .ZN(n170) );
  AND2_X1 U57bar ( .A1(n184bar), .A2(cbar[7]), .ZN(n170bar) );
  OR2_X1 U58 ( .A1(n168), .A2(n222), .ZN(y[6]) );
  AND2_X1 U58bar ( .A1(n168bar), .A2(n222bar), .ZN(ybar[6]) );
  OR2_X1 U59 ( .A1(n166), .A2(n198), .ZN(n167) );
  AND2_X1 U59bar ( .A1(n166bar), .A2(n198bar), .ZN(n167bar) );
  AND2_X1 U60 ( .A1(n198), .A2(n166), .ZN(n168) );
  OR2_X1 U60bar ( .A1(n198bar), .A2(n166bar), .ZN(n168bar) );
  AND2_X1 U61 ( .A1(n165), .A2(n164), .ZN(n166) );
  OR2_X1 U61bar ( .A1(n165bar), .A2(n164bar), .ZN(n166bar) );
  OR2_X1 U62 ( .A1(n221), .A2(b[6]), .ZN(n164) );
  AND2_X1 U62bar ( .A1(n221bar), .A2(bbar[6]), .ZN(n164bar) );
  OR2_X1 U63 ( .A1(n207), .A2(a[6]), .ZN(n165) );
  AND2_X1 U63bar ( .A1(n207bar), .A2(abar[6]), .ZN(n165bar) );
  AND2_X1 U64 ( .A1(n162), .A2(n161), .ZN(n163) );
  OR2_X1 U64bar ( .A1(n162bar), .A2(n161bar), .ZN(n163bar) );
  OR2_X1 U65 ( .A1(n197), .A2(d[6]), .ZN(n161) );
  AND2_X1 U65bar ( .A1(n197bar), .A2(dbar[6]), .ZN(n161bar) );
  OR2_X1 U66 ( .A1(n183), .A2(c[6]), .ZN(n162) );
  AND2_X1 U66bar ( .A1(n183bar), .A2(cbar[6]), .ZN(n162bar) );
  OR2_X1 U67 ( .A1(n160), .A2(n220), .ZN(y[5]) );
  AND2_X1 U67bar ( .A1(n160bar), .A2(n220bar), .ZN(ybar[5]) );
  OR2_X1 U68 ( .A1(n158), .A2(n196), .ZN(n159) );
  AND2_X1 U68bar ( .A1(n158bar), .A2(n196bar), .ZN(n159bar) );
  AND2_X1 U69 ( .A1(n196), .A2(n158), .ZN(n160) );
  OR2_X1 U69bar ( .A1(n196bar), .A2(n158bar), .ZN(n160bar) );
  AND2_X1 U70 ( .A1(n157), .A2(n156), .ZN(n158) );
  OR2_X1 U70bar ( .A1(n157bar), .A2(n156bar), .ZN(n158bar) );
  OR2_X1 U71 ( .A1(n219), .A2(b[5]), .ZN(n156) );
  AND2_X1 U71bar ( .A1(n219bar), .A2(bbar[5]), .ZN(n156bar) );
  OR2_X1 U72 ( .A1(n206), .A2(a[5]), .ZN(n157) );
  AND2_X1 U72bar ( .A1(n206bar), .A2(abar[5]), .ZN(n157bar) );
  AND2_X1 U73 ( .A1(n154), .A2(n153), .ZN(n155) );
  OR2_X1 U73bar ( .A1(n154bar), .A2(n153bar), .ZN(n155bar) );
  OR2_X1 U74 ( .A1(n195), .A2(d[5]), .ZN(n153) );
  AND2_X1 U74bar ( .A1(n195bar), .A2(dbar[5]), .ZN(n153bar) );
  OR2_X1 U75 ( .A1(n182), .A2(c[5]), .ZN(n154) );
  AND2_X1 U75bar ( .A1(n182bar), .A2(cbar[5]), .ZN(n154bar) );
  OR2_X1 U76 ( .A1(n152), .A2(n218), .ZN(y[4]) );
  AND2_X1 U76bar ( .A1(n152bar), .A2(n218bar), .ZN(ybar[4]) );
  OR2_X1 U77 ( .A1(n150), .A2(n194), .ZN(n151) );
  AND2_X1 U77bar ( .A1(n150bar), .A2(n194bar), .ZN(n151bar) );
  AND2_X1 U78 ( .A1(n194), .A2(n150), .ZN(n152) );
  OR2_X1 U78bar ( .A1(n194bar), .A2(n150bar), .ZN(n152bar) );
  AND2_X1 U79 ( .A1(n149), .A2(n148), .ZN(n150) );
  OR2_X1 U79bar ( .A1(n149bar), .A2(n148bar), .ZN(n150bar) );
  OR2_X1 U80 ( .A1(n217), .A2(b[4]), .ZN(n148) );
  AND2_X1 U80bar ( .A1(n217bar), .A2(bbar[4]), .ZN(n148bar) );
  OR2_X1 U81 ( .A1(n205), .A2(a[4]), .ZN(n149) );
  AND2_X1 U81bar ( .A1(n205bar), .A2(abar[4]), .ZN(n149bar) );
  AND2_X1 U82 ( .A1(n146), .A2(n145), .ZN(n147) );
  OR2_X1 U82bar ( .A1(n146bar), .A2(n145bar), .ZN(n147bar) );
  OR2_X1 U83 ( .A1(n193), .A2(d[4]), .ZN(n145) );
  AND2_X1 U83bar ( .A1(n193bar), .A2(dbar[4]), .ZN(n145bar) );
  OR2_X1 U84 ( .A1(n181), .A2(c[4]), .ZN(n146) );
  AND2_X1 U84bar ( .A1(n181bar), .A2(cbar[4]), .ZN(n146bar) );
  OR2_X1 U85 ( .A1(n144), .A2(n216), .ZN(y[3]) );
  AND2_X1 U85bar ( .A1(n144bar), .A2(n216bar), .ZN(ybar[3]) );
  OR2_X1 U86 ( .A1(n142), .A2(n192), .ZN(n143) );
  AND2_X1 U86bar ( .A1(n142bar), .A2(n192bar), .ZN(n143bar) );
  AND2_X1 U87 ( .A1(n192), .A2(n142), .ZN(n144) );
  OR2_X1 U87bar ( .A1(n192bar), .A2(n142bar), .ZN(n144bar) );
  AND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(n142) );
  OR2_X1 U88bar ( .A1(n141bar), .A2(n140bar), .ZN(n142bar) );
  OR2_X1 U89 ( .A1(n215), .A2(b[3]), .ZN(n140) );
  AND2_X1 U89bar ( .A1(n215bar), .A2(bbar[3]), .ZN(n140bar) );
  OR2_X1 U90 ( .A1(n204), .A2(a[3]), .ZN(n141) );
  AND2_X1 U90bar ( .A1(n204bar), .A2(abar[3]), .ZN(n141bar) );
  AND2_X1 U91 ( .A1(n138), .A2(n137), .ZN(n139) );
  OR2_X1 U91bar ( .A1(n138bar), .A2(n137bar), .ZN(n139bar) );
  OR2_X1 U92 ( .A1(n191), .A2(d[3]), .ZN(n137) );
  AND2_X1 U92bar ( .A1(n191bar), .A2(dbar[3]), .ZN(n137bar) );
  OR2_X1 U93 ( .A1(n180), .A2(c[3]), .ZN(n138) );
  AND2_X1 U93bar ( .A1(n180bar), .A2(cbar[3]), .ZN(n138bar) );
  OR2_X1 U94 ( .A1(n136), .A2(n214), .ZN(y[2]) );
  AND2_X1 U94bar ( .A1(n136bar), .A2(n214bar), .ZN(ybar[2]) );
  OR2_X1 U95 ( .A1(n134), .A2(n190), .ZN(n135) );
  AND2_X1 U95bar ( .A1(n134bar), .A2(n190bar), .ZN(n135bar) );
  AND2_X1 U96 ( .A1(n190), .A2(n134), .ZN(n136) );
  OR2_X1 U96bar ( .A1(n190bar), .A2(n134bar), .ZN(n136bar) );
  AND2_X1 U97 ( .A1(n133), .A2(n132), .ZN(n134) );
  OR2_X1 U97bar ( .A1(n133bar), .A2(n132bar), .ZN(n134bar) );
  OR2_X1 U98 ( .A1(n213), .A2(b[2]), .ZN(n132) );
  AND2_X1 U98bar ( .A1(n213bar), .A2(bbar[2]), .ZN(n132bar) );
  OR2_X1 U99 ( .A1(n203), .A2(a[2]), .ZN(n133) );
  AND2_X1 U99bar ( .A1(n203bar), .A2(abar[2]), .ZN(n133bar) );
  AND2_X1 U100 ( .A1(n130), .A2(n129), .ZN(n131) );
  OR2_X1 U100bar ( .A1(n130bar), .A2(n129bar), .ZN(n131bar) );
  OR2_X1 U101 ( .A1(n189), .A2(d[2]), .ZN(n129) );
  AND2_X1 U101bar ( .A1(n189bar), .A2(dbar[2]), .ZN(n129bar) );
  OR2_X1 U102 ( .A1(n179), .A2(c[2]), .ZN(n130) );
  AND2_X1 U102bar ( .A1(n179bar), .A2(cbar[2]), .ZN(n130bar) );
  OR2_X1 U103 ( .A1(n128), .A2(n212), .ZN(y[1]) );
  AND2_X1 U103bar ( .A1(n128bar), .A2(n212bar), .ZN(ybar[1]) );
  OR2_X1 U104 ( .A1(n126), .A2(n188), .ZN(n127) );
  AND2_X1 U104bar ( .A1(n126bar), .A2(n188bar), .ZN(n127bar) );
  AND2_X1 U105 ( .A1(n188), .A2(n126), .ZN(n128) );
  OR2_X1 U105bar ( .A1(n188bar), .A2(n126bar), .ZN(n128bar) );
  AND2_X1 U106 ( .A1(n125), .A2(n124), .ZN(n126) );
  OR2_X1 U106bar ( .A1(n125bar), .A2(n124bar), .ZN(n126bar) );
  OR2_X1 U107 ( .A1(n211), .A2(b[1]), .ZN(n124) );
  AND2_X1 U107bar ( .A1(n211bar), .A2(bbar[1]), .ZN(n124bar) );
  OR2_X1 U108 ( .A1(n202), .A2(a[1]), .ZN(n125) );
  AND2_X1 U108bar ( .A1(n202bar), .A2(abar[1]), .ZN(n125bar) );
  AND2_X1 U109 ( .A1(n122), .A2(n121), .ZN(n123) );
  OR2_X1 U109bar ( .A1(n122bar), .A2(n121bar), .ZN(n123bar) );
  OR2_X1 U110 ( .A1(n187), .A2(d[1]), .ZN(n121) );
  AND2_X1 U110bar ( .A1(n187bar), .A2(dbar[1]), .ZN(n121bar) );
  OR2_X1 U111 ( .A1(n178), .A2(c[1]), .ZN(n122) );
  AND2_X1 U111bar ( .A1(n178bar), .A2(cbar[1]), .ZN(n122bar) );
  OR2_X1 U112 ( .A1(n120), .A2(n210), .ZN(y[0]) );
  AND2_X1 U112bar ( .A1(n120bar), .A2(n210bar), .ZN(ybar[0]) );
  OR2_X1 U113 ( .A1(n118), .A2(n186), .ZN(n119) );
  AND2_X1 U113bar ( .A1(n118bar), .A2(n186bar), .ZN(n119bar) );
  AND2_X1 U114 ( .A1(n186), .A2(n118), .ZN(n120) );
  OR2_X1 U114bar ( .A1(n186bar), .A2(n118bar), .ZN(n120bar) );
  AND2_X1 U115 ( .A1(n117), .A2(n116), .ZN(n118) );
  OR2_X1 U115bar ( .A1(n117bar), .A2(n116bar), .ZN(n118bar) );
  OR2_X1 U116 ( .A1(n209), .A2(b[0]), .ZN(n116) );
  AND2_X1 U116bar ( .A1(n209bar), .A2(bbar[0]), .ZN(n116bar) );
  OR2_X1 U117 ( .A1(n201), .A2(a[0]), .ZN(n117) );
  AND2_X1 U117bar ( .A1(n201bar), .A2(abar[0]), .ZN(n117bar) );
  AND2_X1 U118 ( .A1(n114), .A2(n113), .ZN(n115) );
  OR2_X1 U118bar ( .A1(n114bar), .A2(n113bar), .ZN(n115bar) );
  OR2_X1 U119 ( .A1(n185), .A2(d[0]), .ZN(n113) );
  AND2_X1 U119bar ( .A1(n185bar), .A2(dbar[0]), .ZN(n113bar) );
  OR2_X1 U120 ( .A1(n177), .A2(c[0]), .ZN(n114) );
  AND2_X1 U120bar ( .A1(n177bar), .A2(cbar[0]), .ZN(n114bar) );
endmodule

module byteXor4_12 ( a, abar, b, bbar, c, cbar, d, dbar, y, ybar );

  input wire [7:0] a;
  input wire [7:0] b;
  input wire [7:0] c;
  input wire [7:0] d;
  input wire [7:0] abar;
  input wire [7:0] bbar;
  input wire [7:0] cbar;
  input wire [7:0] dbar;
//input_done

  output wire [7:0] y;
  output wire [7:0] ybar;
//output_done

  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n113bar;
  wire n114bar;
  wire n115bar;
  wire n116bar;
  wire n117bar;
  wire n118bar;
  wire n119bar;
  wire n120bar;
  wire n121bar;
  wire n122bar;
  wire n123bar;
  wire n124bar;
  wire n125bar;
  wire n126bar;
  wire n127bar;
  wire n128bar;
  wire n129bar;
  wire n130bar;
  wire n131bar;
  wire n132bar;
  wire n133bar;
  wire n134bar;
  wire n135bar;
  wire n136bar;
  wire n137bar;
  wire n138bar;
  wire n139bar;
  wire n140bar;
  wire n141bar;
  wire n142bar;
  wire n143bar;
  wire n144bar;
  wire n145bar;
  wire n146bar;
  wire n147bar;
  wire n148bar;
  wire n149bar;
  wire n150bar;
  wire n151bar;
  wire n152bar;
  wire n153bar;
  wire n154bar;
  wire n155bar;
  wire n156bar;
  wire n157bar;
  wire n158bar;
  wire n159bar;
  wire n160bar;
  wire n161bar;
  wire n162bar;
  wire n163bar;
  wire n164bar;
  wire n165bar;
  wire n166bar;
  wire n167bar;
  wire n168bar;
  wire n169bar;
  wire n170bar;
  wire n171bar;
  wire n172bar;
  wire n173bar;
  wire n174bar;
  wire n175bar;
  wire n176bar;
  wire n177bar;
  wire n178bar;
  wire n179bar;
  wire n180bar;
  wire n181bar;
  wire n182bar;
  wire n183bar;
  wire n184bar;
  wire n185bar;
  wire n186bar;
  wire n187bar;
  wire n188bar;
  wire n189bar;
  wire n190bar;
  wire n191bar;
  wire n192bar;
  wire n193bar;
  wire n194bar;
  wire n195bar;
  wire n196bar;
  wire n197bar;
  wire n198bar;
  wire n199bar;
  wire n200bar;
  wire n201bar;
  wire n202bar;
  wire n203bar;
  wire n204bar;
  wire n205bar;
  wire n206bar;
  wire n207bar;
  wire n208bar;
  wire n209bar;
  wire n210bar;
  wire n211bar;
  wire n212bar;
  wire n213bar;
  wire n214bar;
  wire n215bar;
  wire n216bar;
  wire n217bar;
  wire n218bar;
  wire n219bar;
  wire n220bar;
  wire n221bar;
  wire n222bar;
  wire n223bar;
  wire n224bar;
//wire_done

 //assign_done

  assign n224bar = n175;
  assign n224 = n175bar;
  assign n223bar = a[7];
  assign n223 = abar[7];
  assign n222bar = n167;
  assign n222 = n167bar;
  assign n221bar = a[6];
  assign n221 = abar[6];
  assign n220bar = n159;
  assign n220 = n159bar;
  assign n219bar = a[5];
  assign n219 = abar[5];
  assign n218bar = n151;
  assign n218 = n151bar;
  assign n217bar = a[4];
  assign n217 = abar[4];
  assign n216bar = n143;
  assign n216 = n143bar;
  assign n215bar = a[3];
  assign n215 = abar[3];
  assign n214bar = n135;
  assign n214 = n135bar;
  assign n213bar = a[2];
  assign n213 = abar[2];
  assign n212bar = n127;
  assign n212 = n127bar;
  assign n211bar = a[1];
  assign n211 = abar[1];
  assign n210bar = n119;
  assign n210 = n119bar;
  assign n209bar = a[0];
  assign n209 = abar[0];
  assign n208bar = b[7];
  assign n208 = bbar[7];
  assign n207bar = b[6];
  assign n207 = bbar[6];
  assign n206bar = b[5];
  assign n206 = bbar[5];
  assign n205bar = b[4];
  assign n205 = bbar[4];
  assign n204bar = b[3];
  assign n204 = bbar[3];
  assign n203bar = b[2];
  assign n203 = bbar[2];
  assign n202bar = b[1];
  assign n202 = bbar[1];
  assign n201bar = b[0];
  assign n201 = bbar[0];
  assign n200bar = n171;
  assign n200 = n171bar;
  assign n199bar = c[7];
  assign n199 = cbar[7];
  assign n198bar = n163;
  assign n198 = n163bar;
  assign n197bar = c[6];
  assign n197 = cbar[6];
  assign n196bar = n155;
  assign n196 = n155bar;
  assign n195bar = c[5];
  assign n195 = cbar[5];
  assign n194bar = n147;
  assign n194 = n147bar;
  assign n193bar = c[4];
  assign n193 = cbar[4];
  assign n192bar = n139;
  assign n192 = n139bar;
  assign n191bar = c[3];
  assign n191 = cbar[3];
  assign n190bar = n131;
  assign n190 = n131bar;
  assign n189bar = c[2];
  assign n189 = cbar[2];
  assign n188bar = n123;
  assign n188 = n123bar;
  assign n187bar = c[1];
  assign n187 = cbar[1];
  assign n186bar = n115;
  assign n186 = n115bar;
  assign n185bar = c[0];
  assign n185 = cbar[0];
  assign n184bar = d[7];
  assign n184 = dbar[7];
  assign n183bar = d[6];
  assign n183 = dbar[6];
  assign n182bar = d[5];
  assign n182 = dbar[5];
  assign n181bar = d[4];
  assign n181 = dbar[4];
  assign n180bar = d[3];
  assign n180 = dbar[3];
  assign n179bar = d[2];
  assign n179 = dbar[2];
  assign n178bar = d[1];
  assign n178 = dbar[1];
  assign n177bar = d[0];
  assign n177 = dbar[0];
  OR2_X1 U49 ( .A1(n176), .A2(n224), .ZN(y[7]) );
  AND2_X1 U49bar ( .A1(n176bar), .A2(n224bar), .ZN(ybar[7]) );
  OR2_X1 U50 ( .A1(n174), .A2(n200), .ZN(n175) );
  AND2_X1 U50bar ( .A1(n174bar), .A2(n200bar), .ZN(n175bar) );
  AND2_X1 U51 ( .A1(n200), .A2(n174), .ZN(n176) );
  OR2_X1 U51bar ( .A1(n200bar), .A2(n174bar), .ZN(n176bar) );
  AND2_X1 U52 ( .A1(n173), .A2(n172), .ZN(n174) );
  OR2_X1 U52bar ( .A1(n173bar), .A2(n172bar), .ZN(n174bar) );
  OR2_X1 U53 ( .A1(n223), .A2(b[7]), .ZN(n172) );
  AND2_X1 U53bar ( .A1(n223bar), .A2(bbar[7]), .ZN(n172bar) );
  OR2_X1 U54 ( .A1(n208), .A2(a[7]), .ZN(n173) );
  AND2_X1 U54bar ( .A1(n208bar), .A2(abar[7]), .ZN(n173bar) );
  AND2_X1 U55 ( .A1(n170), .A2(n169), .ZN(n171) );
  OR2_X1 U55bar ( .A1(n170bar), .A2(n169bar), .ZN(n171bar) );
  OR2_X1 U56 ( .A1(n199), .A2(d[7]), .ZN(n169) );
  AND2_X1 U56bar ( .A1(n199bar), .A2(dbar[7]), .ZN(n169bar) );
  OR2_X1 U57 ( .A1(n184), .A2(c[7]), .ZN(n170) );
  AND2_X1 U57bar ( .A1(n184bar), .A2(cbar[7]), .ZN(n170bar) );
  OR2_X1 U58 ( .A1(n168), .A2(n222), .ZN(y[6]) );
  AND2_X1 U58bar ( .A1(n168bar), .A2(n222bar), .ZN(ybar[6]) );
  OR2_X1 U59 ( .A1(n166), .A2(n198), .ZN(n167) );
  AND2_X1 U59bar ( .A1(n166bar), .A2(n198bar), .ZN(n167bar) );
  AND2_X1 U60 ( .A1(n198), .A2(n166), .ZN(n168) );
  OR2_X1 U60bar ( .A1(n198bar), .A2(n166bar), .ZN(n168bar) );
  AND2_X1 U61 ( .A1(n165), .A2(n164), .ZN(n166) );
  OR2_X1 U61bar ( .A1(n165bar), .A2(n164bar), .ZN(n166bar) );
  OR2_X1 U62 ( .A1(n221), .A2(b[6]), .ZN(n164) );
  AND2_X1 U62bar ( .A1(n221bar), .A2(bbar[6]), .ZN(n164bar) );
  OR2_X1 U63 ( .A1(n207), .A2(a[6]), .ZN(n165) );
  AND2_X1 U63bar ( .A1(n207bar), .A2(abar[6]), .ZN(n165bar) );
  AND2_X1 U64 ( .A1(n162), .A2(n161), .ZN(n163) );
  OR2_X1 U64bar ( .A1(n162bar), .A2(n161bar), .ZN(n163bar) );
  OR2_X1 U65 ( .A1(n197), .A2(d[6]), .ZN(n161) );
  AND2_X1 U65bar ( .A1(n197bar), .A2(dbar[6]), .ZN(n161bar) );
  OR2_X1 U66 ( .A1(n183), .A2(c[6]), .ZN(n162) );
  AND2_X1 U66bar ( .A1(n183bar), .A2(cbar[6]), .ZN(n162bar) );
  OR2_X1 U67 ( .A1(n160), .A2(n220), .ZN(y[5]) );
  AND2_X1 U67bar ( .A1(n160bar), .A2(n220bar), .ZN(ybar[5]) );
  OR2_X1 U68 ( .A1(n158), .A2(n196), .ZN(n159) );
  AND2_X1 U68bar ( .A1(n158bar), .A2(n196bar), .ZN(n159bar) );
  AND2_X1 U69 ( .A1(n196), .A2(n158), .ZN(n160) );
  OR2_X1 U69bar ( .A1(n196bar), .A2(n158bar), .ZN(n160bar) );
  AND2_X1 U70 ( .A1(n157), .A2(n156), .ZN(n158) );
  OR2_X1 U70bar ( .A1(n157bar), .A2(n156bar), .ZN(n158bar) );
  OR2_X1 U71 ( .A1(n219), .A2(b[5]), .ZN(n156) );
  AND2_X1 U71bar ( .A1(n219bar), .A2(bbar[5]), .ZN(n156bar) );
  OR2_X1 U72 ( .A1(n206), .A2(a[5]), .ZN(n157) );
  AND2_X1 U72bar ( .A1(n206bar), .A2(abar[5]), .ZN(n157bar) );
  AND2_X1 U73 ( .A1(n154), .A2(n153), .ZN(n155) );
  OR2_X1 U73bar ( .A1(n154bar), .A2(n153bar), .ZN(n155bar) );
  OR2_X1 U74 ( .A1(n195), .A2(d[5]), .ZN(n153) );
  AND2_X1 U74bar ( .A1(n195bar), .A2(dbar[5]), .ZN(n153bar) );
  OR2_X1 U75 ( .A1(n182), .A2(c[5]), .ZN(n154) );
  AND2_X1 U75bar ( .A1(n182bar), .A2(cbar[5]), .ZN(n154bar) );
  OR2_X1 U76 ( .A1(n152), .A2(n218), .ZN(y[4]) );
  AND2_X1 U76bar ( .A1(n152bar), .A2(n218bar), .ZN(ybar[4]) );
  OR2_X1 U77 ( .A1(n150), .A2(n194), .ZN(n151) );
  AND2_X1 U77bar ( .A1(n150bar), .A2(n194bar), .ZN(n151bar) );
  AND2_X1 U78 ( .A1(n194), .A2(n150), .ZN(n152) );
  OR2_X1 U78bar ( .A1(n194bar), .A2(n150bar), .ZN(n152bar) );
  AND2_X1 U79 ( .A1(n149), .A2(n148), .ZN(n150) );
  OR2_X1 U79bar ( .A1(n149bar), .A2(n148bar), .ZN(n150bar) );
  OR2_X1 U80 ( .A1(n217), .A2(b[4]), .ZN(n148) );
  AND2_X1 U80bar ( .A1(n217bar), .A2(bbar[4]), .ZN(n148bar) );
  OR2_X1 U81 ( .A1(n205), .A2(a[4]), .ZN(n149) );
  AND2_X1 U81bar ( .A1(n205bar), .A2(abar[4]), .ZN(n149bar) );
  AND2_X1 U82 ( .A1(n146), .A2(n145), .ZN(n147) );
  OR2_X1 U82bar ( .A1(n146bar), .A2(n145bar), .ZN(n147bar) );
  OR2_X1 U83 ( .A1(n193), .A2(d[4]), .ZN(n145) );
  AND2_X1 U83bar ( .A1(n193bar), .A2(dbar[4]), .ZN(n145bar) );
  OR2_X1 U84 ( .A1(n181), .A2(c[4]), .ZN(n146) );
  AND2_X1 U84bar ( .A1(n181bar), .A2(cbar[4]), .ZN(n146bar) );
  OR2_X1 U85 ( .A1(n144), .A2(n216), .ZN(y[3]) );
  AND2_X1 U85bar ( .A1(n144bar), .A2(n216bar), .ZN(ybar[3]) );
  OR2_X1 U86 ( .A1(n142), .A2(n192), .ZN(n143) );
  AND2_X1 U86bar ( .A1(n142bar), .A2(n192bar), .ZN(n143bar) );
  AND2_X1 U87 ( .A1(n192), .A2(n142), .ZN(n144) );
  OR2_X1 U87bar ( .A1(n192bar), .A2(n142bar), .ZN(n144bar) );
  AND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(n142) );
  OR2_X1 U88bar ( .A1(n141bar), .A2(n140bar), .ZN(n142bar) );
  OR2_X1 U89 ( .A1(n215), .A2(b[3]), .ZN(n140) );
  AND2_X1 U89bar ( .A1(n215bar), .A2(bbar[3]), .ZN(n140bar) );
  OR2_X1 U90 ( .A1(n204), .A2(a[3]), .ZN(n141) );
  AND2_X1 U90bar ( .A1(n204bar), .A2(abar[3]), .ZN(n141bar) );
  AND2_X1 U91 ( .A1(n138), .A2(n137), .ZN(n139) );
  OR2_X1 U91bar ( .A1(n138bar), .A2(n137bar), .ZN(n139bar) );
  OR2_X1 U92 ( .A1(n191), .A2(d[3]), .ZN(n137) );
  AND2_X1 U92bar ( .A1(n191bar), .A2(dbar[3]), .ZN(n137bar) );
  OR2_X1 U93 ( .A1(n180), .A2(c[3]), .ZN(n138) );
  AND2_X1 U93bar ( .A1(n180bar), .A2(cbar[3]), .ZN(n138bar) );
  OR2_X1 U94 ( .A1(n136), .A2(n214), .ZN(y[2]) );
  AND2_X1 U94bar ( .A1(n136bar), .A2(n214bar), .ZN(ybar[2]) );
  OR2_X1 U95 ( .A1(n134), .A2(n190), .ZN(n135) );
  AND2_X1 U95bar ( .A1(n134bar), .A2(n190bar), .ZN(n135bar) );
  AND2_X1 U96 ( .A1(n190), .A2(n134), .ZN(n136) );
  OR2_X1 U96bar ( .A1(n190bar), .A2(n134bar), .ZN(n136bar) );
  AND2_X1 U97 ( .A1(n133), .A2(n132), .ZN(n134) );
  OR2_X1 U97bar ( .A1(n133bar), .A2(n132bar), .ZN(n134bar) );
  OR2_X1 U98 ( .A1(n213), .A2(b[2]), .ZN(n132) );
  AND2_X1 U98bar ( .A1(n213bar), .A2(bbar[2]), .ZN(n132bar) );
  OR2_X1 U99 ( .A1(n203), .A2(a[2]), .ZN(n133) );
  AND2_X1 U99bar ( .A1(n203bar), .A2(abar[2]), .ZN(n133bar) );
  AND2_X1 U100 ( .A1(n130), .A2(n129), .ZN(n131) );
  OR2_X1 U100bar ( .A1(n130bar), .A2(n129bar), .ZN(n131bar) );
  OR2_X1 U101 ( .A1(n189), .A2(d[2]), .ZN(n129) );
  AND2_X1 U101bar ( .A1(n189bar), .A2(dbar[2]), .ZN(n129bar) );
  OR2_X1 U102 ( .A1(n179), .A2(c[2]), .ZN(n130) );
  AND2_X1 U102bar ( .A1(n179bar), .A2(cbar[2]), .ZN(n130bar) );
  OR2_X1 U103 ( .A1(n128), .A2(n212), .ZN(y[1]) );
  AND2_X1 U103bar ( .A1(n128bar), .A2(n212bar), .ZN(ybar[1]) );
  OR2_X1 U104 ( .A1(n126), .A2(n188), .ZN(n127) );
  AND2_X1 U104bar ( .A1(n126bar), .A2(n188bar), .ZN(n127bar) );
  AND2_X1 U105 ( .A1(n188), .A2(n126), .ZN(n128) );
  OR2_X1 U105bar ( .A1(n188bar), .A2(n126bar), .ZN(n128bar) );
  AND2_X1 U106 ( .A1(n125), .A2(n124), .ZN(n126) );
  OR2_X1 U106bar ( .A1(n125bar), .A2(n124bar), .ZN(n126bar) );
  OR2_X1 U107 ( .A1(n211), .A2(b[1]), .ZN(n124) );
  AND2_X1 U107bar ( .A1(n211bar), .A2(bbar[1]), .ZN(n124bar) );
  OR2_X1 U108 ( .A1(n202), .A2(a[1]), .ZN(n125) );
  AND2_X1 U108bar ( .A1(n202bar), .A2(abar[1]), .ZN(n125bar) );
  AND2_X1 U109 ( .A1(n122), .A2(n121), .ZN(n123) );
  OR2_X1 U109bar ( .A1(n122bar), .A2(n121bar), .ZN(n123bar) );
  OR2_X1 U110 ( .A1(n187), .A2(d[1]), .ZN(n121) );
  AND2_X1 U110bar ( .A1(n187bar), .A2(dbar[1]), .ZN(n121bar) );
  OR2_X1 U111 ( .A1(n178), .A2(c[1]), .ZN(n122) );
  AND2_X1 U111bar ( .A1(n178bar), .A2(cbar[1]), .ZN(n122bar) );
  OR2_X1 U112 ( .A1(n120), .A2(n210), .ZN(y[0]) );
  AND2_X1 U112bar ( .A1(n120bar), .A2(n210bar), .ZN(ybar[0]) );
  OR2_X1 U113 ( .A1(n118), .A2(n186), .ZN(n119) );
  AND2_X1 U113bar ( .A1(n118bar), .A2(n186bar), .ZN(n119bar) );
  AND2_X1 U114 ( .A1(n186), .A2(n118), .ZN(n120) );
  OR2_X1 U114bar ( .A1(n186bar), .A2(n118bar), .ZN(n120bar) );
  AND2_X1 U115 ( .A1(n117), .A2(n116), .ZN(n118) );
  OR2_X1 U115bar ( .A1(n117bar), .A2(n116bar), .ZN(n118bar) );
  OR2_X1 U116 ( .A1(n209), .A2(b[0]), .ZN(n116) );
  AND2_X1 U116bar ( .A1(n209bar), .A2(bbar[0]), .ZN(n116bar) );
  OR2_X1 U117 ( .A1(n201), .A2(a[0]), .ZN(n117) );
  AND2_X1 U117bar ( .A1(n201bar), .A2(abar[0]), .ZN(n117bar) );
  AND2_X1 U118 ( .A1(n114), .A2(n113), .ZN(n115) );
  OR2_X1 U118bar ( .A1(n114bar), .A2(n113bar), .ZN(n115bar) );
  OR2_X1 U119 ( .A1(n185), .A2(d[0]), .ZN(n113) );
  AND2_X1 U119bar ( .A1(n185bar), .A2(dbar[0]), .ZN(n113bar) );
  OR2_X1 U120 ( .A1(n177), .A2(c[0]), .ZN(n114) );
  AND2_X1 U120bar ( .A1(n177bar), .A2(cbar[0]), .ZN(n114bar) );
endmodule

module mixCol_3 ( in, inbar, out, outbar );

  input wire [31:0] in;
  input wire [31:0] inbar;
//input_done

  output wire [31:0] out;
  output wire [31:0] outbar;
//output_done

  wire [7:0] b0_s2;
  wire [7:0] b1_s2;
  wire [7:0] b2_s2;
  wire [7:0] b3_s2;
  wire [7:0] b0_s3;
  wire [7:0] b1_s3;
  wire [7:0] b2_s3;
  wire [7:0] b3_s3;

  wire [7:0] b0_s2bar;
  wire [7:0] b1_s2bar;
  wire [7:0] b2_s2bar;
  wire [7:0] b3_s2bar;
  wire [7:0] b0_s3bar;
  wire [7:0] b1_s3bar;
  wire [7:0] b2_s3bar;
  wire [7:0] b3_s3bar;
//wire_done

 //assign_done

  scale2_12 b0_scale2 ( .in(in[31:24]), .inbar(inbar[31:24]), .out(b0_s2), .outbar(b0_s2bar) );
  scale2_11 b1_scale2 ( .in(in[23:16]), .inbar(inbar[23:16]), .out(b1_s2), .outbar(b1_s2bar) );
  scale2_10 b2_scale2 ( .in(in[15:8]), .inbar(inbar[15:8]), .out(b2_s2), .outbar(b2_s2bar) );
  scale2_9 b3_scale2 ( .in(in[7:0]), .inbar(inbar[7:0]), .out(b3_s2), .outbar(b3_s2bar) );

  byteXor_13 b0_scale3 ( .a(in[31:24]), .abar(inbar[31:24]), .b(b0_s2), .bbar(b0_s2bar), .y(b0_s3), .ybar(b0_s3bar) );
  byteXor_12 b1_scale3 ( .a(in[23:16]), .abar(inbar[23:16]), .b(b1_s2), .bbar(b1_s2bar), .y(b1_s3), .ybar(b1_s3bar) );
  byteXor_11 b2_scale3 ( .a(in[15:8]), .abar(inbar[15:8]), .b(b2_s2), .bbar(b2_s2bar), .y(b2_s3), .ybar(b2_s3bar) );
  byteXor_10 b3_scale3 ( .a(in[7:0]), .abar(inbar[7:0]), .b(b3_s2), .bbar(b3_s2bar), .y(b3_s3), .ybar(b3_s3bar) );

  byteXor4_12 out0 ( .a(b0_s2), .abar(b0_s2bar), .b(b1_s3), .bbar(b1_s3bar), .c(in[15:8]), .cbar(inbar[15:8]),
       .d(in[7:0]), .dbar(inbar[7:0]), .y(out[31:24]), .ybar(outbar[31:24]) );
  byteXor4_11 out1 ( .a(in[31:24]), .abar(inbar[31:24]), .b(b1_s2), .bbar(b1_s2bar), .c(b2_s3), .cbar(b2_s3bar),
       .d(in[7:0]), .dbar(inbar[7:0]), .y(out[23:16]), .ybar(outbar[23:16]) );
  byteXor4_10 out2 ( .a(in[31:24]), .abar(inbar[31:24]), .b(in[23:16]), .bbar(inbar[23:16]), .c(b2_s2), .cbar(b2_s2bar),
       .d(b3_s3), .dbar(b3_s3bar), .y(out[15:8]), .ybar(outbar[15:8]) );
  byteXor4_9 out3 ( .a(b0_s3), .abar(b0_s3bar), .b(in[23:16]), .bbar(inbar[23:16]), .c(in[15:8]), .cbar(inbar[15:8]),
       .d(b3_s2), .dbar(b3_s2bar), .y(out[7:0]), .ybar(outbar[7:0]) );
endmodule

module mixCol_Precharge ( in, inbar, out, outbar );

  input wire [127:0] in;
  input wire [127:0] inbar;
//input_done

  output [127:0] out;
  output [127:0] outbar;
//output_done

//wire_done

 //assign_done

  mixCol_0 m0( .in(in[127:96]) .inbar(inbar[127:96]), .out(out[127:96]), .outbar(outbar[127:96]) );
  mixCol_3 m1( .in(in[95:64]) .inbar(inbar[95:64]), .out(out[95:64]), .outbar(outbar[95:64]) );
  mixCol_2 m2( .in(in[63:32]) .inbar(inbar[63:32]), .out(out[63:32]), .outbar(outbar[63:32]) );
  mixCol_1 m3( .in(in[31:0]) .inbar(inbar[31:0]), .out(out[31:0]), .outbar(outbar[31:0]) );
endmodule

//done
