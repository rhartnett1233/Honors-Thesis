module AND2_X1( A1, A2, ZN );

  input wire A1;
  input wire A2;
//input_done

  output wire ZN;
//output_done

//wire_done

  assign ZN = A1 & A2;
//assign_done

 endmodule

module OR2_X1( A1, A2, ZN );

  input wire A1;
  input wire A2;
//input_done

  output wire ZN;
//output_done

//wire_done

  assign ZN = A1 | A2;
//assign_done

 endmodule

module INV_X1( A, ZN );

  input wire A;
//input_done

  output wire ZN;
//output_done

//wire_done

  assign ZN = ~A;
//assign_done

 endmodule

module scale2_0 ( in, out );

  input wire [7:0] in;
  wire [7:0] inbar;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
//input_done

  output wire [7:0] out;
  wire [7:0] outbar;
//output_done

  wire in_0;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_1;
  wire in_7;
  wire n1;
  wire n2;
  wire n3;
  wire n4;
  wire n5;
  wire n6;
  wire n7;
  wire n8;
  wire n9;
  wire n10;
  wire in_0bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_1bar;
  wire in_7bar;
  wire n1bar;
  wire n2bar;
  wire n3bar;
  wire n4bar;
  wire n5bar;
  wire n6bar;
  wire n7bar;
  wire n8bar;
  wire n9bar;
  wire n10bar;
//wire_done

  assign in_0 = in[0];
  assign out[7] = in_6;
  assign in_6  = in[6];
  assign out[6] = in_5;
  assign in_5  = in[5];
  assign out[5] = in_4;
  assign in_4  = in[4];
  assign out[2] = in_1;
  assign in_1  = in[1];
  assign out[0] = in_7;
  assign in_7  = in[7];
  assign in_0bar = inbar[0];
  assign outbar[7] = in_6bar;
  assign in_6bar = inbar[6];
  assign outbar[6] = in_5bar;
  assign in_5bar = inbar[5];
  assign outbar[5] = in_4bar;
  assign in_4bar = inbar[4];
  assign outbar[2] = in_1bar;
  assign in_1bar = inbar[1];
  assign outbar[0] = in_7bar;
  assign in_7bar = inbar[7];
//assign_done

  assign n1bar = in_7;
  assign n1 = in_7bar;
  assign n2bar = in[3];
  assign n2 = inbar[3];
  assign n3bar = in[2];
  assign n3 = inbar[2];
  assign n4bar = in_0;
  assign n4 = in_0bar;
  OR2_X1 U5 ( .A1(n5), .A2(n6), .ZN(out[4]) );
  AND2_X1 U5bar ( .A1(n5bar), .A2(n6bar), .ZN(outbar[4]) );
  AND2_X1 U6 ( .A1(in[3]), .A2(n1), .ZN(n6) );
  OR2_X1 U6bar ( .A1(inbar[3]), .A2(n1bar), .ZN(n6bar) );
  AND2_X1 U7 ( .A1(in_7), .A2(n2), .ZN(n5) );
  OR2_X1 U7bar ( .A1(in_7bar), .A2(n2bar), .ZN(n5bar) );
  OR2_X1 U8 ( .A1(n7), .A2(n8), .ZN(out[3]) );
  AND2_X1 U8bar ( .A1(n7bar), .A2(n8bar), .ZN(outbar[3]) );
  AND2_X1 U9 ( .A1(in[2]), .A2(n1), .ZN(n8) );
  OR2_X1 U9bar ( .A1(inbar[2]), .A2(n1bar), .ZN(n8bar) );
  AND2_X1 U10 ( .A1(in_7), .A2(n3), .ZN(n7) );
  OR2_X1 U10bar ( .A1(in_7bar), .A2(n3bar), .ZN(n7bar) );
  OR2_X1 U11 ( .A1(n9), .A2(n10), .ZN(out[1]) );
  AND2_X1 U11bar ( .A1(n9bar), .A2(n10bar), .ZN(outbar[1]) );
  AND2_X1 U12 ( .A1(in_0), .A2(n1), .ZN(n10) );
  OR2_X1 U12bar ( .A1(in_0bar), .A2(n1bar), .ZN(n10bar) );
  AND2_X1 U13 ( .A1(in_7), .A2(n4), .ZN(n9) );
  OR2_X1 U13bar ( .A1(in_7bar), .A2(n4bar), .ZN(n9bar) );
endmodule

module byteXor_0 ( a, b, y );

  input wire [7:0] a;
  input wire [7:0] b;
  wire [7:0] abar;
  wire [7:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
//input_done

  output wire [7:0] y;
  wire [7:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n3;
  wire n4;
  wire n5;
  wire n6;
  wire n7;
  wire n8;
  wire n9;
  wire n10;
  wire n11;
  wire n12;
  wire n13;
  wire n14;
  wire n15;
  wire n16;
  wire n17;
  wire n18;
  wire n19;
  wire n20;
  wire n21;
  wire n22;
  wire n23;
  wire n24;
  wire n25;
  wire n26;
  wire n27;
  wire n28;
  wire n29;
  wire n30;
  wire n31;
  wire n32;
  wire n1bar;
  wire n2bar;
  wire n3bar;
  wire n4bar;
  wire n5bar;
  wire n6bar;
  wire n7bar;
  wire n8bar;
  wire n9bar;
  wire n10bar;
  wire n11bar;
  wire n12bar;
  wire n13bar;
  wire n14bar;
  wire n15bar;
  wire n16bar;
  wire n17bar;
  wire n18bar;
  wire n19bar;
  wire n20bar;
  wire n21bar;
  wire n22bar;
  wire n23bar;
  wire n24bar;
  wire n25bar;
  wire n26bar;
  wire n27bar;
  wire n28bar;
  wire n29bar;
  wire n30bar;
  wire n31bar;
  wire n32bar;
//wire_done

 //assign_done

  assign n1bar = n18;
  assign n1 = n18bar;
  assign n2bar = a[7];
  assign n2 = abar[7];
  assign n3bar = n20;
  assign n3 = n20bar;
  assign n4bar = a[6];
  assign n4 = abar[6];
  assign n5bar = n22;
  assign n5 = n22bar;
  assign n6bar = a[5];
  assign n6 = abar[5];
  assign n7bar = n24;
  assign n7 = n24bar;
  assign n8bar = a[4];
  assign n8 = abar[4];
  assign n9bar = n26;
  assign n9 = n26bar;
  assign n10bar = a[3];
  assign n10 = abar[3];
  assign n11bar = n28;
  assign n11 = n28bar;
  assign n12bar = a[2];
  assign n12 = abar[2];
  assign n13bar = n30;
  assign n13 = n30bar;
  assign n14bar = a[1];
  assign n14 = abar[1];
  assign n15bar = n32;
  assign n15 = n32bar;
  assign n16bar = a[0];
  assign n16 = abar[0];
  OR2_X1 U17 ( .A1(n17), .A2(n1), .ZN(y[7]) );
  AND2_X1 U17bar ( .A1(n17bar), .A2(n1bar), .ZN(ybar[7]) );
  OR2_X1 U18 ( .A1(n2), .A2(b[7]), .ZN(n18) );
  AND2_X1 U18bar ( .A1(n2bar), .A2(bbar[7]), .ZN(n18bar) );
  AND2_X1 U19 ( .A1(b[7]), .A2(n2), .ZN(n17) );
  OR2_X1 U19bar ( .A1(bbar[7]), .A2(n2bar), .ZN(n17bar) );
  OR2_X1 U20 ( .A1(n19), .A2(n3), .ZN(y[6]) );
  AND2_X1 U20bar ( .A1(n19bar), .A2(n3bar), .ZN(ybar[6]) );
  OR2_X1 U21 ( .A1(n4), .A2(b[6]), .ZN(n20) );
  AND2_X1 U21bar ( .A1(n4bar), .A2(bbar[6]), .ZN(n20bar) );
  AND2_X1 U22 ( .A1(b[6]), .A2(n4), .ZN(n19) );
  OR2_X1 U22bar ( .A1(bbar[6]), .A2(n4bar), .ZN(n19bar) );
  OR2_X1 U23 ( .A1(n21), .A2(n5), .ZN(y[5]) );
  AND2_X1 U23bar ( .A1(n21bar), .A2(n5bar), .ZN(ybar[5]) );
  OR2_X1 U24 ( .A1(n6), .A2(b[5]), .ZN(n22) );
  AND2_X1 U24bar ( .A1(n6bar), .A2(bbar[5]), .ZN(n22bar) );
  AND2_X1 U25 ( .A1(b[5]), .A2(n6), .ZN(n21) );
  OR2_X1 U25bar ( .A1(bbar[5]), .A2(n6bar), .ZN(n21bar) );
  OR2_X1 U26 ( .A1(n23), .A2(n7), .ZN(y[4]) );
  AND2_X1 U26bar ( .A1(n23bar), .A2(n7bar), .ZN(ybar[4]) );
  OR2_X1 U27 ( .A1(n8), .A2(b[4]), .ZN(n24) );
  AND2_X1 U27bar ( .A1(n8bar), .A2(bbar[4]), .ZN(n24bar) );
  AND2_X1 U28 ( .A1(b[4]), .A2(n8), .ZN(n23) );
  OR2_X1 U28bar ( .A1(bbar[4]), .A2(n8bar), .ZN(n23bar) );
  OR2_X1 U29 ( .A1(n25), .A2(n9), .ZN(y[3]) );
  AND2_X1 U29bar ( .A1(n25bar), .A2(n9bar), .ZN(ybar[3]) );
  OR2_X1 U30 ( .A1(n10), .A2(b[3]), .ZN(n26) );
  AND2_X1 U30bar ( .A1(n10bar), .A2(bbar[3]), .ZN(n26bar) );
  AND2_X1 U31 ( .A1(b[3]), .A2(n10), .ZN(n25) );
  OR2_X1 U31bar ( .A1(bbar[3]), .A2(n10bar), .ZN(n25bar) );
  OR2_X1 U32 ( .A1(n27), .A2(n11), .ZN(y[2]) );
  AND2_X1 U32bar ( .A1(n27bar), .A2(n11bar), .ZN(ybar[2]) );
  OR2_X1 U33 ( .A1(n12), .A2(b[2]), .ZN(n28) );
  AND2_X1 U33bar ( .A1(n12bar), .A2(bbar[2]), .ZN(n28bar) );
  AND2_X1 U34 ( .A1(b[2]), .A2(n12), .ZN(n27) );
  OR2_X1 U34bar ( .A1(bbar[2]), .A2(n12bar), .ZN(n27bar) );
  OR2_X1 U35 ( .A1(n29), .A2(n13), .ZN(y[1]) );
  AND2_X1 U35bar ( .A1(n29bar), .A2(n13bar), .ZN(ybar[1]) );
  OR2_X1 U36 ( .A1(n14), .A2(b[1]), .ZN(n30) );
  AND2_X1 U36bar ( .A1(n14bar), .A2(bbar[1]), .ZN(n30bar) );
  AND2_X1 U37 ( .A1(b[1]), .A2(n14), .ZN(n29) );
  OR2_X1 U37bar ( .A1(bbar[1]), .A2(n14bar), .ZN(n29bar) );
  OR2_X1 U38 ( .A1(n31), .A2(n15), .ZN(y[0]) );
  AND2_X1 U38bar ( .A1(n31bar), .A2(n15bar), .ZN(ybar[0]) );
  OR2_X1 U39 ( .A1(n16), .A2(b[0]), .ZN(n32) );
  AND2_X1 U39bar ( .A1(n16bar), .A2(bbar[0]), .ZN(n32bar) );
  AND2_X1 U40 ( .A1(b[0]), .A2(n16), .ZN(n31) );
  OR2_X1 U40bar ( .A1(bbar[0]), .A2(n16bar), .ZN(n31bar) );
endmodule

module byteXor4_0 ( a, b, c, d, y );

  input wire [7:0] a;
  input wire [7:0] b;
  input wire [7:0] c;
  input wire [7:0] d;
  wire [7:0] abar;
  wire [7:0] bbar;
  wire [7:0] cbar;
  wire [7:0] dbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign cbar[0] = ~c[0];
  assign cbar[1] = ~c[1];
  assign cbar[2] = ~c[2];
  assign cbar[3] = ~c[3];
  assign cbar[4] = ~c[4];
  assign cbar[5] = ~c[5];
  assign cbar[6] = ~c[6];
  assign cbar[7] = ~c[7];
  assign dbar[0] = ~d[0];
  assign dbar[1] = ~d[1];
  assign dbar[2] = ~d[2];
  assign dbar[3] = ~d[3];
  assign dbar[4] = ~d[4];
  assign dbar[5] = ~d[5];
  assign dbar[6] = ~d[6];
  assign dbar[7] = ~d[7];
//input_done

  output wire [7:0] y;
  wire [7:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n3;
  wire n4;
  wire n5;
  wire n6;
  wire n7;
  wire n8;
  wire n9;
  wire n10;
  wire n11;
  wire n12;
  wire n13;
  wire n14;
  wire n15;
  wire n16;
  wire n17;
  wire n18;
  wire n19;
  wire n20;
  wire n21;
  wire n22;
  wire n23;
  wire n24;
  wire n25;
  wire n26;
  wire n27;
  wire n28;
  wire n29;
  wire n30;
  wire n31;
  wire n32;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n1bar;
  wire n2bar;
  wire n3bar;
  wire n4bar;
  wire n5bar;
  wire n6bar;
  wire n7bar;
  wire n8bar;
  wire n9bar;
  wire n10bar;
  wire n11bar;
  wire n12bar;
  wire n13bar;
  wire n14bar;
  wire n15bar;
  wire n16bar;
  wire n17bar;
  wire n18bar;
  wire n19bar;
  wire n20bar;
  wire n21bar;
  wire n22bar;
  wire n23bar;
  wire n24bar;
  wire n25bar;
  wire n26bar;
  wire n27bar;
  wire n28bar;
  wire n29bar;
  wire n30bar;
  wire n31bar;
  wire n32bar;
  wire n33bar;
  wire n34bar;
  wire n35bar;
  wire n36bar;
  wire n37bar;
  wire n38bar;
  wire n39bar;
  wire n40bar;
  wire n41bar;
  wire n42bar;
  wire n43bar;
  wire n44bar;
  wire n45bar;
  wire n46bar;
  wire n47bar;
  wire n48bar;
  wire n49bar;
  wire n50bar;
  wire n51bar;
  wire n52bar;
  wire n53bar;
  wire n54bar;
  wire n55bar;
  wire n56bar;
  wire n57bar;
  wire n58bar;
  wire n59bar;
  wire n60bar;
  wire n61bar;
  wire n62bar;
  wire n63bar;
  wire n64bar;
  wire n65bar;
  wire n66bar;
  wire n67bar;
  wire n68bar;
  wire n69bar;
  wire n70bar;
  wire n71bar;
  wire n72bar;
  wire n73bar;
  wire n74bar;
  wire n75bar;
  wire n76bar;
  wire n77bar;
  wire n78bar;
  wire n79bar;
  wire n80bar;
  wire n81bar;
  wire n82bar;
  wire n83bar;
  wire n84bar;
  wire n85bar;
  wire n86bar;
  wire n87bar;
  wire n88bar;
  wire n89bar;
  wire n90bar;
  wire n91bar;
  wire n92bar;
  wire n93bar;
  wire n94bar;
  wire n95bar;
  wire n96bar;
  wire n97bar;
  wire n98bar;
  wire n99bar;
  wire n100bar;
  wire n101bar;
  wire n102bar;
  wire n103bar;
  wire n104bar;
  wire n105bar;
  wire n106bar;
  wire n107bar;
  wire n108bar;
  wire n109bar;
  wire n110bar;
  wire n111bar;
  wire n112bar;
//wire_done

 //assign_done

  assign n1bar = n50;
  assign n1 = n50bar;
  assign n2bar = a[7];
  assign n2 = abar[7];
  assign n3bar = n58;
  assign n3 = n58bar;
  assign n4bar = a[6];
  assign n4 = abar[6];
  assign n5bar = n66;
  assign n5 = n66bar;
  assign n6bar = a[5];
  assign n6 = abar[5];
  assign n7bar = n74;
  assign n7 = n74bar;
  assign n8bar = a[4];
  assign n8 = abar[4];
  assign n9bar = n82;
  assign n9 = n82bar;
  assign n10bar = a[3];
  assign n10 = abar[3];
  assign n11bar = n90;
  assign n11 = n90bar;
  assign n12bar = a[2];
  assign n12 = abar[2];
  assign n13bar = n98;
  assign n13 = n98bar;
  assign n14bar = a[1];
  assign n14 = abar[1];
  assign n15bar = n106;
  assign n15 = n106bar;
  assign n16bar = a[0];
  assign n16 = abar[0];
  assign n17bar = b[7];
  assign n17 = bbar[7];
  assign n18bar = b[6];
  assign n18 = bbar[6];
  assign n19bar = b[5];
  assign n19 = bbar[5];
  assign n20bar = b[4];
  assign n20 = bbar[4];
  assign n21bar = b[3];
  assign n21 = bbar[3];
  assign n22bar = b[2];
  assign n22 = bbar[2];
  assign n23bar = b[1];
  assign n23 = bbar[1];
  assign n24bar = b[0];
  assign n24 = bbar[0];
  assign n25bar = n54;
  assign n25 = n54bar;
  assign n26bar = c[7];
  assign n26 = cbar[7];
  assign n27bar = n62;
  assign n27 = n62bar;
  assign n28bar = c[6];
  assign n28 = cbar[6];
  assign n29bar = n70;
  assign n29 = n70bar;
  assign n30bar = c[5];
  assign n30 = cbar[5];
  assign n31bar = n78;
  assign n31 = n78bar;
  assign n32bar = c[4];
  assign n32 = cbar[4];
  assign n33bar = n86;
  assign n33 = n86bar;
  assign n34bar = c[3];
  assign n34 = cbar[3];
  assign n35bar = n94;
  assign n35 = n94bar;
  assign n36bar = c[2];
  assign n36 = cbar[2];
  assign n37bar = n102;
  assign n37 = n102bar;
  assign n38bar = c[1];
  assign n38 = cbar[1];
  assign n39bar = n110;
  assign n39 = n110bar;
  assign n40bar = c[0];
  assign n40 = cbar[0];
  assign n41bar = d[7];
  assign n41 = dbar[7];
  assign n42bar = d[6];
  assign n42 = dbar[6];
  assign n43bar = d[5];
  assign n43 = dbar[5];
  assign n44bar = d[4];
  assign n44 = dbar[4];
  assign n45bar = d[3];
  assign n45 = dbar[3];
  assign n46bar = d[2];
  assign n46 = dbar[2];
  assign n47bar = d[1];
  assign n47 = dbar[1];
  assign n48bar = d[0];
  assign n48 = dbar[0];
  OR2_X1 U49 ( .A1(n49), .A2(n1), .ZN(y[7]) );
  AND2_X1 U49bar ( .A1(n49bar), .A2(n1bar), .ZN(ybar[7]) );
  OR2_X1 U50 ( .A1(n51), .A2(n25), .ZN(n50) );
  AND2_X1 U50bar ( .A1(n51bar), .A2(n25bar), .ZN(n50bar) );
  AND2_X1 U51 ( .A1(n25), .A2(n51), .ZN(n49) );
  OR2_X1 U51bar ( .A1(n25bar), .A2(n51bar), .ZN(n49bar) );
  AND2_X1 U52 ( .A1(n52), .A2(n53), .ZN(n51) );
  OR2_X1 U52bar ( .A1(n52bar), .A2(n53bar), .ZN(n51bar) );
  OR2_X1 U53 ( .A1(n2), .A2(b[7]), .ZN(n53) );
  AND2_X1 U53bar ( .A1(n2bar), .A2(bbar[7]), .ZN(n53bar) );
  OR2_X1 U54 ( .A1(n17), .A2(a[7]), .ZN(n52) );
  AND2_X1 U54bar ( .A1(n17bar), .A2(abar[7]), .ZN(n52bar) );
  AND2_X1 U55 ( .A1(n55), .A2(n56), .ZN(n54) );
  OR2_X1 U55bar ( .A1(n55bar), .A2(n56bar), .ZN(n54bar) );
  OR2_X1 U56 ( .A1(n26), .A2(d[7]), .ZN(n56) );
  AND2_X1 U56bar ( .A1(n26bar), .A2(dbar[7]), .ZN(n56bar) );
  OR2_X1 U57 ( .A1(n41), .A2(c[7]), .ZN(n55) );
  AND2_X1 U57bar ( .A1(n41bar), .A2(cbar[7]), .ZN(n55bar) );
  OR2_X1 U58 ( .A1(n57), .A2(n3), .ZN(y[6]) );
  AND2_X1 U58bar ( .A1(n57bar), .A2(n3bar), .ZN(ybar[6]) );
  OR2_X1 U59 ( .A1(n59), .A2(n27), .ZN(n58) );
  AND2_X1 U59bar ( .A1(n59bar), .A2(n27bar), .ZN(n58bar) );
  AND2_X1 U60 ( .A1(n27), .A2(n59), .ZN(n57) );
  OR2_X1 U60bar ( .A1(n27bar), .A2(n59bar), .ZN(n57bar) );
  AND2_X1 U61 ( .A1(n60), .A2(n61), .ZN(n59) );
  OR2_X1 U61bar ( .A1(n60bar), .A2(n61bar), .ZN(n59bar) );
  OR2_X1 U62 ( .A1(n4), .A2(b[6]), .ZN(n61) );
  AND2_X1 U62bar ( .A1(n4bar), .A2(bbar[6]), .ZN(n61bar) );
  OR2_X1 U63 ( .A1(n18), .A2(a[6]), .ZN(n60) );
  AND2_X1 U63bar ( .A1(n18bar), .A2(abar[6]), .ZN(n60bar) );
  AND2_X1 U64 ( .A1(n63), .A2(n64), .ZN(n62) );
  OR2_X1 U64bar ( .A1(n63bar), .A2(n64bar), .ZN(n62bar) );
  OR2_X1 U65 ( .A1(n28), .A2(d[6]), .ZN(n64) );
  AND2_X1 U65bar ( .A1(n28bar), .A2(dbar[6]), .ZN(n64bar) );
  OR2_X1 U66 ( .A1(n42), .A2(c[6]), .ZN(n63) );
  AND2_X1 U66bar ( .A1(n42bar), .A2(cbar[6]), .ZN(n63bar) );
  OR2_X1 U67 ( .A1(n65), .A2(n5), .ZN(y[5]) );
  AND2_X1 U67bar ( .A1(n65bar), .A2(n5bar), .ZN(ybar[5]) );
  OR2_X1 U68 ( .A1(n67), .A2(n29), .ZN(n66) );
  AND2_X1 U68bar ( .A1(n67bar), .A2(n29bar), .ZN(n66bar) );
  AND2_X1 U69 ( .A1(n29), .A2(n67), .ZN(n65) );
  OR2_X1 U69bar ( .A1(n29bar), .A2(n67bar), .ZN(n65bar) );
  AND2_X1 U70 ( .A1(n68), .A2(n69), .ZN(n67) );
  OR2_X1 U70bar ( .A1(n68bar), .A2(n69bar), .ZN(n67bar) );
  OR2_X1 U71 ( .A1(n6), .A2(b[5]), .ZN(n69) );
  AND2_X1 U71bar ( .A1(n6bar), .A2(bbar[5]), .ZN(n69bar) );
  OR2_X1 U72 ( .A1(n19), .A2(a[5]), .ZN(n68) );
  AND2_X1 U72bar ( .A1(n19bar), .A2(abar[5]), .ZN(n68bar) );
  AND2_X1 U73 ( .A1(n71), .A2(n72), .ZN(n70) );
  OR2_X1 U73bar ( .A1(n71bar), .A2(n72bar), .ZN(n70bar) );
  OR2_X1 U74 ( .A1(n30), .A2(d[5]), .ZN(n72) );
  AND2_X1 U74bar ( .A1(n30bar), .A2(dbar[5]), .ZN(n72bar) );
  OR2_X1 U75 ( .A1(n43), .A2(c[5]), .ZN(n71) );
  AND2_X1 U75bar ( .A1(n43bar), .A2(cbar[5]), .ZN(n71bar) );
  OR2_X1 U76 ( .A1(n73), .A2(n7), .ZN(y[4]) );
  AND2_X1 U76bar ( .A1(n73bar), .A2(n7bar), .ZN(ybar[4]) );
  OR2_X1 U77 ( .A1(n75), .A2(n31), .ZN(n74) );
  AND2_X1 U77bar ( .A1(n75bar), .A2(n31bar), .ZN(n74bar) );
  AND2_X1 U78 ( .A1(n31), .A2(n75), .ZN(n73) );
  OR2_X1 U78bar ( .A1(n31bar), .A2(n75bar), .ZN(n73bar) );
  AND2_X1 U79 ( .A1(n76), .A2(n77), .ZN(n75) );
  OR2_X1 U79bar ( .A1(n76bar), .A2(n77bar), .ZN(n75bar) );
  OR2_X1 U80 ( .A1(n8), .A2(b[4]), .ZN(n77) );
  AND2_X1 U80bar ( .A1(n8bar), .A2(bbar[4]), .ZN(n77bar) );
  OR2_X1 U81 ( .A1(n20), .A2(a[4]), .ZN(n76) );
  AND2_X1 U81bar ( .A1(n20bar), .A2(abar[4]), .ZN(n76bar) );
  AND2_X1 U82 ( .A1(n79), .A2(n80), .ZN(n78) );
  OR2_X1 U82bar ( .A1(n79bar), .A2(n80bar), .ZN(n78bar) );
  OR2_X1 U83 ( .A1(n32), .A2(d[4]), .ZN(n80) );
  AND2_X1 U83bar ( .A1(n32bar), .A2(dbar[4]), .ZN(n80bar) );
  OR2_X1 U84 ( .A1(n44), .A2(c[4]), .ZN(n79) );
  AND2_X1 U84bar ( .A1(n44bar), .A2(cbar[4]), .ZN(n79bar) );
  OR2_X1 U85 ( .A1(n81), .A2(n9), .ZN(y[3]) );
  AND2_X1 U85bar ( .A1(n81bar), .A2(n9bar), .ZN(ybar[3]) );
  OR2_X1 U86 ( .A1(n83), .A2(n33), .ZN(n82) );
  AND2_X1 U86bar ( .A1(n83bar), .A2(n33bar), .ZN(n82bar) );
  AND2_X1 U87 ( .A1(n33), .A2(n83), .ZN(n81) );
  OR2_X1 U87bar ( .A1(n33bar), .A2(n83bar), .ZN(n81bar) );
  AND2_X1 U88 ( .A1(n84), .A2(n85), .ZN(n83) );
  OR2_X1 U88bar ( .A1(n84bar), .A2(n85bar), .ZN(n83bar) );
  OR2_X1 U89 ( .A1(n10), .A2(b[3]), .ZN(n85) );
  AND2_X1 U89bar ( .A1(n10bar), .A2(bbar[3]), .ZN(n85bar) );
  OR2_X1 U90 ( .A1(n21), .A2(a[3]), .ZN(n84) );
  AND2_X1 U90bar ( .A1(n21bar), .A2(abar[3]), .ZN(n84bar) );
  AND2_X1 U91 ( .A1(n87), .A2(n88), .ZN(n86) );
  OR2_X1 U91bar ( .A1(n87bar), .A2(n88bar), .ZN(n86bar) );
  OR2_X1 U92 ( .A1(n34), .A2(d[3]), .ZN(n88) );
  AND2_X1 U92bar ( .A1(n34bar), .A2(dbar[3]), .ZN(n88bar) );
  OR2_X1 U93 ( .A1(n45), .A2(c[3]), .ZN(n87) );
  AND2_X1 U93bar ( .A1(n45bar), .A2(cbar[3]), .ZN(n87bar) );
  OR2_X1 U94 ( .A1(n89), .A2(n11), .ZN(y[2]) );
  AND2_X1 U94bar ( .A1(n89bar), .A2(n11bar), .ZN(ybar[2]) );
  OR2_X1 U95 ( .A1(n91), .A2(n35), .ZN(n90) );
  AND2_X1 U95bar ( .A1(n91bar), .A2(n35bar), .ZN(n90bar) );
  AND2_X1 U96 ( .A1(n35), .A2(n91), .ZN(n89) );
  OR2_X1 U96bar ( .A1(n35bar), .A2(n91bar), .ZN(n89bar) );
  AND2_X1 U97 ( .A1(n92), .A2(n93), .ZN(n91) );
  OR2_X1 U97bar ( .A1(n92bar), .A2(n93bar), .ZN(n91bar) );
  OR2_X1 U98 ( .A1(n12), .A2(b[2]), .ZN(n93) );
  AND2_X1 U98bar ( .A1(n12bar), .A2(bbar[2]), .ZN(n93bar) );
  OR2_X1 U99 ( .A1(n22), .A2(a[2]), .ZN(n92) );
  AND2_X1 U99bar ( .A1(n22bar), .A2(abar[2]), .ZN(n92bar) );
  AND2_X1 U100 ( .A1(n95), .A2(n96), .ZN(n94) );
  OR2_X1 U100bar ( .A1(n95bar), .A2(n96bar), .ZN(n94bar) );
  OR2_X1 U101 ( .A1(n36), .A2(d[2]), .ZN(n96) );
  AND2_X1 U101bar ( .A1(n36bar), .A2(dbar[2]), .ZN(n96bar) );
  OR2_X1 U102 ( .A1(n46), .A2(c[2]), .ZN(n95) );
  AND2_X1 U102bar ( .A1(n46bar), .A2(cbar[2]), .ZN(n95bar) );
  OR2_X1 U103 ( .A1(n97), .A2(n13), .ZN(y[1]) );
  AND2_X1 U103bar ( .A1(n97bar), .A2(n13bar), .ZN(ybar[1]) );
  OR2_X1 U104 ( .A1(n99), .A2(n37), .ZN(n98) );
  AND2_X1 U104bar ( .A1(n99bar), .A2(n37bar), .ZN(n98bar) );
  AND2_X1 U105 ( .A1(n37), .A2(n99), .ZN(n97) );
  OR2_X1 U105bar ( .A1(n37bar), .A2(n99bar), .ZN(n97bar) );
  AND2_X1 U106 ( .A1(n100), .A2(n101), .ZN(n99) );
  OR2_X1 U106bar ( .A1(n100bar), .A2(n101bar), .ZN(n99bar) );
  OR2_X1 U107 ( .A1(n14), .A2(b[1]), .ZN(n101) );
  AND2_X1 U107bar ( .A1(n14bar), .A2(bbar[1]), .ZN(n101bar) );
  OR2_X1 U108 ( .A1(n23), .A2(a[1]), .ZN(n100) );
  AND2_X1 U108bar ( .A1(n23bar), .A2(abar[1]), .ZN(n100bar) );
  AND2_X1 U109 ( .A1(n103), .A2(n104), .ZN(n102) );
  OR2_X1 U109bar ( .A1(n103bar), .A2(n104bar), .ZN(n102bar) );
  OR2_X1 U110 ( .A1(n38), .A2(d[1]), .ZN(n104) );
  AND2_X1 U110bar ( .A1(n38bar), .A2(dbar[1]), .ZN(n104bar) );
  OR2_X1 U111 ( .A1(n47), .A2(c[1]), .ZN(n103) );
  AND2_X1 U111bar ( .A1(n47bar), .A2(cbar[1]), .ZN(n103bar) );
  OR2_X1 U112 ( .A1(n105), .A2(n15), .ZN(y[0]) );
  AND2_X1 U112bar ( .A1(n105bar), .A2(n15bar), .ZN(ybar[0]) );
  OR2_X1 U113 ( .A1(n107), .A2(n39), .ZN(n106) );
  AND2_X1 U113bar ( .A1(n107bar), .A2(n39bar), .ZN(n106bar) );
  AND2_X1 U114 ( .A1(n39), .A2(n107), .ZN(n105) );
  OR2_X1 U114bar ( .A1(n39bar), .A2(n107bar), .ZN(n105bar) );
  AND2_X1 U115 ( .A1(n108), .A2(n109), .ZN(n107) );
  OR2_X1 U115bar ( .A1(n108bar), .A2(n109bar), .ZN(n107bar) );
  OR2_X1 U116 ( .A1(n16), .A2(b[0]), .ZN(n109) );
  AND2_X1 U116bar ( .A1(n16bar), .A2(bbar[0]), .ZN(n109bar) );
  OR2_X1 U117 ( .A1(n24), .A2(a[0]), .ZN(n108) );
  AND2_X1 U117bar ( .A1(n24bar), .A2(abar[0]), .ZN(n108bar) );
  AND2_X1 U118 ( .A1(n111), .A2(n112), .ZN(n110) );
  OR2_X1 U118bar ( .A1(n111bar), .A2(n112bar), .ZN(n110bar) );
  OR2_X1 U119 ( .A1(n40), .A2(d[0]), .ZN(n112) );
  AND2_X1 U119bar ( .A1(n40bar), .A2(dbar[0]), .ZN(n112bar) );
  OR2_X1 U120 ( .A1(n48), .A2(c[0]), .ZN(n111) );
  AND2_X1 U120bar ( .A1(n48bar), .A2(cbar[0]), .ZN(n111bar) );
endmodule

module scale2_13 ( in, out );

  input wire [7:0] in;
  wire [7:0] inbar;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
//input_done

  output wire [7:0] out;
  wire [7:0] outbar;
//output_done

  wire in_0;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_1;
  wire in_7;
  wire n11;
  wire n12;
  wire n13;
  wire n14;
  wire n15;
  wire n16;
  wire n17;
  wire n18;
  wire n19;
  wire n20;
  wire in_0bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_1bar;
  wire in_7bar;
  wire n11bar;
  wire n12bar;
  wire n13bar;
  wire n14bar;
  wire n15bar;
  wire n16bar;
  wire n17bar;
  wire n18bar;
  wire n19bar;
  wire n20bar;
//wire_done

  assign in_0 = in[0];
  assign out[7] = in_6;
  assign in_6  = in[6];
  assign out[6] = in_5;
  assign in_5  = in[5];
  assign out[5] = in_4;
  assign in_4  = in[4];
  assign out[2] = in_1;
  assign in_1  = in[1];
  assign out[0] = in_7;
  assign in_7  = in[7];
  assign in_0bar = inbar[0];
  assign outbar[7] = in_6bar;
  assign in_6bar = inbar[6];
  assign outbar[6] = in_5bar;
  assign in_5bar = inbar[5];
  assign outbar[5] = in_4bar;
  assign in_4bar = inbar[4];
  assign outbar[2] = in_1bar;
  assign in_1bar = inbar[1];
  assign outbar[0] = in_7bar;
  assign in_7bar = inbar[7];
//assign_done

  assign n20bar = in_7;
  assign n20 = in_7bar;
  assign n19bar = in[3];
  assign n19 = inbar[3];
  assign n18bar = in[2];
  assign n18 = inbar[2];
  assign n17bar = in_0;
  assign n17 = in_0bar;
  OR2_X1 U5 ( .A1(n16), .A2(n15), .ZN(out[4]) );
  AND2_X1 U5bar ( .A1(n16bar), .A2(n15bar), .ZN(outbar[4]) );
  AND2_X1 U6 ( .A1(in[3]), .A2(n20), .ZN(n15) );
  OR2_X1 U6bar ( .A1(inbar[3]), .A2(n20bar), .ZN(n15bar) );
  AND2_X1 U7 ( .A1(in_7), .A2(n19), .ZN(n16) );
  OR2_X1 U7bar ( .A1(in_7bar), .A2(n19bar), .ZN(n16bar) );
  OR2_X1 U8 ( .A1(n14), .A2(n13), .ZN(out[3]) );
  AND2_X1 U8bar ( .A1(n14bar), .A2(n13bar), .ZN(outbar[3]) );
  AND2_X1 U9 ( .A1(in[2]), .A2(n20), .ZN(n13) );
  OR2_X1 U9bar ( .A1(inbar[2]), .A2(n20bar), .ZN(n13bar) );
  AND2_X1 U10 ( .A1(in_7), .A2(n18), .ZN(n14) );
  OR2_X1 U10bar ( .A1(in_7bar), .A2(n18bar), .ZN(n14bar) );
  OR2_X1 U11 ( .A1(n12), .A2(n11), .ZN(out[1]) );
  AND2_X1 U11bar ( .A1(n12bar), .A2(n11bar), .ZN(outbar[1]) );
  AND2_X1 U12 ( .A1(in_0), .A2(n20), .ZN(n11) );
  OR2_X1 U12bar ( .A1(in_0bar), .A2(n20bar), .ZN(n11bar) );
  AND2_X1 U13 ( .A1(in_7), .A2(n17), .ZN(n12) );
  OR2_X1 U13bar ( .A1(in_7bar), .A2(n17bar), .ZN(n12bar) );
endmodule

module scale2_14 ( in, out );

  input wire [7:0] in;
  wire [7:0] inbar;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
//input_done

  output wire [7:0] out;
  wire [7:0] outbar;
//output_done

  wire in_0;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_1;
  wire in_7;
  wire n11;
  wire n12;
  wire n13;
  wire n14;
  wire n15;
  wire n16;
  wire n17;
  wire n18;
  wire n19;
  wire n20;
  wire in_0bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_1bar;
  wire in_7bar;
  wire n11bar;
  wire n12bar;
  wire n13bar;
  wire n14bar;
  wire n15bar;
  wire n16bar;
  wire n17bar;
  wire n18bar;
  wire n19bar;
  wire n20bar;
//wire_done

  assign in_0 = in[0];
  assign out[7] = in_6;
  assign in_6  = in[6];
  assign out[6] = in_5;
  assign in_5  = in[5];
  assign out[5] = in_4;
  assign in_4  = in[4];
  assign out[2] = in_1;
  assign in_1  = in[1];
  assign out[0] = in_7;
  assign in_7  = in[7];
  assign in_0bar = inbar[0];
  assign outbar[7] = in_6bar;
  assign in_6bar = inbar[6];
  assign outbar[6] = in_5bar;
  assign in_5bar = inbar[5];
  assign outbar[5] = in_4bar;
  assign in_4bar = inbar[4];
  assign outbar[2] = in_1bar;
  assign in_1bar = inbar[1];
  assign outbar[0] = in_7bar;
  assign in_7bar = inbar[7];
//assign_done

  assign n20bar = in_7;
  assign n20 = in_7bar;
  assign n19bar = in[3];
  assign n19 = inbar[3];
  assign n18bar = in[2];
  assign n18 = inbar[2];
  assign n17bar = in_0;
  assign n17 = in_0bar;
  OR2_X1 U5 ( .A1(n16), .A2(n15), .ZN(out[4]) );
  AND2_X1 U5bar ( .A1(n16bar), .A2(n15bar), .ZN(outbar[4]) );
  AND2_X1 U6 ( .A1(in[3]), .A2(n20), .ZN(n15) );
  OR2_X1 U6bar ( .A1(inbar[3]), .A2(n20bar), .ZN(n15bar) );
  AND2_X1 U7 ( .A1(in_7), .A2(n19), .ZN(n16) );
  OR2_X1 U7bar ( .A1(in_7bar), .A2(n19bar), .ZN(n16bar) );
  OR2_X1 U8 ( .A1(n14), .A2(n13), .ZN(out[3]) );
  AND2_X1 U8bar ( .A1(n14bar), .A2(n13bar), .ZN(outbar[3]) );
  AND2_X1 U9 ( .A1(in[2]), .A2(n20), .ZN(n13) );
  OR2_X1 U9bar ( .A1(inbar[2]), .A2(n20bar), .ZN(n13bar) );
  AND2_X1 U10 ( .A1(in_7), .A2(n18), .ZN(n14) );
  OR2_X1 U10bar ( .A1(in_7bar), .A2(n18bar), .ZN(n14bar) );
  OR2_X1 U11 ( .A1(n12), .A2(n11), .ZN(out[1]) );
  AND2_X1 U11bar ( .A1(n12bar), .A2(n11bar), .ZN(outbar[1]) );
  AND2_X1 U12 ( .A1(in_0), .A2(n20), .ZN(n11) );
  OR2_X1 U12bar ( .A1(in_0bar), .A2(n20bar), .ZN(n11bar) );
  AND2_X1 U13 ( .A1(in_7), .A2(n17), .ZN(n12) );
  OR2_X1 U13bar ( .A1(in_7bar), .A2(n17bar), .ZN(n12bar) );
endmodule

module scale2_15 ( in, out );

  input wire [7:0] in;
  wire [7:0] inbar;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
//input_done

  output wire [7:0] out;
  wire [7:0] outbar;
//output_done

  wire in_0;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_1;
  wire in_7;
  wire n11;
  wire n12;
  wire n13;
  wire n14;
  wire n15;
  wire n16;
  wire n17;
  wire n18;
  wire n19;
  wire n20;
  wire in_0bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_1bar;
  wire in_7bar;
  wire n11bar;
  wire n12bar;
  wire n13bar;
  wire n14bar;
  wire n15bar;
  wire n16bar;
  wire n17bar;
  wire n18bar;
  wire n19bar;
  wire n20bar;
//wire_done

  assign in_0 = in[0];
  assign out[7] = in_6;
  assign in_6  = in[6];
  assign out[6] = in_5;
  assign in_5  = in[5];
  assign out[5] = in_4;
  assign in_4  = in[4];
  assign out[2] = in_1;
  assign in_1  = in[1];
  assign out[0] = in_7;
  assign in_7  = in[7];
  assign in_0bar = inbar[0];
  assign outbar[7] = in_6bar;
  assign in_6bar = inbar[6];
  assign outbar[6] = in_5bar;
  assign in_5bar = inbar[5];
  assign outbar[5] = in_4bar;
  assign in_4bar = inbar[4];
  assign outbar[2] = in_1bar;
  assign in_1bar = inbar[1];
  assign outbar[0] = in_7bar;
  assign in_7bar = inbar[7];
//assign_done

  assign n20bar = in_7;
  assign n20 = in_7bar;
  assign n19bar = in[3];
  assign n19 = inbar[3];
  assign n18bar = in[2];
  assign n18 = inbar[2];
  assign n17bar = in_0;
  assign n17 = in_0bar;
  OR2_X1 U5 ( .A1(n16), .A2(n15), .ZN(out[4]) );
  AND2_X1 U5bar ( .A1(n16bar), .A2(n15bar), .ZN(outbar[4]) );
  AND2_X1 U6 ( .A1(in[3]), .A2(n20), .ZN(n15) );
  OR2_X1 U6bar ( .A1(inbar[3]), .A2(n20bar), .ZN(n15bar) );
  AND2_X1 U7 ( .A1(in_7), .A2(n19), .ZN(n16) );
  OR2_X1 U7bar ( .A1(in_7bar), .A2(n19bar), .ZN(n16bar) );
  OR2_X1 U8 ( .A1(n14), .A2(n13), .ZN(out[3]) );
  AND2_X1 U8bar ( .A1(n14bar), .A2(n13bar), .ZN(outbar[3]) );
  AND2_X1 U9 ( .A1(in[2]), .A2(n20), .ZN(n13) );
  OR2_X1 U9bar ( .A1(inbar[2]), .A2(n20bar), .ZN(n13bar) );
  AND2_X1 U10 ( .A1(in_7), .A2(n18), .ZN(n14) );
  OR2_X1 U10bar ( .A1(in_7bar), .A2(n18bar), .ZN(n14bar) );
  OR2_X1 U11 ( .A1(n12), .A2(n11), .ZN(out[1]) );
  AND2_X1 U11bar ( .A1(n12bar), .A2(n11bar), .ZN(outbar[1]) );
  AND2_X1 U12 ( .A1(in_0), .A2(n20), .ZN(n11) );
  OR2_X1 U12bar ( .A1(in_0bar), .A2(n20bar), .ZN(n11bar) );
  AND2_X1 U13 ( .A1(in_7), .A2(n17), .ZN(n12) );
  OR2_X1 U13bar ( .A1(in_7bar), .A2(n17bar), .ZN(n12bar) );
endmodule

module byteXor_14 ( a, b, y );

  input wire [7:0] a;
  input wire [7:0] b;
  wire [7:0] abar;
  wire [7:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
//input_done

  output wire [7:0] y;
  wire [7:0] ybar;
//output_done

  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n33bar;
  wire n34bar;
  wire n35bar;
  wire n36bar;
  wire n37bar;
  wire n38bar;
  wire n39bar;
  wire n40bar;
  wire n41bar;
  wire n42bar;
  wire n43bar;
  wire n44bar;
  wire n45bar;
  wire n46bar;
  wire n47bar;
  wire n48bar;
  wire n49bar;
  wire n50bar;
  wire n51bar;
  wire n52bar;
  wire n53bar;
  wire n54bar;
  wire n55bar;
  wire n56bar;
  wire n57bar;
  wire n58bar;
  wire n59bar;
  wire n60bar;
  wire n61bar;
  wire n62bar;
  wire n63bar;
  wire n64bar;
//wire_done

 //assign_done

  assign n64bar = n47;
  assign n64 = n47bar;
  assign n63bar = a[7];
  assign n63 = abar[7];
  assign n62bar = n45;
  assign n62 = n45bar;
  assign n61bar = a[6];
  assign n61 = abar[6];
  assign n60bar = n43;
  assign n60 = n43bar;
  assign n59bar = a[5];
  assign n59 = abar[5];
  assign n58bar = n41;
  assign n58 = n41bar;
  assign n57bar = a[4];
  assign n57 = abar[4];
  assign n56bar = n39;
  assign n56 = n39bar;
  assign n55bar = a[3];
  assign n55 = abar[3];
  assign n54bar = n37;
  assign n54 = n37bar;
  assign n53bar = a[2];
  assign n53 = abar[2];
  assign n52bar = n35;
  assign n52 = n35bar;
  assign n51bar = a[1];
  assign n51 = abar[1];
  assign n50bar = n33;
  assign n50 = n33bar;
  assign n49bar = a[0];
  assign n49 = abar[0];
  OR2_X1 U17 ( .A1(n48), .A2(n64), .ZN(y[7]) );
  AND2_X1 U17bar ( .A1(n48bar), .A2(n64bar), .ZN(ybar[7]) );
  OR2_X1 U18 ( .A1(n63), .A2(b[7]), .ZN(n47) );
  AND2_X1 U18bar ( .A1(n63bar), .A2(bbar[7]), .ZN(n47bar) );
  AND2_X1 U19 ( .A1(b[7]), .A2(n63), .ZN(n48) );
  OR2_X1 U19bar ( .A1(bbar[7]), .A2(n63bar), .ZN(n48bar) );
  OR2_X1 U20 ( .A1(n46), .A2(n62), .ZN(y[6]) );
  AND2_X1 U20bar ( .A1(n46bar), .A2(n62bar), .ZN(ybar[6]) );
  OR2_X1 U21 ( .A1(n61), .A2(b[6]), .ZN(n45) );
  AND2_X1 U21bar ( .A1(n61bar), .A2(bbar[6]), .ZN(n45bar) );
  AND2_X1 U22 ( .A1(b[6]), .A2(n61), .ZN(n46) );
  OR2_X1 U22bar ( .A1(bbar[6]), .A2(n61bar), .ZN(n46bar) );
  OR2_X1 U23 ( .A1(n44), .A2(n60), .ZN(y[5]) );
  AND2_X1 U23bar ( .A1(n44bar), .A2(n60bar), .ZN(ybar[5]) );
  OR2_X1 U24 ( .A1(n59), .A2(b[5]), .ZN(n43) );
  AND2_X1 U24bar ( .A1(n59bar), .A2(bbar[5]), .ZN(n43bar) );
  AND2_X1 U25 ( .A1(b[5]), .A2(n59), .ZN(n44) );
  OR2_X1 U25bar ( .A1(bbar[5]), .A2(n59bar), .ZN(n44bar) );
  OR2_X1 U26 ( .A1(n42), .A2(n58), .ZN(y[4]) );
  AND2_X1 U26bar ( .A1(n42bar), .A2(n58bar), .ZN(ybar[4]) );
  OR2_X1 U27 ( .A1(n57), .A2(b[4]), .ZN(n41) );
  AND2_X1 U27bar ( .A1(n57bar), .A2(bbar[4]), .ZN(n41bar) );
  AND2_X1 U28 ( .A1(b[4]), .A2(n57), .ZN(n42) );
  OR2_X1 U28bar ( .A1(bbar[4]), .A2(n57bar), .ZN(n42bar) );
  OR2_X1 U29 ( .A1(n40), .A2(n56), .ZN(y[3]) );
  AND2_X1 U29bar ( .A1(n40bar), .A2(n56bar), .ZN(ybar[3]) );
  OR2_X1 U30 ( .A1(n55), .A2(b[3]), .ZN(n39) );
  AND2_X1 U30bar ( .A1(n55bar), .A2(bbar[3]), .ZN(n39bar) );
  AND2_X1 U31 ( .A1(b[3]), .A2(n55), .ZN(n40) );
  OR2_X1 U31bar ( .A1(bbar[3]), .A2(n55bar), .ZN(n40bar) );
  OR2_X1 U32 ( .A1(n38), .A2(n54), .ZN(y[2]) );
  AND2_X1 U32bar ( .A1(n38bar), .A2(n54bar), .ZN(ybar[2]) );
  OR2_X1 U33 ( .A1(n53), .A2(b[2]), .ZN(n37) );
  AND2_X1 U33bar ( .A1(n53bar), .A2(bbar[2]), .ZN(n37bar) );
  AND2_X1 U34 ( .A1(b[2]), .A2(n53), .ZN(n38) );
  OR2_X1 U34bar ( .A1(bbar[2]), .A2(n53bar), .ZN(n38bar) );
  OR2_X1 U35 ( .A1(n36), .A2(n52), .ZN(y[1]) );
  AND2_X1 U35bar ( .A1(n36bar), .A2(n52bar), .ZN(ybar[1]) );
  OR2_X1 U36 ( .A1(n51), .A2(b[1]), .ZN(n35) );
  AND2_X1 U36bar ( .A1(n51bar), .A2(bbar[1]), .ZN(n35bar) );
  AND2_X1 U37 ( .A1(b[1]), .A2(n51), .ZN(n36) );
  OR2_X1 U37bar ( .A1(bbar[1]), .A2(n51bar), .ZN(n36bar) );
  OR2_X1 U38 ( .A1(n34), .A2(n50), .ZN(y[0]) );
  AND2_X1 U38bar ( .A1(n34bar), .A2(n50bar), .ZN(ybar[0]) );
  OR2_X1 U39 ( .A1(n49), .A2(b[0]), .ZN(n33) );
  AND2_X1 U39bar ( .A1(n49bar), .A2(bbar[0]), .ZN(n33bar) );
  AND2_X1 U40 ( .A1(b[0]), .A2(n49), .ZN(n34) );
  OR2_X1 U40bar ( .A1(bbar[0]), .A2(n49bar), .ZN(n34bar) );
endmodule

module byteXor_15 ( a, b, y );

  input wire [7:0] a;
  input wire [7:0] b;
  wire [7:0] abar;
  wire [7:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
//input_done

  output wire [7:0] y;
  wire [7:0] ybar;
//output_done

  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n33bar;
  wire n34bar;
  wire n35bar;
  wire n36bar;
  wire n37bar;
  wire n38bar;
  wire n39bar;
  wire n40bar;
  wire n41bar;
  wire n42bar;
  wire n43bar;
  wire n44bar;
  wire n45bar;
  wire n46bar;
  wire n47bar;
  wire n48bar;
  wire n49bar;
  wire n50bar;
  wire n51bar;
  wire n52bar;
  wire n53bar;
  wire n54bar;
  wire n55bar;
  wire n56bar;
  wire n57bar;
  wire n58bar;
  wire n59bar;
  wire n60bar;
  wire n61bar;
  wire n62bar;
  wire n63bar;
  wire n64bar;
//wire_done

 //assign_done

  assign n64bar = n47;
  assign n64 = n47bar;
  assign n63bar = a[7];
  assign n63 = abar[7];
  assign n62bar = n45;
  assign n62 = n45bar;
  assign n61bar = a[6];
  assign n61 = abar[6];
  assign n60bar = n43;
  assign n60 = n43bar;
  assign n59bar = a[5];
  assign n59 = abar[5];
  assign n58bar = n41;
  assign n58 = n41bar;
  assign n57bar = a[4];
  assign n57 = abar[4];
  assign n56bar = n39;
  assign n56 = n39bar;
  assign n55bar = a[3];
  assign n55 = abar[3];
  assign n54bar = n37;
  assign n54 = n37bar;
  assign n53bar = a[2];
  assign n53 = abar[2];
  assign n52bar = n35;
  assign n52 = n35bar;
  assign n51bar = a[1];
  assign n51 = abar[1];
  assign n50bar = n33;
  assign n50 = n33bar;
  assign n49bar = a[0];
  assign n49 = abar[0];
  OR2_X1 U17 ( .A1(n48), .A2(n64), .ZN(y[7]) );
  AND2_X1 U17bar ( .A1(n48bar), .A2(n64bar), .ZN(ybar[7]) );
  OR2_X1 U18 ( .A1(n63), .A2(b[7]), .ZN(n47) );
  AND2_X1 U18bar ( .A1(n63bar), .A2(bbar[7]), .ZN(n47bar) );
  AND2_X1 U19 ( .A1(b[7]), .A2(n63), .ZN(n48) );
  OR2_X1 U19bar ( .A1(bbar[7]), .A2(n63bar), .ZN(n48bar) );
  OR2_X1 U20 ( .A1(n46), .A2(n62), .ZN(y[6]) );
  AND2_X1 U20bar ( .A1(n46bar), .A2(n62bar), .ZN(ybar[6]) );
  OR2_X1 U21 ( .A1(n61), .A2(b[6]), .ZN(n45) );
  AND2_X1 U21bar ( .A1(n61bar), .A2(bbar[6]), .ZN(n45bar) );
  AND2_X1 U22 ( .A1(b[6]), .A2(n61), .ZN(n46) );
  OR2_X1 U22bar ( .A1(bbar[6]), .A2(n61bar), .ZN(n46bar) );
  OR2_X1 U23 ( .A1(n44), .A2(n60), .ZN(y[5]) );
  AND2_X1 U23bar ( .A1(n44bar), .A2(n60bar), .ZN(ybar[5]) );
  OR2_X1 U24 ( .A1(n59), .A2(b[5]), .ZN(n43) );
  AND2_X1 U24bar ( .A1(n59bar), .A2(bbar[5]), .ZN(n43bar) );
  AND2_X1 U25 ( .A1(b[5]), .A2(n59), .ZN(n44) );
  OR2_X1 U25bar ( .A1(bbar[5]), .A2(n59bar), .ZN(n44bar) );
  OR2_X1 U26 ( .A1(n42), .A2(n58), .ZN(y[4]) );
  AND2_X1 U26bar ( .A1(n42bar), .A2(n58bar), .ZN(ybar[4]) );
  OR2_X1 U27 ( .A1(n57), .A2(b[4]), .ZN(n41) );
  AND2_X1 U27bar ( .A1(n57bar), .A2(bbar[4]), .ZN(n41bar) );
  AND2_X1 U28 ( .A1(b[4]), .A2(n57), .ZN(n42) );
  OR2_X1 U28bar ( .A1(bbar[4]), .A2(n57bar), .ZN(n42bar) );
  OR2_X1 U29 ( .A1(n40), .A2(n56), .ZN(y[3]) );
  AND2_X1 U29bar ( .A1(n40bar), .A2(n56bar), .ZN(ybar[3]) );
  OR2_X1 U30 ( .A1(n55), .A2(b[3]), .ZN(n39) );
  AND2_X1 U30bar ( .A1(n55bar), .A2(bbar[3]), .ZN(n39bar) );
  AND2_X1 U31 ( .A1(b[3]), .A2(n55), .ZN(n40) );
  OR2_X1 U31bar ( .A1(bbar[3]), .A2(n55bar), .ZN(n40bar) );
  OR2_X1 U32 ( .A1(n38), .A2(n54), .ZN(y[2]) );
  AND2_X1 U32bar ( .A1(n38bar), .A2(n54bar), .ZN(ybar[2]) );
  OR2_X1 U33 ( .A1(n53), .A2(b[2]), .ZN(n37) );
  AND2_X1 U33bar ( .A1(n53bar), .A2(bbar[2]), .ZN(n37bar) );
  AND2_X1 U34 ( .A1(b[2]), .A2(n53), .ZN(n38) );
  OR2_X1 U34bar ( .A1(bbar[2]), .A2(n53bar), .ZN(n38bar) );
  OR2_X1 U35 ( .A1(n36), .A2(n52), .ZN(y[1]) );
  AND2_X1 U35bar ( .A1(n36bar), .A2(n52bar), .ZN(ybar[1]) );
  OR2_X1 U36 ( .A1(n51), .A2(b[1]), .ZN(n35) );
  AND2_X1 U36bar ( .A1(n51bar), .A2(bbar[1]), .ZN(n35bar) );
  AND2_X1 U37 ( .A1(b[1]), .A2(n51), .ZN(n36) );
  OR2_X1 U37bar ( .A1(bbar[1]), .A2(n51bar), .ZN(n36bar) );
  OR2_X1 U38 ( .A1(n34), .A2(n50), .ZN(y[0]) );
  AND2_X1 U38bar ( .A1(n34bar), .A2(n50bar), .ZN(ybar[0]) );
  OR2_X1 U39 ( .A1(n49), .A2(b[0]), .ZN(n33) );
  AND2_X1 U39bar ( .A1(n49bar), .A2(bbar[0]), .ZN(n33bar) );
  AND2_X1 U40 ( .A1(b[0]), .A2(n49), .ZN(n34) );
  OR2_X1 U40bar ( .A1(bbar[0]), .A2(n49bar), .ZN(n34bar) );
endmodule

module byteXor_16 ( a, b, y );

  input wire [7:0] a;
  input wire [7:0] b;
  wire [7:0] abar;
  wire [7:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
//input_done

  output wire [7:0] y;
  wire [7:0] ybar;
//output_done

  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n33bar;
  wire n34bar;
  wire n35bar;
  wire n36bar;
  wire n37bar;
  wire n38bar;
  wire n39bar;
  wire n40bar;
  wire n41bar;
  wire n42bar;
  wire n43bar;
  wire n44bar;
  wire n45bar;
  wire n46bar;
  wire n47bar;
  wire n48bar;
  wire n49bar;
  wire n50bar;
  wire n51bar;
  wire n52bar;
  wire n53bar;
  wire n54bar;
  wire n55bar;
  wire n56bar;
  wire n57bar;
  wire n58bar;
  wire n59bar;
  wire n60bar;
  wire n61bar;
  wire n62bar;
  wire n63bar;
  wire n64bar;
//wire_done

 //assign_done

  assign n64bar = n47;
  assign n64 = n47bar;
  assign n63bar = a[7];
  assign n63 = abar[7];
  assign n62bar = n45;
  assign n62 = n45bar;
  assign n61bar = a[6];
  assign n61 = abar[6];
  assign n60bar = n43;
  assign n60 = n43bar;
  assign n59bar = a[5];
  assign n59 = abar[5];
  assign n58bar = n41;
  assign n58 = n41bar;
  assign n57bar = a[4];
  assign n57 = abar[4];
  assign n56bar = n39;
  assign n56 = n39bar;
  assign n55bar = a[3];
  assign n55 = abar[3];
  assign n54bar = n37;
  assign n54 = n37bar;
  assign n53bar = a[2];
  assign n53 = abar[2];
  assign n52bar = n35;
  assign n52 = n35bar;
  assign n51bar = a[1];
  assign n51 = abar[1];
  assign n50bar = n33;
  assign n50 = n33bar;
  assign n49bar = a[0];
  assign n49 = abar[0];
  OR2_X1 U17 ( .A1(n48), .A2(n64), .ZN(y[7]) );
  AND2_X1 U17bar ( .A1(n48bar), .A2(n64bar), .ZN(ybar[7]) );
  OR2_X1 U18 ( .A1(n63), .A2(b[7]), .ZN(n47) );
  AND2_X1 U18bar ( .A1(n63bar), .A2(bbar[7]), .ZN(n47bar) );
  AND2_X1 U19 ( .A1(b[7]), .A2(n63), .ZN(n48) );
  OR2_X1 U19bar ( .A1(bbar[7]), .A2(n63bar), .ZN(n48bar) );
  OR2_X1 U20 ( .A1(n46), .A2(n62), .ZN(y[6]) );
  AND2_X1 U20bar ( .A1(n46bar), .A2(n62bar), .ZN(ybar[6]) );
  OR2_X1 U21 ( .A1(n61), .A2(b[6]), .ZN(n45) );
  AND2_X1 U21bar ( .A1(n61bar), .A2(bbar[6]), .ZN(n45bar) );
  AND2_X1 U22 ( .A1(b[6]), .A2(n61), .ZN(n46) );
  OR2_X1 U22bar ( .A1(bbar[6]), .A2(n61bar), .ZN(n46bar) );
  OR2_X1 U23 ( .A1(n44), .A2(n60), .ZN(y[5]) );
  AND2_X1 U23bar ( .A1(n44bar), .A2(n60bar), .ZN(ybar[5]) );
  OR2_X1 U24 ( .A1(n59), .A2(b[5]), .ZN(n43) );
  AND2_X1 U24bar ( .A1(n59bar), .A2(bbar[5]), .ZN(n43bar) );
  AND2_X1 U25 ( .A1(b[5]), .A2(n59), .ZN(n44) );
  OR2_X1 U25bar ( .A1(bbar[5]), .A2(n59bar), .ZN(n44bar) );
  OR2_X1 U26 ( .A1(n42), .A2(n58), .ZN(y[4]) );
  AND2_X1 U26bar ( .A1(n42bar), .A2(n58bar), .ZN(ybar[4]) );
  OR2_X1 U27 ( .A1(n57), .A2(b[4]), .ZN(n41) );
  AND2_X1 U27bar ( .A1(n57bar), .A2(bbar[4]), .ZN(n41bar) );
  AND2_X1 U28 ( .A1(b[4]), .A2(n57), .ZN(n42) );
  OR2_X1 U28bar ( .A1(bbar[4]), .A2(n57bar), .ZN(n42bar) );
  OR2_X1 U29 ( .A1(n40), .A2(n56), .ZN(y[3]) );
  AND2_X1 U29bar ( .A1(n40bar), .A2(n56bar), .ZN(ybar[3]) );
  OR2_X1 U30 ( .A1(n55), .A2(b[3]), .ZN(n39) );
  AND2_X1 U30bar ( .A1(n55bar), .A2(bbar[3]), .ZN(n39bar) );
  AND2_X1 U31 ( .A1(b[3]), .A2(n55), .ZN(n40) );
  OR2_X1 U31bar ( .A1(bbar[3]), .A2(n55bar), .ZN(n40bar) );
  OR2_X1 U32 ( .A1(n38), .A2(n54), .ZN(y[2]) );
  AND2_X1 U32bar ( .A1(n38bar), .A2(n54bar), .ZN(ybar[2]) );
  OR2_X1 U33 ( .A1(n53), .A2(b[2]), .ZN(n37) );
  AND2_X1 U33bar ( .A1(n53bar), .A2(bbar[2]), .ZN(n37bar) );
  AND2_X1 U34 ( .A1(b[2]), .A2(n53), .ZN(n38) );
  OR2_X1 U34bar ( .A1(bbar[2]), .A2(n53bar), .ZN(n38bar) );
  OR2_X1 U35 ( .A1(n36), .A2(n52), .ZN(y[1]) );
  AND2_X1 U35bar ( .A1(n36bar), .A2(n52bar), .ZN(ybar[1]) );
  OR2_X1 U36 ( .A1(n51), .A2(b[1]), .ZN(n35) );
  AND2_X1 U36bar ( .A1(n51bar), .A2(bbar[1]), .ZN(n35bar) );
  AND2_X1 U37 ( .A1(b[1]), .A2(n51), .ZN(n36) );
  OR2_X1 U37bar ( .A1(bbar[1]), .A2(n51bar), .ZN(n36bar) );
  OR2_X1 U38 ( .A1(n34), .A2(n50), .ZN(y[0]) );
  AND2_X1 U38bar ( .A1(n34bar), .A2(n50bar), .ZN(ybar[0]) );
  OR2_X1 U39 ( .A1(n49), .A2(b[0]), .ZN(n33) );
  AND2_X1 U39bar ( .A1(n49bar), .A2(bbar[0]), .ZN(n33bar) );
  AND2_X1 U40 ( .A1(b[0]), .A2(n49), .ZN(n34) );
  OR2_X1 U40bar ( .A1(bbar[0]), .A2(n49bar), .ZN(n34bar) );
endmodule

module byteXor4_13 ( a, b, c, d, y );

  input wire [7:0] a;
  input wire [7:0] b;
  input wire [7:0] c;
  input wire [7:0] d;
  wire [7:0] abar;
  wire [7:0] bbar;
  wire [7:0] cbar;
  wire [7:0] dbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign cbar[0] = ~c[0];
  assign cbar[1] = ~c[1];
  assign cbar[2] = ~c[2];
  assign cbar[3] = ~c[3];
  assign cbar[4] = ~c[4];
  assign cbar[5] = ~c[5];
  assign cbar[6] = ~c[6];
  assign cbar[7] = ~c[7];
  assign dbar[0] = ~d[0];
  assign dbar[1] = ~d[1];
  assign dbar[2] = ~d[2];
  assign dbar[3] = ~d[3];
  assign dbar[4] = ~d[4];
  assign dbar[5] = ~d[5];
  assign dbar[6] = ~d[6];
  assign dbar[7] = ~d[7];
//input_done

  output wire [7:0] y;
  wire [7:0] ybar;
//output_done

  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n113bar;
  wire n114bar;
  wire n115bar;
  wire n116bar;
  wire n117bar;
  wire n118bar;
  wire n119bar;
  wire n120bar;
  wire n121bar;
  wire n122bar;
  wire n123bar;
  wire n124bar;
  wire n125bar;
  wire n126bar;
  wire n127bar;
  wire n128bar;
  wire n129bar;
  wire n130bar;
  wire n131bar;
  wire n132bar;
  wire n133bar;
  wire n134bar;
  wire n135bar;
  wire n136bar;
  wire n137bar;
  wire n138bar;
  wire n139bar;
  wire n140bar;
  wire n141bar;
  wire n142bar;
  wire n143bar;
  wire n144bar;
  wire n145bar;
  wire n146bar;
  wire n147bar;
  wire n148bar;
  wire n149bar;
  wire n150bar;
  wire n151bar;
  wire n152bar;
  wire n153bar;
  wire n154bar;
  wire n155bar;
  wire n156bar;
  wire n157bar;
  wire n158bar;
  wire n159bar;
  wire n160bar;
  wire n161bar;
  wire n162bar;
  wire n163bar;
  wire n164bar;
  wire n165bar;
  wire n166bar;
  wire n167bar;
  wire n168bar;
  wire n169bar;
  wire n170bar;
  wire n171bar;
  wire n172bar;
  wire n173bar;
  wire n174bar;
  wire n175bar;
  wire n176bar;
  wire n177bar;
  wire n178bar;
  wire n179bar;
  wire n180bar;
  wire n181bar;
  wire n182bar;
  wire n183bar;
  wire n184bar;
  wire n185bar;
  wire n186bar;
  wire n187bar;
  wire n188bar;
  wire n189bar;
  wire n190bar;
  wire n191bar;
  wire n192bar;
  wire n193bar;
  wire n194bar;
  wire n195bar;
  wire n196bar;
  wire n197bar;
  wire n198bar;
  wire n199bar;
  wire n200bar;
  wire n201bar;
  wire n202bar;
  wire n203bar;
  wire n204bar;
  wire n205bar;
  wire n206bar;
  wire n207bar;
  wire n208bar;
  wire n209bar;
  wire n210bar;
  wire n211bar;
  wire n212bar;
  wire n213bar;
  wire n214bar;
  wire n215bar;
  wire n216bar;
  wire n217bar;
  wire n218bar;
  wire n219bar;
  wire n220bar;
  wire n221bar;
  wire n222bar;
  wire n223bar;
  wire n224bar;
//wire_done

 //assign_done

  assign n224bar = n175;
  assign n224 = n175bar;
  assign n223bar = a[7];
  assign n223 = abar[7];
  assign n222bar = n167;
  assign n222 = n167bar;
  assign n221bar = a[6];
  assign n221 = abar[6];
  assign n220bar = n159;
  assign n220 = n159bar;
  assign n219bar = a[5];
  assign n219 = abar[5];
  assign n218bar = n151;
  assign n218 = n151bar;
  assign n217bar = a[4];
  assign n217 = abar[4];
  assign n216bar = n143;
  assign n216 = n143bar;
  assign n215bar = a[3];
  assign n215 = abar[3];
  assign n214bar = n135;
  assign n214 = n135bar;
  assign n213bar = a[2];
  assign n213 = abar[2];
  assign n212bar = n127;
  assign n212 = n127bar;
  assign n211bar = a[1];
  assign n211 = abar[1];
  assign n210bar = n119;
  assign n210 = n119bar;
  assign n209bar = a[0];
  assign n209 = abar[0];
  assign n208bar = b[7];
  assign n208 = bbar[7];
  assign n207bar = b[6];
  assign n207 = bbar[6];
  assign n206bar = b[5];
  assign n206 = bbar[5];
  assign n205bar = b[4];
  assign n205 = bbar[4];
  assign n204bar = b[3];
  assign n204 = bbar[3];
  assign n203bar = b[2];
  assign n203 = bbar[2];
  assign n202bar = b[1];
  assign n202 = bbar[1];
  assign n201bar = b[0];
  assign n201 = bbar[0];
  assign n200bar = n171;
  assign n200 = n171bar;
  assign n199bar = c[7];
  assign n199 = cbar[7];
  assign n198bar = n163;
  assign n198 = n163bar;
  assign n197bar = c[6];
  assign n197 = cbar[6];
  assign n196bar = n155;
  assign n196 = n155bar;
  assign n195bar = c[5];
  assign n195 = cbar[5];
  assign n194bar = n147;
  assign n194 = n147bar;
  assign n193bar = c[4];
  assign n193 = cbar[4];
  assign n192bar = n139;
  assign n192 = n139bar;
  assign n191bar = c[3];
  assign n191 = cbar[3];
  assign n190bar = n131;
  assign n190 = n131bar;
  assign n189bar = c[2];
  assign n189 = cbar[2];
  assign n188bar = n123;
  assign n188 = n123bar;
  assign n187bar = c[1];
  assign n187 = cbar[1];
  assign n186bar = n115;
  assign n186 = n115bar;
  assign n185bar = c[0];
  assign n185 = cbar[0];
  assign n184bar = d[7];
  assign n184 = dbar[7];
  assign n183bar = d[6];
  assign n183 = dbar[6];
  assign n182bar = d[5];
  assign n182 = dbar[5];
  assign n181bar = d[4];
  assign n181 = dbar[4];
  assign n180bar = d[3];
  assign n180 = dbar[3];
  assign n179bar = d[2];
  assign n179 = dbar[2];
  assign n178bar = d[1];
  assign n178 = dbar[1];
  assign n177bar = d[0];
  assign n177 = dbar[0];
  OR2_X1 U49 ( .A1(n176), .A2(n224), .ZN(y[7]) );
  AND2_X1 U49bar ( .A1(n176bar), .A2(n224bar), .ZN(ybar[7]) );
  OR2_X1 U50 ( .A1(n174), .A2(n200), .ZN(n175) );
  AND2_X1 U50bar ( .A1(n174bar), .A2(n200bar), .ZN(n175bar) );
  AND2_X1 U51 ( .A1(n200), .A2(n174), .ZN(n176) );
  OR2_X1 U51bar ( .A1(n200bar), .A2(n174bar), .ZN(n176bar) );
  AND2_X1 U52 ( .A1(n173), .A2(n172), .ZN(n174) );
  OR2_X1 U52bar ( .A1(n173bar), .A2(n172bar), .ZN(n174bar) );
  OR2_X1 U53 ( .A1(n223), .A2(b[7]), .ZN(n172) );
  AND2_X1 U53bar ( .A1(n223bar), .A2(bbar[7]), .ZN(n172bar) );
  OR2_X1 U54 ( .A1(n208), .A2(a[7]), .ZN(n173) );
  AND2_X1 U54bar ( .A1(n208bar), .A2(abar[7]), .ZN(n173bar) );
  AND2_X1 U55 ( .A1(n170), .A2(n169), .ZN(n171) );
  OR2_X1 U55bar ( .A1(n170bar), .A2(n169bar), .ZN(n171bar) );
  OR2_X1 U56 ( .A1(n199), .A2(d[7]), .ZN(n169) );
  AND2_X1 U56bar ( .A1(n199bar), .A2(dbar[7]), .ZN(n169bar) );
  OR2_X1 U57 ( .A1(n184), .A2(c[7]), .ZN(n170) );
  AND2_X1 U57bar ( .A1(n184bar), .A2(cbar[7]), .ZN(n170bar) );
  OR2_X1 U58 ( .A1(n168), .A2(n222), .ZN(y[6]) );
  AND2_X1 U58bar ( .A1(n168bar), .A2(n222bar), .ZN(ybar[6]) );
  OR2_X1 U59 ( .A1(n166), .A2(n198), .ZN(n167) );
  AND2_X1 U59bar ( .A1(n166bar), .A2(n198bar), .ZN(n167bar) );
  AND2_X1 U60 ( .A1(n198), .A2(n166), .ZN(n168) );
  OR2_X1 U60bar ( .A1(n198bar), .A2(n166bar), .ZN(n168bar) );
  AND2_X1 U61 ( .A1(n165), .A2(n164), .ZN(n166) );
  OR2_X1 U61bar ( .A1(n165bar), .A2(n164bar), .ZN(n166bar) );
  OR2_X1 U62 ( .A1(n221), .A2(b[6]), .ZN(n164) );
  AND2_X1 U62bar ( .A1(n221bar), .A2(bbar[6]), .ZN(n164bar) );
  OR2_X1 U63 ( .A1(n207), .A2(a[6]), .ZN(n165) );
  AND2_X1 U63bar ( .A1(n207bar), .A2(abar[6]), .ZN(n165bar) );
  AND2_X1 U64 ( .A1(n162), .A2(n161), .ZN(n163) );
  OR2_X1 U64bar ( .A1(n162bar), .A2(n161bar), .ZN(n163bar) );
  OR2_X1 U65 ( .A1(n197), .A2(d[6]), .ZN(n161) );
  AND2_X1 U65bar ( .A1(n197bar), .A2(dbar[6]), .ZN(n161bar) );
  OR2_X1 U66 ( .A1(n183), .A2(c[6]), .ZN(n162) );
  AND2_X1 U66bar ( .A1(n183bar), .A2(cbar[6]), .ZN(n162bar) );
  OR2_X1 U67 ( .A1(n160), .A2(n220), .ZN(y[5]) );
  AND2_X1 U67bar ( .A1(n160bar), .A2(n220bar), .ZN(ybar[5]) );
  OR2_X1 U68 ( .A1(n158), .A2(n196), .ZN(n159) );
  AND2_X1 U68bar ( .A1(n158bar), .A2(n196bar), .ZN(n159bar) );
  AND2_X1 U69 ( .A1(n196), .A2(n158), .ZN(n160) );
  OR2_X1 U69bar ( .A1(n196bar), .A2(n158bar), .ZN(n160bar) );
  AND2_X1 U70 ( .A1(n157), .A2(n156), .ZN(n158) );
  OR2_X1 U70bar ( .A1(n157bar), .A2(n156bar), .ZN(n158bar) );
  OR2_X1 U71 ( .A1(n219), .A2(b[5]), .ZN(n156) );
  AND2_X1 U71bar ( .A1(n219bar), .A2(bbar[5]), .ZN(n156bar) );
  OR2_X1 U72 ( .A1(n206), .A2(a[5]), .ZN(n157) );
  AND2_X1 U72bar ( .A1(n206bar), .A2(abar[5]), .ZN(n157bar) );
  AND2_X1 U73 ( .A1(n154), .A2(n153), .ZN(n155) );
  OR2_X1 U73bar ( .A1(n154bar), .A2(n153bar), .ZN(n155bar) );
  OR2_X1 U74 ( .A1(n195), .A2(d[5]), .ZN(n153) );
  AND2_X1 U74bar ( .A1(n195bar), .A2(dbar[5]), .ZN(n153bar) );
  OR2_X1 U75 ( .A1(n182), .A2(c[5]), .ZN(n154) );
  AND2_X1 U75bar ( .A1(n182bar), .A2(cbar[5]), .ZN(n154bar) );
  OR2_X1 U76 ( .A1(n152), .A2(n218), .ZN(y[4]) );
  AND2_X1 U76bar ( .A1(n152bar), .A2(n218bar), .ZN(ybar[4]) );
  OR2_X1 U77 ( .A1(n150), .A2(n194), .ZN(n151) );
  AND2_X1 U77bar ( .A1(n150bar), .A2(n194bar), .ZN(n151bar) );
  AND2_X1 U78 ( .A1(n194), .A2(n150), .ZN(n152) );
  OR2_X1 U78bar ( .A1(n194bar), .A2(n150bar), .ZN(n152bar) );
  AND2_X1 U79 ( .A1(n149), .A2(n148), .ZN(n150) );
  OR2_X1 U79bar ( .A1(n149bar), .A2(n148bar), .ZN(n150bar) );
  OR2_X1 U80 ( .A1(n217), .A2(b[4]), .ZN(n148) );
  AND2_X1 U80bar ( .A1(n217bar), .A2(bbar[4]), .ZN(n148bar) );
  OR2_X1 U81 ( .A1(n205), .A2(a[4]), .ZN(n149) );
  AND2_X1 U81bar ( .A1(n205bar), .A2(abar[4]), .ZN(n149bar) );
  AND2_X1 U82 ( .A1(n146), .A2(n145), .ZN(n147) );
  OR2_X1 U82bar ( .A1(n146bar), .A2(n145bar), .ZN(n147bar) );
  OR2_X1 U83 ( .A1(n193), .A2(d[4]), .ZN(n145) );
  AND2_X1 U83bar ( .A1(n193bar), .A2(dbar[4]), .ZN(n145bar) );
  OR2_X1 U84 ( .A1(n181), .A2(c[4]), .ZN(n146) );
  AND2_X1 U84bar ( .A1(n181bar), .A2(cbar[4]), .ZN(n146bar) );
  OR2_X1 U85 ( .A1(n144), .A2(n216), .ZN(y[3]) );
  AND2_X1 U85bar ( .A1(n144bar), .A2(n216bar), .ZN(ybar[3]) );
  OR2_X1 U86 ( .A1(n142), .A2(n192), .ZN(n143) );
  AND2_X1 U86bar ( .A1(n142bar), .A2(n192bar), .ZN(n143bar) );
  AND2_X1 U87 ( .A1(n192), .A2(n142), .ZN(n144) );
  OR2_X1 U87bar ( .A1(n192bar), .A2(n142bar), .ZN(n144bar) );
  AND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(n142) );
  OR2_X1 U88bar ( .A1(n141bar), .A2(n140bar), .ZN(n142bar) );
  OR2_X1 U89 ( .A1(n215), .A2(b[3]), .ZN(n140) );
  AND2_X1 U89bar ( .A1(n215bar), .A2(bbar[3]), .ZN(n140bar) );
  OR2_X1 U90 ( .A1(n204), .A2(a[3]), .ZN(n141) );
  AND2_X1 U90bar ( .A1(n204bar), .A2(abar[3]), .ZN(n141bar) );
  AND2_X1 U91 ( .A1(n138), .A2(n137), .ZN(n139) );
  OR2_X1 U91bar ( .A1(n138bar), .A2(n137bar), .ZN(n139bar) );
  OR2_X1 U92 ( .A1(n191), .A2(d[3]), .ZN(n137) );
  AND2_X1 U92bar ( .A1(n191bar), .A2(dbar[3]), .ZN(n137bar) );
  OR2_X1 U93 ( .A1(n180), .A2(c[3]), .ZN(n138) );
  AND2_X1 U93bar ( .A1(n180bar), .A2(cbar[3]), .ZN(n138bar) );
  OR2_X1 U94 ( .A1(n136), .A2(n214), .ZN(y[2]) );
  AND2_X1 U94bar ( .A1(n136bar), .A2(n214bar), .ZN(ybar[2]) );
  OR2_X1 U95 ( .A1(n134), .A2(n190), .ZN(n135) );
  AND2_X1 U95bar ( .A1(n134bar), .A2(n190bar), .ZN(n135bar) );
  AND2_X1 U96 ( .A1(n190), .A2(n134), .ZN(n136) );
  OR2_X1 U96bar ( .A1(n190bar), .A2(n134bar), .ZN(n136bar) );
  AND2_X1 U97 ( .A1(n133), .A2(n132), .ZN(n134) );
  OR2_X1 U97bar ( .A1(n133bar), .A2(n132bar), .ZN(n134bar) );
  OR2_X1 U98 ( .A1(n213), .A2(b[2]), .ZN(n132) );
  AND2_X1 U98bar ( .A1(n213bar), .A2(bbar[2]), .ZN(n132bar) );
  OR2_X1 U99 ( .A1(n203), .A2(a[2]), .ZN(n133) );
  AND2_X1 U99bar ( .A1(n203bar), .A2(abar[2]), .ZN(n133bar) );
  AND2_X1 U100 ( .A1(n130), .A2(n129), .ZN(n131) );
  OR2_X1 U100bar ( .A1(n130bar), .A2(n129bar), .ZN(n131bar) );
  OR2_X1 U101 ( .A1(n189), .A2(d[2]), .ZN(n129) );
  AND2_X1 U101bar ( .A1(n189bar), .A2(dbar[2]), .ZN(n129bar) );
  OR2_X1 U102 ( .A1(n179), .A2(c[2]), .ZN(n130) );
  AND2_X1 U102bar ( .A1(n179bar), .A2(cbar[2]), .ZN(n130bar) );
  OR2_X1 U103 ( .A1(n128), .A2(n212), .ZN(y[1]) );
  AND2_X1 U103bar ( .A1(n128bar), .A2(n212bar), .ZN(ybar[1]) );
  OR2_X1 U104 ( .A1(n126), .A2(n188), .ZN(n127) );
  AND2_X1 U104bar ( .A1(n126bar), .A2(n188bar), .ZN(n127bar) );
  AND2_X1 U105 ( .A1(n188), .A2(n126), .ZN(n128) );
  OR2_X1 U105bar ( .A1(n188bar), .A2(n126bar), .ZN(n128bar) );
  AND2_X1 U106 ( .A1(n125), .A2(n124), .ZN(n126) );
  OR2_X1 U106bar ( .A1(n125bar), .A2(n124bar), .ZN(n126bar) );
  OR2_X1 U107 ( .A1(n211), .A2(b[1]), .ZN(n124) );
  AND2_X1 U107bar ( .A1(n211bar), .A2(bbar[1]), .ZN(n124bar) );
  OR2_X1 U108 ( .A1(n202), .A2(a[1]), .ZN(n125) );
  AND2_X1 U108bar ( .A1(n202bar), .A2(abar[1]), .ZN(n125bar) );
  AND2_X1 U109 ( .A1(n122), .A2(n121), .ZN(n123) );
  OR2_X1 U109bar ( .A1(n122bar), .A2(n121bar), .ZN(n123bar) );
  OR2_X1 U110 ( .A1(n187), .A2(d[1]), .ZN(n121) );
  AND2_X1 U110bar ( .A1(n187bar), .A2(dbar[1]), .ZN(n121bar) );
  OR2_X1 U111 ( .A1(n178), .A2(c[1]), .ZN(n122) );
  AND2_X1 U111bar ( .A1(n178bar), .A2(cbar[1]), .ZN(n122bar) );
  OR2_X1 U112 ( .A1(n120), .A2(n210), .ZN(y[0]) );
  AND2_X1 U112bar ( .A1(n120bar), .A2(n210bar), .ZN(ybar[0]) );
  OR2_X1 U113 ( .A1(n118), .A2(n186), .ZN(n119) );
  AND2_X1 U113bar ( .A1(n118bar), .A2(n186bar), .ZN(n119bar) );
  AND2_X1 U114 ( .A1(n186), .A2(n118), .ZN(n120) );
  OR2_X1 U114bar ( .A1(n186bar), .A2(n118bar), .ZN(n120bar) );
  AND2_X1 U115 ( .A1(n117), .A2(n116), .ZN(n118) );
  OR2_X1 U115bar ( .A1(n117bar), .A2(n116bar), .ZN(n118bar) );
  OR2_X1 U116 ( .A1(n209), .A2(b[0]), .ZN(n116) );
  AND2_X1 U116bar ( .A1(n209bar), .A2(bbar[0]), .ZN(n116bar) );
  OR2_X1 U117 ( .A1(n201), .A2(a[0]), .ZN(n117) );
  AND2_X1 U117bar ( .A1(n201bar), .A2(abar[0]), .ZN(n117bar) );
  AND2_X1 U118 ( .A1(n114), .A2(n113), .ZN(n115) );
  OR2_X1 U118bar ( .A1(n114bar), .A2(n113bar), .ZN(n115bar) );
  OR2_X1 U119 ( .A1(n185), .A2(d[0]), .ZN(n113) );
  AND2_X1 U119bar ( .A1(n185bar), .A2(dbar[0]), .ZN(n113bar) );
  OR2_X1 U120 ( .A1(n177), .A2(c[0]), .ZN(n114) );
  AND2_X1 U120bar ( .A1(n177bar), .A2(cbar[0]), .ZN(n114bar) );
endmodule

module byteXor4_14 ( a, b, c, d, y );

  input wire [7:0] a;
  input wire [7:0] b;
  input wire [7:0] c;
  input wire [7:0] d;
  wire [7:0] abar;
  wire [7:0] bbar;
  wire [7:0] cbar;
  wire [7:0] dbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign cbar[0] = ~c[0];
  assign cbar[1] = ~c[1];
  assign cbar[2] = ~c[2];
  assign cbar[3] = ~c[3];
  assign cbar[4] = ~c[4];
  assign cbar[5] = ~c[5];
  assign cbar[6] = ~c[6];
  assign cbar[7] = ~c[7];
  assign dbar[0] = ~d[0];
  assign dbar[1] = ~d[1];
  assign dbar[2] = ~d[2];
  assign dbar[3] = ~d[3];
  assign dbar[4] = ~d[4];
  assign dbar[5] = ~d[5];
  assign dbar[6] = ~d[6];
  assign dbar[7] = ~d[7];
//input_done

  output wire [7:0] y;
  wire [7:0] ybar;
//output_done

  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n113bar;
  wire n114bar;
  wire n115bar;
  wire n116bar;
  wire n117bar;
  wire n118bar;
  wire n119bar;
  wire n120bar;
  wire n121bar;
  wire n122bar;
  wire n123bar;
  wire n124bar;
  wire n125bar;
  wire n126bar;
  wire n127bar;
  wire n128bar;
  wire n129bar;
  wire n130bar;
  wire n131bar;
  wire n132bar;
  wire n133bar;
  wire n134bar;
  wire n135bar;
  wire n136bar;
  wire n137bar;
  wire n138bar;
  wire n139bar;
  wire n140bar;
  wire n141bar;
  wire n142bar;
  wire n143bar;
  wire n144bar;
  wire n145bar;
  wire n146bar;
  wire n147bar;
  wire n148bar;
  wire n149bar;
  wire n150bar;
  wire n151bar;
  wire n152bar;
  wire n153bar;
  wire n154bar;
  wire n155bar;
  wire n156bar;
  wire n157bar;
  wire n158bar;
  wire n159bar;
  wire n160bar;
  wire n161bar;
  wire n162bar;
  wire n163bar;
  wire n164bar;
  wire n165bar;
  wire n166bar;
  wire n167bar;
  wire n168bar;
  wire n169bar;
  wire n170bar;
  wire n171bar;
  wire n172bar;
  wire n173bar;
  wire n174bar;
  wire n175bar;
  wire n176bar;
  wire n177bar;
  wire n178bar;
  wire n179bar;
  wire n180bar;
  wire n181bar;
  wire n182bar;
  wire n183bar;
  wire n184bar;
  wire n185bar;
  wire n186bar;
  wire n187bar;
  wire n188bar;
  wire n189bar;
  wire n190bar;
  wire n191bar;
  wire n192bar;
  wire n193bar;
  wire n194bar;
  wire n195bar;
  wire n196bar;
  wire n197bar;
  wire n198bar;
  wire n199bar;
  wire n200bar;
  wire n201bar;
  wire n202bar;
  wire n203bar;
  wire n204bar;
  wire n205bar;
  wire n206bar;
  wire n207bar;
  wire n208bar;
  wire n209bar;
  wire n210bar;
  wire n211bar;
  wire n212bar;
  wire n213bar;
  wire n214bar;
  wire n215bar;
  wire n216bar;
  wire n217bar;
  wire n218bar;
  wire n219bar;
  wire n220bar;
  wire n221bar;
  wire n222bar;
  wire n223bar;
  wire n224bar;
//wire_done

 //assign_done

  assign n224bar = n175;
  assign n224 = n175bar;
  assign n223bar = a[7];
  assign n223 = abar[7];
  assign n222bar = n167;
  assign n222 = n167bar;
  assign n221bar = a[6];
  assign n221 = abar[6];
  assign n220bar = n159;
  assign n220 = n159bar;
  assign n219bar = a[5];
  assign n219 = abar[5];
  assign n218bar = n151;
  assign n218 = n151bar;
  assign n217bar = a[4];
  assign n217 = abar[4];
  assign n216bar = n143;
  assign n216 = n143bar;
  assign n215bar = a[3];
  assign n215 = abar[3];
  assign n214bar = n135;
  assign n214 = n135bar;
  assign n213bar = a[2];
  assign n213 = abar[2];
  assign n212bar = n127;
  assign n212 = n127bar;
  assign n211bar = a[1];
  assign n211 = abar[1];
  assign n210bar = n119;
  assign n210 = n119bar;
  assign n209bar = a[0];
  assign n209 = abar[0];
  assign n208bar = b[7];
  assign n208 = bbar[7];
  assign n207bar = b[6];
  assign n207 = bbar[6];
  assign n206bar = b[5];
  assign n206 = bbar[5];
  assign n205bar = b[4];
  assign n205 = bbar[4];
  assign n204bar = b[3];
  assign n204 = bbar[3];
  assign n203bar = b[2];
  assign n203 = bbar[2];
  assign n202bar = b[1];
  assign n202 = bbar[1];
  assign n201bar = b[0];
  assign n201 = bbar[0];
  assign n200bar = n171;
  assign n200 = n171bar;
  assign n199bar = c[7];
  assign n199 = cbar[7];
  assign n198bar = n163;
  assign n198 = n163bar;
  assign n197bar = c[6];
  assign n197 = cbar[6];
  assign n196bar = n155;
  assign n196 = n155bar;
  assign n195bar = c[5];
  assign n195 = cbar[5];
  assign n194bar = n147;
  assign n194 = n147bar;
  assign n193bar = c[4];
  assign n193 = cbar[4];
  assign n192bar = n139;
  assign n192 = n139bar;
  assign n191bar = c[3];
  assign n191 = cbar[3];
  assign n190bar = n131;
  assign n190 = n131bar;
  assign n189bar = c[2];
  assign n189 = cbar[2];
  assign n188bar = n123;
  assign n188 = n123bar;
  assign n187bar = c[1];
  assign n187 = cbar[1];
  assign n186bar = n115;
  assign n186 = n115bar;
  assign n185bar = c[0];
  assign n185 = cbar[0];
  assign n184bar = d[7];
  assign n184 = dbar[7];
  assign n183bar = d[6];
  assign n183 = dbar[6];
  assign n182bar = d[5];
  assign n182 = dbar[5];
  assign n181bar = d[4];
  assign n181 = dbar[4];
  assign n180bar = d[3];
  assign n180 = dbar[3];
  assign n179bar = d[2];
  assign n179 = dbar[2];
  assign n178bar = d[1];
  assign n178 = dbar[1];
  assign n177bar = d[0];
  assign n177 = dbar[0];
  OR2_X1 U49 ( .A1(n176), .A2(n224), .ZN(y[7]) );
  AND2_X1 U49bar ( .A1(n176bar), .A2(n224bar), .ZN(ybar[7]) );
  OR2_X1 U50 ( .A1(n174), .A2(n200), .ZN(n175) );
  AND2_X1 U50bar ( .A1(n174bar), .A2(n200bar), .ZN(n175bar) );
  AND2_X1 U51 ( .A1(n200), .A2(n174), .ZN(n176) );
  OR2_X1 U51bar ( .A1(n200bar), .A2(n174bar), .ZN(n176bar) );
  AND2_X1 U52 ( .A1(n173), .A2(n172), .ZN(n174) );
  OR2_X1 U52bar ( .A1(n173bar), .A2(n172bar), .ZN(n174bar) );
  OR2_X1 U53 ( .A1(n223), .A2(b[7]), .ZN(n172) );
  AND2_X1 U53bar ( .A1(n223bar), .A2(bbar[7]), .ZN(n172bar) );
  OR2_X1 U54 ( .A1(n208), .A2(a[7]), .ZN(n173) );
  AND2_X1 U54bar ( .A1(n208bar), .A2(abar[7]), .ZN(n173bar) );
  AND2_X1 U55 ( .A1(n170), .A2(n169), .ZN(n171) );
  OR2_X1 U55bar ( .A1(n170bar), .A2(n169bar), .ZN(n171bar) );
  OR2_X1 U56 ( .A1(n199), .A2(d[7]), .ZN(n169) );
  AND2_X1 U56bar ( .A1(n199bar), .A2(dbar[7]), .ZN(n169bar) );
  OR2_X1 U57 ( .A1(n184), .A2(c[7]), .ZN(n170) );
  AND2_X1 U57bar ( .A1(n184bar), .A2(cbar[7]), .ZN(n170bar) );
  OR2_X1 U58 ( .A1(n168), .A2(n222), .ZN(y[6]) );
  AND2_X1 U58bar ( .A1(n168bar), .A2(n222bar), .ZN(ybar[6]) );
  OR2_X1 U59 ( .A1(n166), .A2(n198), .ZN(n167) );
  AND2_X1 U59bar ( .A1(n166bar), .A2(n198bar), .ZN(n167bar) );
  AND2_X1 U60 ( .A1(n198), .A2(n166), .ZN(n168) );
  OR2_X1 U60bar ( .A1(n198bar), .A2(n166bar), .ZN(n168bar) );
  AND2_X1 U61 ( .A1(n165), .A2(n164), .ZN(n166) );
  OR2_X1 U61bar ( .A1(n165bar), .A2(n164bar), .ZN(n166bar) );
  OR2_X1 U62 ( .A1(n221), .A2(b[6]), .ZN(n164) );
  AND2_X1 U62bar ( .A1(n221bar), .A2(bbar[6]), .ZN(n164bar) );
  OR2_X1 U63 ( .A1(n207), .A2(a[6]), .ZN(n165) );
  AND2_X1 U63bar ( .A1(n207bar), .A2(abar[6]), .ZN(n165bar) );
  AND2_X1 U64 ( .A1(n162), .A2(n161), .ZN(n163) );
  OR2_X1 U64bar ( .A1(n162bar), .A2(n161bar), .ZN(n163bar) );
  OR2_X1 U65 ( .A1(n197), .A2(d[6]), .ZN(n161) );
  AND2_X1 U65bar ( .A1(n197bar), .A2(dbar[6]), .ZN(n161bar) );
  OR2_X1 U66 ( .A1(n183), .A2(c[6]), .ZN(n162) );
  AND2_X1 U66bar ( .A1(n183bar), .A2(cbar[6]), .ZN(n162bar) );
  OR2_X1 U67 ( .A1(n160), .A2(n220), .ZN(y[5]) );
  AND2_X1 U67bar ( .A1(n160bar), .A2(n220bar), .ZN(ybar[5]) );
  OR2_X1 U68 ( .A1(n158), .A2(n196), .ZN(n159) );
  AND2_X1 U68bar ( .A1(n158bar), .A2(n196bar), .ZN(n159bar) );
  AND2_X1 U69 ( .A1(n196), .A2(n158), .ZN(n160) );
  OR2_X1 U69bar ( .A1(n196bar), .A2(n158bar), .ZN(n160bar) );
  AND2_X1 U70 ( .A1(n157), .A2(n156), .ZN(n158) );
  OR2_X1 U70bar ( .A1(n157bar), .A2(n156bar), .ZN(n158bar) );
  OR2_X1 U71 ( .A1(n219), .A2(b[5]), .ZN(n156) );
  AND2_X1 U71bar ( .A1(n219bar), .A2(bbar[5]), .ZN(n156bar) );
  OR2_X1 U72 ( .A1(n206), .A2(a[5]), .ZN(n157) );
  AND2_X1 U72bar ( .A1(n206bar), .A2(abar[5]), .ZN(n157bar) );
  AND2_X1 U73 ( .A1(n154), .A2(n153), .ZN(n155) );
  OR2_X1 U73bar ( .A1(n154bar), .A2(n153bar), .ZN(n155bar) );
  OR2_X1 U74 ( .A1(n195), .A2(d[5]), .ZN(n153) );
  AND2_X1 U74bar ( .A1(n195bar), .A2(dbar[5]), .ZN(n153bar) );
  OR2_X1 U75 ( .A1(n182), .A2(c[5]), .ZN(n154) );
  AND2_X1 U75bar ( .A1(n182bar), .A2(cbar[5]), .ZN(n154bar) );
  OR2_X1 U76 ( .A1(n152), .A2(n218), .ZN(y[4]) );
  AND2_X1 U76bar ( .A1(n152bar), .A2(n218bar), .ZN(ybar[4]) );
  OR2_X1 U77 ( .A1(n150), .A2(n194), .ZN(n151) );
  AND2_X1 U77bar ( .A1(n150bar), .A2(n194bar), .ZN(n151bar) );
  AND2_X1 U78 ( .A1(n194), .A2(n150), .ZN(n152) );
  OR2_X1 U78bar ( .A1(n194bar), .A2(n150bar), .ZN(n152bar) );
  AND2_X1 U79 ( .A1(n149), .A2(n148), .ZN(n150) );
  OR2_X1 U79bar ( .A1(n149bar), .A2(n148bar), .ZN(n150bar) );
  OR2_X1 U80 ( .A1(n217), .A2(b[4]), .ZN(n148) );
  AND2_X1 U80bar ( .A1(n217bar), .A2(bbar[4]), .ZN(n148bar) );
  OR2_X1 U81 ( .A1(n205), .A2(a[4]), .ZN(n149) );
  AND2_X1 U81bar ( .A1(n205bar), .A2(abar[4]), .ZN(n149bar) );
  AND2_X1 U82 ( .A1(n146), .A2(n145), .ZN(n147) );
  OR2_X1 U82bar ( .A1(n146bar), .A2(n145bar), .ZN(n147bar) );
  OR2_X1 U83 ( .A1(n193), .A2(d[4]), .ZN(n145) );
  AND2_X1 U83bar ( .A1(n193bar), .A2(dbar[4]), .ZN(n145bar) );
  OR2_X1 U84 ( .A1(n181), .A2(c[4]), .ZN(n146) );
  AND2_X1 U84bar ( .A1(n181bar), .A2(cbar[4]), .ZN(n146bar) );
  OR2_X1 U85 ( .A1(n144), .A2(n216), .ZN(y[3]) );
  AND2_X1 U85bar ( .A1(n144bar), .A2(n216bar), .ZN(ybar[3]) );
  OR2_X1 U86 ( .A1(n142), .A2(n192), .ZN(n143) );
  AND2_X1 U86bar ( .A1(n142bar), .A2(n192bar), .ZN(n143bar) );
  AND2_X1 U87 ( .A1(n192), .A2(n142), .ZN(n144) );
  OR2_X1 U87bar ( .A1(n192bar), .A2(n142bar), .ZN(n144bar) );
  AND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(n142) );
  OR2_X1 U88bar ( .A1(n141bar), .A2(n140bar), .ZN(n142bar) );
  OR2_X1 U89 ( .A1(n215), .A2(b[3]), .ZN(n140) );
  AND2_X1 U89bar ( .A1(n215bar), .A2(bbar[3]), .ZN(n140bar) );
  OR2_X1 U90 ( .A1(n204), .A2(a[3]), .ZN(n141) );
  AND2_X1 U90bar ( .A1(n204bar), .A2(abar[3]), .ZN(n141bar) );
  AND2_X1 U91 ( .A1(n138), .A2(n137), .ZN(n139) );
  OR2_X1 U91bar ( .A1(n138bar), .A2(n137bar), .ZN(n139bar) );
  OR2_X1 U92 ( .A1(n191), .A2(d[3]), .ZN(n137) );
  AND2_X1 U92bar ( .A1(n191bar), .A2(dbar[3]), .ZN(n137bar) );
  OR2_X1 U93 ( .A1(n180), .A2(c[3]), .ZN(n138) );
  AND2_X1 U93bar ( .A1(n180bar), .A2(cbar[3]), .ZN(n138bar) );
  OR2_X1 U94 ( .A1(n136), .A2(n214), .ZN(y[2]) );
  AND2_X1 U94bar ( .A1(n136bar), .A2(n214bar), .ZN(ybar[2]) );
  OR2_X1 U95 ( .A1(n134), .A2(n190), .ZN(n135) );
  AND2_X1 U95bar ( .A1(n134bar), .A2(n190bar), .ZN(n135bar) );
  AND2_X1 U96 ( .A1(n190), .A2(n134), .ZN(n136) );
  OR2_X1 U96bar ( .A1(n190bar), .A2(n134bar), .ZN(n136bar) );
  AND2_X1 U97 ( .A1(n133), .A2(n132), .ZN(n134) );
  OR2_X1 U97bar ( .A1(n133bar), .A2(n132bar), .ZN(n134bar) );
  OR2_X1 U98 ( .A1(n213), .A2(b[2]), .ZN(n132) );
  AND2_X1 U98bar ( .A1(n213bar), .A2(bbar[2]), .ZN(n132bar) );
  OR2_X1 U99 ( .A1(n203), .A2(a[2]), .ZN(n133) );
  AND2_X1 U99bar ( .A1(n203bar), .A2(abar[2]), .ZN(n133bar) );
  AND2_X1 U100 ( .A1(n130), .A2(n129), .ZN(n131) );
  OR2_X1 U100bar ( .A1(n130bar), .A2(n129bar), .ZN(n131bar) );
  OR2_X1 U101 ( .A1(n189), .A2(d[2]), .ZN(n129) );
  AND2_X1 U101bar ( .A1(n189bar), .A2(dbar[2]), .ZN(n129bar) );
  OR2_X1 U102 ( .A1(n179), .A2(c[2]), .ZN(n130) );
  AND2_X1 U102bar ( .A1(n179bar), .A2(cbar[2]), .ZN(n130bar) );
  OR2_X1 U103 ( .A1(n128), .A2(n212), .ZN(y[1]) );
  AND2_X1 U103bar ( .A1(n128bar), .A2(n212bar), .ZN(ybar[1]) );
  OR2_X1 U104 ( .A1(n126), .A2(n188), .ZN(n127) );
  AND2_X1 U104bar ( .A1(n126bar), .A2(n188bar), .ZN(n127bar) );
  AND2_X1 U105 ( .A1(n188), .A2(n126), .ZN(n128) );
  OR2_X1 U105bar ( .A1(n188bar), .A2(n126bar), .ZN(n128bar) );
  AND2_X1 U106 ( .A1(n125), .A2(n124), .ZN(n126) );
  OR2_X1 U106bar ( .A1(n125bar), .A2(n124bar), .ZN(n126bar) );
  OR2_X1 U107 ( .A1(n211), .A2(b[1]), .ZN(n124) );
  AND2_X1 U107bar ( .A1(n211bar), .A2(bbar[1]), .ZN(n124bar) );
  OR2_X1 U108 ( .A1(n202), .A2(a[1]), .ZN(n125) );
  AND2_X1 U108bar ( .A1(n202bar), .A2(abar[1]), .ZN(n125bar) );
  AND2_X1 U109 ( .A1(n122), .A2(n121), .ZN(n123) );
  OR2_X1 U109bar ( .A1(n122bar), .A2(n121bar), .ZN(n123bar) );
  OR2_X1 U110 ( .A1(n187), .A2(d[1]), .ZN(n121) );
  AND2_X1 U110bar ( .A1(n187bar), .A2(dbar[1]), .ZN(n121bar) );
  OR2_X1 U111 ( .A1(n178), .A2(c[1]), .ZN(n122) );
  AND2_X1 U111bar ( .A1(n178bar), .A2(cbar[1]), .ZN(n122bar) );
  OR2_X1 U112 ( .A1(n120), .A2(n210), .ZN(y[0]) );
  AND2_X1 U112bar ( .A1(n120bar), .A2(n210bar), .ZN(ybar[0]) );
  OR2_X1 U113 ( .A1(n118), .A2(n186), .ZN(n119) );
  AND2_X1 U113bar ( .A1(n118bar), .A2(n186bar), .ZN(n119bar) );
  AND2_X1 U114 ( .A1(n186), .A2(n118), .ZN(n120) );
  OR2_X1 U114bar ( .A1(n186bar), .A2(n118bar), .ZN(n120bar) );
  AND2_X1 U115 ( .A1(n117), .A2(n116), .ZN(n118) );
  OR2_X1 U115bar ( .A1(n117bar), .A2(n116bar), .ZN(n118bar) );
  OR2_X1 U116 ( .A1(n209), .A2(b[0]), .ZN(n116) );
  AND2_X1 U116bar ( .A1(n209bar), .A2(bbar[0]), .ZN(n116bar) );
  OR2_X1 U117 ( .A1(n201), .A2(a[0]), .ZN(n117) );
  AND2_X1 U117bar ( .A1(n201bar), .A2(abar[0]), .ZN(n117bar) );
  AND2_X1 U118 ( .A1(n114), .A2(n113), .ZN(n115) );
  OR2_X1 U118bar ( .A1(n114bar), .A2(n113bar), .ZN(n115bar) );
  OR2_X1 U119 ( .A1(n185), .A2(d[0]), .ZN(n113) );
  AND2_X1 U119bar ( .A1(n185bar), .A2(dbar[0]), .ZN(n113bar) );
  OR2_X1 U120 ( .A1(n177), .A2(c[0]), .ZN(n114) );
  AND2_X1 U120bar ( .A1(n177bar), .A2(cbar[0]), .ZN(n114bar) );
endmodule

module byteXor4_15 ( a, b, c, d, y );

  input wire [7:0] a;
  input wire [7:0] b;
  input wire [7:0] c;
  input wire [7:0] d;
  wire [7:0] abar;
  wire [7:0] bbar;
  wire [7:0] cbar;
  wire [7:0] dbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign cbar[0] = ~c[0];
  assign cbar[1] = ~c[1];
  assign cbar[2] = ~c[2];
  assign cbar[3] = ~c[3];
  assign cbar[4] = ~c[4];
  assign cbar[5] = ~c[5];
  assign cbar[6] = ~c[6];
  assign cbar[7] = ~c[7];
  assign dbar[0] = ~d[0];
  assign dbar[1] = ~d[1];
  assign dbar[2] = ~d[2];
  assign dbar[3] = ~d[3];
  assign dbar[4] = ~d[4];
  assign dbar[5] = ~d[5];
  assign dbar[6] = ~d[6];
  assign dbar[7] = ~d[7];
//input_done

  output wire [7:0] y;
  wire [7:0] ybar;
//output_done

  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n113bar;
  wire n114bar;
  wire n115bar;
  wire n116bar;
  wire n117bar;
  wire n118bar;
  wire n119bar;
  wire n120bar;
  wire n121bar;
  wire n122bar;
  wire n123bar;
  wire n124bar;
  wire n125bar;
  wire n126bar;
  wire n127bar;
  wire n128bar;
  wire n129bar;
  wire n130bar;
  wire n131bar;
  wire n132bar;
  wire n133bar;
  wire n134bar;
  wire n135bar;
  wire n136bar;
  wire n137bar;
  wire n138bar;
  wire n139bar;
  wire n140bar;
  wire n141bar;
  wire n142bar;
  wire n143bar;
  wire n144bar;
  wire n145bar;
  wire n146bar;
  wire n147bar;
  wire n148bar;
  wire n149bar;
  wire n150bar;
  wire n151bar;
  wire n152bar;
  wire n153bar;
  wire n154bar;
  wire n155bar;
  wire n156bar;
  wire n157bar;
  wire n158bar;
  wire n159bar;
  wire n160bar;
  wire n161bar;
  wire n162bar;
  wire n163bar;
  wire n164bar;
  wire n165bar;
  wire n166bar;
  wire n167bar;
  wire n168bar;
  wire n169bar;
  wire n170bar;
  wire n171bar;
  wire n172bar;
  wire n173bar;
  wire n174bar;
  wire n175bar;
  wire n176bar;
  wire n177bar;
  wire n178bar;
  wire n179bar;
  wire n180bar;
  wire n181bar;
  wire n182bar;
  wire n183bar;
  wire n184bar;
  wire n185bar;
  wire n186bar;
  wire n187bar;
  wire n188bar;
  wire n189bar;
  wire n190bar;
  wire n191bar;
  wire n192bar;
  wire n193bar;
  wire n194bar;
  wire n195bar;
  wire n196bar;
  wire n197bar;
  wire n198bar;
  wire n199bar;
  wire n200bar;
  wire n201bar;
  wire n202bar;
  wire n203bar;
  wire n204bar;
  wire n205bar;
  wire n206bar;
  wire n207bar;
  wire n208bar;
  wire n209bar;
  wire n210bar;
  wire n211bar;
  wire n212bar;
  wire n213bar;
  wire n214bar;
  wire n215bar;
  wire n216bar;
  wire n217bar;
  wire n218bar;
  wire n219bar;
  wire n220bar;
  wire n221bar;
  wire n222bar;
  wire n223bar;
  wire n224bar;
//wire_done

 //assign_done

  assign n224bar = n175;
  assign n224 = n175bar;
  assign n223bar = a[7];
  assign n223 = abar[7];
  assign n222bar = n167;
  assign n222 = n167bar;
  assign n221bar = a[6];
  assign n221 = abar[6];
  assign n220bar = n159;
  assign n220 = n159bar;
  assign n219bar = a[5];
  assign n219 = abar[5];
  assign n218bar = n151;
  assign n218 = n151bar;
  assign n217bar = a[4];
  assign n217 = abar[4];
  assign n216bar = n143;
  assign n216 = n143bar;
  assign n215bar = a[3];
  assign n215 = abar[3];
  assign n214bar = n135;
  assign n214 = n135bar;
  assign n213bar = a[2];
  assign n213 = abar[2];
  assign n212bar = n127;
  assign n212 = n127bar;
  assign n211bar = a[1];
  assign n211 = abar[1];
  assign n210bar = n119;
  assign n210 = n119bar;
  assign n209bar = a[0];
  assign n209 = abar[0];
  assign n208bar = b[7];
  assign n208 = bbar[7];
  assign n207bar = b[6];
  assign n207 = bbar[6];
  assign n206bar = b[5];
  assign n206 = bbar[5];
  assign n205bar = b[4];
  assign n205 = bbar[4];
  assign n204bar = b[3];
  assign n204 = bbar[3];
  assign n203bar = b[2];
  assign n203 = bbar[2];
  assign n202bar = b[1];
  assign n202 = bbar[1];
  assign n201bar = b[0];
  assign n201 = bbar[0];
  assign n200bar = n171;
  assign n200 = n171bar;
  assign n199bar = c[7];
  assign n199 = cbar[7];
  assign n198bar = n163;
  assign n198 = n163bar;
  assign n197bar = c[6];
  assign n197 = cbar[6];
  assign n196bar = n155;
  assign n196 = n155bar;
  assign n195bar = c[5];
  assign n195 = cbar[5];
  assign n194bar = n147;
  assign n194 = n147bar;
  assign n193bar = c[4];
  assign n193 = cbar[4];
  assign n192bar = n139;
  assign n192 = n139bar;
  assign n191bar = c[3];
  assign n191 = cbar[3];
  assign n190bar = n131;
  assign n190 = n131bar;
  assign n189bar = c[2];
  assign n189 = cbar[2];
  assign n188bar = n123;
  assign n188 = n123bar;
  assign n187bar = c[1];
  assign n187 = cbar[1];
  assign n186bar = n115;
  assign n186 = n115bar;
  assign n185bar = c[0];
  assign n185 = cbar[0];
  assign n184bar = d[7];
  assign n184 = dbar[7];
  assign n183bar = d[6];
  assign n183 = dbar[6];
  assign n182bar = d[5];
  assign n182 = dbar[5];
  assign n181bar = d[4];
  assign n181 = dbar[4];
  assign n180bar = d[3];
  assign n180 = dbar[3];
  assign n179bar = d[2];
  assign n179 = dbar[2];
  assign n178bar = d[1];
  assign n178 = dbar[1];
  assign n177bar = d[0];
  assign n177 = dbar[0];
  OR2_X1 U49 ( .A1(n176), .A2(n224), .ZN(y[7]) );
  AND2_X1 U49bar ( .A1(n176bar), .A2(n224bar), .ZN(ybar[7]) );
  OR2_X1 U50 ( .A1(n174), .A2(n200), .ZN(n175) );
  AND2_X1 U50bar ( .A1(n174bar), .A2(n200bar), .ZN(n175bar) );
  AND2_X1 U51 ( .A1(n200), .A2(n174), .ZN(n176) );
  OR2_X1 U51bar ( .A1(n200bar), .A2(n174bar), .ZN(n176bar) );
  AND2_X1 U52 ( .A1(n173), .A2(n172), .ZN(n174) );
  OR2_X1 U52bar ( .A1(n173bar), .A2(n172bar), .ZN(n174bar) );
  OR2_X1 U53 ( .A1(n223), .A2(b[7]), .ZN(n172) );
  AND2_X1 U53bar ( .A1(n223bar), .A2(bbar[7]), .ZN(n172bar) );
  OR2_X1 U54 ( .A1(n208), .A2(a[7]), .ZN(n173) );
  AND2_X1 U54bar ( .A1(n208bar), .A2(abar[7]), .ZN(n173bar) );
  AND2_X1 U55 ( .A1(n170), .A2(n169), .ZN(n171) );
  OR2_X1 U55bar ( .A1(n170bar), .A2(n169bar), .ZN(n171bar) );
  OR2_X1 U56 ( .A1(n199), .A2(d[7]), .ZN(n169) );
  AND2_X1 U56bar ( .A1(n199bar), .A2(dbar[7]), .ZN(n169bar) );
  OR2_X1 U57 ( .A1(n184), .A2(c[7]), .ZN(n170) );
  AND2_X1 U57bar ( .A1(n184bar), .A2(cbar[7]), .ZN(n170bar) );
  OR2_X1 U58 ( .A1(n168), .A2(n222), .ZN(y[6]) );
  AND2_X1 U58bar ( .A1(n168bar), .A2(n222bar), .ZN(ybar[6]) );
  OR2_X1 U59 ( .A1(n166), .A2(n198), .ZN(n167) );
  AND2_X1 U59bar ( .A1(n166bar), .A2(n198bar), .ZN(n167bar) );
  AND2_X1 U60 ( .A1(n198), .A2(n166), .ZN(n168) );
  OR2_X1 U60bar ( .A1(n198bar), .A2(n166bar), .ZN(n168bar) );
  AND2_X1 U61 ( .A1(n165), .A2(n164), .ZN(n166) );
  OR2_X1 U61bar ( .A1(n165bar), .A2(n164bar), .ZN(n166bar) );
  OR2_X1 U62 ( .A1(n221), .A2(b[6]), .ZN(n164) );
  AND2_X1 U62bar ( .A1(n221bar), .A2(bbar[6]), .ZN(n164bar) );
  OR2_X1 U63 ( .A1(n207), .A2(a[6]), .ZN(n165) );
  AND2_X1 U63bar ( .A1(n207bar), .A2(abar[6]), .ZN(n165bar) );
  AND2_X1 U64 ( .A1(n162), .A2(n161), .ZN(n163) );
  OR2_X1 U64bar ( .A1(n162bar), .A2(n161bar), .ZN(n163bar) );
  OR2_X1 U65 ( .A1(n197), .A2(d[6]), .ZN(n161) );
  AND2_X1 U65bar ( .A1(n197bar), .A2(dbar[6]), .ZN(n161bar) );
  OR2_X1 U66 ( .A1(n183), .A2(c[6]), .ZN(n162) );
  AND2_X1 U66bar ( .A1(n183bar), .A2(cbar[6]), .ZN(n162bar) );
  OR2_X1 U67 ( .A1(n160), .A2(n220), .ZN(y[5]) );
  AND2_X1 U67bar ( .A1(n160bar), .A2(n220bar), .ZN(ybar[5]) );
  OR2_X1 U68 ( .A1(n158), .A2(n196), .ZN(n159) );
  AND2_X1 U68bar ( .A1(n158bar), .A2(n196bar), .ZN(n159bar) );
  AND2_X1 U69 ( .A1(n196), .A2(n158), .ZN(n160) );
  OR2_X1 U69bar ( .A1(n196bar), .A2(n158bar), .ZN(n160bar) );
  AND2_X1 U70 ( .A1(n157), .A2(n156), .ZN(n158) );
  OR2_X1 U70bar ( .A1(n157bar), .A2(n156bar), .ZN(n158bar) );
  OR2_X1 U71 ( .A1(n219), .A2(b[5]), .ZN(n156) );
  AND2_X1 U71bar ( .A1(n219bar), .A2(bbar[5]), .ZN(n156bar) );
  OR2_X1 U72 ( .A1(n206), .A2(a[5]), .ZN(n157) );
  AND2_X1 U72bar ( .A1(n206bar), .A2(abar[5]), .ZN(n157bar) );
  AND2_X1 U73 ( .A1(n154), .A2(n153), .ZN(n155) );
  OR2_X1 U73bar ( .A1(n154bar), .A2(n153bar), .ZN(n155bar) );
  OR2_X1 U74 ( .A1(n195), .A2(d[5]), .ZN(n153) );
  AND2_X1 U74bar ( .A1(n195bar), .A2(dbar[5]), .ZN(n153bar) );
  OR2_X1 U75 ( .A1(n182), .A2(c[5]), .ZN(n154) );
  AND2_X1 U75bar ( .A1(n182bar), .A2(cbar[5]), .ZN(n154bar) );
  OR2_X1 U76 ( .A1(n152), .A2(n218), .ZN(y[4]) );
  AND2_X1 U76bar ( .A1(n152bar), .A2(n218bar), .ZN(ybar[4]) );
  OR2_X1 U77 ( .A1(n150), .A2(n194), .ZN(n151) );
  AND2_X1 U77bar ( .A1(n150bar), .A2(n194bar), .ZN(n151bar) );
  AND2_X1 U78 ( .A1(n194), .A2(n150), .ZN(n152) );
  OR2_X1 U78bar ( .A1(n194bar), .A2(n150bar), .ZN(n152bar) );
  AND2_X1 U79 ( .A1(n149), .A2(n148), .ZN(n150) );
  OR2_X1 U79bar ( .A1(n149bar), .A2(n148bar), .ZN(n150bar) );
  OR2_X1 U80 ( .A1(n217), .A2(b[4]), .ZN(n148) );
  AND2_X1 U80bar ( .A1(n217bar), .A2(bbar[4]), .ZN(n148bar) );
  OR2_X1 U81 ( .A1(n205), .A2(a[4]), .ZN(n149) );
  AND2_X1 U81bar ( .A1(n205bar), .A2(abar[4]), .ZN(n149bar) );
  AND2_X1 U82 ( .A1(n146), .A2(n145), .ZN(n147) );
  OR2_X1 U82bar ( .A1(n146bar), .A2(n145bar), .ZN(n147bar) );
  OR2_X1 U83 ( .A1(n193), .A2(d[4]), .ZN(n145) );
  AND2_X1 U83bar ( .A1(n193bar), .A2(dbar[4]), .ZN(n145bar) );
  OR2_X1 U84 ( .A1(n181), .A2(c[4]), .ZN(n146) );
  AND2_X1 U84bar ( .A1(n181bar), .A2(cbar[4]), .ZN(n146bar) );
  OR2_X1 U85 ( .A1(n144), .A2(n216), .ZN(y[3]) );
  AND2_X1 U85bar ( .A1(n144bar), .A2(n216bar), .ZN(ybar[3]) );
  OR2_X1 U86 ( .A1(n142), .A2(n192), .ZN(n143) );
  AND2_X1 U86bar ( .A1(n142bar), .A2(n192bar), .ZN(n143bar) );
  AND2_X1 U87 ( .A1(n192), .A2(n142), .ZN(n144) );
  OR2_X1 U87bar ( .A1(n192bar), .A2(n142bar), .ZN(n144bar) );
  AND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(n142) );
  OR2_X1 U88bar ( .A1(n141bar), .A2(n140bar), .ZN(n142bar) );
  OR2_X1 U89 ( .A1(n215), .A2(b[3]), .ZN(n140) );
  AND2_X1 U89bar ( .A1(n215bar), .A2(bbar[3]), .ZN(n140bar) );
  OR2_X1 U90 ( .A1(n204), .A2(a[3]), .ZN(n141) );
  AND2_X1 U90bar ( .A1(n204bar), .A2(abar[3]), .ZN(n141bar) );
  AND2_X1 U91 ( .A1(n138), .A2(n137), .ZN(n139) );
  OR2_X1 U91bar ( .A1(n138bar), .A2(n137bar), .ZN(n139bar) );
  OR2_X1 U92 ( .A1(n191), .A2(d[3]), .ZN(n137) );
  AND2_X1 U92bar ( .A1(n191bar), .A2(dbar[3]), .ZN(n137bar) );
  OR2_X1 U93 ( .A1(n180), .A2(c[3]), .ZN(n138) );
  AND2_X1 U93bar ( .A1(n180bar), .A2(cbar[3]), .ZN(n138bar) );
  OR2_X1 U94 ( .A1(n136), .A2(n214), .ZN(y[2]) );
  AND2_X1 U94bar ( .A1(n136bar), .A2(n214bar), .ZN(ybar[2]) );
  OR2_X1 U95 ( .A1(n134), .A2(n190), .ZN(n135) );
  AND2_X1 U95bar ( .A1(n134bar), .A2(n190bar), .ZN(n135bar) );
  AND2_X1 U96 ( .A1(n190), .A2(n134), .ZN(n136) );
  OR2_X1 U96bar ( .A1(n190bar), .A2(n134bar), .ZN(n136bar) );
  AND2_X1 U97 ( .A1(n133), .A2(n132), .ZN(n134) );
  OR2_X1 U97bar ( .A1(n133bar), .A2(n132bar), .ZN(n134bar) );
  OR2_X1 U98 ( .A1(n213), .A2(b[2]), .ZN(n132) );
  AND2_X1 U98bar ( .A1(n213bar), .A2(bbar[2]), .ZN(n132bar) );
  OR2_X1 U99 ( .A1(n203), .A2(a[2]), .ZN(n133) );
  AND2_X1 U99bar ( .A1(n203bar), .A2(abar[2]), .ZN(n133bar) );
  AND2_X1 U100 ( .A1(n130), .A2(n129), .ZN(n131) );
  OR2_X1 U100bar ( .A1(n130bar), .A2(n129bar), .ZN(n131bar) );
  OR2_X1 U101 ( .A1(n189), .A2(d[2]), .ZN(n129) );
  AND2_X1 U101bar ( .A1(n189bar), .A2(dbar[2]), .ZN(n129bar) );
  OR2_X1 U102 ( .A1(n179), .A2(c[2]), .ZN(n130) );
  AND2_X1 U102bar ( .A1(n179bar), .A2(cbar[2]), .ZN(n130bar) );
  OR2_X1 U103 ( .A1(n128), .A2(n212), .ZN(y[1]) );
  AND2_X1 U103bar ( .A1(n128bar), .A2(n212bar), .ZN(ybar[1]) );
  OR2_X1 U104 ( .A1(n126), .A2(n188), .ZN(n127) );
  AND2_X1 U104bar ( .A1(n126bar), .A2(n188bar), .ZN(n127bar) );
  AND2_X1 U105 ( .A1(n188), .A2(n126), .ZN(n128) );
  OR2_X1 U105bar ( .A1(n188bar), .A2(n126bar), .ZN(n128bar) );
  AND2_X1 U106 ( .A1(n125), .A2(n124), .ZN(n126) );
  OR2_X1 U106bar ( .A1(n125bar), .A2(n124bar), .ZN(n126bar) );
  OR2_X1 U107 ( .A1(n211), .A2(b[1]), .ZN(n124) );
  AND2_X1 U107bar ( .A1(n211bar), .A2(bbar[1]), .ZN(n124bar) );
  OR2_X1 U108 ( .A1(n202), .A2(a[1]), .ZN(n125) );
  AND2_X1 U108bar ( .A1(n202bar), .A2(abar[1]), .ZN(n125bar) );
  AND2_X1 U109 ( .A1(n122), .A2(n121), .ZN(n123) );
  OR2_X1 U109bar ( .A1(n122bar), .A2(n121bar), .ZN(n123bar) );
  OR2_X1 U110 ( .A1(n187), .A2(d[1]), .ZN(n121) );
  AND2_X1 U110bar ( .A1(n187bar), .A2(dbar[1]), .ZN(n121bar) );
  OR2_X1 U111 ( .A1(n178), .A2(c[1]), .ZN(n122) );
  AND2_X1 U111bar ( .A1(n178bar), .A2(cbar[1]), .ZN(n122bar) );
  OR2_X1 U112 ( .A1(n120), .A2(n210), .ZN(y[0]) );
  AND2_X1 U112bar ( .A1(n120bar), .A2(n210bar), .ZN(ybar[0]) );
  OR2_X1 U113 ( .A1(n118), .A2(n186), .ZN(n119) );
  AND2_X1 U113bar ( .A1(n118bar), .A2(n186bar), .ZN(n119bar) );
  AND2_X1 U114 ( .A1(n186), .A2(n118), .ZN(n120) );
  OR2_X1 U114bar ( .A1(n186bar), .A2(n118bar), .ZN(n120bar) );
  AND2_X1 U115 ( .A1(n117), .A2(n116), .ZN(n118) );
  OR2_X1 U115bar ( .A1(n117bar), .A2(n116bar), .ZN(n118bar) );
  OR2_X1 U116 ( .A1(n209), .A2(b[0]), .ZN(n116) );
  AND2_X1 U116bar ( .A1(n209bar), .A2(bbar[0]), .ZN(n116bar) );
  OR2_X1 U117 ( .A1(n201), .A2(a[0]), .ZN(n117) );
  AND2_X1 U117bar ( .A1(n201bar), .A2(abar[0]), .ZN(n117bar) );
  AND2_X1 U118 ( .A1(n114), .A2(n113), .ZN(n115) );
  OR2_X1 U118bar ( .A1(n114bar), .A2(n113bar), .ZN(n115bar) );
  OR2_X1 U119 ( .A1(n185), .A2(d[0]), .ZN(n113) );
  AND2_X1 U119bar ( .A1(n185bar), .A2(dbar[0]), .ZN(n113bar) );
  OR2_X1 U120 ( .A1(n177), .A2(c[0]), .ZN(n114) );
  AND2_X1 U120bar ( .A1(n177bar), .A2(cbar[0]), .ZN(n114bar) );
endmodule

module mixCol_0 ( in, out );

  input wire [31:0] in;
//input_done

  output wire [31:0] out;
//output_done

  wire [7:0] b0_s2;
  wire [7:0] b1_s2;
  wire [7:0] b2_s2;
  wire [7:0] b3_s2;
  wire [7:0] b0_s3;
  wire [7:0] b1_s3;
  wire [7:0] b2_s3;
  wire [7:0] b3_s3;
//wire_done

 //assign_done

  scale2_0 b0_scale2 ( .in(in[31:24]), .out(b0_s2) );
  scale2_15 b1_scale2 ( .in(in[23:16]), .out(b1_s2) );
  scale2_14 b2_scale2 ( .in(in[15:8]), .out(b2_s2) );
  scale2_13 b3_scale2 ( .in(in[7:0]), .out(b3_s2) );
  byteXor_0 b0_scale3 ( .a(in[31:24]), .b(b0_s2), .y(b0_s3) );
  byteXor_16 b1_scale3 ( .a(in[23:16]), .b(b1_s2), .y(b1_s3) );
  byteXor_15 b2_scale3 ( .a(in[15:8]), .b(b2_s2), .y(b2_s3) );
  byteXor_14 b3_scale3 ( .a(in[7:0]), .b(b3_s2), .y(b3_s3) );
  byteXor4_0 out0 ( .a(b0_s2), .b(b1_s3), .c(in[15:8]), .d(in[7:0]), .y(
        out[31:24]) );
  byteXor4_15 out1 ( .a(in[31:24]), .b(b1_s2), .c(b2_s3), .d(in[7:0]), .y(
        out[23:16]) );
  byteXor4_14 out2 ( .a(in[31:24]), .b(in[23:16]), .c(b2_s2), .d(b3_s3), .y(
        out[15:8]) );
  byteXor4_13 out3 ( .a(b0_s3), .b(in[23:16]), .c(in[15:8]), .d(b3_s2), .y(
        out[7:0]) );
endmodule

module scale2_1 ( in, out );

  input wire [7:0] in;
  wire [7:0] inbar;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
//input_done

  output wire [7:0] out;
  wire [7:0] outbar;
//output_done

  wire in_0;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_1;
  wire in_7;
  wire n11;
  wire n12;
  wire n13;
  wire n14;
  wire n15;
  wire n16;
  wire n17;
  wire n18;
  wire n19;
  wire n20;
  wire in_0bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_1bar;
  wire in_7bar;
  wire n11bar;
  wire n12bar;
  wire n13bar;
  wire n14bar;
  wire n15bar;
  wire n16bar;
  wire n17bar;
  wire n18bar;
  wire n19bar;
  wire n20bar;
//wire_done

  assign in_0 = in[0];
  assign out[7] = in_6;
  assign in_6  = in[6];
  assign out[6] = in_5;
  assign in_5  = in[5];
  assign out[5] = in_4;
  assign in_4  = in[4];
  assign out[2] = in_1;
  assign in_1  = in[1];
  assign out[0] = in_7;
  assign in_7  = in[7];
  assign in_0bar = inbar[0];
  assign outbar[7] = in_6bar;
  assign in_6bar = inbar[6];
  assign outbar[6] = in_5bar;
  assign in_5bar = inbar[5];
  assign outbar[5] = in_4bar;
  assign in_4bar = inbar[4];
  assign outbar[2] = in_1bar;
  assign in_1bar = inbar[1];
  assign outbar[0] = in_7bar;
  assign in_7bar = inbar[7];
//assign_done

  assign n20bar = in_7;
  assign n20 = in_7bar;
  assign n19bar = in[3];
  assign n19 = inbar[3];
  assign n18bar = in[2];
  assign n18 = inbar[2];
  assign n17bar = in_0;
  assign n17 = in_0bar;
  OR2_X1 U5 ( .A1(n16), .A2(n15), .ZN(out[4]) );
  AND2_X1 U5bar ( .A1(n16bar), .A2(n15bar), .ZN(outbar[4]) );
  AND2_X1 U6 ( .A1(in[3]), .A2(n20), .ZN(n15) );
  OR2_X1 U6bar ( .A1(inbar[3]), .A2(n20bar), .ZN(n15bar) );
  AND2_X1 U7 ( .A1(in_7), .A2(n19), .ZN(n16) );
  OR2_X1 U7bar ( .A1(in_7bar), .A2(n19bar), .ZN(n16bar) );
  OR2_X1 U8 ( .A1(n14), .A2(n13), .ZN(out[3]) );
  AND2_X1 U8bar ( .A1(n14bar), .A2(n13bar), .ZN(outbar[3]) );
  AND2_X1 U9 ( .A1(in[2]), .A2(n20), .ZN(n13) );
  OR2_X1 U9bar ( .A1(inbar[2]), .A2(n20bar), .ZN(n13bar) );
  AND2_X1 U10 ( .A1(in_7), .A2(n18), .ZN(n14) );
  OR2_X1 U10bar ( .A1(in_7bar), .A2(n18bar), .ZN(n14bar) );
  OR2_X1 U11 ( .A1(n12), .A2(n11), .ZN(out[1]) );
  AND2_X1 U11bar ( .A1(n12bar), .A2(n11bar), .ZN(outbar[1]) );
  AND2_X1 U12 ( .A1(in_0), .A2(n20), .ZN(n11) );
  OR2_X1 U12bar ( .A1(in_0bar), .A2(n20bar), .ZN(n11bar) );
  AND2_X1 U13 ( .A1(in_7), .A2(n17), .ZN(n12) );
  OR2_X1 U13bar ( .A1(in_7bar), .A2(n17bar), .ZN(n12bar) );
endmodule

module scale2_2 ( in, out );

  input wire [7:0] in;
  wire [7:0] inbar;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
//input_done

  output wire [7:0] out;
  wire [7:0] outbar;
//output_done

  wire in_0;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_1;
  wire in_7;
  wire n11;
  wire n12;
  wire n13;
  wire n14;
  wire n15;
  wire n16;
  wire n17;
  wire n18;
  wire n19;
  wire n20;
  wire in_0bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_1bar;
  wire in_7bar;
  wire n11bar;
  wire n12bar;
  wire n13bar;
  wire n14bar;
  wire n15bar;
  wire n16bar;
  wire n17bar;
  wire n18bar;
  wire n19bar;
  wire n20bar;
//wire_done

  assign in_0 = in[0];
  assign out[7] = in_6;
  assign in_6  = in[6];
  assign out[6] = in_5;
  assign in_5  = in[5];
  assign out[5] = in_4;
  assign in_4  = in[4];
  assign out[2] = in_1;
  assign in_1  = in[1];
  assign out[0] = in_7;
  assign in_7  = in[7];
  assign in_0bar = inbar[0];
  assign outbar[7] = in_6bar;
  assign in_6bar = inbar[6];
  assign outbar[6] = in_5bar;
  assign in_5bar = inbar[5];
  assign outbar[5] = in_4bar;
  assign in_4bar = inbar[4];
  assign outbar[2] = in_1bar;
  assign in_1bar = inbar[1];
  assign outbar[0] = in_7bar;
  assign in_7bar = inbar[7];
//assign_done

  assign n20bar = in_7;
  assign n20 = in_7bar;
  assign n19bar = in[3];
  assign n19 = inbar[3];
  assign n18bar = in[2];
  assign n18 = inbar[2];
  assign n17bar = in_0;
  assign n17 = in_0bar;
  OR2_X1 U5 ( .A1(n16), .A2(n15), .ZN(out[4]) );
  AND2_X1 U5bar ( .A1(n16bar), .A2(n15bar), .ZN(outbar[4]) );
  AND2_X1 U6 ( .A1(in[3]), .A2(n20), .ZN(n15) );
  OR2_X1 U6bar ( .A1(inbar[3]), .A2(n20bar), .ZN(n15bar) );
  AND2_X1 U7 ( .A1(in_7), .A2(n19), .ZN(n16) );
  OR2_X1 U7bar ( .A1(in_7bar), .A2(n19bar), .ZN(n16bar) );
  OR2_X1 U8 ( .A1(n14), .A2(n13), .ZN(out[3]) );
  AND2_X1 U8bar ( .A1(n14bar), .A2(n13bar), .ZN(outbar[3]) );
  AND2_X1 U9 ( .A1(in[2]), .A2(n20), .ZN(n13) );
  OR2_X1 U9bar ( .A1(inbar[2]), .A2(n20bar), .ZN(n13bar) );
  AND2_X1 U10 ( .A1(in_7), .A2(n18), .ZN(n14) );
  OR2_X1 U10bar ( .A1(in_7bar), .A2(n18bar), .ZN(n14bar) );
  OR2_X1 U11 ( .A1(n12), .A2(n11), .ZN(out[1]) );
  AND2_X1 U11bar ( .A1(n12bar), .A2(n11bar), .ZN(outbar[1]) );
  AND2_X1 U12 ( .A1(in_0), .A2(n20), .ZN(n11) );
  OR2_X1 U12bar ( .A1(in_0bar), .A2(n20bar), .ZN(n11bar) );
  AND2_X1 U13 ( .A1(in_7), .A2(n17), .ZN(n12) );
  OR2_X1 U13bar ( .A1(in_7bar), .A2(n17bar), .ZN(n12bar) );
endmodule

module scale2_3 ( in, out );

  input wire [7:0] in;
  wire [7:0] inbar;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
//input_done

  output wire [7:0] out;
  wire [7:0] outbar;
//output_done

  wire in_0;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_1;
  wire in_7;
  wire n11;
  wire n12;
  wire n13;
  wire n14;
  wire n15;
  wire n16;
  wire n17;
  wire n18;
  wire n19;
  wire n20;
  wire in_0bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_1bar;
  wire in_7bar;
  wire n11bar;
  wire n12bar;
  wire n13bar;
  wire n14bar;
  wire n15bar;
  wire n16bar;
  wire n17bar;
  wire n18bar;
  wire n19bar;
  wire n20bar;
//wire_done

  assign in_0 = in[0];
  assign out[7] = in_6;
  assign in_6  = in[6];
  assign out[6] = in_5;
  assign in_5  = in[5];
  assign out[5] = in_4;
  assign in_4  = in[4];
  assign out[2] = in_1;
  assign in_1  = in[1];
  assign out[0] = in_7;
  assign in_7  = in[7];
  assign in_0bar = inbar[0];
  assign outbar[7] = in_6bar;
  assign in_6bar = inbar[6];
  assign outbar[6] = in_5bar;
  assign in_5bar = inbar[5];
  assign outbar[5] = in_4bar;
  assign in_4bar = inbar[4];
  assign outbar[2] = in_1bar;
  assign in_1bar = inbar[1];
  assign outbar[0] = in_7bar;
  assign in_7bar = inbar[7];
//assign_done

  assign n20bar = in_7;
  assign n20 = in_7bar;
  assign n19bar = in[3];
  assign n19 = inbar[3];
  assign n18bar = in[2];
  assign n18 = inbar[2];
  assign n17bar = in_0;
  assign n17 = in_0bar;
  OR2_X1 U5 ( .A1(n16), .A2(n15), .ZN(out[4]) );
  AND2_X1 U5bar ( .A1(n16bar), .A2(n15bar), .ZN(outbar[4]) );
  AND2_X1 U6 ( .A1(in[3]), .A2(n20), .ZN(n15) );
  OR2_X1 U6bar ( .A1(inbar[3]), .A2(n20bar), .ZN(n15bar) );
  AND2_X1 U7 ( .A1(in_7), .A2(n19), .ZN(n16) );
  OR2_X1 U7bar ( .A1(in_7bar), .A2(n19bar), .ZN(n16bar) );
  OR2_X1 U8 ( .A1(n14), .A2(n13), .ZN(out[3]) );
  AND2_X1 U8bar ( .A1(n14bar), .A2(n13bar), .ZN(outbar[3]) );
  AND2_X1 U9 ( .A1(in[2]), .A2(n20), .ZN(n13) );
  OR2_X1 U9bar ( .A1(inbar[2]), .A2(n20bar), .ZN(n13bar) );
  AND2_X1 U10 ( .A1(in_7), .A2(n18), .ZN(n14) );
  OR2_X1 U10bar ( .A1(in_7bar), .A2(n18bar), .ZN(n14bar) );
  OR2_X1 U11 ( .A1(n12), .A2(n11), .ZN(out[1]) );
  AND2_X1 U11bar ( .A1(n12bar), .A2(n11bar), .ZN(outbar[1]) );
  AND2_X1 U12 ( .A1(in_0), .A2(n20), .ZN(n11) );
  OR2_X1 U12bar ( .A1(in_0bar), .A2(n20bar), .ZN(n11bar) );
  AND2_X1 U13 ( .A1(in_7), .A2(n17), .ZN(n12) );
  OR2_X1 U13bar ( .A1(in_7bar), .A2(n17bar), .ZN(n12bar) );
endmodule

module scale2_4 ( in, out );

  input wire [7:0] in;
  wire [7:0] inbar;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
//input_done

  output wire [7:0] out;
  wire [7:0] outbar;
//output_done

  wire in_0;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_1;
  wire in_7;
  wire n11;
  wire n12;
  wire n13;
  wire n14;
  wire n15;
  wire n16;
  wire n17;
  wire n18;
  wire n19;
  wire n20;
  wire in_0bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_1bar;
  wire in_7bar;
  wire n11bar;
  wire n12bar;
  wire n13bar;
  wire n14bar;
  wire n15bar;
  wire n16bar;
  wire n17bar;
  wire n18bar;
  wire n19bar;
  wire n20bar;
//wire_done

  assign in_0 = in[0];
  assign out[7] = in_6;
  assign in_6  = in[6];
  assign out[6] = in_5;
  assign in_5  = in[5];
  assign out[5] = in_4;
  assign in_4  = in[4];
  assign out[2] = in_1;
  assign in_1  = in[1];
  assign out[0] = in_7;
  assign in_7  = in[7];
  assign in_0bar = inbar[0];
  assign outbar[7] = in_6bar;
  assign in_6bar = inbar[6];
  assign outbar[6] = in_5bar;
  assign in_5bar = inbar[5];
  assign outbar[5] = in_4bar;
  assign in_4bar = inbar[4];
  assign outbar[2] = in_1bar;
  assign in_1bar = inbar[1];
  assign outbar[0] = in_7bar;
  assign in_7bar = inbar[7];
//assign_done

  assign n20bar = in_7;
  assign n20 = in_7bar;
  assign n19bar = in[3];
  assign n19 = inbar[3];
  assign n18bar = in[2];
  assign n18 = inbar[2];
  assign n17bar = in_0;
  assign n17 = in_0bar;
  OR2_X1 U5 ( .A1(n16), .A2(n15), .ZN(out[4]) );
  AND2_X1 U5bar ( .A1(n16bar), .A2(n15bar), .ZN(outbar[4]) );
  AND2_X1 U6 ( .A1(in[3]), .A2(n20), .ZN(n15) );
  OR2_X1 U6bar ( .A1(inbar[3]), .A2(n20bar), .ZN(n15bar) );
  AND2_X1 U7 ( .A1(in_7), .A2(n19), .ZN(n16) );
  OR2_X1 U7bar ( .A1(in_7bar), .A2(n19bar), .ZN(n16bar) );
  OR2_X1 U8 ( .A1(n14), .A2(n13), .ZN(out[3]) );
  AND2_X1 U8bar ( .A1(n14bar), .A2(n13bar), .ZN(outbar[3]) );
  AND2_X1 U9 ( .A1(in[2]), .A2(n20), .ZN(n13) );
  OR2_X1 U9bar ( .A1(inbar[2]), .A2(n20bar), .ZN(n13bar) );
  AND2_X1 U10 ( .A1(in_7), .A2(n18), .ZN(n14) );
  OR2_X1 U10bar ( .A1(in_7bar), .A2(n18bar), .ZN(n14bar) );
  OR2_X1 U11 ( .A1(n12), .A2(n11), .ZN(out[1]) );
  AND2_X1 U11bar ( .A1(n12bar), .A2(n11bar), .ZN(outbar[1]) );
  AND2_X1 U12 ( .A1(in_0), .A2(n20), .ZN(n11) );
  OR2_X1 U12bar ( .A1(in_0bar), .A2(n20bar), .ZN(n11bar) );
  AND2_X1 U13 ( .A1(in_7), .A2(n17), .ZN(n12) );
  OR2_X1 U13bar ( .A1(in_7bar), .A2(n17bar), .ZN(n12bar) );
endmodule

module byteXor_2 ( a, b, y );

  input wire [7:0] a;
  input wire [7:0] b;
  wire [7:0] abar;
  wire [7:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
//input_done

  output wire [7:0] y;
  wire [7:0] ybar;
//output_done

  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n33bar;
  wire n34bar;
  wire n35bar;
  wire n36bar;
  wire n37bar;
  wire n38bar;
  wire n39bar;
  wire n40bar;
  wire n41bar;
  wire n42bar;
  wire n43bar;
  wire n44bar;
  wire n45bar;
  wire n46bar;
  wire n47bar;
  wire n48bar;
  wire n49bar;
  wire n50bar;
  wire n51bar;
  wire n52bar;
  wire n53bar;
  wire n54bar;
  wire n55bar;
  wire n56bar;
  wire n57bar;
  wire n58bar;
  wire n59bar;
  wire n60bar;
  wire n61bar;
  wire n62bar;
  wire n63bar;
  wire n64bar;
//wire_done

 //assign_done

  assign n64bar = n47;
  assign n64 = n47bar;
  assign n63bar = a[7];
  assign n63 = abar[7];
  assign n62bar = n45;
  assign n62 = n45bar;
  assign n61bar = a[6];
  assign n61 = abar[6];
  assign n60bar = n43;
  assign n60 = n43bar;
  assign n59bar = a[5];
  assign n59 = abar[5];
  assign n58bar = n41;
  assign n58 = n41bar;
  assign n57bar = a[4];
  assign n57 = abar[4];
  assign n56bar = n39;
  assign n56 = n39bar;
  assign n55bar = a[3];
  assign n55 = abar[3];
  assign n54bar = n37;
  assign n54 = n37bar;
  assign n53bar = a[2];
  assign n53 = abar[2];
  assign n52bar = n35;
  assign n52 = n35bar;
  assign n51bar = a[1];
  assign n51 = abar[1];
  assign n50bar = n33;
  assign n50 = n33bar;
  assign n49bar = a[0];
  assign n49 = abar[0];
  OR2_X1 U17 ( .A1(n48), .A2(n64), .ZN(y[7]) );
  AND2_X1 U17bar ( .A1(n48bar), .A2(n64bar), .ZN(ybar[7]) );
  OR2_X1 U18 ( .A1(n63), .A2(b[7]), .ZN(n47) );
  AND2_X1 U18bar ( .A1(n63bar), .A2(bbar[7]), .ZN(n47bar) );
  AND2_X1 U19 ( .A1(b[7]), .A2(n63), .ZN(n48) );
  OR2_X1 U19bar ( .A1(bbar[7]), .A2(n63bar), .ZN(n48bar) );
  OR2_X1 U20 ( .A1(n46), .A2(n62), .ZN(y[6]) );
  AND2_X1 U20bar ( .A1(n46bar), .A2(n62bar), .ZN(ybar[6]) );
  OR2_X1 U21 ( .A1(n61), .A2(b[6]), .ZN(n45) );
  AND2_X1 U21bar ( .A1(n61bar), .A2(bbar[6]), .ZN(n45bar) );
  AND2_X1 U22 ( .A1(b[6]), .A2(n61), .ZN(n46) );
  OR2_X1 U22bar ( .A1(bbar[6]), .A2(n61bar), .ZN(n46bar) );
  OR2_X1 U23 ( .A1(n44), .A2(n60), .ZN(y[5]) );
  AND2_X1 U23bar ( .A1(n44bar), .A2(n60bar), .ZN(ybar[5]) );
  OR2_X1 U24 ( .A1(n59), .A2(b[5]), .ZN(n43) );
  AND2_X1 U24bar ( .A1(n59bar), .A2(bbar[5]), .ZN(n43bar) );
  AND2_X1 U25 ( .A1(b[5]), .A2(n59), .ZN(n44) );
  OR2_X1 U25bar ( .A1(bbar[5]), .A2(n59bar), .ZN(n44bar) );
  OR2_X1 U26 ( .A1(n42), .A2(n58), .ZN(y[4]) );
  AND2_X1 U26bar ( .A1(n42bar), .A2(n58bar), .ZN(ybar[4]) );
  OR2_X1 U27 ( .A1(n57), .A2(b[4]), .ZN(n41) );
  AND2_X1 U27bar ( .A1(n57bar), .A2(bbar[4]), .ZN(n41bar) );
  AND2_X1 U28 ( .A1(b[4]), .A2(n57), .ZN(n42) );
  OR2_X1 U28bar ( .A1(bbar[4]), .A2(n57bar), .ZN(n42bar) );
  OR2_X1 U29 ( .A1(n40), .A2(n56), .ZN(y[3]) );
  AND2_X1 U29bar ( .A1(n40bar), .A2(n56bar), .ZN(ybar[3]) );
  OR2_X1 U30 ( .A1(n55), .A2(b[3]), .ZN(n39) );
  AND2_X1 U30bar ( .A1(n55bar), .A2(bbar[3]), .ZN(n39bar) );
  AND2_X1 U31 ( .A1(b[3]), .A2(n55), .ZN(n40) );
  OR2_X1 U31bar ( .A1(bbar[3]), .A2(n55bar), .ZN(n40bar) );
  OR2_X1 U32 ( .A1(n38), .A2(n54), .ZN(y[2]) );
  AND2_X1 U32bar ( .A1(n38bar), .A2(n54bar), .ZN(ybar[2]) );
  OR2_X1 U33 ( .A1(n53), .A2(b[2]), .ZN(n37) );
  AND2_X1 U33bar ( .A1(n53bar), .A2(bbar[2]), .ZN(n37bar) );
  AND2_X1 U34 ( .A1(b[2]), .A2(n53), .ZN(n38) );
  OR2_X1 U34bar ( .A1(bbar[2]), .A2(n53bar), .ZN(n38bar) );
  OR2_X1 U35 ( .A1(n36), .A2(n52), .ZN(y[1]) );
  AND2_X1 U35bar ( .A1(n36bar), .A2(n52bar), .ZN(ybar[1]) );
  OR2_X1 U36 ( .A1(n51), .A2(b[1]), .ZN(n35) );
  AND2_X1 U36bar ( .A1(n51bar), .A2(bbar[1]), .ZN(n35bar) );
  AND2_X1 U37 ( .A1(b[1]), .A2(n51), .ZN(n36) );
  OR2_X1 U37bar ( .A1(bbar[1]), .A2(n51bar), .ZN(n36bar) );
  OR2_X1 U38 ( .A1(n34), .A2(n50), .ZN(y[0]) );
  AND2_X1 U38bar ( .A1(n34bar), .A2(n50bar), .ZN(ybar[0]) );
  OR2_X1 U39 ( .A1(n49), .A2(b[0]), .ZN(n33) );
  AND2_X1 U39bar ( .A1(n49bar), .A2(bbar[0]), .ZN(n33bar) );
  AND2_X1 U40 ( .A1(b[0]), .A2(n49), .ZN(n34) );
  OR2_X1 U40bar ( .A1(bbar[0]), .A2(n49bar), .ZN(n34bar) );
endmodule

module byteXor_3 ( a, b, y );

  input wire [7:0] a;
  input wire [7:0] b;
  wire [7:0] abar;
  wire [7:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
//input_done

  output wire [7:0] y;
  wire [7:0] ybar;
//output_done

  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n33bar;
  wire n34bar;
  wire n35bar;
  wire n36bar;
  wire n37bar;
  wire n38bar;
  wire n39bar;
  wire n40bar;
  wire n41bar;
  wire n42bar;
  wire n43bar;
  wire n44bar;
  wire n45bar;
  wire n46bar;
  wire n47bar;
  wire n48bar;
  wire n49bar;
  wire n50bar;
  wire n51bar;
  wire n52bar;
  wire n53bar;
  wire n54bar;
  wire n55bar;
  wire n56bar;
  wire n57bar;
  wire n58bar;
  wire n59bar;
  wire n60bar;
  wire n61bar;
  wire n62bar;
  wire n63bar;
  wire n64bar;
//wire_done

 //assign_done

  assign n64bar = n47;
  assign n64 = n47bar;
  assign n63bar = a[7];
  assign n63 = abar[7];
  assign n62bar = n45;
  assign n62 = n45bar;
  assign n61bar = a[6];
  assign n61 = abar[6];
  assign n60bar = n43;
  assign n60 = n43bar;
  assign n59bar = a[5];
  assign n59 = abar[5];
  assign n58bar = n41;
  assign n58 = n41bar;
  assign n57bar = a[4];
  assign n57 = abar[4];
  assign n56bar = n39;
  assign n56 = n39bar;
  assign n55bar = a[3];
  assign n55 = abar[3];
  assign n54bar = n37;
  assign n54 = n37bar;
  assign n53bar = a[2];
  assign n53 = abar[2];
  assign n52bar = n35;
  assign n52 = n35bar;
  assign n51bar = a[1];
  assign n51 = abar[1];
  assign n50bar = n33;
  assign n50 = n33bar;
  assign n49bar = a[0];
  assign n49 = abar[0];
  OR2_X1 U17 ( .A1(n48), .A2(n64), .ZN(y[7]) );
  AND2_X1 U17bar ( .A1(n48bar), .A2(n64bar), .ZN(ybar[7]) );
  OR2_X1 U18 ( .A1(n63), .A2(b[7]), .ZN(n47) );
  AND2_X1 U18bar ( .A1(n63bar), .A2(bbar[7]), .ZN(n47bar) );
  AND2_X1 U19 ( .A1(b[7]), .A2(n63), .ZN(n48) );
  OR2_X1 U19bar ( .A1(bbar[7]), .A2(n63bar), .ZN(n48bar) );
  OR2_X1 U20 ( .A1(n46), .A2(n62), .ZN(y[6]) );
  AND2_X1 U20bar ( .A1(n46bar), .A2(n62bar), .ZN(ybar[6]) );
  OR2_X1 U21 ( .A1(n61), .A2(b[6]), .ZN(n45) );
  AND2_X1 U21bar ( .A1(n61bar), .A2(bbar[6]), .ZN(n45bar) );
  AND2_X1 U22 ( .A1(b[6]), .A2(n61), .ZN(n46) );
  OR2_X1 U22bar ( .A1(bbar[6]), .A2(n61bar), .ZN(n46bar) );
  OR2_X1 U23 ( .A1(n44), .A2(n60), .ZN(y[5]) );
  AND2_X1 U23bar ( .A1(n44bar), .A2(n60bar), .ZN(ybar[5]) );
  OR2_X1 U24 ( .A1(n59), .A2(b[5]), .ZN(n43) );
  AND2_X1 U24bar ( .A1(n59bar), .A2(bbar[5]), .ZN(n43bar) );
  AND2_X1 U25 ( .A1(b[5]), .A2(n59), .ZN(n44) );
  OR2_X1 U25bar ( .A1(bbar[5]), .A2(n59bar), .ZN(n44bar) );
  OR2_X1 U26 ( .A1(n42), .A2(n58), .ZN(y[4]) );
  AND2_X1 U26bar ( .A1(n42bar), .A2(n58bar), .ZN(ybar[4]) );
  OR2_X1 U27 ( .A1(n57), .A2(b[4]), .ZN(n41) );
  AND2_X1 U27bar ( .A1(n57bar), .A2(bbar[4]), .ZN(n41bar) );
  AND2_X1 U28 ( .A1(b[4]), .A2(n57), .ZN(n42) );
  OR2_X1 U28bar ( .A1(bbar[4]), .A2(n57bar), .ZN(n42bar) );
  OR2_X1 U29 ( .A1(n40), .A2(n56), .ZN(y[3]) );
  AND2_X1 U29bar ( .A1(n40bar), .A2(n56bar), .ZN(ybar[3]) );
  OR2_X1 U30 ( .A1(n55), .A2(b[3]), .ZN(n39) );
  AND2_X1 U30bar ( .A1(n55bar), .A2(bbar[3]), .ZN(n39bar) );
  AND2_X1 U31 ( .A1(b[3]), .A2(n55), .ZN(n40) );
  OR2_X1 U31bar ( .A1(bbar[3]), .A2(n55bar), .ZN(n40bar) );
  OR2_X1 U32 ( .A1(n38), .A2(n54), .ZN(y[2]) );
  AND2_X1 U32bar ( .A1(n38bar), .A2(n54bar), .ZN(ybar[2]) );
  OR2_X1 U33 ( .A1(n53), .A2(b[2]), .ZN(n37) );
  AND2_X1 U33bar ( .A1(n53bar), .A2(bbar[2]), .ZN(n37bar) );
  AND2_X1 U34 ( .A1(b[2]), .A2(n53), .ZN(n38) );
  OR2_X1 U34bar ( .A1(bbar[2]), .A2(n53bar), .ZN(n38bar) );
  OR2_X1 U35 ( .A1(n36), .A2(n52), .ZN(y[1]) );
  AND2_X1 U35bar ( .A1(n36bar), .A2(n52bar), .ZN(ybar[1]) );
  OR2_X1 U36 ( .A1(n51), .A2(b[1]), .ZN(n35) );
  AND2_X1 U36bar ( .A1(n51bar), .A2(bbar[1]), .ZN(n35bar) );
  AND2_X1 U37 ( .A1(b[1]), .A2(n51), .ZN(n36) );
  OR2_X1 U37bar ( .A1(bbar[1]), .A2(n51bar), .ZN(n36bar) );
  OR2_X1 U38 ( .A1(n34), .A2(n50), .ZN(y[0]) );
  AND2_X1 U38bar ( .A1(n34bar), .A2(n50bar), .ZN(ybar[0]) );
  OR2_X1 U39 ( .A1(n49), .A2(b[0]), .ZN(n33) );
  AND2_X1 U39bar ( .A1(n49bar), .A2(bbar[0]), .ZN(n33bar) );
  AND2_X1 U40 ( .A1(b[0]), .A2(n49), .ZN(n34) );
  OR2_X1 U40bar ( .A1(bbar[0]), .A2(n49bar), .ZN(n34bar) );
endmodule

module byteXor_4 ( a, b, y );

  input wire [7:0] a;
  input wire [7:0] b;
  wire [7:0] abar;
  wire [7:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
//input_done

  output wire [7:0] y;
  wire [7:0] ybar;
//output_done

  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n33bar;
  wire n34bar;
  wire n35bar;
  wire n36bar;
  wire n37bar;
  wire n38bar;
  wire n39bar;
  wire n40bar;
  wire n41bar;
  wire n42bar;
  wire n43bar;
  wire n44bar;
  wire n45bar;
  wire n46bar;
  wire n47bar;
  wire n48bar;
  wire n49bar;
  wire n50bar;
  wire n51bar;
  wire n52bar;
  wire n53bar;
  wire n54bar;
  wire n55bar;
  wire n56bar;
  wire n57bar;
  wire n58bar;
  wire n59bar;
  wire n60bar;
  wire n61bar;
  wire n62bar;
  wire n63bar;
  wire n64bar;
//wire_done

 //assign_done

  assign n64bar = n47;
  assign n64 = n47bar;
  assign n63bar = a[7];
  assign n63 = abar[7];
  assign n62bar = n45;
  assign n62 = n45bar;
  assign n61bar = a[6];
  assign n61 = abar[6];
  assign n60bar = n43;
  assign n60 = n43bar;
  assign n59bar = a[5];
  assign n59 = abar[5];
  assign n58bar = n41;
  assign n58 = n41bar;
  assign n57bar = a[4];
  assign n57 = abar[4];
  assign n56bar = n39;
  assign n56 = n39bar;
  assign n55bar = a[3];
  assign n55 = abar[3];
  assign n54bar = n37;
  assign n54 = n37bar;
  assign n53bar = a[2];
  assign n53 = abar[2];
  assign n52bar = n35;
  assign n52 = n35bar;
  assign n51bar = a[1];
  assign n51 = abar[1];
  assign n50bar = n33;
  assign n50 = n33bar;
  assign n49bar = a[0];
  assign n49 = abar[0];
  OR2_X1 U17 ( .A1(n48), .A2(n64), .ZN(y[7]) );
  AND2_X1 U17bar ( .A1(n48bar), .A2(n64bar), .ZN(ybar[7]) );
  OR2_X1 U18 ( .A1(n63), .A2(b[7]), .ZN(n47) );
  AND2_X1 U18bar ( .A1(n63bar), .A2(bbar[7]), .ZN(n47bar) );
  AND2_X1 U19 ( .A1(b[7]), .A2(n63), .ZN(n48) );
  OR2_X1 U19bar ( .A1(bbar[7]), .A2(n63bar), .ZN(n48bar) );
  OR2_X1 U20 ( .A1(n46), .A2(n62), .ZN(y[6]) );
  AND2_X1 U20bar ( .A1(n46bar), .A2(n62bar), .ZN(ybar[6]) );
  OR2_X1 U21 ( .A1(n61), .A2(b[6]), .ZN(n45) );
  AND2_X1 U21bar ( .A1(n61bar), .A2(bbar[6]), .ZN(n45bar) );
  AND2_X1 U22 ( .A1(b[6]), .A2(n61), .ZN(n46) );
  OR2_X1 U22bar ( .A1(bbar[6]), .A2(n61bar), .ZN(n46bar) );
  OR2_X1 U23 ( .A1(n44), .A2(n60), .ZN(y[5]) );
  AND2_X1 U23bar ( .A1(n44bar), .A2(n60bar), .ZN(ybar[5]) );
  OR2_X1 U24 ( .A1(n59), .A2(b[5]), .ZN(n43) );
  AND2_X1 U24bar ( .A1(n59bar), .A2(bbar[5]), .ZN(n43bar) );
  AND2_X1 U25 ( .A1(b[5]), .A2(n59), .ZN(n44) );
  OR2_X1 U25bar ( .A1(bbar[5]), .A2(n59bar), .ZN(n44bar) );
  OR2_X1 U26 ( .A1(n42), .A2(n58), .ZN(y[4]) );
  AND2_X1 U26bar ( .A1(n42bar), .A2(n58bar), .ZN(ybar[4]) );
  OR2_X1 U27 ( .A1(n57), .A2(b[4]), .ZN(n41) );
  AND2_X1 U27bar ( .A1(n57bar), .A2(bbar[4]), .ZN(n41bar) );
  AND2_X1 U28 ( .A1(b[4]), .A2(n57), .ZN(n42) );
  OR2_X1 U28bar ( .A1(bbar[4]), .A2(n57bar), .ZN(n42bar) );
  OR2_X1 U29 ( .A1(n40), .A2(n56), .ZN(y[3]) );
  AND2_X1 U29bar ( .A1(n40bar), .A2(n56bar), .ZN(ybar[3]) );
  OR2_X1 U30 ( .A1(n55), .A2(b[3]), .ZN(n39) );
  AND2_X1 U30bar ( .A1(n55bar), .A2(bbar[3]), .ZN(n39bar) );
  AND2_X1 U31 ( .A1(b[3]), .A2(n55), .ZN(n40) );
  OR2_X1 U31bar ( .A1(bbar[3]), .A2(n55bar), .ZN(n40bar) );
  OR2_X1 U32 ( .A1(n38), .A2(n54), .ZN(y[2]) );
  AND2_X1 U32bar ( .A1(n38bar), .A2(n54bar), .ZN(ybar[2]) );
  OR2_X1 U33 ( .A1(n53), .A2(b[2]), .ZN(n37) );
  AND2_X1 U33bar ( .A1(n53bar), .A2(bbar[2]), .ZN(n37bar) );
  AND2_X1 U34 ( .A1(b[2]), .A2(n53), .ZN(n38) );
  OR2_X1 U34bar ( .A1(bbar[2]), .A2(n53bar), .ZN(n38bar) );
  OR2_X1 U35 ( .A1(n36), .A2(n52), .ZN(y[1]) );
  AND2_X1 U35bar ( .A1(n36bar), .A2(n52bar), .ZN(ybar[1]) );
  OR2_X1 U36 ( .A1(n51), .A2(b[1]), .ZN(n35) );
  AND2_X1 U36bar ( .A1(n51bar), .A2(bbar[1]), .ZN(n35bar) );
  AND2_X1 U37 ( .A1(b[1]), .A2(n51), .ZN(n36) );
  OR2_X1 U37bar ( .A1(bbar[1]), .A2(n51bar), .ZN(n36bar) );
  OR2_X1 U38 ( .A1(n34), .A2(n50), .ZN(y[0]) );
  AND2_X1 U38bar ( .A1(n34bar), .A2(n50bar), .ZN(ybar[0]) );
  OR2_X1 U39 ( .A1(n49), .A2(b[0]), .ZN(n33) );
  AND2_X1 U39bar ( .A1(n49bar), .A2(bbar[0]), .ZN(n33bar) );
  AND2_X1 U40 ( .A1(b[0]), .A2(n49), .ZN(n34) );
  OR2_X1 U40bar ( .A1(bbar[0]), .A2(n49bar), .ZN(n34bar) );
endmodule

module byteXor_5 ( a, b, y );

  input wire [7:0] a;
  input wire [7:0] b;
  wire [7:0] abar;
  wire [7:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
//input_done

  output wire [7:0] y;
  wire [7:0] ybar;
//output_done

  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n33bar;
  wire n34bar;
  wire n35bar;
  wire n36bar;
  wire n37bar;
  wire n38bar;
  wire n39bar;
  wire n40bar;
  wire n41bar;
  wire n42bar;
  wire n43bar;
  wire n44bar;
  wire n45bar;
  wire n46bar;
  wire n47bar;
  wire n48bar;
  wire n49bar;
  wire n50bar;
  wire n51bar;
  wire n52bar;
  wire n53bar;
  wire n54bar;
  wire n55bar;
  wire n56bar;
  wire n57bar;
  wire n58bar;
  wire n59bar;
  wire n60bar;
  wire n61bar;
  wire n62bar;
  wire n63bar;
  wire n64bar;
//wire_done

 //assign_done

  assign n64bar = n47;
  assign n64 = n47bar;
  assign n63bar = a[7];
  assign n63 = abar[7];
  assign n62bar = n45;
  assign n62 = n45bar;
  assign n61bar = a[6];
  assign n61 = abar[6];
  assign n60bar = n43;
  assign n60 = n43bar;
  assign n59bar = a[5];
  assign n59 = abar[5];
  assign n58bar = n41;
  assign n58 = n41bar;
  assign n57bar = a[4];
  assign n57 = abar[4];
  assign n56bar = n39;
  assign n56 = n39bar;
  assign n55bar = a[3];
  assign n55 = abar[3];
  assign n54bar = n37;
  assign n54 = n37bar;
  assign n53bar = a[2];
  assign n53 = abar[2];
  assign n52bar = n35;
  assign n52 = n35bar;
  assign n51bar = a[1];
  assign n51 = abar[1];
  assign n50bar = n33;
  assign n50 = n33bar;
  assign n49bar = a[0];
  assign n49 = abar[0];
  OR2_X1 U17 ( .A1(n48), .A2(n64), .ZN(y[7]) );
  AND2_X1 U17bar ( .A1(n48bar), .A2(n64bar), .ZN(ybar[7]) );
  OR2_X1 U18 ( .A1(n63), .A2(b[7]), .ZN(n47) );
  AND2_X1 U18bar ( .A1(n63bar), .A2(bbar[7]), .ZN(n47bar) );
  AND2_X1 U19 ( .A1(b[7]), .A2(n63), .ZN(n48) );
  OR2_X1 U19bar ( .A1(bbar[7]), .A2(n63bar), .ZN(n48bar) );
  OR2_X1 U20 ( .A1(n46), .A2(n62), .ZN(y[6]) );
  AND2_X1 U20bar ( .A1(n46bar), .A2(n62bar), .ZN(ybar[6]) );
  OR2_X1 U21 ( .A1(n61), .A2(b[6]), .ZN(n45) );
  AND2_X1 U21bar ( .A1(n61bar), .A2(bbar[6]), .ZN(n45bar) );
  AND2_X1 U22 ( .A1(b[6]), .A2(n61), .ZN(n46) );
  OR2_X1 U22bar ( .A1(bbar[6]), .A2(n61bar), .ZN(n46bar) );
  OR2_X1 U23 ( .A1(n44), .A2(n60), .ZN(y[5]) );
  AND2_X1 U23bar ( .A1(n44bar), .A2(n60bar), .ZN(ybar[5]) );
  OR2_X1 U24 ( .A1(n59), .A2(b[5]), .ZN(n43) );
  AND2_X1 U24bar ( .A1(n59bar), .A2(bbar[5]), .ZN(n43bar) );
  AND2_X1 U25 ( .A1(b[5]), .A2(n59), .ZN(n44) );
  OR2_X1 U25bar ( .A1(bbar[5]), .A2(n59bar), .ZN(n44bar) );
  OR2_X1 U26 ( .A1(n42), .A2(n58), .ZN(y[4]) );
  AND2_X1 U26bar ( .A1(n42bar), .A2(n58bar), .ZN(ybar[4]) );
  OR2_X1 U27 ( .A1(n57), .A2(b[4]), .ZN(n41) );
  AND2_X1 U27bar ( .A1(n57bar), .A2(bbar[4]), .ZN(n41bar) );
  AND2_X1 U28 ( .A1(b[4]), .A2(n57), .ZN(n42) );
  OR2_X1 U28bar ( .A1(bbar[4]), .A2(n57bar), .ZN(n42bar) );
  OR2_X1 U29 ( .A1(n40), .A2(n56), .ZN(y[3]) );
  AND2_X1 U29bar ( .A1(n40bar), .A2(n56bar), .ZN(ybar[3]) );
  OR2_X1 U30 ( .A1(n55), .A2(b[3]), .ZN(n39) );
  AND2_X1 U30bar ( .A1(n55bar), .A2(bbar[3]), .ZN(n39bar) );
  AND2_X1 U31 ( .A1(b[3]), .A2(n55), .ZN(n40) );
  OR2_X1 U31bar ( .A1(bbar[3]), .A2(n55bar), .ZN(n40bar) );
  OR2_X1 U32 ( .A1(n38), .A2(n54), .ZN(y[2]) );
  AND2_X1 U32bar ( .A1(n38bar), .A2(n54bar), .ZN(ybar[2]) );
  OR2_X1 U33 ( .A1(n53), .A2(b[2]), .ZN(n37) );
  AND2_X1 U33bar ( .A1(n53bar), .A2(bbar[2]), .ZN(n37bar) );
  AND2_X1 U34 ( .A1(b[2]), .A2(n53), .ZN(n38) );
  OR2_X1 U34bar ( .A1(bbar[2]), .A2(n53bar), .ZN(n38bar) );
  OR2_X1 U35 ( .A1(n36), .A2(n52), .ZN(y[1]) );
  AND2_X1 U35bar ( .A1(n36bar), .A2(n52bar), .ZN(ybar[1]) );
  OR2_X1 U36 ( .A1(n51), .A2(b[1]), .ZN(n35) );
  AND2_X1 U36bar ( .A1(n51bar), .A2(bbar[1]), .ZN(n35bar) );
  AND2_X1 U37 ( .A1(b[1]), .A2(n51), .ZN(n36) );
  OR2_X1 U37bar ( .A1(bbar[1]), .A2(n51bar), .ZN(n36bar) );
  OR2_X1 U38 ( .A1(n34), .A2(n50), .ZN(y[0]) );
  AND2_X1 U38bar ( .A1(n34bar), .A2(n50bar), .ZN(ybar[0]) );
  OR2_X1 U39 ( .A1(n49), .A2(b[0]), .ZN(n33) );
  AND2_X1 U39bar ( .A1(n49bar), .A2(bbar[0]), .ZN(n33bar) );
  AND2_X1 U40 ( .A1(b[0]), .A2(n49), .ZN(n34) );
  OR2_X1 U40bar ( .A1(bbar[0]), .A2(n49bar), .ZN(n34bar) );
endmodule

module byteXor4_1 ( a, b, c, d, y );

  input wire [7:0] a;
  input wire [7:0] b;
  input wire [7:0] c;
  input wire [7:0] d;
  wire [7:0] abar;
  wire [7:0] bbar;
  wire [7:0] cbar;
  wire [7:0] dbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign cbar[0] = ~c[0];
  assign cbar[1] = ~c[1];
  assign cbar[2] = ~c[2];
  assign cbar[3] = ~c[3];
  assign cbar[4] = ~c[4];
  assign cbar[5] = ~c[5];
  assign cbar[6] = ~c[6];
  assign cbar[7] = ~c[7];
  assign dbar[0] = ~d[0];
  assign dbar[1] = ~d[1];
  assign dbar[2] = ~d[2];
  assign dbar[3] = ~d[3];
  assign dbar[4] = ~d[4];
  assign dbar[5] = ~d[5];
  assign dbar[6] = ~d[6];
  assign dbar[7] = ~d[7];
//input_done

  output wire [7:0] y;
  wire [7:0] ybar;
//output_done

  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n113bar;
  wire n114bar;
  wire n115bar;
  wire n116bar;
  wire n117bar;
  wire n118bar;
  wire n119bar;
  wire n120bar;
  wire n121bar;
  wire n122bar;
  wire n123bar;
  wire n124bar;
  wire n125bar;
  wire n126bar;
  wire n127bar;
  wire n128bar;
  wire n129bar;
  wire n130bar;
  wire n131bar;
  wire n132bar;
  wire n133bar;
  wire n134bar;
  wire n135bar;
  wire n136bar;
  wire n137bar;
  wire n138bar;
  wire n139bar;
  wire n140bar;
  wire n141bar;
  wire n142bar;
  wire n143bar;
  wire n144bar;
  wire n145bar;
  wire n146bar;
  wire n147bar;
  wire n148bar;
  wire n149bar;
  wire n150bar;
  wire n151bar;
  wire n152bar;
  wire n153bar;
  wire n154bar;
  wire n155bar;
  wire n156bar;
  wire n157bar;
  wire n158bar;
  wire n159bar;
  wire n160bar;
  wire n161bar;
  wire n162bar;
  wire n163bar;
  wire n164bar;
  wire n165bar;
  wire n166bar;
  wire n167bar;
  wire n168bar;
  wire n169bar;
  wire n170bar;
  wire n171bar;
  wire n172bar;
  wire n173bar;
  wire n174bar;
  wire n175bar;
  wire n176bar;
  wire n177bar;
  wire n178bar;
  wire n179bar;
  wire n180bar;
  wire n181bar;
  wire n182bar;
  wire n183bar;
  wire n184bar;
  wire n185bar;
  wire n186bar;
  wire n187bar;
  wire n188bar;
  wire n189bar;
  wire n190bar;
  wire n191bar;
  wire n192bar;
  wire n193bar;
  wire n194bar;
  wire n195bar;
  wire n196bar;
  wire n197bar;
  wire n198bar;
  wire n199bar;
  wire n200bar;
  wire n201bar;
  wire n202bar;
  wire n203bar;
  wire n204bar;
  wire n205bar;
  wire n206bar;
  wire n207bar;
  wire n208bar;
  wire n209bar;
  wire n210bar;
  wire n211bar;
  wire n212bar;
  wire n213bar;
  wire n214bar;
  wire n215bar;
  wire n216bar;
  wire n217bar;
  wire n218bar;
  wire n219bar;
  wire n220bar;
  wire n221bar;
  wire n222bar;
  wire n223bar;
  wire n224bar;
//wire_done

 //assign_done

  assign n224bar = n175;
  assign n224 = n175bar;
  assign n223bar = a[7];
  assign n223 = abar[7];
  assign n222bar = n167;
  assign n222 = n167bar;
  assign n221bar = a[6];
  assign n221 = abar[6];
  assign n220bar = n159;
  assign n220 = n159bar;
  assign n219bar = a[5];
  assign n219 = abar[5];
  assign n218bar = n151;
  assign n218 = n151bar;
  assign n217bar = a[4];
  assign n217 = abar[4];
  assign n216bar = n143;
  assign n216 = n143bar;
  assign n215bar = a[3];
  assign n215 = abar[3];
  assign n214bar = n135;
  assign n214 = n135bar;
  assign n213bar = a[2];
  assign n213 = abar[2];
  assign n212bar = n127;
  assign n212 = n127bar;
  assign n211bar = a[1];
  assign n211 = abar[1];
  assign n210bar = n119;
  assign n210 = n119bar;
  assign n209bar = a[0];
  assign n209 = abar[0];
  assign n208bar = b[7];
  assign n208 = bbar[7];
  assign n207bar = b[6];
  assign n207 = bbar[6];
  assign n206bar = b[5];
  assign n206 = bbar[5];
  assign n205bar = b[4];
  assign n205 = bbar[4];
  assign n204bar = b[3];
  assign n204 = bbar[3];
  assign n203bar = b[2];
  assign n203 = bbar[2];
  assign n202bar = b[1];
  assign n202 = bbar[1];
  assign n201bar = b[0];
  assign n201 = bbar[0];
  assign n200bar = n171;
  assign n200 = n171bar;
  assign n199bar = c[7];
  assign n199 = cbar[7];
  assign n198bar = n163;
  assign n198 = n163bar;
  assign n197bar = c[6];
  assign n197 = cbar[6];
  assign n196bar = n155;
  assign n196 = n155bar;
  assign n195bar = c[5];
  assign n195 = cbar[5];
  assign n194bar = n147;
  assign n194 = n147bar;
  assign n193bar = c[4];
  assign n193 = cbar[4];
  assign n192bar = n139;
  assign n192 = n139bar;
  assign n191bar = c[3];
  assign n191 = cbar[3];
  assign n190bar = n131;
  assign n190 = n131bar;
  assign n189bar = c[2];
  assign n189 = cbar[2];
  assign n188bar = n123;
  assign n188 = n123bar;
  assign n187bar = c[1];
  assign n187 = cbar[1];
  assign n186bar = n115;
  assign n186 = n115bar;
  assign n185bar = c[0];
  assign n185 = cbar[0];
  assign n184bar = d[7];
  assign n184 = dbar[7];
  assign n183bar = d[6];
  assign n183 = dbar[6];
  assign n182bar = d[5];
  assign n182 = dbar[5];
  assign n181bar = d[4];
  assign n181 = dbar[4];
  assign n180bar = d[3];
  assign n180 = dbar[3];
  assign n179bar = d[2];
  assign n179 = dbar[2];
  assign n178bar = d[1];
  assign n178 = dbar[1];
  assign n177bar = d[0];
  assign n177 = dbar[0];
  OR2_X1 U49 ( .A1(n176), .A2(n224), .ZN(y[7]) );
  AND2_X1 U49bar ( .A1(n176bar), .A2(n224bar), .ZN(ybar[7]) );
  OR2_X1 U50 ( .A1(n174), .A2(n200), .ZN(n175) );
  AND2_X1 U50bar ( .A1(n174bar), .A2(n200bar), .ZN(n175bar) );
  AND2_X1 U51 ( .A1(n200), .A2(n174), .ZN(n176) );
  OR2_X1 U51bar ( .A1(n200bar), .A2(n174bar), .ZN(n176bar) );
  AND2_X1 U52 ( .A1(n173), .A2(n172), .ZN(n174) );
  OR2_X1 U52bar ( .A1(n173bar), .A2(n172bar), .ZN(n174bar) );
  OR2_X1 U53 ( .A1(n223), .A2(b[7]), .ZN(n172) );
  AND2_X1 U53bar ( .A1(n223bar), .A2(bbar[7]), .ZN(n172bar) );
  OR2_X1 U54 ( .A1(n208), .A2(a[7]), .ZN(n173) );
  AND2_X1 U54bar ( .A1(n208bar), .A2(abar[7]), .ZN(n173bar) );
  AND2_X1 U55 ( .A1(n170), .A2(n169), .ZN(n171) );
  OR2_X1 U55bar ( .A1(n170bar), .A2(n169bar), .ZN(n171bar) );
  OR2_X1 U56 ( .A1(n199), .A2(d[7]), .ZN(n169) );
  AND2_X1 U56bar ( .A1(n199bar), .A2(dbar[7]), .ZN(n169bar) );
  OR2_X1 U57 ( .A1(n184), .A2(c[7]), .ZN(n170) );
  AND2_X1 U57bar ( .A1(n184bar), .A2(cbar[7]), .ZN(n170bar) );
  OR2_X1 U58 ( .A1(n168), .A2(n222), .ZN(y[6]) );
  AND2_X1 U58bar ( .A1(n168bar), .A2(n222bar), .ZN(ybar[6]) );
  OR2_X1 U59 ( .A1(n166), .A2(n198), .ZN(n167) );
  AND2_X1 U59bar ( .A1(n166bar), .A2(n198bar), .ZN(n167bar) );
  AND2_X1 U60 ( .A1(n198), .A2(n166), .ZN(n168) );
  OR2_X1 U60bar ( .A1(n198bar), .A2(n166bar), .ZN(n168bar) );
  AND2_X1 U61 ( .A1(n165), .A2(n164), .ZN(n166) );
  OR2_X1 U61bar ( .A1(n165bar), .A2(n164bar), .ZN(n166bar) );
  OR2_X1 U62 ( .A1(n221), .A2(b[6]), .ZN(n164) );
  AND2_X1 U62bar ( .A1(n221bar), .A2(bbar[6]), .ZN(n164bar) );
  OR2_X1 U63 ( .A1(n207), .A2(a[6]), .ZN(n165) );
  AND2_X1 U63bar ( .A1(n207bar), .A2(abar[6]), .ZN(n165bar) );
  AND2_X1 U64 ( .A1(n162), .A2(n161), .ZN(n163) );
  OR2_X1 U64bar ( .A1(n162bar), .A2(n161bar), .ZN(n163bar) );
  OR2_X1 U65 ( .A1(n197), .A2(d[6]), .ZN(n161) );
  AND2_X1 U65bar ( .A1(n197bar), .A2(dbar[6]), .ZN(n161bar) );
  OR2_X1 U66 ( .A1(n183), .A2(c[6]), .ZN(n162) );
  AND2_X1 U66bar ( .A1(n183bar), .A2(cbar[6]), .ZN(n162bar) );
  OR2_X1 U67 ( .A1(n160), .A2(n220), .ZN(y[5]) );
  AND2_X1 U67bar ( .A1(n160bar), .A2(n220bar), .ZN(ybar[5]) );
  OR2_X1 U68 ( .A1(n158), .A2(n196), .ZN(n159) );
  AND2_X1 U68bar ( .A1(n158bar), .A2(n196bar), .ZN(n159bar) );
  AND2_X1 U69 ( .A1(n196), .A2(n158), .ZN(n160) );
  OR2_X1 U69bar ( .A1(n196bar), .A2(n158bar), .ZN(n160bar) );
  AND2_X1 U70 ( .A1(n157), .A2(n156), .ZN(n158) );
  OR2_X1 U70bar ( .A1(n157bar), .A2(n156bar), .ZN(n158bar) );
  OR2_X1 U71 ( .A1(n219), .A2(b[5]), .ZN(n156) );
  AND2_X1 U71bar ( .A1(n219bar), .A2(bbar[5]), .ZN(n156bar) );
  OR2_X1 U72 ( .A1(n206), .A2(a[5]), .ZN(n157) );
  AND2_X1 U72bar ( .A1(n206bar), .A2(abar[5]), .ZN(n157bar) );
  AND2_X1 U73 ( .A1(n154), .A2(n153), .ZN(n155) );
  OR2_X1 U73bar ( .A1(n154bar), .A2(n153bar), .ZN(n155bar) );
  OR2_X1 U74 ( .A1(n195), .A2(d[5]), .ZN(n153) );
  AND2_X1 U74bar ( .A1(n195bar), .A2(dbar[5]), .ZN(n153bar) );
  OR2_X1 U75 ( .A1(n182), .A2(c[5]), .ZN(n154) );
  AND2_X1 U75bar ( .A1(n182bar), .A2(cbar[5]), .ZN(n154bar) );
  OR2_X1 U76 ( .A1(n152), .A2(n218), .ZN(y[4]) );
  AND2_X1 U76bar ( .A1(n152bar), .A2(n218bar), .ZN(ybar[4]) );
  OR2_X1 U77 ( .A1(n150), .A2(n194), .ZN(n151) );
  AND2_X1 U77bar ( .A1(n150bar), .A2(n194bar), .ZN(n151bar) );
  AND2_X1 U78 ( .A1(n194), .A2(n150), .ZN(n152) );
  OR2_X1 U78bar ( .A1(n194bar), .A2(n150bar), .ZN(n152bar) );
  AND2_X1 U79 ( .A1(n149), .A2(n148), .ZN(n150) );
  OR2_X1 U79bar ( .A1(n149bar), .A2(n148bar), .ZN(n150bar) );
  OR2_X1 U80 ( .A1(n217), .A2(b[4]), .ZN(n148) );
  AND2_X1 U80bar ( .A1(n217bar), .A2(bbar[4]), .ZN(n148bar) );
  OR2_X1 U81 ( .A1(n205), .A2(a[4]), .ZN(n149) );
  AND2_X1 U81bar ( .A1(n205bar), .A2(abar[4]), .ZN(n149bar) );
  AND2_X1 U82 ( .A1(n146), .A2(n145), .ZN(n147) );
  OR2_X1 U82bar ( .A1(n146bar), .A2(n145bar), .ZN(n147bar) );
  OR2_X1 U83 ( .A1(n193), .A2(d[4]), .ZN(n145) );
  AND2_X1 U83bar ( .A1(n193bar), .A2(dbar[4]), .ZN(n145bar) );
  OR2_X1 U84 ( .A1(n181), .A2(c[4]), .ZN(n146) );
  AND2_X1 U84bar ( .A1(n181bar), .A2(cbar[4]), .ZN(n146bar) );
  OR2_X1 U85 ( .A1(n144), .A2(n216), .ZN(y[3]) );
  AND2_X1 U85bar ( .A1(n144bar), .A2(n216bar), .ZN(ybar[3]) );
  OR2_X1 U86 ( .A1(n142), .A2(n192), .ZN(n143) );
  AND2_X1 U86bar ( .A1(n142bar), .A2(n192bar), .ZN(n143bar) );
  AND2_X1 U87 ( .A1(n192), .A2(n142), .ZN(n144) );
  OR2_X1 U87bar ( .A1(n192bar), .A2(n142bar), .ZN(n144bar) );
  AND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(n142) );
  OR2_X1 U88bar ( .A1(n141bar), .A2(n140bar), .ZN(n142bar) );
  OR2_X1 U89 ( .A1(n215), .A2(b[3]), .ZN(n140) );
  AND2_X1 U89bar ( .A1(n215bar), .A2(bbar[3]), .ZN(n140bar) );
  OR2_X1 U90 ( .A1(n204), .A2(a[3]), .ZN(n141) );
  AND2_X1 U90bar ( .A1(n204bar), .A2(abar[3]), .ZN(n141bar) );
  AND2_X1 U91 ( .A1(n138), .A2(n137), .ZN(n139) );
  OR2_X1 U91bar ( .A1(n138bar), .A2(n137bar), .ZN(n139bar) );
  OR2_X1 U92 ( .A1(n191), .A2(d[3]), .ZN(n137) );
  AND2_X1 U92bar ( .A1(n191bar), .A2(dbar[3]), .ZN(n137bar) );
  OR2_X1 U93 ( .A1(n180), .A2(c[3]), .ZN(n138) );
  AND2_X1 U93bar ( .A1(n180bar), .A2(cbar[3]), .ZN(n138bar) );
  OR2_X1 U94 ( .A1(n136), .A2(n214), .ZN(y[2]) );
  AND2_X1 U94bar ( .A1(n136bar), .A2(n214bar), .ZN(ybar[2]) );
  OR2_X1 U95 ( .A1(n134), .A2(n190), .ZN(n135) );
  AND2_X1 U95bar ( .A1(n134bar), .A2(n190bar), .ZN(n135bar) );
  AND2_X1 U96 ( .A1(n190), .A2(n134), .ZN(n136) );
  OR2_X1 U96bar ( .A1(n190bar), .A2(n134bar), .ZN(n136bar) );
  AND2_X1 U97 ( .A1(n133), .A2(n132), .ZN(n134) );
  OR2_X1 U97bar ( .A1(n133bar), .A2(n132bar), .ZN(n134bar) );
  OR2_X1 U98 ( .A1(n213), .A2(b[2]), .ZN(n132) );
  AND2_X1 U98bar ( .A1(n213bar), .A2(bbar[2]), .ZN(n132bar) );
  OR2_X1 U99 ( .A1(n203), .A2(a[2]), .ZN(n133) );
  AND2_X1 U99bar ( .A1(n203bar), .A2(abar[2]), .ZN(n133bar) );
  AND2_X1 U100 ( .A1(n130), .A2(n129), .ZN(n131) );
  OR2_X1 U100bar ( .A1(n130bar), .A2(n129bar), .ZN(n131bar) );
  OR2_X1 U101 ( .A1(n189), .A2(d[2]), .ZN(n129) );
  AND2_X1 U101bar ( .A1(n189bar), .A2(dbar[2]), .ZN(n129bar) );
  OR2_X1 U102 ( .A1(n179), .A2(c[2]), .ZN(n130) );
  AND2_X1 U102bar ( .A1(n179bar), .A2(cbar[2]), .ZN(n130bar) );
  OR2_X1 U103 ( .A1(n128), .A2(n212), .ZN(y[1]) );
  AND2_X1 U103bar ( .A1(n128bar), .A2(n212bar), .ZN(ybar[1]) );
  OR2_X1 U104 ( .A1(n126), .A2(n188), .ZN(n127) );
  AND2_X1 U104bar ( .A1(n126bar), .A2(n188bar), .ZN(n127bar) );
  AND2_X1 U105 ( .A1(n188), .A2(n126), .ZN(n128) );
  OR2_X1 U105bar ( .A1(n188bar), .A2(n126bar), .ZN(n128bar) );
  AND2_X1 U106 ( .A1(n125), .A2(n124), .ZN(n126) );
  OR2_X1 U106bar ( .A1(n125bar), .A2(n124bar), .ZN(n126bar) );
  OR2_X1 U107 ( .A1(n211), .A2(b[1]), .ZN(n124) );
  AND2_X1 U107bar ( .A1(n211bar), .A2(bbar[1]), .ZN(n124bar) );
  OR2_X1 U108 ( .A1(n202), .A2(a[1]), .ZN(n125) );
  AND2_X1 U108bar ( .A1(n202bar), .A2(abar[1]), .ZN(n125bar) );
  AND2_X1 U109 ( .A1(n122), .A2(n121), .ZN(n123) );
  OR2_X1 U109bar ( .A1(n122bar), .A2(n121bar), .ZN(n123bar) );
  OR2_X1 U110 ( .A1(n187), .A2(d[1]), .ZN(n121) );
  AND2_X1 U110bar ( .A1(n187bar), .A2(dbar[1]), .ZN(n121bar) );
  OR2_X1 U111 ( .A1(n178), .A2(c[1]), .ZN(n122) );
  AND2_X1 U111bar ( .A1(n178bar), .A2(cbar[1]), .ZN(n122bar) );
  OR2_X1 U112 ( .A1(n120), .A2(n210), .ZN(y[0]) );
  AND2_X1 U112bar ( .A1(n120bar), .A2(n210bar), .ZN(ybar[0]) );
  OR2_X1 U113 ( .A1(n118), .A2(n186), .ZN(n119) );
  AND2_X1 U113bar ( .A1(n118bar), .A2(n186bar), .ZN(n119bar) );
  AND2_X1 U114 ( .A1(n186), .A2(n118), .ZN(n120) );
  OR2_X1 U114bar ( .A1(n186bar), .A2(n118bar), .ZN(n120bar) );
  AND2_X1 U115 ( .A1(n117), .A2(n116), .ZN(n118) );
  OR2_X1 U115bar ( .A1(n117bar), .A2(n116bar), .ZN(n118bar) );
  OR2_X1 U116 ( .A1(n209), .A2(b[0]), .ZN(n116) );
  AND2_X1 U116bar ( .A1(n209bar), .A2(bbar[0]), .ZN(n116bar) );
  OR2_X1 U117 ( .A1(n201), .A2(a[0]), .ZN(n117) );
  AND2_X1 U117bar ( .A1(n201bar), .A2(abar[0]), .ZN(n117bar) );
  AND2_X1 U118 ( .A1(n114), .A2(n113), .ZN(n115) );
  OR2_X1 U118bar ( .A1(n114bar), .A2(n113bar), .ZN(n115bar) );
  OR2_X1 U119 ( .A1(n185), .A2(d[0]), .ZN(n113) );
  AND2_X1 U119bar ( .A1(n185bar), .A2(dbar[0]), .ZN(n113bar) );
  OR2_X1 U120 ( .A1(n177), .A2(c[0]), .ZN(n114) );
  AND2_X1 U120bar ( .A1(n177bar), .A2(cbar[0]), .ZN(n114bar) );
endmodule

module byteXor4_2 ( a, b, c, d, y );

  input wire [7:0] a;
  input wire [7:0] b;
  input wire [7:0] c;
  input wire [7:0] d;
  wire [7:0] abar;
  wire [7:0] bbar;
  wire [7:0] cbar;
  wire [7:0] dbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign cbar[0] = ~c[0];
  assign cbar[1] = ~c[1];
  assign cbar[2] = ~c[2];
  assign cbar[3] = ~c[3];
  assign cbar[4] = ~c[4];
  assign cbar[5] = ~c[5];
  assign cbar[6] = ~c[6];
  assign cbar[7] = ~c[7];
  assign dbar[0] = ~d[0];
  assign dbar[1] = ~d[1];
  assign dbar[2] = ~d[2];
  assign dbar[3] = ~d[3];
  assign dbar[4] = ~d[4];
  assign dbar[5] = ~d[5];
  assign dbar[6] = ~d[6];
  assign dbar[7] = ~d[7];
//input_done

  output wire [7:0] y;
  wire [7:0] ybar;
//output_done

  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n113bar;
  wire n114bar;
  wire n115bar;
  wire n116bar;
  wire n117bar;
  wire n118bar;
  wire n119bar;
  wire n120bar;
  wire n121bar;
  wire n122bar;
  wire n123bar;
  wire n124bar;
  wire n125bar;
  wire n126bar;
  wire n127bar;
  wire n128bar;
  wire n129bar;
  wire n130bar;
  wire n131bar;
  wire n132bar;
  wire n133bar;
  wire n134bar;
  wire n135bar;
  wire n136bar;
  wire n137bar;
  wire n138bar;
  wire n139bar;
  wire n140bar;
  wire n141bar;
  wire n142bar;
  wire n143bar;
  wire n144bar;
  wire n145bar;
  wire n146bar;
  wire n147bar;
  wire n148bar;
  wire n149bar;
  wire n150bar;
  wire n151bar;
  wire n152bar;
  wire n153bar;
  wire n154bar;
  wire n155bar;
  wire n156bar;
  wire n157bar;
  wire n158bar;
  wire n159bar;
  wire n160bar;
  wire n161bar;
  wire n162bar;
  wire n163bar;
  wire n164bar;
  wire n165bar;
  wire n166bar;
  wire n167bar;
  wire n168bar;
  wire n169bar;
  wire n170bar;
  wire n171bar;
  wire n172bar;
  wire n173bar;
  wire n174bar;
  wire n175bar;
  wire n176bar;
  wire n177bar;
  wire n178bar;
  wire n179bar;
  wire n180bar;
  wire n181bar;
  wire n182bar;
  wire n183bar;
  wire n184bar;
  wire n185bar;
  wire n186bar;
  wire n187bar;
  wire n188bar;
  wire n189bar;
  wire n190bar;
  wire n191bar;
  wire n192bar;
  wire n193bar;
  wire n194bar;
  wire n195bar;
  wire n196bar;
  wire n197bar;
  wire n198bar;
  wire n199bar;
  wire n200bar;
  wire n201bar;
  wire n202bar;
  wire n203bar;
  wire n204bar;
  wire n205bar;
  wire n206bar;
  wire n207bar;
  wire n208bar;
  wire n209bar;
  wire n210bar;
  wire n211bar;
  wire n212bar;
  wire n213bar;
  wire n214bar;
  wire n215bar;
  wire n216bar;
  wire n217bar;
  wire n218bar;
  wire n219bar;
  wire n220bar;
  wire n221bar;
  wire n222bar;
  wire n223bar;
  wire n224bar;
//wire_done

 //assign_done

  assign n224bar = n175;
  assign n224 = n175bar;
  assign n223bar = a[7];
  assign n223 = abar[7];
  assign n222bar = n167;
  assign n222 = n167bar;
  assign n221bar = a[6];
  assign n221 = abar[6];
  assign n220bar = n159;
  assign n220 = n159bar;
  assign n219bar = a[5];
  assign n219 = abar[5];
  assign n218bar = n151;
  assign n218 = n151bar;
  assign n217bar = a[4];
  assign n217 = abar[4];
  assign n216bar = n143;
  assign n216 = n143bar;
  assign n215bar = a[3];
  assign n215 = abar[3];
  assign n214bar = n135;
  assign n214 = n135bar;
  assign n213bar = a[2];
  assign n213 = abar[2];
  assign n212bar = n127;
  assign n212 = n127bar;
  assign n211bar = a[1];
  assign n211 = abar[1];
  assign n210bar = n119;
  assign n210 = n119bar;
  assign n209bar = a[0];
  assign n209 = abar[0];
  assign n208bar = b[7];
  assign n208 = bbar[7];
  assign n207bar = b[6];
  assign n207 = bbar[6];
  assign n206bar = b[5];
  assign n206 = bbar[5];
  assign n205bar = b[4];
  assign n205 = bbar[4];
  assign n204bar = b[3];
  assign n204 = bbar[3];
  assign n203bar = b[2];
  assign n203 = bbar[2];
  assign n202bar = b[1];
  assign n202 = bbar[1];
  assign n201bar = b[0];
  assign n201 = bbar[0];
  assign n200bar = n171;
  assign n200 = n171bar;
  assign n199bar = c[7];
  assign n199 = cbar[7];
  assign n198bar = n163;
  assign n198 = n163bar;
  assign n197bar = c[6];
  assign n197 = cbar[6];
  assign n196bar = n155;
  assign n196 = n155bar;
  assign n195bar = c[5];
  assign n195 = cbar[5];
  assign n194bar = n147;
  assign n194 = n147bar;
  assign n193bar = c[4];
  assign n193 = cbar[4];
  assign n192bar = n139;
  assign n192 = n139bar;
  assign n191bar = c[3];
  assign n191 = cbar[3];
  assign n190bar = n131;
  assign n190 = n131bar;
  assign n189bar = c[2];
  assign n189 = cbar[2];
  assign n188bar = n123;
  assign n188 = n123bar;
  assign n187bar = c[1];
  assign n187 = cbar[1];
  assign n186bar = n115;
  assign n186 = n115bar;
  assign n185bar = c[0];
  assign n185 = cbar[0];
  assign n184bar = d[7];
  assign n184 = dbar[7];
  assign n183bar = d[6];
  assign n183 = dbar[6];
  assign n182bar = d[5];
  assign n182 = dbar[5];
  assign n181bar = d[4];
  assign n181 = dbar[4];
  assign n180bar = d[3];
  assign n180 = dbar[3];
  assign n179bar = d[2];
  assign n179 = dbar[2];
  assign n178bar = d[1];
  assign n178 = dbar[1];
  assign n177bar = d[0];
  assign n177 = dbar[0];
  OR2_X1 U49 ( .A1(n176), .A2(n224), .ZN(y[7]) );
  AND2_X1 U49bar ( .A1(n176bar), .A2(n224bar), .ZN(ybar[7]) );
  OR2_X1 U50 ( .A1(n174), .A2(n200), .ZN(n175) );
  AND2_X1 U50bar ( .A1(n174bar), .A2(n200bar), .ZN(n175bar) );
  AND2_X1 U51 ( .A1(n200), .A2(n174), .ZN(n176) );
  OR2_X1 U51bar ( .A1(n200bar), .A2(n174bar), .ZN(n176bar) );
  AND2_X1 U52 ( .A1(n173), .A2(n172), .ZN(n174) );
  OR2_X1 U52bar ( .A1(n173bar), .A2(n172bar), .ZN(n174bar) );
  OR2_X1 U53 ( .A1(n223), .A2(b[7]), .ZN(n172) );
  AND2_X1 U53bar ( .A1(n223bar), .A2(bbar[7]), .ZN(n172bar) );
  OR2_X1 U54 ( .A1(n208), .A2(a[7]), .ZN(n173) );
  AND2_X1 U54bar ( .A1(n208bar), .A2(abar[7]), .ZN(n173bar) );
  AND2_X1 U55 ( .A1(n170), .A2(n169), .ZN(n171) );
  OR2_X1 U55bar ( .A1(n170bar), .A2(n169bar), .ZN(n171bar) );
  OR2_X1 U56 ( .A1(n199), .A2(d[7]), .ZN(n169) );
  AND2_X1 U56bar ( .A1(n199bar), .A2(dbar[7]), .ZN(n169bar) );
  OR2_X1 U57 ( .A1(n184), .A2(c[7]), .ZN(n170) );
  AND2_X1 U57bar ( .A1(n184bar), .A2(cbar[7]), .ZN(n170bar) );
  OR2_X1 U58 ( .A1(n168), .A2(n222), .ZN(y[6]) );
  AND2_X1 U58bar ( .A1(n168bar), .A2(n222bar), .ZN(ybar[6]) );
  OR2_X1 U59 ( .A1(n166), .A2(n198), .ZN(n167) );
  AND2_X1 U59bar ( .A1(n166bar), .A2(n198bar), .ZN(n167bar) );
  AND2_X1 U60 ( .A1(n198), .A2(n166), .ZN(n168) );
  OR2_X1 U60bar ( .A1(n198bar), .A2(n166bar), .ZN(n168bar) );
  AND2_X1 U61 ( .A1(n165), .A2(n164), .ZN(n166) );
  OR2_X1 U61bar ( .A1(n165bar), .A2(n164bar), .ZN(n166bar) );
  OR2_X1 U62 ( .A1(n221), .A2(b[6]), .ZN(n164) );
  AND2_X1 U62bar ( .A1(n221bar), .A2(bbar[6]), .ZN(n164bar) );
  OR2_X1 U63 ( .A1(n207), .A2(a[6]), .ZN(n165) );
  AND2_X1 U63bar ( .A1(n207bar), .A2(abar[6]), .ZN(n165bar) );
  AND2_X1 U64 ( .A1(n162), .A2(n161), .ZN(n163) );
  OR2_X1 U64bar ( .A1(n162bar), .A2(n161bar), .ZN(n163bar) );
  OR2_X1 U65 ( .A1(n197), .A2(d[6]), .ZN(n161) );
  AND2_X1 U65bar ( .A1(n197bar), .A2(dbar[6]), .ZN(n161bar) );
  OR2_X1 U66 ( .A1(n183), .A2(c[6]), .ZN(n162) );
  AND2_X1 U66bar ( .A1(n183bar), .A2(cbar[6]), .ZN(n162bar) );
  OR2_X1 U67 ( .A1(n160), .A2(n220), .ZN(y[5]) );
  AND2_X1 U67bar ( .A1(n160bar), .A2(n220bar), .ZN(ybar[5]) );
  OR2_X1 U68 ( .A1(n158), .A2(n196), .ZN(n159) );
  AND2_X1 U68bar ( .A1(n158bar), .A2(n196bar), .ZN(n159bar) );
  AND2_X1 U69 ( .A1(n196), .A2(n158), .ZN(n160) );
  OR2_X1 U69bar ( .A1(n196bar), .A2(n158bar), .ZN(n160bar) );
  AND2_X1 U70 ( .A1(n157), .A2(n156), .ZN(n158) );
  OR2_X1 U70bar ( .A1(n157bar), .A2(n156bar), .ZN(n158bar) );
  OR2_X1 U71 ( .A1(n219), .A2(b[5]), .ZN(n156) );
  AND2_X1 U71bar ( .A1(n219bar), .A2(bbar[5]), .ZN(n156bar) );
  OR2_X1 U72 ( .A1(n206), .A2(a[5]), .ZN(n157) );
  AND2_X1 U72bar ( .A1(n206bar), .A2(abar[5]), .ZN(n157bar) );
  AND2_X1 U73 ( .A1(n154), .A2(n153), .ZN(n155) );
  OR2_X1 U73bar ( .A1(n154bar), .A2(n153bar), .ZN(n155bar) );
  OR2_X1 U74 ( .A1(n195), .A2(d[5]), .ZN(n153) );
  AND2_X1 U74bar ( .A1(n195bar), .A2(dbar[5]), .ZN(n153bar) );
  OR2_X1 U75 ( .A1(n182), .A2(c[5]), .ZN(n154) );
  AND2_X1 U75bar ( .A1(n182bar), .A2(cbar[5]), .ZN(n154bar) );
  OR2_X1 U76 ( .A1(n152), .A2(n218), .ZN(y[4]) );
  AND2_X1 U76bar ( .A1(n152bar), .A2(n218bar), .ZN(ybar[4]) );
  OR2_X1 U77 ( .A1(n150), .A2(n194), .ZN(n151) );
  AND2_X1 U77bar ( .A1(n150bar), .A2(n194bar), .ZN(n151bar) );
  AND2_X1 U78 ( .A1(n194), .A2(n150), .ZN(n152) );
  OR2_X1 U78bar ( .A1(n194bar), .A2(n150bar), .ZN(n152bar) );
  AND2_X1 U79 ( .A1(n149), .A2(n148), .ZN(n150) );
  OR2_X1 U79bar ( .A1(n149bar), .A2(n148bar), .ZN(n150bar) );
  OR2_X1 U80 ( .A1(n217), .A2(b[4]), .ZN(n148) );
  AND2_X1 U80bar ( .A1(n217bar), .A2(bbar[4]), .ZN(n148bar) );
  OR2_X1 U81 ( .A1(n205), .A2(a[4]), .ZN(n149) );
  AND2_X1 U81bar ( .A1(n205bar), .A2(abar[4]), .ZN(n149bar) );
  AND2_X1 U82 ( .A1(n146), .A2(n145), .ZN(n147) );
  OR2_X1 U82bar ( .A1(n146bar), .A2(n145bar), .ZN(n147bar) );
  OR2_X1 U83 ( .A1(n193), .A2(d[4]), .ZN(n145) );
  AND2_X1 U83bar ( .A1(n193bar), .A2(dbar[4]), .ZN(n145bar) );
  OR2_X1 U84 ( .A1(n181), .A2(c[4]), .ZN(n146) );
  AND2_X1 U84bar ( .A1(n181bar), .A2(cbar[4]), .ZN(n146bar) );
  OR2_X1 U85 ( .A1(n144), .A2(n216), .ZN(y[3]) );
  AND2_X1 U85bar ( .A1(n144bar), .A2(n216bar), .ZN(ybar[3]) );
  OR2_X1 U86 ( .A1(n142), .A2(n192), .ZN(n143) );
  AND2_X1 U86bar ( .A1(n142bar), .A2(n192bar), .ZN(n143bar) );
  AND2_X1 U87 ( .A1(n192), .A2(n142), .ZN(n144) );
  OR2_X1 U87bar ( .A1(n192bar), .A2(n142bar), .ZN(n144bar) );
  AND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(n142) );
  OR2_X1 U88bar ( .A1(n141bar), .A2(n140bar), .ZN(n142bar) );
  OR2_X1 U89 ( .A1(n215), .A2(b[3]), .ZN(n140) );
  AND2_X1 U89bar ( .A1(n215bar), .A2(bbar[3]), .ZN(n140bar) );
  OR2_X1 U90 ( .A1(n204), .A2(a[3]), .ZN(n141) );
  AND2_X1 U90bar ( .A1(n204bar), .A2(abar[3]), .ZN(n141bar) );
  AND2_X1 U91 ( .A1(n138), .A2(n137), .ZN(n139) );
  OR2_X1 U91bar ( .A1(n138bar), .A2(n137bar), .ZN(n139bar) );
  OR2_X1 U92 ( .A1(n191), .A2(d[3]), .ZN(n137) );
  AND2_X1 U92bar ( .A1(n191bar), .A2(dbar[3]), .ZN(n137bar) );
  OR2_X1 U93 ( .A1(n180), .A2(c[3]), .ZN(n138) );
  AND2_X1 U93bar ( .A1(n180bar), .A2(cbar[3]), .ZN(n138bar) );
  OR2_X1 U94 ( .A1(n136), .A2(n214), .ZN(y[2]) );
  AND2_X1 U94bar ( .A1(n136bar), .A2(n214bar), .ZN(ybar[2]) );
  OR2_X1 U95 ( .A1(n134), .A2(n190), .ZN(n135) );
  AND2_X1 U95bar ( .A1(n134bar), .A2(n190bar), .ZN(n135bar) );
  AND2_X1 U96 ( .A1(n190), .A2(n134), .ZN(n136) );
  OR2_X1 U96bar ( .A1(n190bar), .A2(n134bar), .ZN(n136bar) );
  AND2_X1 U97 ( .A1(n133), .A2(n132), .ZN(n134) );
  OR2_X1 U97bar ( .A1(n133bar), .A2(n132bar), .ZN(n134bar) );
  OR2_X1 U98 ( .A1(n213), .A2(b[2]), .ZN(n132) );
  AND2_X1 U98bar ( .A1(n213bar), .A2(bbar[2]), .ZN(n132bar) );
  OR2_X1 U99 ( .A1(n203), .A2(a[2]), .ZN(n133) );
  AND2_X1 U99bar ( .A1(n203bar), .A2(abar[2]), .ZN(n133bar) );
  AND2_X1 U100 ( .A1(n130), .A2(n129), .ZN(n131) );
  OR2_X1 U100bar ( .A1(n130bar), .A2(n129bar), .ZN(n131bar) );
  OR2_X1 U101 ( .A1(n189), .A2(d[2]), .ZN(n129) );
  AND2_X1 U101bar ( .A1(n189bar), .A2(dbar[2]), .ZN(n129bar) );
  OR2_X1 U102 ( .A1(n179), .A2(c[2]), .ZN(n130) );
  AND2_X1 U102bar ( .A1(n179bar), .A2(cbar[2]), .ZN(n130bar) );
  OR2_X1 U103 ( .A1(n128), .A2(n212), .ZN(y[1]) );
  AND2_X1 U103bar ( .A1(n128bar), .A2(n212bar), .ZN(ybar[1]) );
  OR2_X1 U104 ( .A1(n126), .A2(n188), .ZN(n127) );
  AND2_X1 U104bar ( .A1(n126bar), .A2(n188bar), .ZN(n127bar) );
  AND2_X1 U105 ( .A1(n188), .A2(n126), .ZN(n128) );
  OR2_X1 U105bar ( .A1(n188bar), .A2(n126bar), .ZN(n128bar) );
  AND2_X1 U106 ( .A1(n125), .A2(n124), .ZN(n126) );
  OR2_X1 U106bar ( .A1(n125bar), .A2(n124bar), .ZN(n126bar) );
  OR2_X1 U107 ( .A1(n211), .A2(b[1]), .ZN(n124) );
  AND2_X1 U107bar ( .A1(n211bar), .A2(bbar[1]), .ZN(n124bar) );
  OR2_X1 U108 ( .A1(n202), .A2(a[1]), .ZN(n125) );
  AND2_X1 U108bar ( .A1(n202bar), .A2(abar[1]), .ZN(n125bar) );
  AND2_X1 U109 ( .A1(n122), .A2(n121), .ZN(n123) );
  OR2_X1 U109bar ( .A1(n122bar), .A2(n121bar), .ZN(n123bar) );
  OR2_X1 U110 ( .A1(n187), .A2(d[1]), .ZN(n121) );
  AND2_X1 U110bar ( .A1(n187bar), .A2(dbar[1]), .ZN(n121bar) );
  OR2_X1 U111 ( .A1(n178), .A2(c[1]), .ZN(n122) );
  AND2_X1 U111bar ( .A1(n178bar), .A2(cbar[1]), .ZN(n122bar) );
  OR2_X1 U112 ( .A1(n120), .A2(n210), .ZN(y[0]) );
  AND2_X1 U112bar ( .A1(n120bar), .A2(n210bar), .ZN(ybar[0]) );
  OR2_X1 U113 ( .A1(n118), .A2(n186), .ZN(n119) );
  AND2_X1 U113bar ( .A1(n118bar), .A2(n186bar), .ZN(n119bar) );
  AND2_X1 U114 ( .A1(n186), .A2(n118), .ZN(n120) );
  OR2_X1 U114bar ( .A1(n186bar), .A2(n118bar), .ZN(n120bar) );
  AND2_X1 U115 ( .A1(n117), .A2(n116), .ZN(n118) );
  OR2_X1 U115bar ( .A1(n117bar), .A2(n116bar), .ZN(n118bar) );
  OR2_X1 U116 ( .A1(n209), .A2(b[0]), .ZN(n116) );
  AND2_X1 U116bar ( .A1(n209bar), .A2(bbar[0]), .ZN(n116bar) );
  OR2_X1 U117 ( .A1(n201), .A2(a[0]), .ZN(n117) );
  AND2_X1 U117bar ( .A1(n201bar), .A2(abar[0]), .ZN(n117bar) );
  AND2_X1 U118 ( .A1(n114), .A2(n113), .ZN(n115) );
  OR2_X1 U118bar ( .A1(n114bar), .A2(n113bar), .ZN(n115bar) );
  OR2_X1 U119 ( .A1(n185), .A2(d[0]), .ZN(n113) );
  AND2_X1 U119bar ( .A1(n185bar), .A2(dbar[0]), .ZN(n113bar) );
  OR2_X1 U120 ( .A1(n177), .A2(c[0]), .ZN(n114) );
  AND2_X1 U120bar ( .A1(n177bar), .A2(cbar[0]), .ZN(n114bar) );
endmodule

module byteXor4_3 ( a, b, c, d, y );

  input wire [7:0] a;
  input wire [7:0] b;
  input wire [7:0] c;
  input wire [7:0] d;
  wire [7:0] abar;
  wire [7:0] bbar;
  wire [7:0] cbar;
  wire [7:0] dbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign cbar[0] = ~c[0];
  assign cbar[1] = ~c[1];
  assign cbar[2] = ~c[2];
  assign cbar[3] = ~c[3];
  assign cbar[4] = ~c[4];
  assign cbar[5] = ~c[5];
  assign cbar[6] = ~c[6];
  assign cbar[7] = ~c[7];
  assign dbar[0] = ~d[0];
  assign dbar[1] = ~d[1];
  assign dbar[2] = ~d[2];
  assign dbar[3] = ~d[3];
  assign dbar[4] = ~d[4];
  assign dbar[5] = ~d[5];
  assign dbar[6] = ~d[6];
  assign dbar[7] = ~d[7];
//input_done

  output wire [7:0] y;
  wire [7:0] ybar;
//output_done

  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n113bar;
  wire n114bar;
  wire n115bar;
  wire n116bar;
  wire n117bar;
  wire n118bar;
  wire n119bar;
  wire n120bar;
  wire n121bar;
  wire n122bar;
  wire n123bar;
  wire n124bar;
  wire n125bar;
  wire n126bar;
  wire n127bar;
  wire n128bar;
  wire n129bar;
  wire n130bar;
  wire n131bar;
  wire n132bar;
  wire n133bar;
  wire n134bar;
  wire n135bar;
  wire n136bar;
  wire n137bar;
  wire n138bar;
  wire n139bar;
  wire n140bar;
  wire n141bar;
  wire n142bar;
  wire n143bar;
  wire n144bar;
  wire n145bar;
  wire n146bar;
  wire n147bar;
  wire n148bar;
  wire n149bar;
  wire n150bar;
  wire n151bar;
  wire n152bar;
  wire n153bar;
  wire n154bar;
  wire n155bar;
  wire n156bar;
  wire n157bar;
  wire n158bar;
  wire n159bar;
  wire n160bar;
  wire n161bar;
  wire n162bar;
  wire n163bar;
  wire n164bar;
  wire n165bar;
  wire n166bar;
  wire n167bar;
  wire n168bar;
  wire n169bar;
  wire n170bar;
  wire n171bar;
  wire n172bar;
  wire n173bar;
  wire n174bar;
  wire n175bar;
  wire n176bar;
  wire n177bar;
  wire n178bar;
  wire n179bar;
  wire n180bar;
  wire n181bar;
  wire n182bar;
  wire n183bar;
  wire n184bar;
  wire n185bar;
  wire n186bar;
  wire n187bar;
  wire n188bar;
  wire n189bar;
  wire n190bar;
  wire n191bar;
  wire n192bar;
  wire n193bar;
  wire n194bar;
  wire n195bar;
  wire n196bar;
  wire n197bar;
  wire n198bar;
  wire n199bar;
  wire n200bar;
  wire n201bar;
  wire n202bar;
  wire n203bar;
  wire n204bar;
  wire n205bar;
  wire n206bar;
  wire n207bar;
  wire n208bar;
  wire n209bar;
  wire n210bar;
  wire n211bar;
  wire n212bar;
  wire n213bar;
  wire n214bar;
  wire n215bar;
  wire n216bar;
  wire n217bar;
  wire n218bar;
  wire n219bar;
  wire n220bar;
  wire n221bar;
  wire n222bar;
  wire n223bar;
  wire n224bar;
//wire_done

 //assign_done

  assign n224bar = n175;
  assign n224 = n175bar;
  assign n223bar = a[7];
  assign n223 = abar[7];
  assign n222bar = n167;
  assign n222 = n167bar;
  assign n221bar = a[6];
  assign n221 = abar[6];
  assign n220bar = n159;
  assign n220 = n159bar;
  assign n219bar = a[5];
  assign n219 = abar[5];
  assign n218bar = n151;
  assign n218 = n151bar;
  assign n217bar = a[4];
  assign n217 = abar[4];
  assign n216bar = n143;
  assign n216 = n143bar;
  assign n215bar = a[3];
  assign n215 = abar[3];
  assign n214bar = n135;
  assign n214 = n135bar;
  assign n213bar = a[2];
  assign n213 = abar[2];
  assign n212bar = n127;
  assign n212 = n127bar;
  assign n211bar = a[1];
  assign n211 = abar[1];
  assign n210bar = n119;
  assign n210 = n119bar;
  assign n209bar = a[0];
  assign n209 = abar[0];
  assign n208bar = b[7];
  assign n208 = bbar[7];
  assign n207bar = b[6];
  assign n207 = bbar[6];
  assign n206bar = b[5];
  assign n206 = bbar[5];
  assign n205bar = b[4];
  assign n205 = bbar[4];
  assign n204bar = b[3];
  assign n204 = bbar[3];
  assign n203bar = b[2];
  assign n203 = bbar[2];
  assign n202bar = b[1];
  assign n202 = bbar[1];
  assign n201bar = b[0];
  assign n201 = bbar[0];
  assign n200bar = n171;
  assign n200 = n171bar;
  assign n199bar = c[7];
  assign n199 = cbar[7];
  assign n198bar = n163;
  assign n198 = n163bar;
  assign n197bar = c[6];
  assign n197 = cbar[6];
  assign n196bar = n155;
  assign n196 = n155bar;
  assign n195bar = c[5];
  assign n195 = cbar[5];
  assign n194bar = n147;
  assign n194 = n147bar;
  assign n193bar = c[4];
  assign n193 = cbar[4];
  assign n192bar = n139;
  assign n192 = n139bar;
  assign n191bar = c[3];
  assign n191 = cbar[3];
  assign n190bar = n131;
  assign n190 = n131bar;
  assign n189bar = c[2];
  assign n189 = cbar[2];
  assign n188bar = n123;
  assign n188 = n123bar;
  assign n187bar = c[1];
  assign n187 = cbar[1];
  assign n186bar = n115;
  assign n186 = n115bar;
  assign n185bar = c[0];
  assign n185 = cbar[0];
  assign n184bar = d[7];
  assign n184 = dbar[7];
  assign n183bar = d[6];
  assign n183 = dbar[6];
  assign n182bar = d[5];
  assign n182 = dbar[5];
  assign n181bar = d[4];
  assign n181 = dbar[4];
  assign n180bar = d[3];
  assign n180 = dbar[3];
  assign n179bar = d[2];
  assign n179 = dbar[2];
  assign n178bar = d[1];
  assign n178 = dbar[1];
  assign n177bar = d[0];
  assign n177 = dbar[0];
  OR2_X1 U49 ( .A1(n176), .A2(n224), .ZN(y[7]) );
  AND2_X1 U49bar ( .A1(n176bar), .A2(n224bar), .ZN(ybar[7]) );
  OR2_X1 U50 ( .A1(n174), .A2(n200), .ZN(n175) );
  AND2_X1 U50bar ( .A1(n174bar), .A2(n200bar), .ZN(n175bar) );
  AND2_X1 U51 ( .A1(n200), .A2(n174), .ZN(n176) );
  OR2_X1 U51bar ( .A1(n200bar), .A2(n174bar), .ZN(n176bar) );
  AND2_X1 U52 ( .A1(n173), .A2(n172), .ZN(n174) );
  OR2_X1 U52bar ( .A1(n173bar), .A2(n172bar), .ZN(n174bar) );
  OR2_X1 U53 ( .A1(n223), .A2(b[7]), .ZN(n172) );
  AND2_X1 U53bar ( .A1(n223bar), .A2(bbar[7]), .ZN(n172bar) );
  OR2_X1 U54 ( .A1(n208), .A2(a[7]), .ZN(n173) );
  AND2_X1 U54bar ( .A1(n208bar), .A2(abar[7]), .ZN(n173bar) );
  AND2_X1 U55 ( .A1(n170), .A2(n169), .ZN(n171) );
  OR2_X1 U55bar ( .A1(n170bar), .A2(n169bar), .ZN(n171bar) );
  OR2_X1 U56 ( .A1(n199), .A2(d[7]), .ZN(n169) );
  AND2_X1 U56bar ( .A1(n199bar), .A2(dbar[7]), .ZN(n169bar) );
  OR2_X1 U57 ( .A1(n184), .A2(c[7]), .ZN(n170) );
  AND2_X1 U57bar ( .A1(n184bar), .A2(cbar[7]), .ZN(n170bar) );
  OR2_X1 U58 ( .A1(n168), .A2(n222), .ZN(y[6]) );
  AND2_X1 U58bar ( .A1(n168bar), .A2(n222bar), .ZN(ybar[6]) );
  OR2_X1 U59 ( .A1(n166), .A2(n198), .ZN(n167) );
  AND2_X1 U59bar ( .A1(n166bar), .A2(n198bar), .ZN(n167bar) );
  AND2_X1 U60 ( .A1(n198), .A2(n166), .ZN(n168) );
  OR2_X1 U60bar ( .A1(n198bar), .A2(n166bar), .ZN(n168bar) );
  AND2_X1 U61 ( .A1(n165), .A2(n164), .ZN(n166) );
  OR2_X1 U61bar ( .A1(n165bar), .A2(n164bar), .ZN(n166bar) );
  OR2_X1 U62 ( .A1(n221), .A2(b[6]), .ZN(n164) );
  AND2_X1 U62bar ( .A1(n221bar), .A2(bbar[6]), .ZN(n164bar) );
  OR2_X1 U63 ( .A1(n207), .A2(a[6]), .ZN(n165) );
  AND2_X1 U63bar ( .A1(n207bar), .A2(abar[6]), .ZN(n165bar) );
  AND2_X1 U64 ( .A1(n162), .A2(n161), .ZN(n163) );
  OR2_X1 U64bar ( .A1(n162bar), .A2(n161bar), .ZN(n163bar) );
  OR2_X1 U65 ( .A1(n197), .A2(d[6]), .ZN(n161) );
  AND2_X1 U65bar ( .A1(n197bar), .A2(dbar[6]), .ZN(n161bar) );
  OR2_X1 U66 ( .A1(n183), .A2(c[6]), .ZN(n162) );
  AND2_X1 U66bar ( .A1(n183bar), .A2(cbar[6]), .ZN(n162bar) );
  OR2_X1 U67 ( .A1(n160), .A2(n220), .ZN(y[5]) );
  AND2_X1 U67bar ( .A1(n160bar), .A2(n220bar), .ZN(ybar[5]) );
  OR2_X1 U68 ( .A1(n158), .A2(n196), .ZN(n159) );
  AND2_X1 U68bar ( .A1(n158bar), .A2(n196bar), .ZN(n159bar) );
  AND2_X1 U69 ( .A1(n196), .A2(n158), .ZN(n160) );
  OR2_X1 U69bar ( .A1(n196bar), .A2(n158bar), .ZN(n160bar) );
  AND2_X1 U70 ( .A1(n157), .A2(n156), .ZN(n158) );
  OR2_X1 U70bar ( .A1(n157bar), .A2(n156bar), .ZN(n158bar) );
  OR2_X1 U71 ( .A1(n219), .A2(b[5]), .ZN(n156) );
  AND2_X1 U71bar ( .A1(n219bar), .A2(bbar[5]), .ZN(n156bar) );
  OR2_X1 U72 ( .A1(n206), .A2(a[5]), .ZN(n157) );
  AND2_X1 U72bar ( .A1(n206bar), .A2(abar[5]), .ZN(n157bar) );
  AND2_X1 U73 ( .A1(n154), .A2(n153), .ZN(n155) );
  OR2_X1 U73bar ( .A1(n154bar), .A2(n153bar), .ZN(n155bar) );
  OR2_X1 U74 ( .A1(n195), .A2(d[5]), .ZN(n153) );
  AND2_X1 U74bar ( .A1(n195bar), .A2(dbar[5]), .ZN(n153bar) );
  OR2_X1 U75 ( .A1(n182), .A2(c[5]), .ZN(n154) );
  AND2_X1 U75bar ( .A1(n182bar), .A2(cbar[5]), .ZN(n154bar) );
  OR2_X1 U76 ( .A1(n152), .A2(n218), .ZN(y[4]) );
  AND2_X1 U76bar ( .A1(n152bar), .A2(n218bar), .ZN(ybar[4]) );
  OR2_X1 U77 ( .A1(n150), .A2(n194), .ZN(n151) );
  AND2_X1 U77bar ( .A1(n150bar), .A2(n194bar), .ZN(n151bar) );
  AND2_X1 U78 ( .A1(n194), .A2(n150), .ZN(n152) );
  OR2_X1 U78bar ( .A1(n194bar), .A2(n150bar), .ZN(n152bar) );
  AND2_X1 U79 ( .A1(n149), .A2(n148), .ZN(n150) );
  OR2_X1 U79bar ( .A1(n149bar), .A2(n148bar), .ZN(n150bar) );
  OR2_X1 U80 ( .A1(n217), .A2(b[4]), .ZN(n148) );
  AND2_X1 U80bar ( .A1(n217bar), .A2(bbar[4]), .ZN(n148bar) );
  OR2_X1 U81 ( .A1(n205), .A2(a[4]), .ZN(n149) );
  AND2_X1 U81bar ( .A1(n205bar), .A2(abar[4]), .ZN(n149bar) );
  AND2_X1 U82 ( .A1(n146), .A2(n145), .ZN(n147) );
  OR2_X1 U82bar ( .A1(n146bar), .A2(n145bar), .ZN(n147bar) );
  OR2_X1 U83 ( .A1(n193), .A2(d[4]), .ZN(n145) );
  AND2_X1 U83bar ( .A1(n193bar), .A2(dbar[4]), .ZN(n145bar) );
  OR2_X1 U84 ( .A1(n181), .A2(c[4]), .ZN(n146) );
  AND2_X1 U84bar ( .A1(n181bar), .A2(cbar[4]), .ZN(n146bar) );
  OR2_X1 U85 ( .A1(n144), .A2(n216), .ZN(y[3]) );
  AND2_X1 U85bar ( .A1(n144bar), .A2(n216bar), .ZN(ybar[3]) );
  OR2_X1 U86 ( .A1(n142), .A2(n192), .ZN(n143) );
  AND2_X1 U86bar ( .A1(n142bar), .A2(n192bar), .ZN(n143bar) );
  AND2_X1 U87 ( .A1(n192), .A2(n142), .ZN(n144) );
  OR2_X1 U87bar ( .A1(n192bar), .A2(n142bar), .ZN(n144bar) );
  AND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(n142) );
  OR2_X1 U88bar ( .A1(n141bar), .A2(n140bar), .ZN(n142bar) );
  OR2_X1 U89 ( .A1(n215), .A2(b[3]), .ZN(n140) );
  AND2_X1 U89bar ( .A1(n215bar), .A2(bbar[3]), .ZN(n140bar) );
  OR2_X1 U90 ( .A1(n204), .A2(a[3]), .ZN(n141) );
  AND2_X1 U90bar ( .A1(n204bar), .A2(abar[3]), .ZN(n141bar) );
  AND2_X1 U91 ( .A1(n138), .A2(n137), .ZN(n139) );
  OR2_X1 U91bar ( .A1(n138bar), .A2(n137bar), .ZN(n139bar) );
  OR2_X1 U92 ( .A1(n191), .A2(d[3]), .ZN(n137) );
  AND2_X1 U92bar ( .A1(n191bar), .A2(dbar[3]), .ZN(n137bar) );
  OR2_X1 U93 ( .A1(n180), .A2(c[3]), .ZN(n138) );
  AND2_X1 U93bar ( .A1(n180bar), .A2(cbar[3]), .ZN(n138bar) );
  OR2_X1 U94 ( .A1(n136), .A2(n214), .ZN(y[2]) );
  AND2_X1 U94bar ( .A1(n136bar), .A2(n214bar), .ZN(ybar[2]) );
  OR2_X1 U95 ( .A1(n134), .A2(n190), .ZN(n135) );
  AND2_X1 U95bar ( .A1(n134bar), .A2(n190bar), .ZN(n135bar) );
  AND2_X1 U96 ( .A1(n190), .A2(n134), .ZN(n136) );
  OR2_X1 U96bar ( .A1(n190bar), .A2(n134bar), .ZN(n136bar) );
  AND2_X1 U97 ( .A1(n133), .A2(n132), .ZN(n134) );
  OR2_X1 U97bar ( .A1(n133bar), .A2(n132bar), .ZN(n134bar) );
  OR2_X1 U98 ( .A1(n213), .A2(b[2]), .ZN(n132) );
  AND2_X1 U98bar ( .A1(n213bar), .A2(bbar[2]), .ZN(n132bar) );
  OR2_X1 U99 ( .A1(n203), .A2(a[2]), .ZN(n133) );
  AND2_X1 U99bar ( .A1(n203bar), .A2(abar[2]), .ZN(n133bar) );
  AND2_X1 U100 ( .A1(n130), .A2(n129), .ZN(n131) );
  OR2_X1 U100bar ( .A1(n130bar), .A2(n129bar), .ZN(n131bar) );
  OR2_X1 U101 ( .A1(n189), .A2(d[2]), .ZN(n129) );
  AND2_X1 U101bar ( .A1(n189bar), .A2(dbar[2]), .ZN(n129bar) );
  OR2_X1 U102 ( .A1(n179), .A2(c[2]), .ZN(n130) );
  AND2_X1 U102bar ( .A1(n179bar), .A2(cbar[2]), .ZN(n130bar) );
  OR2_X1 U103 ( .A1(n128), .A2(n212), .ZN(y[1]) );
  AND2_X1 U103bar ( .A1(n128bar), .A2(n212bar), .ZN(ybar[1]) );
  OR2_X1 U104 ( .A1(n126), .A2(n188), .ZN(n127) );
  AND2_X1 U104bar ( .A1(n126bar), .A2(n188bar), .ZN(n127bar) );
  AND2_X1 U105 ( .A1(n188), .A2(n126), .ZN(n128) );
  OR2_X1 U105bar ( .A1(n188bar), .A2(n126bar), .ZN(n128bar) );
  AND2_X1 U106 ( .A1(n125), .A2(n124), .ZN(n126) );
  OR2_X1 U106bar ( .A1(n125bar), .A2(n124bar), .ZN(n126bar) );
  OR2_X1 U107 ( .A1(n211), .A2(b[1]), .ZN(n124) );
  AND2_X1 U107bar ( .A1(n211bar), .A2(bbar[1]), .ZN(n124bar) );
  OR2_X1 U108 ( .A1(n202), .A2(a[1]), .ZN(n125) );
  AND2_X1 U108bar ( .A1(n202bar), .A2(abar[1]), .ZN(n125bar) );
  AND2_X1 U109 ( .A1(n122), .A2(n121), .ZN(n123) );
  OR2_X1 U109bar ( .A1(n122bar), .A2(n121bar), .ZN(n123bar) );
  OR2_X1 U110 ( .A1(n187), .A2(d[1]), .ZN(n121) );
  AND2_X1 U110bar ( .A1(n187bar), .A2(dbar[1]), .ZN(n121bar) );
  OR2_X1 U111 ( .A1(n178), .A2(c[1]), .ZN(n122) );
  AND2_X1 U111bar ( .A1(n178bar), .A2(cbar[1]), .ZN(n122bar) );
  OR2_X1 U112 ( .A1(n120), .A2(n210), .ZN(y[0]) );
  AND2_X1 U112bar ( .A1(n120bar), .A2(n210bar), .ZN(ybar[0]) );
  OR2_X1 U113 ( .A1(n118), .A2(n186), .ZN(n119) );
  AND2_X1 U113bar ( .A1(n118bar), .A2(n186bar), .ZN(n119bar) );
  AND2_X1 U114 ( .A1(n186), .A2(n118), .ZN(n120) );
  OR2_X1 U114bar ( .A1(n186bar), .A2(n118bar), .ZN(n120bar) );
  AND2_X1 U115 ( .A1(n117), .A2(n116), .ZN(n118) );
  OR2_X1 U115bar ( .A1(n117bar), .A2(n116bar), .ZN(n118bar) );
  OR2_X1 U116 ( .A1(n209), .A2(b[0]), .ZN(n116) );
  AND2_X1 U116bar ( .A1(n209bar), .A2(bbar[0]), .ZN(n116bar) );
  OR2_X1 U117 ( .A1(n201), .A2(a[0]), .ZN(n117) );
  AND2_X1 U117bar ( .A1(n201bar), .A2(abar[0]), .ZN(n117bar) );
  AND2_X1 U118 ( .A1(n114), .A2(n113), .ZN(n115) );
  OR2_X1 U118bar ( .A1(n114bar), .A2(n113bar), .ZN(n115bar) );
  OR2_X1 U119 ( .A1(n185), .A2(d[0]), .ZN(n113) );
  AND2_X1 U119bar ( .A1(n185bar), .A2(dbar[0]), .ZN(n113bar) );
  OR2_X1 U120 ( .A1(n177), .A2(c[0]), .ZN(n114) );
  AND2_X1 U120bar ( .A1(n177bar), .A2(cbar[0]), .ZN(n114bar) );
endmodule

module byteXor4_4 ( a, b, c, d, y );

  input wire [7:0] a;
  input wire [7:0] b;
  input wire [7:0] c;
  input wire [7:0] d;
  wire [7:0] abar;
  wire [7:0] bbar;
  wire [7:0] cbar;
  wire [7:0] dbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign cbar[0] = ~c[0];
  assign cbar[1] = ~c[1];
  assign cbar[2] = ~c[2];
  assign cbar[3] = ~c[3];
  assign cbar[4] = ~c[4];
  assign cbar[5] = ~c[5];
  assign cbar[6] = ~c[6];
  assign cbar[7] = ~c[7];
  assign dbar[0] = ~d[0];
  assign dbar[1] = ~d[1];
  assign dbar[2] = ~d[2];
  assign dbar[3] = ~d[3];
  assign dbar[4] = ~d[4];
  assign dbar[5] = ~d[5];
  assign dbar[6] = ~d[6];
  assign dbar[7] = ~d[7];
//input_done

  output wire [7:0] y;
  wire [7:0] ybar;
//output_done

  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n113bar;
  wire n114bar;
  wire n115bar;
  wire n116bar;
  wire n117bar;
  wire n118bar;
  wire n119bar;
  wire n120bar;
  wire n121bar;
  wire n122bar;
  wire n123bar;
  wire n124bar;
  wire n125bar;
  wire n126bar;
  wire n127bar;
  wire n128bar;
  wire n129bar;
  wire n130bar;
  wire n131bar;
  wire n132bar;
  wire n133bar;
  wire n134bar;
  wire n135bar;
  wire n136bar;
  wire n137bar;
  wire n138bar;
  wire n139bar;
  wire n140bar;
  wire n141bar;
  wire n142bar;
  wire n143bar;
  wire n144bar;
  wire n145bar;
  wire n146bar;
  wire n147bar;
  wire n148bar;
  wire n149bar;
  wire n150bar;
  wire n151bar;
  wire n152bar;
  wire n153bar;
  wire n154bar;
  wire n155bar;
  wire n156bar;
  wire n157bar;
  wire n158bar;
  wire n159bar;
  wire n160bar;
  wire n161bar;
  wire n162bar;
  wire n163bar;
  wire n164bar;
  wire n165bar;
  wire n166bar;
  wire n167bar;
  wire n168bar;
  wire n169bar;
  wire n170bar;
  wire n171bar;
  wire n172bar;
  wire n173bar;
  wire n174bar;
  wire n175bar;
  wire n176bar;
  wire n177bar;
  wire n178bar;
  wire n179bar;
  wire n180bar;
  wire n181bar;
  wire n182bar;
  wire n183bar;
  wire n184bar;
  wire n185bar;
  wire n186bar;
  wire n187bar;
  wire n188bar;
  wire n189bar;
  wire n190bar;
  wire n191bar;
  wire n192bar;
  wire n193bar;
  wire n194bar;
  wire n195bar;
  wire n196bar;
  wire n197bar;
  wire n198bar;
  wire n199bar;
  wire n200bar;
  wire n201bar;
  wire n202bar;
  wire n203bar;
  wire n204bar;
  wire n205bar;
  wire n206bar;
  wire n207bar;
  wire n208bar;
  wire n209bar;
  wire n210bar;
  wire n211bar;
  wire n212bar;
  wire n213bar;
  wire n214bar;
  wire n215bar;
  wire n216bar;
  wire n217bar;
  wire n218bar;
  wire n219bar;
  wire n220bar;
  wire n221bar;
  wire n222bar;
  wire n223bar;
  wire n224bar;
//wire_done

 //assign_done

  assign n224bar = n175;
  assign n224 = n175bar;
  assign n223bar = a[7];
  assign n223 = abar[7];
  assign n222bar = n167;
  assign n222 = n167bar;
  assign n221bar = a[6];
  assign n221 = abar[6];
  assign n220bar = n159;
  assign n220 = n159bar;
  assign n219bar = a[5];
  assign n219 = abar[5];
  assign n218bar = n151;
  assign n218 = n151bar;
  assign n217bar = a[4];
  assign n217 = abar[4];
  assign n216bar = n143;
  assign n216 = n143bar;
  assign n215bar = a[3];
  assign n215 = abar[3];
  assign n214bar = n135;
  assign n214 = n135bar;
  assign n213bar = a[2];
  assign n213 = abar[2];
  assign n212bar = n127;
  assign n212 = n127bar;
  assign n211bar = a[1];
  assign n211 = abar[1];
  assign n210bar = n119;
  assign n210 = n119bar;
  assign n209bar = a[0];
  assign n209 = abar[0];
  assign n208bar = b[7];
  assign n208 = bbar[7];
  assign n207bar = b[6];
  assign n207 = bbar[6];
  assign n206bar = b[5];
  assign n206 = bbar[5];
  assign n205bar = b[4];
  assign n205 = bbar[4];
  assign n204bar = b[3];
  assign n204 = bbar[3];
  assign n203bar = b[2];
  assign n203 = bbar[2];
  assign n202bar = b[1];
  assign n202 = bbar[1];
  assign n201bar = b[0];
  assign n201 = bbar[0];
  assign n200bar = n171;
  assign n200 = n171bar;
  assign n199bar = c[7];
  assign n199 = cbar[7];
  assign n198bar = n163;
  assign n198 = n163bar;
  assign n197bar = c[6];
  assign n197 = cbar[6];
  assign n196bar = n155;
  assign n196 = n155bar;
  assign n195bar = c[5];
  assign n195 = cbar[5];
  assign n194bar = n147;
  assign n194 = n147bar;
  assign n193bar = c[4];
  assign n193 = cbar[4];
  assign n192bar = n139;
  assign n192 = n139bar;
  assign n191bar = c[3];
  assign n191 = cbar[3];
  assign n190bar = n131;
  assign n190 = n131bar;
  assign n189bar = c[2];
  assign n189 = cbar[2];
  assign n188bar = n123;
  assign n188 = n123bar;
  assign n187bar = c[1];
  assign n187 = cbar[1];
  assign n186bar = n115;
  assign n186 = n115bar;
  assign n185bar = c[0];
  assign n185 = cbar[0];
  assign n184bar = d[7];
  assign n184 = dbar[7];
  assign n183bar = d[6];
  assign n183 = dbar[6];
  assign n182bar = d[5];
  assign n182 = dbar[5];
  assign n181bar = d[4];
  assign n181 = dbar[4];
  assign n180bar = d[3];
  assign n180 = dbar[3];
  assign n179bar = d[2];
  assign n179 = dbar[2];
  assign n178bar = d[1];
  assign n178 = dbar[1];
  assign n177bar = d[0];
  assign n177 = dbar[0];
  OR2_X1 U49 ( .A1(n176), .A2(n224), .ZN(y[7]) );
  AND2_X1 U49bar ( .A1(n176bar), .A2(n224bar), .ZN(ybar[7]) );
  OR2_X1 U50 ( .A1(n174), .A2(n200), .ZN(n175) );
  AND2_X1 U50bar ( .A1(n174bar), .A2(n200bar), .ZN(n175bar) );
  AND2_X1 U51 ( .A1(n200), .A2(n174), .ZN(n176) );
  OR2_X1 U51bar ( .A1(n200bar), .A2(n174bar), .ZN(n176bar) );
  AND2_X1 U52 ( .A1(n173), .A2(n172), .ZN(n174) );
  OR2_X1 U52bar ( .A1(n173bar), .A2(n172bar), .ZN(n174bar) );
  OR2_X1 U53 ( .A1(n223), .A2(b[7]), .ZN(n172) );
  AND2_X1 U53bar ( .A1(n223bar), .A2(bbar[7]), .ZN(n172bar) );
  OR2_X1 U54 ( .A1(n208), .A2(a[7]), .ZN(n173) );
  AND2_X1 U54bar ( .A1(n208bar), .A2(abar[7]), .ZN(n173bar) );
  AND2_X1 U55 ( .A1(n170), .A2(n169), .ZN(n171) );
  OR2_X1 U55bar ( .A1(n170bar), .A2(n169bar), .ZN(n171bar) );
  OR2_X1 U56 ( .A1(n199), .A2(d[7]), .ZN(n169) );
  AND2_X1 U56bar ( .A1(n199bar), .A2(dbar[7]), .ZN(n169bar) );
  OR2_X1 U57 ( .A1(n184), .A2(c[7]), .ZN(n170) );
  AND2_X1 U57bar ( .A1(n184bar), .A2(cbar[7]), .ZN(n170bar) );
  OR2_X1 U58 ( .A1(n168), .A2(n222), .ZN(y[6]) );
  AND2_X1 U58bar ( .A1(n168bar), .A2(n222bar), .ZN(ybar[6]) );
  OR2_X1 U59 ( .A1(n166), .A2(n198), .ZN(n167) );
  AND2_X1 U59bar ( .A1(n166bar), .A2(n198bar), .ZN(n167bar) );
  AND2_X1 U60 ( .A1(n198), .A2(n166), .ZN(n168) );
  OR2_X1 U60bar ( .A1(n198bar), .A2(n166bar), .ZN(n168bar) );
  AND2_X1 U61 ( .A1(n165), .A2(n164), .ZN(n166) );
  OR2_X1 U61bar ( .A1(n165bar), .A2(n164bar), .ZN(n166bar) );
  OR2_X1 U62 ( .A1(n221), .A2(b[6]), .ZN(n164) );
  AND2_X1 U62bar ( .A1(n221bar), .A2(bbar[6]), .ZN(n164bar) );
  OR2_X1 U63 ( .A1(n207), .A2(a[6]), .ZN(n165) );
  AND2_X1 U63bar ( .A1(n207bar), .A2(abar[6]), .ZN(n165bar) );
  AND2_X1 U64 ( .A1(n162), .A2(n161), .ZN(n163) );
  OR2_X1 U64bar ( .A1(n162bar), .A2(n161bar), .ZN(n163bar) );
  OR2_X1 U65 ( .A1(n197), .A2(d[6]), .ZN(n161) );
  AND2_X1 U65bar ( .A1(n197bar), .A2(dbar[6]), .ZN(n161bar) );
  OR2_X1 U66 ( .A1(n183), .A2(c[6]), .ZN(n162) );
  AND2_X1 U66bar ( .A1(n183bar), .A2(cbar[6]), .ZN(n162bar) );
  OR2_X1 U67 ( .A1(n160), .A2(n220), .ZN(y[5]) );
  AND2_X1 U67bar ( .A1(n160bar), .A2(n220bar), .ZN(ybar[5]) );
  OR2_X1 U68 ( .A1(n158), .A2(n196), .ZN(n159) );
  AND2_X1 U68bar ( .A1(n158bar), .A2(n196bar), .ZN(n159bar) );
  AND2_X1 U69 ( .A1(n196), .A2(n158), .ZN(n160) );
  OR2_X1 U69bar ( .A1(n196bar), .A2(n158bar), .ZN(n160bar) );
  AND2_X1 U70 ( .A1(n157), .A2(n156), .ZN(n158) );
  OR2_X1 U70bar ( .A1(n157bar), .A2(n156bar), .ZN(n158bar) );
  OR2_X1 U71 ( .A1(n219), .A2(b[5]), .ZN(n156) );
  AND2_X1 U71bar ( .A1(n219bar), .A2(bbar[5]), .ZN(n156bar) );
  OR2_X1 U72 ( .A1(n206), .A2(a[5]), .ZN(n157) );
  AND2_X1 U72bar ( .A1(n206bar), .A2(abar[5]), .ZN(n157bar) );
  AND2_X1 U73 ( .A1(n154), .A2(n153), .ZN(n155) );
  OR2_X1 U73bar ( .A1(n154bar), .A2(n153bar), .ZN(n155bar) );
  OR2_X1 U74 ( .A1(n195), .A2(d[5]), .ZN(n153) );
  AND2_X1 U74bar ( .A1(n195bar), .A2(dbar[5]), .ZN(n153bar) );
  OR2_X1 U75 ( .A1(n182), .A2(c[5]), .ZN(n154) );
  AND2_X1 U75bar ( .A1(n182bar), .A2(cbar[5]), .ZN(n154bar) );
  OR2_X1 U76 ( .A1(n152), .A2(n218), .ZN(y[4]) );
  AND2_X1 U76bar ( .A1(n152bar), .A2(n218bar), .ZN(ybar[4]) );
  OR2_X1 U77 ( .A1(n150), .A2(n194), .ZN(n151) );
  AND2_X1 U77bar ( .A1(n150bar), .A2(n194bar), .ZN(n151bar) );
  AND2_X1 U78 ( .A1(n194), .A2(n150), .ZN(n152) );
  OR2_X1 U78bar ( .A1(n194bar), .A2(n150bar), .ZN(n152bar) );
  AND2_X1 U79 ( .A1(n149), .A2(n148), .ZN(n150) );
  OR2_X1 U79bar ( .A1(n149bar), .A2(n148bar), .ZN(n150bar) );
  OR2_X1 U80 ( .A1(n217), .A2(b[4]), .ZN(n148) );
  AND2_X1 U80bar ( .A1(n217bar), .A2(bbar[4]), .ZN(n148bar) );
  OR2_X1 U81 ( .A1(n205), .A2(a[4]), .ZN(n149) );
  AND2_X1 U81bar ( .A1(n205bar), .A2(abar[4]), .ZN(n149bar) );
  AND2_X1 U82 ( .A1(n146), .A2(n145), .ZN(n147) );
  OR2_X1 U82bar ( .A1(n146bar), .A2(n145bar), .ZN(n147bar) );
  OR2_X1 U83 ( .A1(n193), .A2(d[4]), .ZN(n145) );
  AND2_X1 U83bar ( .A1(n193bar), .A2(dbar[4]), .ZN(n145bar) );
  OR2_X1 U84 ( .A1(n181), .A2(c[4]), .ZN(n146) );
  AND2_X1 U84bar ( .A1(n181bar), .A2(cbar[4]), .ZN(n146bar) );
  OR2_X1 U85 ( .A1(n144), .A2(n216), .ZN(y[3]) );
  AND2_X1 U85bar ( .A1(n144bar), .A2(n216bar), .ZN(ybar[3]) );
  OR2_X1 U86 ( .A1(n142), .A2(n192), .ZN(n143) );
  AND2_X1 U86bar ( .A1(n142bar), .A2(n192bar), .ZN(n143bar) );
  AND2_X1 U87 ( .A1(n192), .A2(n142), .ZN(n144) );
  OR2_X1 U87bar ( .A1(n192bar), .A2(n142bar), .ZN(n144bar) );
  AND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(n142) );
  OR2_X1 U88bar ( .A1(n141bar), .A2(n140bar), .ZN(n142bar) );
  OR2_X1 U89 ( .A1(n215), .A2(b[3]), .ZN(n140) );
  AND2_X1 U89bar ( .A1(n215bar), .A2(bbar[3]), .ZN(n140bar) );
  OR2_X1 U90 ( .A1(n204), .A2(a[3]), .ZN(n141) );
  AND2_X1 U90bar ( .A1(n204bar), .A2(abar[3]), .ZN(n141bar) );
  AND2_X1 U91 ( .A1(n138), .A2(n137), .ZN(n139) );
  OR2_X1 U91bar ( .A1(n138bar), .A2(n137bar), .ZN(n139bar) );
  OR2_X1 U92 ( .A1(n191), .A2(d[3]), .ZN(n137) );
  AND2_X1 U92bar ( .A1(n191bar), .A2(dbar[3]), .ZN(n137bar) );
  OR2_X1 U93 ( .A1(n180), .A2(c[3]), .ZN(n138) );
  AND2_X1 U93bar ( .A1(n180bar), .A2(cbar[3]), .ZN(n138bar) );
  OR2_X1 U94 ( .A1(n136), .A2(n214), .ZN(y[2]) );
  AND2_X1 U94bar ( .A1(n136bar), .A2(n214bar), .ZN(ybar[2]) );
  OR2_X1 U95 ( .A1(n134), .A2(n190), .ZN(n135) );
  AND2_X1 U95bar ( .A1(n134bar), .A2(n190bar), .ZN(n135bar) );
  AND2_X1 U96 ( .A1(n190), .A2(n134), .ZN(n136) );
  OR2_X1 U96bar ( .A1(n190bar), .A2(n134bar), .ZN(n136bar) );
  AND2_X1 U97 ( .A1(n133), .A2(n132), .ZN(n134) );
  OR2_X1 U97bar ( .A1(n133bar), .A2(n132bar), .ZN(n134bar) );
  OR2_X1 U98 ( .A1(n213), .A2(b[2]), .ZN(n132) );
  AND2_X1 U98bar ( .A1(n213bar), .A2(bbar[2]), .ZN(n132bar) );
  OR2_X1 U99 ( .A1(n203), .A2(a[2]), .ZN(n133) );
  AND2_X1 U99bar ( .A1(n203bar), .A2(abar[2]), .ZN(n133bar) );
  AND2_X1 U100 ( .A1(n130), .A2(n129), .ZN(n131) );
  OR2_X1 U100bar ( .A1(n130bar), .A2(n129bar), .ZN(n131bar) );
  OR2_X1 U101 ( .A1(n189), .A2(d[2]), .ZN(n129) );
  AND2_X1 U101bar ( .A1(n189bar), .A2(dbar[2]), .ZN(n129bar) );
  OR2_X1 U102 ( .A1(n179), .A2(c[2]), .ZN(n130) );
  AND2_X1 U102bar ( .A1(n179bar), .A2(cbar[2]), .ZN(n130bar) );
  OR2_X1 U103 ( .A1(n128), .A2(n212), .ZN(y[1]) );
  AND2_X1 U103bar ( .A1(n128bar), .A2(n212bar), .ZN(ybar[1]) );
  OR2_X1 U104 ( .A1(n126), .A2(n188), .ZN(n127) );
  AND2_X1 U104bar ( .A1(n126bar), .A2(n188bar), .ZN(n127bar) );
  AND2_X1 U105 ( .A1(n188), .A2(n126), .ZN(n128) );
  OR2_X1 U105bar ( .A1(n188bar), .A2(n126bar), .ZN(n128bar) );
  AND2_X1 U106 ( .A1(n125), .A2(n124), .ZN(n126) );
  OR2_X1 U106bar ( .A1(n125bar), .A2(n124bar), .ZN(n126bar) );
  OR2_X1 U107 ( .A1(n211), .A2(b[1]), .ZN(n124) );
  AND2_X1 U107bar ( .A1(n211bar), .A2(bbar[1]), .ZN(n124bar) );
  OR2_X1 U108 ( .A1(n202), .A2(a[1]), .ZN(n125) );
  AND2_X1 U108bar ( .A1(n202bar), .A2(abar[1]), .ZN(n125bar) );
  AND2_X1 U109 ( .A1(n122), .A2(n121), .ZN(n123) );
  OR2_X1 U109bar ( .A1(n122bar), .A2(n121bar), .ZN(n123bar) );
  OR2_X1 U110 ( .A1(n187), .A2(d[1]), .ZN(n121) );
  AND2_X1 U110bar ( .A1(n187bar), .A2(dbar[1]), .ZN(n121bar) );
  OR2_X1 U111 ( .A1(n178), .A2(c[1]), .ZN(n122) );
  AND2_X1 U111bar ( .A1(n178bar), .A2(cbar[1]), .ZN(n122bar) );
  OR2_X1 U112 ( .A1(n120), .A2(n210), .ZN(y[0]) );
  AND2_X1 U112bar ( .A1(n120bar), .A2(n210bar), .ZN(ybar[0]) );
  OR2_X1 U113 ( .A1(n118), .A2(n186), .ZN(n119) );
  AND2_X1 U113bar ( .A1(n118bar), .A2(n186bar), .ZN(n119bar) );
  AND2_X1 U114 ( .A1(n186), .A2(n118), .ZN(n120) );
  OR2_X1 U114bar ( .A1(n186bar), .A2(n118bar), .ZN(n120bar) );
  AND2_X1 U115 ( .A1(n117), .A2(n116), .ZN(n118) );
  OR2_X1 U115bar ( .A1(n117bar), .A2(n116bar), .ZN(n118bar) );
  OR2_X1 U116 ( .A1(n209), .A2(b[0]), .ZN(n116) );
  AND2_X1 U116bar ( .A1(n209bar), .A2(bbar[0]), .ZN(n116bar) );
  OR2_X1 U117 ( .A1(n201), .A2(a[0]), .ZN(n117) );
  AND2_X1 U117bar ( .A1(n201bar), .A2(abar[0]), .ZN(n117bar) );
  AND2_X1 U118 ( .A1(n114), .A2(n113), .ZN(n115) );
  OR2_X1 U118bar ( .A1(n114bar), .A2(n113bar), .ZN(n115bar) );
  OR2_X1 U119 ( .A1(n185), .A2(d[0]), .ZN(n113) );
  AND2_X1 U119bar ( .A1(n185bar), .A2(dbar[0]), .ZN(n113bar) );
  OR2_X1 U120 ( .A1(n177), .A2(c[0]), .ZN(n114) );
  AND2_X1 U120bar ( .A1(n177bar), .A2(cbar[0]), .ZN(n114bar) );
endmodule

module mixCol_1 ( in, out );

  input wire [31:0] in;
//input_done

  output wire [31:0] out;
//output_done

  wire [7:0] b0_s2;
  wire [7:0] b1_s2;
  wire [7:0] b2_s2;
  wire [7:0] b3_s2;
  wire [7:0] b0_s3;
  wire [7:0] b1_s3;
  wire [7:0] b2_s3;
  wire [7:0] b3_s3;
//wire_done

 //assign_done

  scale2_4 b0_scale2 ( .in(in[31:24]), .out(b0_s2) );
  scale2_3 b1_scale2 ( .in(in[23:16]), .out(b1_s2) );
  scale2_2 b2_scale2 ( .in(in[15:8]), .out(b2_s2) );
  scale2_1 b3_scale2 ( .in(in[7:0]), .out(b3_s2) );
  byteXor_5 b0_scale3 ( .a(in[31:24]), .b(b0_s2), .y(b0_s3) );
  byteXor_4 b1_scale3 ( .a(in[23:16]), .b(b1_s2), .y(b1_s3) );
  byteXor_3 b2_scale3 ( .a(in[15:8]), .b(b2_s2), .y(b2_s3) );
  byteXor_2 b3_scale3 ( .a(in[7:0]), .b(b3_s2), .y(b3_s3) );
  byteXor4_4 out0 ( .a(b0_s2), .b(b1_s3), .c(in[15:8]), .d(in[7:0]), .y(
        out[31:24]) );
  byteXor4_3 out1 ( .a(in[31:24]), .b(b1_s2), .c(b2_s3), .d(in[7:0]), .y(
        out[23:16]) );
  byteXor4_2 out2 ( .a(in[31:24]), .b(in[23:16]), .c(b2_s2), .d(b3_s3), .y(
        out[15:8]) );
  byteXor4_1 out3 ( .a(b0_s3), .b(in[23:16]), .c(in[15:8]), .d(b3_s2), .y(
        out[7:0]) );
endmodule

module scale2_5 ( in, out );

  input wire [7:0] in;
  wire [7:0] inbar;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
//input_done

  output wire [7:0] out;
  wire [7:0] outbar;
//output_done

  wire in_0;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_1;
  wire in_7;
  wire n11;
  wire n12;
  wire n13;
  wire n14;
  wire n15;
  wire n16;
  wire n17;
  wire n18;
  wire n19;
  wire n20;
  wire in_0bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_1bar;
  wire in_7bar;
  wire n11bar;
  wire n12bar;
  wire n13bar;
  wire n14bar;
  wire n15bar;
  wire n16bar;
  wire n17bar;
  wire n18bar;
  wire n19bar;
  wire n20bar;
//wire_done

  assign in_0 = in[0];
  assign out[7] = in_6;
  assign in_6  = in[6];
  assign out[6] = in_5;
  assign in_5  = in[5];
  assign out[5] = in_4;
  assign in_4  = in[4];
  assign out[2] = in_1;
  assign in_1  = in[1];
  assign out[0] = in_7;
  assign in_7  = in[7];
  assign in_0bar = inbar[0];
  assign outbar[7] = in_6bar;
  assign in_6bar = inbar[6];
  assign outbar[6] = in_5bar;
  assign in_5bar = inbar[5];
  assign outbar[5] = in_4bar;
  assign in_4bar = inbar[4];
  assign outbar[2] = in_1bar;
  assign in_1bar = inbar[1];
  assign outbar[0] = in_7bar;
  assign in_7bar = inbar[7];
//assign_done

  assign n20bar = in_7;
  assign n20 = in_7bar;
  assign n19bar = in[3];
  assign n19 = inbar[3];
  assign n18bar = in[2];
  assign n18 = inbar[2];
  assign n17bar = in_0;
  assign n17 = in_0bar;
  OR2_X1 U5 ( .A1(n16), .A2(n15), .ZN(out[4]) );
  AND2_X1 U5bar ( .A1(n16bar), .A2(n15bar), .ZN(outbar[4]) );
  AND2_X1 U6 ( .A1(in[3]), .A2(n20), .ZN(n15) );
  OR2_X1 U6bar ( .A1(inbar[3]), .A2(n20bar), .ZN(n15bar) );
  AND2_X1 U7 ( .A1(in_7), .A2(n19), .ZN(n16) );
  OR2_X1 U7bar ( .A1(in_7bar), .A2(n19bar), .ZN(n16bar) );
  OR2_X1 U8 ( .A1(n14), .A2(n13), .ZN(out[3]) );
  AND2_X1 U8bar ( .A1(n14bar), .A2(n13bar), .ZN(outbar[3]) );
  AND2_X1 U9 ( .A1(in[2]), .A2(n20), .ZN(n13) );
  OR2_X1 U9bar ( .A1(inbar[2]), .A2(n20bar), .ZN(n13bar) );
  AND2_X1 U10 ( .A1(in_7), .A2(n18), .ZN(n14) );
  OR2_X1 U10bar ( .A1(in_7bar), .A2(n18bar), .ZN(n14bar) );
  OR2_X1 U11 ( .A1(n12), .A2(n11), .ZN(out[1]) );
  AND2_X1 U11bar ( .A1(n12bar), .A2(n11bar), .ZN(outbar[1]) );
  AND2_X1 U12 ( .A1(in_0), .A2(n20), .ZN(n11) );
  OR2_X1 U12bar ( .A1(in_0bar), .A2(n20bar), .ZN(n11bar) );
  AND2_X1 U13 ( .A1(in_7), .A2(n17), .ZN(n12) );
  OR2_X1 U13bar ( .A1(in_7bar), .A2(n17bar), .ZN(n12bar) );
endmodule

module scale2_6 ( in, out );

  input wire [7:0] in;
  wire [7:0] inbar;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
//input_done

  output wire [7:0] out;
  wire [7:0] outbar;
//output_done

  wire in_0;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_1;
  wire in_7;
  wire n11;
  wire n12;
  wire n13;
  wire n14;
  wire n15;
  wire n16;
  wire n17;
  wire n18;
  wire n19;
  wire n20;
  wire in_0bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_1bar;
  wire in_7bar;
  wire n11bar;
  wire n12bar;
  wire n13bar;
  wire n14bar;
  wire n15bar;
  wire n16bar;
  wire n17bar;
  wire n18bar;
  wire n19bar;
  wire n20bar;
//wire_done

  assign in_0 = in[0];
  assign out[7] = in_6;
  assign in_6  = in[6];
  assign out[6] = in_5;
  assign in_5  = in[5];
  assign out[5] = in_4;
  assign in_4  = in[4];
  assign out[2] = in_1;
  assign in_1  = in[1];
  assign out[0] = in_7;
  assign in_7  = in[7];
  assign in_0bar = inbar[0];
  assign outbar[7] = in_6bar;
  assign in_6bar = inbar[6];
  assign outbar[6] = in_5bar;
  assign in_5bar = inbar[5];
  assign outbar[5] = in_4bar;
  assign in_4bar = inbar[4];
  assign outbar[2] = in_1bar;
  assign in_1bar = inbar[1];
  assign outbar[0] = in_7bar;
  assign in_7bar = inbar[7];
//assign_done

  assign n20bar = in_7;
  assign n20 = in_7bar;
  assign n19bar = in[3];
  assign n19 = inbar[3];
  assign n18bar = in[2];
  assign n18 = inbar[2];
  assign n17bar = in_0;
  assign n17 = in_0bar;
  OR2_X1 U5 ( .A1(n16), .A2(n15), .ZN(out[4]) );
  AND2_X1 U5bar ( .A1(n16bar), .A2(n15bar), .ZN(outbar[4]) );
  AND2_X1 U6 ( .A1(in[3]), .A2(n20), .ZN(n15) );
  OR2_X1 U6bar ( .A1(inbar[3]), .A2(n20bar), .ZN(n15bar) );
  AND2_X1 U7 ( .A1(in_7), .A2(n19), .ZN(n16) );
  OR2_X1 U7bar ( .A1(in_7bar), .A2(n19bar), .ZN(n16bar) );
  OR2_X1 U8 ( .A1(n14), .A2(n13), .ZN(out[3]) );
  AND2_X1 U8bar ( .A1(n14bar), .A2(n13bar), .ZN(outbar[3]) );
  AND2_X1 U9 ( .A1(in[2]), .A2(n20), .ZN(n13) );
  OR2_X1 U9bar ( .A1(inbar[2]), .A2(n20bar), .ZN(n13bar) );
  AND2_X1 U10 ( .A1(in_7), .A2(n18), .ZN(n14) );
  OR2_X1 U10bar ( .A1(in_7bar), .A2(n18bar), .ZN(n14bar) );
  OR2_X1 U11 ( .A1(n12), .A2(n11), .ZN(out[1]) );
  AND2_X1 U11bar ( .A1(n12bar), .A2(n11bar), .ZN(outbar[1]) );
  AND2_X1 U12 ( .A1(in_0), .A2(n20), .ZN(n11) );
  OR2_X1 U12bar ( .A1(in_0bar), .A2(n20bar), .ZN(n11bar) );
  AND2_X1 U13 ( .A1(in_7), .A2(n17), .ZN(n12) );
  OR2_X1 U13bar ( .A1(in_7bar), .A2(n17bar), .ZN(n12bar) );
endmodule

module scale2_7 ( in, out );

  input wire [7:0] in;
  wire [7:0] inbar;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
//input_done

  output wire [7:0] out;
  wire [7:0] outbar;
//output_done

  wire in_0;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_1;
  wire in_7;
  wire n11;
  wire n12;
  wire n13;
  wire n14;
  wire n15;
  wire n16;
  wire n17;
  wire n18;
  wire n19;
  wire n20;
  wire in_0bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_1bar;
  wire in_7bar;
  wire n11bar;
  wire n12bar;
  wire n13bar;
  wire n14bar;
  wire n15bar;
  wire n16bar;
  wire n17bar;
  wire n18bar;
  wire n19bar;
  wire n20bar;
//wire_done

  assign in_0 = in[0];
  assign out[7] = in_6;
  assign in_6  = in[6];
  assign out[6] = in_5;
  assign in_5  = in[5];
  assign out[5] = in_4;
  assign in_4  = in[4];
  assign out[2] = in_1;
  assign in_1  = in[1];
  assign out[0] = in_7;
  assign in_7  = in[7];
  assign in_0bar = inbar[0];
  assign outbar[7] = in_6bar;
  assign in_6bar = inbar[6];
  assign outbar[6] = in_5bar;
  assign in_5bar = inbar[5];
  assign outbar[5] = in_4bar;
  assign in_4bar = inbar[4];
  assign outbar[2] = in_1bar;
  assign in_1bar = inbar[1];
  assign outbar[0] = in_7bar;
  assign in_7bar = inbar[7];
//assign_done

  assign n20bar = in_7;
  assign n20 = in_7bar;
  assign n19bar = in[3];
  assign n19 = inbar[3];
  assign n18bar = in[2];
  assign n18 = inbar[2];
  assign n17bar = in_0;
  assign n17 = in_0bar;
  OR2_X1 U5 ( .A1(n16), .A2(n15), .ZN(out[4]) );
  AND2_X1 U5bar ( .A1(n16bar), .A2(n15bar), .ZN(outbar[4]) );
  AND2_X1 U6 ( .A1(in[3]), .A2(n20), .ZN(n15) );
  OR2_X1 U6bar ( .A1(inbar[3]), .A2(n20bar), .ZN(n15bar) );
  AND2_X1 U7 ( .A1(in_7), .A2(n19), .ZN(n16) );
  OR2_X1 U7bar ( .A1(in_7bar), .A2(n19bar), .ZN(n16bar) );
  OR2_X1 U8 ( .A1(n14), .A2(n13), .ZN(out[3]) );
  AND2_X1 U8bar ( .A1(n14bar), .A2(n13bar), .ZN(outbar[3]) );
  AND2_X1 U9 ( .A1(in[2]), .A2(n20), .ZN(n13) );
  OR2_X1 U9bar ( .A1(inbar[2]), .A2(n20bar), .ZN(n13bar) );
  AND2_X1 U10 ( .A1(in_7), .A2(n18), .ZN(n14) );
  OR2_X1 U10bar ( .A1(in_7bar), .A2(n18bar), .ZN(n14bar) );
  OR2_X1 U11 ( .A1(n12), .A2(n11), .ZN(out[1]) );
  AND2_X1 U11bar ( .A1(n12bar), .A2(n11bar), .ZN(outbar[1]) );
  AND2_X1 U12 ( .A1(in_0), .A2(n20), .ZN(n11) );
  OR2_X1 U12bar ( .A1(in_0bar), .A2(n20bar), .ZN(n11bar) );
  AND2_X1 U13 ( .A1(in_7), .A2(n17), .ZN(n12) );
  OR2_X1 U13bar ( .A1(in_7bar), .A2(n17bar), .ZN(n12bar) );
endmodule

module scale2_8 ( in, out );

  input wire [7:0] in;
  wire [7:0] inbar;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
//input_done

  output wire [7:0] out;
  wire [7:0] outbar;
//output_done

  wire in_0;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_1;
  wire in_7;
  wire n11;
  wire n12;
  wire n13;
  wire n14;
  wire n15;
  wire n16;
  wire n17;
  wire n18;
  wire n19;
  wire n20;
  wire in_0bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_1bar;
  wire in_7bar;
  wire n11bar;
  wire n12bar;
  wire n13bar;
  wire n14bar;
  wire n15bar;
  wire n16bar;
  wire n17bar;
  wire n18bar;
  wire n19bar;
  wire n20bar;
//wire_done

  assign in_0 = in[0];
  assign out[7] = in_6;
  assign in_6  = in[6];
  assign out[6] = in_5;
  assign in_5  = in[5];
  assign out[5] = in_4;
  assign in_4  = in[4];
  assign out[2] = in_1;
  assign in_1  = in[1];
  assign out[0] = in_7;
  assign in_7  = in[7];
  assign in_0bar = inbar[0];
  assign outbar[7] = in_6bar;
  assign in_6bar = inbar[6];
  assign outbar[6] = in_5bar;
  assign in_5bar = inbar[5];
  assign outbar[5] = in_4bar;
  assign in_4bar = inbar[4];
  assign outbar[2] = in_1bar;
  assign in_1bar = inbar[1];
  assign outbar[0] = in_7bar;
  assign in_7bar = inbar[7];
//assign_done

  assign n20bar = in_7;
  assign n20 = in_7bar;
  assign n19bar = in[3];
  assign n19 = inbar[3];
  assign n18bar = in[2];
  assign n18 = inbar[2];
  assign n17bar = in_0;
  assign n17 = in_0bar;
  OR2_X1 U5 ( .A1(n16), .A2(n15), .ZN(out[4]) );
  AND2_X1 U5bar ( .A1(n16bar), .A2(n15bar), .ZN(outbar[4]) );
  AND2_X1 U6 ( .A1(in[3]), .A2(n20), .ZN(n15) );
  OR2_X1 U6bar ( .A1(inbar[3]), .A2(n20bar), .ZN(n15bar) );
  AND2_X1 U7 ( .A1(in_7), .A2(n19), .ZN(n16) );
  OR2_X1 U7bar ( .A1(in_7bar), .A2(n19bar), .ZN(n16bar) );
  OR2_X1 U8 ( .A1(n14), .A2(n13), .ZN(out[3]) );
  AND2_X1 U8bar ( .A1(n14bar), .A2(n13bar), .ZN(outbar[3]) );
  AND2_X1 U9 ( .A1(in[2]), .A2(n20), .ZN(n13) );
  OR2_X1 U9bar ( .A1(inbar[2]), .A2(n20bar), .ZN(n13bar) );
  AND2_X1 U10 ( .A1(in_7), .A2(n18), .ZN(n14) );
  OR2_X1 U10bar ( .A1(in_7bar), .A2(n18bar), .ZN(n14bar) );
  OR2_X1 U11 ( .A1(n12), .A2(n11), .ZN(out[1]) );
  AND2_X1 U11bar ( .A1(n12bar), .A2(n11bar), .ZN(outbar[1]) );
  AND2_X1 U12 ( .A1(in_0), .A2(n20), .ZN(n11) );
  OR2_X1 U12bar ( .A1(in_0bar), .A2(n20bar), .ZN(n11bar) );
  AND2_X1 U13 ( .A1(in_7), .A2(n17), .ZN(n12) );
  OR2_X1 U13bar ( .A1(in_7bar), .A2(n17bar), .ZN(n12bar) );
endmodule

module byteXor_6 ( a, b, y );

  input wire [7:0] a;
  input wire [7:0] b;
  wire [7:0] abar;
  wire [7:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
//input_done

  output wire [7:0] y;
  wire [7:0] ybar;
//output_done

  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n33bar;
  wire n34bar;
  wire n35bar;
  wire n36bar;
  wire n37bar;
  wire n38bar;
  wire n39bar;
  wire n40bar;
  wire n41bar;
  wire n42bar;
  wire n43bar;
  wire n44bar;
  wire n45bar;
  wire n46bar;
  wire n47bar;
  wire n48bar;
  wire n49bar;
  wire n50bar;
  wire n51bar;
  wire n52bar;
  wire n53bar;
  wire n54bar;
  wire n55bar;
  wire n56bar;
  wire n57bar;
  wire n58bar;
  wire n59bar;
  wire n60bar;
  wire n61bar;
  wire n62bar;
  wire n63bar;
  wire n64bar;
//wire_done

 //assign_done

  assign n64bar = n47;
  assign n64 = n47bar;
  assign n63bar = a[7];
  assign n63 = abar[7];
  assign n62bar = n45;
  assign n62 = n45bar;
  assign n61bar = a[6];
  assign n61 = abar[6];
  assign n60bar = n43;
  assign n60 = n43bar;
  assign n59bar = a[5];
  assign n59 = abar[5];
  assign n58bar = n41;
  assign n58 = n41bar;
  assign n57bar = a[4];
  assign n57 = abar[4];
  assign n56bar = n39;
  assign n56 = n39bar;
  assign n55bar = a[3];
  assign n55 = abar[3];
  assign n54bar = n37;
  assign n54 = n37bar;
  assign n53bar = a[2];
  assign n53 = abar[2];
  assign n52bar = n35;
  assign n52 = n35bar;
  assign n51bar = a[1];
  assign n51 = abar[1];
  assign n50bar = n33;
  assign n50 = n33bar;
  assign n49bar = a[0];
  assign n49 = abar[0];
  OR2_X1 U17 ( .A1(n48), .A2(n64), .ZN(y[7]) );
  AND2_X1 U17bar ( .A1(n48bar), .A2(n64bar), .ZN(ybar[7]) );
  OR2_X1 U18 ( .A1(n63), .A2(b[7]), .ZN(n47) );
  AND2_X1 U18bar ( .A1(n63bar), .A2(bbar[7]), .ZN(n47bar) );
  AND2_X1 U19 ( .A1(b[7]), .A2(n63), .ZN(n48) );
  OR2_X1 U19bar ( .A1(bbar[7]), .A2(n63bar), .ZN(n48bar) );
  OR2_X1 U20 ( .A1(n46), .A2(n62), .ZN(y[6]) );
  AND2_X1 U20bar ( .A1(n46bar), .A2(n62bar), .ZN(ybar[6]) );
  OR2_X1 U21 ( .A1(n61), .A2(b[6]), .ZN(n45) );
  AND2_X1 U21bar ( .A1(n61bar), .A2(bbar[6]), .ZN(n45bar) );
  AND2_X1 U22 ( .A1(b[6]), .A2(n61), .ZN(n46) );
  OR2_X1 U22bar ( .A1(bbar[6]), .A2(n61bar), .ZN(n46bar) );
  OR2_X1 U23 ( .A1(n44), .A2(n60), .ZN(y[5]) );
  AND2_X1 U23bar ( .A1(n44bar), .A2(n60bar), .ZN(ybar[5]) );
  OR2_X1 U24 ( .A1(n59), .A2(b[5]), .ZN(n43) );
  AND2_X1 U24bar ( .A1(n59bar), .A2(bbar[5]), .ZN(n43bar) );
  AND2_X1 U25 ( .A1(b[5]), .A2(n59), .ZN(n44) );
  OR2_X1 U25bar ( .A1(bbar[5]), .A2(n59bar), .ZN(n44bar) );
  OR2_X1 U26 ( .A1(n42), .A2(n58), .ZN(y[4]) );
  AND2_X1 U26bar ( .A1(n42bar), .A2(n58bar), .ZN(ybar[4]) );
  OR2_X1 U27 ( .A1(n57), .A2(b[4]), .ZN(n41) );
  AND2_X1 U27bar ( .A1(n57bar), .A2(bbar[4]), .ZN(n41bar) );
  AND2_X1 U28 ( .A1(b[4]), .A2(n57), .ZN(n42) );
  OR2_X1 U28bar ( .A1(bbar[4]), .A2(n57bar), .ZN(n42bar) );
  OR2_X1 U29 ( .A1(n40), .A2(n56), .ZN(y[3]) );
  AND2_X1 U29bar ( .A1(n40bar), .A2(n56bar), .ZN(ybar[3]) );
  OR2_X1 U30 ( .A1(n55), .A2(b[3]), .ZN(n39) );
  AND2_X1 U30bar ( .A1(n55bar), .A2(bbar[3]), .ZN(n39bar) );
  AND2_X1 U31 ( .A1(b[3]), .A2(n55), .ZN(n40) );
  OR2_X1 U31bar ( .A1(bbar[3]), .A2(n55bar), .ZN(n40bar) );
  OR2_X1 U32 ( .A1(n38), .A2(n54), .ZN(y[2]) );
  AND2_X1 U32bar ( .A1(n38bar), .A2(n54bar), .ZN(ybar[2]) );
  OR2_X1 U33 ( .A1(n53), .A2(b[2]), .ZN(n37) );
  AND2_X1 U33bar ( .A1(n53bar), .A2(bbar[2]), .ZN(n37bar) );
  AND2_X1 U34 ( .A1(b[2]), .A2(n53), .ZN(n38) );
  OR2_X1 U34bar ( .A1(bbar[2]), .A2(n53bar), .ZN(n38bar) );
  OR2_X1 U35 ( .A1(n36), .A2(n52), .ZN(y[1]) );
  AND2_X1 U35bar ( .A1(n36bar), .A2(n52bar), .ZN(ybar[1]) );
  OR2_X1 U36 ( .A1(n51), .A2(b[1]), .ZN(n35) );
  AND2_X1 U36bar ( .A1(n51bar), .A2(bbar[1]), .ZN(n35bar) );
  AND2_X1 U37 ( .A1(b[1]), .A2(n51), .ZN(n36) );
  OR2_X1 U37bar ( .A1(bbar[1]), .A2(n51bar), .ZN(n36bar) );
  OR2_X1 U38 ( .A1(n34), .A2(n50), .ZN(y[0]) );
  AND2_X1 U38bar ( .A1(n34bar), .A2(n50bar), .ZN(ybar[0]) );
  OR2_X1 U39 ( .A1(n49), .A2(b[0]), .ZN(n33) );
  AND2_X1 U39bar ( .A1(n49bar), .A2(bbar[0]), .ZN(n33bar) );
  AND2_X1 U40 ( .A1(b[0]), .A2(n49), .ZN(n34) );
  OR2_X1 U40bar ( .A1(bbar[0]), .A2(n49bar), .ZN(n34bar) );
endmodule

module byteXor_7 ( a, b, y );

  input wire [7:0] a;
  input wire [7:0] b;
  wire [7:0] abar;
  wire [7:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
//input_done

  output wire [7:0] y;
  wire [7:0] ybar;
//output_done

  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n33bar;
  wire n34bar;
  wire n35bar;
  wire n36bar;
  wire n37bar;
  wire n38bar;
  wire n39bar;
  wire n40bar;
  wire n41bar;
  wire n42bar;
  wire n43bar;
  wire n44bar;
  wire n45bar;
  wire n46bar;
  wire n47bar;
  wire n48bar;
  wire n49bar;
  wire n50bar;
  wire n51bar;
  wire n52bar;
  wire n53bar;
  wire n54bar;
  wire n55bar;
  wire n56bar;
  wire n57bar;
  wire n58bar;
  wire n59bar;
  wire n60bar;
  wire n61bar;
  wire n62bar;
  wire n63bar;
  wire n64bar;
//wire_done

 //assign_done

  assign n64bar = n47;
  assign n64 = n47bar;
  assign n63bar = a[7];
  assign n63 = abar[7];
  assign n62bar = n45;
  assign n62 = n45bar;
  assign n61bar = a[6];
  assign n61 = abar[6];
  assign n60bar = n43;
  assign n60 = n43bar;
  assign n59bar = a[5];
  assign n59 = abar[5];
  assign n58bar = n41;
  assign n58 = n41bar;
  assign n57bar = a[4];
  assign n57 = abar[4];
  assign n56bar = n39;
  assign n56 = n39bar;
  assign n55bar = a[3];
  assign n55 = abar[3];
  assign n54bar = n37;
  assign n54 = n37bar;
  assign n53bar = a[2];
  assign n53 = abar[2];
  assign n52bar = n35;
  assign n52 = n35bar;
  assign n51bar = a[1];
  assign n51 = abar[1];
  assign n50bar = n33;
  assign n50 = n33bar;
  assign n49bar = a[0];
  assign n49 = abar[0];
  OR2_X1 U17 ( .A1(n48), .A2(n64), .ZN(y[7]) );
  AND2_X1 U17bar ( .A1(n48bar), .A2(n64bar), .ZN(ybar[7]) );
  OR2_X1 U18 ( .A1(n63), .A2(b[7]), .ZN(n47) );
  AND2_X1 U18bar ( .A1(n63bar), .A2(bbar[7]), .ZN(n47bar) );
  AND2_X1 U19 ( .A1(b[7]), .A2(n63), .ZN(n48) );
  OR2_X1 U19bar ( .A1(bbar[7]), .A2(n63bar), .ZN(n48bar) );
  OR2_X1 U20 ( .A1(n46), .A2(n62), .ZN(y[6]) );
  AND2_X1 U20bar ( .A1(n46bar), .A2(n62bar), .ZN(ybar[6]) );
  OR2_X1 U21 ( .A1(n61), .A2(b[6]), .ZN(n45) );
  AND2_X1 U21bar ( .A1(n61bar), .A2(bbar[6]), .ZN(n45bar) );
  AND2_X1 U22 ( .A1(b[6]), .A2(n61), .ZN(n46) );
  OR2_X1 U22bar ( .A1(bbar[6]), .A2(n61bar), .ZN(n46bar) );
  OR2_X1 U23 ( .A1(n44), .A2(n60), .ZN(y[5]) );
  AND2_X1 U23bar ( .A1(n44bar), .A2(n60bar), .ZN(ybar[5]) );
  OR2_X1 U24 ( .A1(n59), .A2(b[5]), .ZN(n43) );
  AND2_X1 U24bar ( .A1(n59bar), .A2(bbar[5]), .ZN(n43bar) );
  AND2_X1 U25 ( .A1(b[5]), .A2(n59), .ZN(n44) );
  OR2_X1 U25bar ( .A1(bbar[5]), .A2(n59bar), .ZN(n44bar) );
  OR2_X1 U26 ( .A1(n42), .A2(n58), .ZN(y[4]) );
  AND2_X1 U26bar ( .A1(n42bar), .A2(n58bar), .ZN(ybar[4]) );
  OR2_X1 U27 ( .A1(n57), .A2(b[4]), .ZN(n41) );
  AND2_X1 U27bar ( .A1(n57bar), .A2(bbar[4]), .ZN(n41bar) );
  AND2_X1 U28 ( .A1(b[4]), .A2(n57), .ZN(n42) );
  OR2_X1 U28bar ( .A1(bbar[4]), .A2(n57bar), .ZN(n42bar) );
  OR2_X1 U29 ( .A1(n40), .A2(n56), .ZN(y[3]) );
  AND2_X1 U29bar ( .A1(n40bar), .A2(n56bar), .ZN(ybar[3]) );
  OR2_X1 U30 ( .A1(n55), .A2(b[3]), .ZN(n39) );
  AND2_X1 U30bar ( .A1(n55bar), .A2(bbar[3]), .ZN(n39bar) );
  AND2_X1 U31 ( .A1(b[3]), .A2(n55), .ZN(n40) );
  OR2_X1 U31bar ( .A1(bbar[3]), .A2(n55bar), .ZN(n40bar) );
  OR2_X1 U32 ( .A1(n38), .A2(n54), .ZN(y[2]) );
  AND2_X1 U32bar ( .A1(n38bar), .A2(n54bar), .ZN(ybar[2]) );
  OR2_X1 U33 ( .A1(n53), .A2(b[2]), .ZN(n37) );
  AND2_X1 U33bar ( .A1(n53bar), .A2(bbar[2]), .ZN(n37bar) );
  AND2_X1 U34 ( .A1(b[2]), .A2(n53), .ZN(n38) );
  OR2_X1 U34bar ( .A1(bbar[2]), .A2(n53bar), .ZN(n38bar) );
  OR2_X1 U35 ( .A1(n36), .A2(n52), .ZN(y[1]) );
  AND2_X1 U35bar ( .A1(n36bar), .A2(n52bar), .ZN(ybar[1]) );
  OR2_X1 U36 ( .A1(n51), .A2(b[1]), .ZN(n35) );
  AND2_X1 U36bar ( .A1(n51bar), .A2(bbar[1]), .ZN(n35bar) );
  AND2_X1 U37 ( .A1(b[1]), .A2(n51), .ZN(n36) );
  OR2_X1 U37bar ( .A1(bbar[1]), .A2(n51bar), .ZN(n36bar) );
  OR2_X1 U38 ( .A1(n34), .A2(n50), .ZN(y[0]) );
  AND2_X1 U38bar ( .A1(n34bar), .A2(n50bar), .ZN(ybar[0]) );
  OR2_X1 U39 ( .A1(n49), .A2(b[0]), .ZN(n33) );
  AND2_X1 U39bar ( .A1(n49bar), .A2(bbar[0]), .ZN(n33bar) );
  AND2_X1 U40 ( .A1(b[0]), .A2(n49), .ZN(n34) );
  OR2_X1 U40bar ( .A1(bbar[0]), .A2(n49bar), .ZN(n34bar) );
endmodule

module byteXor_8 ( a, b, y );

  input wire [7:0] a;
  input wire [7:0] b;
  wire [7:0] abar;
  wire [7:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
//input_done

  output wire [7:0] y;
  wire [7:0] ybar;
//output_done

  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n33bar;
  wire n34bar;
  wire n35bar;
  wire n36bar;
  wire n37bar;
  wire n38bar;
  wire n39bar;
  wire n40bar;
  wire n41bar;
  wire n42bar;
  wire n43bar;
  wire n44bar;
  wire n45bar;
  wire n46bar;
  wire n47bar;
  wire n48bar;
  wire n49bar;
  wire n50bar;
  wire n51bar;
  wire n52bar;
  wire n53bar;
  wire n54bar;
  wire n55bar;
  wire n56bar;
  wire n57bar;
  wire n58bar;
  wire n59bar;
  wire n60bar;
  wire n61bar;
  wire n62bar;
  wire n63bar;
  wire n64bar;
//wire_done

 //assign_done

  assign n64bar = n47;
  assign n64 = n47bar;
  assign n63bar = a[7];
  assign n63 = abar[7];
  assign n62bar = n45;
  assign n62 = n45bar;
  assign n61bar = a[6];
  assign n61 = abar[6];
  assign n60bar = n43;
  assign n60 = n43bar;
  assign n59bar = a[5];
  assign n59 = abar[5];
  assign n58bar = n41;
  assign n58 = n41bar;
  assign n57bar = a[4];
  assign n57 = abar[4];
  assign n56bar = n39;
  assign n56 = n39bar;
  assign n55bar = a[3];
  assign n55 = abar[3];
  assign n54bar = n37;
  assign n54 = n37bar;
  assign n53bar = a[2];
  assign n53 = abar[2];
  assign n52bar = n35;
  assign n52 = n35bar;
  assign n51bar = a[1];
  assign n51 = abar[1];
  assign n50bar = n33;
  assign n50 = n33bar;
  assign n49bar = a[0];
  assign n49 = abar[0];
  OR2_X1 U17 ( .A1(n48), .A2(n64), .ZN(y[7]) );
  AND2_X1 U17bar ( .A1(n48bar), .A2(n64bar), .ZN(ybar[7]) );
  OR2_X1 U18 ( .A1(n63), .A2(b[7]), .ZN(n47) );
  AND2_X1 U18bar ( .A1(n63bar), .A2(bbar[7]), .ZN(n47bar) );
  AND2_X1 U19 ( .A1(b[7]), .A2(n63), .ZN(n48) );
  OR2_X1 U19bar ( .A1(bbar[7]), .A2(n63bar), .ZN(n48bar) );
  OR2_X1 U20 ( .A1(n46), .A2(n62), .ZN(y[6]) );
  AND2_X1 U20bar ( .A1(n46bar), .A2(n62bar), .ZN(ybar[6]) );
  OR2_X1 U21 ( .A1(n61), .A2(b[6]), .ZN(n45) );
  AND2_X1 U21bar ( .A1(n61bar), .A2(bbar[6]), .ZN(n45bar) );
  AND2_X1 U22 ( .A1(b[6]), .A2(n61), .ZN(n46) );
  OR2_X1 U22bar ( .A1(bbar[6]), .A2(n61bar), .ZN(n46bar) );
  OR2_X1 U23 ( .A1(n44), .A2(n60), .ZN(y[5]) );
  AND2_X1 U23bar ( .A1(n44bar), .A2(n60bar), .ZN(ybar[5]) );
  OR2_X1 U24 ( .A1(n59), .A2(b[5]), .ZN(n43) );
  AND2_X1 U24bar ( .A1(n59bar), .A2(bbar[5]), .ZN(n43bar) );
  AND2_X1 U25 ( .A1(b[5]), .A2(n59), .ZN(n44) );
  OR2_X1 U25bar ( .A1(bbar[5]), .A2(n59bar), .ZN(n44bar) );
  OR2_X1 U26 ( .A1(n42), .A2(n58), .ZN(y[4]) );
  AND2_X1 U26bar ( .A1(n42bar), .A2(n58bar), .ZN(ybar[4]) );
  OR2_X1 U27 ( .A1(n57), .A2(b[4]), .ZN(n41) );
  AND2_X1 U27bar ( .A1(n57bar), .A2(bbar[4]), .ZN(n41bar) );
  AND2_X1 U28 ( .A1(b[4]), .A2(n57), .ZN(n42) );
  OR2_X1 U28bar ( .A1(bbar[4]), .A2(n57bar), .ZN(n42bar) );
  OR2_X1 U29 ( .A1(n40), .A2(n56), .ZN(y[3]) );
  AND2_X1 U29bar ( .A1(n40bar), .A2(n56bar), .ZN(ybar[3]) );
  OR2_X1 U30 ( .A1(n55), .A2(b[3]), .ZN(n39) );
  AND2_X1 U30bar ( .A1(n55bar), .A2(bbar[3]), .ZN(n39bar) );
  AND2_X1 U31 ( .A1(b[3]), .A2(n55), .ZN(n40) );
  OR2_X1 U31bar ( .A1(bbar[3]), .A2(n55bar), .ZN(n40bar) );
  OR2_X1 U32 ( .A1(n38), .A2(n54), .ZN(y[2]) );
  AND2_X1 U32bar ( .A1(n38bar), .A2(n54bar), .ZN(ybar[2]) );
  OR2_X1 U33 ( .A1(n53), .A2(b[2]), .ZN(n37) );
  AND2_X1 U33bar ( .A1(n53bar), .A2(bbar[2]), .ZN(n37bar) );
  AND2_X1 U34 ( .A1(b[2]), .A2(n53), .ZN(n38) );
  OR2_X1 U34bar ( .A1(bbar[2]), .A2(n53bar), .ZN(n38bar) );
  OR2_X1 U35 ( .A1(n36), .A2(n52), .ZN(y[1]) );
  AND2_X1 U35bar ( .A1(n36bar), .A2(n52bar), .ZN(ybar[1]) );
  OR2_X1 U36 ( .A1(n51), .A2(b[1]), .ZN(n35) );
  AND2_X1 U36bar ( .A1(n51bar), .A2(bbar[1]), .ZN(n35bar) );
  AND2_X1 U37 ( .A1(b[1]), .A2(n51), .ZN(n36) );
  OR2_X1 U37bar ( .A1(bbar[1]), .A2(n51bar), .ZN(n36bar) );
  OR2_X1 U38 ( .A1(n34), .A2(n50), .ZN(y[0]) );
  AND2_X1 U38bar ( .A1(n34bar), .A2(n50bar), .ZN(ybar[0]) );
  OR2_X1 U39 ( .A1(n49), .A2(b[0]), .ZN(n33) );
  AND2_X1 U39bar ( .A1(n49bar), .A2(bbar[0]), .ZN(n33bar) );
  AND2_X1 U40 ( .A1(b[0]), .A2(n49), .ZN(n34) );
  OR2_X1 U40bar ( .A1(bbar[0]), .A2(n49bar), .ZN(n34bar) );
endmodule

module byteXor_9 ( a, b, y );

  input wire [7:0] a;
  input wire [7:0] b;
  wire [7:0] abar;
  wire [7:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
//input_done

  output wire [7:0] y;
  wire [7:0] ybar;
//output_done

  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n33bar;
  wire n34bar;
  wire n35bar;
  wire n36bar;
  wire n37bar;
  wire n38bar;
  wire n39bar;
  wire n40bar;
  wire n41bar;
  wire n42bar;
  wire n43bar;
  wire n44bar;
  wire n45bar;
  wire n46bar;
  wire n47bar;
  wire n48bar;
  wire n49bar;
  wire n50bar;
  wire n51bar;
  wire n52bar;
  wire n53bar;
  wire n54bar;
  wire n55bar;
  wire n56bar;
  wire n57bar;
  wire n58bar;
  wire n59bar;
  wire n60bar;
  wire n61bar;
  wire n62bar;
  wire n63bar;
  wire n64bar;
//wire_done

 //assign_done

  assign n64bar = n47;
  assign n64 = n47bar;
  assign n63bar = a[7];
  assign n63 = abar[7];
  assign n62bar = n45;
  assign n62 = n45bar;
  assign n61bar = a[6];
  assign n61 = abar[6];
  assign n60bar = n43;
  assign n60 = n43bar;
  assign n59bar = a[5];
  assign n59 = abar[5];
  assign n58bar = n41;
  assign n58 = n41bar;
  assign n57bar = a[4];
  assign n57 = abar[4];
  assign n56bar = n39;
  assign n56 = n39bar;
  assign n55bar = a[3];
  assign n55 = abar[3];
  assign n54bar = n37;
  assign n54 = n37bar;
  assign n53bar = a[2];
  assign n53 = abar[2];
  assign n52bar = n35;
  assign n52 = n35bar;
  assign n51bar = a[1];
  assign n51 = abar[1];
  assign n50bar = n33;
  assign n50 = n33bar;
  assign n49bar = a[0];
  assign n49 = abar[0];
  OR2_X1 U17 ( .A1(n48), .A2(n64), .ZN(y[7]) );
  AND2_X1 U17bar ( .A1(n48bar), .A2(n64bar), .ZN(ybar[7]) );
  OR2_X1 U18 ( .A1(n63), .A2(b[7]), .ZN(n47) );
  AND2_X1 U18bar ( .A1(n63bar), .A2(bbar[7]), .ZN(n47bar) );
  AND2_X1 U19 ( .A1(b[7]), .A2(n63), .ZN(n48) );
  OR2_X1 U19bar ( .A1(bbar[7]), .A2(n63bar), .ZN(n48bar) );
  OR2_X1 U20 ( .A1(n46), .A2(n62), .ZN(y[6]) );
  AND2_X1 U20bar ( .A1(n46bar), .A2(n62bar), .ZN(ybar[6]) );
  OR2_X1 U21 ( .A1(n61), .A2(b[6]), .ZN(n45) );
  AND2_X1 U21bar ( .A1(n61bar), .A2(bbar[6]), .ZN(n45bar) );
  AND2_X1 U22 ( .A1(b[6]), .A2(n61), .ZN(n46) );
  OR2_X1 U22bar ( .A1(bbar[6]), .A2(n61bar), .ZN(n46bar) );
  OR2_X1 U23 ( .A1(n44), .A2(n60), .ZN(y[5]) );
  AND2_X1 U23bar ( .A1(n44bar), .A2(n60bar), .ZN(ybar[5]) );
  OR2_X1 U24 ( .A1(n59), .A2(b[5]), .ZN(n43) );
  AND2_X1 U24bar ( .A1(n59bar), .A2(bbar[5]), .ZN(n43bar) );
  AND2_X1 U25 ( .A1(b[5]), .A2(n59), .ZN(n44) );
  OR2_X1 U25bar ( .A1(bbar[5]), .A2(n59bar), .ZN(n44bar) );
  OR2_X1 U26 ( .A1(n42), .A2(n58), .ZN(y[4]) );
  AND2_X1 U26bar ( .A1(n42bar), .A2(n58bar), .ZN(ybar[4]) );
  OR2_X1 U27 ( .A1(n57), .A2(b[4]), .ZN(n41) );
  AND2_X1 U27bar ( .A1(n57bar), .A2(bbar[4]), .ZN(n41bar) );
  AND2_X1 U28 ( .A1(b[4]), .A2(n57), .ZN(n42) );
  OR2_X1 U28bar ( .A1(bbar[4]), .A2(n57bar), .ZN(n42bar) );
  OR2_X1 U29 ( .A1(n40), .A2(n56), .ZN(y[3]) );
  AND2_X1 U29bar ( .A1(n40bar), .A2(n56bar), .ZN(ybar[3]) );
  OR2_X1 U30 ( .A1(n55), .A2(b[3]), .ZN(n39) );
  AND2_X1 U30bar ( .A1(n55bar), .A2(bbar[3]), .ZN(n39bar) );
  AND2_X1 U31 ( .A1(b[3]), .A2(n55), .ZN(n40) );
  OR2_X1 U31bar ( .A1(bbar[3]), .A2(n55bar), .ZN(n40bar) );
  OR2_X1 U32 ( .A1(n38), .A2(n54), .ZN(y[2]) );
  AND2_X1 U32bar ( .A1(n38bar), .A2(n54bar), .ZN(ybar[2]) );
  OR2_X1 U33 ( .A1(n53), .A2(b[2]), .ZN(n37) );
  AND2_X1 U33bar ( .A1(n53bar), .A2(bbar[2]), .ZN(n37bar) );
  AND2_X1 U34 ( .A1(b[2]), .A2(n53), .ZN(n38) );
  OR2_X1 U34bar ( .A1(bbar[2]), .A2(n53bar), .ZN(n38bar) );
  OR2_X1 U35 ( .A1(n36), .A2(n52), .ZN(y[1]) );
  AND2_X1 U35bar ( .A1(n36bar), .A2(n52bar), .ZN(ybar[1]) );
  OR2_X1 U36 ( .A1(n51), .A2(b[1]), .ZN(n35) );
  AND2_X1 U36bar ( .A1(n51bar), .A2(bbar[1]), .ZN(n35bar) );
  AND2_X1 U37 ( .A1(b[1]), .A2(n51), .ZN(n36) );
  OR2_X1 U37bar ( .A1(bbar[1]), .A2(n51bar), .ZN(n36bar) );
  OR2_X1 U38 ( .A1(n34), .A2(n50), .ZN(y[0]) );
  AND2_X1 U38bar ( .A1(n34bar), .A2(n50bar), .ZN(ybar[0]) );
  OR2_X1 U39 ( .A1(n49), .A2(b[0]), .ZN(n33) );
  AND2_X1 U39bar ( .A1(n49bar), .A2(bbar[0]), .ZN(n33bar) );
  AND2_X1 U40 ( .A1(b[0]), .A2(n49), .ZN(n34) );
  OR2_X1 U40bar ( .A1(bbar[0]), .A2(n49bar), .ZN(n34bar) );
endmodule

module byteXor4_5 ( a, b, c, d, y );

  input wire [7:0] a;
  input wire [7:0] b;
  input wire [7:0] c;
  input wire [7:0] d;
  wire [7:0] abar;
  wire [7:0] bbar;
  wire [7:0] cbar;
  wire [7:0] dbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign cbar[0] = ~c[0];
  assign cbar[1] = ~c[1];
  assign cbar[2] = ~c[2];
  assign cbar[3] = ~c[3];
  assign cbar[4] = ~c[4];
  assign cbar[5] = ~c[5];
  assign cbar[6] = ~c[6];
  assign cbar[7] = ~c[7];
  assign dbar[0] = ~d[0];
  assign dbar[1] = ~d[1];
  assign dbar[2] = ~d[2];
  assign dbar[3] = ~d[3];
  assign dbar[4] = ~d[4];
  assign dbar[5] = ~d[5];
  assign dbar[6] = ~d[6];
  assign dbar[7] = ~d[7];
//input_done

  output wire [7:0] y;
  wire [7:0] ybar;
//output_done

  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n113bar;
  wire n114bar;
  wire n115bar;
  wire n116bar;
  wire n117bar;
  wire n118bar;
  wire n119bar;
  wire n120bar;
  wire n121bar;
  wire n122bar;
  wire n123bar;
  wire n124bar;
  wire n125bar;
  wire n126bar;
  wire n127bar;
  wire n128bar;
  wire n129bar;
  wire n130bar;
  wire n131bar;
  wire n132bar;
  wire n133bar;
  wire n134bar;
  wire n135bar;
  wire n136bar;
  wire n137bar;
  wire n138bar;
  wire n139bar;
  wire n140bar;
  wire n141bar;
  wire n142bar;
  wire n143bar;
  wire n144bar;
  wire n145bar;
  wire n146bar;
  wire n147bar;
  wire n148bar;
  wire n149bar;
  wire n150bar;
  wire n151bar;
  wire n152bar;
  wire n153bar;
  wire n154bar;
  wire n155bar;
  wire n156bar;
  wire n157bar;
  wire n158bar;
  wire n159bar;
  wire n160bar;
  wire n161bar;
  wire n162bar;
  wire n163bar;
  wire n164bar;
  wire n165bar;
  wire n166bar;
  wire n167bar;
  wire n168bar;
  wire n169bar;
  wire n170bar;
  wire n171bar;
  wire n172bar;
  wire n173bar;
  wire n174bar;
  wire n175bar;
  wire n176bar;
  wire n177bar;
  wire n178bar;
  wire n179bar;
  wire n180bar;
  wire n181bar;
  wire n182bar;
  wire n183bar;
  wire n184bar;
  wire n185bar;
  wire n186bar;
  wire n187bar;
  wire n188bar;
  wire n189bar;
  wire n190bar;
  wire n191bar;
  wire n192bar;
  wire n193bar;
  wire n194bar;
  wire n195bar;
  wire n196bar;
  wire n197bar;
  wire n198bar;
  wire n199bar;
  wire n200bar;
  wire n201bar;
  wire n202bar;
  wire n203bar;
  wire n204bar;
  wire n205bar;
  wire n206bar;
  wire n207bar;
  wire n208bar;
  wire n209bar;
  wire n210bar;
  wire n211bar;
  wire n212bar;
  wire n213bar;
  wire n214bar;
  wire n215bar;
  wire n216bar;
  wire n217bar;
  wire n218bar;
  wire n219bar;
  wire n220bar;
  wire n221bar;
  wire n222bar;
  wire n223bar;
  wire n224bar;
//wire_done

 //assign_done

  assign n224bar = n175;
  assign n224 = n175bar;
  assign n223bar = a[7];
  assign n223 = abar[7];
  assign n222bar = n167;
  assign n222 = n167bar;
  assign n221bar = a[6];
  assign n221 = abar[6];
  assign n220bar = n159;
  assign n220 = n159bar;
  assign n219bar = a[5];
  assign n219 = abar[5];
  assign n218bar = n151;
  assign n218 = n151bar;
  assign n217bar = a[4];
  assign n217 = abar[4];
  assign n216bar = n143;
  assign n216 = n143bar;
  assign n215bar = a[3];
  assign n215 = abar[3];
  assign n214bar = n135;
  assign n214 = n135bar;
  assign n213bar = a[2];
  assign n213 = abar[2];
  assign n212bar = n127;
  assign n212 = n127bar;
  assign n211bar = a[1];
  assign n211 = abar[1];
  assign n210bar = n119;
  assign n210 = n119bar;
  assign n209bar = a[0];
  assign n209 = abar[0];
  assign n208bar = b[7];
  assign n208 = bbar[7];
  assign n207bar = b[6];
  assign n207 = bbar[6];
  assign n206bar = b[5];
  assign n206 = bbar[5];
  assign n205bar = b[4];
  assign n205 = bbar[4];
  assign n204bar = b[3];
  assign n204 = bbar[3];
  assign n203bar = b[2];
  assign n203 = bbar[2];
  assign n202bar = b[1];
  assign n202 = bbar[1];
  assign n201bar = b[0];
  assign n201 = bbar[0];
  assign n200bar = n171;
  assign n200 = n171bar;
  assign n199bar = c[7];
  assign n199 = cbar[7];
  assign n198bar = n163;
  assign n198 = n163bar;
  assign n197bar = c[6];
  assign n197 = cbar[6];
  assign n196bar = n155;
  assign n196 = n155bar;
  assign n195bar = c[5];
  assign n195 = cbar[5];
  assign n194bar = n147;
  assign n194 = n147bar;
  assign n193bar = c[4];
  assign n193 = cbar[4];
  assign n192bar = n139;
  assign n192 = n139bar;
  assign n191bar = c[3];
  assign n191 = cbar[3];
  assign n190bar = n131;
  assign n190 = n131bar;
  assign n189bar = c[2];
  assign n189 = cbar[2];
  assign n188bar = n123;
  assign n188 = n123bar;
  assign n187bar = c[1];
  assign n187 = cbar[1];
  assign n186bar = n115;
  assign n186 = n115bar;
  assign n185bar = c[0];
  assign n185 = cbar[0];
  assign n184bar = d[7];
  assign n184 = dbar[7];
  assign n183bar = d[6];
  assign n183 = dbar[6];
  assign n182bar = d[5];
  assign n182 = dbar[5];
  assign n181bar = d[4];
  assign n181 = dbar[4];
  assign n180bar = d[3];
  assign n180 = dbar[3];
  assign n179bar = d[2];
  assign n179 = dbar[2];
  assign n178bar = d[1];
  assign n178 = dbar[1];
  assign n177bar = d[0];
  assign n177 = dbar[0];
  OR2_X1 U49 ( .A1(n176), .A2(n224), .ZN(y[7]) );
  AND2_X1 U49bar ( .A1(n176bar), .A2(n224bar), .ZN(ybar[7]) );
  OR2_X1 U50 ( .A1(n174), .A2(n200), .ZN(n175) );
  AND2_X1 U50bar ( .A1(n174bar), .A2(n200bar), .ZN(n175bar) );
  AND2_X1 U51 ( .A1(n200), .A2(n174), .ZN(n176) );
  OR2_X1 U51bar ( .A1(n200bar), .A2(n174bar), .ZN(n176bar) );
  AND2_X1 U52 ( .A1(n173), .A2(n172), .ZN(n174) );
  OR2_X1 U52bar ( .A1(n173bar), .A2(n172bar), .ZN(n174bar) );
  OR2_X1 U53 ( .A1(n223), .A2(b[7]), .ZN(n172) );
  AND2_X1 U53bar ( .A1(n223bar), .A2(bbar[7]), .ZN(n172bar) );
  OR2_X1 U54 ( .A1(n208), .A2(a[7]), .ZN(n173) );
  AND2_X1 U54bar ( .A1(n208bar), .A2(abar[7]), .ZN(n173bar) );
  AND2_X1 U55 ( .A1(n170), .A2(n169), .ZN(n171) );
  OR2_X1 U55bar ( .A1(n170bar), .A2(n169bar), .ZN(n171bar) );
  OR2_X1 U56 ( .A1(n199), .A2(d[7]), .ZN(n169) );
  AND2_X1 U56bar ( .A1(n199bar), .A2(dbar[7]), .ZN(n169bar) );
  OR2_X1 U57 ( .A1(n184), .A2(c[7]), .ZN(n170) );
  AND2_X1 U57bar ( .A1(n184bar), .A2(cbar[7]), .ZN(n170bar) );
  OR2_X1 U58 ( .A1(n168), .A2(n222), .ZN(y[6]) );
  AND2_X1 U58bar ( .A1(n168bar), .A2(n222bar), .ZN(ybar[6]) );
  OR2_X1 U59 ( .A1(n166), .A2(n198), .ZN(n167) );
  AND2_X1 U59bar ( .A1(n166bar), .A2(n198bar), .ZN(n167bar) );
  AND2_X1 U60 ( .A1(n198), .A2(n166), .ZN(n168) );
  OR2_X1 U60bar ( .A1(n198bar), .A2(n166bar), .ZN(n168bar) );
  AND2_X1 U61 ( .A1(n165), .A2(n164), .ZN(n166) );
  OR2_X1 U61bar ( .A1(n165bar), .A2(n164bar), .ZN(n166bar) );
  OR2_X1 U62 ( .A1(n221), .A2(b[6]), .ZN(n164) );
  AND2_X1 U62bar ( .A1(n221bar), .A2(bbar[6]), .ZN(n164bar) );
  OR2_X1 U63 ( .A1(n207), .A2(a[6]), .ZN(n165) );
  AND2_X1 U63bar ( .A1(n207bar), .A2(abar[6]), .ZN(n165bar) );
  AND2_X1 U64 ( .A1(n162), .A2(n161), .ZN(n163) );
  OR2_X1 U64bar ( .A1(n162bar), .A2(n161bar), .ZN(n163bar) );
  OR2_X1 U65 ( .A1(n197), .A2(d[6]), .ZN(n161) );
  AND2_X1 U65bar ( .A1(n197bar), .A2(dbar[6]), .ZN(n161bar) );
  OR2_X1 U66 ( .A1(n183), .A2(c[6]), .ZN(n162) );
  AND2_X1 U66bar ( .A1(n183bar), .A2(cbar[6]), .ZN(n162bar) );
  OR2_X1 U67 ( .A1(n160), .A2(n220), .ZN(y[5]) );
  AND2_X1 U67bar ( .A1(n160bar), .A2(n220bar), .ZN(ybar[5]) );
  OR2_X1 U68 ( .A1(n158), .A2(n196), .ZN(n159) );
  AND2_X1 U68bar ( .A1(n158bar), .A2(n196bar), .ZN(n159bar) );
  AND2_X1 U69 ( .A1(n196), .A2(n158), .ZN(n160) );
  OR2_X1 U69bar ( .A1(n196bar), .A2(n158bar), .ZN(n160bar) );
  AND2_X1 U70 ( .A1(n157), .A2(n156), .ZN(n158) );
  OR2_X1 U70bar ( .A1(n157bar), .A2(n156bar), .ZN(n158bar) );
  OR2_X1 U71 ( .A1(n219), .A2(b[5]), .ZN(n156) );
  AND2_X1 U71bar ( .A1(n219bar), .A2(bbar[5]), .ZN(n156bar) );
  OR2_X1 U72 ( .A1(n206), .A2(a[5]), .ZN(n157) );
  AND2_X1 U72bar ( .A1(n206bar), .A2(abar[5]), .ZN(n157bar) );
  AND2_X1 U73 ( .A1(n154), .A2(n153), .ZN(n155) );
  OR2_X1 U73bar ( .A1(n154bar), .A2(n153bar), .ZN(n155bar) );
  OR2_X1 U74 ( .A1(n195), .A2(d[5]), .ZN(n153) );
  AND2_X1 U74bar ( .A1(n195bar), .A2(dbar[5]), .ZN(n153bar) );
  OR2_X1 U75 ( .A1(n182), .A2(c[5]), .ZN(n154) );
  AND2_X1 U75bar ( .A1(n182bar), .A2(cbar[5]), .ZN(n154bar) );
  OR2_X1 U76 ( .A1(n152), .A2(n218), .ZN(y[4]) );
  AND2_X1 U76bar ( .A1(n152bar), .A2(n218bar), .ZN(ybar[4]) );
  OR2_X1 U77 ( .A1(n150), .A2(n194), .ZN(n151) );
  AND2_X1 U77bar ( .A1(n150bar), .A2(n194bar), .ZN(n151bar) );
  AND2_X1 U78 ( .A1(n194), .A2(n150), .ZN(n152) );
  OR2_X1 U78bar ( .A1(n194bar), .A2(n150bar), .ZN(n152bar) );
  AND2_X1 U79 ( .A1(n149), .A2(n148), .ZN(n150) );
  OR2_X1 U79bar ( .A1(n149bar), .A2(n148bar), .ZN(n150bar) );
  OR2_X1 U80 ( .A1(n217), .A2(b[4]), .ZN(n148) );
  AND2_X1 U80bar ( .A1(n217bar), .A2(bbar[4]), .ZN(n148bar) );
  OR2_X1 U81 ( .A1(n205), .A2(a[4]), .ZN(n149) );
  AND2_X1 U81bar ( .A1(n205bar), .A2(abar[4]), .ZN(n149bar) );
  AND2_X1 U82 ( .A1(n146), .A2(n145), .ZN(n147) );
  OR2_X1 U82bar ( .A1(n146bar), .A2(n145bar), .ZN(n147bar) );
  OR2_X1 U83 ( .A1(n193), .A2(d[4]), .ZN(n145) );
  AND2_X1 U83bar ( .A1(n193bar), .A2(dbar[4]), .ZN(n145bar) );
  OR2_X1 U84 ( .A1(n181), .A2(c[4]), .ZN(n146) );
  AND2_X1 U84bar ( .A1(n181bar), .A2(cbar[4]), .ZN(n146bar) );
  OR2_X1 U85 ( .A1(n144), .A2(n216), .ZN(y[3]) );
  AND2_X1 U85bar ( .A1(n144bar), .A2(n216bar), .ZN(ybar[3]) );
  OR2_X1 U86 ( .A1(n142), .A2(n192), .ZN(n143) );
  AND2_X1 U86bar ( .A1(n142bar), .A2(n192bar), .ZN(n143bar) );
  AND2_X1 U87 ( .A1(n192), .A2(n142), .ZN(n144) );
  OR2_X1 U87bar ( .A1(n192bar), .A2(n142bar), .ZN(n144bar) );
  AND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(n142) );
  OR2_X1 U88bar ( .A1(n141bar), .A2(n140bar), .ZN(n142bar) );
  OR2_X1 U89 ( .A1(n215), .A2(b[3]), .ZN(n140) );
  AND2_X1 U89bar ( .A1(n215bar), .A2(bbar[3]), .ZN(n140bar) );
  OR2_X1 U90 ( .A1(n204), .A2(a[3]), .ZN(n141) );
  AND2_X1 U90bar ( .A1(n204bar), .A2(abar[3]), .ZN(n141bar) );
  AND2_X1 U91 ( .A1(n138), .A2(n137), .ZN(n139) );
  OR2_X1 U91bar ( .A1(n138bar), .A2(n137bar), .ZN(n139bar) );
  OR2_X1 U92 ( .A1(n191), .A2(d[3]), .ZN(n137) );
  AND2_X1 U92bar ( .A1(n191bar), .A2(dbar[3]), .ZN(n137bar) );
  OR2_X1 U93 ( .A1(n180), .A2(c[3]), .ZN(n138) );
  AND2_X1 U93bar ( .A1(n180bar), .A2(cbar[3]), .ZN(n138bar) );
  OR2_X1 U94 ( .A1(n136), .A2(n214), .ZN(y[2]) );
  AND2_X1 U94bar ( .A1(n136bar), .A2(n214bar), .ZN(ybar[2]) );
  OR2_X1 U95 ( .A1(n134), .A2(n190), .ZN(n135) );
  AND2_X1 U95bar ( .A1(n134bar), .A2(n190bar), .ZN(n135bar) );
  AND2_X1 U96 ( .A1(n190), .A2(n134), .ZN(n136) );
  OR2_X1 U96bar ( .A1(n190bar), .A2(n134bar), .ZN(n136bar) );
  AND2_X1 U97 ( .A1(n133), .A2(n132), .ZN(n134) );
  OR2_X1 U97bar ( .A1(n133bar), .A2(n132bar), .ZN(n134bar) );
  OR2_X1 U98 ( .A1(n213), .A2(b[2]), .ZN(n132) );
  AND2_X1 U98bar ( .A1(n213bar), .A2(bbar[2]), .ZN(n132bar) );
  OR2_X1 U99 ( .A1(n203), .A2(a[2]), .ZN(n133) );
  AND2_X1 U99bar ( .A1(n203bar), .A2(abar[2]), .ZN(n133bar) );
  AND2_X1 U100 ( .A1(n130), .A2(n129), .ZN(n131) );
  OR2_X1 U100bar ( .A1(n130bar), .A2(n129bar), .ZN(n131bar) );
  OR2_X1 U101 ( .A1(n189), .A2(d[2]), .ZN(n129) );
  AND2_X1 U101bar ( .A1(n189bar), .A2(dbar[2]), .ZN(n129bar) );
  OR2_X1 U102 ( .A1(n179), .A2(c[2]), .ZN(n130) );
  AND2_X1 U102bar ( .A1(n179bar), .A2(cbar[2]), .ZN(n130bar) );
  OR2_X1 U103 ( .A1(n128), .A2(n212), .ZN(y[1]) );
  AND2_X1 U103bar ( .A1(n128bar), .A2(n212bar), .ZN(ybar[1]) );
  OR2_X1 U104 ( .A1(n126), .A2(n188), .ZN(n127) );
  AND2_X1 U104bar ( .A1(n126bar), .A2(n188bar), .ZN(n127bar) );
  AND2_X1 U105 ( .A1(n188), .A2(n126), .ZN(n128) );
  OR2_X1 U105bar ( .A1(n188bar), .A2(n126bar), .ZN(n128bar) );
  AND2_X1 U106 ( .A1(n125), .A2(n124), .ZN(n126) );
  OR2_X1 U106bar ( .A1(n125bar), .A2(n124bar), .ZN(n126bar) );
  OR2_X1 U107 ( .A1(n211), .A2(b[1]), .ZN(n124) );
  AND2_X1 U107bar ( .A1(n211bar), .A2(bbar[1]), .ZN(n124bar) );
  OR2_X1 U108 ( .A1(n202), .A2(a[1]), .ZN(n125) );
  AND2_X1 U108bar ( .A1(n202bar), .A2(abar[1]), .ZN(n125bar) );
  AND2_X1 U109 ( .A1(n122), .A2(n121), .ZN(n123) );
  OR2_X1 U109bar ( .A1(n122bar), .A2(n121bar), .ZN(n123bar) );
  OR2_X1 U110 ( .A1(n187), .A2(d[1]), .ZN(n121) );
  AND2_X1 U110bar ( .A1(n187bar), .A2(dbar[1]), .ZN(n121bar) );
  OR2_X1 U111 ( .A1(n178), .A2(c[1]), .ZN(n122) );
  AND2_X1 U111bar ( .A1(n178bar), .A2(cbar[1]), .ZN(n122bar) );
  OR2_X1 U112 ( .A1(n120), .A2(n210), .ZN(y[0]) );
  AND2_X1 U112bar ( .A1(n120bar), .A2(n210bar), .ZN(ybar[0]) );
  OR2_X1 U113 ( .A1(n118), .A2(n186), .ZN(n119) );
  AND2_X1 U113bar ( .A1(n118bar), .A2(n186bar), .ZN(n119bar) );
  AND2_X1 U114 ( .A1(n186), .A2(n118), .ZN(n120) );
  OR2_X1 U114bar ( .A1(n186bar), .A2(n118bar), .ZN(n120bar) );
  AND2_X1 U115 ( .A1(n117), .A2(n116), .ZN(n118) );
  OR2_X1 U115bar ( .A1(n117bar), .A2(n116bar), .ZN(n118bar) );
  OR2_X1 U116 ( .A1(n209), .A2(b[0]), .ZN(n116) );
  AND2_X1 U116bar ( .A1(n209bar), .A2(bbar[0]), .ZN(n116bar) );
  OR2_X1 U117 ( .A1(n201), .A2(a[0]), .ZN(n117) );
  AND2_X1 U117bar ( .A1(n201bar), .A2(abar[0]), .ZN(n117bar) );
  AND2_X1 U118 ( .A1(n114), .A2(n113), .ZN(n115) );
  OR2_X1 U118bar ( .A1(n114bar), .A2(n113bar), .ZN(n115bar) );
  OR2_X1 U119 ( .A1(n185), .A2(d[0]), .ZN(n113) );
  AND2_X1 U119bar ( .A1(n185bar), .A2(dbar[0]), .ZN(n113bar) );
  OR2_X1 U120 ( .A1(n177), .A2(c[0]), .ZN(n114) );
  AND2_X1 U120bar ( .A1(n177bar), .A2(cbar[0]), .ZN(n114bar) );
endmodule

module byteXor4_6 ( a, b, c, d, y );

  input wire [7:0] a;
  input wire [7:0] b;
  input wire [7:0] c;
  input wire [7:0] d;
  wire [7:0] abar;
  wire [7:0] bbar;
  wire [7:0] cbar;
  wire [7:0] dbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign cbar[0] = ~c[0];
  assign cbar[1] = ~c[1];
  assign cbar[2] = ~c[2];
  assign cbar[3] = ~c[3];
  assign cbar[4] = ~c[4];
  assign cbar[5] = ~c[5];
  assign cbar[6] = ~c[6];
  assign cbar[7] = ~c[7];
  assign dbar[0] = ~d[0];
  assign dbar[1] = ~d[1];
  assign dbar[2] = ~d[2];
  assign dbar[3] = ~d[3];
  assign dbar[4] = ~d[4];
  assign dbar[5] = ~d[5];
  assign dbar[6] = ~d[6];
  assign dbar[7] = ~d[7];
//input_done

  output wire [7:0] y;
  wire [7:0] ybar;
//output_done

  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n113bar;
  wire n114bar;
  wire n115bar;
  wire n116bar;
  wire n117bar;
  wire n118bar;
  wire n119bar;
  wire n120bar;
  wire n121bar;
  wire n122bar;
  wire n123bar;
  wire n124bar;
  wire n125bar;
  wire n126bar;
  wire n127bar;
  wire n128bar;
  wire n129bar;
  wire n130bar;
  wire n131bar;
  wire n132bar;
  wire n133bar;
  wire n134bar;
  wire n135bar;
  wire n136bar;
  wire n137bar;
  wire n138bar;
  wire n139bar;
  wire n140bar;
  wire n141bar;
  wire n142bar;
  wire n143bar;
  wire n144bar;
  wire n145bar;
  wire n146bar;
  wire n147bar;
  wire n148bar;
  wire n149bar;
  wire n150bar;
  wire n151bar;
  wire n152bar;
  wire n153bar;
  wire n154bar;
  wire n155bar;
  wire n156bar;
  wire n157bar;
  wire n158bar;
  wire n159bar;
  wire n160bar;
  wire n161bar;
  wire n162bar;
  wire n163bar;
  wire n164bar;
  wire n165bar;
  wire n166bar;
  wire n167bar;
  wire n168bar;
  wire n169bar;
  wire n170bar;
  wire n171bar;
  wire n172bar;
  wire n173bar;
  wire n174bar;
  wire n175bar;
  wire n176bar;
  wire n177bar;
  wire n178bar;
  wire n179bar;
  wire n180bar;
  wire n181bar;
  wire n182bar;
  wire n183bar;
  wire n184bar;
  wire n185bar;
  wire n186bar;
  wire n187bar;
  wire n188bar;
  wire n189bar;
  wire n190bar;
  wire n191bar;
  wire n192bar;
  wire n193bar;
  wire n194bar;
  wire n195bar;
  wire n196bar;
  wire n197bar;
  wire n198bar;
  wire n199bar;
  wire n200bar;
  wire n201bar;
  wire n202bar;
  wire n203bar;
  wire n204bar;
  wire n205bar;
  wire n206bar;
  wire n207bar;
  wire n208bar;
  wire n209bar;
  wire n210bar;
  wire n211bar;
  wire n212bar;
  wire n213bar;
  wire n214bar;
  wire n215bar;
  wire n216bar;
  wire n217bar;
  wire n218bar;
  wire n219bar;
  wire n220bar;
  wire n221bar;
  wire n222bar;
  wire n223bar;
  wire n224bar;
//wire_done

 //assign_done

  assign n224bar = n175;
  assign n224 = n175bar;
  assign n223bar = a[7];
  assign n223 = abar[7];
  assign n222bar = n167;
  assign n222 = n167bar;
  assign n221bar = a[6];
  assign n221 = abar[6];
  assign n220bar = n159;
  assign n220 = n159bar;
  assign n219bar = a[5];
  assign n219 = abar[5];
  assign n218bar = n151;
  assign n218 = n151bar;
  assign n217bar = a[4];
  assign n217 = abar[4];
  assign n216bar = n143;
  assign n216 = n143bar;
  assign n215bar = a[3];
  assign n215 = abar[3];
  assign n214bar = n135;
  assign n214 = n135bar;
  assign n213bar = a[2];
  assign n213 = abar[2];
  assign n212bar = n127;
  assign n212 = n127bar;
  assign n211bar = a[1];
  assign n211 = abar[1];
  assign n210bar = n119;
  assign n210 = n119bar;
  assign n209bar = a[0];
  assign n209 = abar[0];
  assign n208bar = b[7];
  assign n208 = bbar[7];
  assign n207bar = b[6];
  assign n207 = bbar[6];
  assign n206bar = b[5];
  assign n206 = bbar[5];
  assign n205bar = b[4];
  assign n205 = bbar[4];
  assign n204bar = b[3];
  assign n204 = bbar[3];
  assign n203bar = b[2];
  assign n203 = bbar[2];
  assign n202bar = b[1];
  assign n202 = bbar[1];
  assign n201bar = b[0];
  assign n201 = bbar[0];
  assign n200bar = n171;
  assign n200 = n171bar;
  assign n199bar = c[7];
  assign n199 = cbar[7];
  assign n198bar = n163;
  assign n198 = n163bar;
  assign n197bar = c[6];
  assign n197 = cbar[6];
  assign n196bar = n155;
  assign n196 = n155bar;
  assign n195bar = c[5];
  assign n195 = cbar[5];
  assign n194bar = n147;
  assign n194 = n147bar;
  assign n193bar = c[4];
  assign n193 = cbar[4];
  assign n192bar = n139;
  assign n192 = n139bar;
  assign n191bar = c[3];
  assign n191 = cbar[3];
  assign n190bar = n131;
  assign n190 = n131bar;
  assign n189bar = c[2];
  assign n189 = cbar[2];
  assign n188bar = n123;
  assign n188 = n123bar;
  assign n187bar = c[1];
  assign n187 = cbar[1];
  assign n186bar = n115;
  assign n186 = n115bar;
  assign n185bar = c[0];
  assign n185 = cbar[0];
  assign n184bar = d[7];
  assign n184 = dbar[7];
  assign n183bar = d[6];
  assign n183 = dbar[6];
  assign n182bar = d[5];
  assign n182 = dbar[5];
  assign n181bar = d[4];
  assign n181 = dbar[4];
  assign n180bar = d[3];
  assign n180 = dbar[3];
  assign n179bar = d[2];
  assign n179 = dbar[2];
  assign n178bar = d[1];
  assign n178 = dbar[1];
  assign n177bar = d[0];
  assign n177 = dbar[0];
  OR2_X1 U49 ( .A1(n176), .A2(n224), .ZN(y[7]) );
  AND2_X1 U49bar ( .A1(n176bar), .A2(n224bar), .ZN(ybar[7]) );
  OR2_X1 U50 ( .A1(n174), .A2(n200), .ZN(n175) );
  AND2_X1 U50bar ( .A1(n174bar), .A2(n200bar), .ZN(n175bar) );
  AND2_X1 U51 ( .A1(n200), .A2(n174), .ZN(n176) );
  OR2_X1 U51bar ( .A1(n200bar), .A2(n174bar), .ZN(n176bar) );
  AND2_X1 U52 ( .A1(n173), .A2(n172), .ZN(n174) );
  OR2_X1 U52bar ( .A1(n173bar), .A2(n172bar), .ZN(n174bar) );
  OR2_X1 U53 ( .A1(n223), .A2(b[7]), .ZN(n172) );
  AND2_X1 U53bar ( .A1(n223bar), .A2(bbar[7]), .ZN(n172bar) );
  OR2_X1 U54 ( .A1(n208), .A2(a[7]), .ZN(n173) );
  AND2_X1 U54bar ( .A1(n208bar), .A2(abar[7]), .ZN(n173bar) );
  AND2_X1 U55 ( .A1(n170), .A2(n169), .ZN(n171) );
  OR2_X1 U55bar ( .A1(n170bar), .A2(n169bar), .ZN(n171bar) );
  OR2_X1 U56 ( .A1(n199), .A2(d[7]), .ZN(n169) );
  AND2_X1 U56bar ( .A1(n199bar), .A2(dbar[7]), .ZN(n169bar) );
  OR2_X1 U57 ( .A1(n184), .A2(c[7]), .ZN(n170) );
  AND2_X1 U57bar ( .A1(n184bar), .A2(cbar[7]), .ZN(n170bar) );
  OR2_X1 U58 ( .A1(n168), .A2(n222), .ZN(y[6]) );
  AND2_X1 U58bar ( .A1(n168bar), .A2(n222bar), .ZN(ybar[6]) );
  OR2_X1 U59 ( .A1(n166), .A2(n198), .ZN(n167) );
  AND2_X1 U59bar ( .A1(n166bar), .A2(n198bar), .ZN(n167bar) );
  AND2_X1 U60 ( .A1(n198), .A2(n166), .ZN(n168) );
  OR2_X1 U60bar ( .A1(n198bar), .A2(n166bar), .ZN(n168bar) );
  AND2_X1 U61 ( .A1(n165), .A2(n164), .ZN(n166) );
  OR2_X1 U61bar ( .A1(n165bar), .A2(n164bar), .ZN(n166bar) );
  OR2_X1 U62 ( .A1(n221), .A2(b[6]), .ZN(n164) );
  AND2_X1 U62bar ( .A1(n221bar), .A2(bbar[6]), .ZN(n164bar) );
  OR2_X1 U63 ( .A1(n207), .A2(a[6]), .ZN(n165) );
  AND2_X1 U63bar ( .A1(n207bar), .A2(abar[6]), .ZN(n165bar) );
  AND2_X1 U64 ( .A1(n162), .A2(n161), .ZN(n163) );
  OR2_X1 U64bar ( .A1(n162bar), .A2(n161bar), .ZN(n163bar) );
  OR2_X1 U65 ( .A1(n197), .A2(d[6]), .ZN(n161) );
  AND2_X1 U65bar ( .A1(n197bar), .A2(dbar[6]), .ZN(n161bar) );
  OR2_X1 U66 ( .A1(n183), .A2(c[6]), .ZN(n162) );
  AND2_X1 U66bar ( .A1(n183bar), .A2(cbar[6]), .ZN(n162bar) );
  OR2_X1 U67 ( .A1(n160), .A2(n220), .ZN(y[5]) );
  AND2_X1 U67bar ( .A1(n160bar), .A2(n220bar), .ZN(ybar[5]) );
  OR2_X1 U68 ( .A1(n158), .A2(n196), .ZN(n159) );
  AND2_X1 U68bar ( .A1(n158bar), .A2(n196bar), .ZN(n159bar) );
  AND2_X1 U69 ( .A1(n196), .A2(n158), .ZN(n160) );
  OR2_X1 U69bar ( .A1(n196bar), .A2(n158bar), .ZN(n160bar) );
  AND2_X1 U70 ( .A1(n157), .A2(n156), .ZN(n158) );
  OR2_X1 U70bar ( .A1(n157bar), .A2(n156bar), .ZN(n158bar) );
  OR2_X1 U71 ( .A1(n219), .A2(b[5]), .ZN(n156) );
  AND2_X1 U71bar ( .A1(n219bar), .A2(bbar[5]), .ZN(n156bar) );
  OR2_X1 U72 ( .A1(n206), .A2(a[5]), .ZN(n157) );
  AND2_X1 U72bar ( .A1(n206bar), .A2(abar[5]), .ZN(n157bar) );
  AND2_X1 U73 ( .A1(n154), .A2(n153), .ZN(n155) );
  OR2_X1 U73bar ( .A1(n154bar), .A2(n153bar), .ZN(n155bar) );
  OR2_X1 U74 ( .A1(n195), .A2(d[5]), .ZN(n153) );
  AND2_X1 U74bar ( .A1(n195bar), .A2(dbar[5]), .ZN(n153bar) );
  OR2_X1 U75 ( .A1(n182), .A2(c[5]), .ZN(n154) );
  AND2_X1 U75bar ( .A1(n182bar), .A2(cbar[5]), .ZN(n154bar) );
  OR2_X1 U76 ( .A1(n152), .A2(n218), .ZN(y[4]) );
  AND2_X1 U76bar ( .A1(n152bar), .A2(n218bar), .ZN(ybar[4]) );
  OR2_X1 U77 ( .A1(n150), .A2(n194), .ZN(n151) );
  AND2_X1 U77bar ( .A1(n150bar), .A2(n194bar), .ZN(n151bar) );
  AND2_X1 U78 ( .A1(n194), .A2(n150), .ZN(n152) );
  OR2_X1 U78bar ( .A1(n194bar), .A2(n150bar), .ZN(n152bar) );
  AND2_X1 U79 ( .A1(n149), .A2(n148), .ZN(n150) );
  OR2_X1 U79bar ( .A1(n149bar), .A2(n148bar), .ZN(n150bar) );
  OR2_X1 U80 ( .A1(n217), .A2(b[4]), .ZN(n148) );
  AND2_X1 U80bar ( .A1(n217bar), .A2(bbar[4]), .ZN(n148bar) );
  OR2_X1 U81 ( .A1(n205), .A2(a[4]), .ZN(n149) );
  AND2_X1 U81bar ( .A1(n205bar), .A2(abar[4]), .ZN(n149bar) );
  AND2_X1 U82 ( .A1(n146), .A2(n145), .ZN(n147) );
  OR2_X1 U82bar ( .A1(n146bar), .A2(n145bar), .ZN(n147bar) );
  OR2_X1 U83 ( .A1(n193), .A2(d[4]), .ZN(n145) );
  AND2_X1 U83bar ( .A1(n193bar), .A2(dbar[4]), .ZN(n145bar) );
  OR2_X1 U84 ( .A1(n181), .A2(c[4]), .ZN(n146) );
  AND2_X1 U84bar ( .A1(n181bar), .A2(cbar[4]), .ZN(n146bar) );
  OR2_X1 U85 ( .A1(n144), .A2(n216), .ZN(y[3]) );
  AND2_X1 U85bar ( .A1(n144bar), .A2(n216bar), .ZN(ybar[3]) );
  OR2_X1 U86 ( .A1(n142), .A2(n192), .ZN(n143) );
  AND2_X1 U86bar ( .A1(n142bar), .A2(n192bar), .ZN(n143bar) );
  AND2_X1 U87 ( .A1(n192), .A2(n142), .ZN(n144) );
  OR2_X1 U87bar ( .A1(n192bar), .A2(n142bar), .ZN(n144bar) );
  AND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(n142) );
  OR2_X1 U88bar ( .A1(n141bar), .A2(n140bar), .ZN(n142bar) );
  OR2_X1 U89 ( .A1(n215), .A2(b[3]), .ZN(n140) );
  AND2_X1 U89bar ( .A1(n215bar), .A2(bbar[3]), .ZN(n140bar) );
  OR2_X1 U90 ( .A1(n204), .A2(a[3]), .ZN(n141) );
  AND2_X1 U90bar ( .A1(n204bar), .A2(abar[3]), .ZN(n141bar) );
  AND2_X1 U91 ( .A1(n138), .A2(n137), .ZN(n139) );
  OR2_X1 U91bar ( .A1(n138bar), .A2(n137bar), .ZN(n139bar) );
  OR2_X1 U92 ( .A1(n191), .A2(d[3]), .ZN(n137) );
  AND2_X1 U92bar ( .A1(n191bar), .A2(dbar[3]), .ZN(n137bar) );
  OR2_X1 U93 ( .A1(n180), .A2(c[3]), .ZN(n138) );
  AND2_X1 U93bar ( .A1(n180bar), .A2(cbar[3]), .ZN(n138bar) );
  OR2_X1 U94 ( .A1(n136), .A2(n214), .ZN(y[2]) );
  AND2_X1 U94bar ( .A1(n136bar), .A2(n214bar), .ZN(ybar[2]) );
  OR2_X1 U95 ( .A1(n134), .A2(n190), .ZN(n135) );
  AND2_X1 U95bar ( .A1(n134bar), .A2(n190bar), .ZN(n135bar) );
  AND2_X1 U96 ( .A1(n190), .A2(n134), .ZN(n136) );
  OR2_X1 U96bar ( .A1(n190bar), .A2(n134bar), .ZN(n136bar) );
  AND2_X1 U97 ( .A1(n133), .A2(n132), .ZN(n134) );
  OR2_X1 U97bar ( .A1(n133bar), .A2(n132bar), .ZN(n134bar) );
  OR2_X1 U98 ( .A1(n213), .A2(b[2]), .ZN(n132) );
  AND2_X1 U98bar ( .A1(n213bar), .A2(bbar[2]), .ZN(n132bar) );
  OR2_X1 U99 ( .A1(n203), .A2(a[2]), .ZN(n133) );
  AND2_X1 U99bar ( .A1(n203bar), .A2(abar[2]), .ZN(n133bar) );
  AND2_X1 U100 ( .A1(n130), .A2(n129), .ZN(n131) );
  OR2_X1 U100bar ( .A1(n130bar), .A2(n129bar), .ZN(n131bar) );
  OR2_X1 U101 ( .A1(n189), .A2(d[2]), .ZN(n129) );
  AND2_X1 U101bar ( .A1(n189bar), .A2(dbar[2]), .ZN(n129bar) );
  OR2_X1 U102 ( .A1(n179), .A2(c[2]), .ZN(n130) );
  AND2_X1 U102bar ( .A1(n179bar), .A2(cbar[2]), .ZN(n130bar) );
  OR2_X1 U103 ( .A1(n128), .A2(n212), .ZN(y[1]) );
  AND2_X1 U103bar ( .A1(n128bar), .A2(n212bar), .ZN(ybar[1]) );
  OR2_X1 U104 ( .A1(n126), .A2(n188), .ZN(n127) );
  AND2_X1 U104bar ( .A1(n126bar), .A2(n188bar), .ZN(n127bar) );
  AND2_X1 U105 ( .A1(n188), .A2(n126), .ZN(n128) );
  OR2_X1 U105bar ( .A1(n188bar), .A2(n126bar), .ZN(n128bar) );
  AND2_X1 U106 ( .A1(n125), .A2(n124), .ZN(n126) );
  OR2_X1 U106bar ( .A1(n125bar), .A2(n124bar), .ZN(n126bar) );
  OR2_X1 U107 ( .A1(n211), .A2(b[1]), .ZN(n124) );
  AND2_X1 U107bar ( .A1(n211bar), .A2(bbar[1]), .ZN(n124bar) );
  OR2_X1 U108 ( .A1(n202), .A2(a[1]), .ZN(n125) );
  AND2_X1 U108bar ( .A1(n202bar), .A2(abar[1]), .ZN(n125bar) );
  AND2_X1 U109 ( .A1(n122), .A2(n121), .ZN(n123) );
  OR2_X1 U109bar ( .A1(n122bar), .A2(n121bar), .ZN(n123bar) );
  OR2_X1 U110 ( .A1(n187), .A2(d[1]), .ZN(n121) );
  AND2_X1 U110bar ( .A1(n187bar), .A2(dbar[1]), .ZN(n121bar) );
  OR2_X1 U111 ( .A1(n178), .A2(c[1]), .ZN(n122) );
  AND2_X1 U111bar ( .A1(n178bar), .A2(cbar[1]), .ZN(n122bar) );
  OR2_X1 U112 ( .A1(n120), .A2(n210), .ZN(y[0]) );
  AND2_X1 U112bar ( .A1(n120bar), .A2(n210bar), .ZN(ybar[0]) );
  OR2_X1 U113 ( .A1(n118), .A2(n186), .ZN(n119) );
  AND2_X1 U113bar ( .A1(n118bar), .A2(n186bar), .ZN(n119bar) );
  AND2_X1 U114 ( .A1(n186), .A2(n118), .ZN(n120) );
  OR2_X1 U114bar ( .A1(n186bar), .A2(n118bar), .ZN(n120bar) );
  AND2_X1 U115 ( .A1(n117), .A2(n116), .ZN(n118) );
  OR2_X1 U115bar ( .A1(n117bar), .A2(n116bar), .ZN(n118bar) );
  OR2_X1 U116 ( .A1(n209), .A2(b[0]), .ZN(n116) );
  AND2_X1 U116bar ( .A1(n209bar), .A2(bbar[0]), .ZN(n116bar) );
  OR2_X1 U117 ( .A1(n201), .A2(a[0]), .ZN(n117) );
  AND2_X1 U117bar ( .A1(n201bar), .A2(abar[0]), .ZN(n117bar) );
  AND2_X1 U118 ( .A1(n114), .A2(n113), .ZN(n115) );
  OR2_X1 U118bar ( .A1(n114bar), .A2(n113bar), .ZN(n115bar) );
  OR2_X1 U119 ( .A1(n185), .A2(d[0]), .ZN(n113) );
  AND2_X1 U119bar ( .A1(n185bar), .A2(dbar[0]), .ZN(n113bar) );
  OR2_X1 U120 ( .A1(n177), .A2(c[0]), .ZN(n114) );
  AND2_X1 U120bar ( .A1(n177bar), .A2(cbar[0]), .ZN(n114bar) );
endmodule

module byteXor4_7 ( a, b, c, d, y );

  input wire [7:0] a;
  input wire [7:0] b;
  input wire [7:0] c;
  input wire [7:0] d;
  wire [7:0] abar;
  wire [7:0] bbar;
  wire [7:0] cbar;
  wire [7:0] dbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign cbar[0] = ~c[0];
  assign cbar[1] = ~c[1];
  assign cbar[2] = ~c[2];
  assign cbar[3] = ~c[3];
  assign cbar[4] = ~c[4];
  assign cbar[5] = ~c[5];
  assign cbar[6] = ~c[6];
  assign cbar[7] = ~c[7];
  assign dbar[0] = ~d[0];
  assign dbar[1] = ~d[1];
  assign dbar[2] = ~d[2];
  assign dbar[3] = ~d[3];
  assign dbar[4] = ~d[4];
  assign dbar[5] = ~d[5];
  assign dbar[6] = ~d[6];
  assign dbar[7] = ~d[7];
//input_done

  output wire [7:0] y;
  wire [7:0] ybar;
//output_done

  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n113bar;
  wire n114bar;
  wire n115bar;
  wire n116bar;
  wire n117bar;
  wire n118bar;
  wire n119bar;
  wire n120bar;
  wire n121bar;
  wire n122bar;
  wire n123bar;
  wire n124bar;
  wire n125bar;
  wire n126bar;
  wire n127bar;
  wire n128bar;
  wire n129bar;
  wire n130bar;
  wire n131bar;
  wire n132bar;
  wire n133bar;
  wire n134bar;
  wire n135bar;
  wire n136bar;
  wire n137bar;
  wire n138bar;
  wire n139bar;
  wire n140bar;
  wire n141bar;
  wire n142bar;
  wire n143bar;
  wire n144bar;
  wire n145bar;
  wire n146bar;
  wire n147bar;
  wire n148bar;
  wire n149bar;
  wire n150bar;
  wire n151bar;
  wire n152bar;
  wire n153bar;
  wire n154bar;
  wire n155bar;
  wire n156bar;
  wire n157bar;
  wire n158bar;
  wire n159bar;
  wire n160bar;
  wire n161bar;
  wire n162bar;
  wire n163bar;
  wire n164bar;
  wire n165bar;
  wire n166bar;
  wire n167bar;
  wire n168bar;
  wire n169bar;
  wire n170bar;
  wire n171bar;
  wire n172bar;
  wire n173bar;
  wire n174bar;
  wire n175bar;
  wire n176bar;
  wire n177bar;
  wire n178bar;
  wire n179bar;
  wire n180bar;
  wire n181bar;
  wire n182bar;
  wire n183bar;
  wire n184bar;
  wire n185bar;
  wire n186bar;
  wire n187bar;
  wire n188bar;
  wire n189bar;
  wire n190bar;
  wire n191bar;
  wire n192bar;
  wire n193bar;
  wire n194bar;
  wire n195bar;
  wire n196bar;
  wire n197bar;
  wire n198bar;
  wire n199bar;
  wire n200bar;
  wire n201bar;
  wire n202bar;
  wire n203bar;
  wire n204bar;
  wire n205bar;
  wire n206bar;
  wire n207bar;
  wire n208bar;
  wire n209bar;
  wire n210bar;
  wire n211bar;
  wire n212bar;
  wire n213bar;
  wire n214bar;
  wire n215bar;
  wire n216bar;
  wire n217bar;
  wire n218bar;
  wire n219bar;
  wire n220bar;
  wire n221bar;
  wire n222bar;
  wire n223bar;
  wire n224bar;
//wire_done

 //assign_done

  assign n224bar = n175;
  assign n224 = n175bar;
  assign n223bar = a[7];
  assign n223 = abar[7];
  assign n222bar = n167;
  assign n222 = n167bar;
  assign n221bar = a[6];
  assign n221 = abar[6];
  assign n220bar = n159;
  assign n220 = n159bar;
  assign n219bar = a[5];
  assign n219 = abar[5];
  assign n218bar = n151;
  assign n218 = n151bar;
  assign n217bar = a[4];
  assign n217 = abar[4];
  assign n216bar = n143;
  assign n216 = n143bar;
  assign n215bar = a[3];
  assign n215 = abar[3];
  assign n214bar = n135;
  assign n214 = n135bar;
  assign n213bar = a[2];
  assign n213 = abar[2];
  assign n212bar = n127;
  assign n212 = n127bar;
  assign n211bar = a[1];
  assign n211 = abar[1];
  assign n210bar = n119;
  assign n210 = n119bar;
  assign n209bar = a[0];
  assign n209 = abar[0];
  assign n208bar = b[7];
  assign n208 = bbar[7];
  assign n207bar = b[6];
  assign n207 = bbar[6];
  assign n206bar = b[5];
  assign n206 = bbar[5];
  assign n205bar = b[4];
  assign n205 = bbar[4];
  assign n204bar = b[3];
  assign n204 = bbar[3];
  assign n203bar = b[2];
  assign n203 = bbar[2];
  assign n202bar = b[1];
  assign n202 = bbar[1];
  assign n201bar = b[0];
  assign n201 = bbar[0];
  assign n200bar = n171;
  assign n200 = n171bar;
  assign n199bar = c[7];
  assign n199 = cbar[7];
  assign n198bar = n163;
  assign n198 = n163bar;
  assign n197bar = c[6];
  assign n197 = cbar[6];
  assign n196bar = n155;
  assign n196 = n155bar;
  assign n195bar = c[5];
  assign n195 = cbar[5];
  assign n194bar = n147;
  assign n194 = n147bar;
  assign n193bar = c[4];
  assign n193 = cbar[4];
  assign n192bar = n139;
  assign n192 = n139bar;
  assign n191bar = c[3];
  assign n191 = cbar[3];
  assign n190bar = n131;
  assign n190 = n131bar;
  assign n189bar = c[2];
  assign n189 = cbar[2];
  assign n188bar = n123;
  assign n188 = n123bar;
  assign n187bar = c[1];
  assign n187 = cbar[1];
  assign n186bar = n115;
  assign n186 = n115bar;
  assign n185bar = c[0];
  assign n185 = cbar[0];
  assign n184bar = d[7];
  assign n184 = dbar[7];
  assign n183bar = d[6];
  assign n183 = dbar[6];
  assign n182bar = d[5];
  assign n182 = dbar[5];
  assign n181bar = d[4];
  assign n181 = dbar[4];
  assign n180bar = d[3];
  assign n180 = dbar[3];
  assign n179bar = d[2];
  assign n179 = dbar[2];
  assign n178bar = d[1];
  assign n178 = dbar[1];
  assign n177bar = d[0];
  assign n177 = dbar[0];
  OR2_X1 U49 ( .A1(n176), .A2(n224), .ZN(y[7]) );
  AND2_X1 U49bar ( .A1(n176bar), .A2(n224bar), .ZN(ybar[7]) );
  OR2_X1 U50 ( .A1(n174), .A2(n200), .ZN(n175) );
  AND2_X1 U50bar ( .A1(n174bar), .A2(n200bar), .ZN(n175bar) );
  AND2_X1 U51 ( .A1(n200), .A2(n174), .ZN(n176) );
  OR2_X1 U51bar ( .A1(n200bar), .A2(n174bar), .ZN(n176bar) );
  AND2_X1 U52 ( .A1(n173), .A2(n172), .ZN(n174) );
  OR2_X1 U52bar ( .A1(n173bar), .A2(n172bar), .ZN(n174bar) );
  OR2_X1 U53 ( .A1(n223), .A2(b[7]), .ZN(n172) );
  AND2_X1 U53bar ( .A1(n223bar), .A2(bbar[7]), .ZN(n172bar) );
  OR2_X1 U54 ( .A1(n208), .A2(a[7]), .ZN(n173) );
  AND2_X1 U54bar ( .A1(n208bar), .A2(abar[7]), .ZN(n173bar) );
  AND2_X1 U55 ( .A1(n170), .A2(n169), .ZN(n171) );
  OR2_X1 U55bar ( .A1(n170bar), .A2(n169bar), .ZN(n171bar) );
  OR2_X1 U56 ( .A1(n199), .A2(d[7]), .ZN(n169) );
  AND2_X1 U56bar ( .A1(n199bar), .A2(dbar[7]), .ZN(n169bar) );
  OR2_X1 U57 ( .A1(n184), .A2(c[7]), .ZN(n170) );
  AND2_X1 U57bar ( .A1(n184bar), .A2(cbar[7]), .ZN(n170bar) );
  OR2_X1 U58 ( .A1(n168), .A2(n222), .ZN(y[6]) );
  AND2_X1 U58bar ( .A1(n168bar), .A2(n222bar), .ZN(ybar[6]) );
  OR2_X1 U59 ( .A1(n166), .A2(n198), .ZN(n167) );
  AND2_X1 U59bar ( .A1(n166bar), .A2(n198bar), .ZN(n167bar) );
  AND2_X1 U60 ( .A1(n198), .A2(n166), .ZN(n168) );
  OR2_X1 U60bar ( .A1(n198bar), .A2(n166bar), .ZN(n168bar) );
  AND2_X1 U61 ( .A1(n165), .A2(n164), .ZN(n166) );
  OR2_X1 U61bar ( .A1(n165bar), .A2(n164bar), .ZN(n166bar) );
  OR2_X1 U62 ( .A1(n221), .A2(b[6]), .ZN(n164) );
  AND2_X1 U62bar ( .A1(n221bar), .A2(bbar[6]), .ZN(n164bar) );
  OR2_X1 U63 ( .A1(n207), .A2(a[6]), .ZN(n165) );
  AND2_X1 U63bar ( .A1(n207bar), .A2(abar[6]), .ZN(n165bar) );
  AND2_X1 U64 ( .A1(n162), .A2(n161), .ZN(n163) );
  OR2_X1 U64bar ( .A1(n162bar), .A2(n161bar), .ZN(n163bar) );
  OR2_X1 U65 ( .A1(n197), .A2(d[6]), .ZN(n161) );
  AND2_X1 U65bar ( .A1(n197bar), .A2(dbar[6]), .ZN(n161bar) );
  OR2_X1 U66 ( .A1(n183), .A2(c[6]), .ZN(n162) );
  AND2_X1 U66bar ( .A1(n183bar), .A2(cbar[6]), .ZN(n162bar) );
  OR2_X1 U67 ( .A1(n160), .A2(n220), .ZN(y[5]) );
  AND2_X1 U67bar ( .A1(n160bar), .A2(n220bar), .ZN(ybar[5]) );
  OR2_X1 U68 ( .A1(n158), .A2(n196), .ZN(n159) );
  AND2_X1 U68bar ( .A1(n158bar), .A2(n196bar), .ZN(n159bar) );
  AND2_X1 U69 ( .A1(n196), .A2(n158), .ZN(n160) );
  OR2_X1 U69bar ( .A1(n196bar), .A2(n158bar), .ZN(n160bar) );
  AND2_X1 U70 ( .A1(n157), .A2(n156), .ZN(n158) );
  OR2_X1 U70bar ( .A1(n157bar), .A2(n156bar), .ZN(n158bar) );
  OR2_X1 U71 ( .A1(n219), .A2(b[5]), .ZN(n156) );
  AND2_X1 U71bar ( .A1(n219bar), .A2(bbar[5]), .ZN(n156bar) );
  OR2_X1 U72 ( .A1(n206), .A2(a[5]), .ZN(n157) );
  AND2_X1 U72bar ( .A1(n206bar), .A2(abar[5]), .ZN(n157bar) );
  AND2_X1 U73 ( .A1(n154), .A2(n153), .ZN(n155) );
  OR2_X1 U73bar ( .A1(n154bar), .A2(n153bar), .ZN(n155bar) );
  OR2_X1 U74 ( .A1(n195), .A2(d[5]), .ZN(n153) );
  AND2_X1 U74bar ( .A1(n195bar), .A2(dbar[5]), .ZN(n153bar) );
  OR2_X1 U75 ( .A1(n182), .A2(c[5]), .ZN(n154) );
  AND2_X1 U75bar ( .A1(n182bar), .A2(cbar[5]), .ZN(n154bar) );
  OR2_X1 U76 ( .A1(n152), .A2(n218), .ZN(y[4]) );
  AND2_X1 U76bar ( .A1(n152bar), .A2(n218bar), .ZN(ybar[4]) );
  OR2_X1 U77 ( .A1(n150), .A2(n194), .ZN(n151) );
  AND2_X1 U77bar ( .A1(n150bar), .A2(n194bar), .ZN(n151bar) );
  AND2_X1 U78 ( .A1(n194), .A2(n150), .ZN(n152) );
  OR2_X1 U78bar ( .A1(n194bar), .A2(n150bar), .ZN(n152bar) );
  AND2_X1 U79 ( .A1(n149), .A2(n148), .ZN(n150) );
  OR2_X1 U79bar ( .A1(n149bar), .A2(n148bar), .ZN(n150bar) );
  OR2_X1 U80 ( .A1(n217), .A2(b[4]), .ZN(n148) );
  AND2_X1 U80bar ( .A1(n217bar), .A2(bbar[4]), .ZN(n148bar) );
  OR2_X1 U81 ( .A1(n205), .A2(a[4]), .ZN(n149) );
  AND2_X1 U81bar ( .A1(n205bar), .A2(abar[4]), .ZN(n149bar) );
  AND2_X1 U82 ( .A1(n146), .A2(n145), .ZN(n147) );
  OR2_X1 U82bar ( .A1(n146bar), .A2(n145bar), .ZN(n147bar) );
  OR2_X1 U83 ( .A1(n193), .A2(d[4]), .ZN(n145) );
  AND2_X1 U83bar ( .A1(n193bar), .A2(dbar[4]), .ZN(n145bar) );
  OR2_X1 U84 ( .A1(n181), .A2(c[4]), .ZN(n146) );
  AND2_X1 U84bar ( .A1(n181bar), .A2(cbar[4]), .ZN(n146bar) );
  OR2_X1 U85 ( .A1(n144), .A2(n216), .ZN(y[3]) );
  AND2_X1 U85bar ( .A1(n144bar), .A2(n216bar), .ZN(ybar[3]) );
  OR2_X1 U86 ( .A1(n142), .A2(n192), .ZN(n143) );
  AND2_X1 U86bar ( .A1(n142bar), .A2(n192bar), .ZN(n143bar) );
  AND2_X1 U87 ( .A1(n192), .A2(n142), .ZN(n144) );
  OR2_X1 U87bar ( .A1(n192bar), .A2(n142bar), .ZN(n144bar) );
  AND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(n142) );
  OR2_X1 U88bar ( .A1(n141bar), .A2(n140bar), .ZN(n142bar) );
  OR2_X1 U89 ( .A1(n215), .A2(b[3]), .ZN(n140) );
  AND2_X1 U89bar ( .A1(n215bar), .A2(bbar[3]), .ZN(n140bar) );
  OR2_X1 U90 ( .A1(n204), .A2(a[3]), .ZN(n141) );
  AND2_X1 U90bar ( .A1(n204bar), .A2(abar[3]), .ZN(n141bar) );
  AND2_X1 U91 ( .A1(n138), .A2(n137), .ZN(n139) );
  OR2_X1 U91bar ( .A1(n138bar), .A2(n137bar), .ZN(n139bar) );
  OR2_X1 U92 ( .A1(n191), .A2(d[3]), .ZN(n137) );
  AND2_X1 U92bar ( .A1(n191bar), .A2(dbar[3]), .ZN(n137bar) );
  OR2_X1 U93 ( .A1(n180), .A2(c[3]), .ZN(n138) );
  AND2_X1 U93bar ( .A1(n180bar), .A2(cbar[3]), .ZN(n138bar) );
  OR2_X1 U94 ( .A1(n136), .A2(n214), .ZN(y[2]) );
  AND2_X1 U94bar ( .A1(n136bar), .A2(n214bar), .ZN(ybar[2]) );
  OR2_X1 U95 ( .A1(n134), .A2(n190), .ZN(n135) );
  AND2_X1 U95bar ( .A1(n134bar), .A2(n190bar), .ZN(n135bar) );
  AND2_X1 U96 ( .A1(n190), .A2(n134), .ZN(n136) );
  OR2_X1 U96bar ( .A1(n190bar), .A2(n134bar), .ZN(n136bar) );
  AND2_X1 U97 ( .A1(n133), .A2(n132), .ZN(n134) );
  OR2_X1 U97bar ( .A1(n133bar), .A2(n132bar), .ZN(n134bar) );
  OR2_X1 U98 ( .A1(n213), .A2(b[2]), .ZN(n132) );
  AND2_X1 U98bar ( .A1(n213bar), .A2(bbar[2]), .ZN(n132bar) );
  OR2_X1 U99 ( .A1(n203), .A2(a[2]), .ZN(n133) );
  AND2_X1 U99bar ( .A1(n203bar), .A2(abar[2]), .ZN(n133bar) );
  AND2_X1 U100 ( .A1(n130), .A2(n129), .ZN(n131) );
  OR2_X1 U100bar ( .A1(n130bar), .A2(n129bar), .ZN(n131bar) );
  OR2_X1 U101 ( .A1(n189), .A2(d[2]), .ZN(n129) );
  AND2_X1 U101bar ( .A1(n189bar), .A2(dbar[2]), .ZN(n129bar) );
  OR2_X1 U102 ( .A1(n179), .A2(c[2]), .ZN(n130) );
  AND2_X1 U102bar ( .A1(n179bar), .A2(cbar[2]), .ZN(n130bar) );
  OR2_X1 U103 ( .A1(n128), .A2(n212), .ZN(y[1]) );
  AND2_X1 U103bar ( .A1(n128bar), .A2(n212bar), .ZN(ybar[1]) );
  OR2_X1 U104 ( .A1(n126), .A2(n188), .ZN(n127) );
  AND2_X1 U104bar ( .A1(n126bar), .A2(n188bar), .ZN(n127bar) );
  AND2_X1 U105 ( .A1(n188), .A2(n126), .ZN(n128) );
  OR2_X1 U105bar ( .A1(n188bar), .A2(n126bar), .ZN(n128bar) );
  AND2_X1 U106 ( .A1(n125), .A2(n124), .ZN(n126) );
  OR2_X1 U106bar ( .A1(n125bar), .A2(n124bar), .ZN(n126bar) );
  OR2_X1 U107 ( .A1(n211), .A2(b[1]), .ZN(n124) );
  AND2_X1 U107bar ( .A1(n211bar), .A2(bbar[1]), .ZN(n124bar) );
  OR2_X1 U108 ( .A1(n202), .A2(a[1]), .ZN(n125) );
  AND2_X1 U108bar ( .A1(n202bar), .A2(abar[1]), .ZN(n125bar) );
  AND2_X1 U109 ( .A1(n122), .A2(n121), .ZN(n123) );
  OR2_X1 U109bar ( .A1(n122bar), .A2(n121bar), .ZN(n123bar) );
  OR2_X1 U110 ( .A1(n187), .A2(d[1]), .ZN(n121) );
  AND2_X1 U110bar ( .A1(n187bar), .A2(dbar[1]), .ZN(n121bar) );
  OR2_X1 U111 ( .A1(n178), .A2(c[1]), .ZN(n122) );
  AND2_X1 U111bar ( .A1(n178bar), .A2(cbar[1]), .ZN(n122bar) );
  OR2_X1 U112 ( .A1(n120), .A2(n210), .ZN(y[0]) );
  AND2_X1 U112bar ( .A1(n120bar), .A2(n210bar), .ZN(ybar[0]) );
  OR2_X1 U113 ( .A1(n118), .A2(n186), .ZN(n119) );
  AND2_X1 U113bar ( .A1(n118bar), .A2(n186bar), .ZN(n119bar) );
  AND2_X1 U114 ( .A1(n186), .A2(n118), .ZN(n120) );
  OR2_X1 U114bar ( .A1(n186bar), .A2(n118bar), .ZN(n120bar) );
  AND2_X1 U115 ( .A1(n117), .A2(n116), .ZN(n118) );
  OR2_X1 U115bar ( .A1(n117bar), .A2(n116bar), .ZN(n118bar) );
  OR2_X1 U116 ( .A1(n209), .A2(b[0]), .ZN(n116) );
  AND2_X1 U116bar ( .A1(n209bar), .A2(bbar[0]), .ZN(n116bar) );
  OR2_X1 U117 ( .A1(n201), .A2(a[0]), .ZN(n117) );
  AND2_X1 U117bar ( .A1(n201bar), .A2(abar[0]), .ZN(n117bar) );
  AND2_X1 U118 ( .A1(n114), .A2(n113), .ZN(n115) );
  OR2_X1 U118bar ( .A1(n114bar), .A2(n113bar), .ZN(n115bar) );
  OR2_X1 U119 ( .A1(n185), .A2(d[0]), .ZN(n113) );
  AND2_X1 U119bar ( .A1(n185bar), .A2(dbar[0]), .ZN(n113bar) );
  OR2_X1 U120 ( .A1(n177), .A2(c[0]), .ZN(n114) );
  AND2_X1 U120bar ( .A1(n177bar), .A2(cbar[0]), .ZN(n114bar) );
endmodule

module byteXor4_8 ( a, b, c, d, y );

  input wire [7:0] a;
  input wire [7:0] b;
  input wire [7:0] c;
  input wire [7:0] d;
  wire [7:0] abar;
  wire [7:0] bbar;
  wire [7:0] cbar;
  wire [7:0] dbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign cbar[0] = ~c[0];
  assign cbar[1] = ~c[1];
  assign cbar[2] = ~c[2];
  assign cbar[3] = ~c[3];
  assign cbar[4] = ~c[4];
  assign cbar[5] = ~c[5];
  assign cbar[6] = ~c[6];
  assign cbar[7] = ~c[7];
  assign dbar[0] = ~d[0];
  assign dbar[1] = ~d[1];
  assign dbar[2] = ~d[2];
  assign dbar[3] = ~d[3];
  assign dbar[4] = ~d[4];
  assign dbar[5] = ~d[5];
  assign dbar[6] = ~d[6];
  assign dbar[7] = ~d[7];
//input_done

  output wire [7:0] y;
  wire [7:0] ybar;
//output_done

  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n113bar;
  wire n114bar;
  wire n115bar;
  wire n116bar;
  wire n117bar;
  wire n118bar;
  wire n119bar;
  wire n120bar;
  wire n121bar;
  wire n122bar;
  wire n123bar;
  wire n124bar;
  wire n125bar;
  wire n126bar;
  wire n127bar;
  wire n128bar;
  wire n129bar;
  wire n130bar;
  wire n131bar;
  wire n132bar;
  wire n133bar;
  wire n134bar;
  wire n135bar;
  wire n136bar;
  wire n137bar;
  wire n138bar;
  wire n139bar;
  wire n140bar;
  wire n141bar;
  wire n142bar;
  wire n143bar;
  wire n144bar;
  wire n145bar;
  wire n146bar;
  wire n147bar;
  wire n148bar;
  wire n149bar;
  wire n150bar;
  wire n151bar;
  wire n152bar;
  wire n153bar;
  wire n154bar;
  wire n155bar;
  wire n156bar;
  wire n157bar;
  wire n158bar;
  wire n159bar;
  wire n160bar;
  wire n161bar;
  wire n162bar;
  wire n163bar;
  wire n164bar;
  wire n165bar;
  wire n166bar;
  wire n167bar;
  wire n168bar;
  wire n169bar;
  wire n170bar;
  wire n171bar;
  wire n172bar;
  wire n173bar;
  wire n174bar;
  wire n175bar;
  wire n176bar;
  wire n177bar;
  wire n178bar;
  wire n179bar;
  wire n180bar;
  wire n181bar;
  wire n182bar;
  wire n183bar;
  wire n184bar;
  wire n185bar;
  wire n186bar;
  wire n187bar;
  wire n188bar;
  wire n189bar;
  wire n190bar;
  wire n191bar;
  wire n192bar;
  wire n193bar;
  wire n194bar;
  wire n195bar;
  wire n196bar;
  wire n197bar;
  wire n198bar;
  wire n199bar;
  wire n200bar;
  wire n201bar;
  wire n202bar;
  wire n203bar;
  wire n204bar;
  wire n205bar;
  wire n206bar;
  wire n207bar;
  wire n208bar;
  wire n209bar;
  wire n210bar;
  wire n211bar;
  wire n212bar;
  wire n213bar;
  wire n214bar;
  wire n215bar;
  wire n216bar;
  wire n217bar;
  wire n218bar;
  wire n219bar;
  wire n220bar;
  wire n221bar;
  wire n222bar;
  wire n223bar;
  wire n224bar;
//wire_done

 //assign_done

  assign n224bar = n175;
  assign n224 = n175bar;
  assign n223bar = a[7];
  assign n223 = abar[7];
  assign n222bar = n167;
  assign n222 = n167bar;
  assign n221bar = a[6];
  assign n221 = abar[6];
  assign n220bar = n159;
  assign n220 = n159bar;
  assign n219bar = a[5];
  assign n219 = abar[5];
  assign n218bar = n151;
  assign n218 = n151bar;
  assign n217bar = a[4];
  assign n217 = abar[4];
  assign n216bar = n143;
  assign n216 = n143bar;
  assign n215bar = a[3];
  assign n215 = abar[3];
  assign n214bar = n135;
  assign n214 = n135bar;
  assign n213bar = a[2];
  assign n213 = abar[2];
  assign n212bar = n127;
  assign n212 = n127bar;
  assign n211bar = a[1];
  assign n211 = abar[1];
  assign n210bar = n119;
  assign n210 = n119bar;
  assign n209bar = a[0];
  assign n209 = abar[0];
  assign n208bar = b[7];
  assign n208 = bbar[7];
  assign n207bar = b[6];
  assign n207 = bbar[6];
  assign n206bar = b[5];
  assign n206 = bbar[5];
  assign n205bar = b[4];
  assign n205 = bbar[4];
  assign n204bar = b[3];
  assign n204 = bbar[3];
  assign n203bar = b[2];
  assign n203 = bbar[2];
  assign n202bar = b[1];
  assign n202 = bbar[1];
  assign n201bar = b[0];
  assign n201 = bbar[0];
  assign n200bar = n171;
  assign n200 = n171bar;
  assign n199bar = c[7];
  assign n199 = cbar[7];
  assign n198bar = n163;
  assign n198 = n163bar;
  assign n197bar = c[6];
  assign n197 = cbar[6];
  assign n196bar = n155;
  assign n196 = n155bar;
  assign n195bar = c[5];
  assign n195 = cbar[5];
  assign n194bar = n147;
  assign n194 = n147bar;
  assign n193bar = c[4];
  assign n193 = cbar[4];
  assign n192bar = n139;
  assign n192 = n139bar;
  assign n191bar = c[3];
  assign n191 = cbar[3];
  assign n190bar = n131;
  assign n190 = n131bar;
  assign n189bar = c[2];
  assign n189 = cbar[2];
  assign n188bar = n123;
  assign n188 = n123bar;
  assign n187bar = c[1];
  assign n187 = cbar[1];
  assign n186bar = n115;
  assign n186 = n115bar;
  assign n185bar = c[0];
  assign n185 = cbar[0];
  assign n184bar = d[7];
  assign n184 = dbar[7];
  assign n183bar = d[6];
  assign n183 = dbar[6];
  assign n182bar = d[5];
  assign n182 = dbar[5];
  assign n181bar = d[4];
  assign n181 = dbar[4];
  assign n180bar = d[3];
  assign n180 = dbar[3];
  assign n179bar = d[2];
  assign n179 = dbar[2];
  assign n178bar = d[1];
  assign n178 = dbar[1];
  assign n177bar = d[0];
  assign n177 = dbar[0];
  OR2_X1 U49 ( .A1(n176), .A2(n224), .ZN(y[7]) );
  AND2_X1 U49bar ( .A1(n176bar), .A2(n224bar), .ZN(ybar[7]) );
  OR2_X1 U50 ( .A1(n174), .A2(n200), .ZN(n175) );
  AND2_X1 U50bar ( .A1(n174bar), .A2(n200bar), .ZN(n175bar) );
  AND2_X1 U51 ( .A1(n200), .A2(n174), .ZN(n176) );
  OR2_X1 U51bar ( .A1(n200bar), .A2(n174bar), .ZN(n176bar) );
  AND2_X1 U52 ( .A1(n173), .A2(n172), .ZN(n174) );
  OR2_X1 U52bar ( .A1(n173bar), .A2(n172bar), .ZN(n174bar) );
  OR2_X1 U53 ( .A1(n223), .A2(b[7]), .ZN(n172) );
  AND2_X1 U53bar ( .A1(n223bar), .A2(bbar[7]), .ZN(n172bar) );
  OR2_X1 U54 ( .A1(n208), .A2(a[7]), .ZN(n173) );
  AND2_X1 U54bar ( .A1(n208bar), .A2(abar[7]), .ZN(n173bar) );
  AND2_X1 U55 ( .A1(n170), .A2(n169), .ZN(n171) );
  OR2_X1 U55bar ( .A1(n170bar), .A2(n169bar), .ZN(n171bar) );
  OR2_X1 U56 ( .A1(n199), .A2(d[7]), .ZN(n169) );
  AND2_X1 U56bar ( .A1(n199bar), .A2(dbar[7]), .ZN(n169bar) );
  OR2_X1 U57 ( .A1(n184), .A2(c[7]), .ZN(n170) );
  AND2_X1 U57bar ( .A1(n184bar), .A2(cbar[7]), .ZN(n170bar) );
  OR2_X1 U58 ( .A1(n168), .A2(n222), .ZN(y[6]) );
  AND2_X1 U58bar ( .A1(n168bar), .A2(n222bar), .ZN(ybar[6]) );
  OR2_X1 U59 ( .A1(n166), .A2(n198), .ZN(n167) );
  AND2_X1 U59bar ( .A1(n166bar), .A2(n198bar), .ZN(n167bar) );
  AND2_X1 U60 ( .A1(n198), .A2(n166), .ZN(n168) );
  OR2_X1 U60bar ( .A1(n198bar), .A2(n166bar), .ZN(n168bar) );
  AND2_X1 U61 ( .A1(n165), .A2(n164), .ZN(n166) );
  OR2_X1 U61bar ( .A1(n165bar), .A2(n164bar), .ZN(n166bar) );
  OR2_X1 U62 ( .A1(n221), .A2(b[6]), .ZN(n164) );
  AND2_X1 U62bar ( .A1(n221bar), .A2(bbar[6]), .ZN(n164bar) );
  OR2_X1 U63 ( .A1(n207), .A2(a[6]), .ZN(n165) );
  AND2_X1 U63bar ( .A1(n207bar), .A2(abar[6]), .ZN(n165bar) );
  AND2_X1 U64 ( .A1(n162), .A2(n161), .ZN(n163) );
  OR2_X1 U64bar ( .A1(n162bar), .A2(n161bar), .ZN(n163bar) );
  OR2_X1 U65 ( .A1(n197), .A2(d[6]), .ZN(n161) );
  AND2_X1 U65bar ( .A1(n197bar), .A2(dbar[6]), .ZN(n161bar) );
  OR2_X1 U66 ( .A1(n183), .A2(c[6]), .ZN(n162) );
  AND2_X1 U66bar ( .A1(n183bar), .A2(cbar[6]), .ZN(n162bar) );
  OR2_X1 U67 ( .A1(n160), .A2(n220), .ZN(y[5]) );
  AND2_X1 U67bar ( .A1(n160bar), .A2(n220bar), .ZN(ybar[5]) );
  OR2_X1 U68 ( .A1(n158), .A2(n196), .ZN(n159) );
  AND2_X1 U68bar ( .A1(n158bar), .A2(n196bar), .ZN(n159bar) );
  AND2_X1 U69 ( .A1(n196), .A2(n158), .ZN(n160) );
  OR2_X1 U69bar ( .A1(n196bar), .A2(n158bar), .ZN(n160bar) );
  AND2_X1 U70 ( .A1(n157), .A2(n156), .ZN(n158) );
  OR2_X1 U70bar ( .A1(n157bar), .A2(n156bar), .ZN(n158bar) );
  OR2_X1 U71 ( .A1(n219), .A2(b[5]), .ZN(n156) );
  AND2_X1 U71bar ( .A1(n219bar), .A2(bbar[5]), .ZN(n156bar) );
  OR2_X1 U72 ( .A1(n206), .A2(a[5]), .ZN(n157) );
  AND2_X1 U72bar ( .A1(n206bar), .A2(abar[5]), .ZN(n157bar) );
  AND2_X1 U73 ( .A1(n154), .A2(n153), .ZN(n155) );
  OR2_X1 U73bar ( .A1(n154bar), .A2(n153bar), .ZN(n155bar) );
  OR2_X1 U74 ( .A1(n195), .A2(d[5]), .ZN(n153) );
  AND2_X1 U74bar ( .A1(n195bar), .A2(dbar[5]), .ZN(n153bar) );
  OR2_X1 U75 ( .A1(n182), .A2(c[5]), .ZN(n154) );
  AND2_X1 U75bar ( .A1(n182bar), .A2(cbar[5]), .ZN(n154bar) );
  OR2_X1 U76 ( .A1(n152), .A2(n218), .ZN(y[4]) );
  AND2_X1 U76bar ( .A1(n152bar), .A2(n218bar), .ZN(ybar[4]) );
  OR2_X1 U77 ( .A1(n150), .A2(n194), .ZN(n151) );
  AND2_X1 U77bar ( .A1(n150bar), .A2(n194bar), .ZN(n151bar) );
  AND2_X1 U78 ( .A1(n194), .A2(n150), .ZN(n152) );
  OR2_X1 U78bar ( .A1(n194bar), .A2(n150bar), .ZN(n152bar) );
  AND2_X1 U79 ( .A1(n149), .A2(n148), .ZN(n150) );
  OR2_X1 U79bar ( .A1(n149bar), .A2(n148bar), .ZN(n150bar) );
  OR2_X1 U80 ( .A1(n217), .A2(b[4]), .ZN(n148) );
  AND2_X1 U80bar ( .A1(n217bar), .A2(bbar[4]), .ZN(n148bar) );
  OR2_X1 U81 ( .A1(n205), .A2(a[4]), .ZN(n149) );
  AND2_X1 U81bar ( .A1(n205bar), .A2(abar[4]), .ZN(n149bar) );
  AND2_X1 U82 ( .A1(n146), .A2(n145), .ZN(n147) );
  OR2_X1 U82bar ( .A1(n146bar), .A2(n145bar), .ZN(n147bar) );
  OR2_X1 U83 ( .A1(n193), .A2(d[4]), .ZN(n145) );
  AND2_X1 U83bar ( .A1(n193bar), .A2(dbar[4]), .ZN(n145bar) );
  OR2_X1 U84 ( .A1(n181), .A2(c[4]), .ZN(n146) );
  AND2_X1 U84bar ( .A1(n181bar), .A2(cbar[4]), .ZN(n146bar) );
  OR2_X1 U85 ( .A1(n144), .A2(n216), .ZN(y[3]) );
  AND2_X1 U85bar ( .A1(n144bar), .A2(n216bar), .ZN(ybar[3]) );
  OR2_X1 U86 ( .A1(n142), .A2(n192), .ZN(n143) );
  AND2_X1 U86bar ( .A1(n142bar), .A2(n192bar), .ZN(n143bar) );
  AND2_X1 U87 ( .A1(n192), .A2(n142), .ZN(n144) );
  OR2_X1 U87bar ( .A1(n192bar), .A2(n142bar), .ZN(n144bar) );
  AND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(n142) );
  OR2_X1 U88bar ( .A1(n141bar), .A2(n140bar), .ZN(n142bar) );
  OR2_X1 U89 ( .A1(n215), .A2(b[3]), .ZN(n140) );
  AND2_X1 U89bar ( .A1(n215bar), .A2(bbar[3]), .ZN(n140bar) );
  OR2_X1 U90 ( .A1(n204), .A2(a[3]), .ZN(n141) );
  AND2_X1 U90bar ( .A1(n204bar), .A2(abar[3]), .ZN(n141bar) );
  AND2_X1 U91 ( .A1(n138), .A2(n137), .ZN(n139) );
  OR2_X1 U91bar ( .A1(n138bar), .A2(n137bar), .ZN(n139bar) );
  OR2_X1 U92 ( .A1(n191), .A2(d[3]), .ZN(n137) );
  AND2_X1 U92bar ( .A1(n191bar), .A2(dbar[3]), .ZN(n137bar) );
  OR2_X1 U93 ( .A1(n180), .A2(c[3]), .ZN(n138) );
  AND2_X1 U93bar ( .A1(n180bar), .A2(cbar[3]), .ZN(n138bar) );
  OR2_X1 U94 ( .A1(n136), .A2(n214), .ZN(y[2]) );
  AND2_X1 U94bar ( .A1(n136bar), .A2(n214bar), .ZN(ybar[2]) );
  OR2_X1 U95 ( .A1(n134), .A2(n190), .ZN(n135) );
  AND2_X1 U95bar ( .A1(n134bar), .A2(n190bar), .ZN(n135bar) );
  AND2_X1 U96 ( .A1(n190), .A2(n134), .ZN(n136) );
  OR2_X1 U96bar ( .A1(n190bar), .A2(n134bar), .ZN(n136bar) );
  AND2_X1 U97 ( .A1(n133), .A2(n132), .ZN(n134) );
  OR2_X1 U97bar ( .A1(n133bar), .A2(n132bar), .ZN(n134bar) );
  OR2_X1 U98 ( .A1(n213), .A2(b[2]), .ZN(n132) );
  AND2_X1 U98bar ( .A1(n213bar), .A2(bbar[2]), .ZN(n132bar) );
  OR2_X1 U99 ( .A1(n203), .A2(a[2]), .ZN(n133) );
  AND2_X1 U99bar ( .A1(n203bar), .A2(abar[2]), .ZN(n133bar) );
  AND2_X1 U100 ( .A1(n130), .A2(n129), .ZN(n131) );
  OR2_X1 U100bar ( .A1(n130bar), .A2(n129bar), .ZN(n131bar) );
  OR2_X1 U101 ( .A1(n189), .A2(d[2]), .ZN(n129) );
  AND2_X1 U101bar ( .A1(n189bar), .A2(dbar[2]), .ZN(n129bar) );
  OR2_X1 U102 ( .A1(n179), .A2(c[2]), .ZN(n130) );
  AND2_X1 U102bar ( .A1(n179bar), .A2(cbar[2]), .ZN(n130bar) );
  OR2_X1 U103 ( .A1(n128), .A2(n212), .ZN(y[1]) );
  AND2_X1 U103bar ( .A1(n128bar), .A2(n212bar), .ZN(ybar[1]) );
  OR2_X1 U104 ( .A1(n126), .A2(n188), .ZN(n127) );
  AND2_X1 U104bar ( .A1(n126bar), .A2(n188bar), .ZN(n127bar) );
  AND2_X1 U105 ( .A1(n188), .A2(n126), .ZN(n128) );
  OR2_X1 U105bar ( .A1(n188bar), .A2(n126bar), .ZN(n128bar) );
  AND2_X1 U106 ( .A1(n125), .A2(n124), .ZN(n126) );
  OR2_X1 U106bar ( .A1(n125bar), .A2(n124bar), .ZN(n126bar) );
  OR2_X1 U107 ( .A1(n211), .A2(b[1]), .ZN(n124) );
  AND2_X1 U107bar ( .A1(n211bar), .A2(bbar[1]), .ZN(n124bar) );
  OR2_X1 U108 ( .A1(n202), .A2(a[1]), .ZN(n125) );
  AND2_X1 U108bar ( .A1(n202bar), .A2(abar[1]), .ZN(n125bar) );
  AND2_X1 U109 ( .A1(n122), .A2(n121), .ZN(n123) );
  OR2_X1 U109bar ( .A1(n122bar), .A2(n121bar), .ZN(n123bar) );
  OR2_X1 U110 ( .A1(n187), .A2(d[1]), .ZN(n121) );
  AND2_X1 U110bar ( .A1(n187bar), .A2(dbar[1]), .ZN(n121bar) );
  OR2_X1 U111 ( .A1(n178), .A2(c[1]), .ZN(n122) );
  AND2_X1 U111bar ( .A1(n178bar), .A2(cbar[1]), .ZN(n122bar) );
  OR2_X1 U112 ( .A1(n120), .A2(n210), .ZN(y[0]) );
  AND2_X1 U112bar ( .A1(n120bar), .A2(n210bar), .ZN(ybar[0]) );
  OR2_X1 U113 ( .A1(n118), .A2(n186), .ZN(n119) );
  AND2_X1 U113bar ( .A1(n118bar), .A2(n186bar), .ZN(n119bar) );
  AND2_X1 U114 ( .A1(n186), .A2(n118), .ZN(n120) );
  OR2_X1 U114bar ( .A1(n186bar), .A2(n118bar), .ZN(n120bar) );
  AND2_X1 U115 ( .A1(n117), .A2(n116), .ZN(n118) );
  OR2_X1 U115bar ( .A1(n117bar), .A2(n116bar), .ZN(n118bar) );
  OR2_X1 U116 ( .A1(n209), .A2(b[0]), .ZN(n116) );
  AND2_X1 U116bar ( .A1(n209bar), .A2(bbar[0]), .ZN(n116bar) );
  OR2_X1 U117 ( .A1(n201), .A2(a[0]), .ZN(n117) );
  AND2_X1 U117bar ( .A1(n201bar), .A2(abar[0]), .ZN(n117bar) );
  AND2_X1 U118 ( .A1(n114), .A2(n113), .ZN(n115) );
  OR2_X1 U118bar ( .A1(n114bar), .A2(n113bar), .ZN(n115bar) );
  OR2_X1 U119 ( .A1(n185), .A2(d[0]), .ZN(n113) );
  AND2_X1 U119bar ( .A1(n185bar), .A2(dbar[0]), .ZN(n113bar) );
  OR2_X1 U120 ( .A1(n177), .A2(c[0]), .ZN(n114) );
  AND2_X1 U120bar ( .A1(n177bar), .A2(cbar[0]), .ZN(n114bar) );
endmodule

module mixCol_2 ( in, out );

  input wire [31:0] in;
//input_done

  output wire [31:0] out;
//output_done

  wire [7:0] b0_s2;
  wire [7:0] b1_s2;
  wire [7:0] b2_s2;
  wire [7:0] b3_s2;
  wire [7:0] b0_s3;
  wire [7:0] b1_s3;
  wire [7:0] b2_s3;
  wire [7:0] b3_s3;
//wire_done

 //assign_done

  scale2_8 b0_scale2 ( .in(in[31:24]), .out(b0_s2) );
  scale2_7 b1_scale2 ( .in(in[23:16]), .out(b1_s2) );
  scale2_6 b2_scale2 ( .in(in[15:8]), .out(b2_s2) );
  scale2_5 b3_scale2 ( .in(in[7:0]), .out(b3_s2) );
  byteXor_9 b0_scale3 ( .a(in[31:24]), .b(b0_s2), .y(b0_s3) );
  byteXor_8 b1_scale3 ( .a(in[23:16]), .b(b1_s2), .y(b1_s3) );
  byteXor_7 b2_scale3 ( .a(in[15:8]), .b(b2_s2), .y(b2_s3) );
  byteXor_6 b3_scale3 ( .a(in[7:0]), .b(b3_s2), .y(b3_s3) );
  byteXor4_8 out0 ( .a(b0_s2), .b(b1_s3), .c(in[15:8]), .d(in[7:0]), .y(
        out[31:24]) );
  byteXor4_7 out1 ( .a(in[31:24]), .b(b1_s2), .c(b2_s3), .d(in[7:0]), .y(
        out[23:16]) );
  byteXor4_6 out2 ( .a(in[31:24]), .b(in[23:16]), .c(b2_s2), .d(b3_s3), .y(
        out[15:8]) );
  byteXor4_5 out3 ( .a(b0_s3), .b(in[23:16]), .c(in[15:8]), .d(b3_s2), .y(
        out[7:0]) );
endmodule

module scale2_9 ( in, out );

  input wire [7:0] in;
  wire [7:0] inbar;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
//input_done

  output wire [7:0] out;
  wire [7:0] outbar;
//output_done

  wire in_0;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_1;
  wire in_7;
  wire n11;
  wire n12;
  wire n13;
  wire n14;
  wire n15;
  wire n16;
  wire n17;
  wire n18;
  wire n19;
  wire n20;
  wire in_0bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_1bar;
  wire in_7bar;
  wire n11bar;
  wire n12bar;
  wire n13bar;
  wire n14bar;
  wire n15bar;
  wire n16bar;
  wire n17bar;
  wire n18bar;
  wire n19bar;
  wire n20bar;
//wire_done

  assign in_0 = in[0];
  assign out[7] = in_6;
  assign in_6  = in[6];
  assign out[6] = in_5;
  assign in_5  = in[5];
  assign out[5] = in_4;
  assign in_4  = in[4];
  assign out[2] = in_1;
  assign in_1  = in[1];
  assign out[0] = in_7;
  assign in_7  = in[7];
  assign in_0bar = inbar[0];
  assign outbar[7] = in_6bar;
  assign in_6bar = inbar[6];
  assign outbar[6] = in_5bar;
  assign in_5bar = inbar[5];
  assign outbar[5] = in_4bar;
  assign in_4bar = inbar[4];
  assign outbar[2] = in_1bar;
  assign in_1bar = inbar[1];
  assign outbar[0] = in_7bar;
  assign in_7bar = inbar[7];
//assign_done

  assign n20bar = in_7;
  assign n20 = in_7bar;
  assign n19bar = in[3];
  assign n19 = inbar[3];
  assign n18bar = in[2];
  assign n18 = inbar[2];
  assign n17bar = in_0;
  assign n17 = in_0bar;
  OR2_X1 U5 ( .A1(n16), .A2(n15), .ZN(out[4]) );
  AND2_X1 U5bar ( .A1(n16bar), .A2(n15bar), .ZN(outbar[4]) );
  AND2_X1 U6 ( .A1(in[3]), .A2(n20), .ZN(n15) );
  OR2_X1 U6bar ( .A1(inbar[3]), .A2(n20bar), .ZN(n15bar) );
  AND2_X1 U7 ( .A1(in_7), .A2(n19), .ZN(n16) );
  OR2_X1 U7bar ( .A1(in_7bar), .A2(n19bar), .ZN(n16bar) );
  OR2_X1 U8 ( .A1(n14), .A2(n13), .ZN(out[3]) );
  AND2_X1 U8bar ( .A1(n14bar), .A2(n13bar), .ZN(outbar[3]) );
  AND2_X1 U9 ( .A1(in[2]), .A2(n20), .ZN(n13) );
  OR2_X1 U9bar ( .A1(inbar[2]), .A2(n20bar), .ZN(n13bar) );
  AND2_X1 U10 ( .A1(in_7), .A2(n18), .ZN(n14) );
  OR2_X1 U10bar ( .A1(in_7bar), .A2(n18bar), .ZN(n14bar) );
  OR2_X1 U11 ( .A1(n12), .A2(n11), .ZN(out[1]) );
  AND2_X1 U11bar ( .A1(n12bar), .A2(n11bar), .ZN(outbar[1]) );
  AND2_X1 U12 ( .A1(in_0), .A2(n20), .ZN(n11) );
  OR2_X1 U12bar ( .A1(in_0bar), .A2(n20bar), .ZN(n11bar) );
  AND2_X1 U13 ( .A1(in_7), .A2(n17), .ZN(n12) );
  OR2_X1 U13bar ( .A1(in_7bar), .A2(n17bar), .ZN(n12bar) );
endmodule

module scale2_10 ( in, out );

  input wire [7:0] in;
  wire [7:0] inbar;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
//input_done

  output wire [7:0] out;
  wire [7:0] outbar;
//output_done

  wire in_0;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_1;
  wire in_7;
  wire n11;
  wire n12;
  wire n13;
  wire n14;
  wire n15;
  wire n16;
  wire n17;
  wire n18;
  wire n19;
  wire n20;
  wire in_0bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_1bar;
  wire in_7bar;
  wire n11bar;
  wire n12bar;
  wire n13bar;
  wire n14bar;
  wire n15bar;
  wire n16bar;
  wire n17bar;
  wire n18bar;
  wire n19bar;
  wire n20bar;
//wire_done

  assign in_0 = in[0];
  assign out[7] = in_6;
  assign in_6  = in[6];
  assign out[6] = in_5;
  assign in_5  = in[5];
  assign out[5] = in_4;
  assign in_4  = in[4];
  assign out[2] = in_1;
  assign in_1  = in[1];
  assign out[0] = in_7;
  assign in_7  = in[7];
  assign in_0bar = inbar[0];
  assign outbar[7] = in_6bar;
  assign in_6bar = inbar[6];
  assign outbar[6] = in_5bar;
  assign in_5bar = inbar[5];
  assign outbar[5] = in_4bar;
  assign in_4bar = inbar[4];
  assign outbar[2] = in_1bar;
  assign in_1bar = inbar[1];
  assign outbar[0] = in_7bar;
  assign in_7bar = inbar[7];
//assign_done

  assign n20bar = in_7;
  assign n20 = in_7bar;
  assign n19bar = in[3];
  assign n19 = inbar[3];
  assign n18bar = in[2];
  assign n18 = inbar[2];
  assign n17bar = in_0;
  assign n17 = in_0bar;
  OR2_X1 U5 ( .A1(n16), .A2(n15), .ZN(out[4]) );
  AND2_X1 U5bar ( .A1(n16bar), .A2(n15bar), .ZN(outbar[4]) );
  AND2_X1 U6 ( .A1(in[3]), .A2(n20), .ZN(n15) );
  OR2_X1 U6bar ( .A1(inbar[3]), .A2(n20bar), .ZN(n15bar) );
  AND2_X1 U7 ( .A1(in_7), .A2(n19), .ZN(n16) );
  OR2_X1 U7bar ( .A1(in_7bar), .A2(n19bar), .ZN(n16bar) );
  OR2_X1 U8 ( .A1(n14), .A2(n13), .ZN(out[3]) );
  AND2_X1 U8bar ( .A1(n14bar), .A2(n13bar), .ZN(outbar[3]) );
  AND2_X1 U9 ( .A1(in[2]), .A2(n20), .ZN(n13) );
  OR2_X1 U9bar ( .A1(inbar[2]), .A2(n20bar), .ZN(n13bar) );
  AND2_X1 U10 ( .A1(in_7), .A2(n18), .ZN(n14) );
  OR2_X1 U10bar ( .A1(in_7bar), .A2(n18bar), .ZN(n14bar) );
  OR2_X1 U11 ( .A1(n12), .A2(n11), .ZN(out[1]) );
  AND2_X1 U11bar ( .A1(n12bar), .A2(n11bar), .ZN(outbar[1]) );
  AND2_X1 U12 ( .A1(in_0), .A2(n20), .ZN(n11) );
  OR2_X1 U12bar ( .A1(in_0bar), .A2(n20bar), .ZN(n11bar) );
  AND2_X1 U13 ( .A1(in_7), .A2(n17), .ZN(n12) );
  OR2_X1 U13bar ( .A1(in_7bar), .A2(n17bar), .ZN(n12bar) );
endmodule

module scale2_11 ( in, out );

  input wire [7:0] in;
  wire [7:0] inbar;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
//input_done

  output wire [7:0] out;
  wire [7:0] outbar;
//output_done

  wire in_0;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_1;
  wire in_7;
  wire n11;
  wire n12;
  wire n13;
  wire n14;
  wire n15;
  wire n16;
  wire n17;
  wire n18;
  wire n19;
  wire n20;
  wire in_0bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_1bar;
  wire in_7bar;
  wire n11bar;
  wire n12bar;
  wire n13bar;
  wire n14bar;
  wire n15bar;
  wire n16bar;
  wire n17bar;
  wire n18bar;
  wire n19bar;
  wire n20bar;
//wire_done

  assign in_0 = in[0];
  assign out[7] = in_6;
  assign in_6  = in[6];
  assign out[6] = in_5;
  assign in_5  = in[5];
  assign out[5] = in_4;
  assign in_4  = in[4];
  assign out[2] = in_1;
  assign in_1  = in[1];
  assign out[0] = in_7;
  assign in_7  = in[7];
  assign in_0bar = inbar[0];
  assign outbar[7] = in_6bar;
  assign in_6bar = inbar[6];
  assign outbar[6] = in_5bar;
  assign in_5bar = inbar[5];
  assign outbar[5] = in_4bar;
  assign in_4bar = inbar[4];
  assign outbar[2] = in_1bar;
  assign in_1bar = inbar[1];
  assign outbar[0] = in_7bar;
  assign in_7bar = inbar[7];
//assign_done

  assign n20bar = in_7;
  assign n20 = in_7bar;
  assign n19bar = in[3];
  assign n19 = inbar[3];
  assign n18bar = in[2];
  assign n18 = inbar[2];
  assign n17bar = in_0;
  assign n17 = in_0bar;
  OR2_X1 U5 ( .A1(n16), .A2(n15), .ZN(out[4]) );
  AND2_X1 U5bar ( .A1(n16bar), .A2(n15bar), .ZN(outbar[4]) );
  AND2_X1 U6 ( .A1(in[3]), .A2(n20), .ZN(n15) );
  OR2_X1 U6bar ( .A1(inbar[3]), .A2(n20bar), .ZN(n15bar) );
  AND2_X1 U7 ( .A1(in_7), .A2(n19), .ZN(n16) );
  OR2_X1 U7bar ( .A1(in_7bar), .A2(n19bar), .ZN(n16bar) );
  OR2_X1 U8 ( .A1(n14), .A2(n13), .ZN(out[3]) );
  AND2_X1 U8bar ( .A1(n14bar), .A2(n13bar), .ZN(outbar[3]) );
  AND2_X1 U9 ( .A1(in[2]), .A2(n20), .ZN(n13) );
  OR2_X1 U9bar ( .A1(inbar[2]), .A2(n20bar), .ZN(n13bar) );
  AND2_X1 U10 ( .A1(in_7), .A2(n18), .ZN(n14) );
  OR2_X1 U10bar ( .A1(in_7bar), .A2(n18bar), .ZN(n14bar) );
  OR2_X1 U11 ( .A1(n12), .A2(n11), .ZN(out[1]) );
  AND2_X1 U11bar ( .A1(n12bar), .A2(n11bar), .ZN(outbar[1]) );
  AND2_X1 U12 ( .A1(in_0), .A2(n20), .ZN(n11) );
  OR2_X1 U12bar ( .A1(in_0bar), .A2(n20bar), .ZN(n11bar) );
  AND2_X1 U13 ( .A1(in_7), .A2(n17), .ZN(n12) );
  OR2_X1 U13bar ( .A1(in_7bar), .A2(n17bar), .ZN(n12bar) );
endmodule

module scale2_12 ( in, out );

  input wire [7:0] in;
  wire [7:0] inbar;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
//input_done

  output wire [7:0] out;
  wire [7:0] outbar;
//output_done

  wire in_0;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_1;
  wire in_7;
  wire n11;
  wire n12;
  wire n13;
  wire n14;
  wire n15;
  wire n16;
  wire n17;
  wire n18;
  wire n19;
  wire n20;
  wire in_0bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_1bar;
  wire in_7bar;
  wire n11bar;
  wire n12bar;
  wire n13bar;
  wire n14bar;
  wire n15bar;
  wire n16bar;
  wire n17bar;
  wire n18bar;
  wire n19bar;
  wire n20bar;
//wire_done

  assign in_0 = in[0];
  assign out[7] = in_6;
  assign in_6  = in[6];
  assign out[6] = in_5;
  assign in_5  = in[5];
  assign out[5] = in_4;
  assign in_4  = in[4];
  assign out[2] = in_1;
  assign in_1  = in[1];
  assign out[0] = in_7;
  assign in_7  = in[7];
  assign in_0bar = inbar[0];
  assign outbar[7] = in_6bar;
  assign in_6bar = inbar[6];
  assign outbar[6] = in_5bar;
  assign in_5bar = inbar[5];
  assign outbar[5] = in_4bar;
  assign in_4bar = inbar[4];
  assign outbar[2] = in_1bar;
  assign in_1bar = inbar[1];
  assign outbar[0] = in_7bar;
  assign in_7bar = inbar[7];
//assign_done

  assign n20bar = in_7;
  assign n20 = in_7bar;
  assign n19bar = in[3];
  assign n19 = inbar[3];
  assign n18bar = in[2];
  assign n18 = inbar[2];
  assign n17bar = in_0;
  assign n17 = in_0bar;
  OR2_X1 U5 ( .A1(n16), .A2(n15), .ZN(out[4]) );
  AND2_X1 U5bar ( .A1(n16bar), .A2(n15bar), .ZN(outbar[4]) );
  AND2_X1 U6 ( .A1(in[3]), .A2(n20), .ZN(n15) );
  OR2_X1 U6bar ( .A1(inbar[3]), .A2(n20bar), .ZN(n15bar) );
  AND2_X1 U7 ( .A1(in_7), .A2(n19), .ZN(n16) );
  OR2_X1 U7bar ( .A1(in_7bar), .A2(n19bar), .ZN(n16bar) );
  OR2_X1 U8 ( .A1(n14), .A2(n13), .ZN(out[3]) );
  AND2_X1 U8bar ( .A1(n14bar), .A2(n13bar), .ZN(outbar[3]) );
  AND2_X1 U9 ( .A1(in[2]), .A2(n20), .ZN(n13) );
  OR2_X1 U9bar ( .A1(inbar[2]), .A2(n20bar), .ZN(n13bar) );
  AND2_X1 U10 ( .A1(in_7), .A2(n18), .ZN(n14) );
  OR2_X1 U10bar ( .A1(in_7bar), .A2(n18bar), .ZN(n14bar) );
  OR2_X1 U11 ( .A1(n12), .A2(n11), .ZN(out[1]) );
  AND2_X1 U11bar ( .A1(n12bar), .A2(n11bar), .ZN(outbar[1]) );
  AND2_X1 U12 ( .A1(in_0), .A2(n20), .ZN(n11) );
  OR2_X1 U12bar ( .A1(in_0bar), .A2(n20bar), .ZN(n11bar) );
  AND2_X1 U13 ( .A1(in_7), .A2(n17), .ZN(n12) );
  OR2_X1 U13bar ( .A1(in_7bar), .A2(n17bar), .ZN(n12bar) );
endmodule

module byteXor_10 ( a, b, y );

  input wire [7:0] a;
  input wire [7:0] b;
  wire [7:0] abar;
  wire [7:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
//input_done

  output wire [7:0] y;
  wire [7:0] ybar;
//output_done

  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n33bar;
  wire n34bar;
  wire n35bar;
  wire n36bar;
  wire n37bar;
  wire n38bar;
  wire n39bar;
  wire n40bar;
  wire n41bar;
  wire n42bar;
  wire n43bar;
  wire n44bar;
  wire n45bar;
  wire n46bar;
  wire n47bar;
  wire n48bar;
  wire n49bar;
  wire n50bar;
  wire n51bar;
  wire n52bar;
  wire n53bar;
  wire n54bar;
  wire n55bar;
  wire n56bar;
  wire n57bar;
  wire n58bar;
  wire n59bar;
  wire n60bar;
  wire n61bar;
  wire n62bar;
  wire n63bar;
  wire n64bar;
//wire_done

 //assign_done

  assign n64bar = n47;
  assign n64 = n47bar;
  assign n63bar = a[7];
  assign n63 = abar[7];
  assign n62bar = n45;
  assign n62 = n45bar;
  assign n61bar = a[6];
  assign n61 = abar[6];
  assign n60bar = n43;
  assign n60 = n43bar;
  assign n59bar = a[5];
  assign n59 = abar[5];
  assign n58bar = n41;
  assign n58 = n41bar;
  assign n57bar = a[4];
  assign n57 = abar[4];
  assign n56bar = n39;
  assign n56 = n39bar;
  assign n55bar = a[3];
  assign n55 = abar[3];
  assign n54bar = n37;
  assign n54 = n37bar;
  assign n53bar = a[2];
  assign n53 = abar[2];
  assign n52bar = n35;
  assign n52 = n35bar;
  assign n51bar = a[1];
  assign n51 = abar[1];
  assign n50bar = n33;
  assign n50 = n33bar;
  assign n49bar = a[0];
  assign n49 = abar[0];
  OR2_X1 U17 ( .A1(n48), .A2(n64), .ZN(y[7]) );
  AND2_X1 U17bar ( .A1(n48bar), .A2(n64bar), .ZN(ybar[7]) );
  OR2_X1 U18 ( .A1(n63), .A2(b[7]), .ZN(n47) );
  AND2_X1 U18bar ( .A1(n63bar), .A2(bbar[7]), .ZN(n47bar) );
  AND2_X1 U19 ( .A1(b[7]), .A2(n63), .ZN(n48) );
  OR2_X1 U19bar ( .A1(bbar[7]), .A2(n63bar), .ZN(n48bar) );
  OR2_X1 U20 ( .A1(n46), .A2(n62), .ZN(y[6]) );
  AND2_X1 U20bar ( .A1(n46bar), .A2(n62bar), .ZN(ybar[6]) );
  OR2_X1 U21 ( .A1(n61), .A2(b[6]), .ZN(n45) );
  AND2_X1 U21bar ( .A1(n61bar), .A2(bbar[6]), .ZN(n45bar) );
  AND2_X1 U22 ( .A1(b[6]), .A2(n61), .ZN(n46) );
  OR2_X1 U22bar ( .A1(bbar[6]), .A2(n61bar), .ZN(n46bar) );
  OR2_X1 U23 ( .A1(n44), .A2(n60), .ZN(y[5]) );
  AND2_X1 U23bar ( .A1(n44bar), .A2(n60bar), .ZN(ybar[5]) );
  OR2_X1 U24 ( .A1(n59), .A2(b[5]), .ZN(n43) );
  AND2_X1 U24bar ( .A1(n59bar), .A2(bbar[5]), .ZN(n43bar) );
  AND2_X1 U25 ( .A1(b[5]), .A2(n59), .ZN(n44) );
  OR2_X1 U25bar ( .A1(bbar[5]), .A2(n59bar), .ZN(n44bar) );
  OR2_X1 U26 ( .A1(n42), .A2(n58), .ZN(y[4]) );
  AND2_X1 U26bar ( .A1(n42bar), .A2(n58bar), .ZN(ybar[4]) );
  OR2_X1 U27 ( .A1(n57), .A2(b[4]), .ZN(n41) );
  AND2_X1 U27bar ( .A1(n57bar), .A2(bbar[4]), .ZN(n41bar) );
  AND2_X1 U28 ( .A1(b[4]), .A2(n57), .ZN(n42) );
  OR2_X1 U28bar ( .A1(bbar[4]), .A2(n57bar), .ZN(n42bar) );
  OR2_X1 U29 ( .A1(n40), .A2(n56), .ZN(y[3]) );
  AND2_X1 U29bar ( .A1(n40bar), .A2(n56bar), .ZN(ybar[3]) );
  OR2_X1 U30 ( .A1(n55), .A2(b[3]), .ZN(n39) );
  AND2_X1 U30bar ( .A1(n55bar), .A2(bbar[3]), .ZN(n39bar) );
  AND2_X1 U31 ( .A1(b[3]), .A2(n55), .ZN(n40) );
  OR2_X1 U31bar ( .A1(bbar[3]), .A2(n55bar), .ZN(n40bar) );
  OR2_X1 U32 ( .A1(n38), .A2(n54), .ZN(y[2]) );
  AND2_X1 U32bar ( .A1(n38bar), .A2(n54bar), .ZN(ybar[2]) );
  OR2_X1 U33 ( .A1(n53), .A2(b[2]), .ZN(n37) );
  AND2_X1 U33bar ( .A1(n53bar), .A2(bbar[2]), .ZN(n37bar) );
  AND2_X1 U34 ( .A1(b[2]), .A2(n53), .ZN(n38) );
  OR2_X1 U34bar ( .A1(bbar[2]), .A2(n53bar), .ZN(n38bar) );
  OR2_X1 U35 ( .A1(n36), .A2(n52), .ZN(y[1]) );
  AND2_X1 U35bar ( .A1(n36bar), .A2(n52bar), .ZN(ybar[1]) );
  OR2_X1 U36 ( .A1(n51), .A2(b[1]), .ZN(n35) );
  AND2_X1 U36bar ( .A1(n51bar), .A2(bbar[1]), .ZN(n35bar) );
  AND2_X1 U37 ( .A1(b[1]), .A2(n51), .ZN(n36) );
  OR2_X1 U37bar ( .A1(bbar[1]), .A2(n51bar), .ZN(n36bar) );
  OR2_X1 U38 ( .A1(n34), .A2(n50), .ZN(y[0]) );
  AND2_X1 U38bar ( .A1(n34bar), .A2(n50bar), .ZN(ybar[0]) );
  OR2_X1 U39 ( .A1(n49), .A2(b[0]), .ZN(n33) );
  AND2_X1 U39bar ( .A1(n49bar), .A2(bbar[0]), .ZN(n33bar) );
  AND2_X1 U40 ( .A1(b[0]), .A2(n49), .ZN(n34) );
  OR2_X1 U40bar ( .A1(bbar[0]), .A2(n49bar), .ZN(n34bar) );
endmodule

module byteXor_11 ( a, b, y );

  input wire [7:0] a;
  input wire [7:0] b;
  wire [7:0] abar;
  wire [7:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
//input_done

  output wire [7:0] y;
  wire [7:0] ybar;
//output_done

  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n33bar;
  wire n34bar;
  wire n35bar;
  wire n36bar;
  wire n37bar;
  wire n38bar;
  wire n39bar;
  wire n40bar;
  wire n41bar;
  wire n42bar;
  wire n43bar;
  wire n44bar;
  wire n45bar;
  wire n46bar;
  wire n47bar;
  wire n48bar;
  wire n49bar;
  wire n50bar;
  wire n51bar;
  wire n52bar;
  wire n53bar;
  wire n54bar;
  wire n55bar;
  wire n56bar;
  wire n57bar;
  wire n58bar;
  wire n59bar;
  wire n60bar;
  wire n61bar;
  wire n62bar;
  wire n63bar;
  wire n64bar;
//wire_done

 //assign_done

  assign n64bar = n47;
  assign n64 = n47bar;
  assign n63bar = a[7];
  assign n63 = abar[7];
  assign n62bar = n45;
  assign n62 = n45bar;
  assign n61bar = a[6];
  assign n61 = abar[6];
  assign n60bar = n43;
  assign n60 = n43bar;
  assign n59bar = a[5];
  assign n59 = abar[5];
  assign n58bar = n41;
  assign n58 = n41bar;
  assign n57bar = a[4];
  assign n57 = abar[4];
  assign n56bar = n39;
  assign n56 = n39bar;
  assign n55bar = a[3];
  assign n55 = abar[3];
  assign n54bar = n37;
  assign n54 = n37bar;
  assign n53bar = a[2];
  assign n53 = abar[2];
  assign n52bar = n35;
  assign n52 = n35bar;
  assign n51bar = a[1];
  assign n51 = abar[1];
  assign n50bar = n33;
  assign n50 = n33bar;
  assign n49bar = a[0];
  assign n49 = abar[0];
  OR2_X1 U17 ( .A1(n48), .A2(n64), .ZN(y[7]) );
  AND2_X1 U17bar ( .A1(n48bar), .A2(n64bar), .ZN(ybar[7]) );
  OR2_X1 U18 ( .A1(n63), .A2(b[7]), .ZN(n47) );
  AND2_X1 U18bar ( .A1(n63bar), .A2(bbar[7]), .ZN(n47bar) );
  AND2_X1 U19 ( .A1(b[7]), .A2(n63), .ZN(n48) );
  OR2_X1 U19bar ( .A1(bbar[7]), .A2(n63bar), .ZN(n48bar) );
  OR2_X1 U20 ( .A1(n46), .A2(n62), .ZN(y[6]) );
  AND2_X1 U20bar ( .A1(n46bar), .A2(n62bar), .ZN(ybar[6]) );
  OR2_X1 U21 ( .A1(n61), .A2(b[6]), .ZN(n45) );
  AND2_X1 U21bar ( .A1(n61bar), .A2(bbar[6]), .ZN(n45bar) );
  AND2_X1 U22 ( .A1(b[6]), .A2(n61), .ZN(n46) );
  OR2_X1 U22bar ( .A1(bbar[6]), .A2(n61bar), .ZN(n46bar) );
  OR2_X1 U23 ( .A1(n44), .A2(n60), .ZN(y[5]) );
  AND2_X1 U23bar ( .A1(n44bar), .A2(n60bar), .ZN(ybar[5]) );
  OR2_X1 U24 ( .A1(n59), .A2(b[5]), .ZN(n43) );
  AND2_X1 U24bar ( .A1(n59bar), .A2(bbar[5]), .ZN(n43bar) );
  AND2_X1 U25 ( .A1(b[5]), .A2(n59), .ZN(n44) );
  OR2_X1 U25bar ( .A1(bbar[5]), .A2(n59bar), .ZN(n44bar) );
  OR2_X1 U26 ( .A1(n42), .A2(n58), .ZN(y[4]) );
  AND2_X1 U26bar ( .A1(n42bar), .A2(n58bar), .ZN(ybar[4]) );
  OR2_X1 U27 ( .A1(n57), .A2(b[4]), .ZN(n41) );
  AND2_X1 U27bar ( .A1(n57bar), .A2(bbar[4]), .ZN(n41bar) );
  AND2_X1 U28 ( .A1(b[4]), .A2(n57), .ZN(n42) );
  OR2_X1 U28bar ( .A1(bbar[4]), .A2(n57bar), .ZN(n42bar) );
  OR2_X1 U29 ( .A1(n40), .A2(n56), .ZN(y[3]) );
  AND2_X1 U29bar ( .A1(n40bar), .A2(n56bar), .ZN(ybar[3]) );
  OR2_X1 U30 ( .A1(n55), .A2(b[3]), .ZN(n39) );
  AND2_X1 U30bar ( .A1(n55bar), .A2(bbar[3]), .ZN(n39bar) );
  AND2_X1 U31 ( .A1(b[3]), .A2(n55), .ZN(n40) );
  OR2_X1 U31bar ( .A1(bbar[3]), .A2(n55bar), .ZN(n40bar) );
  OR2_X1 U32 ( .A1(n38), .A2(n54), .ZN(y[2]) );
  AND2_X1 U32bar ( .A1(n38bar), .A2(n54bar), .ZN(ybar[2]) );
  OR2_X1 U33 ( .A1(n53), .A2(b[2]), .ZN(n37) );
  AND2_X1 U33bar ( .A1(n53bar), .A2(bbar[2]), .ZN(n37bar) );
  AND2_X1 U34 ( .A1(b[2]), .A2(n53), .ZN(n38) );
  OR2_X1 U34bar ( .A1(bbar[2]), .A2(n53bar), .ZN(n38bar) );
  OR2_X1 U35 ( .A1(n36), .A2(n52), .ZN(y[1]) );
  AND2_X1 U35bar ( .A1(n36bar), .A2(n52bar), .ZN(ybar[1]) );
  OR2_X1 U36 ( .A1(n51), .A2(b[1]), .ZN(n35) );
  AND2_X1 U36bar ( .A1(n51bar), .A2(bbar[1]), .ZN(n35bar) );
  AND2_X1 U37 ( .A1(b[1]), .A2(n51), .ZN(n36) );
  OR2_X1 U37bar ( .A1(bbar[1]), .A2(n51bar), .ZN(n36bar) );
  OR2_X1 U38 ( .A1(n34), .A2(n50), .ZN(y[0]) );
  AND2_X1 U38bar ( .A1(n34bar), .A2(n50bar), .ZN(ybar[0]) );
  OR2_X1 U39 ( .A1(n49), .A2(b[0]), .ZN(n33) );
  AND2_X1 U39bar ( .A1(n49bar), .A2(bbar[0]), .ZN(n33bar) );
  AND2_X1 U40 ( .A1(b[0]), .A2(n49), .ZN(n34) );
  OR2_X1 U40bar ( .A1(bbar[0]), .A2(n49bar), .ZN(n34bar) );
endmodule

module byteXor_12 ( a, b, y );

  input wire [7:0] a;
  input wire [7:0] b;
  wire [7:0] abar;
  wire [7:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
//input_done

  output wire [7:0] y;
  wire [7:0] ybar;
//output_done

  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n33bar;
  wire n34bar;
  wire n35bar;
  wire n36bar;
  wire n37bar;
  wire n38bar;
  wire n39bar;
  wire n40bar;
  wire n41bar;
  wire n42bar;
  wire n43bar;
  wire n44bar;
  wire n45bar;
  wire n46bar;
  wire n47bar;
  wire n48bar;
  wire n49bar;
  wire n50bar;
  wire n51bar;
  wire n52bar;
  wire n53bar;
  wire n54bar;
  wire n55bar;
  wire n56bar;
  wire n57bar;
  wire n58bar;
  wire n59bar;
  wire n60bar;
  wire n61bar;
  wire n62bar;
  wire n63bar;
  wire n64bar;
//wire_done

 //assign_done

  assign n64bar = n47;
  assign n64 = n47bar;
  assign n63bar = a[7];
  assign n63 = abar[7];
  assign n62bar = n45;
  assign n62 = n45bar;
  assign n61bar = a[6];
  assign n61 = abar[6];
  assign n60bar = n43;
  assign n60 = n43bar;
  assign n59bar = a[5];
  assign n59 = abar[5];
  assign n58bar = n41;
  assign n58 = n41bar;
  assign n57bar = a[4];
  assign n57 = abar[4];
  assign n56bar = n39;
  assign n56 = n39bar;
  assign n55bar = a[3];
  assign n55 = abar[3];
  assign n54bar = n37;
  assign n54 = n37bar;
  assign n53bar = a[2];
  assign n53 = abar[2];
  assign n52bar = n35;
  assign n52 = n35bar;
  assign n51bar = a[1];
  assign n51 = abar[1];
  assign n50bar = n33;
  assign n50 = n33bar;
  assign n49bar = a[0];
  assign n49 = abar[0];
  OR2_X1 U17 ( .A1(n48), .A2(n64), .ZN(y[7]) );
  AND2_X1 U17bar ( .A1(n48bar), .A2(n64bar), .ZN(ybar[7]) );
  OR2_X1 U18 ( .A1(n63), .A2(b[7]), .ZN(n47) );
  AND2_X1 U18bar ( .A1(n63bar), .A2(bbar[7]), .ZN(n47bar) );
  AND2_X1 U19 ( .A1(b[7]), .A2(n63), .ZN(n48) );
  OR2_X1 U19bar ( .A1(bbar[7]), .A2(n63bar), .ZN(n48bar) );
  OR2_X1 U20 ( .A1(n46), .A2(n62), .ZN(y[6]) );
  AND2_X1 U20bar ( .A1(n46bar), .A2(n62bar), .ZN(ybar[6]) );
  OR2_X1 U21 ( .A1(n61), .A2(b[6]), .ZN(n45) );
  AND2_X1 U21bar ( .A1(n61bar), .A2(bbar[6]), .ZN(n45bar) );
  AND2_X1 U22 ( .A1(b[6]), .A2(n61), .ZN(n46) );
  OR2_X1 U22bar ( .A1(bbar[6]), .A2(n61bar), .ZN(n46bar) );
  OR2_X1 U23 ( .A1(n44), .A2(n60), .ZN(y[5]) );
  AND2_X1 U23bar ( .A1(n44bar), .A2(n60bar), .ZN(ybar[5]) );
  OR2_X1 U24 ( .A1(n59), .A2(b[5]), .ZN(n43) );
  AND2_X1 U24bar ( .A1(n59bar), .A2(bbar[5]), .ZN(n43bar) );
  AND2_X1 U25 ( .A1(b[5]), .A2(n59), .ZN(n44) );
  OR2_X1 U25bar ( .A1(bbar[5]), .A2(n59bar), .ZN(n44bar) );
  OR2_X1 U26 ( .A1(n42), .A2(n58), .ZN(y[4]) );
  AND2_X1 U26bar ( .A1(n42bar), .A2(n58bar), .ZN(ybar[4]) );
  OR2_X1 U27 ( .A1(n57), .A2(b[4]), .ZN(n41) );
  AND2_X1 U27bar ( .A1(n57bar), .A2(bbar[4]), .ZN(n41bar) );
  AND2_X1 U28 ( .A1(b[4]), .A2(n57), .ZN(n42) );
  OR2_X1 U28bar ( .A1(bbar[4]), .A2(n57bar), .ZN(n42bar) );
  OR2_X1 U29 ( .A1(n40), .A2(n56), .ZN(y[3]) );
  AND2_X1 U29bar ( .A1(n40bar), .A2(n56bar), .ZN(ybar[3]) );
  OR2_X1 U30 ( .A1(n55), .A2(b[3]), .ZN(n39) );
  AND2_X1 U30bar ( .A1(n55bar), .A2(bbar[3]), .ZN(n39bar) );
  AND2_X1 U31 ( .A1(b[3]), .A2(n55), .ZN(n40) );
  OR2_X1 U31bar ( .A1(bbar[3]), .A2(n55bar), .ZN(n40bar) );
  OR2_X1 U32 ( .A1(n38), .A2(n54), .ZN(y[2]) );
  AND2_X1 U32bar ( .A1(n38bar), .A2(n54bar), .ZN(ybar[2]) );
  OR2_X1 U33 ( .A1(n53), .A2(b[2]), .ZN(n37) );
  AND2_X1 U33bar ( .A1(n53bar), .A2(bbar[2]), .ZN(n37bar) );
  AND2_X1 U34 ( .A1(b[2]), .A2(n53), .ZN(n38) );
  OR2_X1 U34bar ( .A1(bbar[2]), .A2(n53bar), .ZN(n38bar) );
  OR2_X1 U35 ( .A1(n36), .A2(n52), .ZN(y[1]) );
  AND2_X1 U35bar ( .A1(n36bar), .A2(n52bar), .ZN(ybar[1]) );
  OR2_X1 U36 ( .A1(n51), .A2(b[1]), .ZN(n35) );
  AND2_X1 U36bar ( .A1(n51bar), .A2(bbar[1]), .ZN(n35bar) );
  AND2_X1 U37 ( .A1(b[1]), .A2(n51), .ZN(n36) );
  OR2_X1 U37bar ( .A1(bbar[1]), .A2(n51bar), .ZN(n36bar) );
  OR2_X1 U38 ( .A1(n34), .A2(n50), .ZN(y[0]) );
  AND2_X1 U38bar ( .A1(n34bar), .A2(n50bar), .ZN(ybar[0]) );
  OR2_X1 U39 ( .A1(n49), .A2(b[0]), .ZN(n33) );
  AND2_X1 U39bar ( .A1(n49bar), .A2(bbar[0]), .ZN(n33bar) );
  AND2_X1 U40 ( .A1(b[0]), .A2(n49), .ZN(n34) );
  OR2_X1 U40bar ( .A1(bbar[0]), .A2(n49bar), .ZN(n34bar) );
endmodule

module byteXor_13 ( a, b, y );

  input wire [7:0] a;
  input wire [7:0] b;
  wire [7:0] abar;
  wire [7:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
//input_done

  output wire [7:0] y;
  wire [7:0] ybar;
//output_done

  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n33bar;
  wire n34bar;
  wire n35bar;
  wire n36bar;
  wire n37bar;
  wire n38bar;
  wire n39bar;
  wire n40bar;
  wire n41bar;
  wire n42bar;
  wire n43bar;
  wire n44bar;
  wire n45bar;
  wire n46bar;
  wire n47bar;
  wire n48bar;
  wire n49bar;
  wire n50bar;
  wire n51bar;
  wire n52bar;
  wire n53bar;
  wire n54bar;
  wire n55bar;
  wire n56bar;
  wire n57bar;
  wire n58bar;
  wire n59bar;
  wire n60bar;
  wire n61bar;
  wire n62bar;
  wire n63bar;
  wire n64bar;
//wire_done

 //assign_done

  assign n64bar = n47;
  assign n64 = n47bar;
  assign n63bar = a[7];
  assign n63 = abar[7];
  assign n62bar = n45;
  assign n62 = n45bar;
  assign n61bar = a[6];
  assign n61 = abar[6];
  assign n60bar = n43;
  assign n60 = n43bar;
  assign n59bar = a[5];
  assign n59 = abar[5];
  assign n58bar = n41;
  assign n58 = n41bar;
  assign n57bar = a[4];
  assign n57 = abar[4];
  assign n56bar = n39;
  assign n56 = n39bar;
  assign n55bar = a[3];
  assign n55 = abar[3];
  assign n54bar = n37;
  assign n54 = n37bar;
  assign n53bar = a[2];
  assign n53 = abar[2];
  assign n52bar = n35;
  assign n52 = n35bar;
  assign n51bar = a[1];
  assign n51 = abar[1];
  assign n50bar = n33;
  assign n50 = n33bar;
  assign n49bar = a[0];
  assign n49 = abar[0];
  OR2_X1 U17 ( .A1(n48), .A2(n64), .ZN(y[7]) );
  AND2_X1 U17bar ( .A1(n48bar), .A2(n64bar), .ZN(ybar[7]) );
  OR2_X1 U18 ( .A1(n63), .A2(b[7]), .ZN(n47) );
  AND2_X1 U18bar ( .A1(n63bar), .A2(bbar[7]), .ZN(n47bar) );
  AND2_X1 U19 ( .A1(b[7]), .A2(n63), .ZN(n48) );
  OR2_X1 U19bar ( .A1(bbar[7]), .A2(n63bar), .ZN(n48bar) );
  OR2_X1 U20 ( .A1(n46), .A2(n62), .ZN(y[6]) );
  AND2_X1 U20bar ( .A1(n46bar), .A2(n62bar), .ZN(ybar[6]) );
  OR2_X1 U21 ( .A1(n61), .A2(b[6]), .ZN(n45) );
  AND2_X1 U21bar ( .A1(n61bar), .A2(bbar[6]), .ZN(n45bar) );
  AND2_X1 U22 ( .A1(b[6]), .A2(n61), .ZN(n46) );
  OR2_X1 U22bar ( .A1(bbar[6]), .A2(n61bar), .ZN(n46bar) );
  OR2_X1 U23 ( .A1(n44), .A2(n60), .ZN(y[5]) );
  AND2_X1 U23bar ( .A1(n44bar), .A2(n60bar), .ZN(ybar[5]) );
  OR2_X1 U24 ( .A1(n59), .A2(b[5]), .ZN(n43) );
  AND2_X1 U24bar ( .A1(n59bar), .A2(bbar[5]), .ZN(n43bar) );
  AND2_X1 U25 ( .A1(b[5]), .A2(n59), .ZN(n44) );
  OR2_X1 U25bar ( .A1(bbar[5]), .A2(n59bar), .ZN(n44bar) );
  OR2_X1 U26 ( .A1(n42), .A2(n58), .ZN(y[4]) );
  AND2_X1 U26bar ( .A1(n42bar), .A2(n58bar), .ZN(ybar[4]) );
  OR2_X1 U27 ( .A1(n57), .A2(b[4]), .ZN(n41) );
  AND2_X1 U27bar ( .A1(n57bar), .A2(bbar[4]), .ZN(n41bar) );
  AND2_X1 U28 ( .A1(b[4]), .A2(n57), .ZN(n42) );
  OR2_X1 U28bar ( .A1(bbar[4]), .A2(n57bar), .ZN(n42bar) );
  OR2_X1 U29 ( .A1(n40), .A2(n56), .ZN(y[3]) );
  AND2_X1 U29bar ( .A1(n40bar), .A2(n56bar), .ZN(ybar[3]) );
  OR2_X1 U30 ( .A1(n55), .A2(b[3]), .ZN(n39) );
  AND2_X1 U30bar ( .A1(n55bar), .A2(bbar[3]), .ZN(n39bar) );
  AND2_X1 U31 ( .A1(b[3]), .A2(n55), .ZN(n40) );
  OR2_X1 U31bar ( .A1(bbar[3]), .A2(n55bar), .ZN(n40bar) );
  OR2_X1 U32 ( .A1(n38), .A2(n54), .ZN(y[2]) );
  AND2_X1 U32bar ( .A1(n38bar), .A2(n54bar), .ZN(ybar[2]) );
  OR2_X1 U33 ( .A1(n53), .A2(b[2]), .ZN(n37) );
  AND2_X1 U33bar ( .A1(n53bar), .A2(bbar[2]), .ZN(n37bar) );
  AND2_X1 U34 ( .A1(b[2]), .A2(n53), .ZN(n38) );
  OR2_X1 U34bar ( .A1(bbar[2]), .A2(n53bar), .ZN(n38bar) );
  OR2_X1 U35 ( .A1(n36), .A2(n52), .ZN(y[1]) );
  AND2_X1 U35bar ( .A1(n36bar), .A2(n52bar), .ZN(ybar[1]) );
  OR2_X1 U36 ( .A1(n51), .A2(b[1]), .ZN(n35) );
  AND2_X1 U36bar ( .A1(n51bar), .A2(bbar[1]), .ZN(n35bar) );
  AND2_X1 U37 ( .A1(b[1]), .A2(n51), .ZN(n36) );
  OR2_X1 U37bar ( .A1(bbar[1]), .A2(n51bar), .ZN(n36bar) );
  OR2_X1 U38 ( .A1(n34), .A2(n50), .ZN(y[0]) );
  AND2_X1 U38bar ( .A1(n34bar), .A2(n50bar), .ZN(ybar[0]) );
  OR2_X1 U39 ( .A1(n49), .A2(b[0]), .ZN(n33) );
  AND2_X1 U39bar ( .A1(n49bar), .A2(bbar[0]), .ZN(n33bar) );
  AND2_X1 U40 ( .A1(b[0]), .A2(n49), .ZN(n34) );
  OR2_X1 U40bar ( .A1(bbar[0]), .A2(n49bar), .ZN(n34bar) );
endmodule

module byteXor4_9 ( a, b, c, d, y );

  input wire [7:0] a;
  input wire [7:0] b;
  input wire [7:0] c;
  input wire [7:0] d;
  wire [7:0] abar;
  wire [7:0] bbar;
  wire [7:0] cbar;
  wire [7:0] dbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign cbar[0] = ~c[0];
  assign cbar[1] = ~c[1];
  assign cbar[2] = ~c[2];
  assign cbar[3] = ~c[3];
  assign cbar[4] = ~c[4];
  assign cbar[5] = ~c[5];
  assign cbar[6] = ~c[6];
  assign cbar[7] = ~c[7];
  assign dbar[0] = ~d[0];
  assign dbar[1] = ~d[1];
  assign dbar[2] = ~d[2];
  assign dbar[3] = ~d[3];
  assign dbar[4] = ~d[4];
  assign dbar[5] = ~d[5];
  assign dbar[6] = ~d[6];
  assign dbar[7] = ~d[7];
//input_done

  output wire [7:0] y;
  wire [7:0] ybar;
//output_done

  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n113bar;
  wire n114bar;
  wire n115bar;
  wire n116bar;
  wire n117bar;
  wire n118bar;
  wire n119bar;
  wire n120bar;
  wire n121bar;
  wire n122bar;
  wire n123bar;
  wire n124bar;
  wire n125bar;
  wire n126bar;
  wire n127bar;
  wire n128bar;
  wire n129bar;
  wire n130bar;
  wire n131bar;
  wire n132bar;
  wire n133bar;
  wire n134bar;
  wire n135bar;
  wire n136bar;
  wire n137bar;
  wire n138bar;
  wire n139bar;
  wire n140bar;
  wire n141bar;
  wire n142bar;
  wire n143bar;
  wire n144bar;
  wire n145bar;
  wire n146bar;
  wire n147bar;
  wire n148bar;
  wire n149bar;
  wire n150bar;
  wire n151bar;
  wire n152bar;
  wire n153bar;
  wire n154bar;
  wire n155bar;
  wire n156bar;
  wire n157bar;
  wire n158bar;
  wire n159bar;
  wire n160bar;
  wire n161bar;
  wire n162bar;
  wire n163bar;
  wire n164bar;
  wire n165bar;
  wire n166bar;
  wire n167bar;
  wire n168bar;
  wire n169bar;
  wire n170bar;
  wire n171bar;
  wire n172bar;
  wire n173bar;
  wire n174bar;
  wire n175bar;
  wire n176bar;
  wire n177bar;
  wire n178bar;
  wire n179bar;
  wire n180bar;
  wire n181bar;
  wire n182bar;
  wire n183bar;
  wire n184bar;
  wire n185bar;
  wire n186bar;
  wire n187bar;
  wire n188bar;
  wire n189bar;
  wire n190bar;
  wire n191bar;
  wire n192bar;
  wire n193bar;
  wire n194bar;
  wire n195bar;
  wire n196bar;
  wire n197bar;
  wire n198bar;
  wire n199bar;
  wire n200bar;
  wire n201bar;
  wire n202bar;
  wire n203bar;
  wire n204bar;
  wire n205bar;
  wire n206bar;
  wire n207bar;
  wire n208bar;
  wire n209bar;
  wire n210bar;
  wire n211bar;
  wire n212bar;
  wire n213bar;
  wire n214bar;
  wire n215bar;
  wire n216bar;
  wire n217bar;
  wire n218bar;
  wire n219bar;
  wire n220bar;
  wire n221bar;
  wire n222bar;
  wire n223bar;
  wire n224bar;
//wire_done

 //assign_done

  assign n224bar = n175;
  assign n224 = n175bar;
  assign n223bar = a[7];
  assign n223 = abar[7];
  assign n222bar = n167;
  assign n222 = n167bar;
  assign n221bar = a[6];
  assign n221 = abar[6];
  assign n220bar = n159;
  assign n220 = n159bar;
  assign n219bar = a[5];
  assign n219 = abar[5];
  assign n218bar = n151;
  assign n218 = n151bar;
  assign n217bar = a[4];
  assign n217 = abar[4];
  assign n216bar = n143;
  assign n216 = n143bar;
  assign n215bar = a[3];
  assign n215 = abar[3];
  assign n214bar = n135;
  assign n214 = n135bar;
  assign n213bar = a[2];
  assign n213 = abar[2];
  assign n212bar = n127;
  assign n212 = n127bar;
  assign n211bar = a[1];
  assign n211 = abar[1];
  assign n210bar = n119;
  assign n210 = n119bar;
  assign n209bar = a[0];
  assign n209 = abar[0];
  assign n208bar = b[7];
  assign n208 = bbar[7];
  assign n207bar = b[6];
  assign n207 = bbar[6];
  assign n206bar = b[5];
  assign n206 = bbar[5];
  assign n205bar = b[4];
  assign n205 = bbar[4];
  assign n204bar = b[3];
  assign n204 = bbar[3];
  assign n203bar = b[2];
  assign n203 = bbar[2];
  assign n202bar = b[1];
  assign n202 = bbar[1];
  assign n201bar = b[0];
  assign n201 = bbar[0];
  assign n200bar = n171;
  assign n200 = n171bar;
  assign n199bar = c[7];
  assign n199 = cbar[7];
  assign n198bar = n163;
  assign n198 = n163bar;
  assign n197bar = c[6];
  assign n197 = cbar[6];
  assign n196bar = n155;
  assign n196 = n155bar;
  assign n195bar = c[5];
  assign n195 = cbar[5];
  assign n194bar = n147;
  assign n194 = n147bar;
  assign n193bar = c[4];
  assign n193 = cbar[4];
  assign n192bar = n139;
  assign n192 = n139bar;
  assign n191bar = c[3];
  assign n191 = cbar[3];
  assign n190bar = n131;
  assign n190 = n131bar;
  assign n189bar = c[2];
  assign n189 = cbar[2];
  assign n188bar = n123;
  assign n188 = n123bar;
  assign n187bar = c[1];
  assign n187 = cbar[1];
  assign n186bar = n115;
  assign n186 = n115bar;
  assign n185bar = c[0];
  assign n185 = cbar[0];
  assign n184bar = d[7];
  assign n184 = dbar[7];
  assign n183bar = d[6];
  assign n183 = dbar[6];
  assign n182bar = d[5];
  assign n182 = dbar[5];
  assign n181bar = d[4];
  assign n181 = dbar[4];
  assign n180bar = d[3];
  assign n180 = dbar[3];
  assign n179bar = d[2];
  assign n179 = dbar[2];
  assign n178bar = d[1];
  assign n178 = dbar[1];
  assign n177bar = d[0];
  assign n177 = dbar[0];
  OR2_X1 U49 ( .A1(n176), .A2(n224), .ZN(y[7]) );
  AND2_X1 U49bar ( .A1(n176bar), .A2(n224bar), .ZN(ybar[7]) );
  OR2_X1 U50 ( .A1(n174), .A2(n200), .ZN(n175) );
  AND2_X1 U50bar ( .A1(n174bar), .A2(n200bar), .ZN(n175bar) );
  AND2_X1 U51 ( .A1(n200), .A2(n174), .ZN(n176) );
  OR2_X1 U51bar ( .A1(n200bar), .A2(n174bar), .ZN(n176bar) );
  AND2_X1 U52 ( .A1(n173), .A2(n172), .ZN(n174) );
  OR2_X1 U52bar ( .A1(n173bar), .A2(n172bar), .ZN(n174bar) );
  OR2_X1 U53 ( .A1(n223), .A2(b[7]), .ZN(n172) );
  AND2_X1 U53bar ( .A1(n223bar), .A2(bbar[7]), .ZN(n172bar) );
  OR2_X1 U54 ( .A1(n208), .A2(a[7]), .ZN(n173) );
  AND2_X1 U54bar ( .A1(n208bar), .A2(abar[7]), .ZN(n173bar) );
  AND2_X1 U55 ( .A1(n170), .A2(n169), .ZN(n171) );
  OR2_X1 U55bar ( .A1(n170bar), .A2(n169bar), .ZN(n171bar) );
  OR2_X1 U56 ( .A1(n199), .A2(d[7]), .ZN(n169) );
  AND2_X1 U56bar ( .A1(n199bar), .A2(dbar[7]), .ZN(n169bar) );
  OR2_X1 U57 ( .A1(n184), .A2(c[7]), .ZN(n170) );
  AND2_X1 U57bar ( .A1(n184bar), .A2(cbar[7]), .ZN(n170bar) );
  OR2_X1 U58 ( .A1(n168), .A2(n222), .ZN(y[6]) );
  AND2_X1 U58bar ( .A1(n168bar), .A2(n222bar), .ZN(ybar[6]) );
  OR2_X1 U59 ( .A1(n166), .A2(n198), .ZN(n167) );
  AND2_X1 U59bar ( .A1(n166bar), .A2(n198bar), .ZN(n167bar) );
  AND2_X1 U60 ( .A1(n198), .A2(n166), .ZN(n168) );
  OR2_X1 U60bar ( .A1(n198bar), .A2(n166bar), .ZN(n168bar) );
  AND2_X1 U61 ( .A1(n165), .A2(n164), .ZN(n166) );
  OR2_X1 U61bar ( .A1(n165bar), .A2(n164bar), .ZN(n166bar) );
  OR2_X1 U62 ( .A1(n221), .A2(b[6]), .ZN(n164) );
  AND2_X1 U62bar ( .A1(n221bar), .A2(bbar[6]), .ZN(n164bar) );
  OR2_X1 U63 ( .A1(n207), .A2(a[6]), .ZN(n165) );
  AND2_X1 U63bar ( .A1(n207bar), .A2(abar[6]), .ZN(n165bar) );
  AND2_X1 U64 ( .A1(n162), .A2(n161), .ZN(n163) );
  OR2_X1 U64bar ( .A1(n162bar), .A2(n161bar), .ZN(n163bar) );
  OR2_X1 U65 ( .A1(n197), .A2(d[6]), .ZN(n161) );
  AND2_X1 U65bar ( .A1(n197bar), .A2(dbar[6]), .ZN(n161bar) );
  OR2_X1 U66 ( .A1(n183), .A2(c[6]), .ZN(n162) );
  AND2_X1 U66bar ( .A1(n183bar), .A2(cbar[6]), .ZN(n162bar) );
  OR2_X1 U67 ( .A1(n160), .A2(n220), .ZN(y[5]) );
  AND2_X1 U67bar ( .A1(n160bar), .A2(n220bar), .ZN(ybar[5]) );
  OR2_X1 U68 ( .A1(n158), .A2(n196), .ZN(n159) );
  AND2_X1 U68bar ( .A1(n158bar), .A2(n196bar), .ZN(n159bar) );
  AND2_X1 U69 ( .A1(n196), .A2(n158), .ZN(n160) );
  OR2_X1 U69bar ( .A1(n196bar), .A2(n158bar), .ZN(n160bar) );
  AND2_X1 U70 ( .A1(n157), .A2(n156), .ZN(n158) );
  OR2_X1 U70bar ( .A1(n157bar), .A2(n156bar), .ZN(n158bar) );
  OR2_X1 U71 ( .A1(n219), .A2(b[5]), .ZN(n156) );
  AND2_X1 U71bar ( .A1(n219bar), .A2(bbar[5]), .ZN(n156bar) );
  OR2_X1 U72 ( .A1(n206), .A2(a[5]), .ZN(n157) );
  AND2_X1 U72bar ( .A1(n206bar), .A2(abar[5]), .ZN(n157bar) );
  AND2_X1 U73 ( .A1(n154), .A2(n153), .ZN(n155) );
  OR2_X1 U73bar ( .A1(n154bar), .A2(n153bar), .ZN(n155bar) );
  OR2_X1 U74 ( .A1(n195), .A2(d[5]), .ZN(n153) );
  AND2_X1 U74bar ( .A1(n195bar), .A2(dbar[5]), .ZN(n153bar) );
  OR2_X1 U75 ( .A1(n182), .A2(c[5]), .ZN(n154) );
  AND2_X1 U75bar ( .A1(n182bar), .A2(cbar[5]), .ZN(n154bar) );
  OR2_X1 U76 ( .A1(n152), .A2(n218), .ZN(y[4]) );
  AND2_X1 U76bar ( .A1(n152bar), .A2(n218bar), .ZN(ybar[4]) );
  OR2_X1 U77 ( .A1(n150), .A2(n194), .ZN(n151) );
  AND2_X1 U77bar ( .A1(n150bar), .A2(n194bar), .ZN(n151bar) );
  AND2_X1 U78 ( .A1(n194), .A2(n150), .ZN(n152) );
  OR2_X1 U78bar ( .A1(n194bar), .A2(n150bar), .ZN(n152bar) );
  AND2_X1 U79 ( .A1(n149), .A2(n148), .ZN(n150) );
  OR2_X1 U79bar ( .A1(n149bar), .A2(n148bar), .ZN(n150bar) );
  OR2_X1 U80 ( .A1(n217), .A2(b[4]), .ZN(n148) );
  AND2_X1 U80bar ( .A1(n217bar), .A2(bbar[4]), .ZN(n148bar) );
  OR2_X1 U81 ( .A1(n205), .A2(a[4]), .ZN(n149) );
  AND2_X1 U81bar ( .A1(n205bar), .A2(abar[4]), .ZN(n149bar) );
  AND2_X1 U82 ( .A1(n146), .A2(n145), .ZN(n147) );
  OR2_X1 U82bar ( .A1(n146bar), .A2(n145bar), .ZN(n147bar) );
  OR2_X1 U83 ( .A1(n193), .A2(d[4]), .ZN(n145) );
  AND2_X1 U83bar ( .A1(n193bar), .A2(dbar[4]), .ZN(n145bar) );
  OR2_X1 U84 ( .A1(n181), .A2(c[4]), .ZN(n146) );
  AND2_X1 U84bar ( .A1(n181bar), .A2(cbar[4]), .ZN(n146bar) );
  OR2_X1 U85 ( .A1(n144), .A2(n216), .ZN(y[3]) );
  AND2_X1 U85bar ( .A1(n144bar), .A2(n216bar), .ZN(ybar[3]) );
  OR2_X1 U86 ( .A1(n142), .A2(n192), .ZN(n143) );
  AND2_X1 U86bar ( .A1(n142bar), .A2(n192bar), .ZN(n143bar) );
  AND2_X1 U87 ( .A1(n192), .A2(n142), .ZN(n144) );
  OR2_X1 U87bar ( .A1(n192bar), .A2(n142bar), .ZN(n144bar) );
  AND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(n142) );
  OR2_X1 U88bar ( .A1(n141bar), .A2(n140bar), .ZN(n142bar) );
  OR2_X1 U89 ( .A1(n215), .A2(b[3]), .ZN(n140) );
  AND2_X1 U89bar ( .A1(n215bar), .A2(bbar[3]), .ZN(n140bar) );
  OR2_X1 U90 ( .A1(n204), .A2(a[3]), .ZN(n141) );
  AND2_X1 U90bar ( .A1(n204bar), .A2(abar[3]), .ZN(n141bar) );
  AND2_X1 U91 ( .A1(n138), .A2(n137), .ZN(n139) );
  OR2_X1 U91bar ( .A1(n138bar), .A2(n137bar), .ZN(n139bar) );
  OR2_X1 U92 ( .A1(n191), .A2(d[3]), .ZN(n137) );
  AND2_X1 U92bar ( .A1(n191bar), .A2(dbar[3]), .ZN(n137bar) );
  OR2_X1 U93 ( .A1(n180), .A2(c[3]), .ZN(n138) );
  AND2_X1 U93bar ( .A1(n180bar), .A2(cbar[3]), .ZN(n138bar) );
  OR2_X1 U94 ( .A1(n136), .A2(n214), .ZN(y[2]) );
  AND2_X1 U94bar ( .A1(n136bar), .A2(n214bar), .ZN(ybar[2]) );
  OR2_X1 U95 ( .A1(n134), .A2(n190), .ZN(n135) );
  AND2_X1 U95bar ( .A1(n134bar), .A2(n190bar), .ZN(n135bar) );
  AND2_X1 U96 ( .A1(n190), .A2(n134), .ZN(n136) );
  OR2_X1 U96bar ( .A1(n190bar), .A2(n134bar), .ZN(n136bar) );
  AND2_X1 U97 ( .A1(n133), .A2(n132), .ZN(n134) );
  OR2_X1 U97bar ( .A1(n133bar), .A2(n132bar), .ZN(n134bar) );
  OR2_X1 U98 ( .A1(n213), .A2(b[2]), .ZN(n132) );
  AND2_X1 U98bar ( .A1(n213bar), .A2(bbar[2]), .ZN(n132bar) );
  OR2_X1 U99 ( .A1(n203), .A2(a[2]), .ZN(n133) );
  AND2_X1 U99bar ( .A1(n203bar), .A2(abar[2]), .ZN(n133bar) );
  AND2_X1 U100 ( .A1(n130), .A2(n129), .ZN(n131) );
  OR2_X1 U100bar ( .A1(n130bar), .A2(n129bar), .ZN(n131bar) );
  OR2_X1 U101 ( .A1(n189), .A2(d[2]), .ZN(n129) );
  AND2_X1 U101bar ( .A1(n189bar), .A2(dbar[2]), .ZN(n129bar) );
  OR2_X1 U102 ( .A1(n179), .A2(c[2]), .ZN(n130) );
  AND2_X1 U102bar ( .A1(n179bar), .A2(cbar[2]), .ZN(n130bar) );
  OR2_X1 U103 ( .A1(n128), .A2(n212), .ZN(y[1]) );
  AND2_X1 U103bar ( .A1(n128bar), .A2(n212bar), .ZN(ybar[1]) );
  OR2_X1 U104 ( .A1(n126), .A2(n188), .ZN(n127) );
  AND2_X1 U104bar ( .A1(n126bar), .A2(n188bar), .ZN(n127bar) );
  AND2_X1 U105 ( .A1(n188), .A2(n126), .ZN(n128) );
  OR2_X1 U105bar ( .A1(n188bar), .A2(n126bar), .ZN(n128bar) );
  AND2_X1 U106 ( .A1(n125), .A2(n124), .ZN(n126) );
  OR2_X1 U106bar ( .A1(n125bar), .A2(n124bar), .ZN(n126bar) );
  OR2_X1 U107 ( .A1(n211), .A2(b[1]), .ZN(n124) );
  AND2_X1 U107bar ( .A1(n211bar), .A2(bbar[1]), .ZN(n124bar) );
  OR2_X1 U108 ( .A1(n202), .A2(a[1]), .ZN(n125) );
  AND2_X1 U108bar ( .A1(n202bar), .A2(abar[1]), .ZN(n125bar) );
  AND2_X1 U109 ( .A1(n122), .A2(n121), .ZN(n123) );
  OR2_X1 U109bar ( .A1(n122bar), .A2(n121bar), .ZN(n123bar) );
  OR2_X1 U110 ( .A1(n187), .A2(d[1]), .ZN(n121) );
  AND2_X1 U110bar ( .A1(n187bar), .A2(dbar[1]), .ZN(n121bar) );
  OR2_X1 U111 ( .A1(n178), .A2(c[1]), .ZN(n122) );
  AND2_X1 U111bar ( .A1(n178bar), .A2(cbar[1]), .ZN(n122bar) );
  OR2_X1 U112 ( .A1(n120), .A2(n210), .ZN(y[0]) );
  AND2_X1 U112bar ( .A1(n120bar), .A2(n210bar), .ZN(ybar[0]) );
  OR2_X1 U113 ( .A1(n118), .A2(n186), .ZN(n119) );
  AND2_X1 U113bar ( .A1(n118bar), .A2(n186bar), .ZN(n119bar) );
  AND2_X1 U114 ( .A1(n186), .A2(n118), .ZN(n120) );
  OR2_X1 U114bar ( .A1(n186bar), .A2(n118bar), .ZN(n120bar) );
  AND2_X1 U115 ( .A1(n117), .A2(n116), .ZN(n118) );
  OR2_X1 U115bar ( .A1(n117bar), .A2(n116bar), .ZN(n118bar) );
  OR2_X1 U116 ( .A1(n209), .A2(b[0]), .ZN(n116) );
  AND2_X1 U116bar ( .A1(n209bar), .A2(bbar[0]), .ZN(n116bar) );
  OR2_X1 U117 ( .A1(n201), .A2(a[0]), .ZN(n117) );
  AND2_X1 U117bar ( .A1(n201bar), .A2(abar[0]), .ZN(n117bar) );
  AND2_X1 U118 ( .A1(n114), .A2(n113), .ZN(n115) );
  OR2_X1 U118bar ( .A1(n114bar), .A2(n113bar), .ZN(n115bar) );
  OR2_X1 U119 ( .A1(n185), .A2(d[0]), .ZN(n113) );
  AND2_X1 U119bar ( .A1(n185bar), .A2(dbar[0]), .ZN(n113bar) );
  OR2_X1 U120 ( .A1(n177), .A2(c[0]), .ZN(n114) );
  AND2_X1 U120bar ( .A1(n177bar), .A2(cbar[0]), .ZN(n114bar) );
endmodule

module byteXor4_10 ( a, b, c, d, y );

  input wire [7:0] a;
  input wire [7:0] b;
  input wire [7:0] c;
  input wire [7:0] d;
  wire [7:0] abar;
  wire [7:0] bbar;
  wire [7:0] cbar;
  wire [7:0] dbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign cbar[0] = ~c[0];
  assign cbar[1] = ~c[1];
  assign cbar[2] = ~c[2];
  assign cbar[3] = ~c[3];
  assign cbar[4] = ~c[4];
  assign cbar[5] = ~c[5];
  assign cbar[6] = ~c[6];
  assign cbar[7] = ~c[7];
  assign dbar[0] = ~d[0];
  assign dbar[1] = ~d[1];
  assign dbar[2] = ~d[2];
  assign dbar[3] = ~d[3];
  assign dbar[4] = ~d[4];
  assign dbar[5] = ~d[5];
  assign dbar[6] = ~d[6];
  assign dbar[7] = ~d[7];
//input_done

  output wire [7:0] y;
  wire [7:0] ybar;
//output_done

  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n113bar;
  wire n114bar;
  wire n115bar;
  wire n116bar;
  wire n117bar;
  wire n118bar;
  wire n119bar;
  wire n120bar;
  wire n121bar;
  wire n122bar;
  wire n123bar;
  wire n124bar;
  wire n125bar;
  wire n126bar;
  wire n127bar;
  wire n128bar;
  wire n129bar;
  wire n130bar;
  wire n131bar;
  wire n132bar;
  wire n133bar;
  wire n134bar;
  wire n135bar;
  wire n136bar;
  wire n137bar;
  wire n138bar;
  wire n139bar;
  wire n140bar;
  wire n141bar;
  wire n142bar;
  wire n143bar;
  wire n144bar;
  wire n145bar;
  wire n146bar;
  wire n147bar;
  wire n148bar;
  wire n149bar;
  wire n150bar;
  wire n151bar;
  wire n152bar;
  wire n153bar;
  wire n154bar;
  wire n155bar;
  wire n156bar;
  wire n157bar;
  wire n158bar;
  wire n159bar;
  wire n160bar;
  wire n161bar;
  wire n162bar;
  wire n163bar;
  wire n164bar;
  wire n165bar;
  wire n166bar;
  wire n167bar;
  wire n168bar;
  wire n169bar;
  wire n170bar;
  wire n171bar;
  wire n172bar;
  wire n173bar;
  wire n174bar;
  wire n175bar;
  wire n176bar;
  wire n177bar;
  wire n178bar;
  wire n179bar;
  wire n180bar;
  wire n181bar;
  wire n182bar;
  wire n183bar;
  wire n184bar;
  wire n185bar;
  wire n186bar;
  wire n187bar;
  wire n188bar;
  wire n189bar;
  wire n190bar;
  wire n191bar;
  wire n192bar;
  wire n193bar;
  wire n194bar;
  wire n195bar;
  wire n196bar;
  wire n197bar;
  wire n198bar;
  wire n199bar;
  wire n200bar;
  wire n201bar;
  wire n202bar;
  wire n203bar;
  wire n204bar;
  wire n205bar;
  wire n206bar;
  wire n207bar;
  wire n208bar;
  wire n209bar;
  wire n210bar;
  wire n211bar;
  wire n212bar;
  wire n213bar;
  wire n214bar;
  wire n215bar;
  wire n216bar;
  wire n217bar;
  wire n218bar;
  wire n219bar;
  wire n220bar;
  wire n221bar;
  wire n222bar;
  wire n223bar;
  wire n224bar;
//wire_done

 //assign_done

  assign n224bar = n175;
  assign n224 = n175bar;
  assign n223bar = a[7];
  assign n223 = abar[7];
  assign n222bar = n167;
  assign n222 = n167bar;
  assign n221bar = a[6];
  assign n221 = abar[6];
  assign n220bar = n159;
  assign n220 = n159bar;
  assign n219bar = a[5];
  assign n219 = abar[5];
  assign n218bar = n151;
  assign n218 = n151bar;
  assign n217bar = a[4];
  assign n217 = abar[4];
  assign n216bar = n143;
  assign n216 = n143bar;
  assign n215bar = a[3];
  assign n215 = abar[3];
  assign n214bar = n135;
  assign n214 = n135bar;
  assign n213bar = a[2];
  assign n213 = abar[2];
  assign n212bar = n127;
  assign n212 = n127bar;
  assign n211bar = a[1];
  assign n211 = abar[1];
  assign n210bar = n119;
  assign n210 = n119bar;
  assign n209bar = a[0];
  assign n209 = abar[0];
  assign n208bar = b[7];
  assign n208 = bbar[7];
  assign n207bar = b[6];
  assign n207 = bbar[6];
  assign n206bar = b[5];
  assign n206 = bbar[5];
  assign n205bar = b[4];
  assign n205 = bbar[4];
  assign n204bar = b[3];
  assign n204 = bbar[3];
  assign n203bar = b[2];
  assign n203 = bbar[2];
  assign n202bar = b[1];
  assign n202 = bbar[1];
  assign n201bar = b[0];
  assign n201 = bbar[0];
  assign n200bar = n171;
  assign n200 = n171bar;
  assign n199bar = c[7];
  assign n199 = cbar[7];
  assign n198bar = n163;
  assign n198 = n163bar;
  assign n197bar = c[6];
  assign n197 = cbar[6];
  assign n196bar = n155;
  assign n196 = n155bar;
  assign n195bar = c[5];
  assign n195 = cbar[5];
  assign n194bar = n147;
  assign n194 = n147bar;
  assign n193bar = c[4];
  assign n193 = cbar[4];
  assign n192bar = n139;
  assign n192 = n139bar;
  assign n191bar = c[3];
  assign n191 = cbar[3];
  assign n190bar = n131;
  assign n190 = n131bar;
  assign n189bar = c[2];
  assign n189 = cbar[2];
  assign n188bar = n123;
  assign n188 = n123bar;
  assign n187bar = c[1];
  assign n187 = cbar[1];
  assign n186bar = n115;
  assign n186 = n115bar;
  assign n185bar = c[0];
  assign n185 = cbar[0];
  assign n184bar = d[7];
  assign n184 = dbar[7];
  assign n183bar = d[6];
  assign n183 = dbar[6];
  assign n182bar = d[5];
  assign n182 = dbar[5];
  assign n181bar = d[4];
  assign n181 = dbar[4];
  assign n180bar = d[3];
  assign n180 = dbar[3];
  assign n179bar = d[2];
  assign n179 = dbar[2];
  assign n178bar = d[1];
  assign n178 = dbar[1];
  assign n177bar = d[0];
  assign n177 = dbar[0];
  OR2_X1 U49 ( .A1(n176), .A2(n224), .ZN(y[7]) );
  AND2_X1 U49bar ( .A1(n176bar), .A2(n224bar), .ZN(ybar[7]) );
  OR2_X1 U50 ( .A1(n174), .A2(n200), .ZN(n175) );
  AND2_X1 U50bar ( .A1(n174bar), .A2(n200bar), .ZN(n175bar) );
  AND2_X1 U51 ( .A1(n200), .A2(n174), .ZN(n176) );
  OR2_X1 U51bar ( .A1(n200bar), .A2(n174bar), .ZN(n176bar) );
  AND2_X1 U52 ( .A1(n173), .A2(n172), .ZN(n174) );
  OR2_X1 U52bar ( .A1(n173bar), .A2(n172bar), .ZN(n174bar) );
  OR2_X1 U53 ( .A1(n223), .A2(b[7]), .ZN(n172) );
  AND2_X1 U53bar ( .A1(n223bar), .A2(bbar[7]), .ZN(n172bar) );
  OR2_X1 U54 ( .A1(n208), .A2(a[7]), .ZN(n173) );
  AND2_X1 U54bar ( .A1(n208bar), .A2(abar[7]), .ZN(n173bar) );
  AND2_X1 U55 ( .A1(n170), .A2(n169), .ZN(n171) );
  OR2_X1 U55bar ( .A1(n170bar), .A2(n169bar), .ZN(n171bar) );
  OR2_X1 U56 ( .A1(n199), .A2(d[7]), .ZN(n169) );
  AND2_X1 U56bar ( .A1(n199bar), .A2(dbar[7]), .ZN(n169bar) );
  OR2_X1 U57 ( .A1(n184), .A2(c[7]), .ZN(n170) );
  AND2_X1 U57bar ( .A1(n184bar), .A2(cbar[7]), .ZN(n170bar) );
  OR2_X1 U58 ( .A1(n168), .A2(n222), .ZN(y[6]) );
  AND2_X1 U58bar ( .A1(n168bar), .A2(n222bar), .ZN(ybar[6]) );
  OR2_X1 U59 ( .A1(n166), .A2(n198), .ZN(n167) );
  AND2_X1 U59bar ( .A1(n166bar), .A2(n198bar), .ZN(n167bar) );
  AND2_X1 U60 ( .A1(n198), .A2(n166), .ZN(n168) );
  OR2_X1 U60bar ( .A1(n198bar), .A2(n166bar), .ZN(n168bar) );
  AND2_X1 U61 ( .A1(n165), .A2(n164), .ZN(n166) );
  OR2_X1 U61bar ( .A1(n165bar), .A2(n164bar), .ZN(n166bar) );
  OR2_X1 U62 ( .A1(n221), .A2(b[6]), .ZN(n164) );
  AND2_X1 U62bar ( .A1(n221bar), .A2(bbar[6]), .ZN(n164bar) );
  OR2_X1 U63 ( .A1(n207), .A2(a[6]), .ZN(n165) );
  AND2_X1 U63bar ( .A1(n207bar), .A2(abar[6]), .ZN(n165bar) );
  AND2_X1 U64 ( .A1(n162), .A2(n161), .ZN(n163) );
  OR2_X1 U64bar ( .A1(n162bar), .A2(n161bar), .ZN(n163bar) );
  OR2_X1 U65 ( .A1(n197), .A2(d[6]), .ZN(n161) );
  AND2_X1 U65bar ( .A1(n197bar), .A2(dbar[6]), .ZN(n161bar) );
  OR2_X1 U66 ( .A1(n183), .A2(c[6]), .ZN(n162) );
  AND2_X1 U66bar ( .A1(n183bar), .A2(cbar[6]), .ZN(n162bar) );
  OR2_X1 U67 ( .A1(n160), .A2(n220), .ZN(y[5]) );
  AND2_X1 U67bar ( .A1(n160bar), .A2(n220bar), .ZN(ybar[5]) );
  OR2_X1 U68 ( .A1(n158), .A2(n196), .ZN(n159) );
  AND2_X1 U68bar ( .A1(n158bar), .A2(n196bar), .ZN(n159bar) );
  AND2_X1 U69 ( .A1(n196), .A2(n158), .ZN(n160) );
  OR2_X1 U69bar ( .A1(n196bar), .A2(n158bar), .ZN(n160bar) );
  AND2_X1 U70 ( .A1(n157), .A2(n156), .ZN(n158) );
  OR2_X1 U70bar ( .A1(n157bar), .A2(n156bar), .ZN(n158bar) );
  OR2_X1 U71 ( .A1(n219), .A2(b[5]), .ZN(n156) );
  AND2_X1 U71bar ( .A1(n219bar), .A2(bbar[5]), .ZN(n156bar) );
  OR2_X1 U72 ( .A1(n206), .A2(a[5]), .ZN(n157) );
  AND2_X1 U72bar ( .A1(n206bar), .A2(abar[5]), .ZN(n157bar) );
  AND2_X1 U73 ( .A1(n154), .A2(n153), .ZN(n155) );
  OR2_X1 U73bar ( .A1(n154bar), .A2(n153bar), .ZN(n155bar) );
  OR2_X1 U74 ( .A1(n195), .A2(d[5]), .ZN(n153) );
  AND2_X1 U74bar ( .A1(n195bar), .A2(dbar[5]), .ZN(n153bar) );
  OR2_X1 U75 ( .A1(n182), .A2(c[5]), .ZN(n154) );
  AND2_X1 U75bar ( .A1(n182bar), .A2(cbar[5]), .ZN(n154bar) );
  OR2_X1 U76 ( .A1(n152), .A2(n218), .ZN(y[4]) );
  AND2_X1 U76bar ( .A1(n152bar), .A2(n218bar), .ZN(ybar[4]) );
  OR2_X1 U77 ( .A1(n150), .A2(n194), .ZN(n151) );
  AND2_X1 U77bar ( .A1(n150bar), .A2(n194bar), .ZN(n151bar) );
  AND2_X1 U78 ( .A1(n194), .A2(n150), .ZN(n152) );
  OR2_X1 U78bar ( .A1(n194bar), .A2(n150bar), .ZN(n152bar) );
  AND2_X1 U79 ( .A1(n149), .A2(n148), .ZN(n150) );
  OR2_X1 U79bar ( .A1(n149bar), .A2(n148bar), .ZN(n150bar) );
  OR2_X1 U80 ( .A1(n217), .A2(b[4]), .ZN(n148) );
  AND2_X1 U80bar ( .A1(n217bar), .A2(bbar[4]), .ZN(n148bar) );
  OR2_X1 U81 ( .A1(n205), .A2(a[4]), .ZN(n149) );
  AND2_X1 U81bar ( .A1(n205bar), .A2(abar[4]), .ZN(n149bar) );
  AND2_X1 U82 ( .A1(n146), .A2(n145), .ZN(n147) );
  OR2_X1 U82bar ( .A1(n146bar), .A2(n145bar), .ZN(n147bar) );
  OR2_X1 U83 ( .A1(n193), .A2(d[4]), .ZN(n145) );
  AND2_X1 U83bar ( .A1(n193bar), .A2(dbar[4]), .ZN(n145bar) );
  OR2_X1 U84 ( .A1(n181), .A2(c[4]), .ZN(n146) );
  AND2_X1 U84bar ( .A1(n181bar), .A2(cbar[4]), .ZN(n146bar) );
  OR2_X1 U85 ( .A1(n144), .A2(n216), .ZN(y[3]) );
  AND2_X1 U85bar ( .A1(n144bar), .A2(n216bar), .ZN(ybar[3]) );
  OR2_X1 U86 ( .A1(n142), .A2(n192), .ZN(n143) );
  AND2_X1 U86bar ( .A1(n142bar), .A2(n192bar), .ZN(n143bar) );
  AND2_X1 U87 ( .A1(n192), .A2(n142), .ZN(n144) );
  OR2_X1 U87bar ( .A1(n192bar), .A2(n142bar), .ZN(n144bar) );
  AND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(n142) );
  OR2_X1 U88bar ( .A1(n141bar), .A2(n140bar), .ZN(n142bar) );
  OR2_X1 U89 ( .A1(n215), .A2(b[3]), .ZN(n140) );
  AND2_X1 U89bar ( .A1(n215bar), .A2(bbar[3]), .ZN(n140bar) );
  OR2_X1 U90 ( .A1(n204), .A2(a[3]), .ZN(n141) );
  AND2_X1 U90bar ( .A1(n204bar), .A2(abar[3]), .ZN(n141bar) );
  AND2_X1 U91 ( .A1(n138), .A2(n137), .ZN(n139) );
  OR2_X1 U91bar ( .A1(n138bar), .A2(n137bar), .ZN(n139bar) );
  OR2_X1 U92 ( .A1(n191), .A2(d[3]), .ZN(n137) );
  AND2_X1 U92bar ( .A1(n191bar), .A2(dbar[3]), .ZN(n137bar) );
  OR2_X1 U93 ( .A1(n180), .A2(c[3]), .ZN(n138) );
  AND2_X1 U93bar ( .A1(n180bar), .A2(cbar[3]), .ZN(n138bar) );
  OR2_X1 U94 ( .A1(n136), .A2(n214), .ZN(y[2]) );
  AND2_X1 U94bar ( .A1(n136bar), .A2(n214bar), .ZN(ybar[2]) );
  OR2_X1 U95 ( .A1(n134), .A2(n190), .ZN(n135) );
  AND2_X1 U95bar ( .A1(n134bar), .A2(n190bar), .ZN(n135bar) );
  AND2_X1 U96 ( .A1(n190), .A2(n134), .ZN(n136) );
  OR2_X1 U96bar ( .A1(n190bar), .A2(n134bar), .ZN(n136bar) );
  AND2_X1 U97 ( .A1(n133), .A2(n132), .ZN(n134) );
  OR2_X1 U97bar ( .A1(n133bar), .A2(n132bar), .ZN(n134bar) );
  OR2_X1 U98 ( .A1(n213), .A2(b[2]), .ZN(n132) );
  AND2_X1 U98bar ( .A1(n213bar), .A2(bbar[2]), .ZN(n132bar) );
  OR2_X1 U99 ( .A1(n203), .A2(a[2]), .ZN(n133) );
  AND2_X1 U99bar ( .A1(n203bar), .A2(abar[2]), .ZN(n133bar) );
  AND2_X1 U100 ( .A1(n130), .A2(n129), .ZN(n131) );
  OR2_X1 U100bar ( .A1(n130bar), .A2(n129bar), .ZN(n131bar) );
  OR2_X1 U101 ( .A1(n189), .A2(d[2]), .ZN(n129) );
  AND2_X1 U101bar ( .A1(n189bar), .A2(dbar[2]), .ZN(n129bar) );
  OR2_X1 U102 ( .A1(n179), .A2(c[2]), .ZN(n130) );
  AND2_X1 U102bar ( .A1(n179bar), .A2(cbar[2]), .ZN(n130bar) );
  OR2_X1 U103 ( .A1(n128), .A2(n212), .ZN(y[1]) );
  AND2_X1 U103bar ( .A1(n128bar), .A2(n212bar), .ZN(ybar[1]) );
  OR2_X1 U104 ( .A1(n126), .A2(n188), .ZN(n127) );
  AND2_X1 U104bar ( .A1(n126bar), .A2(n188bar), .ZN(n127bar) );
  AND2_X1 U105 ( .A1(n188), .A2(n126), .ZN(n128) );
  OR2_X1 U105bar ( .A1(n188bar), .A2(n126bar), .ZN(n128bar) );
  AND2_X1 U106 ( .A1(n125), .A2(n124), .ZN(n126) );
  OR2_X1 U106bar ( .A1(n125bar), .A2(n124bar), .ZN(n126bar) );
  OR2_X1 U107 ( .A1(n211), .A2(b[1]), .ZN(n124) );
  AND2_X1 U107bar ( .A1(n211bar), .A2(bbar[1]), .ZN(n124bar) );
  OR2_X1 U108 ( .A1(n202), .A2(a[1]), .ZN(n125) );
  AND2_X1 U108bar ( .A1(n202bar), .A2(abar[1]), .ZN(n125bar) );
  AND2_X1 U109 ( .A1(n122), .A2(n121), .ZN(n123) );
  OR2_X1 U109bar ( .A1(n122bar), .A2(n121bar), .ZN(n123bar) );
  OR2_X1 U110 ( .A1(n187), .A2(d[1]), .ZN(n121) );
  AND2_X1 U110bar ( .A1(n187bar), .A2(dbar[1]), .ZN(n121bar) );
  OR2_X1 U111 ( .A1(n178), .A2(c[1]), .ZN(n122) );
  AND2_X1 U111bar ( .A1(n178bar), .A2(cbar[1]), .ZN(n122bar) );
  OR2_X1 U112 ( .A1(n120), .A2(n210), .ZN(y[0]) );
  AND2_X1 U112bar ( .A1(n120bar), .A2(n210bar), .ZN(ybar[0]) );
  OR2_X1 U113 ( .A1(n118), .A2(n186), .ZN(n119) );
  AND2_X1 U113bar ( .A1(n118bar), .A2(n186bar), .ZN(n119bar) );
  AND2_X1 U114 ( .A1(n186), .A2(n118), .ZN(n120) );
  OR2_X1 U114bar ( .A1(n186bar), .A2(n118bar), .ZN(n120bar) );
  AND2_X1 U115 ( .A1(n117), .A2(n116), .ZN(n118) );
  OR2_X1 U115bar ( .A1(n117bar), .A2(n116bar), .ZN(n118bar) );
  OR2_X1 U116 ( .A1(n209), .A2(b[0]), .ZN(n116) );
  AND2_X1 U116bar ( .A1(n209bar), .A2(bbar[0]), .ZN(n116bar) );
  OR2_X1 U117 ( .A1(n201), .A2(a[0]), .ZN(n117) );
  AND2_X1 U117bar ( .A1(n201bar), .A2(abar[0]), .ZN(n117bar) );
  AND2_X1 U118 ( .A1(n114), .A2(n113), .ZN(n115) );
  OR2_X1 U118bar ( .A1(n114bar), .A2(n113bar), .ZN(n115bar) );
  OR2_X1 U119 ( .A1(n185), .A2(d[0]), .ZN(n113) );
  AND2_X1 U119bar ( .A1(n185bar), .A2(dbar[0]), .ZN(n113bar) );
  OR2_X1 U120 ( .A1(n177), .A2(c[0]), .ZN(n114) );
  AND2_X1 U120bar ( .A1(n177bar), .A2(cbar[0]), .ZN(n114bar) );
endmodule

module byteXor4_11 ( a, b, c, d, y );

  input wire [7:0] a;
  input wire [7:0] b;
  input wire [7:0] c;
  input wire [7:0] d;
  wire [7:0] abar;
  wire [7:0] bbar;
  wire [7:0] cbar;
  wire [7:0] dbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign cbar[0] = ~c[0];
  assign cbar[1] = ~c[1];
  assign cbar[2] = ~c[2];
  assign cbar[3] = ~c[3];
  assign cbar[4] = ~c[4];
  assign cbar[5] = ~c[5];
  assign cbar[6] = ~c[6];
  assign cbar[7] = ~c[7];
  assign dbar[0] = ~d[0];
  assign dbar[1] = ~d[1];
  assign dbar[2] = ~d[2];
  assign dbar[3] = ~d[3];
  assign dbar[4] = ~d[4];
  assign dbar[5] = ~d[5];
  assign dbar[6] = ~d[6];
  assign dbar[7] = ~d[7];
//input_done

  output wire [7:0] y;
  wire [7:0] ybar;
//output_done

  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n113bar;
  wire n114bar;
  wire n115bar;
  wire n116bar;
  wire n117bar;
  wire n118bar;
  wire n119bar;
  wire n120bar;
  wire n121bar;
  wire n122bar;
  wire n123bar;
  wire n124bar;
  wire n125bar;
  wire n126bar;
  wire n127bar;
  wire n128bar;
  wire n129bar;
  wire n130bar;
  wire n131bar;
  wire n132bar;
  wire n133bar;
  wire n134bar;
  wire n135bar;
  wire n136bar;
  wire n137bar;
  wire n138bar;
  wire n139bar;
  wire n140bar;
  wire n141bar;
  wire n142bar;
  wire n143bar;
  wire n144bar;
  wire n145bar;
  wire n146bar;
  wire n147bar;
  wire n148bar;
  wire n149bar;
  wire n150bar;
  wire n151bar;
  wire n152bar;
  wire n153bar;
  wire n154bar;
  wire n155bar;
  wire n156bar;
  wire n157bar;
  wire n158bar;
  wire n159bar;
  wire n160bar;
  wire n161bar;
  wire n162bar;
  wire n163bar;
  wire n164bar;
  wire n165bar;
  wire n166bar;
  wire n167bar;
  wire n168bar;
  wire n169bar;
  wire n170bar;
  wire n171bar;
  wire n172bar;
  wire n173bar;
  wire n174bar;
  wire n175bar;
  wire n176bar;
  wire n177bar;
  wire n178bar;
  wire n179bar;
  wire n180bar;
  wire n181bar;
  wire n182bar;
  wire n183bar;
  wire n184bar;
  wire n185bar;
  wire n186bar;
  wire n187bar;
  wire n188bar;
  wire n189bar;
  wire n190bar;
  wire n191bar;
  wire n192bar;
  wire n193bar;
  wire n194bar;
  wire n195bar;
  wire n196bar;
  wire n197bar;
  wire n198bar;
  wire n199bar;
  wire n200bar;
  wire n201bar;
  wire n202bar;
  wire n203bar;
  wire n204bar;
  wire n205bar;
  wire n206bar;
  wire n207bar;
  wire n208bar;
  wire n209bar;
  wire n210bar;
  wire n211bar;
  wire n212bar;
  wire n213bar;
  wire n214bar;
  wire n215bar;
  wire n216bar;
  wire n217bar;
  wire n218bar;
  wire n219bar;
  wire n220bar;
  wire n221bar;
  wire n222bar;
  wire n223bar;
  wire n224bar;
//wire_done

 //assign_done

  assign n224bar = n175;
  assign n224 = n175bar;
  assign n223bar = a[7];
  assign n223 = abar[7];
  assign n222bar = n167;
  assign n222 = n167bar;
  assign n221bar = a[6];
  assign n221 = abar[6];
  assign n220bar = n159;
  assign n220 = n159bar;
  assign n219bar = a[5];
  assign n219 = abar[5];
  assign n218bar = n151;
  assign n218 = n151bar;
  assign n217bar = a[4];
  assign n217 = abar[4];
  assign n216bar = n143;
  assign n216 = n143bar;
  assign n215bar = a[3];
  assign n215 = abar[3];
  assign n214bar = n135;
  assign n214 = n135bar;
  assign n213bar = a[2];
  assign n213 = abar[2];
  assign n212bar = n127;
  assign n212 = n127bar;
  assign n211bar = a[1];
  assign n211 = abar[1];
  assign n210bar = n119;
  assign n210 = n119bar;
  assign n209bar = a[0];
  assign n209 = abar[0];
  assign n208bar = b[7];
  assign n208 = bbar[7];
  assign n207bar = b[6];
  assign n207 = bbar[6];
  assign n206bar = b[5];
  assign n206 = bbar[5];
  assign n205bar = b[4];
  assign n205 = bbar[4];
  assign n204bar = b[3];
  assign n204 = bbar[3];
  assign n203bar = b[2];
  assign n203 = bbar[2];
  assign n202bar = b[1];
  assign n202 = bbar[1];
  assign n201bar = b[0];
  assign n201 = bbar[0];
  assign n200bar = n171;
  assign n200 = n171bar;
  assign n199bar = c[7];
  assign n199 = cbar[7];
  assign n198bar = n163;
  assign n198 = n163bar;
  assign n197bar = c[6];
  assign n197 = cbar[6];
  assign n196bar = n155;
  assign n196 = n155bar;
  assign n195bar = c[5];
  assign n195 = cbar[5];
  assign n194bar = n147;
  assign n194 = n147bar;
  assign n193bar = c[4];
  assign n193 = cbar[4];
  assign n192bar = n139;
  assign n192 = n139bar;
  assign n191bar = c[3];
  assign n191 = cbar[3];
  assign n190bar = n131;
  assign n190 = n131bar;
  assign n189bar = c[2];
  assign n189 = cbar[2];
  assign n188bar = n123;
  assign n188 = n123bar;
  assign n187bar = c[1];
  assign n187 = cbar[1];
  assign n186bar = n115;
  assign n186 = n115bar;
  assign n185bar = c[0];
  assign n185 = cbar[0];
  assign n184bar = d[7];
  assign n184 = dbar[7];
  assign n183bar = d[6];
  assign n183 = dbar[6];
  assign n182bar = d[5];
  assign n182 = dbar[5];
  assign n181bar = d[4];
  assign n181 = dbar[4];
  assign n180bar = d[3];
  assign n180 = dbar[3];
  assign n179bar = d[2];
  assign n179 = dbar[2];
  assign n178bar = d[1];
  assign n178 = dbar[1];
  assign n177bar = d[0];
  assign n177 = dbar[0];
  OR2_X1 U49 ( .A1(n176), .A2(n224), .ZN(y[7]) );
  AND2_X1 U49bar ( .A1(n176bar), .A2(n224bar), .ZN(ybar[7]) );
  OR2_X1 U50 ( .A1(n174), .A2(n200), .ZN(n175) );
  AND2_X1 U50bar ( .A1(n174bar), .A2(n200bar), .ZN(n175bar) );
  AND2_X1 U51 ( .A1(n200), .A2(n174), .ZN(n176) );
  OR2_X1 U51bar ( .A1(n200bar), .A2(n174bar), .ZN(n176bar) );
  AND2_X1 U52 ( .A1(n173), .A2(n172), .ZN(n174) );
  OR2_X1 U52bar ( .A1(n173bar), .A2(n172bar), .ZN(n174bar) );
  OR2_X1 U53 ( .A1(n223), .A2(b[7]), .ZN(n172) );
  AND2_X1 U53bar ( .A1(n223bar), .A2(bbar[7]), .ZN(n172bar) );
  OR2_X1 U54 ( .A1(n208), .A2(a[7]), .ZN(n173) );
  AND2_X1 U54bar ( .A1(n208bar), .A2(abar[7]), .ZN(n173bar) );
  AND2_X1 U55 ( .A1(n170), .A2(n169), .ZN(n171) );
  OR2_X1 U55bar ( .A1(n170bar), .A2(n169bar), .ZN(n171bar) );
  OR2_X1 U56 ( .A1(n199), .A2(d[7]), .ZN(n169) );
  AND2_X1 U56bar ( .A1(n199bar), .A2(dbar[7]), .ZN(n169bar) );
  OR2_X1 U57 ( .A1(n184), .A2(c[7]), .ZN(n170) );
  AND2_X1 U57bar ( .A1(n184bar), .A2(cbar[7]), .ZN(n170bar) );
  OR2_X1 U58 ( .A1(n168), .A2(n222), .ZN(y[6]) );
  AND2_X1 U58bar ( .A1(n168bar), .A2(n222bar), .ZN(ybar[6]) );
  OR2_X1 U59 ( .A1(n166), .A2(n198), .ZN(n167) );
  AND2_X1 U59bar ( .A1(n166bar), .A2(n198bar), .ZN(n167bar) );
  AND2_X1 U60 ( .A1(n198), .A2(n166), .ZN(n168) );
  OR2_X1 U60bar ( .A1(n198bar), .A2(n166bar), .ZN(n168bar) );
  AND2_X1 U61 ( .A1(n165), .A2(n164), .ZN(n166) );
  OR2_X1 U61bar ( .A1(n165bar), .A2(n164bar), .ZN(n166bar) );
  OR2_X1 U62 ( .A1(n221), .A2(b[6]), .ZN(n164) );
  AND2_X1 U62bar ( .A1(n221bar), .A2(bbar[6]), .ZN(n164bar) );
  OR2_X1 U63 ( .A1(n207), .A2(a[6]), .ZN(n165) );
  AND2_X1 U63bar ( .A1(n207bar), .A2(abar[6]), .ZN(n165bar) );
  AND2_X1 U64 ( .A1(n162), .A2(n161), .ZN(n163) );
  OR2_X1 U64bar ( .A1(n162bar), .A2(n161bar), .ZN(n163bar) );
  OR2_X1 U65 ( .A1(n197), .A2(d[6]), .ZN(n161) );
  AND2_X1 U65bar ( .A1(n197bar), .A2(dbar[6]), .ZN(n161bar) );
  OR2_X1 U66 ( .A1(n183), .A2(c[6]), .ZN(n162) );
  AND2_X1 U66bar ( .A1(n183bar), .A2(cbar[6]), .ZN(n162bar) );
  OR2_X1 U67 ( .A1(n160), .A2(n220), .ZN(y[5]) );
  AND2_X1 U67bar ( .A1(n160bar), .A2(n220bar), .ZN(ybar[5]) );
  OR2_X1 U68 ( .A1(n158), .A2(n196), .ZN(n159) );
  AND2_X1 U68bar ( .A1(n158bar), .A2(n196bar), .ZN(n159bar) );
  AND2_X1 U69 ( .A1(n196), .A2(n158), .ZN(n160) );
  OR2_X1 U69bar ( .A1(n196bar), .A2(n158bar), .ZN(n160bar) );
  AND2_X1 U70 ( .A1(n157), .A2(n156), .ZN(n158) );
  OR2_X1 U70bar ( .A1(n157bar), .A2(n156bar), .ZN(n158bar) );
  OR2_X1 U71 ( .A1(n219), .A2(b[5]), .ZN(n156) );
  AND2_X1 U71bar ( .A1(n219bar), .A2(bbar[5]), .ZN(n156bar) );
  OR2_X1 U72 ( .A1(n206), .A2(a[5]), .ZN(n157) );
  AND2_X1 U72bar ( .A1(n206bar), .A2(abar[5]), .ZN(n157bar) );
  AND2_X1 U73 ( .A1(n154), .A2(n153), .ZN(n155) );
  OR2_X1 U73bar ( .A1(n154bar), .A2(n153bar), .ZN(n155bar) );
  OR2_X1 U74 ( .A1(n195), .A2(d[5]), .ZN(n153) );
  AND2_X1 U74bar ( .A1(n195bar), .A2(dbar[5]), .ZN(n153bar) );
  OR2_X1 U75 ( .A1(n182), .A2(c[5]), .ZN(n154) );
  AND2_X1 U75bar ( .A1(n182bar), .A2(cbar[5]), .ZN(n154bar) );
  OR2_X1 U76 ( .A1(n152), .A2(n218), .ZN(y[4]) );
  AND2_X1 U76bar ( .A1(n152bar), .A2(n218bar), .ZN(ybar[4]) );
  OR2_X1 U77 ( .A1(n150), .A2(n194), .ZN(n151) );
  AND2_X1 U77bar ( .A1(n150bar), .A2(n194bar), .ZN(n151bar) );
  AND2_X1 U78 ( .A1(n194), .A2(n150), .ZN(n152) );
  OR2_X1 U78bar ( .A1(n194bar), .A2(n150bar), .ZN(n152bar) );
  AND2_X1 U79 ( .A1(n149), .A2(n148), .ZN(n150) );
  OR2_X1 U79bar ( .A1(n149bar), .A2(n148bar), .ZN(n150bar) );
  OR2_X1 U80 ( .A1(n217), .A2(b[4]), .ZN(n148) );
  AND2_X1 U80bar ( .A1(n217bar), .A2(bbar[4]), .ZN(n148bar) );
  OR2_X1 U81 ( .A1(n205), .A2(a[4]), .ZN(n149) );
  AND2_X1 U81bar ( .A1(n205bar), .A2(abar[4]), .ZN(n149bar) );
  AND2_X1 U82 ( .A1(n146), .A2(n145), .ZN(n147) );
  OR2_X1 U82bar ( .A1(n146bar), .A2(n145bar), .ZN(n147bar) );
  OR2_X1 U83 ( .A1(n193), .A2(d[4]), .ZN(n145) );
  AND2_X1 U83bar ( .A1(n193bar), .A2(dbar[4]), .ZN(n145bar) );
  OR2_X1 U84 ( .A1(n181), .A2(c[4]), .ZN(n146) );
  AND2_X1 U84bar ( .A1(n181bar), .A2(cbar[4]), .ZN(n146bar) );
  OR2_X1 U85 ( .A1(n144), .A2(n216), .ZN(y[3]) );
  AND2_X1 U85bar ( .A1(n144bar), .A2(n216bar), .ZN(ybar[3]) );
  OR2_X1 U86 ( .A1(n142), .A2(n192), .ZN(n143) );
  AND2_X1 U86bar ( .A1(n142bar), .A2(n192bar), .ZN(n143bar) );
  AND2_X1 U87 ( .A1(n192), .A2(n142), .ZN(n144) );
  OR2_X1 U87bar ( .A1(n192bar), .A2(n142bar), .ZN(n144bar) );
  AND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(n142) );
  OR2_X1 U88bar ( .A1(n141bar), .A2(n140bar), .ZN(n142bar) );
  OR2_X1 U89 ( .A1(n215), .A2(b[3]), .ZN(n140) );
  AND2_X1 U89bar ( .A1(n215bar), .A2(bbar[3]), .ZN(n140bar) );
  OR2_X1 U90 ( .A1(n204), .A2(a[3]), .ZN(n141) );
  AND2_X1 U90bar ( .A1(n204bar), .A2(abar[3]), .ZN(n141bar) );
  AND2_X1 U91 ( .A1(n138), .A2(n137), .ZN(n139) );
  OR2_X1 U91bar ( .A1(n138bar), .A2(n137bar), .ZN(n139bar) );
  OR2_X1 U92 ( .A1(n191), .A2(d[3]), .ZN(n137) );
  AND2_X1 U92bar ( .A1(n191bar), .A2(dbar[3]), .ZN(n137bar) );
  OR2_X1 U93 ( .A1(n180), .A2(c[3]), .ZN(n138) );
  AND2_X1 U93bar ( .A1(n180bar), .A2(cbar[3]), .ZN(n138bar) );
  OR2_X1 U94 ( .A1(n136), .A2(n214), .ZN(y[2]) );
  AND2_X1 U94bar ( .A1(n136bar), .A2(n214bar), .ZN(ybar[2]) );
  OR2_X1 U95 ( .A1(n134), .A2(n190), .ZN(n135) );
  AND2_X1 U95bar ( .A1(n134bar), .A2(n190bar), .ZN(n135bar) );
  AND2_X1 U96 ( .A1(n190), .A2(n134), .ZN(n136) );
  OR2_X1 U96bar ( .A1(n190bar), .A2(n134bar), .ZN(n136bar) );
  AND2_X1 U97 ( .A1(n133), .A2(n132), .ZN(n134) );
  OR2_X1 U97bar ( .A1(n133bar), .A2(n132bar), .ZN(n134bar) );
  OR2_X1 U98 ( .A1(n213), .A2(b[2]), .ZN(n132) );
  AND2_X1 U98bar ( .A1(n213bar), .A2(bbar[2]), .ZN(n132bar) );
  OR2_X1 U99 ( .A1(n203), .A2(a[2]), .ZN(n133) );
  AND2_X1 U99bar ( .A1(n203bar), .A2(abar[2]), .ZN(n133bar) );
  AND2_X1 U100 ( .A1(n130), .A2(n129), .ZN(n131) );
  OR2_X1 U100bar ( .A1(n130bar), .A2(n129bar), .ZN(n131bar) );
  OR2_X1 U101 ( .A1(n189), .A2(d[2]), .ZN(n129) );
  AND2_X1 U101bar ( .A1(n189bar), .A2(dbar[2]), .ZN(n129bar) );
  OR2_X1 U102 ( .A1(n179), .A2(c[2]), .ZN(n130) );
  AND2_X1 U102bar ( .A1(n179bar), .A2(cbar[2]), .ZN(n130bar) );
  OR2_X1 U103 ( .A1(n128), .A2(n212), .ZN(y[1]) );
  AND2_X1 U103bar ( .A1(n128bar), .A2(n212bar), .ZN(ybar[1]) );
  OR2_X1 U104 ( .A1(n126), .A2(n188), .ZN(n127) );
  AND2_X1 U104bar ( .A1(n126bar), .A2(n188bar), .ZN(n127bar) );
  AND2_X1 U105 ( .A1(n188), .A2(n126), .ZN(n128) );
  OR2_X1 U105bar ( .A1(n188bar), .A2(n126bar), .ZN(n128bar) );
  AND2_X1 U106 ( .A1(n125), .A2(n124), .ZN(n126) );
  OR2_X1 U106bar ( .A1(n125bar), .A2(n124bar), .ZN(n126bar) );
  OR2_X1 U107 ( .A1(n211), .A2(b[1]), .ZN(n124) );
  AND2_X1 U107bar ( .A1(n211bar), .A2(bbar[1]), .ZN(n124bar) );
  OR2_X1 U108 ( .A1(n202), .A2(a[1]), .ZN(n125) );
  AND2_X1 U108bar ( .A1(n202bar), .A2(abar[1]), .ZN(n125bar) );
  AND2_X1 U109 ( .A1(n122), .A2(n121), .ZN(n123) );
  OR2_X1 U109bar ( .A1(n122bar), .A2(n121bar), .ZN(n123bar) );
  OR2_X1 U110 ( .A1(n187), .A2(d[1]), .ZN(n121) );
  AND2_X1 U110bar ( .A1(n187bar), .A2(dbar[1]), .ZN(n121bar) );
  OR2_X1 U111 ( .A1(n178), .A2(c[1]), .ZN(n122) );
  AND2_X1 U111bar ( .A1(n178bar), .A2(cbar[1]), .ZN(n122bar) );
  OR2_X1 U112 ( .A1(n120), .A2(n210), .ZN(y[0]) );
  AND2_X1 U112bar ( .A1(n120bar), .A2(n210bar), .ZN(ybar[0]) );
  OR2_X1 U113 ( .A1(n118), .A2(n186), .ZN(n119) );
  AND2_X1 U113bar ( .A1(n118bar), .A2(n186bar), .ZN(n119bar) );
  AND2_X1 U114 ( .A1(n186), .A2(n118), .ZN(n120) );
  OR2_X1 U114bar ( .A1(n186bar), .A2(n118bar), .ZN(n120bar) );
  AND2_X1 U115 ( .A1(n117), .A2(n116), .ZN(n118) );
  OR2_X1 U115bar ( .A1(n117bar), .A2(n116bar), .ZN(n118bar) );
  OR2_X1 U116 ( .A1(n209), .A2(b[0]), .ZN(n116) );
  AND2_X1 U116bar ( .A1(n209bar), .A2(bbar[0]), .ZN(n116bar) );
  OR2_X1 U117 ( .A1(n201), .A2(a[0]), .ZN(n117) );
  AND2_X1 U117bar ( .A1(n201bar), .A2(abar[0]), .ZN(n117bar) );
  AND2_X1 U118 ( .A1(n114), .A2(n113), .ZN(n115) );
  OR2_X1 U118bar ( .A1(n114bar), .A2(n113bar), .ZN(n115bar) );
  OR2_X1 U119 ( .A1(n185), .A2(d[0]), .ZN(n113) );
  AND2_X1 U119bar ( .A1(n185bar), .A2(dbar[0]), .ZN(n113bar) );
  OR2_X1 U120 ( .A1(n177), .A2(c[0]), .ZN(n114) );
  AND2_X1 U120bar ( .A1(n177bar), .A2(cbar[0]), .ZN(n114bar) );
endmodule

module byteXor4_12 ( a, b, c, d, y );

  input wire [7:0] a;
  input wire [7:0] b;
  input wire [7:0] c;
  input wire [7:0] d;
  wire [7:0] abar;
  wire [7:0] bbar;
  wire [7:0] cbar;
  wire [7:0] dbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign cbar[0] = ~c[0];
  assign cbar[1] = ~c[1];
  assign cbar[2] = ~c[2];
  assign cbar[3] = ~c[3];
  assign cbar[4] = ~c[4];
  assign cbar[5] = ~c[5];
  assign cbar[6] = ~c[6];
  assign cbar[7] = ~c[7];
  assign dbar[0] = ~d[0];
  assign dbar[1] = ~d[1];
  assign dbar[2] = ~d[2];
  assign dbar[3] = ~d[3];
  assign dbar[4] = ~d[4];
  assign dbar[5] = ~d[5];
  assign dbar[6] = ~d[6];
  assign dbar[7] = ~d[7];
//input_done

  output wire [7:0] y;
  wire [7:0] ybar;
//output_done

  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n113bar;
  wire n114bar;
  wire n115bar;
  wire n116bar;
  wire n117bar;
  wire n118bar;
  wire n119bar;
  wire n120bar;
  wire n121bar;
  wire n122bar;
  wire n123bar;
  wire n124bar;
  wire n125bar;
  wire n126bar;
  wire n127bar;
  wire n128bar;
  wire n129bar;
  wire n130bar;
  wire n131bar;
  wire n132bar;
  wire n133bar;
  wire n134bar;
  wire n135bar;
  wire n136bar;
  wire n137bar;
  wire n138bar;
  wire n139bar;
  wire n140bar;
  wire n141bar;
  wire n142bar;
  wire n143bar;
  wire n144bar;
  wire n145bar;
  wire n146bar;
  wire n147bar;
  wire n148bar;
  wire n149bar;
  wire n150bar;
  wire n151bar;
  wire n152bar;
  wire n153bar;
  wire n154bar;
  wire n155bar;
  wire n156bar;
  wire n157bar;
  wire n158bar;
  wire n159bar;
  wire n160bar;
  wire n161bar;
  wire n162bar;
  wire n163bar;
  wire n164bar;
  wire n165bar;
  wire n166bar;
  wire n167bar;
  wire n168bar;
  wire n169bar;
  wire n170bar;
  wire n171bar;
  wire n172bar;
  wire n173bar;
  wire n174bar;
  wire n175bar;
  wire n176bar;
  wire n177bar;
  wire n178bar;
  wire n179bar;
  wire n180bar;
  wire n181bar;
  wire n182bar;
  wire n183bar;
  wire n184bar;
  wire n185bar;
  wire n186bar;
  wire n187bar;
  wire n188bar;
  wire n189bar;
  wire n190bar;
  wire n191bar;
  wire n192bar;
  wire n193bar;
  wire n194bar;
  wire n195bar;
  wire n196bar;
  wire n197bar;
  wire n198bar;
  wire n199bar;
  wire n200bar;
  wire n201bar;
  wire n202bar;
  wire n203bar;
  wire n204bar;
  wire n205bar;
  wire n206bar;
  wire n207bar;
  wire n208bar;
  wire n209bar;
  wire n210bar;
  wire n211bar;
  wire n212bar;
  wire n213bar;
  wire n214bar;
  wire n215bar;
  wire n216bar;
  wire n217bar;
  wire n218bar;
  wire n219bar;
  wire n220bar;
  wire n221bar;
  wire n222bar;
  wire n223bar;
  wire n224bar;
//wire_done

 //assign_done

  assign n224bar = n175;
  assign n224 = n175bar;
  assign n223bar = a[7];
  assign n223 = abar[7];
  assign n222bar = n167;
  assign n222 = n167bar;
  assign n221bar = a[6];
  assign n221 = abar[6];
  assign n220bar = n159;
  assign n220 = n159bar;
  assign n219bar = a[5];
  assign n219 = abar[5];
  assign n218bar = n151;
  assign n218 = n151bar;
  assign n217bar = a[4];
  assign n217 = abar[4];
  assign n216bar = n143;
  assign n216 = n143bar;
  assign n215bar = a[3];
  assign n215 = abar[3];
  assign n214bar = n135;
  assign n214 = n135bar;
  assign n213bar = a[2];
  assign n213 = abar[2];
  assign n212bar = n127;
  assign n212 = n127bar;
  assign n211bar = a[1];
  assign n211 = abar[1];
  assign n210bar = n119;
  assign n210 = n119bar;
  assign n209bar = a[0];
  assign n209 = abar[0];
  assign n208bar = b[7];
  assign n208 = bbar[7];
  assign n207bar = b[6];
  assign n207 = bbar[6];
  assign n206bar = b[5];
  assign n206 = bbar[5];
  assign n205bar = b[4];
  assign n205 = bbar[4];
  assign n204bar = b[3];
  assign n204 = bbar[3];
  assign n203bar = b[2];
  assign n203 = bbar[2];
  assign n202bar = b[1];
  assign n202 = bbar[1];
  assign n201bar = b[0];
  assign n201 = bbar[0];
  assign n200bar = n171;
  assign n200 = n171bar;
  assign n199bar = c[7];
  assign n199 = cbar[7];
  assign n198bar = n163;
  assign n198 = n163bar;
  assign n197bar = c[6];
  assign n197 = cbar[6];
  assign n196bar = n155;
  assign n196 = n155bar;
  assign n195bar = c[5];
  assign n195 = cbar[5];
  assign n194bar = n147;
  assign n194 = n147bar;
  assign n193bar = c[4];
  assign n193 = cbar[4];
  assign n192bar = n139;
  assign n192 = n139bar;
  assign n191bar = c[3];
  assign n191 = cbar[3];
  assign n190bar = n131;
  assign n190 = n131bar;
  assign n189bar = c[2];
  assign n189 = cbar[2];
  assign n188bar = n123;
  assign n188 = n123bar;
  assign n187bar = c[1];
  assign n187 = cbar[1];
  assign n186bar = n115;
  assign n186 = n115bar;
  assign n185bar = c[0];
  assign n185 = cbar[0];
  assign n184bar = d[7];
  assign n184 = dbar[7];
  assign n183bar = d[6];
  assign n183 = dbar[6];
  assign n182bar = d[5];
  assign n182 = dbar[5];
  assign n181bar = d[4];
  assign n181 = dbar[4];
  assign n180bar = d[3];
  assign n180 = dbar[3];
  assign n179bar = d[2];
  assign n179 = dbar[2];
  assign n178bar = d[1];
  assign n178 = dbar[1];
  assign n177bar = d[0];
  assign n177 = dbar[0];
  OR2_X1 U49 ( .A1(n176), .A2(n224), .ZN(y[7]) );
  AND2_X1 U49bar ( .A1(n176bar), .A2(n224bar), .ZN(ybar[7]) );
  OR2_X1 U50 ( .A1(n174), .A2(n200), .ZN(n175) );
  AND2_X1 U50bar ( .A1(n174bar), .A2(n200bar), .ZN(n175bar) );
  AND2_X1 U51 ( .A1(n200), .A2(n174), .ZN(n176) );
  OR2_X1 U51bar ( .A1(n200bar), .A2(n174bar), .ZN(n176bar) );
  AND2_X1 U52 ( .A1(n173), .A2(n172), .ZN(n174) );
  OR2_X1 U52bar ( .A1(n173bar), .A2(n172bar), .ZN(n174bar) );
  OR2_X1 U53 ( .A1(n223), .A2(b[7]), .ZN(n172) );
  AND2_X1 U53bar ( .A1(n223bar), .A2(bbar[7]), .ZN(n172bar) );
  OR2_X1 U54 ( .A1(n208), .A2(a[7]), .ZN(n173) );
  AND2_X1 U54bar ( .A1(n208bar), .A2(abar[7]), .ZN(n173bar) );
  AND2_X1 U55 ( .A1(n170), .A2(n169), .ZN(n171) );
  OR2_X1 U55bar ( .A1(n170bar), .A2(n169bar), .ZN(n171bar) );
  OR2_X1 U56 ( .A1(n199), .A2(d[7]), .ZN(n169) );
  AND2_X1 U56bar ( .A1(n199bar), .A2(dbar[7]), .ZN(n169bar) );
  OR2_X1 U57 ( .A1(n184), .A2(c[7]), .ZN(n170) );
  AND2_X1 U57bar ( .A1(n184bar), .A2(cbar[7]), .ZN(n170bar) );
  OR2_X1 U58 ( .A1(n168), .A2(n222), .ZN(y[6]) );
  AND2_X1 U58bar ( .A1(n168bar), .A2(n222bar), .ZN(ybar[6]) );
  OR2_X1 U59 ( .A1(n166), .A2(n198), .ZN(n167) );
  AND2_X1 U59bar ( .A1(n166bar), .A2(n198bar), .ZN(n167bar) );
  AND2_X1 U60 ( .A1(n198), .A2(n166), .ZN(n168) );
  OR2_X1 U60bar ( .A1(n198bar), .A2(n166bar), .ZN(n168bar) );
  AND2_X1 U61 ( .A1(n165), .A2(n164), .ZN(n166) );
  OR2_X1 U61bar ( .A1(n165bar), .A2(n164bar), .ZN(n166bar) );
  OR2_X1 U62 ( .A1(n221), .A2(b[6]), .ZN(n164) );
  AND2_X1 U62bar ( .A1(n221bar), .A2(bbar[6]), .ZN(n164bar) );
  OR2_X1 U63 ( .A1(n207), .A2(a[6]), .ZN(n165) );
  AND2_X1 U63bar ( .A1(n207bar), .A2(abar[6]), .ZN(n165bar) );
  AND2_X1 U64 ( .A1(n162), .A2(n161), .ZN(n163) );
  OR2_X1 U64bar ( .A1(n162bar), .A2(n161bar), .ZN(n163bar) );
  OR2_X1 U65 ( .A1(n197), .A2(d[6]), .ZN(n161) );
  AND2_X1 U65bar ( .A1(n197bar), .A2(dbar[6]), .ZN(n161bar) );
  OR2_X1 U66 ( .A1(n183), .A2(c[6]), .ZN(n162) );
  AND2_X1 U66bar ( .A1(n183bar), .A2(cbar[6]), .ZN(n162bar) );
  OR2_X1 U67 ( .A1(n160), .A2(n220), .ZN(y[5]) );
  AND2_X1 U67bar ( .A1(n160bar), .A2(n220bar), .ZN(ybar[5]) );
  OR2_X1 U68 ( .A1(n158), .A2(n196), .ZN(n159) );
  AND2_X1 U68bar ( .A1(n158bar), .A2(n196bar), .ZN(n159bar) );
  AND2_X1 U69 ( .A1(n196), .A2(n158), .ZN(n160) );
  OR2_X1 U69bar ( .A1(n196bar), .A2(n158bar), .ZN(n160bar) );
  AND2_X1 U70 ( .A1(n157), .A2(n156), .ZN(n158) );
  OR2_X1 U70bar ( .A1(n157bar), .A2(n156bar), .ZN(n158bar) );
  OR2_X1 U71 ( .A1(n219), .A2(b[5]), .ZN(n156) );
  AND2_X1 U71bar ( .A1(n219bar), .A2(bbar[5]), .ZN(n156bar) );
  OR2_X1 U72 ( .A1(n206), .A2(a[5]), .ZN(n157) );
  AND2_X1 U72bar ( .A1(n206bar), .A2(abar[5]), .ZN(n157bar) );
  AND2_X1 U73 ( .A1(n154), .A2(n153), .ZN(n155) );
  OR2_X1 U73bar ( .A1(n154bar), .A2(n153bar), .ZN(n155bar) );
  OR2_X1 U74 ( .A1(n195), .A2(d[5]), .ZN(n153) );
  AND2_X1 U74bar ( .A1(n195bar), .A2(dbar[5]), .ZN(n153bar) );
  OR2_X1 U75 ( .A1(n182), .A2(c[5]), .ZN(n154) );
  AND2_X1 U75bar ( .A1(n182bar), .A2(cbar[5]), .ZN(n154bar) );
  OR2_X1 U76 ( .A1(n152), .A2(n218), .ZN(y[4]) );
  AND2_X1 U76bar ( .A1(n152bar), .A2(n218bar), .ZN(ybar[4]) );
  OR2_X1 U77 ( .A1(n150), .A2(n194), .ZN(n151) );
  AND2_X1 U77bar ( .A1(n150bar), .A2(n194bar), .ZN(n151bar) );
  AND2_X1 U78 ( .A1(n194), .A2(n150), .ZN(n152) );
  OR2_X1 U78bar ( .A1(n194bar), .A2(n150bar), .ZN(n152bar) );
  AND2_X1 U79 ( .A1(n149), .A2(n148), .ZN(n150) );
  OR2_X1 U79bar ( .A1(n149bar), .A2(n148bar), .ZN(n150bar) );
  OR2_X1 U80 ( .A1(n217), .A2(b[4]), .ZN(n148) );
  AND2_X1 U80bar ( .A1(n217bar), .A2(bbar[4]), .ZN(n148bar) );
  OR2_X1 U81 ( .A1(n205), .A2(a[4]), .ZN(n149) );
  AND2_X1 U81bar ( .A1(n205bar), .A2(abar[4]), .ZN(n149bar) );
  AND2_X1 U82 ( .A1(n146), .A2(n145), .ZN(n147) );
  OR2_X1 U82bar ( .A1(n146bar), .A2(n145bar), .ZN(n147bar) );
  OR2_X1 U83 ( .A1(n193), .A2(d[4]), .ZN(n145) );
  AND2_X1 U83bar ( .A1(n193bar), .A2(dbar[4]), .ZN(n145bar) );
  OR2_X1 U84 ( .A1(n181), .A2(c[4]), .ZN(n146) );
  AND2_X1 U84bar ( .A1(n181bar), .A2(cbar[4]), .ZN(n146bar) );
  OR2_X1 U85 ( .A1(n144), .A2(n216), .ZN(y[3]) );
  AND2_X1 U85bar ( .A1(n144bar), .A2(n216bar), .ZN(ybar[3]) );
  OR2_X1 U86 ( .A1(n142), .A2(n192), .ZN(n143) );
  AND2_X1 U86bar ( .A1(n142bar), .A2(n192bar), .ZN(n143bar) );
  AND2_X1 U87 ( .A1(n192), .A2(n142), .ZN(n144) );
  OR2_X1 U87bar ( .A1(n192bar), .A2(n142bar), .ZN(n144bar) );
  AND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(n142) );
  OR2_X1 U88bar ( .A1(n141bar), .A2(n140bar), .ZN(n142bar) );
  OR2_X1 U89 ( .A1(n215), .A2(b[3]), .ZN(n140) );
  AND2_X1 U89bar ( .A1(n215bar), .A2(bbar[3]), .ZN(n140bar) );
  OR2_X1 U90 ( .A1(n204), .A2(a[3]), .ZN(n141) );
  AND2_X1 U90bar ( .A1(n204bar), .A2(abar[3]), .ZN(n141bar) );
  AND2_X1 U91 ( .A1(n138), .A2(n137), .ZN(n139) );
  OR2_X1 U91bar ( .A1(n138bar), .A2(n137bar), .ZN(n139bar) );
  OR2_X1 U92 ( .A1(n191), .A2(d[3]), .ZN(n137) );
  AND2_X1 U92bar ( .A1(n191bar), .A2(dbar[3]), .ZN(n137bar) );
  OR2_X1 U93 ( .A1(n180), .A2(c[3]), .ZN(n138) );
  AND2_X1 U93bar ( .A1(n180bar), .A2(cbar[3]), .ZN(n138bar) );
  OR2_X1 U94 ( .A1(n136), .A2(n214), .ZN(y[2]) );
  AND2_X1 U94bar ( .A1(n136bar), .A2(n214bar), .ZN(ybar[2]) );
  OR2_X1 U95 ( .A1(n134), .A2(n190), .ZN(n135) );
  AND2_X1 U95bar ( .A1(n134bar), .A2(n190bar), .ZN(n135bar) );
  AND2_X1 U96 ( .A1(n190), .A2(n134), .ZN(n136) );
  OR2_X1 U96bar ( .A1(n190bar), .A2(n134bar), .ZN(n136bar) );
  AND2_X1 U97 ( .A1(n133), .A2(n132), .ZN(n134) );
  OR2_X1 U97bar ( .A1(n133bar), .A2(n132bar), .ZN(n134bar) );
  OR2_X1 U98 ( .A1(n213), .A2(b[2]), .ZN(n132) );
  AND2_X1 U98bar ( .A1(n213bar), .A2(bbar[2]), .ZN(n132bar) );
  OR2_X1 U99 ( .A1(n203), .A2(a[2]), .ZN(n133) );
  AND2_X1 U99bar ( .A1(n203bar), .A2(abar[2]), .ZN(n133bar) );
  AND2_X1 U100 ( .A1(n130), .A2(n129), .ZN(n131) );
  OR2_X1 U100bar ( .A1(n130bar), .A2(n129bar), .ZN(n131bar) );
  OR2_X1 U101 ( .A1(n189), .A2(d[2]), .ZN(n129) );
  AND2_X1 U101bar ( .A1(n189bar), .A2(dbar[2]), .ZN(n129bar) );
  OR2_X1 U102 ( .A1(n179), .A2(c[2]), .ZN(n130) );
  AND2_X1 U102bar ( .A1(n179bar), .A2(cbar[2]), .ZN(n130bar) );
  OR2_X1 U103 ( .A1(n128), .A2(n212), .ZN(y[1]) );
  AND2_X1 U103bar ( .A1(n128bar), .A2(n212bar), .ZN(ybar[1]) );
  OR2_X1 U104 ( .A1(n126), .A2(n188), .ZN(n127) );
  AND2_X1 U104bar ( .A1(n126bar), .A2(n188bar), .ZN(n127bar) );
  AND2_X1 U105 ( .A1(n188), .A2(n126), .ZN(n128) );
  OR2_X1 U105bar ( .A1(n188bar), .A2(n126bar), .ZN(n128bar) );
  AND2_X1 U106 ( .A1(n125), .A2(n124), .ZN(n126) );
  OR2_X1 U106bar ( .A1(n125bar), .A2(n124bar), .ZN(n126bar) );
  OR2_X1 U107 ( .A1(n211), .A2(b[1]), .ZN(n124) );
  AND2_X1 U107bar ( .A1(n211bar), .A2(bbar[1]), .ZN(n124bar) );
  OR2_X1 U108 ( .A1(n202), .A2(a[1]), .ZN(n125) );
  AND2_X1 U108bar ( .A1(n202bar), .A2(abar[1]), .ZN(n125bar) );
  AND2_X1 U109 ( .A1(n122), .A2(n121), .ZN(n123) );
  OR2_X1 U109bar ( .A1(n122bar), .A2(n121bar), .ZN(n123bar) );
  OR2_X1 U110 ( .A1(n187), .A2(d[1]), .ZN(n121) );
  AND2_X1 U110bar ( .A1(n187bar), .A2(dbar[1]), .ZN(n121bar) );
  OR2_X1 U111 ( .A1(n178), .A2(c[1]), .ZN(n122) );
  AND2_X1 U111bar ( .A1(n178bar), .A2(cbar[1]), .ZN(n122bar) );
  OR2_X1 U112 ( .A1(n120), .A2(n210), .ZN(y[0]) );
  AND2_X1 U112bar ( .A1(n120bar), .A2(n210bar), .ZN(ybar[0]) );
  OR2_X1 U113 ( .A1(n118), .A2(n186), .ZN(n119) );
  AND2_X1 U113bar ( .A1(n118bar), .A2(n186bar), .ZN(n119bar) );
  AND2_X1 U114 ( .A1(n186), .A2(n118), .ZN(n120) );
  OR2_X1 U114bar ( .A1(n186bar), .A2(n118bar), .ZN(n120bar) );
  AND2_X1 U115 ( .A1(n117), .A2(n116), .ZN(n118) );
  OR2_X1 U115bar ( .A1(n117bar), .A2(n116bar), .ZN(n118bar) );
  OR2_X1 U116 ( .A1(n209), .A2(b[0]), .ZN(n116) );
  AND2_X1 U116bar ( .A1(n209bar), .A2(bbar[0]), .ZN(n116bar) );
  OR2_X1 U117 ( .A1(n201), .A2(a[0]), .ZN(n117) );
  AND2_X1 U117bar ( .A1(n201bar), .A2(abar[0]), .ZN(n117bar) );
  AND2_X1 U118 ( .A1(n114), .A2(n113), .ZN(n115) );
  OR2_X1 U118bar ( .A1(n114bar), .A2(n113bar), .ZN(n115bar) );
  OR2_X1 U119 ( .A1(n185), .A2(d[0]), .ZN(n113) );
  AND2_X1 U119bar ( .A1(n185bar), .A2(dbar[0]), .ZN(n113bar) );
  OR2_X1 U120 ( .A1(n177), .A2(c[0]), .ZN(n114) );
  AND2_X1 U120bar ( .A1(n177bar), .A2(cbar[0]), .ZN(n114bar) );
endmodule

module mixCol_3 ( in, out );

  input wire [31:0] in;
//input_done

  output wire [31:0] out;
//output_done

  wire [7:0] b0_s2;
  wire [7:0] b1_s2;
  wire [7:0] b2_s2;
  wire [7:0] b3_s2;
  wire [7:0] b0_s3;
  wire [7:0] b1_s3;
  wire [7:0] b2_s3;
  wire [7:0] b3_s3;
//wire_done

 //assign_done

  scale2_12 b0_scale2 ( .in(in[31:24]), .out(b0_s2) );
  scale2_11 b1_scale2 ( .in(in[23:16]), .out(b1_s2) );
  scale2_10 b2_scale2 ( .in(in[15:8]), .out(b2_s2) );
  scale2_9 b3_scale2 ( .in(in[7:0]), .out(b3_s2) );
  byteXor_13 b0_scale3 ( .a(in[31:24]), .b(b0_s2), .y(b0_s3) );
  byteXor_12 b1_scale3 ( .a(in[23:16]), .b(b1_s2), .y(b1_s3) );
  byteXor_11 b2_scale3 ( .a(in[15:8]), .b(b2_s2), .y(b2_s3) );
  byteXor_10 b3_scale3 ( .a(in[7:0]), .b(b3_s2), .y(b3_s3) );
  byteXor4_12 out0 ( .a(b0_s2), .b(b1_s3), .c(in[15:8]), .d(in[7:0]), .y(
        out[31:24]) );
  byteXor4_11 out1 ( .a(in[31:24]), .b(b1_s2), .c(b2_s3), .d(in[7:0]), .y(
        out[23:16]) );
  byteXor4_10 out2 ( .a(in[31:24]), .b(in[23:16]), .c(b2_s2), .d(b3_s3), .y(
        out[15:8]) );
  byteXor4_9 out3 ( .a(b0_s3), .b(in[23:16]), .c(in[15:8]), .d(b3_s2), .y(
        out[7:0]) );
endmodule

module mixCol_WDDL ( in, out );

  input wire [127:0] in;
//input_done

  output [127:0] out;
//output_done

//wire_done

 //assign_done

  mixCol_0 m0( .in(in[127:96]), .out(out[127:96]) );
  mixCol_3 m1( .in(in[95:64]), .out(out[95:64]) );
  mixCol_2 m2( .in(in[63:32]), .out(out[63:32]) );
  mixCol_1 m3( .in(in[31:0]), .out(out[31:0]) );
endmodule

//done
