
module CD2_0 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n2)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n2bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n1)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n1bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n1),
    .I1(n2)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n1bar),
    .I1(n2bar)
  );
endmodule

module CD4_0 ( a, b, y );

  input wire [3:0] a;
  input wire [3:0] b;
  wire [3:0] abar;
  wire [3:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
//input_done

  output wire [15:0] y;
  wire [15:0] ybar;
//output_done

//wire_done

  //AND U1
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1 (
    .O(y[9]),
    .I0(b[1]),
    .I1(a[2])
  );
  //OR U1bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1bar (
    .O(ybar[9]),
    .I0(bbar[1]),
    .I1(abar[2])
  );
  //AND U2
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2 (
    .O(y[8]),
    .I0(b[0]),
    .I1(a[2])
  );
  //OR U2bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2bar (
    .O(ybar[8]),
    .I0(bbar[0]),
    .I1(abar[2])
  );
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[7]),
    .I0(b[3]),
    .I1(a[1])
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[7]),
    .I0(bbar[3]),
    .I1(abar[1])
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[6]),
    .I0(b[2]),
    .I1(a[1])
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[6]),
    .I0(bbar[2]),
    .I1(abar[1])
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[5]),
    .I0(a[1]),
    .I1(b[1])
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[5]),
    .I0(abar[1]),
    .I1(bbar[1])
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[4]),
    .I0(a[1]),
    .I1(b[0])
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[4]),
    .I0(abar[1]),
    .I1(bbar[0])
  );
  //AND U7
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7 (
    .O(y[3]),
    .I0(a[0]),
    .I1(b[3])
  );
  //OR U7bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7bar (
    .O(ybar[3]),
    .I0(abar[0]),
    .I1(bbar[3])
  );
  //AND U8
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8 (
    .O(y[2]),
    .I0(a[0]),
    .I1(b[2])
  );
  //OR U8bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8bar (
    .O(ybar[2]),
    .I0(abar[0]),
    .I1(bbar[2])
  );
  //AND U9
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9 (
    .O(y[1]),
    .I0(a[0]),
    .I1(b[1])
  );
  //OR U9bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9bar (
    .O(ybar[1]),
    .I0(abar[0]),
    .I1(bbar[1])
  );
  //AND U10
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10 (
    .O(y[15]),
    .I0(a[3]),
    .I1(b[3])
  );
  //OR U10bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10bar (
    .O(ybar[15]),
    .I0(abar[3]),
    .I1(bbar[3])
  );
  //AND U11
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11 (
    .O(y[14]),
    .I0(a[3]),
    .I1(b[2])
  );
  //OR U11bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11bar (
    .O(ybar[14]),
    .I0(abar[3]),
    .I1(bbar[2])
  );
  //AND U12
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12 (
    .O(y[13]),
    .I0(a[3]),
    .I1(b[1])
  );
  //OR U12bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12bar (
    .O(ybar[13]),
    .I0(abar[3]),
    .I1(bbar[1])
  );
  //AND U13
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13 (
    .O(y[12]),
    .I0(a[3]),
    .I1(b[0])
  );
  //OR U13bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13bar (
    .O(ybar[12]),
    .I0(abar[3]),
    .I1(bbar[0])
  );
  //AND U14
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14 (
    .O(y[11]),
    .I0(b[3]),
    .I1(a[2])
  );
  //OR U14bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14bar (
    .O(ybar[11]),
    .I0(bbar[3]),
    .I1(abar[2])
  );
  //AND U15
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15 (
    .O(y[10]),
    .I0(b[2]),
    .I1(a[2])
  );
  //OR U15bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15bar (
    .O(ybar[10]),
    .I0(bbar[2]),
    .I1(abar[2])
  );
  //AND U16
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16 (
    .O(y[0]),
    .I0(a[0]),
    .I1(b[0])
  );
  //OR U16bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16bar (
    .O(ybar[0]),
    .I0(abar[0]),
    .I1(bbar[0])
  );
endmodule

module CD16_0 ( a, b, y );

  input wire [15:0] a;
  input wire [15:0] b;
  wire [15:0] abar;
  wire [15:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign abar[8] = ~a[8];
  assign abar[9] = ~a[9];
  assign abar[10] = ~a[10];
  assign abar[11] = ~a[11];
  assign abar[12] = ~a[12];
  assign abar[13] = ~a[13];
  assign abar[14] = ~a[14];
  assign abar[15] = ~a[15];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign bbar[8] = ~b[8];
  assign bbar[9] = ~b[9];
  assign bbar[10] = ~b[10];
  assign bbar[11] = ~b[11];
  assign bbar[12] = ~b[12];
  assign bbar[13] = ~b[13];
  assign bbar[14] = ~b[14];
  assign bbar[15] = ~b[15];
//input_done

  output wire [255:0] y;
  wire [255:0] ybar;
//output_done

//wire_done

  //AND U1
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1 (
    .O(y[9]),
    .I0(b[9]),
    .I1(a[0])
  );
  //OR U1bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1bar (
    .O(ybar[9]),
    .I0(bbar[9]),
    .I1(abar[0])
  );
  //AND U2
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2 (
    .O(y[99]),
    .I0(b[3]),
    .I1(a[6])
  );
  //OR U2bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2bar (
    .O(ybar[99]),
    .I0(bbar[3]),
    .I1(abar[6])
  );
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[98]),
    .I0(b[2]),
    .I1(a[6])
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[98]),
    .I0(bbar[2]),
    .I1(abar[6])
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[97]),
    .I0(b[1]),
    .I1(a[6])
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[97]),
    .I0(bbar[1]),
    .I1(abar[6])
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[96]),
    .I0(b[0]),
    .I1(a[6])
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[96]),
    .I0(bbar[0]),
    .I1(abar[6])
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[95]),
    .I0(b[15]),
    .I1(a[5])
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[95]),
    .I0(bbar[15]),
    .I1(abar[5])
  );
  //AND U7
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7 (
    .O(y[94]),
    .I0(b[14]),
    .I1(a[5])
  );
  //OR U7bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7bar (
    .O(ybar[94]),
    .I0(bbar[14]),
    .I1(abar[5])
  );
  //AND U8
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8 (
    .O(y[93]),
    .I0(b[13]),
    .I1(a[5])
  );
  //OR U8bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8bar (
    .O(ybar[93]),
    .I0(bbar[13]),
    .I1(abar[5])
  );
  //AND U9
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9 (
    .O(y[92]),
    .I0(b[12]),
    .I1(a[5])
  );
  //OR U9bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9bar (
    .O(ybar[92]),
    .I0(bbar[12]),
    .I1(abar[5])
  );
  //AND U10
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10 (
    .O(y[91]),
    .I0(b[11]),
    .I1(a[5])
  );
  //OR U10bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10bar (
    .O(ybar[91]),
    .I0(bbar[11]),
    .I1(abar[5])
  );
  //AND U11
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11 (
    .O(y[90]),
    .I0(b[10]),
    .I1(a[5])
  );
  //OR U11bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11bar (
    .O(ybar[90]),
    .I0(bbar[10]),
    .I1(abar[5])
  );
  //AND U12
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12 (
    .O(y[8]),
    .I0(b[8]),
    .I1(a[0])
  );
  //OR U12bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12bar (
    .O(ybar[8]),
    .I0(bbar[8]),
    .I1(abar[0])
  );
  //AND U13
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13 (
    .O(y[89]),
    .I0(a[5]),
    .I1(b[9])
  );
  //OR U13bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13bar (
    .O(ybar[89]),
    .I0(abar[5]),
    .I1(bbar[9])
  );
  //AND U14
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14 (
    .O(y[88]),
    .I0(b[8]),
    .I1(a[5])
  );
  //OR U14bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14bar (
    .O(ybar[88]),
    .I0(bbar[8]),
    .I1(abar[5])
  );
  //AND U15
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15 (
    .O(y[87]),
    .I0(b[7]),
    .I1(a[5])
  );
  //OR U15bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15bar (
    .O(ybar[87]),
    .I0(bbar[7]),
    .I1(abar[5])
  );
  //AND U16
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16 (
    .O(y[86]),
    .I0(b[6]),
    .I1(a[5])
  );
  //OR U16bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16bar (
    .O(ybar[86]),
    .I0(bbar[6]),
    .I1(abar[5])
  );
  //AND U17
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U17 (
    .O(y[85]),
    .I0(b[5]),
    .I1(a[5])
  );
  //OR U17bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U17bar (
    .O(ybar[85]),
    .I0(bbar[5]),
    .I1(abar[5])
  );
  //AND U18
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U18 (
    .O(y[84]),
    .I0(b[4]),
    .I1(a[5])
  );
  //OR U18bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U18bar (
    .O(ybar[84]),
    .I0(bbar[4]),
    .I1(abar[5])
  );
  //AND U19
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U19 (
    .O(y[83]),
    .I0(a[5]),
    .I1(b[3])
  );
  //OR U19bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U19bar (
    .O(ybar[83]),
    .I0(abar[5]),
    .I1(bbar[3])
  );
  //AND U20
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U20 (
    .O(y[82]),
    .I0(a[5]),
    .I1(b[2])
  );
  //OR U20bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U20bar (
    .O(ybar[82]),
    .I0(abar[5]),
    .I1(bbar[2])
  );
  //AND U21
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U21 (
    .O(y[81]),
    .I0(a[5]),
    .I1(b[1])
  );
  //OR U21bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U21bar (
    .O(ybar[81]),
    .I0(abar[5]),
    .I1(bbar[1])
  );
  //AND U22
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U22 (
    .O(y[80]),
    .I0(a[5]),
    .I1(b[0])
  );
  //OR U22bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U22bar (
    .O(ybar[80]),
    .I0(abar[5]),
    .I1(bbar[0])
  );
  //AND U23
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U23 (
    .O(y[7]),
    .I0(b[7]),
    .I1(a[0])
  );
  //OR U23bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U23bar (
    .O(ybar[7]),
    .I0(bbar[7]),
    .I1(abar[0])
  );
  //AND U24
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U24 (
    .O(y[79]),
    .I0(a[4]),
    .I1(b[15])
  );
  //OR U24bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U24bar (
    .O(ybar[79]),
    .I0(abar[4]),
    .I1(bbar[15])
  );
  //AND U25
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U25 (
    .O(y[78]),
    .I0(a[4]),
    .I1(b[14])
  );
  //OR U25bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U25bar (
    .O(ybar[78]),
    .I0(abar[4]),
    .I1(bbar[14])
  );
  //AND U26
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U26 (
    .O(y[77]),
    .I0(a[4]),
    .I1(b[13])
  );
  //OR U26bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U26bar (
    .O(ybar[77]),
    .I0(abar[4]),
    .I1(bbar[13])
  );
  //AND U27
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U27 (
    .O(y[76]),
    .I0(a[4]),
    .I1(b[12])
  );
  //OR U27bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U27bar (
    .O(ybar[76]),
    .I0(abar[4]),
    .I1(bbar[12])
  );
  //AND U28
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U28 (
    .O(y[75]),
    .I0(a[4]),
    .I1(b[11])
  );
  //OR U28bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U28bar (
    .O(ybar[75]),
    .I0(abar[4]),
    .I1(bbar[11])
  );
  //AND U29
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U29 (
    .O(y[74]),
    .I0(a[4]),
    .I1(b[10])
  );
  //OR U29bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U29bar (
    .O(ybar[74]),
    .I0(abar[4]),
    .I1(bbar[10])
  );
  //AND U30
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U30 (
    .O(y[73]),
    .I0(a[4]),
    .I1(b[9])
  );
  //OR U30bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U30bar (
    .O(ybar[73]),
    .I0(abar[4]),
    .I1(bbar[9])
  );
  //AND U31
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U31 (
    .O(y[72]),
    .I0(a[4]),
    .I1(b[8])
  );
  //OR U31bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U31bar (
    .O(ybar[72]),
    .I0(abar[4]),
    .I1(bbar[8])
  );
  //AND U32
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U32 (
    .O(y[71]),
    .I0(a[4]),
    .I1(b[7])
  );
  //OR U32bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U32bar (
    .O(ybar[71]),
    .I0(abar[4]),
    .I1(bbar[7])
  );
  //AND U33
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U33 (
    .O(y[70]),
    .I0(a[4]),
    .I1(b[6])
  );
  //OR U33bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U33bar (
    .O(ybar[70]),
    .I0(abar[4]),
    .I1(bbar[6])
  );
  //AND U34
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U34 (
    .O(y[6]),
    .I0(b[6]),
    .I1(a[0])
  );
  //OR U34bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U34bar (
    .O(ybar[6]),
    .I0(bbar[6]),
    .I1(abar[0])
  );
  //AND U35
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U35 (
    .O(y[69]),
    .I0(a[4]),
    .I1(b[5])
  );
  //OR U35bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U35bar (
    .O(ybar[69]),
    .I0(abar[4]),
    .I1(bbar[5])
  );
  //AND U36
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U36 (
    .O(y[68]),
    .I0(a[4]),
    .I1(b[4])
  );
  //OR U36bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U36bar (
    .O(ybar[68]),
    .I0(abar[4]),
    .I1(bbar[4])
  );
  //AND U37
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U37 (
    .O(y[67]),
    .I0(a[4]),
    .I1(b[3])
  );
  //OR U37bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U37bar (
    .O(ybar[67]),
    .I0(abar[4]),
    .I1(bbar[3])
  );
  //AND U38
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U38 (
    .O(y[66]),
    .I0(a[4]),
    .I1(b[2])
  );
  //OR U38bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U38bar (
    .O(ybar[66]),
    .I0(abar[4]),
    .I1(bbar[2])
  );
  //AND U39
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U39 (
    .O(y[65]),
    .I0(a[4]),
    .I1(b[1])
  );
  //OR U39bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U39bar (
    .O(ybar[65]),
    .I0(abar[4]),
    .I1(bbar[1])
  );
  //AND U40
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U40 (
    .O(y[64]),
    .I0(a[4]),
    .I1(b[0])
  );
  //OR U40bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U40bar (
    .O(ybar[64]),
    .I0(abar[4]),
    .I1(bbar[0])
  );
  //AND U41
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U41 (
    .O(y[63]),
    .I0(a[3]),
    .I1(b[15])
  );
  //OR U41bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U41bar (
    .O(ybar[63]),
    .I0(abar[3]),
    .I1(bbar[15])
  );
  //AND U42
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U42 (
    .O(y[62]),
    .I0(a[3]),
    .I1(b[14])
  );
  //OR U42bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U42bar (
    .O(ybar[62]),
    .I0(abar[3]),
    .I1(bbar[14])
  );
  //AND U43
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U43 (
    .O(y[61]),
    .I0(a[3]),
    .I1(b[13])
  );
  //OR U43bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U43bar (
    .O(ybar[61]),
    .I0(abar[3]),
    .I1(bbar[13])
  );
  //AND U44
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U44 (
    .O(y[60]),
    .I0(a[3]),
    .I1(b[12])
  );
  //OR U44bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U44bar (
    .O(ybar[60]),
    .I0(abar[3]),
    .I1(bbar[12])
  );
  //AND U45
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U45 (
    .O(y[5]),
    .I0(b[5]),
    .I1(a[0])
  );
  //OR U45bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U45bar (
    .O(ybar[5]),
    .I0(bbar[5]),
    .I1(abar[0])
  );
  //AND U46
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U46 (
    .O(y[59]),
    .I0(a[3]),
    .I1(b[11])
  );
  //OR U46bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U46bar (
    .O(ybar[59]),
    .I0(abar[3]),
    .I1(bbar[11])
  );
  //AND U47
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U47 (
    .O(y[58]),
    .I0(a[3]),
    .I1(b[10])
  );
  //OR U47bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U47bar (
    .O(ybar[58]),
    .I0(abar[3]),
    .I1(bbar[10])
  );
  //AND U48
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U48 (
    .O(y[57]),
    .I0(a[3]),
    .I1(b[9])
  );
  //OR U48bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U48bar (
    .O(ybar[57]),
    .I0(abar[3]),
    .I1(bbar[9])
  );
  //AND U49
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U49 (
    .O(y[56]),
    .I0(a[3]),
    .I1(b[8])
  );
  //OR U49bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U49bar (
    .O(ybar[56]),
    .I0(abar[3]),
    .I1(bbar[8])
  );
  //AND U50
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U50 (
    .O(y[55]),
    .I0(a[3]),
    .I1(b[7])
  );
  //OR U50bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U50bar (
    .O(ybar[55]),
    .I0(abar[3]),
    .I1(bbar[7])
  );
  //AND U51
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U51 (
    .O(y[54]),
    .I0(a[3]),
    .I1(b[6])
  );
  //OR U51bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U51bar (
    .O(ybar[54]),
    .I0(abar[3]),
    .I1(bbar[6])
  );
  //AND U52
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U52 (
    .O(y[53]),
    .I0(a[3]),
    .I1(b[5])
  );
  //OR U52bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U52bar (
    .O(ybar[53]),
    .I0(abar[3]),
    .I1(bbar[5])
  );
  //AND U53
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U53 (
    .O(y[52]),
    .I0(a[3]),
    .I1(b[4])
  );
  //OR U53bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U53bar (
    .O(ybar[52]),
    .I0(abar[3]),
    .I1(bbar[4])
  );
  //AND U54
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U54 (
    .O(y[51]),
    .I0(a[3]),
    .I1(b[3])
  );
  //OR U54bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U54bar (
    .O(ybar[51]),
    .I0(abar[3]),
    .I1(bbar[3])
  );
  //AND U55
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U55 (
    .O(y[50]),
    .I0(a[3]),
    .I1(b[2])
  );
  //OR U55bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U55bar (
    .O(ybar[50]),
    .I0(abar[3]),
    .I1(bbar[2])
  );
  //AND U56
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U56 (
    .O(y[4]),
    .I0(b[4]),
    .I1(a[0])
  );
  //OR U56bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U56bar (
    .O(ybar[4]),
    .I0(bbar[4]),
    .I1(abar[0])
  );
  //AND U57
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U57 (
    .O(y[49]),
    .I0(a[3]),
    .I1(b[1])
  );
  //OR U57bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U57bar (
    .O(ybar[49]),
    .I0(abar[3]),
    .I1(bbar[1])
  );
  //AND U58
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U58 (
    .O(y[48]),
    .I0(a[3]),
    .I1(b[0])
  );
  //OR U58bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U58bar (
    .O(ybar[48]),
    .I0(abar[3]),
    .I1(bbar[0])
  );
  //AND U59
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U59 (
    .O(y[47]),
    .I0(a[2]),
    .I1(b[15])
  );
  //OR U59bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U59bar (
    .O(ybar[47]),
    .I0(abar[2]),
    .I1(bbar[15])
  );
  //AND U60
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U60 (
    .O(y[46]),
    .I0(a[2]),
    .I1(b[14])
  );
  //OR U60bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U60bar (
    .O(ybar[46]),
    .I0(abar[2]),
    .I1(bbar[14])
  );
  //AND U61
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U61 (
    .O(y[45]),
    .I0(a[2]),
    .I1(b[13])
  );
  //OR U61bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U61bar (
    .O(ybar[45]),
    .I0(abar[2]),
    .I1(bbar[13])
  );
  //AND U62
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U62 (
    .O(y[44]),
    .I0(a[2]),
    .I1(b[12])
  );
  //OR U62bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U62bar (
    .O(ybar[44]),
    .I0(abar[2]),
    .I1(bbar[12])
  );
  //AND U63
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U63 (
    .O(y[43]),
    .I0(a[2]),
    .I1(b[11])
  );
  //OR U63bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U63bar (
    .O(ybar[43]),
    .I0(abar[2]),
    .I1(bbar[11])
  );
  //AND U64
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U64 (
    .O(y[42]),
    .I0(a[2]),
    .I1(b[10])
  );
  //OR U64bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U64bar (
    .O(ybar[42]),
    .I0(abar[2]),
    .I1(bbar[10])
  );
  //AND U65
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U65 (
    .O(y[41]),
    .I0(a[2]),
    .I1(b[9])
  );
  //OR U65bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U65bar (
    .O(ybar[41]),
    .I0(abar[2]),
    .I1(bbar[9])
  );
  //AND U66
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U66 (
    .O(y[40]),
    .I0(a[2]),
    .I1(b[8])
  );
  //OR U66bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U66bar (
    .O(ybar[40]),
    .I0(abar[2]),
    .I1(bbar[8])
  );
  //AND U67
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U67 (
    .O(y[3]),
    .I0(b[3]),
    .I1(a[0])
  );
  //OR U67bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U67bar (
    .O(ybar[3]),
    .I0(bbar[3]),
    .I1(abar[0])
  );
  //AND U68
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U68 (
    .O(y[39]),
    .I0(a[2]),
    .I1(b[7])
  );
  //OR U68bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U68bar (
    .O(ybar[39]),
    .I0(abar[2]),
    .I1(bbar[7])
  );
  //AND U69
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U69 (
    .O(y[38]),
    .I0(a[2]),
    .I1(b[6])
  );
  //OR U69bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U69bar (
    .O(ybar[38]),
    .I0(abar[2]),
    .I1(bbar[6])
  );
  //AND U70
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U70 (
    .O(y[37]),
    .I0(a[2]),
    .I1(b[5])
  );
  //OR U70bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U70bar (
    .O(ybar[37]),
    .I0(abar[2]),
    .I1(bbar[5])
  );
  //AND U71
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U71 (
    .O(y[36]),
    .I0(a[2]),
    .I1(b[4])
  );
  //OR U71bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U71bar (
    .O(ybar[36]),
    .I0(abar[2]),
    .I1(bbar[4])
  );
  //AND U72
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U72 (
    .O(y[35]),
    .I0(a[2]),
    .I1(b[3])
  );
  //OR U72bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U72bar (
    .O(ybar[35]),
    .I0(abar[2]),
    .I1(bbar[3])
  );
  //AND U73
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U73 (
    .O(y[34]),
    .I0(a[2]),
    .I1(b[2])
  );
  //OR U73bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U73bar (
    .O(ybar[34]),
    .I0(abar[2]),
    .I1(bbar[2])
  );
  //AND U74
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U74 (
    .O(y[33]),
    .I0(a[2]),
    .I1(b[1])
  );
  //OR U74bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U74bar (
    .O(ybar[33]),
    .I0(abar[2]),
    .I1(bbar[1])
  );
  //AND U75
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U75 (
    .O(y[32]),
    .I0(a[2]),
    .I1(b[0])
  );
  //OR U75bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U75bar (
    .O(ybar[32]),
    .I0(abar[2]),
    .I1(bbar[0])
  );
  //AND U76
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U76 (
    .O(y[31]),
    .I0(a[1]),
    .I1(b[15])
  );
  //OR U76bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U76bar (
    .O(ybar[31]),
    .I0(abar[1]),
    .I1(bbar[15])
  );
  //AND U77
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U77 (
    .O(y[30]),
    .I0(a[1]),
    .I1(b[14])
  );
  //OR U77bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U77bar (
    .O(ybar[30]),
    .I0(abar[1]),
    .I1(bbar[14])
  );
  //AND U78
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U78 (
    .O(y[2]),
    .I0(b[2]),
    .I1(a[0])
  );
  //OR U78bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U78bar (
    .O(ybar[2]),
    .I0(bbar[2]),
    .I1(abar[0])
  );
  //AND U79
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U79 (
    .O(y[29]),
    .I0(a[1]),
    .I1(b[13])
  );
  //OR U79bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U79bar (
    .O(ybar[29]),
    .I0(abar[1]),
    .I1(bbar[13])
  );
  //AND U80
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U80 (
    .O(y[28]),
    .I0(a[1]),
    .I1(b[12])
  );
  //OR U80bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U80bar (
    .O(ybar[28]),
    .I0(abar[1]),
    .I1(bbar[12])
  );
  //AND U81
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U81 (
    .O(y[27]),
    .I0(a[1]),
    .I1(b[11])
  );
  //OR U81bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U81bar (
    .O(ybar[27]),
    .I0(abar[1]),
    .I1(bbar[11])
  );
  //AND U82
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U82 (
    .O(y[26]),
    .I0(a[1]),
    .I1(b[10])
  );
  //OR U82bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U82bar (
    .O(ybar[26]),
    .I0(abar[1]),
    .I1(bbar[10])
  );
  //AND U83
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U83 (
    .O(y[25]),
    .I0(a[1]),
    .I1(b[9])
  );
  //OR U83bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U83bar (
    .O(ybar[25]),
    .I0(abar[1]),
    .I1(bbar[9])
  );
  //AND U84
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U84 (
    .O(y[255]),
    .I0(a[15]),
    .I1(b[15])
  );
  //OR U84bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U84bar (
    .O(ybar[255]),
    .I0(abar[15]),
    .I1(bbar[15])
  );
  //AND U85
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U85 (
    .O(y[254]),
    .I0(a[15]),
    .I1(b[14])
  );
  //OR U85bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U85bar (
    .O(ybar[254]),
    .I0(abar[15]),
    .I1(bbar[14])
  );
  //AND U86
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U86 (
    .O(y[253]),
    .I0(a[15]),
    .I1(b[13])
  );
  //OR U86bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U86bar (
    .O(ybar[253]),
    .I0(abar[15]),
    .I1(bbar[13])
  );
  //AND U87
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U87 (
    .O(y[252]),
    .I0(a[15]),
    .I1(b[12])
  );
  //OR U87bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U87bar (
    .O(ybar[252]),
    .I0(abar[15]),
    .I1(bbar[12])
  );
  //AND U88
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U88 (
    .O(y[251]),
    .I0(a[15]),
    .I1(b[11])
  );
  //OR U88bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U88bar (
    .O(ybar[251]),
    .I0(abar[15]),
    .I1(bbar[11])
  );
  //AND U89
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U89 (
    .O(y[250]),
    .I0(a[15]),
    .I1(b[10])
  );
  //OR U89bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U89bar (
    .O(ybar[250]),
    .I0(abar[15]),
    .I1(bbar[10])
  );
  //AND U90
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U90 (
    .O(y[24]),
    .I0(a[1]),
    .I1(b[8])
  );
  //OR U90bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U90bar (
    .O(ybar[24]),
    .I0(abar[1]),
    .I1(bbar[8])
  );
  //AND U91
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U91 (
    .O(y[249]),
    .I0(a[15]),
    .I1(b[9])
  );
  //OR U91bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U91bar (
    .O(ybar[249]),
    .I0(abar[15]),
    .I1(bbar[9])
  );
  //AND U92
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U92 (
    .O(y[248]),
    .I0(a[15]),
    .I1(b[8])
  );
  //OR U92bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U92bar (
    .O(ybar[248]),
    .I0(abar[15]),
    .I1(bbar[8])
  );
  //AND U93
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U93 (
    .O(y[247]),
    .I0(a[15]),
    .I1(b[7])
  );
  //OR U93bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U93bar (
    .O(ybar[247]),
    .I0(abar[15]),
    .I1(bbar[7])
  );
  //AND U94
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U94 (
    .O(y[246]),
    .I0(a[15]),
    .I1(b[6])
  );
  //OR U94bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U94bar (
    .O(ybar[246]),
    .I0(abar[15]),
    .I1(bbar[6])
  );
  //AND U95
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U95 (
    .O(y[245]),
    .I0(a[15]),
    .I1(b[5])
  );
  //OR U95bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U95bar (
    .O(ybar[245]),
    .I0(abar[15]),
    .I1(bbar[5])
  );
  //AND U96
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U96 (
    .O(y[244]),
    .I0(a[15]),
    .I1(b[4])
  );
  //OR U96bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U96bar (
    .O(ybar[244]),
    .I0(abar[15]),
    .I1(bbar[4])
  );
  //AND U97
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U97 (
    .O(y[243]),
    .I0(a[15]),
    .I1(b[3])
  );
  //OR U97bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U97bar (
    .O(ybar[243]),
    .I0(abar[15]),
    .I1(bbar[3])
  );
  //AND U98
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U98 (
    .O(y[242]),
    .I0(a[15]),
    .I1(b[2])
  );
  //OR U98bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U98bar (
    .O(ybar[242]),
    .I0(abar[15]),
    .I1(bbar[2])
  );
  //AND U99
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U99 (
    .O(y[241]),
    .I0(a[15]),
    .I1(b[1])
  );
  //OR U99bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U99bar (
    .O(ybar[241]),
    .I0(abar[15]),
    .I1(bbar[1])
  );
  //AND U100
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U100 (
    .O(y[240]),
    .I0(a[15]),
    .I1(b[0])
  );
  //OR U100bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U100bar (
    .O(ybar[240]),
    .I0(abar[15]),
    .I1(bbar[0])
  );
  //AND U101
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U101 (
    .O(y[23]),
    .I0(a[1]),
    .I1(b[7])
  );
  //OR U101bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U101bar (
    .O(ybar[23]),
    .I0(abar[1]),
    .I1(bbar[7])
  );
  //AND U102
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U102 (
    .O(y[239]),
    .I0(a[14]),
    .I1(b[15])
  );
  //OR U102bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U102bar (
    .O(ybar[239]),
    .I0(abar[14]),
    .I1(bbar[15])
  );
  //AND U103
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U103 (
    .O(y[238]),
    .I0(a[14]),
    .I1(b[14])
  );
  //OR U103bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U103bar (
    .O(ybar[238]),
    .I0(abar[14]),
    .I1(bbar[14])
  );
  //AND U104
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U104 (
    .O(y[237]),
    .I0(a[14]),
    .I1(b[13])
  );
  //OR U104bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U104bar (
    .O(ybar[237]),
    .I0(abar[14]),
    .I1(bbar[13])
  );
  //AND U105
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U105 (
    .O(y[236]),
    .I0(a[14]),
    .I1(b[12])
  );
  //OR U105bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U105bar (
    .O(ybar[236]),
    .I0(abar[14]),
    .I1(bbar[12])
  );
  //AND U106
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U106 (
    .O(y[235]),
    .I0(a[14]),
    .I1(b[11])
  );
  //OR U106bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U106bar (
    .O(ybar[235]),
    .I0(abar[14]),
    .I1(bbar[11])
  );
  //AND U107
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U107 (
    .O(y[234]),
    .I0(a[14]),
    .I1(b[10])
  );
  //OR U107bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U107bar (
    .O(ybar[234]),
    .I0(abar[14]),
    .I1(bbar[10])
  );
  //AND U108
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U108 (
    .O(y[233]),
    .I0(a[14]),
    .I1(b[9])
  );
  //OR U108bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U108bar (
    .O(ybar[233]),
    .I0(abar[14]),
    .I1(bbar[9])
  );
  //AND U109
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U109 (
    .O(y[232]),
    .I0(a[14]),
    .I1(b[8])
  );
  //OR U109bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U109bar (
    .O(ybar[232]),
    .I0(abar[14]),
    .I1(bbar[8])
  );
  //AND U110
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U110 (
    .O(y[231]),
    .I0(a[14]),
    .I1(b[7])
  );
  //OR U110bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U110bar (
    .O(ybar[231]),
    .I0(abar[14]),
    .I1(bbar[7])
  );
  //AND U111
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U111 (
    .O(y[230]),
    .I0(a[14]),
    .I1(b[6])
  );
  //OR U111bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U111bar (
    .O(ybar[230]),
    .I0(abar[14]),
    .I1(bbar[6])
  );
  //AND U112
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U112 (
    .O(y[22]),
    .I0(a[1]),
    .I1(b[6])
  );
  //OR U112bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U112bar (
    .O(ybar[22]),
    .I0(abar[1]),
    .I1(bbar[6])
  );
  //AND U113
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U113 (
    .O(y[229]),
    .I0(a[14]),
    .I1(b[5])
  );
  //OR U113bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U113bar (
    .O(ybar[229]),
    .I0(abar[14]),
    .I1(bbar[5])
  );
  //AND U114
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U114 (
    .O(y[228]),
    .I0(a[14]),
    .I1(b[4])
  );
  //OR U114bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U114bar (
    .O(ybar[228]),
    .I0(abar[14]),
    .I1(bbar[4])
  );
  //AND U115
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U115 (
    .O(y[227]),
    .I0(a[14]),
    .I1(b[3])
  );
  //OR U115bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U115bar (
    .O(ybar[227]),
    .I0(abar[14]),
    .I1(bbar[3])
  );
  //AND U116
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U116 (
    .O(y[226]),
    .I0(a[14]),
    .I1(b[2])
  );
  //OR U116bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U116bar (
    .O(ybar[226]),
    .I0(abar[14]),
    .I1(bbar[2])
  );
  //AND U117
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U117 (
    .O(y[225]),
    .I0(a[14]),
    .I1(b[1])
  );
  //OR U117bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U117bar (
    .O(ybar[225]),
    .I0(abar[14]),
    .I1(bbar[1])
  );
  //AND U118
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U118 (
    .O(y[224]),
    .I0(a[14]),
    .I1(b[0])
  );
  //OR U118bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U118bar (
    .O(ybar[224]),
    .I0(abar[14]),
    .I1(bbar[0])
  );
  //AND U119
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U119 (
    .O(y[223]),
    .I0(a[13]),
    .I1(b[15])
  );
  //OR U119bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U119bar (
    .O(ybar[223]),
    .I0(abar[13]),
    .I1(bbar[15])
  );
  //AND U120
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U120 (
    .O(y[222]),
    .I0(a[13]),
    .I1(b[14])
  );
  //OR U120bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U120bar (
    .O(ybar[222]),
    .I0(abar[13]),
    .I1(bbar[14])
  );
  //AND U121
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U121 (
    .O(y[221]),
    .I0(a[13]),
    .I1(b[13])
  );
  //OR U121bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U121bar (
    .O(ybar[221]),
    .I0(abar[13]),
    .I1(bbar[13])
  );
  //AND U122
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U122 (
    .O(y[220]),
    .I0(a[13]),
    .I1(b[12])
  );
  //OR U122bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U122bar (
    .O(ybar[220]),
    .I0(abar[13]),
    .I1(bbar[12])
  );
  //AND U123
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U123 (
    .O(y[21]),
    .I0(a[1]),
    .I1(b[5])
  );
  //OR U123bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U123bar (
    .O(ybar[21]),
    .I0(abar[1]),
    .I1(bbar[5])
  );
  //AND U124
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U124 (
    .O(y[219]),
    .I0(a[13]),
    .I1(b[11])
  );
  //OR U124bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U124bar (
    .O(ybar[219]),
    .I0(abar[13]),
    .I1(bbar[11])
  );
  //AND U125
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U125 (
    .O(y[218]),
    .I0(a[13]),
    .I1(b[10])
  );
  //OR U125bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U125bar (
    .O(ybar[218]),
    .I0(abar[13]),
    .I1(bbar[10])
  );
  //AND U126
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U126 (
    .O(y[217]),
    .I0(a[13]),
    .I1(b[9])
  );
  //OR U126bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U126bar (
    .O(ybar[217]),
    .I0(abar[13]),
    .I1(bbar[9])
  );
  //AND U127
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U127 (
    .O(y[216]),
    .I0(a[13]),
    .I1(b[8])
  );
  //OR U127bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U127bar (
    .O(ybar[216]),
    .I0(abar[13]),
    .I1(bbar[8])
  );
  //AND U128
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U128 (
    .O(y[215]),
    .I0(a[13]),
    .I1(b[7])
  );
  //OR U128bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U128bar (
    .O(ybar[215]),
    .I0(abar[13]),
    .I1(bbar[7])
  );
  //AND U129
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U129 (
    .O(y[214]),
    .I0(a[13]),
    .I1(b[6])
  );
  //OR U129bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U129bar (
    .O(ybar[214]),
    .I0(abar[13]),
    .I1(bbar[6])
  );
  //AND U130
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U130 (
    .O(y[213]),
    .I0(a[13]),
    .I1(b[5])
  );
  //OR U130bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U130bar (
    .O(ybar[213]),
    .I0(abar[13]),
    .I1(bbar[5])
  );
  //AND U131
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U131 (
    .O(y[212]),
    .I0(a[13]),
    .I1(b[4])
  );
  //OR U131bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U131bar (
    .O(ybar[212]),
    .I0(abar[13]),
    .I1(bbar[4])
  );
  //AND U132
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U132 (
    .O(y[211]),
    .I0(a[13]),
    .I1(b[3])
  );
  //OR U132bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U132bar (
    .O(ybar[211]),
    .I0(abar[13]),
    .I1(bbar[3])
  );
  //AND U133
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U133 (
    .O(y[210]),
    .I0(a[13]),
    .I1(b[2])
  );
  //OR U133bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U133bar (
    .O(ybar[210]),
    .I0(abar[13]),
    .I1(bbar[2])
  );
  //AND U134
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U134 (
    .O(y[20]),
    .I0(a[1]),
    .I1(b[4])
  );
  //OR U134bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U134bar (
    .O(ybar[20]),
    .I0(abar[1]),
    .I1(bbar[4])
  );
  //AND U135
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U135 (
    .O(y[209]),
    .I0(a[13]),
    .I1(b[1])
  );
  //OR U135bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U135bar (
    .O(ybar[209]),
    .I0(abar[13]),
    .I1(bbar[1])
  );
  //AND U136
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U136 (
    .O(y[208]),
    .I0(a[13]),
    .I1(b[0])
  );
  //OR U136bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U136bar (
    .O(ybar[208]),
    .I0(abar[13]),
    .I1(bbar[0])
  );
  //AND U137
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U137 (
    .O(y[207]),
    .I0(a[12]),
    .I1(b[15])
  );
  //OR U137bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U137bar (
    .O(ybar[207]),
    .I0(abar[12]),
    .I1(bbar[15])
  );
  //AND U138
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U138 (
    .O(y[206]),
    .I0(a[12]),
    .I1(b[14])
  );
  //OR U138bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U138bar (
    .O(ybar[206]),
    .I0(abar[12]),
    .I1(bbar[14])
  );
  //AND U139
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U139 (
    .O(y[205]),
    .I0(a[12]),
    .I1(b[13])
  );
  //OR U139bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U139bar (
    .O(ybar[205]),
    .I0(abar[12]),
    .I1(bbar[13])
  );
  //AND U140
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U140 (
    .O(y[204]),
    .I0(a[12]),
    .I1(b[12])
  );
  //OR U140bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U140bar (
    .O(ybar[204]),
    .I0(abar[12]),
    .I1(bbar[12])
  );
  //AND U141
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U141 (
    .O(y[203]),
    .I0(a[12]),
    .I1(b[11])
  );
  //OR U141bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U141bar (
    .O(ybar[203]),
    .I0(abar[12]),
    .I1(bbar[11])
  );
  //AND U142
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U142 (
    .O(y[202]),
    .I0(a[12]),
    .I1(b[10])
  );
  //OR U142bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U142bar (
    .O(ybar[202]),
    .I0(abar[12]),
    .I1(bbar[10])
  );
  //AND U143
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U143 (
    .O(y[201]),
    .I0(a[12]),
    .I1(b[9])
  );
  //OR U143bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U143bar (
    .O(ybar[201]),
    .I0(abar[12]),
    .I1(bbar[9])
  );
  //AND U144
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U144 (
    .O(y[200]),
    .I0(a[12]),
    .I1(b[8])
  );
  //OR U144bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U144bar (
    .O(ybar[200]),
    .I0(abar[12]),
    .I1(bbar[8])
  );
  //AND U145
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U145 (
    .O(y[1]),
    .I0(b[1]),
    .I1(a[0])
  );
  //OR U145bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U145bar (
    .O(ybar[1]),
    .I0(bbar[1]),
    .I1(abar[0])
  );
  //AND U146
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U146 (
    .O(y[19]),
    .I0(a[1]),
    .I1(b[3])
  );
  //OR U146bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U146bar (
    .O(ybar[19]),
    .I0(abar[1]),
    .I1(bbar[3])
  );
  //AND U147
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U147 (
    .O(y[199]),
    .I0(a[12]),
    .I1(b[7])
  );
  //OR U147bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U147bar (
    .O(ybar[199]),
    .I0(abar[12]),
    .I1(bbar[7])
  );
  //AND U148
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U148 (
    .O(y[198]),
    .I0(a[12]),
    .I1(b[6])
  );
  //OR U148bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U148bar (
    .O(ybar[198]),
    .I0(abar[12]),
    .I1(bbar[6])
  );
  //AND U149
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U149 (
    .O(y[197]),
    .I0(a[12]),
    .I1(b[5])
  );
  //OR U149bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U149bar (
    .O(ybar[197]),
    .I0(abar[12]),
    .I1(bbar[5])
  );
  //AND U150
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U150 (
    .O(y[196]),
    .I0(a[12]),
    .I1(b[4])
  );
  //OR U150bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U150bar (
    .O(ybar[196]),
    .I0(abar[12]),
    .I1(bbar[4])
  );
  //AND U151
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U151 (
    .O(y[195]),
    .I0(a[12]),
    .I1(b[3])
  );
  //OR U151bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U151bar (
    .O(ybar[195]),
    .I0(abar[12]),
    .I1(bbar[3])
  );
  //AND U152
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U152 (
    .O(y[194]),
    .I0(a[12]),
    .I1(b[2])
  );
  //OR U152bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U152bar (
    .O(ybar[194]),
    .I0(abar[12]),
    .I1(bbar[2])
  );
  //AND U153
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U153 (
    .O(y[193]),
    .I0(a[12]),
    .I1(b[1])
  );
  //OR U153bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U153bar (
    .O(ybar[193]),
    .I0(abar[12]),
    .I1(bbar[1])
  );
  //AND U154
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U154 (
    .O(y[192]),
    .I0(a[12]),
    .I1(b[0])
  );
  //OR U154bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U154bar (
    .O(ybar[192]),
    .I0(abar[12]),
    .I1(bbar[0])
  );
  //AND U155
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U155 (
    .O(y[191]),
    .I0(a[11]),
    .I1(b[15])
  );
  //OR U155bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U155bar (
    .O(ybar[191]),
    .I0(abar[11]),
    .I1(bbar[15])
  );
  //AND U156
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U156 (
    .O(y[190]),
    .I0(a[11]),
    .I1(b[14])
  );
  //OR U156bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U156bar (
    .O(ybar[190]),
    .I0(abar[11]),
    .I1(bbar[14])
  );
  //AND U157
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U157 (
    .O(y[18]),
    .I0(a[1]),
    .I1(b[2])
  );
  //OR U157bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U157bar (
    .O(ybar[18]),
    .I0(abar[1]),
    .I1(bbar[2])
  );
  //AND U158
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U158 (
    .O(y[189]),
    .I0(a[11]),
    .I1(b[13])
  );
  //OR U158bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U158bar (
    .O(ybar[189]),
    .I0(abar[11]),
    .I1(bbar[13])
  );
  //AND U159
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U159 (
    .O(y[188]),
    .I0(a[11]),
    .I1(b[12])
  );
  //OR U159bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U159bar (
    .O(ybar[188]),
    .I0(abar[11]),
    .I1(bbar[12])
  );
  //AND U160
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U160 (
    .O(y[187]),
    .I0(a[11]),
    .I1(b[11])
  );
  //OR U160bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U160bar (
    .O(ybar[187]),
    .I0(abar[11]),
    .I1(bbar[11])
  );
  //AND U161
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U161 (
    .O(y[186]),
    .I0(a[11]),
    .I1(b[10])
  );
  //OR U161bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U161bar (
    .O(ybar[186]),
    .I0(abar[11]),
    .I1(bbar[10])
  );
  //AND U162
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U162 (
    .O(y[185]),
    .I0(a[11]),
    .I1(b[9])
  );
  //OR U162bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U162bar (
    .O(ybar[185]),
    .I0(abar[11]),
    .I1(bbar[9])
  );
  //AND U163
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U163 (
    .O(y[184]),
    .I0(a[11]),
    .I1(b[8])
  );
  //OR U163bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U163bar (
    .O(ybar[184]),
    .I0(abar[11]),
    .I1(bbar[8])
  );
  //AND U164
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U164 (
    .O(y[183]),
    .I0(a[11]),
    .I1(b[7])
  );
  //OR U164bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U164bar (
    .O(ybar[183]),
    .I0(abar[11]),
    .I1(bbar[7])
  );
  //AND U165
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U165 (
    .O(y[182]),
    .I0(a[11]),
    .I1(b[6])
  );
  //OR U165bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U165bar (
    .O(ybar[182]),
    .I0(abar[11]),
    .I1(bbar[6])
  );
  //AND U166
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U166 (
    .O(y[181]),
    .I0(a[11]),
    .I1(b[5])
  );
  //OR U166bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U166bar (
    .O(ybar[181]),
    .I0(abar[11]),
    .I1(bbar[5])
  );
  //AND U167
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U167 (
    .O(y[180]),
    .I0(a[11]),
    .I1(b[4])
  );
  //OR U167bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U167bar (
    .O(ybar[180]),
    .I0(abar[11]),
    .I1(bbar[4])
  );
  //AND U168
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U168 (
    .O(y[17]),
    .I0(a[1]),
    .I1(b[1])
  );
  //OR U168bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U168bar (
    .O(ybar[17]),
    .I0(abar[1]),
    .I1(bbar[1])
  );
  //AND U169
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U169 (
    .O(y[179]),
    .I0(a[11]),
    .I1(b[3])
  );
  //OR U169bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U169bar (
    .O(ybar[179]),
    .I0(abar[11]),
    .I1(bbar[3])
  );
  //AND U170
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U170 (
    .O(y[178]),
    .I0(a[11]),
    .I1(b[2])
  );
  //OR U170bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U170bar (
    .O(ybar[178]),
    .I0(abar[11]),
    .I1(bbar[2])
  );
  //AND U171
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U171 (
    .O(y[177]),
    .I0(a[11]),
    .I1(b[1])
  );
  //OR U171bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U171bar (
    .O(ybar[177]),
    .I0(abar[11]),
    .I1(bbar[1])
  );
  //AND U172
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U172 (
    .O(y[176]),
    .I0(a[11]),
    .I1(b[0])
  );
  //OR U172bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U172bar (
    .O(ybar[176]),
    .I0(abar[11]),
    .I1(bbar[0])
  );
  //AND U173
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U173 (
    .O(y[175]),
    .I0(a[10]),
    .I1(b[15])
  );
  //OR U173bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U173bar (
    .O(ybar[175]),
    .I0(abar[10]),
    .I1(bbar[15])
  );
  //AND U174
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U174 (
    .O(y[174]),
    .I0(a[10]),
    .I1(b[14])
  );
  //OR U174bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U174bar (
    .O(ybar[174]),
    .I0(abar[10]),
    .I1(bbar[14])
  );
  //AND U175
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U175 (
    .O(y[173]),
    .I0(a[10]),
    .I1(b[13])
  );
  //OR U175bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U175bar (
    .O(ybar[173]),
    .I0(abar[10]),
    .I1(bbar[13])
  );
  //AND U176
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U176 (
    .O(y[172]),
    .I0(a[10]),
    .I1(b[12])
  );
  //OR U176bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U176bar (
    .O(ybar[172]),
    .I0(abar[10]),
    .I1(bbar[12])
  );
  //AND U177
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U177 (
    .O(y[171]),
    .I0(a[10]),
    .I1(b[11])
  );
  //OR U177bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U177bar (
    .O(ybar[171]),
    .I0(abar[10]),
    .I1(bbar[11])
  );
  //AND U178
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U178 (
    .O(y[170]),
    .I0(a[10]),
    .I1(b[10])
  );
  //OR U178bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U178bar (
    .O(ybar[170]),
    .I0(abar[10]),
    .I1(bbar[10])
  );
  //AND U179
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U179 (
    .O(y[16]),
    .I0(a[1]),
    .I1(b[0])
  );
  //OR U179bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U179bar (
    .O(ybar[16]),
    .I0(abar[1]),
    .I1(bbar[0])
  );
  //AND U180
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U180 (
    .O(y[169]),
    .I0(a[10]),
    .I1(b[9])
  );
  //OR U180bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U180bar (
    .O(ybar[169]),
    .I0(abar[10]),
    .I1(bbar[9])
  );
  //AND U181
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U181 (
    .O(y[168]),
    .I0(a[10]),
    .I1(b[8])
  );
  //OR U181bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U181bar (
    .O(ybar[168]),
    .I0(abar[10]),
    .I1(bbar[8])
  );
  //AND U182
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U182 (
    .O(y[167]),
    .I0(a[10]),
    .I1(b[7])
  );
  //OR U182bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U182bar (
    .O(ybar[167]),
    .I0(abar[10]),
    .I1(bbar[7])
  );
  //AND U183
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U183 (
    .O(y[166]),
    .I0(a[10]),
    .I1(b[6])
  );
  //OR U183bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U183bar (
    .O(ybar[166]),
    .I0(abar[10]),
    .I1(bbar[6])
  );
  //AND U184
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U184 (
    .O(y[165]),
    .I0(a[10]),
    .I1(b[5])
  );
  //OR U184bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U184bar (
    .O(ybar[165]),
    .I0(abar[10]),
    .I1(bbar[5])
  );
  //AND U185
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U185 (
    .O(y[164]),
    .I0(a[10]),
    .I1(b[4])
  );
  //OR U185bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U185bar (
    .O(ybar[164]),
    .I0(abar[10]),
    .I1(bbar[4])
  );
  //AND U186
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U186 (
    .O(y[163]),
    .I0(a[10]),
    .I1(b[3])
  );
  //OR U186bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U186bar (
    .O(ybar[163]),
    .I0(abar[10]),
    .I1(bbar[3])
  );
  //AND U187
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U187 (
    .O(y[162]),
    .I0(a[10]),
    .I1(b[2])
  );
  //OR U187bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U187bar (
    .O(ybar[162]),
    .I0(abar[10]),
    .I1(bbar[2])
  );
  //AND U188
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U188 (
    .O(y[161]),
    .I0(a[10]),
    .I1(b[1])
  );
  //OR U188bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U188bar (
    .O(ybar[161]),
    .I0(abar[10]),
    .I1(bbar[1])
  );
  //AND U189
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U189 (
    .O(y[160]),
    .I0(a[10]),
    .I1(b[0])
  );
  //OR U189bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U189bar (
    .O(ybar[160]),
    .I0(abar[10]),
    .I1(bbar[0])
  );
  //AND U190
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U190 (
    .O(y[15]),
    .I0(b[15]),
    .I1(a[0])
  );
  //OR U190bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U190bar (
    .O(ybar[15]),
    .I0(bbar[15]),
    .I1(abar[0])
  );
  //AND U191
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U191 (
    .O(y[159]),
    .I0(a[9]),
    .I1(b[15])
  );
  //OR U191bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U191bar (
    .O(ybar[159]),
    .I0(abar[9]),
    .I1(bbar[15])
  );
  //AND U192
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U192 (
    .O(y[158]),
    .I0(a[9]),
    .I1(b[14])
  );
  //OR U192bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U192bar (
    .O(ybar[158]),
    .I0(abar[9]),
    .I1(bbar[14])
  );
  //AND U193
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U193 (
    .O(y[157]),
    .I0(a[9]),
    .I1(b[13])
  );
  //OR U193bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U193bar (
    .O(ybar[157]),
    .I0(abar[9]),
    .I1(bbar[13])
  );
  //AND U194
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U194 (
    .O(y[156]),
    .I0(a[9]),
    .I1(b[12])
  );
  //OR U194bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U194bar (
    .O(ybar[156]),
    .I0(abar[9]),
    .I1(bbar[12])
  );
  //AND U195
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U195 (
    .O(y[155]),
    .I0(a[9]),
    .I1(b[11])
  );
  //OR U195bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U195bar (
    .O(ybar[155]),
    .I0(abar[9]),
    .I1(bbar[11])
  );
  //AND U196
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U196 (
    .O(y[154]),
    .I0(a[9]),
    .I1(b[10])
  );
  //OR U196bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U196bar (
    .O(ybar[154]),
    .I0(abar[9]),
    .I1(bbar[10])
  );
  //AND U197
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U197 (
    .O(y[153]),
    .I0(a[9]),
    .I1(b[9])
  );
  //OR U197bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U197bar (
    .O(ybar[153]),
    .I0(abar[9]),
    .I1(bbar[9])
  );
  //AND U198
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U198 (
    .O(y[152]),
    .I0(a[9]),
    .I1(b[8])
  );
  //OR U198bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U198bar (
    .O(ybar[152]),
    .I0(abar[9]),
    .I1(bbar[8])
  );
  //AND U199
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U199 (
    .O(y[151]),
    .I0(a[9]),
    .I1(b[7])
  );
  //OR U199bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U199bar (
    .O(ybar[151]),
    .I0(abar[9]),
    .I1(bbar[7])
  );
  //AND U200
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U200 (
    .O(y[150]),
    .I0(a[9]),
    .I1(b[6])
  );
  //OR U200bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U200bar (
    .O(ybar[150]),
    .I0(abar[9]),
    .I1(bbar[6])
  );
  //AND U201
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U201 (
    .O(y[14]),
    .I0(b[14]),
    .I1(a[0])
  );
  //OR U201bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U201bar (
    .O(ybar[14]),
    .I0(bbar[14]),
    .I1(abar[0])
  );
  //AND U202
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U202 (
    .O(y[149]),
    .I0(a[9]),
    .I1(b[5])
  );
  //OR U202bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U202bar (
    .O(ybar[149]),
    .I0(abar[9]),
    .I1(bbar[5])
  );
  //AND U203
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U203 (
    .O(y[148]),
    .I0(a[9]),
    .I1(b[4])
  );
  //OR U203bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U203bar (
    .O(ybar[148]),
    .I0(abar[9]),
    .I1(bbar[4])
  );
  //AND U204
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U204 (
    .O(y[147]),
    .I0(a[9]),
    .I1(b[3])
  );
  //OR U204bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U204bar (
    .O(ybar[147]),
    .I0(abar[9]),
    .I1(bbar[3])
  );
  //AND U205
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U205 (
    .O(y[146]),
    .I0(a[9]),
    .I1(b[2])
  );
  //OR U205bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U205bar (
    .O(ybar[146]),
    .I0(abar[9]),
    .I1(bbar[2])
  );
  //AND U206
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U206 (
    .O(y[145]),
    .I0(a[9]),
    .I1(b[1])
  );
  //OR U206bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U206bar (
    .O(ybar[145]),
    .I0(abar[9]),
    .I1(bbar[1])
  );
  //AND U207
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U207 (
    .O(y[144]),
    .I0(a[9]),
    .I1(b[0])
  );
  //OR U207bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U207bar (
    .O(ybar[144]),
    .I0(abar[9]),
    .I1(bbar[0])
  );
  //AND U208
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U208 (
    .O(y[143]),
    .I0(a[8]),
    .I1(b[15])
  );
  //OR U208bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U208bar (
    .O(ybar[143]),
    .I0(abar[8]),
    .I1(bbar[15])
  );
  //AND U209
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U209 (
    .O(y[142]),
    .I0(a[8]),
    .I1(b[14])
  );
  //OR U209bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U209bar (
    .O(ybar[142]),
    .I0(abar[8]),
    .I1(bbar[14])
  );
  //AND U210
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U210 (
    .O(y[141]),
    .I0(a[8]),
    .I1(b[13])
  );
  //OR U210bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U210bar (
    .O(ybar[141]),
    .I0(abar[8]),
    .I1(bbar[13])
  );
  //AND U211
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U211 (
    .O(y[140]),
    .I0(a[8]),
    .I1(b[12])
  );
  //OR U211bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U211bar (
    .O(ybar[140]),
    .I0(abar[8]),
    .I1(bbar[12])
  );
  //AND U212
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U212 (
    .O(y[13]),
    .I0(b[13]),
    .I1(a[0])
  );
  //OR U212bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U212bar (
    .O(ybar[13]),
    .I0(bbar[13]),
    .I1(abar[0])
  );
  //AND U213
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U213 (
    .O(y[139]),
    .I0(a[8]),
    .I1(b[11])
  );
  //OR U213bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U213bar (
    .O(ybar[139]),
    .I0(abar[8]),
    .I1(bbar[11])
  );
  //AND U214
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U214 (
    .O(y[138]),
    .I0(a[8]),
    .I1(b[10])
  );
  //OR U214bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U214bar (
    .O(ybar[138]),
    .I0(abar[8]),
    .I1(bbar[10])
  );
  //AND U215
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U215 (
    .O(y[137]),
    .I0(a[8]),
    .I1(b[9])
  );
  //OR U215bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U215bar (
    .O(ybar[137]),
    .I0(abar[8]),
    .I1(bbar[9])
  );
  //AND U216
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U216 (
    .O(y[136]),
    .I0(a[8]),
    .I1(b[8])
  );
  //OR U216bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U216bar (
    .O(ybar[136]),
    .I0(abar[8]),
    .I1(bbar[8])
  );
  //AND U217
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U217 (
    .O(y[135]),
    .I0(a[8]),
    .I1(b[7])
  );
  //OR U217bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U217bar (
    .O(ybar[135]),
    .I0(abar[8]),
    .I1(bbar[7])
  );
  //AND U218
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U218 (
    .O(y[134]),
    .I0(a[8]),
    .I1(b[6])
  );
  //OR U218bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U218bar (
    .O(ybar[134]),
    .I0(abar[8]),
    .I1(bbar[6])
  );
  //AND U219
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U219 (
    .O(y[133]),
    .I0(a[8]),
    .I1(b[5])
  );
  //OR U219bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U219bar (
    .O(ybar[133]),
    .I0(abar[8]),
    .I1(bbar[5])
  );
  //AND U220
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U220 (
    .O(y[132]),
    .I0(a[8]),
    .I1(b[4])
  );
  //OR U220bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U220bar (
    .O(ybar[132]),
    .I0(abar[8]),
    .I1(bbar[4])
  );
  //AND U221
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U221 (
    .O(y[131]),
    .I0(a[8]),
    .I1(b[3])
  );
  //OR U221bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U221bar (
    .O(ybar[131]),
    .I0(abar[8]),
    .I1(bbar[3])
  );
  //AND U222
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U222 (
    .O(y[130]),
    .I0(a[8]),
    .I1(b[2])
  );
  //OR U222bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U222bar (
    .O(ybar[130]),
    .I0(abar[8]),
    .I1(bbar[2])
  );
  //AND U223
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U223 (
    .O(y[12]),
    .I0(b[12]),
    .I1(a[0])
  );
  //OR U223bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U223bar (
    .O(ybar[12]),
    .I0(bbar[12]),
    .I1(abar[0])
  );
  //AND U224
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U224 (
    .O(y[129]),
    .I0(a[8]),
    .I1(b[1])
  );
  //OR U224bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U224bar (
    .O(ybar[129]),
    .I0(abar[8]),
    .I1(bbar[1])
  );
  //AND U225
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U225 (
    .O(y[128]),
    .I0(a[8]),
    .I1(b[0])
  );
  //OR U225bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U225bar (
    .O(ybar[128]),
    .I0(abar[8]),
    .I1(bbar[0])
  );
  //AND U226
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U226 (
    .O(y[127]),
    .I0(a[7]),
    .I1(b[15])
  );
  //OR U226bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U226bar (
    .O(ybar[127]),
    .I0(abar[7]),
    .I1(bbar[15])
  );
  //AND U227
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U227 (
    .O(y[126]),
    .I0(a[7]),
    .I1(b[14])
  );
  //OR U227bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U227bar (
    .O(ybar[126]),
    .I0(abar[7]),
    .I1(bbar[14])
  );
  //AND U228
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U228 (
    .O(y[125]),
    .I0(a[7]),
    .I1(b[13])
  );
  //OR U228bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U228bar (
    .O(ybar[125]),
    .I0(abar[7]),
    .I1(bbar[13])
  );
  //AND U229
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U229 (
    .O(y[124]),
    .I0(a[7]),
    .I1(b[12])
  );
  //OR U229bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U229bar (
    .O(ybar[124]),
    .I0(abar[7]),
    .I1(bbar[12])
  );
  //AND U230
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U230 (
    .O(y[123]),
    .I0(a[7]),
    .I1(b[11])
  );
  //OR U230bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U230bar (
    .O(ybar[123]),
    .I0(abar[7]),
    .I1(bbar[11])
  );
  //AND U231
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U231 (
    .O(y[122]),
    .I0(a[7]),
    .I1(b[10])
  );
  //OR U231bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U231bar (
    .O(ybar[122]),
    .I0(abar[7]),
    .I1(bbar[10])
  );
  //AND U232
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U232 (
    .O(y[121]),
    .I0(a[7]),
    .I1(b[9])
  );
  //OR U232bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U232bar (
    .O(ybar[121]),
    .I0(abar[7]),
    .I1(bbar[9])
  );
  //AND U233
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U233 (
    .O(y[120]),
    .I0(a[7]),
    .I1(b[8])
  );
  //OR U233bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U233bar (
    .O(ybar[120]),
    .I0(abar[7]),
    .I1(bbar[8])
  );
  //AND U234
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U234 (
    .O(y[11]),
    .I0(b[11]),
    .I1(a[0])
  );
  //OR U234bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U234bar (
    .O(ybar[11]),
    .I0(bbar[11]),
    .I1(abar[0])
  );
  //AND U235
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U235 (
    .O(y[119]),
    .I0(a[7]),
    .I1(b[7])
  );
  //OR U235bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U235bar (
    .O(ybar[119]),
    .I0(abar[7]),
    .I1(bbar[7])
  );
  //AND U236
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U236 (
    .O(y[118]),
    .I0(a[7]),
    .I1(b[6])
  );
  //OR U236bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U236bar (
    .O(ybar[118]),
    .I0(abar[7]),
    .I1(bbar[6])
  );
  //AND U237
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U237 (
    .O(y[117]),
    .I0(a[7]),
    .I1(b[5])
  );
  //OR U237bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U237bar (
    .O(ybar[117]),
    .I0(abar[7]),
    .I1(bbar[5])
  );
  //AND U238
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U238 (
    .O(y[116]),
    .I0(a[7]),
    .I1(b[4])
  );
  //OR U238bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U238bar (
    .O(ybar[116]),
    .I0(abar[7]),
    .I1(bbar[4])
  );
  //AND U239
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U239 (
    .O(y[115]),
    .I0(a[7]),
    .I1(b[3])
  );
  //OR U239bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U239bar (
    .O(ybar[115]),
    .I0(abar[7]),
    .I1(bbar[3])
  );
  //AND U240
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U240 (
    .O(y[114]),
    .I0(a[7]),
    .I1(b[2])
  );
  //OR U240bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U240bar (
    .O(ybar[114]),
    .I0(abar[7]),
    .I1(bbar[2])
  );
  //AND U241
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U241 (
    .O(y[113]),
    .I0(a[7]),
    .I1(b[1])
  );
  //OR U241bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U241bar (
    .O(ybar[113]),
    .I0(abar[7]),
    .I1(bbar[1])
  );
  //AND U242
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U242 (
    .O(y[112]),
    .I0(a[7]),
    .I1(b[0])
  );
  //OR U242bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U242bar (
    .O(ybar[112]),
    .I0(abar[7]),
    .I1(bbar[0])
  );
  //AND U243
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U243 (
    .O(y[111]),
    .I0(b[15]),
    .I1(a[6])
  );
  //OR U243bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U243bar (
    .O(ybar[111]),
    .I0(bbar[15]),
    .I1(abar[6])
  );
  //AND U244
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U244 (
    .O(y[110]),
    .I0(b[14]),
    .I1(a[6])
  );
  //OR U244bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U244bar (
    .O(ybar[110]),
    .I0(bbar[14]),
    .I1(abar[6])
  );
  //AND U245
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U245 (
    .O(y[10]),
    .I0(b[10]),
    .I1(a[0])
  );
  //OR U245bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U245bar (
    .O(ybar[10]),
    .I0(bbar[10]),
    .I1(abar[0])
  );
  //AND U246
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U246 (
    .O(y[109]),
    .I0(b[13]),
    .I1(a[6])
  );
  //OR U246bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U246bar (
    .O(ybar[109]),
    .I0(bbar[13]),
    .I1(abar[6])
  );
  //AND U247
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U247 (
    .O(y[108]),
    .I0(b[12]),
    .I1(a[6])
  );
  //OR U247bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U247bar (
    .O(ybar[108]),
    .I0(bbar[12]),
    .I1(abar[6])
  );
  //AND U248
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U248 (
    .O(y[107]),
    .I0(b[11]),
    .I1(a[6])
  );
  //OR U248bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U248bar (
    .O(ybar[107]),
    .I0(bbar[11]),
    .I1(abar[6])
  );
  //AND U249
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U249 (
    .O(y[106]),
    .I0(b[10]),
    .I1(a[6])
  );
  //OR U249bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U249bar (
    .O(ybar[106]),
    .I0(bbar[10]),
    .I1(abar[6])
  );
  //AND U250
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U250 (
    .O(y[105]),
    .I0(a[6]),
    .I1(b[9])
  );
  //OR U250bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U250bar (
    .O(ybar[105]),
    .I0(abar[6]),
    .I1(bbar[9])
  );
  //AND U251
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U251 (
    .O(y[104]),
    .I0(b[8]),
    .I1(a[6])
  );
  //OR U251bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U251bar (
    .O(ybar[104]),
    .I0(bbar[8]),
    .I1(abar[6])
  );
  //AND U252
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U252 (
    .O(y[103]),
    .I0(b[7]),
    .I1(a[6])
  );
  //OR U252bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U252bar (
    .O(ybar[103]),
    .I0(bbar[7]),
    .I1(abar[6])
  );
  //AND U253
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U253 (
    .O(y[102]),
    .I0(b[6]),
    .I1(a[6])
  );
  //OR U253bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U253bar (
    .O(ybar[102]),
    .I0(bbar[6]),
    .I1(abar[6])
  );
  //AND U254
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U254 (
    .O(y[101]),
    .I0(b[5]),
    .I1(a[6])
  );
  //OR U254bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U254bar (
    .O(ybar[101]),
    .I0(bbar[5]),
    .I1(abar[6])
  );
  //AND U255
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U255 (
    .O(y[100]),
    .I0(b[4]),
    .I1(a[6])
  );
  //OR U255bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U255bar (
    .O(ybar[100]),
    .I0(bbar[4]),
    .I1(abar[6])
  );
  //AND U256
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U256 (
    .O(y[0]),
    .I0(b[0]),
    .I1(a[0])
  );
  //OR U256bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U256bar (
    .O(ybar[0]),
    .I0(bbar[0]),
    .I1(abar[0])
  );
endmodule

module CD2_77 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD2_78 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD2_79 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD4_39 ( a, b, y );

  input wire [3:0] a;
  input wire [3:0] b;
  wire [3:0] abar;
  wire [3:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
//input_done

  output wire [15:0] y;
  wire [15:0] ybar;
//output_done

//wire_done

  //AND U1
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1 (
    .O(y[9]),
    .I0(b[1]),
    .I1(a[2])
  );
  //OR U1bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1bar (
    .O(ybar[9]),
    .I0(bbar[1]),
    .I1(abar[2])
  );
  //AND U2
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2 (
    .O(y[8]),
    .I0(b[0]),
    .I1(a[2])
  );
  //OR U2bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2bar (
    .O(ybar[8]),
    .I0(bbar[0]),
    .I1(abar[2])
  );
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[7]),
    .I0(b[3]),
    .I1(a[1])
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[7]),
    .I0(bbar[3]),
    .I1(abar[1])
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[6]),
    .I0(b[2]),
    .I1(a[1])
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[6]),
    .I0(bbar[2]),
    .I1(abar[1])
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[5]),
    .I0(a[1]),
    .I1(b[1])
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[5]),
    .I0(abar[1]),
    .I1(bbar[1])
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[4]),
    .I0(a[1]),
    .I1(b[0])
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[4]),
    .I0(abar[1]),
    .I1(bbar[0])
  );
  //AND U7
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7 (
    .O(y[3]),
    .I0(a[0]),
    .I1(b[3])
  );
  //OR U7bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7bar (
    .O(ybar[3]),
    .I0(abar[0]),
    .I1(bbar[3])
  );
  //AND U8
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8 (
    .O(y[2]),
    .I0(a[0]),
    .I1(b[2])
  );
  //OR U8bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8bar (
    .O(ybar[2]),
    .I0(abar[0]),
    .I1(bbar[2])
  );
  //AND U9
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9 (
    .O(y[1]),
    .I0(a[0]),
    .I1(b[1])
  );
  //OR U9bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9bar (
    .O(ybar[1]),
    .I0(abar[0]),
    .I1(bbar[1])
  );
  //AND U10
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10 (
    .O(y[15]),
    .I0(a[3]),
    .I1(b[3])
  );
  //OR U10bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10bar (
    .O(ybar[15]),
    .I0(abar[3]),
    .I1(bbar[3])
  );
  //AND U11
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11 (
    .O(y[14]),
    .I0(a[3]),
    .I1(b[2])
  );
  //OR U11bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11bar (
    .O(ybar[14]),
    .I0(abar[3]),
    .I1(bbar[2])
  );
  //AND U12
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12 (
    .O(y[13]),
    .I0(a[3]),
    .I1(b[1])
  );
  //OR U12bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12bar (
    .O(ybar[13]),
    .I0(abar[3]),
    .I1(bbar[1])
  );
  //AND U13
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13 (
    .O(y[12]),
    .I0(a[3]),
    .I1(b[0])
  );
  //OR U13bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13bar (
    .O(ybar[12]),
    .I0(abar[3]),
    .I1(bbar[0])
  );
  //AND U14
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14 (
    .O(y[11]),
    .I0(b[3]),
    .I1(a[2])
  );
  //OR U14bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14bar (
    .O(ybar[11]),
    .I0(bbar[3]),
    .I1(abar[2])
  );
  //AND U15
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15 (
    .O(y[10]),
    .I0(b[2]),
    .I1(a[2])
  );
  //OR U15bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15bar (
    .O(ybar[10]),
    .I0(bbar[2]),
    .I1(abar[2])
  );
  //AND U16
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16 (
    .O(y[0]),
    .I0(a[0]),
    .I1(b[0])
  );
  //OR U16bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16bar (
    .O(ybar[0]),
    .I0(abar[0]),
    .I1(bbar[0])
  );
endmodule

module decode_0 ( in, out );

  input wire [7:0] in;
//input_done

  output wire [255:0] out;
//output_done

  wire [15:0] level1;
  wire [31:0] level2;
//wire_done

  CD2_0 cd_l1_1 ( .a(in[1]), .b(in[0]), .y(level1[3:0]) );
  CD2_79 cd_l1_2 ( .a(in[3]), .b(in[2]), .y(level1[7:4]) );
  CD2_78 cd_l1_3 ( .a(in[5]), .b(in[4]), .y(level1[11:8]) );
  CD2_77 cd_l1_4 ( .a(in[7]), .b(in[6]), .y(level1[15:12]) );
  CD4_0 cd_l2_1 ( .a(level1[7:4]), .b(level1[3:0]), .y(level2[15:0]) );
  CD4_39 cd_l2_2 ( .a(level1[15:12]), .b(level1[11:8]), .y(level2[31:16]) );
  CD16_0 cd_l3 ( .a(level2[31:16]), .b(level2[15:0]), .y(out) );
endmodule

module encode_0 ( in, out );

  input wire [255:0] in;
  wire [255:0] inbar;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
  assign inbar[8] = ~in[8];
  assign inbar[9] = ~in[9];
  assign inbar[10] = ~in[10];
  assign inbar[11] = ~in[11];
  assign inbar[12] = ~in[12];
  assign inbar[13] = ~in[13];
  assign inbar[14] = ~in[14];
  assign inbar[15] = ~in[15];
  assign inbar[16] = ~in[16];
  assign inbar[17] = ~in[17];
  assign inbar[18] = ~in[18];
  assign inbar[19] = ~in[19];
  assign inbar[20] = ~in[20];
  assign inbar[21] = ~in[21];
  assign inbar[22] = ~in[22];
  assign inbar[23] = ~in[23];
  assign inbar[24] = ~in[24];
  assign inbar[25] = ~in[25];
  assign inbar[26] = ~in[26];
  assign inbar[27] = ~in[27];
  assign inbar[28] = ~in[28];
  assign inbar[29] = ~in[29];
  assign inbar[30] = ~in[30];
  assign inbar[31] = ~in[31];
  assign inbar[32] = ~in[32];
  assign inbar[33] = ~in[33];
  assign inbar[34] = ~in[34];
  assign inbar[35] = ~in[35];
  assign inbar[36] = ~in[36];
  assign inbar[37] = ~in[37];
  assign inbar[38] = ~in[38];
  assign inbar[39] = ~in[39];
  assign inbar[40] = ~in[40];
  assign inbar[41] = ~in[41];
  assign inbar[42] = ~in[42];
  assign inbar[43] = ~in[43];
  assign inbar[44] = ~in[44];
  assign inbar[45] = ~in[45];
  assign inbar[46] = ~in[46];
  assign inbar[47] = ~in[47];
  assign inbar[48] = ~in[48];
  assign inbar[49] = ~in[49];
  assign inbar[50] = ~in[50];
  assign inbar[51] = ~in[51];
  assign inbar[52] = ~in[52];
  assign inbar[53] = ~in[53];
  assign inbar[54] = ~in[54];
  assign inbar[55] = ~in[55];
  assign inbar[56] = ~in[56];
  assign inbar[57] = ~in[57];
  assign inbar[58] = ~in[58];
  assign inbar[59] = ~in[59];
  assign inbar[60] = ~in[60];
  assign inbar[61] = ~in[61];
  assign inbar[62] = ~in[62];
  assign inbar[63] = ~in[63];
  assign inbar[64] = ~in[64];
  assign inbar[65] = ~in[65];
  assign inbar[66] = ~in[66];
  assign inbar[67] = ~in[67];
  assign inbar[68] = ~in[68];
  assign inbar[69] = ~in[69];
  assign inbar[70] = ~in[70];
  assign inbar[71] = ~in[71];
  assign inbar[72] = ~in[72];
  assign inbar[73] = ~in[73];
  assign inbar[74] = ~in[74];
  assign inbar[75] = ~in[75];
  assign inbar[76] = ~in[76];
  assign inbar[77] = ~in[77];
  assign inbar[78] = ~in[78];
  assign inbar[79] = ~in[79];
  assign inbar[80] = ~in[80];
  assign inbar[81] = ~in[81];
  assign inbar[82] = ~in[82];
  assign inbar[83] = ~in[83];
  assign inbar[84] = ~in[84];
  assign inbar[85] = ~in[85];
  assign inbar[86] = ~in[86];
  assign inbar[87] = ~in[87];
  assign inbar[88] = ~in[88];
  assign inbar[89] = ~in[89];
  assign inbar[90] = ~in[90];
  assign inbar[91] = ~in[91];
  assign inbar[92] = ~in[92];
  assign inbar[93] = ~in[93];
  assign inbar[94] = ~in[94];
  assign inbar[95] = ~in[95];
  assign inbar[96] = ~in[96];
  assign inbar[97] = ~in[97];
  assign inbar[98] = ~in[98];
  assign inbar[99] = ~in[99];
  assign inbar[100] = ~in[100];
  assign inbar[101] = ~in[101];
  assign inbar[102] = ~in[102];
  assign inbar[103] = ~in[103];
  assign inbar[104] = ~in[104];
  assign inbar[105] = ~in[105];
  assign inbar[106] = ~in[106];
  assign inbar[107] = ~in[107];
  assign inbar[108] = ~in[108];
  assign inbar[109] = ~in[109];
  assign inbar[110] = ~in[110];
  assign inbar[111] = ~in[111];
  assign inbar[112] = ~in[112];
  assign inbar[113] = ~in[113];
  assign inbar[114] = ~in[114];
  assign inbar[115] = ~in[115];
  assign inbar[116] = ~in[116];
  assign inbar[117] = ~in[117];
  assign inbar[118] = ~in[118];
  assign inbar[119] = ~in[119];
  assign inbar[120] = ~in[120];
  assign inbar[121] = ~in[121];
  assign inbar[122] = ~in[122];
  assign inbar[123] = ~in[123];
  assign inbar[124] = ~in[124];
  assign inbar[125] = ~in[125];
  assign inbar[126] = ~in[126];
  assign inbar[127] = ~in[127];
  assign inbar[128] = ~in[128];
  assign inbar[129] = ~in[129];
  assign inbar[130] = ~in[130];
  assign inbar[131] = ~in[131];
  assign inbar[132] = ~in[132];
  assign inbar[133] = ~in[133];
  assign inbar[134] = ~in[134];
  assign inbar[135] = ~in[135];
  assign inbar[136] = ~in[136];
  assign inbar[137] = ~in[137];
  assign inbar[138] = ~in[138];
  assign inbar[139] = ~in[139];
  assign inbar[140] = ~in[140];
  assign inbar[141] = ~in[141];
  assign inbar[142] = ~in[142];
  assign inbar[143] = ~in[143];
  assign inbar[144] = ~in[144];
  assign inbar[145] = ~in[145];
  assign inbar[146] = ~in[146];
  assign inbar[147] = ~in[147];
  assign inbar[148] = ~in[148];
  assign inbar[149] = ~in[149];
  assign inbar[150] = ~in[150];
  assign inbar[151] = ~in[151];
  assign inbar[152] = ~in[152];
  assign inbar[153] = ~in[153];
  assign inbar[154] = ~in[154];
  assign inbar[155] = ~in[155];
  assign inbar[156] = ~in[156];
  assign inbar[157] = ~in[157];
  assign inbar[158] = ~in[158];
  assign inbar[159] = ~in[159];
  assign inbar[160] = ~in[160];
  assign inbar[161] = ~in[161];
  assign inbar[162] = ~in[162];
  assign inbar[163] = ~in[163];
  assign inbar[164] = ~in[164];
  assign inbar[165] = ~in[165];
  assign inbar[166] = ~in[166];
  assign inbar[167] = ~in[167];
  assign inbar[168] = ~in[168];
  assign inbar[169] = ~in[169];
  assign inbar[170] = ~in[170];
  assign inbar[171] = ~in[171];
  assign inbar[172] = ~in[172];
  assign inbar[173] = ~in[173];
  assign inbar[174] = ~in[174];
  assign inbar[175] = ~in[175];
  assign inbar[176] = ~in[176];
  assign inbar[177] = ~in[177];
  assign inbar[178] = ~in[178];
  assign inbar[179] = ~in[179];
  assign inbar[180] = ~in[180];
  assign inbar[181] = ~in[181];
  assign inbar[182] = ~in[182];
  assign inbar[183] = ~in[183];
  assign inbar[184] = ~in[184];
  assign inbar[185] = ~in[185];
  assign inbar[186] = ~in[186];
  assign inbar[187] = ~in[187];
  assign inbar[188] = ~in[188];
  assign inbar[189] = ~in[189];
  assign inbar[190] = ~in[190];
  assign inbar[191] = ~in[191];
  assign inbar[192] = ~in[192];
  assign inbar[193] = ~in[193];
  assign inbar[194] = ~in[194];
  assign inbar[195] = ~in[195];
  assign inbar[196] = ~in[196];
  assign inbar[197] = ~in[197];
  assign inbar[198] = ~in[198];
  assign inbar[199] = ~in[199];
  assign inbar[200] = ~in[200];
  assign inbar[201] = ~in[201];
  assign inbar[202] = ~in[202];
  assign inbar[203] = ~in[203];
  assign inbar[204] = ~in[204];
  assign inbar[205] = ~in[205];
  assign inbar[206] = ~in[206];
  assign inbar[207] = ~in[207];
  assign inbar[208] = ~in[208];
  assign inbar[209] = ~in[209];
  assign inbar[210] = ~in[210];
  assign inbar[211] = ~in[211];
  assign inbar[212] = ~in[212];
  assign inbar[213] = ~in[213];
  assign inbar[214] = ~in[214];
  assign inbar[215] = ~in[215];
  assign inbar[216] = ~in[216];
  assign inbar[217] = ~in[217];
  assign inbar[218] = ~in[218];
  assign inbar[219] = ~in[219];
  assign inbar[220] = ~in[220];
  assign inbar[221] = ~in[221];
  assign inbar[222] = ~in[222];
  assign inbar[223] = ~in[223];
  assign inbar[224] = ~in[224];
  assign inbar[225] = ~in[225];
  assign inbar[226] = ~in[226];
  assign inbar[227] = ~in[227];
  assign inbar[228] = ~in[228];
  assign inbar[229] = ~in[229];
  assign inbar[230] = ~in[230];
  assign inbar[231] = ~in[231];
  assign inbar[232] = ~in[232];
  assign inbar[233] = ~in[233];
  assign inbar[234] = ~in[234];
  assign inbar[235] = ~in[235];
  assign inbar[236] = ~in[236];
  assign inbar[237] = ~in[237];
  assign inbar[238] = ~in[238];
  assign inbar[239] = ~in[239];
  assign inbar[240] = ~in[240];
  assign inbar[241] = ~in[241];
  assign inbar[242] = ~in[242];
  assign inbar[243] = ~in[243];
  assign inbar[244] = ~in[244];
  assign inbar[245] = ~in[245];
  assign inbar[246] = ~in[246];
  assign inbar[247] = ~in[247];
  assign inbar[248] = ~in[248];
  assign inbar[249] = ~in[249];
  assign inbar[250] = ~in[250];
  assign inbar[251] = ~in[251];
  assign inbar[252] = ~in[252];
  assign inbar[253] = ~in[253];
  assign inbar[254] = ~in[254];
  assign inbar[255] = ~in[255];
//input_done

  output wire [7:0] out;
  wire [7:0] outbar;
//output_done

  wire in_81;
  wire in_80;
  wire in_79;
  wire in_78;
  wire in_77;
  wire in_76;
  wire in_75;
  wire in_74;
  wire in_73;
  wire in_72;
  wire in_71;
  wire in_70;
  wire in_69;
  wire in_68;
  wire in_67;
  wire in_66;
  wire in_65;
  wire in_64;
  wire in_63;
  wire in_62;
  wire in_61;
  wire in_60;
  wire in_59;
  wire in_58;
  wire in_57;
  wire in_56;
  wire in_55;
  wire in_54;
  wire in_53;
  wire in_52;
  wire in_51;
  wire in_50;
  wire in_49;
  wire in_48;
  wire in_47;
  wire in_46;
  wire in_45;
  wire in_44;
  wire in_43;
  wire in_42;
  wire in_41;
  wire in_40;
  wire in_39;
  wire in_38;
  wire in_37;
  wire in_36;
  wire in_35;
  wire in_34;
  wire in_33;
  wire in_32;
  wire in_31;
  wire in_30;
  wire in_29;
  wire in_28;
  wire in_27;
  wire in_26;
  wire in_25;
  wire in_24;
  wire in_23;
  wire in_22;
  wire in_21;
  wire in_20;
  wire in_19;
  wire in_18;
  wire in_17;
  wire in_16;
  wire in_15;
  wire in_14;
  wire in_13;
  wire in_12;
  wire in_11;
  wire in_10;
  wire in_9;
  wire in_8;
  wire in_7;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_3;
  wire in_2;
  wire in_1;
  wire in_0;
  wire n1;
  wire n2;
  wire n3;
  wire n4;
  wire n5;
  wire n6;
  wire n7;
  wire n8;
  wire n9;
  wire n10;
  wire n11;
  wire n12;
  wire n13;
  wire n14;
  wire n15;
  wire n16;
  wire n17;
  wire n18;
  wire n19;
  wire n20;
  wire n21;
  wire n22;
  wire n23;
  wire n24;
  wire n25;
  wire n26;
  wire n27;
  wire n28;
  wire n29;
  wire n30;
  wire n31;
  wire n32;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire in_81bar;
  wire in_80bar;
  wire in_79bar;
  wire in_78bar;
  wire in_77bar;
  wire in_76bar;
  wire in_75bar;
  wire in_74bar;
  wire in_73bar;
  wire in_72bar;
  wire in_71bar;
  wire in_70bar;
  wire in_69bar;
  wire in_68bar;
  wire in_67bar;
  wire in_66bar;
  wire in_65bar;
  wire in_64bar;
  wire in_63bar;
  wire in_62bar;
  wire in_61bar;
  wire in_60bar;
  wire in_59bar;
  wire in_58bar;
  wire in_57bar;
  wire in_56bar;
  wire in_55bar;
  wire in_54bar;
  wire in_53bar;
  wire in_52bar;
  wire in_51bar;
  wire in_50bar;
  wire in_49bar;
  wire in_48bar;
  wire in_47bar;
  wire in_46bar;
  wire in_45bar;
  wire in_44bar;
  wire in_43bar;
  wire in_42bar;
  wire in_41bar;
  wire in_40bar;
  wire in_39bar;
  wire in_38bar;
  wire in_37bar;
  wire in_36bar;
  wire in_35bar;
  wire in_34bar;
  wire in_33bar;
  wire in_32bar;
  wire in_31bar;
  wire in_30bar;
  wire in_29bar;
  wire in_28bar;
  wire in_27bar;
  wire in_26bar;
  wire in_25bar;
  wire in_24bar;
  wire in_23bar;
  wire in_22bar;
  wire in_21bar;
  wire in_20bar;
  wire in_19bar;
  wire in_18bar;
  wire in_17bar;
  wire in_16bar;
  wire in_15bar;
  wire in_14bar;
  wire in_13bar;
  wire in_12bar;
  wire in_11bar;
  wire in_10bar;
  wire in_9bar;
  wire in_8bar;
  wire in_7bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_3bar;
  wire in_2bar;
  wire in_1bar;
  wire in_0bar;
  wire n1bar;
  wire n2bar;
  wire n3bar;
  wire n4bar;
  wire n5bar;
  wire n6bar;
  wire n7bar;
  wire n8bar;
  wire n9bar;
  wire n10bar;
  wire n11bar;
  wire n12bar;
  wire n13bar;
  wire n14bar;
  wire n15bar;
  wire n16bar;
  wire n17bar;
  wire n18bar;
  wire n19bar;
  wire n20bar;
  wire n21bar;
  wire n22bar;
  wire n23bar;
  wire n24bar;
  wire n25bar;
  wire n26bar;
  wire n27bar;
  wire n28bar;
  wire n29bar;
  wire n30bar;
  wire n31bar;
  wire n32bar;
  wire n33bar;
  wire n34bar;
  wire n35bar;
  wire n36bar;
  wire n37bar;
  wire n38bar;
  wire n39bar;
  wire n40bar;
  wire n41bar;
  wire n42bar;
  wire n43bar;
  wire n44bar;
  wire n45bar;
  wire n46bar;
  wire n47bar;
  wire n48bar;
  wire n49bar;
  wire n50bar;
  wire n51bar;
  wire n52bar;
  wire n53bar;
  wire n54bar;
  wire n55bar;
  wire n56bar;
  wire n57bar;
  wire n58bar;
  wire n59bar;
  wire n60bar;
  wire n61bar;
  wire n62bar;
  wire n63bar;
  wire n64bar;
  wire n65bar;
  wire n66bar;
  wire n67bar;
  wire n68bar;
  wire n69bar;
  wire n70bar;
  wire n71bar;
  wire n72bar;
  wire n73bar;
  wire n74bar;
  wire n75bar;
  wire n76bar;
  wire n77bar;
  wire n78bar;
  wire n79bar;
  wire n80bar;
  wire n81bar;
  wire n82bar;
  wire n83bar;
  wire n84bar;
  wire n85bar;
  wire n86bar;
  wire n87bar;
  wire n88bar;
  wire n89bar;
  wire n90bar;
  wire n91bar;
  wire n92bar;
  wire n93bar;
  wire n94bar;
  wire n95bar;
  wire n96bar;
  wire n97bar;
  wire n98bar;
  wire n99bar;
  wire n100bar;
  wire n101bar;
  wire n102bar;
  wire n103bar;
  wire n104bar;
  wire n105bar;
  wire n106bar;
  wire n107bar;
  wire n108bar;
  wire n109bar;
  wire n110bar;
  wire n111bar;
  wire n112bar;
  wire n113bar;
  wire n114bar;
  wire n115bar;
  wire n116bar;
  wire n117bar;
  wire n118bar;
  wire n119bar;
  wire n120bar;
  wire n121bar;
  wire n122bar;
  wire n123bar;
  wire n124bar;
  wire n125bar;
  wire n126bar;
  wire n127bar;
  wire n128bar;
  wire n129bar;
  wire n130bar;
  wire n131bar;
  wire n132bar;
  wire n133bar;
  wire n134bar;
  wire n135bar;
  wire n136bar;
  wire n137bar;
  wire n138bar;
  wire n139bar;
  wire n140bar;
  wire n141bar;
  wire n142bar;
  wire n143bar;
  wire n144bar;
  wire n145bar;
  wire n146bar;
  wire n147bar;
  wire n148bar;
  wire n149bar;
  wire n150bar;
  wire n151bar;
  wire n152bar;
  wire n153bar;
  wire n154bar;
  wire n155bar;
  wire n156bar;
  wire n157bar;
  wire n158bar;
  wire n159bar;
  wire n160bar;
  wire n161bar;
  wire n162bar;
  wire n163bar;
  wire n164bar;
  wire n165bar;
  wire n166bar;
  wire n167bar;
  wire n168bar;
  wire n169bar;
  wire n170bar;
  wire n171bar;
  wire n172bar;
  wire n173bar;
  wire n174bar;
  wire n175bar;
  wire n176bar;
  wire n177bar;
  wire n178bar;
  wire n179bar;
  wire n180bar;
  wire n181bar;
  wire n182bar;
  wire n183bar;
  wire n184bar;
  wire n185bar;
  wire n186bar;
  wire n187bar;
  wire n188bar;
  wire n189bar;
  wire n190bar;
  wire n191bar;
  wire n192bar;
  wire n193bar;
  wire n194bar;
  wire n195bar;
  wire n196bar;
  wire n197bar;
  wire n198bar;
  wire n199bar;
  wire n200bar;
  wire n201bar;
  wire n202bar;
  wire n203bar;
  wire n204bar;
  wire n205bar;
  wire n206bar;
  wire n207bar;
  wire n208bar;
  wire n209bar;
  wire n210bar;
  wire n211bar;
  wire n212bar;
  wire n213bar;
  wire n214bar;
  wire n215bar;
  wire n216bar;
  wire n217bar;
  wire n218bar;
  wire n219bar;
  wire n220bar;
  wire n221bar;
  wire n222bar;
  wire n223bar;
  wire n224bar;
  wire n225bar;
  wire n226bar;
  wire n227bar;
  wire n228bar;
  wire n229bar;
  wire n230bar;
  wire n231bar;
  wire n232bar;
  wire n233bar;
  wire n234bar;
  wire n235bar;
  wire n236bar;
  wire n237bar;
  wire n238bar;
  wire n239bar;
  wire n240bar;
  wire n241bar;
  wire n242bar;
  wire n243bar;
  wire n244bar;
  wire n245bar;
  wire n246bar;
  wire n247bar;
  wire n248bar;
  wire n249bar;
  wire n250bar;
  wire n251bar;
  wire n252bar;
  wire n253bar;
  wire n254bar;
  wire n255bar;
  wire n256bar;
  wire n257bar;
  wire n258bar;
  wire n259bar;
  wire n260bar;
  wire n261bar;
  wire n262bar;
  wire n263bar;
  wire n264bar;
  wire n265bar;
  wire n266bar;
  wire n267bar;
  wire n268bar;
  wire n269bar;
  wire n270bar;
  wire n271bar;
  wire n272bar;
  wire n273bar;
  wire n274bar;
  wire n275bar;
  wire n276bar;
  wire n277bar;
  wire n278bar;
  wire n279bar;
  wire n280bar;
  wire n281bar;
  wire n282bar;
  wire n283bar;
  wire n284bar;
  wire n285bar;
  wire n286bar;
  wire n287bar;
  wire n288bar;
  wire n289bar;
  wire n290bar;
  wire n291bar;
  wire n292bar;
  wire n293bar;
  wire n294bar;
  wire n295bar;
  wire n296bar;
  wire n297bar;
  wire n298bar;
  wire n299bar;
  wire n300bar;
  wire n301bar;
  wire n302bar;
  wire n303bar;
  wire n304bar;
  wire n305bar;
  wire n306bar;
  wire n307bar;
  wire n308bar;
  wire n309bar;
  wire n310bar;
  wire n311bar;
  wire n312bar;
  wire n313bar;
  wire n314bar;
  wire n315bar;
  wire n316bar;
  wire n317bar;
  wire n318bar;
  wire n319bar;
  wire n320bar;
  wire n321bar;
  wire n322bar;
  wire n323bar;
  wire n324bar;
  wire n325bar;
  wire n326bar;
  wire n327bar;
  wire n328bar;
  wire n329bar;
  wire n330bar;
  wire n331bar;
  wire n332bar;
  wire n333bar;
  wire n334bar;
  wire n335bar;
  wire n336bar;
  wire n337bar;
  wire n338bar;
  wire n339bar;
  wire n340bar;
  wire n341bar;
  wire n342bar;
  wire n343bar;
  wire n344bar;
  wire n345bar;
  wire n346bar;
  wire n347bar;
  wire n348bar;
  wire n349bar;
  wire n350bar;
  wire n351bar;
  wire n352bar;
  wire n353bar;
  wire n354bar;
  wire n355bar;
  wire n356bar;
  wire n357bar;
  wire n358bar;
  wire n359bar;
  wire n360bar;
  wire n361bar;
  wire n362bar;
  wire n363bar;
  wire n364bar;
  wire n365bar;
  wire n366bar;
  wire n367bar;
  wire n368bar;
  wire n369bar;
  wire n370bar;
  wire n371bar;
  wire n372bar;
  wire n373bar;
  wire n374bar;
  wire n375bar;
  wire n376bar;
  wire n377bar;
  wire n378bar;
  wire n379bar;
  wire n380bar;
  wire n381bar;
  wire n382bar;
  wire n383bar;
  wire n384bar;
  wire n385bar;
  wire n386bar;
  wire n387bar;
  wire n388bar;
  wire n389bar;
  wire n390bar;
  wire n391bar;
  wire n392bar;
  wire n393bar;
  wire n394bar;
  wire n395bar;
  wire n396bar;
  wire n397bar;
  wire n398bar;
  wire n399bar;
  wire n400bar;
  wire n401bar;
  wire n402bar;
  wire n403bar;
  wire n404bar;
  wire n405bar;
  wire n406bar;
  wire n407bar;
  wire n408bar;
  wire n409bar;
  wire n410bar;
  wire n411bar;
  wire n412bar;
  wire n413bar;
  wire n414bar;
  wire n415bar;
  wire n416bar;
  wire n417bar;
  wire n418bar;
  wire n419bar;
  wire n420bar;
  wire n421bar;
  wire n422bar;
  wire n423bar;
  wire n424bar;
  wire n425bar;
  wire n426bar;
  wire n427bar;
  wire n428bar;
  wire n429bar;
  wire n430bar;
  wire n431bar;
  wire n432bar;
  wire n433bar;
  wire n434bar;
  wire n435bar;
  wire n436bar;
  wire n437bar;
  wire n438bar;
  wire n439bar;
  wire n440bar;
  wire n441bar;
  wire n442bar;
  wire n443bar;
  wire n444bar;
  wire n445bar;
  wire n446bar;
  wire n447bar;
  wire n448bar;
  wire n449bar;
  wire n450bar;
  wire n451bar;
  wire n452bar;
  wire n453bar;
  wire n454bar;
  wire n455bar;
  wire n456bar;
  wire n457bar;
  wire n458bar;
  wire n459bar;
  wire n460bar;
  wire n461bar;
  wire n462bar;
  wire n463bar;
  wire n464bar;
  wire n465bar;
  wire n466bar;
  wire n467bar;
  wire n468bar;
  wire n469bar;
  wire n470bar;
  wire n471bar;
  wire n472bar;
  wire n473bar;
  wire n474bar;
  wire n475bar;
  wire n476bar;
  wire n477bar;
  wire n478bar;
  wire n479bar;
  wire n480bar;
  wire n481bar;
  wire n482bar;
  wire n483bar;
  wire n484bar;
  wire n485bar;
  wire n486bar;
//wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];
  //OR U1
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1 (
    .O(out[7]),
    .I0(n1),
    .I1(n2)
  );
  //AND U1bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1bar (
    .O(outbar[7]),
    .I0(n1bar),
    .I1(n2bar)
  );
  //OR U2
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2 (
    .O(n2),
    .I0(n3),
    .I1(n4)
  );
  //AND U2bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2bar (
    .O(n2bar),
    .I0(n3bar),
    .I1(n4bar)
  );
  //OR U3
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3 (
    .O(n4),
    .I0(n5),
    .I1(n6)
  );
  //AND U3bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3bar (
    .O(n4bar),
    .I0(n5bar),
    .I1(n6bar)
  );
  //OR U4
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4 (
    .O(n6),
    .I0(n7),
    .I1(n8)
  );
  //AND U4bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4bar (
    .O(n6bar),
    .I0(n7bar),
    .I1(n8bar)
  );
  //OR U5
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5 (
    .O(n5),
    .I0(n9),
    .I1(n10)
  );
  //AND U5bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5bar (
    .O(n5bar),
    .I0(n9bar),
    .I1(n10bar)
  );
  //OR U6
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6 (
    .O(n10),
    .I0(in[116]),
    .I1(n11)
  );
  //AND U6bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6bar (
    .O(n10bar),
    .I0(inbar[116]),
    .I1(n11bar)
  );
  //OR U7
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7 (
    .O(n3),
    .I0(n12),
    .I1(n13)
  );
  //AND U7bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7bar (
    .O(n3bar),
    .I0(n12bar),
    .I1(n13bar)
  );
  //OR U8
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8 (
    .O(n13),
    .I0(in[150]),
    .I1(in[127])
  );
  //AND U8bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8bar (
    .O(n13bar),
    .I0(inbar[150]),
    .I1(inbar[127])
  );
  //OR U9
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9 (
    .O(n12),
    .I0(in[160]),
    .I1(n14)
  );
  //AND U9bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9bar (
    .O(n12bar),
    .I0(inbar[160]),
    .I1(n14bar)
  );
  //OR U10
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10 (
    .O(n14),
    .I0(in[252]),
    .I1(in[168])
  );
  //AND U10bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10bar (
    .O(n14bar),
    .I0(inbar[252]),
    .I1(inbar[168])
  );
  //OR U11
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11 (
    .O(n1),
    .I0(n15),
    .I1(n16)
  );
  //AND U11bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11bar (
    .O(n1bar),
    .I0(n15bar),
    .I1(n16bar)
  );
  //OR U12
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12 (
    .O(n16),
    .I0(n17),
    .I1(n18)
  );
  //AND U12bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12bar (
    .O(n16bar),
    .I0(n17bar),
    .I1(n18bar)
  );
  //OR U13
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13 (
    .O(n18),
    .I0(in_17),
    .I1(in[96])
  );
  //AND U13bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13bar (
    .O(n18bar),
    .I0(in_17bar),
    .I1(inbar[96])
  );
  //OR U14
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14 (
    .O(n17),
    .I0(in_23),
    .I1(n19)
  );
  //AND U14bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14bar (
    .O(n17bar),
    .I0(in_23bar),
    .I1(n19bar)
  );
  //OR U15
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15 (
    .O(n19),
    .I0(in_31),
    .I1(in_26)
  );
  //AND U15bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15bar (
    .O(n19bar),
    .I0(in_31bar),
    .I1(in_26bar)
  );
  //OR U16
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16 (
    .O(n15),
    .I0(n20),
    .I1(n21)
  );
  //AND U16bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16bar (
    .O(n15bar),
    .I0(n20bar),
    .I1(n21bar)
  );
  //OR U17
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U17 (
    .O(n21),
    .I0(in_58),
    .I1(in_4)
  );
  //AND U17bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U17bar (
    .O(n21bar),
    .I0(in_58bar),
    .I1(in_4bar)
  );
  //OR U18
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U18 (
    .O(n20),
    .I0(in_59),
    .I1(n22)
  );
  //AND U18bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U18bar (
    .O(n20bar),
    .I0(in_59bar),
    .I1(n22bar)
  );
  //OR U19
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U19 (
    .O(n22),
    .I0(in_71),
    .I1(in_62)
  );
  //AND U19bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U19bar (
    .O(n22bar),
    .I0(in_71bar),
    .I1(in_62bar)
  );
  //OR U20
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U20 (
    .O(out[6]),
    .I0(n23),
    .I1(n24)
  );
  //AND U20bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U20bar (
    .O(outbar[6]),
    .I0(n23bar),
    .I1(n24bar)
  );
  //OR U21
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U21 (
    .O(n24),
    .I0(n25),
    .I1(n26)
  );
  //AND U21bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U21bar (
    .O(n24bar),
    .I0(n25bar),
    .I1(n26bar)
  );
  //OR U22
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U22 (
    .O(n26),
    .I0(n27),
    .I1(n28)
  );
  //AND U22bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U22bar (
    .O(n26bar),
    .I0(n27bar),
    .I1(n28bar)
  );
  //OR U23
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U23 (
    .O(n28),
    .I0(n29),
    .I1(n30)
  );
  //AND U23bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U23bar (
    .O(n28bar),
    .I0(n29bar),
    .I1(n30bar)
  );
  //OR U24
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U24 (
    .O(n27),
    .I0(n31),
    .I1(n32)
  );
  //AND U24bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U24bar (
    .O(n27bar),
    .I0(n31bar),
    .I1(n32bar)
  );
  //OR U25
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U25 (
    .O(n32),
    .I0(in[101]),
    .I1(n33)
  );
  //AND U25bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U25bar (
    .O(n32bar),
    .I0(inbar[101]),
    .I1(n33bar)
  );
  //OR U26
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U26 (
    .O(n25),
    .I0(n34),
    .I1(n35)
  );
  //AND U26bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U26bar (
    .O(n25bar),
    .I0(n34bar),
    .I1(n35bar)
  );
  //OR U27
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U27 (
    .O(n35),
    .I0(in[114]),
    .I1(in[104])
  );
  //AND U27bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U27bar (
    .O(n35bar),
    .I0(inbar[114]),
    .I1(inbar[104])
  );
  //OR U28
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U28 (
    .O(n34),
    .I0(in[128]),
    .I1(n36)
  );
  //AND U28bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U28bar (
    .O(n34bar),
    .I0(inbar[128]),
    .I1(n36bar)
  );
  //OR U29
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U29 (
    .O(n36),
    .I0(in[136]),
    .I1(in[134])
  );
  //AND U29bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U29bar (
    .O(n36bar),
    .I0(inbar[136]),
    .I1(inbar[134])
  );
  //OR U30
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U30 (
    .O(n23),
    .I0(n37),
    .I1(n38)
  );
  //AND U30bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U30bar (
    .O(n23bar),
    .I0(n37bar),
    .I1(n38bar)
  );
  //OR U31
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U31 (
    .O(n38),
    .I0(n39),
    .I1(n40)
  );
  //AND U31bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U31bar (
    .O(n38bar),
    .I0(n39bar),
    .I1(n40bar)
  );
  //OR U32
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U32 (
    .O(n40),
    .I0(in[177]),
    .I1(in[164])
  );
  //AND U32bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U32bar (
    .O(n40bar),
    .I0(inbar[177]),
    .I1(inbar[164])
  );
  //OR U33
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U33 (
    .O(n39),
    .I0(in[212]),
    .I1(n41)
  );
  //AND U33bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U33bar (
    .O(n39bar),
    .I0(inbar[212]),
    .I1(n41bar)
  );
  //OR U34
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U34 (
    .O(n41),
    .I0(in[248]),
    .I1(in[221])
  );
  //AND U34bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U34bar (
    .O(n41bar),
    .I0(inbar[248]),
    .I1(inbar[221])
  );
  //OR U35
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U35 (
    .O(n37),
    .I0(n42),
    .I1(n43)
  );
  //AND U35bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U35bar (
    .O(n37bar),
    .I0(n42bar),
    .I1(n43bar)
  );
  //OR U36
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U36 (
    .O(n43),
    .I0(in_18),
    .I1(in[93])
  );
  //AND U36bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U36bar (
    .O(n43bar),
    .I0(in_18bar),
    .I1(inbar[93])
  );
  //OR U37
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U37 (
    .O(n42),
    .I0(in_31),
    .I1(n44)
  );
  //AND U37bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U37bar (
    .O(n42bar),
    .I0(in_31bar),
    .I1(n44bar)
  );
  //OR U38
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U38 (
    .O(n44),
    .I0(in_7),
    .I1(in_39)
  );
  //AND U38bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U38bar (
    .O(n44bar),
    .I0(in_7bar),
    .I1(in_39bar)
  );
  //OR U39
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U39 (
    .O(out[5]),
    .I0(n45),
    .I1(n46)
  );
  //AND U39bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U39bar (
    .O(outbar[5]),
    .I0(n45bar),
    .I1(n46bar)
  );
  //OR U40
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U40 (
    .O(n46),
    .I0(n47),
    .I1(n48)
  );
  //AND U40bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U40bar (
    .O(n46bar),
    .I0(n47bar),
    .I1(n48bar)
  );
  //OR U41
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U41 (
    .O(n48),
    .I0(n49),
    .I1(n50)
  );
  //AND U41bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U41bar (
    .O(n48bar),
    .I0(n49bar),
    .I1(n50bar)
  );
  //OR U42
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U42 (
    .O(n50),
    .I0(n51),
    .I1(n52)
  );
  //AND U42bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U42bar (
    .O(n50bar),
    .I0(n51bar),
    .I1(n52bar)
  );
  //OR U43
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U43 (
    .O(n49),
    .I0(n33),
    .I1(n53)
  );
  //AND U43bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U43bar (
    .O(n49bar),
    .I0(n33bar),
    .I1(n53bar)
  );
  //OR U44
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U44 (
    .O(n53),
    .I0(in[111]),
    .I1(n54)
  );
  //AND U44bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U44bar (
    .O(n53bar),
    .I0(inbar[111]),
    .I1(n54bar)
  );
  //OR U45
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U45 (
    .O(n33),
    .I0(n55),
    .I1(n56)
  );
  //AND U45bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U45bar (
    .O(n33bar),
    .I0(n55bar),
    .I1(n56bar)
  );
  //OR U46
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U46 (
    .O(n56),
    .I0(n57),
    .I1(n58)
  );
  //AND U46bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U46bar (
    .O(n56bar),
    .I0(n57bar),
    .I1(n58bar)
  );
  //OR U47
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U47 (
    .O(n58),
    .I0(n59),
    .I1(n60)
  );
  //AND U47bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U47bar (
    .O(n58bar),
    .I0(n59bar),
    .I1(n60bar)
  );
  //OR U48
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U48 (
    .O(n60),
    .I0(in[140]),
    .I1(in[131])
  );
  //AND U48bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U48bar (
    .O(n60bar),
    .I0(inbar[140]),
    .I1(inbar[131])
  );
  //OR U49
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U49 (
    .O(n59),
    .I0(in[160]),
    .I1(in[144])
  );
  //AND U49bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U49bar (
    .O(n59bar),
    .I0(inbar[160]),
    .I1(inbar[144])
  );
  //OR U50
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U50 (
    .O(n57),
    .I0(n61),
    .I1(n62)
  );
  //AND U50bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U50bar (
    .O(n57bar),
    .I0(n61bar),
    .I1(n62bar)
  );
  //OR U51
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U51 (
    .O(n62),
    .I0(in[179]),
    .I1(in[174])
  );
  //AND U51bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U51bar (
    .O(n62bar),
    .I0(inbar[179]),
    .I1(inbar[174])
  );
  //OR U52
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U52 (
    .O(n61),
    .I0(in[188]),
    .I1(in[184])
  );
  //AND U52bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U52bar (
    .O(n61bar),
    .I0(inbar[188]),
    .I1(inbar[184])
  );
  //OR U53
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U53 (
    .O(n55),
    .I0(n63),
    .I1(n64)
  );
  //AND U53bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U53bar (
    .O(n55bar),
    .I0(n63bar),
    .I1(n64bar)
  );
  //OR U54
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U54 (
    .O(n64),
    .I0(n65),
    .I1(n66)
  );
  //AND U54bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U54bar (
    .O(n64bar),
    .I0(n65bar),
    .I1(n66bar)
  );
  //OR U55
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U55 (
    .O(n66),
    .I0(in[216]),
    .I1(in[200])
  );
  //AND U55bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U55bar (
    .O(n66bar),
    .I0(inbar[216]),
    .I1(inbar[200])
  );
  //OR U56
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U56 (
    .O(n65),
    .I0(in[228]),
    .I1(in[224])
  );
  //AND U56bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U56bar (
    .O(n65bar),
    .I0(inbar[228]),
    .I1(inbar[224])
  );
  //OR U57
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U57 (
    .O(n63),
    .I0(n67),
    .I1(n68)
  );
  //AND U57bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U57bar (
    .O(n63bar),
    .I0(n67bar),
    .I1(n68bar)
  );
  //OR U58
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U58 (
    .O(n68),
    .I0(in[247]),
    .I1(in[235])
  );
  //AND U58bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U58bar (
    .O(n68bar),
    .I0(inbar[247]),
    .I1(inbar[235])
  );
  //OR U59
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U59 (
    .O(n67),
    .I0(in_42),
    .I1(in[83])
  );
  //AND U59bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U59bar (
    .O(n67bar),
    .I0(in_42bar),
    .I1(inbar[83])
  );
  //OR U60
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U60 (
    .O(n47),
    .I0(n69),
    .I1(n70)
  );
  //AND U60bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U60bar (
    .O(n47bar),
    .I0(n69bar),
    .I1(n70bar)
  );
  //OR U61
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U61 (
    .O(n70),
    .I0(in[166]),
    .I1(in[123])
  );
  //AND U61bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U61bar (
    .O(n70bar),
    .I0(inbar[166]),
    .I1(inbar[123])
  );
  //OR U62
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U62 (
    .O(n69),
    .I0(in[170]),
    .I1(n71)
  );
  //AND U62bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U62bar (
    .O(n69bar),
    .I0(inbar[170]),
    .I1(n71bar)
  );
  //OR U63
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U63 (
    .O(n71),
    .I0(in[194]),
    .I1(in[183])
  );
  //AND U63bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U63bar (
    .O(n71bar),
    .I0(inbar[194]),
    .I1(inbar[183])
  );
  //OR U64
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U64 (
    .O(n45),
    .I0(n72),
    .I1(n73)
  );
  //AND U64bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U64bar (
    .O(n45bar),
    .I0(n72bar),
    .I1(n73bar)
  );
  //OR U65
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U65 (
    .O(n73),
    .I0(n74),
    .I1(n75)
  );
  //AND U65bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U65bar (
    .O(n73bar),
    .I0(n74bar),
    .I1(n75bar)
  );
  //OR U66
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U66 (
    .O(n75),
    .I0(in[241]),
    .I1(in[238])
  );
  //AND U66bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U66bar (
    .O(n75bar),
    .I0(inbar[241]),
    .I1(inbar[238])
  );
  //OR U67
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U67 (
    .O(n74),
    .I0(in[250]),
    .I1(n76)
  );
  //AND U67bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U67bar (
    .O(n74bar),
    .I0(inbar[250]),
    .I1(n76bar)
  );
  //OR U68
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U68 (
    .O(n76),
    .I0(in_24),
    .I1(in[84])
  );
  //AND U68bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U68bar (
    .O(n76bar),
    .I0(in_24bar),
    .I1(inbar[84])
  );
  //OR U69
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U69 (
    .O(n72),
    .I0(n77),
    .I1(n78)
  );
  //AND U69bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U69bar (
    .O(n72bar),
    .I0(n77bar),
    .I1(n78bar)
  );
  //OR U70
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U70 (
    .O(n78),
    .I0(in_41),
    .I1(in_29)
  );
  //AND U70bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U70bar (
    .O(n78bar),
    .I0(in_41bar),
    .I1(in_29bar)
  );
  //OR U71
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U71 (
    .O(n77),
    .I0(in_66),
    .I1(n79)
  );
  //AND U71bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U71bar (
    .O(n77bar),
    .I0(in_66bar),
    .I1(n79bar)
  );
  //OR U72
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U72 (
    .O(n79),
    .I0(in_76),
    .I1(in_71)
  );
  //AND U72bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U72bar (
    .O(n79bar),
    .I0(in_76bar),
    .I1(in_71bar)
  );
  //OR U73
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U73 (
    .O(out[4]),
    .I0(n80),
    .I1(n81)
  );
  //AND U73bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U73bar (
    .O(outbar[4]),
    .I0(n80bar),
    .I1(n81bar)
  );
  //OR U74
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U74 (
    .O(n81),
    .I0(n82),
    .I1(n83)
  );
  //AND U74bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U74bar (
    .O(n81bar),
    .I0(n82bar),
    .I1(n83bar)
  );
  //OR U75
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U75 (
    .O(n83),
    .I0(n84),
    .I1(n85)
  );
  //AND U75bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U75bar (
    .O(n83bar),
    .I0(n84bar),
    .I1(n85bar)
  );
  //OR U76
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U76 (
    .O(n85),
    .I0(n51),
    .I1(n86)
  );
  //AND U76bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U76bar (
    .O(n85bar),
    .I0(n51bar),
    .I1(n86bar)
  );
  //OR U77
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U77 (
    .O(n51),
    .I0(n87),
    .I1(n88)
  );
  //AND U77bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U77bar (
    .O(n51bar),
    .I0(n87bar),
    .I1(n88bar)
  );
  //OR U78
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U78 (
    .O(n88),
    .I0(n89),
    .I1(n90)
  );
  //AND U78bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U78bar (
    .O(n88bar),
    .I0(n89bar),
    .I1(n90bar)
  );
  //OR U79
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U79 (
    .O(n90),
    .I0(n91),
    .I1(n92)
  );
  //AND U79bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U79bar (
    .O(n90bar),
    .I0(n91bar),
    .I1(n92bar)
  );
  //OR U80
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U80 (
    .O(n92),
    .I0(in[118]),
    .I1(in[109])
  );
  //AND U80bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U80bar (
    .O(n92bar),
    .I0(inbar[118]),
    .I1(inbar[109])
  );
  //OR U81
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U81 (
    .O(n91),
    .I0(in[139]),
    .I1(in[120])
  );
  //AND U81bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U81bar (
    .O(n91bar),
    .I0(inbar[139]),
    .I1(inbar[120])
  );
  //OR U82
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U82 (
    .O(n89),
    .I0(n93),
    .I1(n94)
  );
  //AND U82bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U82bar (
    .O(n89bar),
    .I0(n93bar),
    .I1(n94bar)
  );
  //OR U83
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U83 (
    .O(n94),
    .I0(in[198]),
    .I1(in[154])
  );
  //AND U83bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U83bar (
    .O(n94bar),
    .I0(inbar[198]),
    .I1(inbar[154])
  );
  //OR U84
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U84 (
    .O(n93),
    .I0(in[210]),
    .I1(in[205])
  );
  //AND U84bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U84bar (
    .O(n93bar),
    .I0(inbar[210]),
    .I1(inbar[205])
  );
  //OR U85
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U85 (
    .O(n87),
    .I0(n95),
    .I1(n96)
  );
  //AND U85bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U85bar (
    .O(n87bar),
    .I0(n95bar),
    .I1(n96bar)
  );
  //OR U86
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U86 (
    .O(n96),
    .I0(n97),
    .I1(n98)
  );
  //AND U86bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U86bar (
    .O(n96bar),
    .I0(n97bar),
    .I1(n98bar)
  );
  //OR U87
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U87 (
    .O(n98),
    .I0(in[219]),
    .I1(in[217])
  );
  //AND U87bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U87bar (
    .O(n98bar),
    .I0(inbar[219]),
    .I1(inbar[217])
  );
  //OR U88
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U88 (
    .O(n97),
    .I0(in[86]),
    .I1(in[252])
  );
  //AND U88bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U88bar (
    .O(n97bar),
    .I0(inbar[86]),
    .I1(inbar[252])
  );
  //OR U89
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U89 (
    .O(n95),
    .I0(n99),
    .I1(n100)
  );
  //AND U89bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U89bar (
    .O(n95bar),
    .I0(n99bar),
    .I1(n100bar)
  );
  //OR U90
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U90 (
    .O(n100),
    .I0(in_40),
    .I1(in[91])
  );
  //AND U90bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U90bar (
    .O(n100bar),
    .I0(in_40bar),
    .I1(inbar[91])
  );
  //OR U91
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U91 (
    .O(n99),
    .I0(in_8),
    .I1(in_46)
  );
  //AND U91bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U91bar (
    .O(n99bar),
    .I0(in_8bar),
    .I1(in_46bar)
  );
  //OR U92
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U92 (
    .O(n84),
    .I0(n101),
    .I1(n102)
  );
  //AND U92bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U92bar (
    .O(n84bar),
    .I0(n101bar),
    .I1(n102bar)
  );
  //OR U93
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U93 (
    .O(n102),
    .I0(in[117]),
    .I1(n30)
  );
  //AND U93bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U93bar (
    .O(n102bar),
    .I0(inbar[117]),
    .I1(n30bar)
  );
  //OR U94
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U94 (
    .O(n30),
    .I0(n103),
    .I1(n104)
  );
  //AND U94bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U94bar (
    .O(n30bar),
    .I0(n103bar),
    .I1(n104bar)
  );
  //OR U95
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U95 (
    .O(n104),
    .I0(n105),
    .I1(n106)
  );
  //AND U95bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U95bar (
    .O(n104bar),
    .I0(n105bar),
    .I1(n106bar)
  );
  //OR U96
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U96 (
    .O(n106),
    .I0(n107),
    .I1(n108)
  );
  //AND U96bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U96bar (
    .O(n106bar),
    .I0(n107bar),
    .I1(n108bar)
  );
  //OR U97
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U97 (
    .O(n108),
    .I0(n109),
    .I1(n110)
  );
  //AND U97bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U97bar (
    .O(n108bar),
    .I0(n109bar),
    .I1(n110bar)
  );
  //OR U98
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U98 (
    .O(n107),
    .I0(in[108]),
    .I1(n54)
  );
  //AND U98bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U98bar (
    .O(n107bar),
    .I0(inbar[108]),
    .I1(n54bar)
  );
  //OR U99
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U99 (
    .O(n54),
    .I0(n111),
    .I1(n112)
  );
  //AND U99bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U99bar (
    .O(n54bar),
    .I0(n111bar),
    .I1(n112bar)
  );
  //OR U100
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U100 (
    .O(n112),
    .I0(n113),
    .I1(n114)
  );
  //AND U100bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U100bar (
    .O(n112bar),
    .I0(n113bar),
    .I1(n114bar)
  );
  //OR U101
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U101 (
    .O(n114),
    .I0(n115),
    .I1(n116)
  );
  //AND U101bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U101bar (
    .O(n114bar),
    .I0(n115bar),
    .I1(n116bar)
  );
  //OR U102
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U102 (
    .O(n116),
    .I0(in[119]),
    .I1(in[105])
  );
  //AND U102bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U102bar (
    .O(n116bar),
    .I0(inbar[119]),
    .I1(inbar[105])
  );
  //OR U103
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U103 (
    .O(n115),
    .I0(in[186]),
    .I1(in[175])
  );
  //AND U103bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U103bar (
    .O(n115bar),
    .I0(inbar[186]),
    .I1(inbar[175])
  );
  //OR U104
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U104 (
    .O(n113),
    .I0(n117),
    .I1(n118)
  );
  //AND U104bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U104bar (
    .O(n113bar),
    .I0(n117bar),
    .I1(n118bar)
  );
  //OR U105
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U105 (
    .O(n118),
    .I0(in[202]),
    .I1(in[193])
  );
  //AND U105bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U105bar (
    .O(n118bar),
    .I0(inbar[202]),
    .I1(inbar[193])
  );
  //OR U106
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U106 (
    .O(n117),
    .I0(in[225]),
    .I1(in[208])
  );
  //AND U106bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U106bar (
    .O(n117bar),
    .I0(inbar[225]),
    .I1(inbar[208])
  );
  //OR U107
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U107 (
    .O(n111),
    .I0(n119),
    .I1(n120)
  );
  //AND U107bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U107bar (
    .O(n111bar),
    .I0(n119bar),
    .I1(n120bar)
  );
  //OR U108
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U108 (
    .O(n120),
    .I0(n121),
    .I1(n122)
  );
  //AND U108bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U108bar (
    .O(n120bar),
    .I0(n121bar),
    .I1(n122bar)
  );
  //OR U109
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U109 (
    .O(n122),
    .I0(in_1),
    .I1(in[85])
  );
  //AND U109bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U109bar (
    .O(n122bar),
    .I0(in_1bar),
    .I1(inbar[85])
  );
  //OR U110
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U110 (
    .O(n121),
    .I0(in_23),
    .I1(in_19)
  );
  //AND U110bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U110bar (
    .O(n121bar),
    .I0(in_23bar),
    .I1(in_19bar)
  );
  //OR U111
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U111 (
    .O(n119),
    .I0(n123),
    .I1(n124)
  );
  //AND U111bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U111bar (
    .O(n119bar),
    .I0(n123bar),
    .I1(n124bar)
  );
  //OR U112
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U112 (
    .O(n124),
    .I0(in_43),
    .I1(in_33)
  );
  //AND U112bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U112bar (
    .O(n124bar),
    .I0(in_43bar),
    .I1(in_33bar)
  );
  //OR U113
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U113 (
    .O(n123),
    .I0(in_63),
    .I1(in_44)
  );
  //AND U113bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U113bar (
    .O(n123bar),
    .I0(in_63bar),
    .I1(in_44bar)
  );
  //OR U114
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U114 (
    .O(n105),
    .I0(n125),
    .I1(n126)
  );
  //AND U114bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U114bar (
    .O(n105bar),
    .I0(n125bar),
    .I1(n126bar)
  );
  //OR U115
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U115 (
    .O(n126),
    .I0(in[141]),
    .I1(in[112])
  );
  //AND U115bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U115bar (
    .O(n126bar),
    .I0(inbar[141]),
    .I1(inbar[112])
  );
  //OR U116
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U116 (
    .O(n125),
    .I0(in[147]),
    .I1(n127)
  );
  //AND U116bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U116bar (
    .O(n125bar),
    .I0(inbar[147]),
    .I1(n127bar)
  );
  //OR U117
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U117 (
    .O(n127),
    .I0(in[181]),
    .I1(in[167])
  );
  //AND U117bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U117bar (
    .O(n127bar),
    .I0(inbar[181]),
    .I1(inbar[167])
  );
  //OR U118
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U118 (
    .O(n103),
    .I0(n128),
    .I1(n129)
  );
  //AND U118bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U118bar (
    .O(n103bar),
    .I0(n128bar),
    .I1(n129bar)
  );
  //OR U119
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U119 (
    .O(n129),
    .I0(n130),
    .I1(n131)
  );
  //AND U119bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U119bar (
    .O(n129bar),
    .I0(n130bar),
    .I1(n131bar)
  );
  //OR U120
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U120 (
    .O(n131),
    .I0(in[229]),
    .I1(in[201])
  );
  //AND U120bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U120bar (
    .O(n131bar),
    .I0(inbar[229]),
    .I1(inbar[201])
  );
  //OR U121
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U121 (
    .O(n130),
    .I0(in[237]),
    .I1(n132)
  );
  //AND U121bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U121bar (
    .O(n130bar),
    .I0(inbar[237]),
    .I1(n132bar)
  );
  //OR U122
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U122 (
    .O(n132),
    .I0(in[94]),
    .I1(in[253])
  );
  //AND U122bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U122bar (
    .O(n132bar),
    .I0(inbar[94]),
    .I1(inbar[253])
  );
  //OR U123
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U123 (
    .O(n128),
    .I0(n133),
    .I1(n134)
  );
  //AND U123bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U123bar (
    .O(n128bar),
    .I0(n133bar),
    .I1(n134bar)
  );
  //OR U124
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U124 (
    .O(n134),
    .I0(in_21),
    .I1(in[96])
  );
  //AND U124bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U124bar (
    .O(n134bar),
    .I0(in_21bar),
    .I1(inbar[96])
  );
  //OR U125
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U125 (
    .O(n133),
    .I0(in_25),
    .I1(n135)
  );
  //AND U125bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U125bar (
    .O(n133bar),
    .I0(in_25bar),
    .I1(n135bar)
  );
  //OR U126
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U126 (
    .O(n135),
    .I0(in_81),
    .I1(in_45)
  );
  //AND U126bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U126bar (
    .O(n135bar),
    .I0(in_81bar),
    .I1(in_45bar)
  );
  //OR U127
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U127 (
    .O(n82),
    .I0(n136),
    .I1(n137)
  );
  //AND U127bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U127bar (
    .O(n82bar),
    .I0(n136bar),
    .I1(n137bar)
  );
  //OR U128
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U128 (
    .O(n137),
    .I0(in[142]),
    .I1(in[124])
  );
  //AND U128bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U128bar (
    .O(n137bar),
    .I0(inbar[142]),
    .I1(inbar[124])
  );
  //OR U129
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U129 (
    .O(n136),
    .I0(in[150]),
    .I1(n138)
  );
  //AND U129bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U129bar (
    .O(n136bar),
    .I0(inbar[150]),
    .I1(n138bar)
  );
  //OR U130
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U130 (
    .O(n138),
    .I0(in[172]),
    .I1(in[155])
  );
  //AND U130bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U130bar (
    .O(n138bar),
    .I0(inbar[172]),
    .I1(inbar[155])
  );
  //OR U131
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U131 (
    .O(n80),
    .I0(n139),
    .I1(n140)
  );
  //AND U131bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U131bar (
    .O(n80bar),
    .I0(n139bar),
    .I1(n140bar)
  );
  //OR U132
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U132 (
    .O(n140),
    .I0(n141),
    .I1(n142)
  );
  //AND U132bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U132bar (
    .O(n140bar),
    .I0(n141bar),
    .I1(n142bar)
  );
  //OR U133
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U133 (
    .O(n142),
    .I0(in[196]),
    .I1(in[173])
  );
  //AND U133bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U133bar (
    .O(n142bar),
    .I0(inbar[196]),
    .I1(inbar[173])
  );
  //OR U134
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U134 (
    .O(n141),
    .I0(in[222]),
    .I1(n143)
  );
  //AND U134bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U134bar (
    .O(n141bar),
    .I0(inbar[222]),
    .I1(n143bar)
  );
  //OR U135
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U135 (
    .O(n143),
    .I0(in[227]),
    .I1(in[226])
  );
  //AND U135bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U135bar (
    .O(n143bar),
    .I0(inbar[227]),
    .I1(inbar[226])
  );
  //OR U136
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U136 (
    .O(n139),
    .I0(n144),
    .I1(n145)
  );
  //AND U136bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U136bar (
    .O(n139bar),
    .I0(n144bar),
    .I1(n145bar)
  );
  //OR U137
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U137 (
    .O(n145),
    .I0(in[249]),
    .I1(in[231])
  );
  //AND U137bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U137bar (
    .O(n145bar),
    .I0(inbar[249]),
    .I1(inbar[231])
  );
  //OR U138
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U138 (
    .O(n144),
    .I0(in_28),
    .I1(n146)
  );
  //AND U138bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U138bar (
    .O(n144bar),
    .I0(in_28bar),
    .I1(n146bar)
  );
  //OR U139
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U139 (
    .O(n146),
    .I0(in_52),
    .I1(in_47)
  );
  //AND U139bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U139bar (
    .O(n146bar),
    .I0(in_52bar),
    .I1(in_47bar)
  );
  //OR U140
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U140 (
    .O(out[3]),
    .I0(n147),
    .I1(n148)
  );
  //AND U140bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U140bar (
    .O(outbar[3]),
    .I0(n147bar),
    .I1(n148bar)
  );
  //OR U141
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U141 (
    .O(n148),
    .I0(n149),
    .I1(n150)
  );
  //AND U141bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U141bar (
    .O(n148bar),
    .I0(n149bar),
    .I1(n150bar)
  );
  //OR U142
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U142 (
    .O(n150),
    .I0(n151),
    .I1(n152)
  );
  //AND U142bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U142bar (
    .O(n150bar),
    .I0(n151bar),
    .I1(n152bar)
  );
  //OR U143
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U143 (
    .O(n152),
    .I0(n153),
    .I1(n154)
  );
  //AND U143bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U143bar (
    .O(n152bar),
    .I0(n153bar),
    .I1(n154bar)
  );
  //OR U144
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U144 (
    .O(n151),
    .I0(n9),
    .I1(n155)
  );
  //AND U144bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U144bar (
    .O(n151bar),
    .I0(n9bar),
    .I1(n155bar)
  );
  //OR U145
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U145 (
    .O(n155),
    .I0(in[118]),
    .I1(n156)
  );
  //AND U145bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U145bar (
    .O(n155bar),
    .I0(inbar[118]),
    .I1(n156bar)
  );
  //OR U146
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U146 (
    .O(n9),
    .I0(n157),
    .I1(n158)
  );
  //AND U146bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U146bar (
    .O(n9bar),
    .I0(n157bar),
    .I1(n158bar)
  );
  //OR U147
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U147 (
    .O(n158),
    .I0(n159),
    .I1(n160)
  );
  //AND U147bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U147bar (
    .O(n158bar),
    .I0(n159bar),
    .I1(n160bar)
  );
  //OR U148
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U148 (
    .O(n160),
    .I0(n161),
    .I1(n162)
  );
  //AND U148bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U148bar (
    .O(n160bar),
    .I0(n161bar),
    .I1(n162bar)
  );
  //OR U149
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U149 (
    .O(n162),
    .I0(in[122]),
    .I1(in[111])
  );
  //AND U149bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U149bar (
    .O(n162bar),
    .I0(inbar[122]),
    .I1(inbar[111])
  );
  //OR U150
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U150 (
    .O(n161),
    .I0(in[154]),
    .I1(in[151])
  );
  //AND U150bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U150bar (
    .O(n161bar),
    .I0(inbar[154]),
    .I1(inbar[151])
  );
  //OR U151
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U151 (
    .O(n159),
    .I0(n163),
    .I1(n164)
  );
  //AND U151bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U151bar (
    .O(n159bar),
    .I0(n163bar),
    .I1(n164bar)
  );
  //OR U152
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U152 (
    .O(n164),
    .I0(in[187]),
    .I1(in[177])
  );
  //AND U152bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U152bar (
    .O(n164bar),
    .I0(inbar[187]),
    .I1(inbar[177])
  );
  //OR U153
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U153 (
    .O(n163),
    .I0(in[200]),
    .I1(in[192])
  );
  //AND U153bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U153bar (
    .O(n163bar),
    .I0(inbar[200]),
    .I1(inbar[192])
  );
  //OR U154
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U154 (
    .O(n157),
    .I0(n165),
    .I1(n166)
  );
  //AND U154bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U154bar (
    .O(n157bar),
    .I0(n165bar),
    .I1(n166bar)
  );
  //OR U155
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U155 (
    .O(n166),
    .I0(n167),
    .I1(n168)
  );
  //AND U155bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U155bar (
    .O(n166bar),
    .I0(n167bar),
    .I1(n168bar)
  );
  //OR U156
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U156 (
    .O(n168),
    .I0(in[225]),
    .I1(in[207])
  );
  //AND U156bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U156bar (
    .O(n168bar),
    .I0(inbar[225]),
    .I1(inbar[207])
  );
  //OR U157
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U157 (
    .O(n167),
    .I0(in[98]),
    .I1(in[226])
  );
  //AND U157bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U157bar (
    .O(n167bar),
    .I0(inbar[98]),
    .I1(inbar[226])
  );
  //OR U158
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U158 (
    .O(n165),
    .I0(n169),
    .I1(n170)
  );
  //AND U158bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U158bar (
    .O(n165bar),
    .I0(n169bar),
    .I1(n170bar)
  );
  //OR U159
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U159 (
    .O(n170),
    .I0(in_20),
    .I1(in_16)
  );
  //AND U159bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U159bar (
    .O(n170bar),
    .I0(in_20bar),
    .I1(in_16bar)
  );
  //OR U160
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U160 (
    .O(n169),
    .I0(in_55),
    .I1(in_45)
  );
  //AND U160bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U160bar (
    .O(n169bar),
    .I0(in_55bar),
    .I1(in_45bar)
  );
  //OR U161
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U161 (
    .O(n149),
    .I0(n171),
    .I1(n172)
  );
  //AND U161bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U161bar (
    .O(n149bar),
    .I0(n171bar),
    .I1(n172bar)
  );
  //OR U162
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U162 (
    .O(n172),
    .I0(in[162]),
    .I1(in[149])
  );
  //AND U162bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U162bar (
    .O(n172bar),
    .I0(inbar[162]),
    .I1(inbar[149])
  );
  //OR U163
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U163 (
    .O(n171),
    .I0(in[163]),
    .I1(n173)
  );
  //AND U163bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U163bar (
    .O(n171bar),
    .I0(inbar[163]),
    .I1(n173bar)
  );
  //OR U164
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U164 (
    .O(n173),
    .I0(in[191]),
    .I1(in[189])
  );
  //AND U164bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U164bar (
    .O(n173bar),
    .I0(inbar[191]),
    .I1(inbar[189])
  );
  //OR U165
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U165 (
    .O(n147),
    .I0(n174),
    .I1(n175)
  );
  //AND U165bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U165bar (
    .O(n147bar),
    .I0(n174bar),
    .I1(n175bar)
  );
  //OR U166
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U166 (
    .O(n175),
    .I0(n176),
    .I1(n177)
  );
  //AND U166bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U166bar (
    .O(n175bar),
    .I0(n176bar),
    .I1(n177bar)
  );
  //OR U167
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U167 (
    .O(n177),
    .I0(in[212]),
    .I1(in[193])
  );
  //AND U167bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U167bar (
    .O(n177bar),
    .I0(inbar[212]),
    .I1(inbar[193])
  );
  //OR U168
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U168 (
    .O(n176),
    .I0(in[238]),
    .I1(n178)
  );
  //AND U168bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U168bar (
    .O(n176bar),
    .I0(inbar[238]),
    .I1(n178bar)
  );
  //OR U169
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U169 (
    .O(n178),
    .I0(in[88]),
    .I1(in[247])
  );
  //AND U169bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U169bar (
    .O(n178bar),
    .I0(inbar[88]),
    .I1(inbar[247])
  );
  //OR U170
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U170 (
    .O(n174),
    .I0(n179),
    .I1(n180)
  );
  //AND U170bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U170bar (
    .O(n174bar),
    .I0(n179bar),
    .I1(n180bar)
  );
  //OR U171
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U171 (
    .O(n180),
    .I0(in[94]),
    .I1(in[92])
  );
  //AND U171bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U171bar (
    .O(n180bar),
    .I0(inbar[94]),
    .I1(inbar[92])
  );
  //OR U172
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U172 (
    .O(n179),
    .I0(in_52),
    .I1(n181)
  );
  //AND U172bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U172bar (
    .O(n179bar),
    .I0(in_52bar),
    .I1(n181bar)
  );
  //OR U173
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U173 (
    .O(n181),
    .I0(in_70),
    .I1(in_67)
  );
  //AND U173bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U173bar (
    .O(n181bar),
    .I0(in_70bar),
    .I1(in_67bar)
  );
  //OR U174
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U174 (
    .O(out[2]),
    .I0(n182),
    .I1(n183)
  );
  //AND U174bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U174bar (
    .O(outbar[2]),
    .I0(n182bar),
    .I1(n183bar)
  );
  //OR U175
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U175 (
    .O(n183),
    .I0(n184),
    .I1(n185)
  );
  //AND U175bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U175bar (
    .O(n183bar),
    .I0(n184bar),
    .I1(n185bar)
  );
  //OR U176
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U176 (
    .O(n185),
    .I0(n186),
    .I1(n187)
  );
  //AND U176bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U176bar (
    .O(n185bar),
    .I0(n186bar),
    .I1(n187bar)
  );
  //OR U177
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U177 (
    .O(n187),
    .I0(n154),
    .I1(n188)
  );
  //AND U177bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U177bar (
    .O(n187bar),
    .I0(n154bar),
    .I1(n188bar)
  );
  //OR U178
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U178 (
    .O(n154),
    .I0(n189),
    .I1(n190)
  );
  //AND U178bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U178bar (
    .O(n154bar),
    .I0(n189bar),
    .I1(n190bar)
  );
  //OR U179
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U179 (
    .O(n190),
    .I0(n191),
    .I1(n192)
  );
  //AND U179bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U179bar (
    .O(n190bar),
    .I0(n191bar),
    .I1(n192bar)
  );
  //OR U180
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U180 (
    .O(n192),
    .I0(n193),
    .I1(n194)
  );
  //AND U180bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U180bar (
    .O(n192bar),
    .I0(n193bar),
    .I1(n194bar)
  );
  //OR U181
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U181 (
    .O(n194),
    .I0(n11),
    .I1(n195)
  );
  //AND U181bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U181bar (
    .O(n194bar),
    .I0(n11bar),
    .I1(n195bar)
  );
  //OR U182
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U182 (
    .O(n11),
    .I0(n196),
    .I1(n197)
  );
  //AND U182bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U182bar (
    .O(n11bar),
    .I0(n196bar),
    .I1(n197bar)
  );
  //OR U183
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U183 (
    .O(n197),
    .I0(n198),
    .I1(n199)
  );
  //AND U183bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U183bar (
    .O(n197bar),
    .I0(n198bar),
    .I1(n199bar)
  );
  //OR U184
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U184 (
    .O(n199),
    .I0(n200),
    .I1(n201)
  );
  //AND U184bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U184bar (
    .O(n199bar),
    .I0(n200bar),
    .I1(n201bar)
  );
  //OR U185
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U185 (
    .O(n201),
    .I0(in[131]),
    .I1(in[120])
  );
  //AND U185bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U185bar (
    .O(n201bar),
    .I0(inbar[131]),
    .I1(inbar[120])
  );
  //OR U186
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U186 (
    .O(n200),
    .I0(in[153]),
    .I1(in[147])
  );
  //AND U186bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U186bar (
    .O(n200bar),
    .I0(inbar[153]),
    .I1(inbar[147])
  );
  //OR U187
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U187 (
    .O(n198),
    .I0(n202),
    .I1(n203)
  );
  //AND U187bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U187bar (
    .O(n198bar),
    .I0(n202bar),
    .I1(n203bar)
  );
  //OR U188
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U188 (
    .O(n203),
    .I0(in[170]),
    .I1(in[156])
  );
  //AND U188bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U188bar (
    .O(n203bar),
    .I0(inbar[170]),
    .I1(inbar[156])
  );
  //OR U189
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U189 (
    .O(n202),
    .I0(in[223]),
    .I1(in[190])
  );
  //AND U189bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U189bar (
    .O(n202bar),
    .I0(inbar[223]),
    .I1(inbar[190])
  );
  //OR U190
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U190 (
    .O(n196),
    .I0(n204),
    .I1(n205)
  );
  //AND U190bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U190bar (
    .O(n196bar),
    .I0(n204bar),
    .I1(n205bar)
  );
  //OR U191
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U191 (
    .O(n205),
    .I0(n206),
    .I1(n207)
  );
  //AND U191bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U191bar (
    .O(n205bar),
    .I0(n206bar),
    .I1(n207bar)
  );
  //OR U192
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U192 (
    .O(n207),
    .I0(in[236]),
    .I1(in[230])
  );
  //AND U192bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U192bar (
    .O(n207bar),
    .I0(inbar[236]),
    .I1(inbar[230])
  );
  //OR U193
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U193 (
    .O(n206),
    .I0(in[85]),
    .I1(in[240])
  );
  //AND U193bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U193bar (
    .O(n206bar),
    .I0(inbar[85]),
    .I1(inbar[240])
  );
  //OR U194
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U194 (
    .O(n204),
    .I0(n208),
    .I1(n209)
  );
  //AND U194bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U194bar (
    .O(n204bar),
    .I0(n208bar),
    .I1(n209bar)
  );
  //OR U195
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U195 (
    .O(n209),
    .I0(in_12),
    .I1(in[90])
  );
  //AND U195bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U195bar (
    .O(n209bar),
    .I0(in_12bar),
    .I1(inbar[90])
  );
  //OR U196
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U196 (
    .O(n208),
    .I0(in_39),
    .I1(in_28)
  );
  //AND U196bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U196bar (
    .O(n208bar),
    .I0(in_39bar),
    .I1(in_28bar)
  );
  //OR U197
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U197 (
    .O(n193),
    .I0(in[109]),
    .I1(n210)
  );
  //AND U197bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U197bar (
    .O(n193bar),
    .I0(inbar[109]),
    .I1(n210bar)
  );
  //OR U198
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U198 (
    .O(n191),
    .I0(n211),
    .I1(n212)
  );
  //AND U198bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U198bar (
    .O(n191bar),
    .I0(n211bar),
    .I1(n212bar)
  );
  //OR U199
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U199 (
    .O(n212),
    .I0(in[138]),
    .I1(in[129])
  );
  //AND U199bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U199bar (
    .O(n212bar),
    .I0(inbar[138]),
    .I1(inbar[129])
  );
  //OR U200
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U200 (
    .O(n211),
    .I0(in[157]),
    .I1(n213)
  );
  //AND U200bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U200bar (
    .O(n211bar),
    .I0(inbar[157]),
    .I1(n213bar)
  );
  //OR U201
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U201 (
    .O(n213),
    .I0(in[182]),
    .I1(in[167])
  );
  //AND U201bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U201bar (
    .O(n213bar),
    .I0(inbar[182]),
    .I1(inbar[167])
  );
  //OR U202
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U202 (
    .O(n189),
    .I0(n214),
    .I1(n215)
  );
  //AND U202bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U202bar (
    .O(n189bar),
    .I0(n214bar),
    .I1(n215bar)
  );
  //OR U203
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U203 (
    .O(n215),
    .I0(n216),
    .I1(n217)
  );
  //AND U203bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U203bar (
    .O(n215bar),
    .I0(n216bar),
    .I1(n217bar)
  );
  //OR U204
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U204 (
    .O(n217),
    .I0(in[195]),
    .I1(in[184])
  );
  //AND U204bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U204bar (
    .O(n217bar),
    .I0(inbar[195]),
    .I1(inbar[184])
  );
  //OR U205
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U205 (
    .O(n216),
    .I0(in[196]),
    .I1(n218)
  );
  //AND U205bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U205bar (
    .O(n216bar),
    .I0(inbar[196]),
    .I1(n218bar)
  );
  //OR U206
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U206 (
    .O(n218),
    .I0(in[215]),
    .I1(in[209])
  );
  //AND U206bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U206bar (
    .O(n218bar),
    .I0(inbar[215]),
    .I1(inbar[209])
  );
  //OR U207
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U207 (
    .O(n214),
    .I0(n219),
    .I1(n220)
  );
  //AND U207bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U207bar (
    .O(n214bar),
    .I0(n219bar),
    .I1(n220bar)
  );
  //OR U208
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U208 (
    .O(n220),
    .I0(in[93]),
    .I1(in[233])
  );
  //AND U208bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U208bar (
    .O(n220bar),
    .I0(inbar[93]),
    .I1(inbar[233])
  );
  //OR U209
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U209 (
    .O(n219),
    .I0(in_1),
    .I1(n221)
  );
  //AND U209bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U209bar (
    .O(n219bar),
    .I0(in_1bar),
    .I1(n221bar)
  );
  //OR U210
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U210 (
    .O(n221),
    .I0(in_69),
    .I1(in_66)
  );
  //AND U210bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U210bar (
    .O(n221bar),
    .I0(in_69bar),
    .I1(in_66bar)
  );
  //OR U211
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U211 (
    .O(n186),
    .I0(n7),
    .I1(n222)
  );
  //AND U211bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U211bar (
    .O(n186bar),
    .I0(n7bar),
    .I1(n222bar)
  );
  //OR U212
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U212 (
    .O(n222),
    .I0(in[134]),
    .I1(n223)
  );
  //AND U212bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U212bar (
    .O(n222bar),
    .I0(inbar[134]),
    .I1(n223bar)
  );
  //OR U213
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U213 (
    .O(n7),
    .I0(n224),
    .I1(n225)
  );
  //AND U213bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U213bar (
    .O(n7bar),
    .I0(n224bar),
    .I1(n225bar)
  );
  //OR U214
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U214 (
    .O(n225),
    .I0(n226),
    .I1(n227)
  );
  //AND U214bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U214bar (
    .O(n225bar),
    .I0(n226bar),
    .I1(n227bar)
  );
  //OR U215
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U215 (
    .O(n227),
    .I0(n228),
    .I1(n229)
  );
  //AND U215bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U215bar (
    .O(n227bar),
    .I0(n228bar),
    .I1(n229bar)
  );
  //OR U216
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U216 (
    .O(n229),
    .I0(in[136]),
    .I1(in[121])
  );
  //AND U216bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U216bar (
    .O(n229bar),
    .I0(inbar[136]),
    .I1(inbar[121])
  );
  //OR U217
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U217 (
    .O(n228),
    .I0(in[186]),
    .I1(in[174])
  );
  //AND U217bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U217bar (
    .O(n228bar),
    .I0(inbar[186]),
    .I1(inbar[174])
  );
  //OR U218
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U218 (
    .O(n226),
    .I0(n230),
    .I1(n231)
  );
  //AND U218bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U218bar (
    .O(n226bar),
    .I0(n230bar),
    .I1(n231bar)
  );
  //OR U219
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U219 (
    .O(n231),
    .I0(in[198]),
    .I1(in[197])
  );
  //AND U219bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U219bar (
    .O(n231bar),
    .I0(inbar[198]),
    .I1(inbar[197])
  );
  //OR U220
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U220 (
    .O(n230),
    .I0(in[214]),
    .I1(in[199])
  );
  //AND U220bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U220bar (
    .O(n230bar),
    .I0(inbar[214]),
    .I1(inbar[199])
  );
  //OR U221
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U221 (
    .O(n224),
    .I0(n232),
    .I1(n233)
  );
  //AND U221bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U221bar (
    .O(n224bar),
    .I0(n232bar),
    .I1(n233bar)
  );
  //OR U222
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U222 (
    .O(n233),
    .I0(n234),
    .I1(n235)
  );
  //AND U222bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U222bar (
    .O(n233bar),
    .I0(n234bar),
    .I1(n235bar)
  );
  //OR U223
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U223 (
    .O(n235),
    .I0(in[231]),
    .I1(in[220])
  );
  //AND U223bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U223bar (
    .O(n235bar),
    .I0(inbar[231]),
    .I1(inbar[220])
  );
  //OR U224
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U224 (
    .O(n234),
    .I0(in_25),
    .I1(in[245])
  );
  //AND U224bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U224bar (
    .O(n234bar),
    .I0(in_25bar),
    .I1(inbar[245])
  );
  //OR U225
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U225 (
    .O(n232),
    .I0(n236),
    .I1(n237)
  );
  //AND U225bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U225bar (
    .O(n232bar),
    .I0(n236bar),
    .I1(n237bar)
  );
  //OR U226
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U226 (
    .O(n237),
    .I0(in_53),
    .I1(in_29)
  );
  //AND U226bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U226bar (
    .O(n237bar),
    .I0(in_53bar),
    .I1(in_29bar)
  );
  //OR U227
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U227 (
    .O(n236),
    .I0(in_79),
    .I1(in_74)
  );
  //AND U227bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U227bar (
    .O(n236bar),
    .I0(in_79bar),
    .I1(in_74bar)
  );
  //OR U228
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U228 (
    .O(n184),
    .I0(n238),
    .I1(n239)
  );
  //AND U228bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U228bar (
    .O(n184bar),
    .I0(n238bar),
    .I1(n239bar)
  );
  //OR U229
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U229 (
    .O(n239),
    .I0(in[152]),
    .I1(in[140])
  );
  //AND U229bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U229bar (
    .O(n239bar),
    .I0(inbar[152]),
    .I1(inbar[140])
  );
  //OR U230
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U230 (
    .O(n238),
    .I0(in[155]),
    .I1(n240)
  );
  //AND U230bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U230bar (
    .O(n238bar),
    .I0(inbar[155]),
    .I1(n240bar)
  );
  //OR U231
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U231 (
    .O(n240),
    .I0(in[166]),
    .I1(in[165])
  );
  //AND U231bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U231bar (
    .O(n240bar),
    .I0(inbar[166]),
    .I1(inbar[165])
  );
  //OR U232
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U232 (
    .O(n182),
    .I0(n241),
    .I1(n242)
  );
  //AND U232bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U232bar (
    .O(n182bar),
    .I0(n241bar),
    .I1(n242bar)
  );
  //OR U233
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U233 (
    .O(n242),
    .I0(n243),
    .I1(n244)
  );
  //AND U233bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U233bar (
    .O(n242bar),
    .I0(n243bar),
    .I1(n244bar)
  );
  //OR U234
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U234 (
    .O(n244),
    .I0(in[202]),
    .I1(in[185])
  );
  //AND U234bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U234bar (
    .O(n244bar),
    .I0(inbar[202]),
    .I1(inbar[185])
  );
  //OR U235
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U235 (
    .O(n243),
    .I0(in[211]),
    .I1(n245)
  );
  //AND U235bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U235bar (
    .O(n243bar),
    .I0(inbar[211]),
    .I1(n245bar)
  );
  //OR U236
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U236 (
    .O(n245),
    .I0(in[255]),
    .I1(in[253])
  );
  //AND U236bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U236bar (
    .O(n245bar),
    .I0(inbar[255]),
    .I1(inbar[253])
  );
  //OR U237
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U237 (
    .O(n241),
    .I0(n246),
    .I1(n247)
  );
  //AND U237bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U237bar (
    .O(n241bar),
    .I0(n246bar),
    .I1(n247bar)
  );
  //OR U238
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U238 (
    .O(n247),
    .I0(in_35),
    .I1(in_15)
  );
  //AND U238bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U238bar (
    .O(n247bar),
    .I0(in_35bar),
    .I1(in_15bar)
  );
  //OR U239
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U239 (
    .O(n246),
    .I0(in_36),
    .I1(n248)
  );
  //AND U239bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U239bar (
    .O(n246bar),
    .I0(in_36bar),
    .I1(n248bar)
  );
  //OR U240
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U240 (
    .O(n248),
    .I0(in_48),
    .I1(in_40)
  );
  //AND U240bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U240bar (
    .O(n248bar),
    .I0(in_48bar),
    .I1(in_40bar)
  );
  //OR U241
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U241 (
    .O(out[1]),
    .I0(n249),
    .I1(n250)
  );
  //AND U241bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U241bar (
    .O(outbar[1]),
    .I0(n249bar),
    .I1(n250bar)
  );
  //OR U242
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U242 (
    .O(n250),
    .I0(n251),
    .I1(n252)
  );
  //AND U242bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U242bar (
    .O(n250bar),
    .I0(n251bar),
    .I1(n252bar)
  );
  //OR U243
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U243 (
    .O(n252),
    .I0(n253),
    .I1(n254)
  );
  //AND U243bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U243bar (
    .O(n252bar),
    .I0(n253bar),
    .I1(n254bar)
  );
  //OR U244
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U244 (
    .O(n254),
    .I0(n52),
    .I1(n86)
  );
  //AND U244bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U244bar (
    .O(n254bar),
    .I0(n52bar),
    .I1(n86bar)
  );
  //OR U245
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U245 (
    .O(n86),
    .I0(n255),
    .I1(n256)
  );
  //AND U245bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U245bar (
    .O(n86bar),
    .I0(n255bar),
    .I1(n256bar)
  );
  //OR U246
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U246 (
    .O(n256),
    .I0(n257),
    .I1(n258)
  );
  //AND U246bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U246bar (
    .O(n256bar),
    .I0(n257bar),
    .I1(n258bar)
  );
  //OR U247
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U247 (
    .O(n258),
    .I0(n259),
    .I1(n260)
  );
  //AND U247bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U247bar (
    .O(n258bar),
    .I0(n259bar),
    .I1(n260bar)
  );
  //OR U248
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U248 (
    .O(n260),
    .I0(in[116]),
    .I1(in[110])
  );
  //AND U248bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U248bar (
    .O(n260bar),
    .I0(inbar[116]),
    .I1(inbar[110])
  );
  //OR U249
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U249 (
    .O(n259),
    .I0(in[133]),
    .I1(in[130])
  );
  //AND U249bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U249bar (
    .O(n259bar),
    .I0(inbar[133]),
    .I1(inbar[130])
  );
  //OR U250
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U250 (
    .O(n257),
    .I0(n261),
    .I1(n262)
  );
  //AND U250bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U250bar (
    .O(n257bar),
    .I0(n261bar),
    .I1(n262bar)
  );
  //OR U251
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U251 (
    .O(n262),
    .I0(in[203]),
    .I1(in[135])
  );
  //AND U251bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U251bar (
    .O(n262bar),
    .I0(inbar[203]),
    .I1(inbar[135])
  );
  //OR U252
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U252 (
    .O(n261),
    .I0(in[232]),
    .I1(in[223])
  );
  //AND U252bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U252bar (
    .O(n261bar),
    .I0(inbar[232]),
    .I1(inbar[223])
  );
  //OR U253
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U253 (
    .O(n255),
    .I0(n263),
    .I1(n264)
  );
  //AND U253bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U253bar (
    .O(n255bar),
    .I0(n263bar),
    .I1(n264bar)
  );
  //OR U254
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U254 (
    .O(n264),
    .I0(n265),
    .I1(n266)
  );
  //AND U254bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U254bar (
    .O(n264bar),
    .I0(n265bar),
    .I1(n266bar)
  );
  //OR U255
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U255 (
    .O(n266),
    .I0(in[255]),
    .I1(in[233])
  );
  //AND U255bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U255bar (
    .O(n266bar),
    .I0(inbar[255]),
    .I1(inbar[233])
  );
  //OR U256
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U256 (
    .O(n265),
    .I0(in_53),
    .I1(in_34)
  );
  //AND U256bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U256bar (
    .O(n265bar),
    .I0(in_53bar),
    .I1(in_34bar)
  );
  //OR U257
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U257 (
    .O(n263),
    .I0(n267),
    .I1(n268)
  );
  //AND U257bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U257bar (
    .O(n263bar),
    .I0(n267bar),
    .I1(n268bar)
  );
  //OR U258
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U258 (
    .O(n268),
    .I0(in_57),
    .I1(in_55)
  );
  //AND U258bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U258bar (
    .O(n268bar),
    .I0(in_57bar),
    .I1(in_55bar)
  );
  //OR U259
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U259 (
    .O(n267),
    .I0(in_68),
    .I1(in_67)
  );
  //AND U259bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U259bar (
    .O(n267bar),
    .I0(in_68bar),
    .I1(in_67bar)
  );
  //OR U260
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U260 (
    .O(n52),
    .I0(n269),
    .I1(n270)
  );
  //AND U260bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U260bar (
    .O(n52bar),
    .I0(n269bar),
    .I1(n270bar)
  );
  //OR U261
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U261 (
    .O(n270),
    .I0(n271),
    .I1(n272)
  );
  //AND U261bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U261bar (
    .O(n270bar),
    .I0(n271bar),
    .I1(n272bar)
  );
  //OR U262
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U262 (
    .O(n272),
    .I0(n273),
    .I1(n274)
  );
  //AND U262bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U262bar (
    .O(n272bar),
    .I0(n273bar),
    .I1(n274bar)
  );
  //OR U263
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U263 (
    .O(n274),
    .I0(n29),
    .I1(n101)
  );
  //AND U263bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U263bar (
    .O(n274bar),
    .I0(n29bar),
    .I1(n101bar)
  );
  //OR U264
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U264 (
    .O(n101),
    .I0(n275),
    .I1(n276)
  );
  //AND U264bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U264bar (
    .O(n101bar),
    .I0(n275bar),
    .I1(n276bar)
  );
  //OR U265
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U265 (
    .O(n276),
    .I0(n277),
    .I1(n278)
  );
  //AND U265bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U265bar (
    .O(n276bar),
    .I0(n277bar),
    .I1(n278bar)
  );
  //OR U266
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U266 (
    .O(n278),
    .I0(n279),
    .I1(n280)
  );
  //AND U266bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U266bar (
    .O(n278bar),
    .I0(n279bar),
    .I1(n280bar)
  );
  //OR U267
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U267 (
    .O(n280),
    .I0(in[121]),
    .I1(in[102])
  );
  //AND U267bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U267bar (
    .O(n280bar),
    .I0(inbar[121]),
    .I1(inbar[102])
  );
  //OR U268
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U268 (
    .O(n279),
    .I0(in[162]),
    .I1(in[161])
  );
  //AND U268bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U268bar (
    .O(n279bar),
    .I0(inbar[162]),
    .I1(inbar[161])
  );
  //OR U269
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U269 (
    .O(n277),
    .I0(n281),
    .I1(n282)
  );
  //AND U269bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U269bar (
    .O(n277bar),
    .I0(n281bar),
    .I1(n282bar)
  );
  //OR U270
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U270 (
    .O(n282),
    .I0(in[192]),
    .I1(in[178])
  );
  //AND U270bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U270bar (
    .O(n282bar),
    .I0(inbar[192]),
    .I1(inbar[178])
  );
  //OR U271
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U271 (
    .O(n281),
    .I0(in[244]),
    .I1(in[209])
  );
  //AND U271bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U271bar (
    .O(n281bar),
    .I0(inbar[244]),
    .I1(inbar[209])
  );
  //OR U272
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U272 (
    .O(n275),
    .I0(n283),
    .I1(n284)
  );
  //AND U272bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U272bar (
    .O(n275bar),
    .I0(n283bar),
    .I1(n284bar)
  );
  //OR U273
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U273 (
    .O(n284),
    .I0(n285),
    .I1(n286)
  );
  //AND U273bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U273bar (
    .O(n284bar),
    .I0(n285bar),
    .I1(n286bar)
  );
  //OR U274
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U274 (
    .O(n286),
    .I0(in[90]),
    .I1(in[254])
  );
  //AND U274bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U274bar (
    .O(n286bar),
    .I0(inbar[90]),
    .I1(inbar[254])
  );
  //OR U275
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U275 (
    .O(n285),
    .I0(in_36),
    .I1(in_32)
  );
  //AND U275bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U275bar (
    .O(n285bar),
    .I0(in_36bar),
    .I1(in_32bar)
  );
  //OR U276
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U276 (
    .O(n283),
    .I0(n287),
    .I1(n288)
  );
  //AND U276bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U276bar (
    .O(n283bar),
    .I0(n287bar),
    .I1(n288bar)
  );
  //OR U277
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U277 (
    .O(n288),
    .I0(in_62),
    .I1(in_37)
  );
  //AND U277bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U277bar (
    .O(n288bar),
    .I0(in_62bar),
    .I1(in_37bar)
  );
  //OR U278
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U278 (
    .O(n287),
    .I0(in_75),
    .I1(in_73)
  );
  //AND U278bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U278bar (
    .O(n287bar),
    .I0(in_75bar),
    .I1(in_73bar)
  );
  //OR U279
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U279 (
    .O(n29),
    .I0(n289),
    .I1(n290)
  );
  //AND U279bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U279bar (
    .O(n29bar),
    .I0(n289bar),
    .I1(n290bar)
  );
  //OR U280
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U280 (
    .O(n290),
    .I0(n291),
    .I1(n292)
  );
  //AND U280bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U280bar (
    .O(n290bar),
    .I0(n291bar),
    .I1(n292bar)
  );
  //OR U281
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U281 (
    .O(n292),
    .I0(n293),
    .I1(n294)
  );
  //AND U281bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U281bar (
    .O(n292bar),
    .I0(n293bar),
    .I1(n294bar)
  );
  //OR U282
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U282 (
    .O(n294),
    .I0(in[171]),
    .I1(in[153])
  );
  //AND U282bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U282bar (
    .O(n294bar),
    .I0(inbar[171]),
    .I1(inbar[153])
  );
  //OR U283
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U283 (
    .O(n293),
    .I0(in[187]),
    .I1(in[176])
  );
  //AND U283bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U283bar (
    .O(n293bar),
    .I0(inbar[187]),
    .I1(inbar[176])
  );
  //OR U284
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U284 (
    .O(n291),
    .I0(n295),
    .I1(n296)
  );
  //AND U284bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U284bar (
    .O(n291bar),
    .I0(n295bar),
    .I1(n296bar)
  );
  //OR U285
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U285 (
    .O(n296),
    .I0(in[245]),
    .I1(in[211])
  );
  //AND U285bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U285bar (
    .O(n296bar),
    .I0(inbar[245]),
    .I1(inbar[211])
  );
  //OR U286
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U286 (
    .O(n295),
    .I0(in[97]),
    .I1(in[88])
  );
  //AND U286bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U286bar (
    .O(n295bar),
    .I0(inbar[97]),
    .I1(inbar[88])
  );
  //OR U287
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U287 (
    .O(n289),
    .I0(n297),
    .I1(n298)
  );
  //AND U287bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U287bar (
    .O(n289bar),
    .I0(n297bar),
    .I1(n298bar)
  );
  //OR U288
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U288 (
    .O(n298),
    .I0(n299),
    .I1(n300)
  );
  //AND U288bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U288bar (
    .O(n298bar),
    .I0(n299bar),
    .I1(n300bar)
  );
  //OR U289
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U289 (
    .O(n300),
    .I0(in_10),
    .I1(in_0)
  );
  //AND U289bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U289bar (
    .O(n300bar),
    .I0(in_10bar),
    .I1(in_0bar)
  );
  //OR U290
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U290 (
    .O(n299),
    .I0(in_59),
    .I1(in_5)
  );
  //AND U290bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U290bar (
    .O(n299bar),
    .I0(in_59bar),
    .I1(in_5bar)
  );
  //OR U291
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U291 (
    .O(n297),
    .I0(n301),
    .I1(n302)
  );
  //AND U291bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U291bar (
    .O(n297bar),
    .I0(n301bar),
    .I1(n302bar)
  );
  //OR U292
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U292 (
    .O(n302),
    .I0(in_60),
    .I1(in_6)
  );
  //AND U292bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U292bar (
    .O(n302bar),
    .I0(in_60bar),
    .I1(in_6bar)
  );
  //OR U293
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U293 (
    .O(n301),
    .I0(in_77),
    .I1(in_69)
  );
  //AND U293bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U293bar (
    .O(n301bar),
    .I0(in_77bar),
    .I1(in_69bar)
  );
  //OR U294
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U294 (
    .O(n273),
    .I0(in[113]),
    .I1(n109)
  );
  //AND U294bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U294bar (
    .O(n273bar),
    .I0(inbar[113]),
    .I1(n109bar)
  );
  //OR U295
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U295 (
    .O(n109),
    .I0(n303),
    .I1(n304)
  );
  //AND U295bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U295bar (
    .O(n109bar),
    .I0(n303bar),
    .I1(n304bar)
  );
  //OR U296
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U296 (
    .O(n304),
    .I0(n305),
    .I1(n306)
  );
  //AND U296bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U296bar (
    .O(n304bar),
    .I0(n305bar),
    .I1(n306bar)
  );
  //OR U297
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U297 (
    .O(n306),
    .I0(n307),
    .I1(n308)
  );
  //AND U297bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U297bar (
    .O(n306bar),
    .I0(n307bar),
    .I1(n308bar)
  );
  //OR U298
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U298 (
    .O(n308),
    .I0(in[125]),
    .I1(in[107])
  );
  //AND U298bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U298bar (
    .O(n308bar),
    .I0(inbar[125]),
    .I1(inbar[107])
  );
  //OR U299
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U299 (
    .O(n307),
    .I0(in[138]),
    .I1(in[126])
  );
  //AND U299bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U299bar (
    .O(n307bar),
    .I0(inbar[138]),
    .I1(inbar[126])
  );
  //OR U300
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U300 (
    .O(n305),
    .I0(n309),
    .I1(n310)
  );
  //AND U300bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U300bar (
    .O(n305bar),
    .I0(n309bar),
    .I1(n310bar)
  );
  //OR U301
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U301 (
    .O(n310),
    .I0(in[189]),
    .I1(in[143])
  );
  //AND U301bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U301bar (
    .O(n310bar),
    .I0(inbar[189]),
    .I1(inbar[143])
  );
  //OR U302
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U302 (
    .O(n309),
    .I0(in[99]),
    .I1(in[214])
  );
  //AND U302bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U302bar (
    .O(n309bar),
    .I0(inbar[99]),
    .I1(inbar[214])
  );
  //OR U303
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U303 (
    .O(n303),
    .I0(n311),
    .I1(n312)
  );
  //AND U303bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U303bar (
    .O(n303bar),
    .I0(n311bar),
    .I1(n312bar)
  );
  //OR U304
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U304 (
    .O(n312),
    .I0(n313),
    .I1(n314)
  );
  //AND U304bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U304bar (
    .O(n312bar),
    .I0(n313bar),
    .I1(n314bar)
  );
  //OR U305
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U305 (
    .O(n314),
    .I0(in_15),
    .I1(in_12)
  );
  //AND U305bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U305bar (
    .O(n314bar),
    .I0(in_15bar),
    .I1(in_12bar)
  );
  //OR U306
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U306 (
    .O(n313),
    .I0(in_20),
    .I1(in_2)
  );
  //AND U306bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U306bar (
    .O(n313bar),
    .I0(in_20bar),
    .I1(in_2bar)
  );
  //OR U307
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U307 (
    .O(n311),
    .I0(n315),
    .I1(n316)
  );
  //AND U307bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U307bar (
    .O(n311bar),
    .I0(n315bar),
    .I1(n316bar)
  );
  //OR U308
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U308 (
    .O(n316),
    .I0(in_30),
    .I1(in_3)
  );
  //AND U308bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U308bar (
    .O(n316bar),
    .I0(in_30bar),
    .I1(in_3bar)
  );
  //OR U309
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U309 (
    .O(n315),
    .I0(in_4),
    .I1(in_38)
  );
  //AND U309bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U309bar (
    .O(n315bar),
    .I0(in_4bar),
    .I1(in_38bar)
  );
  //OR U310
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U310 (
    .O(n271),
    .I0(n317),
    .I1(n318)
  );
  //AND U310bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U310bar (
    .O(n271bar),
    .I0(n317bar),
    .I1(n318bar)
  );
  //OR U311
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U311 (
    .O(n318),
    .I0(in[148]),
    .I1(in[137])
  );
  //AND U311bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U311bar (
    .O(n318bar),
    .I0(inbar[148]),
    .I1(inbar[137])
  );
  //OR U312
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U312 (
    .O(n317),
    .I0(in[149]),
    .I1(n319)
  );
  //AND U312bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U312bar (
    .O(n317bar),
    .I0(inbar[149]),
    .I1(n319bar)
  );
  //OR U313
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U313 (
    .O(n319),
    .I0(in[195]),
    .I1(in[190])
  );
  //AND U313bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U313bar (
    .O(n319bar),
    .I0(inbar[195]),
    .I1(inbar[190])
  );
  //OR U314
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U314 (
    .O(n269),
    .I0(n320),
    .I1(n321)
  );
  //AND U314bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U314bar (
    .O(n269bar),
    .I0(n320bar),
    .I1(n321bar)
  );
  //OR U315
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U315 (
    .O(n321),
    .I0(n322),
    .I1(n323)
  );
  //AND U315bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U315bar (
    .O(n321bar),
    .I0(n322bar),
    .I1(n323bar)
  );
  //OR U316
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U316 (
    .O(n323),
    .I0(in[98]),
    .I1(in[197])
  );
  //AND U316bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U316bar (
    .O(n323bar),
    .I0(inbar[98]),
    .I1(inbar[197])
  );
  //OR U317
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U317 (
    .O(n322),
    .I0(in_11),
    .I1(n324)
  );
  //AND U317bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U317bar (
    .O(n322bar),
    .I0(in_11bar),
    .I1(n324bar)
  );
  //OR U318
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U318 (
    .O(n324),
    .I0(in_26),
    .I1(in_14)
  );
  //AND U318bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U318bar (
    .O(n324bar),
    .I0(in_26bar),
    .I1(in_14bar)
  );
  //OR U319
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U319 (
    .O(n320),
    .I0(n325),
    .I1(n326)
  );
  //AND U319bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U319bar (
    .O(n320bar),
    .I0(n325bar),
    .I1(n326bar)
  );
  //OR U320
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U320 (
    .O(n326),
    .I0(in_35),
    .I1(in_27)
  );
  //AND U320bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U320bar (
    .O(n326bar),
    .I0(in_35bar),
    .I1(in_27bar)
  );
  //OR U321
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U321 (
    .O(n325),
    .I0(in_50),
    .I1(n327)
  );
  //AND U321bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U321bar (
    .O(n325bar),
    .I0(in_50bar),
    .I1(n327bar)
  );
  //OR U322
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U322 (
    .O(n327),
    .I0(in_78),
    .I1(in_61)
  );
  //AND U322bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U322bar (
    .O(n327bar),
    .I0(in_78bar),
    .I1(in_61bar)
  );
  //OR U323
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U323 (
    .O(n253),
    .I0(n31),
    .I1(n328)
  );
  //AND U323bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U323bar (
    .O(n253bar),
    .I0(n31bar),
    .I1(n328bar)
  );
  //OR U324
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U324 (
    .O(n328),
    .I0(in[106]),
    .I1(n110)
  );
  //AND U324bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U324bar (
    .O(n328bar),
    .I0(inbar[106]),
    .I1(n110bar)
  );
  //OR U325
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U325 (
    .O(n110),
    .I0(n329),
    .I1(n330)
  );
  //AND U325bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U325bar (
    .O(n110bar),
    .I0(n329bar),
    .I1(n330bar)
  );
  //OR U326
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U326 (
    .O(n330),
    .I0(n331),
    .I1(n332)
  );
  //AND U326bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U326bar (
    .O(n330bar),
    .I0(n331bar),
    .I1(n332bar)
  );
  //OR U327
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U327 (
    .O(n332),
    .I0(n333),
    .I1(n334)
  );
  //AND U327bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U327bar (
    .O(n332bar),
    .I0(n333bar),
    .I1(n334bar)
  );
  //OR U328
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U328 (
    .O(n334),
    .I0(in[127]),
    .I1(in[122])
  );
  //AND U328bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U328bar (
    .O(n334bar),
    .I0(inbar[127]),
    .I1(inbar[122])
  );
  //OR U329
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U329 (
    .O(n333),
    .I0(in[156]),
    .I1(in[132])
  );
  //AND U329bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U329bar (
    .O(n333bar),
    .I0(inbar[156]),
    .I1(inbar[132])
  );
  //OR U330
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U330 (
    .O(n331),
    .I0(n335),
    .I1(n336)
  );
  //AND U330bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U330bar (
    .O(n331bar),
    .I0(n335bar),
    .I1(n336bar)
  );
  //OR U331
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U331 (
    .O(n336),
    .I0(in[159]),
    .I1(in[157])
  );
  //AND U331bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U331bar (
    .O(n336bar),
    .I0(inbar[159]),
    .I1(inbar[157])
  );
  //OR U332
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U332 (
    .O(n335),
    .I0(in[185]),
    .I1(in[169])
  );
  //AND U332bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U332bar (
    .O(n335bar),
    .I0(inbar[185]),
    .I1(inbar[169])
  );
  //OR U333
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U333 (
    .O(n329),
    .I0(n337),
    .I1(n338)
  );
  //AND U333bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U333bar (
    .O(n329bar),
    .I0(n337bar),
    .I1(n338bar)
  );
  //OR U334
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U334 (
    .O(n338),
    .I0(n339),
    .I1(n340)
  );
  //AND U334bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U334bar (
    .O(n338bar),
    .I0(n339bar),
    .I1(n340bar)
  );
  //OR U335
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U335 (
    .O(n340),
    .I0(in[239]),
    .I1(in[218])
  );
  //AND U335bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U335bar (
    .O(n340bar),
    .I0(inbar[239]),
    .I1(inbar[218])
  );
  //OR U336
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U336 (
    .O(n339),
    .I0(in_13),
    .I1(in[87])
  );
  //AND U336bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U336bar (
    .O(n339bar),
    .I0(in_13bar),
    .I1(inbar[87])
  );
  //OR U337
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U337 (
    .O(n337),
    .I0(n341),
    .I1(n342)
  );
  //AND U337bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U337bar (
    .O(n337bar),
    .I0(n341bar),
    .I1(n342bar)
  );
  //OR U338
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U338 (
    .O(n342),
    .I0(in_72),
    .I1(in_70)
  );
  //AND U338bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U338bar (
    .O(n342bar),
    .I0(in_72bar),
    .I1(in_70bar)
  );
  //OR U339
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U339 (
    .O(n341),
    .I0(in_80),
    .I1(in_74)
  );
  //AND U339bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U339bar (
    .O(n341bar),
    .I0(in_80bar),
    .I1(in_74bar)
  );
  //OR U340
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U340 (
    .O(n31),
    .I0(n343),
    .I1(n344)
  );
  //AND U340bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U340bar (
    .O(n31bar),
    .I0(n343bar),
    .I1(n344bar)
  );
  //OR U341
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U341 (
    .O(n344),
    .I0(n345),
    .I1(n346)
  );
  //AND U341bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U341bar (
    .O(n344bar),
    .I0(n345bar),
    .I1(n346bar)
  );
  //OR U342
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U342 (
    .O(n346),
    .I0(n347),
    .I1(n348)
  );
  //AND U342bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U342bar (
    .O(n346bar),
    .I0(n347bar),
    .I1(n348bar)
  );
  //OR U343
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U343 (
    .O(n348),
    .I0(in[146]),
    .I1(in[100])
  );
  //AND U343bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U343bar (
    .O(n348bar),
    .I0(inbar[146]),
    .I1(inbar[100])
  );
  //OR U344
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U344 (
    .O(n347),
    .I0(in[168]),
    .I1(in[152])
  );
  //AND U344bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U344bar (
    .O(n347bar),
    .I0(inbar[168]),
    .I1(inbar[152])
  );
  //OR U345
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U345 (
    .O(n345),
    .I0(n349),
    .I1(n350)
  );
  //AND U345bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U345bar (
    .O(n345bar),
    .I0(n349bar),
    .I1(n350bar)
  );
  //OR U346
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U346 (
    .O(n350),
    .I0(in[199]),
    .I1(in[182])
  );
  //AND U346bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U346bar (
    .O(n350bar),
    .I0(inbar[199]),
    .I1(inbar[182])
  );
  //OR U347
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U347 (
    .O(n349),
    .I0(in[236]),
    .I1(in[204])
  );
  //AND U347bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U347bar (
    .O(n349bar),
    .I0(inbar[236]),
    .I1(inbar[204])
  );
  //OR U348
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U348 (
    .O(n343),
    .I0(n351),
    .I1(n352)
  );
  //AND U348bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U348bar (
    .O(n343bar),
    .I0(n351bar),
    .I1(n352bar)
  );
  //OR U349
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U349 (
    .O(n352),
    .I0(n353),
    .I1(n354)
  );
  //AND U349bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U349bar (
    .O(n352bar),
    .I0(n353bar),
    .I1(n354bar)
  );
  //OR U350
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U350 (
    .O(n354),
    .I0(in[89]),
    .I1(in[246])
  );
  //AND U350bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U350bar (
    .O(n354bar),
    .I0(inbar[89]),
    .I1(inbar[246])
  );
  //OR U351
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U351 (
    .O(n353),
    .I0(in[95]),
    .I1(in[92])
  );
  //AND U351bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U351bar (
    .O(n353bar),
    .I0(inbar[95]),
    .I1(inbar[92])
  );
  //OR U352
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U352 (
    .O(n351),
    .I0(n355),
    .I1(n356)
  );
  //AND U352bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U352bar (
    .O(n351bar),
    .I0(n355bar),
    .I1(n356bar)
  );
  //OR U353
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U353 (
    .O(n356),
    .I0(in_22),
    .I1(in_16)
  );
  //AND U353bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U353bar (
    .O(n356bar),
    .I0(in_22bar),
    .I1(in_16bar)
  );
  //OR U354
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U354 (
    .O(n355),
    .I0(in_51),
    .I1(in_49)
  );
  //AND U354bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U354bar (
    .O(n355bar),
    .I0(in_51bar),
    .I1(in_49bar)
  );
  //OR U355
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U355 (
    .O(n251),
    .I0(n357),
    .I1(n358)
  );
  //AND U355bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U355bar (
    .O(n251bar),
    .I0(n357bar),
    .I1(n358bar)
  );
  //OR U356
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U356 (
    .O(n358),
    .I0(in[158]),
    .I1(in[115])
  );
  //AND U356bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U356bar (
    .O(n358bar),
    .I0(inbar[158]),
    .I1(inbar[115])
  );
  //OR U357
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U357 (
    .O(n357),
    .I0(in[163]),
    .I1(n359)
  );
  //AND U357bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U357bar (
    .O(n357bar),
    .I0(inbar[163]),
    .I1(n359bar)
  );
  //OR U358
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U358 (
    .O(n359),
    .I0(in[206]),
    .I1(in[165])
  );
  //AND U358bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U358bar (
    .O(n359bar),
    .I0(inbar[206]),
    .I1(inbar[165])
  );
  //OR U359
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U359 (
    .O(n249),
    .I0(n360),
    .I1(n361)
  );
  //AND U359bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U359bar (
    .O(n249bar),
    .I0(n360bar),
    .I1(n361bar)
  );
  //OR U360
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U360 (
    .O(n361),
    .I0(n362),
    .I1(n363)
  );
  //AND U360bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U360bar (
    .O(n361bar),
    .I0(n362bar),
    .I1(n363bar)
  );
  //OR U361
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U361 (
    .O(n363),
    .I0(in[213]),
    .I1(in[207])
  );
  //AND U361bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U361bar (
    .O(n363bar),
    .I0(inbar[213]),
    .I1(inbar[207])
  );
  //OR U362
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U362 (
    .O(n362),
    .I0(in[215]),
    .I1(n364)
  );
  //AND U362bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U362bar (
    .O(n362bar),
    .I0(inbar[215]),
    .I1(n364bar)
  );
  //OR U363
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U363 (
    .O(n364),
    .I0(in[230]),
    .I1(in[220])
  );
  //AND U363bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U363bar (
    .O(n364bar),
    .I0(inbar[230]),
    .I1(inbar[220])
  );
  //OR U364
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U364 (
    .O(n360),
    .I0(n365),
    .I1(n366)
  );
  //AND U364bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U364bar (
    .O(n360bar),
    .I0(n365bar),
    .I1(n366bar)
  );
  //OR U365
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U365 (
    .O(n366),
    .I0(in[251]),
    .I1(in[234])
  );
  //AND U365bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U365bar (
    .O(n366bar),
    .I0(inbar[251]),
    .I1(inbar[234])
  );
  //OR U366
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U366 (
    .O(n365),
    .I0(in_17),
    .I1(n367)
  );
  //AND U366bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U366bar (
    .O(n365bar),
    .I0(in_17bar),
    .I1(n367bar)
  );
  //OR U367
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U367 (
    .O(n367),
    .I0(in_65),
    .I1(in_56)
  );
  //AND U367bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U367bar (
    .O(n367bar),
    .I0(in_65bar),
    .I1(in_56bar)
  );
  //OR U368
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U368 (
    .O(out[0]),
    .I0(n368),
    .I1(n369)
  );
  //AND U368bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U368bar (
    .O(outbar[0]),
    .I0(n368bar),
    .I1(n369bar)
  );
  //OR U369
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U369 (
    .O(n369),
    .I0(n370),
    .I1(n371)
  );
  //AND U369bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U369bar (
    .O(n369bar),
    .I0(n370bar),
    .I1(n371bar)
  );
  //OR U370
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U370 (
    .O(n371),
    .I0(n372),
    .I1(n373)
  );
  //AND U370bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U370bar (
    .O(n371bar),
    .I0(n372bar),
    .I1(n373bar)
  );
  //OR U371
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U371 (
    .O(n373),
    .I0(n153),
    .I1(n188)
  );
  //AND U371bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U371bar (
    .O(n373bar),
    .I0(n153bar),
    .I1(n188bar)
  );
  //OR U372
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U372 (
    .O(n188),
    .I0(n374),
    .I1(n375)
  );
  //AND U372bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U372bar (
    .O(n188bar),
    .I0(n374bar),
    .I1(n375bar)
  );
  //OR U373
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U373 (
    .O(n375),
    .I0(n376),
    .I1(n377)
  );
  //AND U373bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U373bar (
    .O(n375bar),
    .I0(n376bar),
    .I1(n377bar)
  );
  //OR U374
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U374 (
    .O(n377),
    .I0(n378),
    .I1(n379)
  );
  //AND U374bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U374bar (
    .O(n377bar),
    .I0(n378bar),
    .I1(n379bar)
  );
  //OR U375
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U375 (
    .O(n379),
    .I0(in[135]),
    .I1(in[104])
  );
  //AND U375bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U375bar (
    .O(n379bar),
    .I0(inbar[135]),
    .I1(inbar[104])
  );
  //OR U376
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U376 (
    .O(n378),
    .I0(in[188]),
    .I1(in[178])
  );
  //AND U376bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U376bar (
    .O(n378bar),
    .I0(inbar[188]),
    .I1(inbar[178])
  );
  //OR U377
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U377 (
    .O(n376),
    .I0(n380),
    .I1(n381)
  );
  //AND U377bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U377bar (
    .O(n376bar),
    .I0(n380bar),
    .I1(n381bar)
  );
  //OR U378
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U378 (
    .O(n381),
    .I0(in[217]),
    .I1(in[194])
  );
  //AND U378bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U378bar (
    .O(n381bar),
    .I0(inbar[217]),
    .I1(inbar[194])
  );
  //OR U379
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U379 (
    .O(n380),
    .I0(in[237]),
    .I1(in[218])
  );
  //AND U379bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U379bar (
    .O(n380bar),
    .I0(inbar[237]),
    .I1(inbar[218])
  );
  //OR U380
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U380 (
    .O(n374),
    .I0(n382),
    .I1(n383)
  );
  //AND U380bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U380bar (
    .O(n374bar),
    .I0(n382bar),
    .I1(n383bar)
  );
  //OR U381
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U381 (
    .O(n383),
    .I0(n384),
    .I1(n385)
  );
  //AND U381bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U381bar (
    .O(n383bar),
    .I0(n384bar),
    .I1(n385bar)
  );
  //OR U382
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U382 (
    .O(n385),
    .I0(in_2),
    .I1(in_10)
  );
  //AND U382bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U382bar (
    .O(n385bar),
    .I0(in_2bar),
    .I1(in_10bar)
  );
  //OR U383
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U383 (
    .O(n384),
    .I0(in_47),
    .I1(in_22)
  );
  //AND U383bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U383bar (
    .O(n384bar),
    .I0(in_47bar),
    .I1(in_22bar)
  );
  //OR U384
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U384 (
    .O(n382),
    .I0(n386),
    .I1(n387)
  );
  //AND U384bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U384bar (
    .O(n382bar),
    .I0(n386bar),
    .I1(n387bar)
  );
  //OR U385
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U385 (
    .O(n387),
    .I0(in_56),
    .I1(in_54)
  );
  //AND U385bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U385bar (
    .O(n387bar),
    .I0(in_56bar),
    .I1(in_54bar)
  );
  //OR U386
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U386 (
    .O(n386),
    .I0(in_63),
    .I1(in_61)
  );
  //AND U386bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U386bar (
    .O(n386bar),
    .I0(in_63bar),
    .I1(in_61bar)
  );
  //OR U387
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U387 (
    .O(n153),
    .I0(n388),
    .I1(n389)
  );
  //AND U387bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U387bar (
    .O(n153bar),
    .I0(n388bar),
    .I1(n389bar)
  );
  //OR U388
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U388 (
    .O(n389),
    .I0(n390),
    .I1(n391)
  );
  //AND U388bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U388bar (
    .O(n389bar),
    .I0(n390bar),
    .I1(n391bar)
  );
  //OR U389
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U389 (
    .O(n391),
    .I0(n392),
    .I1(n393)
  );
  //AND U389bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U389bar (
    .O(n391bar),
    .I0(n392bar),
    .I1(n393bar)
  );
  //OR U390
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U390 (
    .O(n393),
    .I0(in[158]),
    .I1(in[142])
  );
  //AND U390bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U390bar (
    .O(n393bar),
    .I0(inbar[158]),
    .I1(inbar[142])
  );
  //OR U391
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U391 (
    .O(n392),
    .I0(in[175]),
    .I1(in[164])
  );
  //AND U391bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U391bar (
    .O(n392bar),
    .I0(inbar[175]),
    .I1(inbar[164])
  );
  //OR U392
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U392 (
    .O(n390),
    .I0(n394),
    .I1(n395)
  );
  //AND U392bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U392bar (
    .O(n390bar),
    .I0(n394bar),
    .I1(n395bar)
  );
  //OR U393
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U393 (
    .O(n395),
    .I0(in[228]),
    .I1(in[204])
  );
  //AND U393bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U393bar (
    .O(n395bar),
    .I0(inbar[228]),
    .I1(inbar[204])
  );
  //OR U394
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U394 (
    .O(n394),
    .I0(in[91]),
    .I1(in[87])
  );
  //AND U394bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U394bar (
    .O(n394bar),
    .I0(inbar[91]),
    .I1(inbar[87])
  );
  //OR U395
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U395 (
    .O(n388),
    .I0(n396),
    .I1(n397)
  );
  //AND U395bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U395bar (
    .O(n388bar),
    .I0(n396bar),
    .I1(n397bar)
  );
  //OR U396
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U396 (
    .O(n397),
    .I0(n398),
    .I1(n399)
  );
  //AND U396bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U396bar (
    .O(n397bar),
    .I0(n398bar),
    .I1(n399bar)
  );
  //OR U397
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U397 (
    .O(n399),
    .I0(in_21),
    .I1(in_11)
  );
  //AND U397bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U397bar (
    .O(n399bar),
    .I0(in_21bar),
    .I1(in_11bar)
  );
  //OR U398
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U398 (
    .O(n398),
    .I0(in_5),
    .I1(in_3)
  );
  //AND U398bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U398bar (
    .O(n398bar),
    .I0(in_5bar),
    .I1(in_3bar)
  );
  //OR U399
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U399 (
    .O(n396),
    .I0(n400),
    .I1(n401)
  );
  //AND U399bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U399bar (
    .O(n396bar),
    .I0(n400bar),
    .I1(n401bar)
  );
  //OR U400
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U400 (
    .O(n401),
    .I0(in_68),
    .I1(in_64)
  );
  //AND U400bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U400bar (
    .O(n401bar),
    .I0(in_68bar),
    .I1(in_64bar)
  );
  //OR U401
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U401 (
    .O(n400),
    .I0(in_76),
    .I1(in_73)
  );
  //AND U401bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U401bar (
    .O(n400bar),
    .I0(in_76bar),
    .I1(in_73bar)
  );
  //OR U402
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U402 (
    .O(n372),
    .I0(n195),
    .I1(n402)
  );
  //AND U402bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U402bar (
    .O(n372bar),
    .I0(n195bar),
    .I1(n402bar)
  );
  //OR U403
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U403 (
    .O(n402),
    .I0(in[100]),
    .I1(n8)
  );
  //AND U403bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U403bar (
    .O(n402bar),
    .I0(inbar[100]),
    .I1(n8bar)
  );
  //OR U404
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U404 (
    .O(n8),
    .I0(n403),
    .I1(n404)
  );
  //AND U404bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U404bar (
    .O(n8bar),
    .I0(n403bar),
    .I1(n404bar)
  );
  //OR U405
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U405 (
    .O(n404),
    .I0(n405),
    .I1(n406)
  );
  //AND U405bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U405bar (
    .O(n404bar),
    .I0(n405bar),
    .I1(n406bar)
  );
  //OR U406
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U406 (
    .O(n406),
    .I0(n407),
    .I1(n408)
  );
  //AND U406bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U406bar (
    .O(n406bar),
    .I0(n407bar),
    .I1(n408bar)
  );
  //OR U407
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U407 (
    .O(n408),
    .I0(n156),
    .I1(n223)
  );
  //AND U407bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U407bar (
    .O(n408bar),
    .I0(n156bar),
    .I1(n223bar)
  );
  //OR U408
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U408 (
    .O(n223),
    .I0(n409),
    .I1(n410)
  );
  //AND U408bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U408bar (
    .O(n223bar),
    .I0(n409bar),
    .I1(n410bar)
  );
  //OR U409
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U409 (
    .O(n410),
    .I0(n411),
    .I1(n412)
  );
  //AND U409bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U409bar (
    .O(n410bar),
    .I0(n411bar),
    .I1(n412bar)
  );
  //OR U410
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U410 (
    .O(n412),
    .I0(n413),
    .I1(n414)
  );
  //AND U410bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U410bar (
    .O(n412bar),
    .I0(n413bar),
    .I1(n414bar)
  );
  //OR U411
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U411 (
    .O(n414),
    .I0(in[119]),
    .I1(in[103])
  );
  //AND U411bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U411bar (
    .O(n414bar),
    .I0(inbar[119]),
    .I1(inbar[103])
  );
  //OR U412
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U412 (
    .O(n413),
    .I0(in[137]),
    .I1(in[133])
  );
  //AND U412bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U412bar (
    .O(n413bar),
    .I0(inbar[137]),
    .I1(inbar[133])
  );
  //OR U413
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U413 (
    .O(n411),
    .I0(n415),
    .I1(n416)
  );
  //AND U413bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U413bar (
    .O(n411bar),
    .I0(n415bar),
    .I1(n416bar)
  );
  //OR U414
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U414 (
    .O(n416),
    .I0(in[176]),
    .I1(in[173])
  );
  //AND U414bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U414bar (
    .O(n416bar),
    .I0(inbar[176]),
    .I1(inbar[173])
  );
  //OR U415
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U415 (
    .O(n415),
    .I0(in[210]),
    .I1(in[181])
  );
  //AND U415bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U415bar (
    .O(n415bar),
    .I0(inbar[210]),
    .I1(inbar[181])
  );
  //OR U416
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U416 (
    .O(n409),
    .I0(n417),
    .I1(n418)
  );
  //AND U416bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U416bar (
    .O(n409bar),
    .I0(n417bar),
    .I1(n418bar)
  );
  //OR U417
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U417 (
    .O(n418),
    .I0(n419),
    .I1(n420)
  );
  //AND U417bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U417bar (
    .O(n418bar),
    .I0(n419bar),
    .I1(n420bar)
  );
  //OR U418
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U418 (
    .O(n420),
    .I0(in_13),
    .I1(in[234])
  );
  //AND U418bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U418bar (
    .O(n420bar),
    .I0(in_13bar),
    .I1(inbar[234])
  );
  //OR U419
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U419 (
    .O(n419),
    .I0(in_38),
    .I1(in_32)
  );
  //AND U419bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U419bar (
    .O(n419bar),
    .I0(in_38bar),
    .I1(in_32bar)
  );
  //OR U420
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U420 (
    .O(n417),
    .I0(n421),
    .I1(n422)
  );
  //AND U420bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U420bar (
    .O(n417bar),
    .I0(n421bar),
    .I1(n422bar)
  );
  //OR U421
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U421 (
    .O(n422),
    .I0(in_42),
    .I1(in_41)
  );
  //AND U421bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U421bar (
    .O(n422bar),
    .I0(in_42bar),
    .I1(in_41bar)
  );
  //OR U422
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U422 (
    .O(n421),
    .I0(in_7),
    .I1(in_49)
  );
  //AND U422bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U422bar (
    .O(n421bar),
    .I0(in_7bar),
    .I1(in_49bar)
  );
  //OR U423
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U423 (
    .O(n156),
    .I0(n423),
    .I1(n424)
  );
  //AND U423bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U423bar (
    .O(n156bar),
    .I0(n423bar),
    .I1(n424bar)
  );
  //OR U424
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U424 (
    .O(n424),
    .I0(n425),
    .I1(n426)
  );
  //AND U424bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U424bar (
    .O(n424bar),
    .I0(n425bar),
    .I1(n426bar)
  );
  //OR U425
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U425 (
    .O(n426),
    .I0(n427),
    .I1(n428)
  );
  //AND U425bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U425bar (
    .O(n426bar),
    .I0(n427bar),
    .I1(n428bar)
  );
  //OR U426
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U426 (
    .O(n428),
    .I0(in[159]),
    .I1(in[105])
  );
  //AND U426bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U426bar (
    .O(n428bar),
    .I0(inbar[159]),
    .I1(inbar[105])
  );
  //OR U427
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U427 (
    .O(n427),
    .I0(in[206]),
    .I1(in[183])
  );
  //AND U427bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U427bar (
    .O(n427bar),
    .I0(inbar[206]),
    .I1(inbar[183])
  );
  //OR U428
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U428 (
    .O(n425),
    .I0(n429),
    .I1(n430)
  );
  //AND U428bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U428bar (
    .O(n425bar),
    .I0(n429bar),
    .I1(n430bar)
  );
  //OR U429
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U429 (
    .O(n430),
    .I0(in[229]),
    .I1(in[219])
  );
  //AND U429bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U429bar (
    .O(n430bar),
    .I0(inbar[229]),
    .I1(inbar[219])
  );
  //OR U430
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U430 (
    .O(n429),
    .I0(in[235]),
    .I1(in[232])
  );
  //AND U430bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U430bar (
    .O(n429bar),
    .I0(inbar[235]),
    .I1(inbar[232])
  );
  //OR U431
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U431 (
    .O(n423),
    .I0(n431),
    .I1(n432)
  );
  //AND U431bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U431bar (
    .O(n423bar),
    .I0(n431bar),
    .I1(n432bar)
  );
  //OR U432
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U432 (
    .O(n432),
    .I0(n433),
    .I1(n434)
  );
  //AND U432bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U432bar (
    .O(n432bar),
    .I0(n433bar),
    .I1(n434bar)
  );
  //OR U433
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U433 (
    .O(n434),
    .I0(in[249]),
    .I1(in[242])
  );
  //AND U433bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U433bar (
    .O(n434bar),
    .I0(inbar[249]),
    .I1(inbar[242])
  );
  //OR U434
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U434 (
    .O(n433),
    .I0(in[89]),
    .I1(in[254])
  );
  //AND U434bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U434bar (
    .O(n433bar),
    .I0(inbar[89]),
    .I1(inbar[254])
  );
  //OR U435
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U435 (
    .O(n431),
    .I0(n435),
    .I1(n436)
  );
  //AND U435bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U435bar (
    .O(n431bar),
    .I0(n435bar),
    .I1(n436bar)
  );
  //OR U436
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U436 (
    .O(n436),
    .I0(in_14),
    .I1(in[99])
  );
  //AND U436bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U436bar (
    .O(n436bar),
    .I0(in_14bar),
    .I1(inbar[99])
  );
  //OR U437
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U437 (
    .O(n435),
    .I0(in_60),
    .I1(in_18)
  );
  //AND U437bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U437bar (
    .O(n435bar),
    .I0(in_60bar),
    .I1(in_18bar)
  );
  //OR U438
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U438 (
    .O(n407),
    .I0(in[113]),
    .I1(n210)
  );
  //AND U438bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U438bar (
    .O(n407bar),
    .I0(inbar[113]),
    .I1(n210bar)
  );
  //OR U439
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U439 (
    .O(n210),
    .I0(n437),
    .I1(n438)
  );
  //AND U439bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U439bar (
    .O(n210bar),
    .I0(n437bar),
    .I1(n438bar)
  );
  //OR U440
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U440 (
    .O(n438),
    .I0(n439),
    .I1(n440)
  );
  //AND U440bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U440bar (
    .O(n438bar),
    .I0(n439bar),
    .I1(n440bar)
  );
  //OR U441
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U441 (
    .O(n440),
    .I0(n441),
    .I1(n442)
  );
  //AND U441bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U441bar (
    .O(n440bar),
    .I0(n441bar),
    .I1(n442bar)
  );
  //OR U442
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U442 (
    .O(n442),
    .I0(in[115]),
    .I1(in[110])
  );
  //AND U442bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U442bar (
    .O(n442bar),
    .I0(inbar[115]),
    .I1(inbar[110])
  );
  //OR U443
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U443 (
    .O(n441),
    .I0(in[125]),
    .I1(in[117])
  );
  //AND U443bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U443bar (
    .O(n441bar),
    .I0(inbar[125]),
    .I1(inbar[117])
  );
  //OR U444
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U444 (
    .O(n439),
    .I0(n443),
    .I1(n444)
  );
  //AND U444bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U444bar (
    .O(n439bar),
    .I0(n443bar),
    .I1(n444bar)
  );
  //OR U445
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U445 (
    .O(n444),
    .I0(in[180]),
    .I1(in[128])
  );
  //AND U445bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U445bar (
    .O(n444bar),
    .I0(inbar[180]),
    .I1(inbar[128])
  );
  //OR U446
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U446 (
    .O(n443),
    .I0(in[205]),
    .I1(in[201])
  );
  //AND U446bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U446bar (
    .O(n443bar),
    .I0(inbar[205]),
    .I1(inbar[201])
  );
  //OR U447
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U447 (
    .O(n437),
    .I0(n445),
    .I1(n446)
  );
  //AND U447bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U447bar (
    .O(n437bar),
    .I0(n445bar),
    .I1(n446bar)
  );
  //OR U448
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U448 (
    .O(n446),
    .I0(n447),
    .I1(n448)
  );
  //AND U448bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U448bar (
    .O(n446bar),
    .I0(n447bar),
    .I1(n448bar)
  );
  //OR U449
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U449 (
    .O(n448),
    .I0(in[244]),
    .I1(in[239])
  );
  //AND U449bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U449bar (
    .O(n448bar),
    .I0(inbar[244]),
    .I1(inbar[239])
  );
  //OR U450
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U450 (
    .O(n447),
    .I0(in[95]),
    .I1(in[83])
  );
  //AND U450bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U450bar (
    .O(n447bar),
    .I0(inbar[95]),
    .I1(inbar[83])
  );
  //OR U451
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U451 (
    .O(n445),
    .I0(n449),
    .I1(n450)
  );
  //AND U451bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U451bar (
    .O(n445bar),
    .I0(n449bar),
    .I1(n450bar)
  );
  //OR U452
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U452 (
    .O(n450),
    .I0(in_24),
    .I1(in[97])
  );
  //AND U452bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U452bar (
    .O(n450bar),
    .I0(in_24bar),
    .I1(inbar[97])
  );
  //OR U453
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U453 (
    .O(n449),
    .I0(in_33),
    .I1(in_27)
  );
  //AND U453bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U453bar (
    .O(n449bar),
    .I0(in_33bar),
    .I1(in_27bar)
  );
  //OR U454
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U454 (
    .O(n405),
    .I0(n451),
    .I1(n452)
  );
  //AND U454bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U454bar (
    .O(n405bar),
    .I0(n451bar),
    .I1(n452bar)
  );
  //OR U455
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U455 (
    .O(n452),
    .I0(in[145]),
    .I1(in[126])
  );
  //AND U455bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U455bar (
    .O(n452bar),
    .I0(inbar[145]),
    .I1(inbar[126])
  );
  //OR U456
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U456 (
    .O(n451),
    .I0(in[169]),
    .I1(n453)
  );
  //AND U456bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U456bar (
    .O(n451bar),
    .I0(inbar[169]),
    .I1(n453bar)
  );
  //OR U457
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U457 (
    .O(n453),
    .I0(in[221]),
    .I1(in[172])
  );
  //AND U457bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U457bar (
    .O(n453bar),
    .I0(inbar[221]),
    .I1(inbar[172])
  );
  //OR U458
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U458 (
    .O(n403),
    .I0(n454),
    .I1(n455)
  );
  //AND U458bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U458bar (
    .O(n403bar),
    .I0(n454bar),
    .I1(n455bar)
  );
  //OR U459
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U459 (
    .O(n455),
    .I0(n456),
    .I1(n457)
  );
  //AND U459bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U459bar (
    .O(n455bar),
    .I0(n456bar),
    .I1(n457bar)
  );
  //OR U460
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U460 (
    .O(n457),
    .I0(in[241]),
    .I1(in[224])
  );
  //AND U460bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U460bar (
    .O(n457bar),
    .I0(inbar[241]),
    .I1(inbar[224])
  );
  //OR U461
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U461 (
    .O(n456),
    .I0(in[86]),
    .I1(n458)
  );
  //AND U461bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U461bar (
    .O(n456bar),
    .I0(inbar[86]),
    .I1(n458bar)
  );
  //OR U462
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U462 (
    .O(n458),
    .I0(in_43),
    .I1(in_34)
  );
  //AND U462bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U462bar (
    .O(n458bar),
    .I0(in_43bar),
    .I1(in_34bar)
  );
  //OR U463
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U463 (
    .O(n454),
    .I0(n459),
    .I1(n460)
  );
  //AND U463bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U463bar (
    .O(n454bar),
    .I0(n459bar),
    .I1(n460bar)
  );
  //OR U464
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U464 (
    .O(n460),
    .I0(in_65),
    .I1(in_51)
  );
  //AND U464bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U464bar (
    .O(n460bar),
    .I0(in_65bar),
    .I1(in_51bar)
  );
  //OR U465
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U465 (
    .O(n459),
    .I0(in_75),
    .I1(n461)
  );
  //AND U465bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U465bar (
    .O(n459bar),
    .I0(in_75bar),
    .I1(n461bar)
  );
  //OR U466
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U466 (
    .O(n461),
    .I0(in_81),
    .I1(in_77)
  );
  //AND U466bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U466bar (
    .O(n461bar),
    .I0(in_81bar),
    .I1(in_77bar)
  );
  //OR U467
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U467 (
    .O(n195),
    .I0(n462),
    .I1(n463)
  );
  //AND U467bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U467bar (
    .O(n195bar),
    .I0(n462bar),
    .I1(n463bar)
  );
  //OR U468
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U468 (
    .O(n463),
    .I0(n464),
    .I1(n465)
  );
  //AND U468bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U468bar (
    .O(n463bar),
    .I0(n464bar),
    .I1(n465bar)
  );
  //OR U469
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U469 (
    .O(n465),
    .I0(n466),
    .I1(n467)
  );
  //AND U469bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U469bar (
    .O(n465bar),
    .I0(n466bar),
    .I1(n467bar)
  );
  //OR U470
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U470 (
    .O(n467),
    .I0(in[107]),
    .I1(in[101])
  );
  //AND U470bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U470bar (
    .O(n467bar),
    .I0(inbar[107]),
    .I1(inbar[101])
  );
  //OR U471
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U471 (
    .O(n466),
    .I0(in[139]),
    .I1(in[132])
  );
  //AND U471bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U471bar (
    .O(n466bar),
    .I0(inbar[139]),
    .I1(inbar[132])
  );
  //OR U472
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U472 (
    .O(n464),
    .I0(n468),
    .I1(n469)
  );
  //AND U472bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U472bar (
    .O(n464bar),
    .I0(n468bar),
    .I1(n469bar)
  );
  //OR U473
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U473 (
    .O(n469),
    .I0(in[146]),
    .I1(in[141])
  );
  //AND U473bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U473bar (
    .O(n469bar),
    .I0(inbar[146]),
    .I1(inbar[141])
  );
  //OR U474
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U474 (
    .O(n468),
    .I0(in[203]),
    .I1(in[179])
  );
  //AND U474bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U474bar (
    .O(n468bar),
    .I0(inbar[203]),
    .I1(inbar[179])
  );
  //OR U475
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U475 (
    .O(n462),
    .I0(n470),
    .I1(n471)
  );
  //AND U475bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U475bar (
    .O(n462bar),
    .I0(n470bar),
    .I1(n471bar)
  );
  //OR U476
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U476 (
    .O(n471),
    .I0(n472),
    .I1(n473)
  );
  //AND U476bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U476bar (
    .O(n471bar),
    .I0(n472bar),
    .I1(n473bar)
  );
  //OR U477
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U477 (
    .O(n473),
    .I0(in[243]),
    .I1(in[222])
  );
  //AND U477bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U477bar (
    .O(n473bar),
    .I0(inbar[243]),
    .I1(inbar[222])
  );
  //OR U478
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U478 (
    .O(n472),
    .I0(in[251]),
    .I1(in[250])
  );
  //AND U478bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U478bar (
    .O(n472bar),
    .I0(inbar[251]),
    .I1(inbar[250])
  );
  //OR U479
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U479 (
    .O(n470),
    .I0(n474),
    .I1(n475)
  );
  //AND U479bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U479bar (
    .O(n470bar),
    .I0(n474bar),
    .I1(n475bar)
  );
  //OR U480
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U480 (
    .O(n475),
    .I0(in_37),
    .I1(in_19)
  );
  //AND U480bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U480bar (
    .O(n475bar),
    .I0(in_37bar),
    .I1(in_19bar)
  );
  //OR U481
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U481 (
    .O(n474),
    .I0(in_78),
    .I1(in_6)
  );
  //AND U481bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U481bar (
    .O(n474bar),
    .I0(in_78bar),
    .I1(in_6bar)
  );
  //OR U482
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U482 (
    .O(n370),
    .I0(n476),
    .I1(n477)
  );
  //AND U482bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U482bar (
    .O(n370bar),
    .I0(n476bar),
    .I1(n477bar)
  );
  //OR U483
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U483 (
    .O(n477),
    .I0(in[112]),
    .I1(in[102])
  );
  //AND U483bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U483bar (
    .O(n477bar),
    .I0(inbar[112]),
    .I1(inbar[102])
  );
  //OR U484
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U484 (
    .O(n476),
    .I0(in[123]),
    .I1(n478)
  );
  //AND U484bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U484bar (
    .O(n476bar),
    .I0(inbar[123]),
    .I1(n478bar)
  );
  //OR U485
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U485 (
    .O(n478),
    .I0(in[143]),
    .I1(in[130])
  );
  //AND U485bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U485bar (
    .O(n478bar),
    .I0(inbar[143]),
    .I1(inbar[130])
  );
  //OR U486
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U486 (
    .O(n368),
    .I0(n479),
    .I1(n480)
  );
  //AND U486bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U486bar (
    .O(n368bar),
    .I0(n479bar),
    .I1(n480bar)
  );
  //OR U487
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U487 (
    .O(n480),
    .I0(n481),
    .I1(n482)
  );
  //AND U487bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U487bar (
    .O(n480bar),
    .I0(n481bar),
    .I1(n482bar)
  );
  //OR U488
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U488 (
    .O(n482),
    .I0(in[216]),
    .I1(in[213])
  );
  //AND U488bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U488bar (
    .O(n482bar),
    .I0(inbar[216]),
    .I1(inbar[213])
  );
  //OR U489
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U489 (
    .O(n481),
    .I0(in[227]),
    .I1(n483)
  );
  //AND U489bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U489bar (
    .O(n481bar),
    .I0(inbar[227]),
    .I1(n483bar)
  );
  //OR U490
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U490 (
    .O(n483),
    .I0(in_0),
    .I1(in[248])
  );
  //AND U490bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U490bar (
    .O(n483bar),
    .I0(in_0bar),
    .I1(inbar[248])
  );
  //OR U491
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U491 (
    .O(n479),
    .I0(n484),
    .I1(n485)
  );
  //AND U491bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U491bar (
    .O(n479bar),
    .I0(n484bar),
    .I1(n485bar)
  );
  //OR U492
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U492 (
    .O(n485),
    .I0(in_46),
    .I1(in_44)
  );
  //AND U492bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U492bar (
    .O(n485bar),
    .I0(in_46bar),
    .I1(in_44bar)
  );
  //OR U493
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U493 (
    .O(n484),
    .I0(in_50),
    .I1(n486)
  );
  //AND U493bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U493bar (
    .O(n484bar),
    .I0(in_50bar),
    .I1(n486bar)
  );
  //OR U494
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U494 (
    .O(n486),
    .I0(in_9),
    .I1(in_80)
  );
  //AND U494bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U494bar (
    .O(n486bar),
    .I0(in_9bar),
    .I1(in_80bar)
  );
endmodule

module sBox_0 ( in, out );

  input wire [7:0] in;
//input_done

  output wire [7:0] out;
//output_done

  wire [255:0] decodeOut;
//wire_done

  decode_0 dec ( .in(in), .out(decodeOut) );
  encode_0 enc ( .in(decodeOut), .out(out) );
endmodule

module CD2_1 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD2_2 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD2_3 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD2_4 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD4_1 ( a, b, y );

  input wire [3:0] a;
  input wire [3:0] b;
  wire [3:0] abar;
  wire [3:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
//input_done

  output wire [15:0] y;
  wire [15:0] ybar;
//output_done

//wire_done

  //AND U1
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1 (
    .O(y[9]),
    .I0(b[1]),
    .I1(a[2])
  );
  //OR U1bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1bar (
    .O(ybar[9]),
    .I0(bbar[1]),
    .I1(abar[2])
  );
  //AND U2
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2 (
    .O(y[8]),
    .I0(b[0]),
    .I1(a[2])
  );
  //OR U2bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2bar (
    .O(ybar[8]),
    .I0(bbar[0]),
    .I1(abar[2])
  );
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[7]),
    .I0(b[3]),
    .I1(a[1])
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[7]),
    .I0(bbar[3]),
    .I1(abar[1])
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[6]),
    .I0(b[2]),
    .I1(a[1])
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[6]),
    .I0(bbar[2]),
    .I1(abar[1])
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[5]),
    .I0(a[1]),
    .I1(b[1])
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[5]),
    .I0(abar[1]),
    .I1(bbar[1])
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[4]),
    .I0(a[1]),
    .I1(b[0])
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[4]),
    .I0(abar[1]),
    .I1(bbar[0])
  );
  //AND U7
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7 (
    .O(y[3]),
    .I0(a[0]),
    .I1(b[3])
  );
  //OR U7bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7bar (
    .O(ybar[3]),
    .I0(abar[0]),
    .I1(bbar[3])
  );
  //AND U8
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8 (
    .O(y[2]),
    .I0(a[0]),
    .I1(b[2])
  );
  //OR U8bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8bar (
    .O(ybar[2]),
    .I0(abar[0]),
    .I1(bbar[2])
  );
  //AND U9
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9 (
    .O(y[1]),
    .I0(a[0]),
    .I1(b[1])
  );
  //OR U9bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9bar (
    .O(ybar[1]),
    .I0(abar[0]),
    .I1(bbar[1])
  );
  //AND U10
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10 (
    .O(y[15]),
    .I0(a[3]),
    .I1(b[3])
  );
  //OR U10bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10bar (
    .O(ybar[15]),
    .I0(abar[3]),
    .I1(bbar[3])
  );
  //AND U11
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11 (
    .O(y[14]),
    .I0(a[3]),
    .I1(b[2])
  );
  //OR U11bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11bar (
    .O(ybar[14]),
    .I0(abar[3]),
    .I1(bbar[2])
  );
  //AND U12
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12 (
    .O(y[13]),
    .I0(a[3]),
    .I1(b[1])
  );
  //OR U12bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12bar (
    .O(ybar[13]),
    .I0(abar[3]),
    .I1(bbar[1])
  );
  //AND U13
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13 (
    .O(y[12]),
    .I0(a[3]),
    .I1(b[0])
  );
  //OR U13bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13bar (
    .O(ybar[12]),
    .I0(abar[3]),
    .I1(bbar[0])
  );
  //AND U14
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14 (
    .O(y[11]),
    .I0(b[3]),
    .I1(a[2])
  );
  //OR U14bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14bar (
    .O(ybar[11]),
    .I0(bbar[3]),
    .I1(abar[2])
  );
  //AND U15
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15 (
    .O(y[10]),
    .I0(b[2]),
    .I1(a[2])
  );
  //OR U15bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15bar (
    .O(ybar[10]),
    .I0(bbar[2]),
    .I1(abar[2])
  );
  //AND U16
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16 (
    .O(y[0]),
    .I0(a[0]),
    .I1(b[0])
  );
  //OR U16bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16bar (
    .O(ybar[0]),
    .I0(abar[0]),
    .I1(bbar[0])
  );
endmodule

module CD4_2 ( a, b, y );

  input wire [3:0] a;
  input wire [3:0] b;
  wire [3:0] abar;
  wire [3:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
//input_done

  output wire [15:0] y;
  wire [15:0] ybar;
//output_done

//wire_done

  //AND U1
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1 (
    .O(y[9]),
    .I0(b[1]),
    .I1(a[2])
  );
  //OR U1bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1bar (
    .O(ybar[9]),
    .I0(bbar[1]),
    .I1(abar[2])
  );
  //AND U2
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2 (
    .O(y[8]),
    .I0(b[0]),
    .I1(a[2])
  );
  //OR U2bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2bar (
    .O(ybar[8]),
    .I0(bbar[0]),
    .I1(abar[2])
  );
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[7]),
    .I0(b[3]),
    .I1(a[1])
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[7]),
    .I0(bbar[3]),
    .I1(abar[1])
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[6]),
    .I0(b[2]),
    .I1(a[1])
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[6]),
    .I0(bbar[2]),
    .I1(abar[1])
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[5]),
    .I0(a[1]),
    .I1(b[1])
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[5]),
    .I0(abar[1]),
    .I1(bbar[1])
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[4]),
    .I0(a[1]),
    .I1(b[0])
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[4]),
    .I0(abar[1]),
    .I1(bbar[0])
  );
  //AND U7
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7 (
    .O(y[3]),
    .I0(a[0]),
    .I1(b[3])
  );
  //OR U7bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7bar (
    .O(ybar[3]),
    .I0(abar[0]),
    .I1(bbar[3])
  );
  //AND U8
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8 (
    .O(y[2]),
    .I0(a[0]),
    .I1(b[2])
  );
  //OR U8bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8bar (
    .O(ybar[2]),
    .I0(abar[0]),
    .I1(bbar[2])
  );
  //AND U9
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9 (
    .O(y[1]),
    .I0(a[0]),
    .I1(b[1])
  );
  //OR U9bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9bar (
    .O(ybar[1]),
    .I0(abar[0]),
    .I1(bbar[1])
  );
  //AND U10
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10 (
    .O(y[15]),
    .I0(a[3]),
    .I1(b[3])
  );
  //OR U10bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10bar (
    .O(ybar[15]),
    .I0(abar[3]),
    .I1(bbar[3])
  );
  //AND U11
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11 (
    .O(y[14]),
    .I0(a[3]),
    .I1(b[2])
  );
  //OR U11bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11bar (
    .O(ybar[14]),
    .I0(abar[3]),
    .I1(bbar[2])
  );
  //AND U12
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12 (
    .O(y[13]),
    .I0(a[3]),
    .I1(b[1])
  );
  //OR U12bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12bar (
    .O(ybar[13]),
    .I0(abar[3]),
    .I1(bbar[1])
  );
  //AND U13
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13 (
    .O(y[12]),
    .I0(a[3]),
    .I1(b[0])
  );
  //OR U13bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13bar (
    .O(ybar[12]),
    .I0(abar[3]),
    .I1(bbar[0])
  );
  //AND U14
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14 (
    .O(y[11]),
    .I0(b[3]),
    .I1(a[2])
  );
  //OR U14bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14bar (
    .O(ybar[11]),
    .I0(bbar[3]),
    .I1(abar[2])
  );
  //AND U15
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15 (
    .O(y[10]),
    .I0(b[2]),
    .I1(a[2])
  );
  //OR U15bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15bar (
    .O(ybar[10]),
    .I0(bbar[2]),
    .I1(abar[2])
  );
  //AND U16
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16 (
    .O(y[0]),
    .I0(a[0]),
    .I1(b[0])
  );
  //OR U16bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16bar (
    .O(ybar[0]),
    .I0(abar[0]),
    .I1(bbar[0])
  );
endmodule

module CD16_1 ( a, b, y );

  input wire [15:0] a;
  input wire [15:0] b;
  wire [15:0] abar;
  wire [15:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign abar[8] = ~a[8];
  assign abar[9] = ~a[9];
  assign abar[10] = ~a[10];
  assign abar[11] = ~a[11];
  assign abar[12] = ~a[12];
  assign abar[13] = ~a[13];
  assign abar[14] = ~a[14];
  assign abar[15] = ~a[15];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign bbar[8] = ~b[8];
  assign bbar[9] = ~b[9];
  assign bbar[10] = ~b[10];
  assign bbar[11] = ~b[11];
  assign bbar[12] = ~b[12];
  assign bbar[13] = ~b[13];
  assign bbar[14] = ~b[14];
  assign bbar[15] = ~b[15];
//input_done

  output wire [255:0] y;
  wire [255:0] ybar;
//output_done

//wire_done

  //AND U1
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1 (
    .O(y[9]),
    .I0(b[9]),
    .I1(a[0])
  );
  //OR U1bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1bar (
    .O(ybar[9]),
    .I0(bbar[9]),
    .I1(abar[0])
  );
  //AND U2
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2 (
    .O(y[99]),
    .I0(b[3]),
    .I1(a[6])
  );
  //OR U2bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2bar (
    .O(ybar[99]),
    .I0(bbar[3]),
    .I1(abar[6])
  );
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[98]),
    .I0(b[2]),
    .I1(a[6])
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[98]),
    .I0(bbar[2]),
    .I1(abar[6])
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[97]),
    .I0(b[1]),
    .I1(a[6])
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[97]),
    .I0(bbar[1]),
    .I1(abar[6])
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[96]),
    .I0(b[0]),
    .I1(a[6])
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[96]),
    .I0(bbar[0]),
    .I1(abar[6])
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[95]),
    .I0(b[15]),
    .I1(a[5])
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[95]),
    .I0(bbar[15]),
    .I1(abar[5])
  );
  //AND U7
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7 (
    .O(y[94]),
    .I0(b[14]),
    .I1(a[5])
  );
  //OR U7bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7bar (
    .O(ybar[94]),
    .I0(bbar[14]),
    .I1(abar[5])
  );
  //AND U8
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8 (
    .O(y[93]),
    .I0(b[13]),
    .I1(a[5])
  );
  //OR U8bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8bar (
    .O(ybar[93]),
    .I0(bbar[13]),
    .I1(abar[5])
  );
  //AND U9
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9 (
    .O(y[92]),
    .I0(b[12]),
    .I1(a[5])
  );
  //OR U9bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9bar (
    .O(ybar[92]),
    .I0(bbar[12]),
    .I1(abar[5])
  );
  //AND U10
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10 (
    .O(y[91]),
    .I0(b[11]),
    .I1(a[5])
  );
  //OR U10bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10bar (
    .O(ybar[91]),
    .I0(bbar[11]),
    .I1(abar[5])
  );
  //AND U11
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11 (
    .O(y[90]),
    .I0(b[10]),
    .I1(a[5])
  );
  //OR U11bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11bar (
    .O(ybar[90]),
    .I0(bbar[10]),
    .I1(abar[5])
  );
  //AND U12
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12 (
    .O(y[8]),
    .I0(b[8]),
    .I1(a[0])
  );
  //OR U12bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12bar (
    .O(ybar[8]),
    .I0(bbar[8]),
    .I1(abar[0])
  );
  //AND U13
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13 (
    .O(y[89]),
    .I0(a[5]),
    .I1(b[9])
  );
  //OR U13bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13bar (
    .O(ybar[89]),
    .I0(abar[5]),
    .I1(bbar[9])
  );
  //AND U14
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14 (
    .O(y[88]),
    .I0(b[8]),
    .I1(a[5])
  );
  //OR U14bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14bar (
    .O(ybar[88]),
    .I0(bbar[8]),
    .I1(abar[5])
  );
  //AND U15
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15 (
    .O(y[87]),
    .I0(b[7]),
    .I1(a[5])
  );
  //OR U15bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15bar (
    .O(ybar[87]),
    .I0(bbar[7]),
    .I1(abar[5])
  );
  //AND U16
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16 (
    .O(y[86]),
    .I0(b[6]),
    .I1(a[5])
  );
  //OR U16bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16bar (
    .O(ybar[86]),
    .I0(bbar[6]),
    .I1(abar[5])
  );
  //AND U17
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U17 (
    .O(y[85]),
    .I0(b[5]),
    .I1(a[5])
  );
  //OR U17bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U17bar (
    .O(ybar[85]),
    .I0(bbar[5]),
    .I1(abar[5])
  );
  //AND U18
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U18 (
    .O(y[84]),
    .I0(b[4]),
    .I1(a[5])
  );
  //OR U18bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U18bar (
    .O(ybar[84]),
    .I0(bbar[4]),
    .I1(abar[5])
  );
  //AND U19
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U19 (
    .O(y[83]),
    .I0(a[5]),
    .I1(b[3])
  );
  //OR U19bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U19bar (
    .O(ybar[83]),
    .I0(abar[5]),
    .I1(bbar[3])
  );
  //AND U20
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U20 (
    .O(y[82]),
    .I0(a[5]),
    .I1(b[2])
  );
  //OR U20bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U20bar (
    .O(ybar[82]),
    .I0(abar[5]),
    .I1(bbar[2])
  );
  //AND U21
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U21 (
    .O(y[81]),
    .I0(a[5]),
    .I1(b[1])
  );
  //OR U21bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U21bar (
    .O(ybar[81]),
    .I0(abar[5]),
    .I1(bbar[1])
  );
  //AND U22
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U22 (
    .O(y[80]),
    .I0(a[5]),
    .I1(b[0])
  );
  //OR U22bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U22bar (
    .O(ybar[80]),
    .I0(abar[5]),
    .I1(bbar[0])
  );
  //AND U23
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U23 (
    .O(y[7]),
    .I0(b[7]),
    .I1(a[0])
  );
  //OR U23bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U23bar (
    .O(ybar[7]),
    .I0(bbar[7]),
    .I1(abar[0])
  );
  //AND U24
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U24 (
    .O(y[79]),
    .I0(a[4]),
    .I1(b[15])
  );
  //OR U24bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U24bar (
    .O(ybar[79]),
    .I0(abar[4]),
    .I1(bbar[15])
  );
  //AND U25
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U25 (
    .O(y[78]),
    .I0(a[4]),
    .I1(b[14])
  );
  //OR U25bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U25bar (
    .O(ybar[78]),
    .I0(abar[4]),
    .I1(bbar[14])
  );
  //AND U26
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U26 (
    .O(y[77]),
    .I0(a[4]),
    .I1(b[13])
  );
  //OR U26bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U26bar (
    .O(ybar[77]),
    .I0(abar[4]),
    .I1(bbar[13])
  );
  //AND U27
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U27 (
    .O(y[76]),
    .I0(a[4]),
    .I1(b[12])
  );
  //OR U27bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U27bar (
    .O(ybar[76]),
    .I0(abar[4]),
    .I1(bbar[12])
  );
  //AND U28
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U28 (
    .O(y[75]),
    .I0(a[4]),
    .I1(b[11])
  );
  //OR U28bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U28bar (
    .O(ybar[75]),
    .I0(abar[4]),
    .I1(bbar[11])
  );
  //AND U29
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U29 (
    .O(y[74]),
    .I0(a[4]),
    .I1(b[10])
  );
  //OR U29bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U29bar (
    .O(ybar[74]),
    .I0(abar[4]),
    .I1(bbar[10])
  );
  //AND U30
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U30 (
    .O(y[73]),
    .I0(a[4]),
    .I1(b[9])
  );
  //OR U30bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U30bar (
    .O(ybar[73]),
    .I0(abar[4]),
    .I1(bbar[9])
  );
  //AND U31
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U31 (
    .O(y[72]),
    .I0(a[4]),
    .I1(b[8])
  );
  //OR U31bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U31bar (
    .O(ybar[72]),
    .I0(abar[4]),
    .I1(bbar[8])
  );
  //AND U32
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U32 (
    .O(y[71]),
    .I0(a[4]),
    .I1(b[7])
  );
  //OR U32bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U32bar (
    .O(ybar[71]),
    .I0(abar[4]),
    .I1(bbar[7])
  );
  //AND U33
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U33 (
    .O(y[70]),
    .I0(a[4]),
    .I1(b[6])
  );
  //OR U33bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U33bar (
    .O(ybar[70]),
    .I0(abar[4]),
    .I1(bbar[6])
  );
  //AND U34
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U34 (
    .O(y[6]),
    .I0(b[6]),
    .I1(a[0])
  );
  //OR U34bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U34bar (
    .O(ybar[6]),
    .I0(bbar[6]),
    .I1(abar[0])
  );
  //AND U35
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U35 (
    .O(y[69]),
    .I0(a[4]),
    .I1(b[5])
  );
  //OR U35bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U35bar (
    .O(ybar[69]),
    .I0(abar[4]),
    .I1(bbar[5])
  );
  //AND U36
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U36 (
    .O(y[68]),
    .I0(a[4]),
    .I1(b[4])
  );
  //OR U36bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U36bar (
    .O(ybar[68]),
    .I0(abar[4]),
    .I1(bbar[4])
  );
  //AND U37
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U37 (
    .O(y[67]),
    .I0(a[4]),
    .I1(b[3])
  );
  //OR U37bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U37bar (
    .O(ybar[67]),
    .I0(abar[4]),
    .I1(bbar[3])
  );
  //AND U38
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U38 (
    .O(y[66]),
    .I0(a[4]),
    .I1(b[2])
  );
  //OR U38bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U38bar (
    .O(ybar[66]),
    .I0(abar[4]),
    .I1(bbar[2])
  );
  //AND U39
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U39 (
    .O(y[65]),
    .I0(a[4]),
    .I1(b[1])
  );
  //OR U39bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U39bar (
    .O(ybar[65]),
    .I0(abar[4]),
    .I1(bbar[1])
  );
  //AND U40
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U40 (
    .O(y[64]),
    .I0(a[4]),
    .I1(b[0])
  );
  //OR U40bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U40bar (
    .O(ybar[64]),
    .I0(abar[4]),
    .I1(bbar[0])
  );
  //AND U41
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U41 (
    .O(y[63]),
    .I0(a[3]),
    .I1(b[15])
  );
  //OR U41bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U41bar (
    .O(ybar[63]),
    .I0(abar[3]),
    .I1(bbar[15])
  );
  //AND U42
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U42 (
    .O(y[62]),
    .I0(a[3]),
    .I1(b[14])
  );
  //OR U42bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U42bar (
    .O(ybar[62]),
    .I0(abar[3]),
    .I1(bbar[14])
  );
  //AND U43
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U43 (
    .O(y[61]),
    .I0(a[3]),
    .I1(b[13])
  );
  //OR U43bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U43bar (
    .O(ybar[61]),
    .I0(abar[3]),
    .I1(bbar[13])
  );
  //AND U44
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U44 (
    .O(y[60]),
    .I0(a[3]),
    .I1(b[12])
  );
  //OR U44bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U44bar (
    .O(ybar[60]),
    .I0(abar[3]),
    .I1(bbar[12])
  );
  //AND U45
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U45 (
    .O(y[5]),
    .I0(b[5]),
    .I1(a[0])
  );
  //OR U45bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U45bar (
    .O(ybar[5]),
    .I0(bbar[5]),
    .I1(abar[0])
  );
  //AND U46
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U46 (
    .O(y[59]),
    .I0(a[3]),
    .I1(b[11])
  );
  //OR U46bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U46bar (
    .O(ybar[59]),
    .I0(abar[3]),
    .I1(bbar[11])
  );
  //AND U47
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U47 (
    .O(y[58]),
    .I0(a[3]),
    .I1(b[10])
  );
  //OR U47bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U47bar (
    .O(ybar[58]),
    .I0(abar[3]),
    .I1(bbar[10])
  );
  //AND U48
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U48 (
    .O(y[57]),
    .I0(a[3]),
    .I1(b[9])
  );
  //OR U48bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U48bar (
    .O(ybar[57]),
    .I0(abar[3]),
    .I1(bbar[9])
  );
  //AND U49
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U49 (
    .O(y[56]),
    .I0(a[3]),
    .I1(b[8])
  );
  //OR U49bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U49bar (
    .O(ybar[56]),
    .I0(abar[3]),
    .I1(bbar[8])
  );
  //AND U50
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U50 (
    .O(y[55]),
    .I0(a[3]),
    .I1(b[7])
  );
  //OR U50bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U50bar (
    .O(ybar[55]),
    .I0(abar[3]),
    .I1(bbar[7])
  );
  //AND U51
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U51 (
    .O(y[54]),
    .I0(a[3]),
    .I1(b[6])
  );
  //OR U51bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U51bar (
    .O(ybar[54]),
    .I0(abar[3]),
    .I1(bbar[6])
  );
  //AND U52
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U52 (
    .O(y[53]),
    .I0(a[3]),
    .I1(b[5])
  );
  //OR U52bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U52bar (
    .O(ybar[53]),
    .I0(abar[3]),
    .I1(bbar[5])
  );
  //AND U53
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U53 (
    .O(y[52]),
    .I0(a[3]),
    .I1(b[4])
  );
  //OR U53bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U53bar (
    .O(ybar[52]),
    .I0(abar[3]),
    .I1(bbar[4])
  );
  //AND U54
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U54 (
    .O(y[51]),
    .I0(a[3]),
    .I1(b[3])
  );
  //OR U54bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U54bar (
    .O(ybar[51]),
    .I0(abar[3]),
    .I1(bbar[3])
  );
  //AND U55
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U55 (
    .O(y[50]),
    .I0(a[3]),
    .I1(b[2])
  );
  //OR U55bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U55bar (
    .O(ybar[50]),
    .I0(abar[3]),
    .I1(bbar[2])
  );
  //AND U56
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U56 (
    .O(y[4]),
    .I0(b[4]),
    .I1(a[0])
  );
  //OR U56bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U56bar (
    .O(ybar[4]),
    .I0(bbar[4]),
    .I1(abar[0])
  );
  //AND U57
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U57 (
    .O(y[49]),
    .I0(a[3]),
    .I1(b[1])
  );
  //OR U57bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U57bar (
    .O(ybar[49]),
    .I0(abar[3]),
    .I1(bbar[1])
  );
  //AND U58
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U58 (
    .O(y[48]),
    .I0(a[3]),
    .I1(b[0])
  );
  //OR U58bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U58bar (
    .O(ybar[48]),
    .I0(abar[3]),
    .I1(bbar[0])
  );
  //AND U59
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U59 (
    .O(y[47]),
    .I0(a[2]),
    .I1(b[15])
  );
  //OR U59bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U59bar (
    .O(ybar[47]),
    .I0(abar[2]),
    .I1(bbar[15])
  );
  //AND U60
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U60 (
    .O(y[46]),
    .I0(a[2]),
    .I1(b[14])
  );
  //OR U60bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U60bar (
    .O(ybar[46]),
    .I0(abar[2]),
    .I1(bbar[14])
  );
  //AND U61
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U61 (
    .O(y[45]),
    .I0(a[2]),
    .I1(b[13])
  );
  //OR U61bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U61bar (
    .O(ybar[45]),
    .I0(abar[2]),
    .I1(bbar[13])
  );
  //AND U62
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U62 (
    .O(y[44]),
    .I0(a[2]),
    .I1(b[12])
  );
  //OR U62bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U62bar (
    .O(ybar[44]),
    .I0(abar[2]),
    .I1(bbar[12])
  );
  //AND U63
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U63 (
    .O(y[43]),
    .I0(a[2]),
    .I1(b[11])
  );
  //OR U63bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U63bar (
    .O(ybar[43]),
    .I0(abar[2]),
    .I1(bbar[11])
  );
  //AND U64
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U64 (
    .O(y[42]),
    .I0(a[2]),
    .I1(b[10])
  );
  //OR U64bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U64bar (
    .O(ybar[42]),
    .I0(abar[2]),
    .I1(bbar[10])
  );
  //AND U65
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U65 (
    .O(y[41]),
    .I0(a[2]),
    .I1(b[9])
  );
  //OR U65bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U65bar (
    .O(ybar[41]),
    .I0(abar[2]),
    .I1(bbar[9])
  );
  //AND U66
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U66 (
    .O(y[40]),
    .I0(a[2]),
    .I1(b[8])
  );
  //OR U66bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U66bar (
    .O(ybar[40]),
    .I0(abar[2]),
    .I1(bbar[8])
  );
  //AND U67
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U67 (
    .O(y[3]),
    .I0(b[3]),
    .I1(a[0])
  );
  //OR U67bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U67bar (
    .O(ybar[3]),
    .I0(bbar[3]),
    .I1(abar[0])
  );
  //AND U68
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U68 (
    .O(y[39]),
    .I0(a[2]),
    .I1(b[7])
  );
  //OR U68bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U68bar (
    .O(ybar[39]),
    .I0(abar[2]),
    .I1(bbar[7])
  );
  //AND U69
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U69 (
    .O(y[38]),
    .I0(a[2]),
    .I1(b[6])
  );
  //OR U69bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U69bar (
    .O(ybar[38]),
    .I0(abar[2]),
    .I1(bbar[6])
  );
  //AND U70
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U70 (
    .O(y[37]),
    .I0(a[2]),
    .I1(b[5])
  );
  //OR U70bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U70bar (
    .O(ybar[37]),
    .I0(abar[2]),
    .I1(bbar[5])
  );
  //AND U71
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U71 (
    .O(y[36]),
    .I0(a[2]),
    .I1(b[4])
  );
  //OR U71bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U71bar (
    .O(ybar[36]),
    .I0(abar[2]),
    .I1(bbar[4])
  );
  //AND U72
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U72 (
    .O(y[35]),
    .I0(a[2]),
    .I1(b[3])
  );
  //OR U72bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U72bar (
    .O(ybar[35]),
    .I0(abar[2]),
    .I1(bbar[3])
  );
  //AND U73
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U73 (
    .O(y[34]),
    .I0(a[2]),
    .I1(b[2])
  );
  //OR U73bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U73bar (
    .O(ybar[34]),
    .I0(abar[2]),
    .I1(bbar[2])
  );
  //AND U74
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U74 (
    .O(y[33]),
    .I0(a[2]),
    .I1(b[1])
  );
  //OR U74bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U74bar (
    .O(ybar[33]),
    .I0(abar[2]),
    .I1(bbar[1])
  );
  //AND U75
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U75 (
    .O(y[32]),
    .I0(a[2]),
    .I1(b[0])
  );
  //OR U75bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U75bar (
    .O(ybar[32]),
    .I0(abar[2]),
    .I1(bbar[0])
  );
  //AND U76
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U76 (
    .O(y[31]),
    .I0(a[1]),
    .I1(b[15])
  );
  //OR U76bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U76bar (
    .O(ybar[31]),
    .I0(abar[1]),
    .I1(bbar[15])
  );
  //AND U77
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U77 (
    .O(y[30]),
    .I0(a[1]),
    .I1(b[14])
  );
  //OR U77bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U77bar (
    .O(ybar[30]),
    .I0(abar[1]),
    .I1(bbar[14])
  );
  //AND U78
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U78 (
    .O(y[2]),
    .I0(b[2]),
    .I1(a[0])
  );
  //OR U78bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U78bar (
    .O(ybar[2]),
    .I0(bbar[2]),
    .I1(abar[0])
  );
  //AND U79
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U79 (
    .O(y[29]),
    .I0(a[1]),
    .I1(b[13])
  );
  //OR U79bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U79bar (
    .O(ybar[29]),
    .I0(abar[1]),
    .I1(bbar[13])
  );
  //AND U80
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U80 (
    .O(y[28]),
    .I0(a[1]),
    .I1(b[12])
  );
  //OR U80bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U80bar (
    .O(ybar[28]),
    .I0(abar[1]),
    .I1(bbar[12])
  );
  //AND U81
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U81 (
    .O(y[27]),
    .I0(a[1]),
    .I1(b[11])
  );
  //OR U81bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U81bar (
    .O(ybar[27]),
    .I0(abar[1]),
    .I1(bbar[11])
  );
  //AND U82
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U82 (
    .O(y[26]),
    .I0(a[1]),
    .I1(b[10])
  );
  //OR U82bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U82bar (
    .O(ybar[26]),
    .I0(abar[1]),
    .I1(bbar[10])
  );
  //AND U83
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U83 (
    .O(y[25]),
    .I0(a[1]),
    .I1(b[9])
  );
  //OR U83bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U83bar (
    .O(ybar[25]),
    .I0(abar[1]),
    .I1(bbar[9])
  );
  //AND U84
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U84 (
    .O(y[255]),
    .I0(a[15]),
    .I1(b[15])
  );
  //OR U84bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U84bar (
    .O(ybar[255]),
    .I0(abar[15]),
    .I1(bbar[15])
  );
  //AND U85
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U85 (
    .O(y[254]),
    .I0(a[15]),
    .I1(b[14])
  );
  //OR U85bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U85bar (
    .O(ybar[254]),
    .I0(abar[15]),
    .I1(bbar[14])
  );
  //AND U86
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U86 (
    .O(y[253]),
    .I0(a[15]),
    .I1(b[13])
  );
  //OR U86bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U86bar (
    .O(ybar[253]),
    .I0(abar[15]),
    .I1(bbar[13])
  );
  //AND U87
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U87 (
    .O(y[252]),
    .I0(a[15]),
    .I1(b[12])
  );
  //OR U87bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U87bar (
    .O(ybar[252]),
    .I0(abar[15]),
    .I1(bbar[12])
  );
  //AND U88
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U88 (
    .O(y[251]),
    .I0(a[15]),
    .I1(b[11])
  );
  //OR U88bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U88bar (
    .O(ybar[251]),
    .I0(abar[15]),
    .I1(bbar[11])
  );
  //AND U89
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U89 (
    .O(y[250]),
    .I0(a[15]),
    .I1(b[10])
  );
  //OR U89bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U89bar (
    .O(ybar[250]),
    .I0(abar[15]),
    .I1(bbar[10])
  );
  //AND U90
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U90 (
    .O(y[24]),
    .I0(a[1]),
    .I1(b[8])
  );
  //OR U90bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U90bar (
    .O(ybar[24]),
    .I0(abar[1]),
    .I1(bbar[8])
  );
  //AND U91
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U91 (
    .O(y[249]),
    .I0(a[15]),
    .I1(b[9])
  );
  //OR U91bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U91bar (
    .O(ybar[249]),
    .I0(abar[15]),
    .I1(bbar[9])
  );
  //AND U92
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U92 (
    .O(y[248]),
    .I0(a[15]),
    .I1(b[8])
  );
  //OR U92bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U92bar (
    .O(ybar[248]),
    .I0(abar[15]),
    .I1(bbar[8])
  );
  //AND U93
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U93 (
    .O(y[247]),
    .I0(a[15]),
    .I1(b[7])
  );
  //OR U93bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U93bar (
    .O(ybar[247]),
    .I0(abar[15]),
    .I1(bbar[7])
  );
  //AND U94
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U94 (
    .O(y[246]),
    .I0(a[15]),
    .I1(b[6])
  );
  //OR U94bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U94bar (
    .O(ybar[246]),
    .I0(abar[15]),
    .I1(bbar[6])
  );
  //AND U95
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U95 (
    .O(y[245]),
    .I0(a[15]),
    .I1(b[5])
  );
  //OR U95bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U95bar (
    .O(ybar[245]),
    .I0(abar[15]),
    .I1(bbar[5])
  );
  //AND U96
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U96 (
    .O(y[244]),
    .I0(a[15]),
    .I1(b[4])
  );
  //OR U96bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U96bar (
    .O(ybar[244]),
    .I0(abar[15]),
    .I1(bbar[4])
  );
  //AND U97
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U97 (
    .O(y[243]),
    .I0(a[15]),
    .I1(b[3])
  );
  //OR U97bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U97bar (
    .O(ybar[243]),
    .I0(abar[15]),
    .I1(bbar[3])
  );
  //AND U98
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U98 (
    .O(y[242]),
    .I0(a[15]),
    .I1(b[2])
  );
  //OR U98bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U98bar (
    .O(ybar[242]),
    .I0(abar[15]),
    .I1(bbar[2])
  );
  //AND U99
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U99 (
    .O(y[241]),
    .I0(a[15]),
    .I1(b[1])
  );
  //OR U99bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U99bar (
    .O(ybar[241]),
    .I0(abar[15]),
    .I1(bbar[1])
  );
  //AND U100
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U100 (
    .O(y[240]),
    .I0(a[15]),
    .I1(b[0])
  );
  //OR U100bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U100bar (
    .O(ybar[240]),
    .I0(abar[15]),
    .I1(bbar[0])
  );
  //AND U101
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U101 (
    .O(y[23]),
    .I0(a[1]),
    .I1(b[7])
  );
  //OR U101bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U101bar (
    .O(ybar[23]),
    .I0(abar[1]),
    .I1(bbar[7])
  );
  //AND U102
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U102 (
    .O(y[239]),
    .I0(a[14]),
    .I1(b[15])
  );
  //OR U102bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U102bar (
    .O(ybar[239]),
    .I0(abar[14]),
    .I1(bbar[15])
  );
  //AND U103
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U103 (
    .O(y[238]),
    .I0(a[14]),
    .I1(b[14])
  );
  //OR U103bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U103bar (
    .O(ybar[238]),
    .I0(abar[14]),
    .I1(bbar[14])
  );
  //AND U104
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U104 (
    .O(y[237]),
    .I0(a[14]),
    .I1(b[13])
  );
  //OR U104bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U104bar (
    .O(ybar[237]),
    .I0(abar[14]),
    .I1(bbar[13])
  );
  //AND U105
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U105 (
    .O(y[236]),
    .I0(a[14]),
    .I1(b[12])
  );
  //OR U105bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U105bar (
    .O(ybar[236]),
    .I0(abar[14]),
    .I1(bbar[12])
  );
  //AND U106
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U106 (
    .O(y[235]),
    .I0(a[14]),
    .I1(b[11])
  );
  //OR U106bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U106bar (
    .O(ybar[235]),
    .I0(abar[14]),
    .I1(bbar[11])
  );
  //AND U107
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U107 (
    .O(y[234]),
    .I0(a[14]),
    .I1(b[10])
  );
  //OR U107bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U107bar (
    .O(ybar[234]),
    .I0(abar[14]),
    .I1(bbar[10])
  );
  //AND U108
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U108 (
    .O(y[233]),
    .I0(a[14]),
    .I1(b[9])
  );
  //OR U108bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U108bar (
    .O(ybar[233]),
    .I0(abar[14]),
    .I1(bbar[9])
  );
  //AND U109
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U109 (
    .O(y[232]),
    .I0(a[14]),
    .I1(b[8])
  );
  //OR U109bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U109bar (
    .O(ybar[232]),
    .I0(abar[14]),
    .I1(bbar[8])
  );
  //AND U110
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U110 (
    .O(y[231]),
    .I0(a[14]),
    .I1(b[7])
  );
  //OR U110bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U110bar (
    .O(ybar[231]),
    .I0(abar[14]),
    .I1(bbar[7])
  );
  //AND U111
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U111 (
    .O(y[230]),
    .I0(a[14]),
    .I1(b[6])
  );
  //OR U111bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U111bar (
    .O(ybar[230]),
    .I0(abar[14]),
    .I1(bbar[6])
  );
  //AND U112
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U112 (
    .O(y[22]),
    .I0(a[1]),
    .I1(b[6])
  );
  //OR U112bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U112bar (
    .O(ybar[22]),
    .I0(abar[1]),
    .I1(bbar[6])
  );
  //AND U113
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U113 (
    .O(y[229]),
    .I0(a[14]),
    .I1(b[5])
  );
  //OR U113bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U113bar (
    .O(ybar[229]),
    .I0(abar[14]),
    .I1(bbar[5])
  );
  //AND U114
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U114 (
    .O(y[228]),
    .I0(a[14]),
    .I1(b[4])
  );
  //OR U114bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U114bar (
    .O(ybar[228]),
    .I0(abar[14]),
    .I1(bbar[4])
  );
  //AND U115
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U115 (
    .O(y[227]),
    .I0(a[14]),
    .I1(b[3])
  );
  //OR U115bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U115bar (
    .O(ybar[227]),
    .I0(abar[14]),
    .I1(bbar[3])
  );
  //AND U116
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U116 (
    .O(y[226]),
    .I0(a[14]),
    .I1(b[2])
  );
  //OR U116bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U116bar (
    .O(ybar[226]),
    .I0(abar[14]),
    .I1(bbar[2])
  );
  //AND U117
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U117 (
    .O(y[225]),
    .I0(a[14]),
    .I1(b[1])
  );
  //OR U117bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U117bar (
    .O(ybar[225]),
    .I0(abar[14]),
    .I1(bbar[1])
  );
  //AND U118
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U118 (
    .O(y[224]),
    .I0(a[14]),
    .I1(b[0])
  );
  //OR U118bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U118bar (
    .O(ybar[224]),
    .I0(abar[14]),
    .I1(bbar[0])
  );
  //AND U119
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U119 (
    .O(y[223]),
    .I0(a[13]),
    .I1(b[15])
  );
  //OR U119bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U119bar (
    .O(ybar[223]),
    .I0(abar[13]),
    .I1(bbar[15])
  );
  //AND U120
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U120 (
    .O(y[222]),
    .I0(a[13]),
    .I1(b[14])
  );
  //OR U120bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U120bar (
    .O(ybar[222]),
    .I0(abar[13]),
    .I1(bbar[14])
  );
  //AND U121
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U121 (
    .O(y[221]),
    .I0(a[13]),
    .I1(b[13])
  );
  //OR U121bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U121bar (
    .O(ybar[221]),
    .I0(abar[13]),
    .I1(bbar[13])
  );
  //AND U122
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U122 (
    .O(y[220]),
    .I0(a[13]),
    .I1(b[12])
  );
  //OR U122bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U122bar (
    .O(ybar[220]),
    .I0(abar[13]),
    .I1(bbar[12])
  );
  //AND U123
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U123 (
    .O(y[21]),
    .I0(a[1]),
    .I1(b[5])
  );
  //OR U123bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U123bar (
    .O(ybar[21]),
    .I0(abar[1]),
    .I1(bbar[5])
  );
  //AND U124
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U124 (
    .O(y[219]),
    .I0(a[13]),
    .I1(b[11])
  );
  //OR U124bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U124bar (
    .O(ybar[219]),
    .I0(abar[13]),
    .I1(bbar[11])
  );
  //AND U125
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U125 (
    .O(y[218]),
    .I0(a[13]),
    .I1(b[10])
  );
  //OR U125bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U125bar (
    .O(ybar[218]),
    .I0(abar[13]),
    .I1(bbar[10])
  );
  //AND U126
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U126 (
    .O(y[217]),
    .I0(a[13]),
    .I1(b[9])
  );
  //OR U126bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U126bar (
    .O(ybar[217]),
    .I0(abar[13]),
    .I1(bbar[9])
  );
  //AND U127
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U127 (
    .O(y[216]),
    .I0(a[13]),
    .I1(b[8])
  );
  //OR U127bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U127bar (
    .O(ybar[216]),
    .I0(abar[13]),
    .I1(bbar[8])
  );
  //AND U128
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U128 (
    .O(y[215]),
    .I0(a[13]),
    .I1(b[7])
  );
  //OR U128bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U128bar (
    .O(ybar[215]),
    .I0(abar[13]),
    .I1(bbar[7])
  );
  //AND U129
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U129 (
    .O(y[214]),
    .I0(a[13]),
    .I1(b[6])
  );
  //OR U129bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U129bar (
    .O(ybar[214]),
    .I0(abar[13]),
    .I1(bbar[6])
  );
  //AND U130
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U130 (
    .O(y[213]),
    .I0(a[13]),
    .I1(b[5])
  );
  //OR U130bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U130bar (
    .O(ybar[213]),
    .I0(abar[13]),
    .I1(bbar[5])
  );
  //AND U131
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U131 (
    .O(y[212]),
    .I0(a[13]),
    .I1(b[4])
  );
  //OR U131bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U131bar (
    .O(ybar[212]),
    .I0(abar[13]),
    .I1(bbar[4])
  );
  //AND U132
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U132 (
    .O(y[211]),
    .I0(a[13]),
    .I1(b[3])
  );
  //OR U132bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U132bar (
    .O(ybar[211]),
    .I0(abar[13]),
    .I1(bbar[3])
  );
  //AND U133
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U133 (
    .O(y[210]),
    .I0(a[13]),
    .I1(b[2])
  );
  //OR U133bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U133bar (
    .O(ybar[210]),
    .I0(abar[13]),
    .I1(bbar[2])
  );
  //AND U134
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U134 (
    .O(y[20]),
    .I0(a[1]),
    .I1(b[4])
  );
  //OR U134bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U134bar (
    .O(ybar[20]),
    .I0(abar[1]),
    .I1(bbar[4])
  );
  //AND U135
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U135 (
    .O(y[209]),
    .I0(a[13]),
    .I1(b[1])
  );
  //OR U135bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U135bar (
    .O(ybar[209]),
    .I0(abar[13]),
    .I1(bbar[1])
  );
  //AND U136
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U136 (
    .O(y[208]),
    .I0(a[13]),
    .I1(b[0])
  );
  //OR U136bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U136bar (
    .O(ybar[208]),
    .I0(abar[13]),
    .I1(bbar[0])
  );
  //AND U137
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U137 (
    .O(y[207]),
    .I0(a[12]),
    .I1(b[15])
  );
  //OR U137bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U137bar (
    .O(ybar[207]),
    .I0(abar[12]),
    .I1(bbar[15])
  );
  //AND U138
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U138 (
    .O(y[206]),
    .I0(a[12]),
    .I1(b[14])
  );
  //OR U138bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U138bar (
    .O(ybar[206]),
    .I0(abar[12]),
    .I1(bbar[14])
  );
  //AND U139
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U139 (
    .O(y[205]),
    .I0(a[12]),
    .I1(b[13])
  );
  //OR U139bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U139bar (
    .O(ybar[205]),
    .I0(abar[12]),
    .I1(bbar[13])
  );
  //AND U140
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U140 (
    .O(y[204]),
    .I0(a[12]),
    .I1(b[12])
  );
  //OR U140bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U140bar (
    .O(ybar[204]),
    .I0(abar[12]),
    .I1(bbar[12])
  );
  //AND U141
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U141 (
    .O(y[203]),
    .I0(a[12]),
    .I1(b[11])
  );
  //OR U141bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U141bar (
    .O(ybar[203]),
    .I0(abar[12]),
    .I1(bbar[11])
  );
  //AND U142
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U142 (
    .O(y[202]),
    .I0(a[12]),
    .I1(b[10])
  );
  //OR U142bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U142bar (
    .O(ybar[202]),
    .I0(abar[12]),
    .I1(bbar[10])
  );
  //AND U143
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U143 (
    .O(y[201]),
    .I0(a[12]),
    .I1(b[9])
  );
  //OR U143bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U143bar (
    .O(ybar[201]),
    .I0(abar[12]),
    .I1(bbar[9])
  );
  //AND U144
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U144 (
    .O(y[200]),
    .I0(a[12]),
    .I1(b[8])
  );
  //OR U144bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U144bar (
    .O(ybar[200]),
    .I0(abar[12]),
    .I1(bbar[8])
  );
  //AND U145
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U145 (
    .O(y[1]),
    .I0(b[1]),
    .I1(a[0])
  );
  //OR U145bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U145bar (
    .O(ybar[1]),
    .I0(bbar[1]),
    .I1(abar[0])
  );
  //AND U146
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U146 (
    .O(y[19]),
    .I0(a[1]),
    .I1(b[3])
  );
  //OR U146bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U146bar (
    .O(ybar[19]),
    .I0(abar[1]),
    .I1(bbar[3])
  );
  //AND U147
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U147 (
    .O(y[199]),
    .I0(a[12]),
    .I1(b[7])
  );
  //OR U147bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U147bar (
    .O(ybar[199]),
    .I0(abar[12]),
    .I1(bbar[7])
  );
  //AND U148
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U148 (
    .O(y[198]),
    .I0(a[12]),
    .I1(b[6])
  );
  //OR U148bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U148bar (
    .O(ybar[198]),
    .I0(abar[12]),
    .I1(bbar[6])
  );
  //AND U149
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U149 (
    .O(y[197]),
    .I0(a[12]),
    .I1(b[5])
  );
  //OR U149bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U149bar (
    .O(ybar[197]),
    .I0(abar[12]),
    .I1(bbar[5])
  );
  //AND U150
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U150 (
    .O(y[196]),
    .I0(a[12]),
    .I1(b[4])
  );
  //OR U150bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U150bar (
    .O(ybar[196]),
    .I0(abar[12]),
    .I1(bbar[4])
  );
  //AND U151
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U151 (
    .O(y[195]),
    .I0(a[12]),
    .I1(b[3])
  );
  //OR U151bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U151bar (
    .O(ybar[195]),
    .I0(abar[12]),
    .I1(bbar[3])
  );
  //AND U152
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U152 (
    .O(y[194]),
    .I0(a[12]),
    .I1(b[2])
  );
  //OR U152bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U152bar (
    .O(ybar[194]),
    .I0(abar[12]),
    .I1(bbar[2])
  );
  //AND U153
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U153 (
    .O(y[193]),
    .I0(a[12]),
    .I1(b[1])
  );
  //OR U153bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U153bar (
    .O(ybar[193]),
    .I0(abar[12]),
    .I1(bbar[1])
  );
  //AND U154
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U154 (
    .O(y[192]),
    .I0(a[12]),
    .I1(b[0])
  );
  //OR U154bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U154bar (
    .O(ybar[192]),
    .I0(abar[12]),
    .I1(bbar[0])
  );
  //AND U155
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U155 (
    .O(y[191]),
    .I0(a[11]),
    .I1(b[15])
  );
  //OR U155bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U155bar (
    .O(ybar[191]),
    .I0(abar[11]),
    .I1(bbar[15])
  );
  //AND U156
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U156 (
    .O(y[190]),
    .I0(a[11]),
    .I1(b[14])
  );
  //OR U156bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U156bar (
    .O(ybar[190]),
    .I0(abar[11]),
    .I1(bbar[14])
  );
  //AND U157
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U157 (
    .O(y[18]),
    .I0(a[1]),
    .I1(b[2])
  );
  //OR U157bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U157bar (
    .O(ybar[18]),
    .I0(abar[1]),
    .I1(bbar[2])
  );
  //AND U158
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U158 (
    .O(y[189]),
    .I0(a[11]),
    .I1(b[13])
  );
  //OR U158bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U158bar (
    .O(ybar[189]),
    .I0(abar[11]),
    .I1(bbar[13])
  );
  //AND U159
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U159 (
    .O(y[188]),
    .I0(a[11]),
    .I1(b[12])
  );
  //OR U159bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U159bar (
    .O(ybar[188]),
    .I0(abar[11]),
    .I1(bbar[12])
  );
  //AND U160
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U160 (
    .O(y[187]),
    .I0(a[11]),
    .I1(b[11])
  );
  //OR U160bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U160bar (
    .O(ybar[187]),
    .I0(abar[11]),
    .I1(bbar[11])
  );
  //AND U161
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U161 (
    .O(y[186]),
    .I0(a[11]),
    .I1(b[10])
  );
  //OR U161bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U161bar (
    .O(ybar[186]),
    .I0(abar[11]),
    .I1(bbar[10])
  );
  //AND U162
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U162 (
    .O(y[185]),
    .I0(a[11]),
    .I1(b[9])
  );
  //OR U162bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U162bar (
    .O(ybar[185]),
    .I0(abar[11]),
    .I1(bbar[9])
  );
  //AND U163
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U163 (
    .O(y[184]),
    .I0(a[11]),
    .I1(b[8])
  );
  //OR U163bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U163bar (
    .O(ybar[184]),
    .I0(abar[11]),
    .I1(bbar[8])
  );
  //AND U164
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U164 (
    .O(y[183]),
    .I0(a[11]),
    .I1(b[7])
  );
  //OR U164bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U164bar (
    .O(ybar[183]),
    .I0(abar[11]),
    .I1(bbar[7])
  );
  //AND U165
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U165 (
    .O(y[182]),
    .I0(a[11]),
    .I1(b[6])
  );
  //OR U165bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U165bar (
    .O(ybar[182]),
    .I0(abar[11]),
    .I1(bbar[6])
  );
  //AND U166
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U166 (
    .O(y[181]),
    .I0(a[11]),
    .I1(b[5])
  );
  //OR U166bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U166bar (
    .O(ybar[181]),
    .I0(abar[11]),
    .I1(bbar[5])
  );
  //AND U167
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U167 (
    .O(y[180]),
    .I0(a[11]),
    .I1(b[4])
  );
  //OR U167bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U167bar (
    .O(ybar[180]),
    .I0(abar[11]),
    .I1(bbar[4])
  );
  //AND U168
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U168 (
    .O(y[17]),
    .I0(a[1]),
    .I1(b[1])
  );
  //OR U168bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U168bar (
    .O(ybar[17]),
    .I0(abar[1]),
    .I1(bbar[1])
  );
  //AND U169
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U169 (
    .O(y[179]),
    .I0(a[11]),
    .I1(b[3])
  );
  //OR U169bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U169bar (
    .O(ybar[179]),
    .I0(abar[11]),
    .I1(bbar[3])
  );
  //AND U170
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U170 (
    .O(y[178]),
    .I0(a[11]),
    .I1(b[2])
  );
  //OR U170bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U170bar (
    .O(ybar[178]),
    .I0(abar[11]),
    .I1(bbar[2])
  );
  //AND U171
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U171 (
    .O(y[177]),
    .I0(a[11]),
    .I1(b[1])
  );
  //OR U171bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U171bar (
    .O(ybar[177]),
    .I0(abar[11]),
    .I1(bbar[1])
  );
  //AND U172
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U172 (
    .O(y[176]),
    .I0(a[11]),
    .I1(b[0])
  );
  //OR U172bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U172bar (
    .O(ybar[176]),
    .I0(abar[11]),
    .I1(bbar[0])
  );
  //AND U173
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U173 (
    .O(y[175]),
    .I0(a[10]),
    .I1(b[15])
  );
  //OR U173bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U173bar (
    .O(ybar[175]),
    .I0(abar[10]),
    .I1(bbar[15])
  );
  //AND U174
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U174 (
    .O(y[174]),
    .I0(a[10]),
    .I1(b[14])
  );
  //OR U174bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U174bar (
    .O(ybar[174]),
    .I0(abar[10]),
    .I1(bbar[14])
  );
  //AND U175
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U175 (
    .O(y[173]),
    .I0(a[10]),
    .I1(b[13])
  );
  //OR U175bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U175bar (
    .O(ybar[173]),
    .I0(abar[10]),
    .I1(bbar[13])
  );
  //AND U176
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U176 (
    .O(y[172]),
    .I0(a[10]),
    .I1(b[12])
  );
  //OR U176bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U176bar (
    .O(ybar[172]),
    .I0(abar[10]),
    .I1(bbar[12])
  );
  //AND U177
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U177 (
    .O(y[171]),
    .I0(a[10]),
    .I1(b[11])
  );
  //OR U177bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U177bar (
    .O(ybar[171]),
    .I0(abar[10]),
    .I1(bbar[11])
  );
  //AND U178
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U178 (
    .O(y[170]),
    .I0(a[10]),
    .I1(b[10])
  );
  //OR U178bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U178bar (
    .O(ybar[170]),
    .I0(abar[10]),
    .I1(bbar[10])
  );
  //AND U179
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U179 (
    .O(y[16]),
    .I0(a[1]),
    .I1(b[0])
  );
  //OR U179bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U179bar (
    .O(ybar[16]),
    .I0(abar[1]),
    .I1(bbar[0])
  );
  //AND U180
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U180 (
    .O(y[169]),
    .I0(a[10]),
    .I1(b[9])
  );
  //OR U180bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U180bar (
    .O(ybar[169]),
    .I0(abar[10]),
    .I1(bbar[9])
  );
  //AND U181
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U181 (
    .O(y[168]),
    .I0(a[10]),
    .I1(b[8])
  );
  //OR U181bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U181bar (
    .O(ybar[168]),
    .I0(abar[10]),
    .I1(bbar[8])
  );
  //AND U182
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U182 (
    .O(y[167]),
    .I0(a[10]),
    .I1(b[7])
  );
  //OR U182bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U182bar (
    .O(ybar[167]),
    .I0(abar[10]),
    .I1(bbar[7])
  );
  //AND U183
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U183 (
    .O(y[166]),
    .I0(a[10]),
    .I1(b[6])
  );
  //OR U183bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U183bar (
    .O(ybar[166]),
    .I0(abar[10]),
    .I1(bbar[6])
  );
  //AND U184
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U184 (
    .O(y[165]),
    .I0(a[10]),
    .I1(b[5])
  );
  //OR U184bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U184bar (
    .O(ybar[165]),
    .I0(abar[10]),
    .I1(bbar[5])
  );
  //AND U185
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U185 (
    .O(y[164]),
    .I0(a[10]),
    .I1(b[4])
  );
  //OR U185bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U185bar (
    .O(ybar[164]),
    .I0(abar[10]),
    .I1(bbar[4])
  );
  //AND U186
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U186 (
    .O(y[163]),
    .I0(a[10]),
    .I1(b[3])
  );
  //OR U186bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U186bar (
    .O(ybar[163]),
    .I0(abar[10]),
    .I1(bbar[3])
  );
  //AND U187
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U187 (
    .O(y[162]),
    .I0(a[10]),
    .I1(b[2])
  );
  //OR U187bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U187bar (
    .O(ybar[162]),
    .I0(abar[10]),
    .I1(bbar[2])
  );
  //AND U188
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U188 (
    .O(y[161]),
    .I0(a[10]),
    .I1(b[1])
  );
  //OR U188bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U188bar (
    .O(ybar[161]),
    .I0(abar[10]),
    .I1(bbar[1])
  );
  //AND U189
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U189 (
    .O(y[160]),
    .I0(a[10]),
    .I1(b[0])
  );
  //OR U189bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U189bar (
    .O(ybar[160]),
    .I0(abar[10]),
    .I1(bbar[0])
  );
  //AND U190
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U190 (
    .O(y[15]),
    .I0(b[15]),
    .I1(a[0])
  );
  //OR U190bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U190bar (
    .O(ybar[15]),
    .I0(bbar[15]),
    .I1(abar[0])
  );
  //AND U191
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U191 (
    .O(y[159]),
    .I0(a[9]),
    .I1(b[15])
  );
  //OR U191bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U191bar (
    .O(ybar[159]),
    .I0(abar[9]),
    .I1(bbar[15])
  );
  //AND U192
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U192 (
    .O(y[158]),
    .I0(a[9]),
    .I1(b[14])
  );
  //OR U192bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U192bar (
    .O(ybar[158]),
    .I0(abar[9]),
    .I1(bbar[14])
  );
  //AND U193
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U193 (
    .O(y[157]),
    .I0(a[9]),
    .I1(b[13])
  );
  //OR U193bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U193bar (
    .O(ybar[157]),
    .I0(abar[9]),
    .I1(bbar[13])
  );
  //AND U194
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U194 (
    .O(y[156]),
    .I0(a[9]),
    .I1(b[12])
  );
  //OR U194bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U194bar (
    .O(ybar[156]),
    .I0(abar[9]),
    .I1(bbar[12])
  );
  //AND U195
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U195 (
    .O(y[155]),
    .I0(a[9]),
    .I1(b[11])
  );
  //OR U195bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U195bar (
    .O(ybar[155]),
    .I0(abar[9]),
    .I1(bbar[11])
  );
  //AND U196
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U196 (
    .O(y[154]),
    .I0(a[9]),
    .I1(b[10])
  );
  //OR U196bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U196bar (
    .O(ybar[154]),
    .I0(abar[9]),
    .I1(bbar[10])
  );
  //AND U197
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U197 (
    .O(y[153]),
    .I0(a[9]),
    .I1(b[9])
  );
  //OR U197bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U197bar (
    .O(ybar[153]),
    .I0(abar[9]),
    .I1(bbar[9])
  );
  //AND U198
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U198 (
    .O(y[152]),
    .I0(a[9]),
    .I1(b[8])
  );
  //OR U198bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U198bar (
    .O(ybar[152]),
    .I0(abar[9]),
    .I1(bbar[8])
  );
  //AND U199
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U199 (
    .O(y[151]),
    .I0(a[9]),
    .I1(b[7])
  );
  //OR U199bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U199bar (
    .O(ybar[151]),
    .I0(abar[9]),
    .I1(bbar[7])
  );
  //AND U200
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U200 (
    .O(y[150]),
    .I0(a[9]),
    .I1(b[6])
  );
  //OR U200bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U200bar (
    .O(ybar[150]),
    .I0(abar[9]),
    .I1(bbar[6])
  );
  //AND U201
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U201 (
    .O(y[14]),
    .I0(b[14]),
    .I1(a[0])
  );
  //OR U201bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U201bar (
    .O(ybar[14]),
    .I0(bbar[14]),
    .I1(abar[0])
  );
  //AND U202
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U202 (
    .O(y[149]),
    .I0(a[9]),
    .I1(b[5])
  );
  //OR U202bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U202bar (
    .O(ybar[149]),
    .I0(abar[9]),
    .I1(bbar[5])
  );
  //AND U203
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U203 (
    .O(y[148]),
    .I0(a[9]),
    .I1(b[4])
  );
  //OR U203bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U203bar (
    .O(ybar[148]),
    .I0(abar[9]),
    .I1(bbar[4])
  );
  //AND U204
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U204 (
    .O(y[147]),
    .I0(a[9]),
    .I1(b[3])
  );
  //OR U204bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U204bar (
    .O(ybar[147]),
    .I0(abar[9]),
    .I1(bbar[3])
  );
  //AND U205
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U205 (
    .O(y[146]),
    .I0(a[9]),
    .I1(b[2])
  );
  //OR U205bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U205bar (
    .O(ybar[146]),
    .I0(abar[9]),
    .I1(bbar[2])
  );
  //AND U206
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U206 (
    .O(y[145]),
    .I0(a[9]),
    .I1(b[1])
  );
  //OR U206bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U206bar (
    .O(ybar[145]),
    .I0(abar[9]),
    .I1(bbar[1])
  );
  //AND U207
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U207 (
    .O(y[144]),
    .I0(a[9]),
    .I1(b[0])
  );
  //OR U207bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U207bar (
    .O(ybar[144]),
    .I0(abar[9]),
    .I1(bbar[0])
  );
  //AND U208
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U208 (
    .O(y[143]),
    .I0(a[8]),
    .I1(b[15])
  );
  //OR U208bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U208bar (
    .O(ybar[143]),
    .I0(abar[8]),
    .I1(bbar[15])
  );
  //AND U209
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U209 (
    .O(y[142]),
    .I0(a[8]),
    .I1(b[14])
  );
  //OR U209bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U209bar (
    .O(ybar[142]),
    .I0(abar[8]),
    .I1(bbar[14])
  );
  //AND U210
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U210 (
    .O(y[141]),
    .I0(a[8]),
    .I1(b[13])
  );
  //OR U210bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U210bar (
    .O(ybar[141]),
    .I0(abar[8]),
    .I1(bbar[13])
  );
  //AND U211
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U211 (
    .O(y[140]),
    .I0(a[8]),
    .I1(b[12])
  );
  //OR U211bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U211bar (
    .O(ybar[140]),
    .I0(abar[8]),
    .I1(bbar[12])
  );
  //AND U212
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U212 (
    .O(y[13]),
    .I0(b[13]),
    .I1(a[0])
  );
  //OR U212bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U212bar (
    .O(ybar[13]),
    .I0(bbar[13]),
    .I1(abar[0])
  );
  //AND U213
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U213 (
    .O(y[139]),
    .I0(a[8]),
    .I1(b[11])
  );
  //OR U213bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U213bar (
    .O(ybar[139]),
    .I0(abar[8]),
    .I1(bbar[11])
  );
  //AND U214
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U214 (
    .O(y[138]),
    .I0(a[8]),
    .I1(b[10])
  );
  //OR U214bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U214bar (
    .O(ybar[138]),
    .I0(abar[8]),
    .I1(bbar[10])
  );
  //AND U215
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U215 (
    .O(y[137]),
    .I0(a[8]),
    .I1(b[9])
  );
  //OR U215bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U215bar (
    .O(ybar[137]),
    .I0(abar[8]),
    .I1(bbar[9])
  );
  //AND U216
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U216 (
    .O(y[136]),
    .I0(a[8]),
    .I1(b[8])
  );
  //OR U216bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U216bar (
    .O(ybar[136]),
    .I0(abar[8]),
    .I1(bbar[8])
  );
  //AND U217
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U217 (
    .O(y[135]),
    .I0(a[8]),
    .I1(b[7])
  );
  //OR U217bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U217bar (
    .O(ybar[135]),
    .I0(abar[8]),
    .I1(bbar[7])
  );
  //AND U218
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U218 (
    .O(y[134]),
    .I0(a[8]),
    .I1(b[6])
  );
  //OR U218bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U218bar (
    .O(ybar[134]),
    .I0(abar[8]),
    .I1(bbar[6])
  );
  //AND U219
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U219 (
    .O(y[133]),
    .I0(a[8]),
    .I1(b[5])
  );
  //OR U219bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U219bar (
    .O(ybar[133]),
    .I0(abar[8]),
    .I1(bbar[5])
  );
  //AND U220
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U220 (
    .O(y[132]),
    .I0(a[8]),
    .I1(b[4])
  );
  //OR U220bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U220bar (
    .O(ybar[132]),
    .I0(abar[8]),
    .I1(bbar[4])
  );
  //AND U221
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U221 (
    .O(y[131]),
    .I0(a[8]),
    .I1(b[3])
  );
  //OR U221bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U221bar (
    .O(ybar[131]),
    .I0(abar[8]),
    .I1(bbar[3])
  );
  //AND U222
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U222 (
    .O(y[130]),
    .I0(a[8]),
    .I1(b[2])
  );
  //OR U222bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U222bar (
    .O(ybar[130]),
    .I0(abar[8]),
    .I1(bbar[2])
  );
  //AND U223
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U223 (
    .O(y[12]),
    .I0(b[12]),
    .I1(a[0])
  );
  //OR U223bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U223bar (
    .O(ybar[12]),
    .I0(bbar[12]),
    .I1(abar[0])
  );
  //AND U224
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U224 (
    .O(y[129]),
    .I0(a[8]),
    .I1(b[1])
  );
  //OR U224bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U224bar (
    .O(ybar[129]),
    .I0(abar[8]),
    .I1(bbar[1])
  );
  //AND U225
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U225 (
    .O(y[128]),
    .I0(a[8]),
    .I1(b[0])
  );
  //OR U225bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U225bar (
    .O(ybar[128]),
    .I0(abar[8]),
    .I1(bbar[0])
  );
  //AND U226
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U226 (
    .O(y[127]),
    .I0(a[7]),
    .I1(b[15])
  );
  //OR U226bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U226bar (
    .O(ybar[127]),
    .I0(abar[7]),
    .I1(bbar[15])
  );
  //AND U227
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U227 (
    .O(y[126]),
    .I0(a[7]),
    .I1(b[14])
  );
  //OR U227bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U227bar (
    .O(ybar[126]),
    .I0(abar[7]),
    .I1(bbar[14])
  );
  //AND U228
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U228 (
    .O(y[125]),
    .I0(a[7]),
    .I1(b[13])
  );
  //OR U228bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U228bar (
    .O(ybar[125]),
    .I0(abar[7]),
    .I1(bbar[13])
  );
  //AND U229
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U229 (
    .O(y[124]),
    .I0(a[7]),
    .I1(b[12])
  );
  //OR U229bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U229bar (
    .O(ybar[124]),
    .I0(abar[7]),
    .I1(bbar[12])
  );
  //AND U230
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U230 (
    .O(y[123]),
    .I0(a[7]),
    .I1(b[11])
  );
  //OR U230bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U230bar (
    .O(ybar[123]),
    .I0(abar[7]),
    .I1(bbar[11])
  );
  //AND U231
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U231 (
    .O(y[122]),
    .I0(a[7]),
    .I1(b[10])
  );
  //OR U231bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U231bar (
    .O(ybar[122]),
    .I0(abar[7]),
    .I1(bbar[10])
  );
  //AND U232
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U232 (
    .O(y[121]),
    .I0(a[7]),
    .I1(b[9])
  );
  //OR U232bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U232bar (
    .O(ybar[121]),
    .I0(abar[7]),
    .I1(bbar[9])
  );
  //AND U233
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U233 (
    .O(y[120]),
    .I0(a[7]),
    .I1(b[8])
  );
  //OR U233bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U233bar (
    .O(ybar[120]),
    .I0(abar[7]),
    .I1(bbar[8])
  );
  //AND U234
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U234 (
    .O(y[11]),
    .I0(b[11]),
    .I1(a[0])
  );
  //OR U234bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U234bar (
    .O(ybar[11]),
    .I0(bbar[11]),
    .I1(abar[0])
  );
  //AND U235
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U235 (
    .O(y[119]),
    .I0(a[7]),
    .I1(b[7])
  );
  //OR U235bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U235bar (
    .O(ybar[119]),
    .I0(abar[7]),
    .I1(bbar[7])
  );
  //AND U236
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U236 (
    .O(y[118]),
    .I0(a[7]),
    .I1(b[6])
  );
  //OR U236bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U236bar (
    .O(ybar[118]),
    .I0(abar[7]),
    .I1(bbar[6])
  );
  //AND U237
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U237 (
    .O(y[117]),
    .I0(a[7]),
    .I1(b[5])
  );
  //OR U237bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U237bar (
    .O(ybar[117]),
    .I0(abar[7]),
    .I1(bbar[5])
  );
  //AND U238
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U238 (
    .O(y[116]),
    .I0(a[7]),
    .I1(b[4])
  );
  //OR U238bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U238bar (
    .O(ybar[116]),
    .I0(abar[7]),
    .I1(bbar[4])
  );
  //AND U239
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U239 (
    .O(y[115]),
    .I0(a[7]),
    .I1(b[3])
  );
  //OR U239bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U239bar (
    .O(ybar[115]),
    .I0(abar[7]),
    .I1(bbar[3])
  );
  //AND U240
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U240 (
    .O(y[114]),
    .I0(a[7]),
    .I1(b[2])
  );
  //OR U240bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U240bar (
    .O(ybar[114]),
    .I0(abar[7]),
    .I1(bbar[2])
  );
  //AND U241
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U241 (
    .O(y[113]),
    .I0(a[7]),
    .I1(b[1])
  );
  //OR U241bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U241bar (
    .O(ybar[113]),
    .I0(abar[7]),
    .I1(bbar[1])
  );
  //AND U242
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U242 (
    .O(y[112]),
    .I0(a[7]),
    .I1(b[0])
  );
  //OR U242bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U242bar (
    .O(ybar[112]),
    .I0(abar[7]),
    .I1(bbar[0])
  );
  //AND U243
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U243 (
    .O(y[111]),
    .I0(b[15]),
    .I1(a[6])
  );
  //OR U243bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U243bar (
    .O(ybar[111]),
    .I0(bbar[15]),
    .I1(abar[6])
  );
  //AND U244
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U244 (
    .O(y[110]),
    .I0(b[14]),
    .I1(a[6])
  );
  //OR U244bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U244bar (
    .O(ybar[110]),
    .I0(bbar[14]),
    .I1(abar[6])
  );
  //AND U245
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U245 (
    .O(y[10]),
    .I0(b[10]),
    .I1(a[0])
  );
  //OR U245bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U245bar (
    .O(ybar[10]),
    .I0(bbar[10]),
    .I1(abar[0])
  );
  //AND U246
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U246 (
    .O(y[109]),
    .I0(b[13]),
    .I1(a[6])
  );
  //OR U246bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U246bar (
    .O(ybar[109]),
    .I0(bbar[13]),
    .I1(abar[6])
  );
  //AND U247
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U247 (
    .O(y[108]),
    .I0(b[12]),
    .I1(a[6])
  );
  //OR U247bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U247bar (
    .O(ybar[108]),
    .I0(bbar[12]),
    .I1(abar[6])
  );
  //AND U248
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U248 (
    .O(y[107]),
    .I0(b[11]),
    .I1(a[6])
  );
  //OR U248bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U248bar (
    .O(ybar[107]),
    .I0(bbar[11]),
    .I1(abar[6])
  );
  //AND U249
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U249 (
    .O(y[106]),
    .I0(b[10]),
    .I1(a[6])
  );
  //OR U249bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U249bar (
    .O(ybar[106]),
    .I0(bbar[10]),
    .I1(abar[6])
  );
  //AND U250
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U250 (
    .O(y[105]),
    .I0(a[6]),
    .I1(b[9])
  );
  //OR U250bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U250bar (
    .O(ybar[105]),
    .I0(abar[6]),
    .I1(bbar[9])
  );
  //AND U251
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U251 (
    .O(y[104]),
    .I0(b[8]),
    .I1(a[6])
  );
  //OR U251bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U251bar (
    .O(ybar[104]),
    .I0(bbar[8]),
    .I1(abar[6])
  );
  //AND U252
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U252 (
    .O(y[103]),
    .I0(b[7]),
    .I1(a[6])
  );
  //OR U252bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U252bar (
    .O(ybar[103]),
    .I0(bbar[7]),
    .I1(abar[6])
  );
  //AND U253
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U253 (
    .O(y[102]),
    .I0(b[6]),
    .I1(a[6])
  );
  //OR U253bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U253bar (
    .O(ybar[102]),
    .I0(bbar[6]),
    .I1(abar[6])
  );
  //AND U254
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U254 (
    .O(y[101]),
    .I0(b[5]),
    .I1(a[6])
  );
  //OR U254bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U254bar (
    .O(ybar[101]),
    .I0(bbar[5]),
    .I1(abar[6])
  );
  //AND U255
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U255 (
    .O(y[100]),
    .I0(b[4]),
    .I1(a[6])
  );
  //OR U255bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U255bar (
    .O(ybar[100]),
    .I0(bbar[4]),
    .I1(abar[6])
  );
  //AND U256
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U256 (
    .O(y[0]),
    .I0(b[0]),
    .I1(a[0])
  );
  //OR U256bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U256bar (
    .O(ybar[0]),
    .I0(bbar[0]),
    .I1(abar[0])
  );
endmodule

module decode_1 ( in, out );

  input wire [7:0] in;
//input_done

  output wire [255:0] out;
//output_done

  wire [15:0] level1;
  wire [31:0] level2;
//wire_done

  CD2_4 cd_l1_1 ( .a(in[1]), .b(in[0]), .y(level1[3:0]) );
  CD2_3 cd_l1_2 ( .a(in[3]), .b(in[2]), .y(level1[7:4]) );
  CD2_2 cd_l1_3 ( .a(in[5]), .b(in[4]), .y(level1[11:8]) );
  CD2_1 cd_l1_4 ( .a(in[7]), .b(in[6]), .y(level1[15:12]) );
  CD4_2 cd_l2_1 ( .a(level1[7:4]), .b(level1[3:0]), .y(level2[15:0]) );
  CD4_1 cd_l2_2 ( .a(level1[15:12]), .b(level1[11:8]), .y(level2[31:16]) );
  CD16_1 cd_l3 ( .a(level2[31:16]), .b(level2[15:0]), .y(out) );
endmodule

module encode_1 ( in, out );

  input wire [255:0] in;
  wire [255:0] inbar;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
  assign inbar[8] = ~in[8];
  assign inbar[9] = ~in[9];
  assign inbar[10] = ~in[10];
  assign inbar[11] = ~in[11];
  assign inbar[12] = ~in[12];
  assign inbar[13] = ~in[13];
  assign inbar[14] = ~in[14];
  assign inbar[15] = ~in[15];
  assign inbar[16] = ~in[16];
  assign inbar[17] = ~in[17];
  assign inbar[18] = ~in[18];
  assign inbar[19] = ~in[19];
  assign inbar[20] = ~in[20];
  assign inbar[21] = ~in[21];
  assign inbar[22] = ~in[22];
  assign inbar[23] = ~in[23];
  assign inbar[24] = ~in[24];
  assign inbar[25] = ~in[25];
  assign inbar[26] = ~in[26];
  assign inbar[27] = ~in[27];
  assign inbar[28] = ~in[28];
  assign inbar[29] = ~in[29];
  assign inbar[30] = ~in[30];
  assign inbar[31] = ~in[31];
  assign inbar[32] = ~in[32];
  assign inbar[33] = ~in[33];
  assign inbar[34] = ~in[34];
  assign inbar[35] = ~in[35];
  assign inbar[36] = ~in[36];
  assign inbar[37] = ~in[37];
  assign inbar[38] = ~in[38];
  assign inbar[39] = ~in[39];
  assign inbar[40] = ~in[40];
  assign inbar[41] = ~in[41];
  assign inbar[42] = ~in[42];
  assign inbar[43] = ~in[43];
  assign inbar[44] = ~in[44];
  assign inbar[45] = ~in[45];
  assign inbar[46] = ~in[46];
  assign inbar[47] = ~in[47];
  assign inbar[48] = ~in[48];
  assign inbar[49] = ~in[49];
  assign inbar[50] = ~in[50];
  assign inbar[51] = ~in[51];
  assign inbar[52] = ~in[52];
  assign inbar[53] = ~in[53];
  assign inbar[54] = ~in[54];
  assign inbar[55] = ~in[55];
  assign inbar[56] = ~in[56];
  assign inbar[57] = ~in[57];
  assign inbar[58] = ~in[58];
  assign inbar[59] = ~in[59];
  assign inbar[60] = ~in[60];
  assign inbar[61] = ~in[61];
  assign inbar[62] = ~in[62];
  assign inbar[63] = ~in[63];
  assign inbar[64] = ~in[64];
  assign inbar[65] = ~in[65];
  assign inbar[66] = ~in[66];
  assign inbar[67] = ~in[67];
  assign inbar[68] = ~in[68];
  assign inbar[69] = ~in[69];
  assign inbar[70] = ~in[70];
  assign inbar[71] = ~in[71];
  assign inbar[72] = ~in[72];
  assign inbar[73] = ~in[73];
  assign inbar[74] = ~in[74];
  assign inbar[75] = ~in[75];
  assign inbar[76] = ~in[76];
  assign inbar[77] = ~in[77];
  assign inbar[78] = ~in[78];
  assign inbar[79] = ~in[79];
  assign inbar[80] = ~in[80];
  assign inbar[81] = ~in[81];
  assign inbar[82] = ~in[82];
  assign inbar[83] = ~in[83];
  assign inbar[84] = ~in[84];
  assign inbar[85] = ~in[85];
  assign inbar[86] = ~in[86];
  assign inbar[87] = ~in[87];
  assign inbar[88] = ~in[88];
  assign inbar[89] = ~in[89];
  assign inbar[90] = ~in[90];
  assign inbar[91] = ~in[91];
  assign inbar[92] = ~in[92];
  assign inbar[93] = ~in[93];
  assign inbar[94] = ~in[94];
  assign inbar[95] = ~in[95];
  assign inbar[96] = ~in[96];
  assign inbar[97] = ~in[97];
  assign inbar[98] = ~in[98];
  assign inbar[99] = ~in[99];
  assign inbar[100] = ~in[100];
  assign inbar[101] = ~in[101];
  assign inbar[102] = ~in[102];
  assign inbar[103] = ~in[103];
  assign inbar[104] = ~in[104];
  assign inbar[105] = ~in[105];
  assign inbar[106] = ~in[106];
  assign inbar[107] = ~in[107];
  assign inbar[108] = ~in[108];
  assign inbar[109] = ~in[109];
  assign inbar[110] = ~in[110];
  assign inbar[111] = ~in[111];
  assign inbar[112] = ~in[112];
  assign inbar[113] = ~in[113];
  assign inbar[114] = ~in[114];
  assign inbar[115] = ~in[115];
  assign inbar[116] = ~in[116];
  assign inbar[117] = ~in[117];
  assign inbar[118] = ~in[118];
  assign inbar[119] = ~in[119];
  assign inbar[120] = ~in[120];
  assign inbar[121] = ~in[121];
  assign inbar[122] = ~in[122];
  assign inbar[123] = ~in[123];
  assign inbar[124] = ~in[124];
  assign inbar[125] = ~in[125];
  assign inbar[126] = ~in[126];
  assign inbar[127] = ~in[127];
  assign inbar[128] = ~in[128];
  assign inbar[129] = ~in[129];
  assign inbar[130] = ~in[130];
  assign inbar[131] = ~in[131];
  assign inbar[132] = ~in[132];
  assign inbar[133] = ~in[133];
  assign inbar[134] = ~in[134];
  assign inbar[135] = ~in[135];
  assign inbar[136] = ~in[136];
  assign inbar[137] = ~in[137];
  assign inbar[138] = ~in[138];
  assign inbar[139] = ~in[139];
  assign inbar[140] = ~in[140];
  assign inbar[141] = ~in[141];
  assign inbar[142] = ~in[142];
  assign inbar[143] = ~in[143];
  assign inbar[144] = ~in[144];
  assign inbar[145] = ~in[145];
  assign inbar[146] = ~in[146];
  assign inbar[147] = ~in[147];
  assign inbar[148] = ~in[148];
  assign inbar[149] = ~in[149];
  assign inbar[150] = ~in[150];
  assign inbar[151] = ~in[151];
  assign inbar[152] = ~in[152];
  assign inbar[153] = ~in[153];
  assign inbar[154] = ~in[154];
  assign inbar[155] = ~in[155];
  assign inbar[156] = ~in[156];
  assign inbar[157] = ~in[157];
  assign inbar[158] = ~in[158];
  assign inbar[159] = ~in[159];
  assign inbar[160] = ~in[160];
  assign inbar[161] = ~in[161];
  assign inbar[162] = ~in[162];
  assign inbar[163] = ~in[163];
  assign inbar[164] = ~in[164];
  assign inbar[165] = ~in[165];
  assign inbar[166] = ~in[166];
  assign inbar[167] = ~in[167];
  assign inbar[168] = ~in[168];
  assign inbar[169] = ~in[169];
  assign inbar[170] = ~in[170];
  assign inbar[171] = ~in[171];
  assign inbar[172] = ~in[172];
  assign inbar[173] = ~in[173];
  assign inbar[174] = ~in[174];
  assign inbar[175] = ~in[175];
  assign inbar[176] = ~in[176];
  assign inbar[177] = ~in[177];
  assign inbar[178] = ~in[178];
  assign inbar[179] = ~in[179];
  assign inbar[180] = ~in[180];
  assign inbar[181] = ~in[181];
  assign inbar[182] = ~in[182];
  assign inbar[183] = ~in[183];
  assign inbar[184] = ~in[184];
  assign inbar[185] = ~in[185];
  assign inbar[186] = ~in[186];
  assign inbar[187] = ~in[187];
  assign inbar[188] = ~in[188];
  assign inbar[189] = ~in[189];
  assign inbar[190] = ~in[190];
  assign inbar[191] = ~in[191];
  assign inbar[192] = ~in[192];
  assign inbar[193] = ~in[193];
  assign inbar[194] = ~in[194];
  assign inbar[195] = ~in[195];
  assign inbar[196] = ~in[196];
  assign inbar[197] = ~in[197];
  assign inbar[198] = ~in[198];
  assign inbar[199] = ~in[199];
  assign inbar[200] = ~in[200];
  assign inbar[201] = ~in[201];
  assign inbar[202] = ~in[202];
  assign inbar[203] = ~in[203];
  assign inbar[204] = ~in[204];
  assign inbar[205] = ~in[205];
  assign inbar[206] = ~in[206];
  assign inbar[207] = ~in[207];
  assign inbar[208] = ~in[208];
  assign inbar[209] = ~in[209];
  assign inbar[210] = ~in[210];
  assign inbar[211] = ~in[211];
  assign inbar[212] = ~in[212];
  assign inbar[213] = ~in[213];
  assign inbar[214] = ~in[214];
  assign inbar[215] = ~in[215];
  assign inbar[216] = ~in[216];
  assign inbar[217] = ~in[217];
  assign inbar[218] = ~in[218];
  assign inbar[219] = ~in[219];
  assign inbar[220] = ~in[220];
  assign inbar[221] = ~in[221];
  assign inbar[222] = ~in[222];
  assign inbar[223] = ~in[223];
  assign inbar[224] = ~in[224];
  assign inbar[225] = ~in[225];
  assign inbar[226] = ~in[226];
  assign inbar[227] = ~in[227];
  assign inbar[228] = ~in[228];
  assign inbar[229] = ~in[229];
  assign inbar[230] = ~in[230];
  assign inbar[231] = ~in[231];
  assign inbar[232] = ~in[232];
  assign inbar[233] = ~in[233];
  assign inbar[234] = ~in[234];
  assign inbar[235] = ~in[235];
  assign inbar[236] = ~in[236];
  assign inbar[237] = ~in[237];
  assign inbar[238] = ~in[238];
  assign inbar[239] = ~in[239];
  assign inbar[240] = ~in[240];
  assign inbar[241] = ~in[241];
  assign inbar[242] = ~in[242];
  assign inbar[243] = ~in[243];
  assign inbar[244] = ~in[244];
  assign inbar[245] = ~in[245];
  assign inbar[246] = ~in[246];
  assign inbar[247] = ~in[247];
  assign inbar[248] = ~in[248];
  assign inbar[249] = ~in[249];
  assign inbar[250] = ~in[250];
  assign inbar[251] = ~in[251];
  assign inbar[252] = ~in[252];
  assign inbar[253] = ~in[253];
  assign inbar[254] = ~in[254];
  assign inbar[255] = ~in[255];
//input_done

  output wire [7:0] out;
  wire [7:0] outbar;
//output_done

  wire in_81;
  wire in_80;
  wire in_79;
  wire in_78;
  wire in_77;
  wire in_76;
  wire in_75;
  wire in_74;
  wire in_73;
  wire in_72;
  wire in_71;
  wire in_70;
  wire in_69;
  wire in_68;
  wire in_67;
  wire in_66;
  wire in_65;
  wire in_64;
  wire in_63;
  wire in_62;
  wire in_61;
  wire in_60;
  wire in_59;
  wire in_58;
  wire in_57;
  wire in_56;
  wire in_55;
  wire in_54;
  wire in_53;
  wire in_52;
  wire in_51;
  wire in_50;
  wire in_49;
  wire in_48;
  wire in_47;
  wire in_46;
  wire in_45;
  wire in_44;
  wire in_43;
  wire in_42;
  wire in_41;
  wire in_40;
  wire in_39;
  wire in_38;
  wire in_37;
  wire in_36;
  wire in_35;
  wire in_34;
  wire in_33;
  wire in_32;
  wire in_31;
  wire in_30;
  wire in_29;
  wire in_28;
  wire in_27;
  wire in_26;
  wire in_25;
  wire in_24;
  wire in_23;
  wire in_22;
  wire in_21;
  wire in_20;
  wire in_19;
  wire in_18;
  wire in_17;
  wire in_16;
  wire in_15;
  wire in_14;
  wire in_13;
  wire in_12;
  wire in_11;
  wire in_10;
  wire in_9;
  wire in_8;
  wire in_7;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_3;
  wire in_2;
  wire in_1;
  wire in_0;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire in_81bar;
  wire in_80bar;
  wire in_79bar;
  wire in_78bar;
  wire in_77bar;
  wire in_76bar;
  wire in_75bar;
  wire in_74bar;
  wire in_73bar;
  wire in_72bar;
  wire in_71bar;
  wire in_70bar;
  wire in_69bar;
  wire in_68bar;
  wire in_67bar;
  wire in_66bar;
  wire in_65bar;
  wire in_64bar;
  wire in_63bar;
  wire in_62bar;
  wire in_61bar;
  wire in_60bar;
  wire in_59bar;
  wire in_58bar;
  wire in_57bar;
  wire in_56bar;
  wire in_55bar;
  wire in_54bar;
  wire in_53bar;
  wire in_52bar;
  wire in_51bar;
  wire in_50bar;
  wire in_49bar;
  wire in_48bar;
  wire in_47bar;
  wire in_46bar;
  wire in_45bar;
  wire in_44bar;
  wire in_43bar;
  wire in_42bar;
  wire in_41bar;
  wire in_40bar;
  wire in_39bar;
  wire in_38bar;
  wire in_37bar;
  wire in_36bar;
  wire in_35bar;
  wire in_34bar;
  wire in_33bar;
  wire in_32bar;
  wire in_31bar;
  wire in_30bar;
  wire in_29bar;
  wire in_28bar;
  wire in_27bar;
  wire in_26bar;
  wire in_25bar;
  wire in_24bar;
  wire in_23bar;
  wire in_22bar;
  wire in_21bar;
  wire in_20bar;
  wire in_19bar;
  wire in_18bar;
  wire in_17bar;
  wire in_16bar;
  wire in_15bar;
  wire in_14bar;
  wire in_13bar;
  wire in_12bar;
  wire in_11bar;
  wire in_10bar;
  wire in_9bar;
  wire in_8bar;
  wire in_7bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_3bar;
  wire in_2bar;
  wire in_1bar;
  wire in_0bar;
  wire n487bar;
  wire n488bar;
  wire n489bar;
  wire n490bar;
  wire n491bar;
  wire n492bar;
  wire n493bar;
  wire n494bar;
  wire n495bar;
  wire n496bar;
  wire n497bar;
  wire n498bar;
  wire n499bar;
  wire n500bar;
  wire n501bar;
  wire n502bar;
  wire n503bar;
  wire n504bar;
  wire n505bar;
  wire n506bar;
  wire n507bar;
  wire n508bar;
  wire n509bar;
  wire n510bar;
  wire n511bar;
  wire n512bar;
  wire n513bar;
  wire n514bar;
  wire n515bar;
  wire n516bar;
  wire n517bar;
  wire n518bar;
  wire n519bar;
  wire n520bar;
  wire n521bar;
  wire n522bar;
  wire n523bar;
  wire n524bar;
  wire n525bar;
  wire n526bar;
  wire n527bar;
  wire n528bar;
  wire n529bar;
  wire n530bar;
  wire n531bar;
  wire n532bar;
  wire n533bar;
  wire n534bar;
  wire n535bar;
  wire n536bar;
  wire n537bar;
  wire n538bar;
  wire n539bar;
  wire n540bar;
  wire n541bar;
  wire n542bar;
  wire n543bar;
  wire n544bar;
  wire n545bar;
  wire n546bar;
  wire n547bar;
  wire n548bar;
  wire n549bar;
  wire n550bar;
  wire n551bar;
  wire n552bar;
  wire n553bar;
  wire n554bar;
  wire n555bar;
  wire n556bar;
  wire n557bar;
  wire n558bar;
  wire n559bar;
  wire n560bar;
  wire n561bar;
  wire n562bar;
  wire n563bar;
  wire n564bar;
  wire n565bar;
  wire n566bar;
  wire n567bar;
  wire n568bar;
  wire n569bar;
  wire n570bar;
  wire n571bar;
  wire n572bar;
  wire n573bar;
  wire n574bar;
  wire n575bar;
  wire n576bar;
  wire n577bar;
  wire n578bar;
  wire n579bar;
  wire n580bar;
  wire n581bar;
  wire n582bar;
  wire n583bar;
  wire n584bar;
  wire n585bar;
  wire n586bar;
  wire n587bar;
  wire n588bar;
  wire n589bar;
  wire n590bar;
  wire n591bar;
  wire n592bar;
  wire n593bar;
  wire n594bar;
  wire n595bar;
  wire n596bar;
  wire n597bar;
  wire n598bar;
  wire n599bar;
  wire n600bar;
  wire n601bar;
  wire n602bar;
  wire n603bar;
  wire n604bar;
  wire n605bar;
  wire n606bar;
  wire n607bar;
  wire n608bar;
  wire n609bar;
  wire n610bar;
  wire n611bar;
  wire n612bar;
  wire n613bar;
  wire n614bar;
  wire n615bar;
  wire n616bar;
  wire n617bar;
  wire n618bar;
  wire n619bar;
  wire n620bar;
  wire n621bar;
  wire n622bar;
  wire n623bar;
  wire n624bar;
  wire n625bar;
  wire n626bar;
  wire n627bar;
  wire n628bar;
  wire n629bar;
  wire n630bar;
  wire n631bar;
  wire n632bar;
  wire n633bar;
  wire n634bar;
  wire n635bar;
  wire n636bar;
  wire n637bar;
  wire n638bar;
  wire n639bar;
  wire n640bar;
  wire n641bar;
  wire n642bar;
  wire n643bar;
  wire n644bar;
  wire n645bar;
  wire n646bar;
  wire n647bar;
  wire n648bar;
  wire n649bar;
  wire n650bar;
  wire n651bar;
  wire n652bar;
  wire n653bar;
  wire n654bar;
  wire n655bar;
  wire n656bar;
  wire n657bar;
  wire n658bar;
  wire n659bar;
  wire n660bar;
  wire n661bar;
  wire n662bar;
  wire n663bar;
  wire n664bar;
  wire n665bar;
  wire n666bar;
  wire n667bar;
  wire n668bar;
  wire n669bar;
  wire n670bar;
  wire n671bar;
  wire n672bar;
  wire n673bar;
  wire n674bar;
  wire n675bar;
  wire n676bar;
  wire n677bar;
  wire n678bar;
  wire n679bar;
  wire n680bar;
  wire n681bar;
  wire n682bar;
  wire n683bar;
  wire n684bar;
  wire n685bar;
  wire n686bar;
  wire n687bar;
  wire n688bar;
  wire n689bar;
  wire n690bar;
  wire n691bar;
  wire n692bar;
  wire n693bar;
  wire n694bar;
  wire n695bar;
  wire n696bar;
  wire n697bar;
  wire n698bar;
  wire n699bar;
  wire n700bar;
  wire n701bar;
  wire n702bar;
  wire n703bar;
  wire n704bar;
  wire n705bar;
  wire n706bar;
  wire n707bar;
  wire n708bar;
  wire n709bar;
  wire n710bar;
  wire n711bar;
  wire n712bar;
  wire n713bar;
  wire n714bar;
  wire n715bar;
  wire n716bar;
  wire n717bar;
  wire n718bar;
  wire n719bar;
  wire n720bar;
  wire n721bar;
  wire n722bar;
  wire n723bar;
  wire n724bar;
  wire n725bar;
  wire n726bar;
  wire n727bar;
  wire n728bar;
  wire n729bar;
  wire n730bar;
  wire n731bar;
  wire n732bar;
  wire n733bar;
  wire n734bar;
  wire n735bar;
  wire n736bar;
  wire n737bar;
  wire n738bar;
  wire n739bar;
  wire n740bar;
  wire n741bar;
  wire n742bar;
  wire n743bar;
  wire n744bar;
  wire n745bar;
  wire n746bar;
  wire n747bar;
  wire n748bar;
  wire n749bar;
  wire n750bar;
  wire n751bar;
  wire n752bar;
  wire n753bar;
  wire n754bar;
  wire n755bar;
  wire n756bar;
  wire n757bar;
  wire n758bar;
  wire n759bar;
  wire n760bar;
  wire n761bar;
  wire n762bar;
  wire n763bar;
  wire n764bar;
  wire n765bar;
  wire n766bar;
  wire n767bar;
  wire n768bar;
  wire n769bar;
  wire n770bar;
  wire n771bar;
  wire n772bar;
  wire n773bar;
  wire n774bar;
  wire n775bar;
  wire n776bar;
  wire n777bar;
  wire n778bar;
  wire n779bar;
  wire n780bar;
  wire n781bar;
  wire n782bar;
  wire n783bar;
  wire n784bar;
  wire n785bar;
  wire n786bar;
  wire n787bar;
  wire n788bar;
  wire n789bar;
  wire n790bar;
  wire n791bar;
  wire n792bar;
  wire n793bar;
  wire n794bar;
  wire n795bar;
  wire n796bar;
  wire n797bar;
  wire n798bar;
  wire n799bar;
  wire n800bar;
  wire n801bar;
  wire n802bar;
  wire n803bar;
  wire n804bar;
  wire n805bar;
  wire n806bar;
  wire n807bar;
  wire n808bar;
  wire n809bar;
  wire n810bar;
  wire n811bar;
  wire n812bar;
  wire n813bar;
  wire n814bar;
  wire n815bar;
  wire n816bar;
  wire n817bar;
  wire n818bar;
  wire n819bar;
  wire n820bar;
  wire n821bar;
  wire n822bar;
  wire n823bar;
  wire n824bar;
  wire n825bar;
  wire n826bar;
  wire n827bar;
  wire n828bar;
  wire n829bar;
  wire n830bar;
  wire n831bar;
  wire n832bar;
  wire n833bar;
  wire n834bar;
  wire n835bar;
  wire n836bar;
  wire n837bar;
  wire n838bar;
  wire n839bar;
  wire n840bar;
  wire n841bar;
  wire n842bar;
  wire n843bar;
  wire n844bar;
  wire n845bar;
  wire n846bar;
  wire n847bar;
  wire n848bar;
  wire n849bar;
  wire n850bar;
  wire n851bar;
  wire n852bar;
  wire n853bar;
  wire n854bar;
  wire n855bar;
  wire n856bar;
  wire n857bar;
  wire n858bar;
  wire n859bar;
  wire n860bar;
  wire n861bar;
  wire n862bar;
  wire n863bar;
  wire n864bar;
  wire n865bar;
  wire n866bar;
  wire n867bar;
  wire n868bar;
  wire n869bar;
  wire n870bar;
  wire n871bar;
  wire n872bar;
  wire n873bar;
  wire n874bar;
  wire n875bar;
  wire n876bar;
  wire n877bar;
  wire n878bar;
  wire n879bar;
  wire n880bar;
  wire n881bar;
  wire n882bar;
  wire n883bar;
  wire n884bar;
  wire n885bar;
  wire n886bar;
  wire n887bar;
  wire n888bar;
  wire n889bar;
  wire n890bar;
  wire n891bar;
  wire n892bar;
  wire n893bar;
  wire n894bar;
  wire n895bar;
  wire n896bar;
  wire n897bar;
  wire n898bar;
  wire n899bar;
  wire n900bar;
  wire n901bar;
  wire n902bar;
  wire n903bar;
  wire n904bar;
  wire n905bar;
  wire n906bar;
  wire n907bar;
  wire n908bar;
  wire n909bar;
  wire n910bar;
  wire n911bar;
  wire n912bar;
  wire n913bar;
  wire n914bar;
  wire n915bar;
  wire n916bar;
  wire n917bar;
  wire n918bar;
  wire n919bar;
  wire n920bar;
  wire n921bar;
  wire n922bar;
  wire n923bar;
  wire n924bar;
  wire n925bar;
  wire n926bar;
  wire n927bar;
  wire n928bar;
  wire n929bar;
  wire n930bar;
  wire n931bar;
  wire n932bar;
  wire n933bar;
  wire n934bar;
  wire n935bar;
  wire n936bar;
  wire n937bar;
  wire n938bar;
  wire n939bar;
  wire n940bar;
  wire n941bar;
  wire n942bar;
  wire n943bar;
  wire n944bar;
  wire n945bar;
  wire n946bar;
  wire n947bar;
  wire n948bar;
  wire n949bar;
  wire n950bar;
  wire n951bar;
  wire n952bar;
  wire n953bar;
  wire n954bar;
  wire n955bar;
  wire n956bar;
  wire n957bar;
  wire n958bar;
  wire n959bar;
  wire n960bar;
  wire n961bar;
  wire n962bar;
  wire n963bar;
  wire n964bar;
  wire n965bar;
  wire n966bar;
  wire n967bar;
  wire n968bar;
  wire n969bar;
  wire n970bar;
  wire n971bar;
  wire n972bar;
//wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];
  //OR U1
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1 (
    .O(out[7]),
    .I0(n972),
    .I1(n971)
  );
  //AND U1bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1bar (
    .O(outbar[7]),
    .I0(n972bar),
    .I1(n971bar)
  );
  //OR U2
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2 (
    .O(n971),
    .I0(n970),
    .I1(n969)
  );
  //AND U2bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2bar (
    .O(n971bar),
    .I0(n970bar),
    .I1(n969bar)
  );
  //OR U3
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3 (
    .O(n969),
    .I0(n968),
    .I1(n967)
  );
  //AND U3bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3bar (
    .O(n969bar),
    .I0(n968bar),
    .I1(n967bar)
  );
  //OR U4
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4 (
    .O(n967),
    .I0(n966),
    .I1(n965)
  );
  //AND U4bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4bar (
    .O(n967bar),
    .I0(n966bar),
    .I1(n965bar)
  );
  //OR U5
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5 (
    .O(n968),
    .I0(n964),
    .I1(n963)
  );
  //AND U5bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5bar (
    .O(n968bar),
    .I0(n964bar),
    .I1(n963bar)
  );
  //OR U6
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6 (
    .O(n963),
    .I0(in[116]),
    .I1(n962)
  );
  //AND U6bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6bar (
    .O(n963bar),
    .I0(inbar[116]),
    .I1(n962bar)
  );
  //OR U7
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7 (
    .O(n970),
    .I0(n961),
    .I1(n960)
  );
  //AND U7bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7bar (
    .O(n970bar),
    .I0(n961bar),
    .I1(n960bar)
  );
  //OR U8
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8 (
    .O(n960),
    .I0(in[150]),
    .I1(in[127])
  );
  //AND U8bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8bar (
    .O(n960bar),
    .I0(inbar[150]),
    .I1(inbar[127])
  );
  //OR U9
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9 (
    .O(n961),
    .I0(in[160]),
    .I1(n959)
  );
  //AND U9bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9bar (
    .O(n961bar),
    .I0(inbar[160]),
    .I1(n959bar)
  );
  //OR U10
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10 (
    .O(n959),
    .I0(in[252]),
    .I1(in[168])
  );
  //AND U10bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10bar (
    .O(n959bar),
    .I0(inbar[252]),
    .I1(inbar[168])
  );
  //OR U11
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11 (
    .O(n972),
    .I0(n958),
    .I1(n957)
  );
  //AND U11bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11bar (
    .O(n972bar),
    .I0(n958bar),
    .I1(n957bar)
  );
  //OR U12
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12 (
    .O(n957),
    .I0(n956),
    .I1(n955)
  );
  //AND U12bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12bar (
    .O(n957bar),
    .I0(n956bar),
    .I1(n955bar)
  );
  //OR U13
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13 (
    .O(n955),
    .I0(in_17),
    .I1(in[96])
  );
  //AND U13bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13bar (
    .O(n955bar),
    .I0(in_17bar),
    .I1(inbar[96])
  );
  //OR U14
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14 (
    .O(n956),
    .I0(in_23),
    .I1(n954)
  );
  //AND U14bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14bar (
    .O(n956bar),
    .I0(in_23bar),
    .I1(n954bar)
  );
  //OR U15
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15 (
    .O(n954),
    .I0(in_31),
    .I1(in_26)
  );
  //AND U15bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15bar (
    .O(n954bar),
    .I0(in_31bar),
    .I1(in_26bar)
  );
  //OR U16
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16 (
    .O(n958),
    .I0(n953),
    .I1(n952)
  );
  //AND U16bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16bar (
    .O(n958bar),
    .I0(n953bar),
    .I1(n952bar)
  );
  //OR U17
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U17 (
    .O(n952),
    .I0(in_58),
    .I1(in_4)
  );
  //AND U17bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U17bar (
    .O(n952bar),
    .I0(in_58bar),
    .I1(in_4bar)
  );
  //OR U18
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U18 (
    .O(n953),
    .I0(in_59),
    .I1(n951)
  );
  //AND U18bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U18bar (
    .O(n953bar),
    .I0(in_59bar),
    .I1(n951bar)
  );
  //OR U19
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U19 (
    .O(n951),
    .I0(in_71),
    .I1(in_62)
  );
  //AND U19bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U19bar (
    .O(n951bar),
    .I0(in_71bar),
    .I1(in_62bar)
  );
  //OR U20
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U20 (
    .O(out[6]),
    .I0(n950),
    .I1(n949)
  );
  //AND U20bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U20bar (
    .O(outbar[6]),
    .I0(n950bar),
    .I1(n949bar)
  );
  //OR U21
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U21 (
    .O(n949),
    .I0(n948),
    .I1(n947)
  );
  //AND U21bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U21bar (
    .O(n949bar),
    .I0(n948bar),
    .I1(n947bar)
  );
  //OR U22
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U22 (
    .O(n947),
    .I0(n946),
    .I1(n945)
  );
  //AND U22bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U22bar (
    .O(n947bar),
    .I0(n946bar),
    .I1(n945bar)
  );
  //OR U23
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U23 (
    .O(n945),
    .I0(n944),
    .I1(n943)
  );
  //AND U23bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U23bar (
    .O(n945bar),
    .I0(n944bar),
    .I1(n943bar)
  );
  //OR U24
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U24 (
    .O(n946),
    .I0(n942),
    .I1(n941)
  );
  //AND U24bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U24bar (
    .O(n946bar),
    .I0(n942bar),
    .I1(n941bar)
  );
  //OR U25
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U25 (
    .O(n941),
    .I0(in[101]),
    .I1(n940)
  );
  //AND U25bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U25bar (
    .O(n941bar),
    .I0(inbar[101]),
    .I1(n940bar)
  );
  //OR U26
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U26 (
    .O(n948),
    .I0(n939),
    .I1(n938)
  );
  //AND U26bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U26bar (
    .O(n948bar),
    .I0(n939bar),
    .I1(n938bar)
  );
  //OR U27
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U27 (
    .O(n938),
    .I0(in[114]),
    .I1(in[104])
  );
  //AND U27bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U27bar (
    .O(n938bar),
    .I0(inbar[114]),
    .I1(inbar[104])
  );
  //OR U28
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U28 (
    .O(n939),
    .I0(in[128]),
    .I1(n937)
  );
  //AND U28bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U28bar (
    .O(n939bar),
    .I0(inbar[128]),
    .I1(n937bar)
  );
  //OR U29
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U29 (
    .O(n937),
    .I0(in[136]),
    .I1(in[134])
  );
  //AND U29bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U29bar (
    .O(n937bar),
    .I0(inbar[136]),
    .I1(inbar[134])
  );
  //OR U30
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U30 (
    .O(n950),
    .I0(n936),
    .I1(n935)
  );
  //AND U30bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U30bar (
    .O(n950bar),
    .I0(n936bar),
    .I1(n935bar)
  );
  //OR U31
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U31 (
    .O(n935),
    .I0(n934),
    .I1(n933)
  );
  //AND U31bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U31bar (
    .O(n935bar),
    .I0(n934bar),
    .I1(n933bar)
  );
  //OR U32
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U32 (
    .O(n933),
    .I0(in[177]),
    .I1(in[164])
  );
  //AND U32bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U32bar (
    .O(n933bar),
    .I0(inbar[177]),
    .I1(inbar[164])
  );
  //OR U33
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U33 (
    .O(n934),
    .I0(in[212]),
    .I1(n932)
  );
  //AND U33bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U33bar (
    .O(n934bar),
    .I0(inbar[212]),
    .I1(n932bar)
  );
  //OR U34
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U34 (
    .O(n932),
    .I0(in[248]),
    .I1(in[221])
  );
  //AND U34bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U34bar (
    .O(n932bar),
    .I0(inbar[248]),
    .I1(inbar[221])
  );
  //OR U35
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U35 (
    .O(n936),
    .I0(n931),
    .I1(n930)
  );
  //AND U35bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U35bar (
    .O(n936bar),
    .I0(n931bar),
    .I1(n930bar)
  );
  //OR U36
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U36 (
    .O(n930),
    .I0(in_18),
    .I1(in[93])
  );
  //AND U36bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U36bar (
    .O(n930bar),
    .I0(in_18bar),
    .I1(inbar[93])
  );
  //OR U37
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U37 (
    .O(n931),
    .I0(in_31),
    .I1(n929)
  );
  //AND U37bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U37bar (
    .O(n931bar),
    .I0(in_31bar),
    .I1(n929bar)
  );
  //OR U38
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U38 (
    .O(n929),
    .I0(in_7),
    .I1(in_39)
  );
  //AND U38bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U38bar (
    .O(n929bar),
    .I0(in_7bar),
    .I1(in_39bar)
  );
  //OR U39
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U39 (
    .O(out[5]),
    .I0(n928),
    .I1(n927)
  );
  //AND U39bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U39bar (
    .O(outbar[5]),
    .I0(n928bar),
    .I1(n927bar)
  );
  //OR U40
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U40 (
    .O(n927),
    .I0(n926),
    .I1(n925)
  );
  //AND U40bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U40bar (
    .O(n927bar),
    .I0(n926bar),
    .I1(n925bar)
  );
  //OR U41
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U41 (
    .O(n925),
    .I0(n924),
    .I1(n923)
  );
  //AND U41bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U41bar (
    .O(n925bar),
    .I0(n924bar),
    .I1(n923bar)
  );
  //OR U42
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U42 (
    .O(n923),
    .I0(n922),
    .I1(n921)
  );
  //AND U42bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U42bar (
    .O(n923bar),
    .I0(n922bar),
    .I1(n921bar)
  );
  //OR U43
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U43 (
    .O(n924),
    .I0(n940),
    .I1(n920)
  );
  //AND U43bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U43bar (
    .O(n924bar),
    .I0(n940bar),
    .I1(n920bar)
  );
  //OR U44
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U44 (
    .O(n920),
    .I0(in[111]),
    .I1(n919)
  );
  //AND U44bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U44bar (
    .O(n920bar),
    .I0(inbar[111]),
    .I1(n919bar)
  );
  //OR U45
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U45 (
    .O(n940),
    .I0(n918),
    .I1(n917)
  );
  //AND U45bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U45bar (
    .O(n940bar),
    .I0(n918bar),
    .I1(n917bar)
  );
  //OR U46
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U46 (
    .O(n917),
    .I0(n916),
    .I1(n915)
  );
  //AND U46bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U46bar (
    .O(n917bar),
    .I0(n916bar),
    .I1(n915bar)
  );
  //OR U47
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U47 (
    .O(n915),
    .I0(n914),
    .I1(n913)
  );
  //AND U47bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U47bar (
    .O(n915bar),
    .I0(n914bar),
    .I1(n913bar)
  );
  //OR U48
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U48 (
    .O(n913),
    .I0(in[140]),
    .I1(in[131])
  );
  //AND U48bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U48bar (
    .O(n913bar),
    .I0(inbar[140]),
    .I1(inbar[131])
  );
  //OR U49
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U49 (
    .O(n914),
    .I0(in[160]),
    .I1(in[144])
  );
  //AND U49bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U49bar (
    .O(n914bar),
    .I0(inbar[160]),
    .I1(inbar[144])
  );
  //OR U50
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U50 (
    .O(n916),
    .I0(n912),
    .I1(n911)
  );
  //AND U50bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U50bar (
    .O(n916bar),
    .I0(n912bar),
    .I1(n911bar)
  );
  //OR U51
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U51 (
    .O(n911),
    .I0(in[179]),
    .I1(in[174])
  );
  //AND U51bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U51bar (
    .O(n911bar),
    .I0(inbar[179]),
    .I1(inbar[174])
  );
  //OR U52
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U52 (
    .O(n912),
    .I0(in[188]),
    .I1(in[184])
  );
  //AND U52bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U52bar (
    .O(n912bar),
    .I0(inbar[188]),
    .I1(inbar[184])
  );
  //OR U53
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U53 (
    .O(n918),
    .I0(n910),
    .I1(n909)
  );
  //AND U53bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U53bar (
    .O(n918bar),
    .I0(n910bar),
    .I1(n909bar)
  );
  //OR U54
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U54 (
    .O(n909),
    .I0(n908),
    .I1(n907)
  );
  //AND U54bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U54bar (
    .O(n909bar),
    .I0(n908bar),
    .I1(n907bar)
  );
  //OR U55
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U55 (
    .O(n907),
    .I0(in[216]),
    .I1(in[200])
  );
  //AND U55bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U55bar (
    .O(n907bar),
    .I0(inbar[216]),
    .I1(inbar[200])
  );
  //OR U56
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U56 (
    .O(n908),
    .I0(in[228]),
    .I1(in[224])
  );
  //AND U56bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U56bar (
    .O(n908bar),
    .I0(inbar[228]),
    .I1(inbar[224])
  );
  //OR U57
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U57 (
    .O(n910),
    .I0(n906),
    .I1(n905)
  );
  //AND U57bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U57bar (
    .O(n910bar),
    .I0(n906bar),
    .I1(n905bar)
  );
  //OR U58
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U58 (
    .O(n905),
    .I0(in[247]),
    .I1(in[235])
  );
  //AND U58bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U58bar (
    .O(n905bar),
    .I0(inbar[247]),
    .I1(inbar[235])
  );
  //OR U59
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U59 (
    .O(n906),
    .I0(in_42),
    .I1(in[83])
  );
  //AND U59bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U59bar (
    .O(n906bar),
    .I0(in_42bar),
    .I1(inbar[83])
  );
  //OR U60
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U60 (
    .O(n926),
    .I0(n904),
    .I1(n903)
  );
  //AND U60bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U60bar (
    .O(n926bar),
    .I0(n904bar),
    .I1(n903bar)
  );
  //OR U61
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U61 (
    .O(n903),
    .I0(in[166]),
    .I1(in[123])
  );
  //AND U61bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U61bar (
    .O(n903bar),
    .I0(inbar[166]),
    .I1(inbar[123])
  );
  //OR U62
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U62 (
    .O(n904),
    .I0(in[170]),
    .I1(n902)
  );
  //AND U62bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U62bar (
    .O(n904bar),
    .I0(inbar[170]),
    .I1(n902bar)
  );
  //OR U63
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U63 (
    .O(n902),
    .I0(in[194]),
    .I1(in[183])
  );
  //AND U63bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U63bar (
    .O(n902bar),
    .I0(inbar[194]),
    .I1(inbar[183])
  );
  //OR U64
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U64 (
    .O(n928),
    .I0(n901),
    .I1(n900)
  );
  //AND U64bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U64bar (
    .O(n928bar),
    .I0(n901bar),
    .I1(n900bar)
  );
  //OR U65
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U65 (
    .O(n900),
    .I0(n899),
    .I1(n898)
  );
  //AND U65bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U65bar (
    .O(n900bar),
    .I0(n899bar),
    .I1(n898bar)
  );
  //OR U66
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U66 (
    .O(n898),
    .I0(in[241]),
    .I1(in[238])
  );
  //AND U66bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U66bar (
    .O(n898bar),
    .I0(inbar[241]),
    .I1(inbar[238])
  );
  //OR U67
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U67 (
    .O(n899),
    .I0(in[250]),
    .I1(n897)
  );
  //AND U67bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U67bar (
    .O(n899bar),
    .I0(inbar[250]),
    .I1(n897bar)
  );
  //OR U68
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U68 (
    .O(n897),
    .I0(in_24),
    .I1(in[84])
  );
  //AND U68bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U68bar (
    .O(n897bar),
    .I0(in_24bar),
    .I1(inbar[84])
  );
  //OR U69
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U69 (
    .O(n901),
    .I0(n896),
    .I1(n895)
  );
  //AND U69bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U69bar (
    .O(n901bar),
    .I0(n896bar),
    .I1(n895bar)
  );
  //OR U70
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U70 (
    .O(n895),
    .I0(in_41),
    .I1(in_29)
  );
  //AND U70bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U70bar (
    .O(n895bar),
    .I0(in_41bar),
    .I1(in_29bar)
  );
  //OR U71
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U71 (
    .O(n896),
    .I0(in_66),
    .I1(n894)
  );
  //AND U71bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U71bar (
    .O(n896bar),
    .I0(in_66bar),
    .I1(n894bar)
  );
  //OR U72
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U72 (
    .O(n894),
    .I0(in_76),
    .I1(in_71)
  );
  //AND U72bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U72bar (
    .O(n894bar),
    .I0(in_76bar),
    .I1(in_71bar)
  );
  //OR U73
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U73 (
    .O(out[4]),
    .I0(n893),
    .I1(n892)
  );
  //AND U73bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U73bar (
    .O(outbar[4]),
    .I0(n893bar),
    .I1(n892bar)
  );
  //OR U74
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U74 (
    .O(n892),
    .I0(n891),
    .I1(n890)
  );
  //AND U74bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U74bar (
    .O(n892bar),
    .I0(n891bar),
    .I1(n890bar)
  );
  //OR U75
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U75 (
    .O(n890),
    .I0(n889),
    .I1(n888)
  );
  //AND U75bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U75bar (
    .O(n890bar),
    .I0(n889bar),
    .I1(n888bar)
  );
  //OR U76
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U76 (
    .O(n888),
    .I0(n922),
    .I1(n887)
  );
  //AND U76bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U76bar (
    .O(n888bar),
    .I0(n922bar),
    .I1(n887bar)
  );
  //OR U77
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U77 (
    .O(n922),
    .I0(n886),
    .I1(n885)
  );
  //AND U77bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U77bar (
    .O(n922bar),
    .I0(n886bar),
    .I1(n885bar)
  );
  //OR U78
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U78 (
    .O(n885),
    .I0(n884),
    .I1(n883)
  );
  //AND U78bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U78bar (
    .O(n885bar),
    .I0(n884bar),
    .I1(n883bar)
  );
  //OR U79
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U79 (
    .O(n883),
    .I0(n882),
    .I1(n881)
  );
  //AND U79bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U79bar (
    .O(n883bar),
    .I0(n882bar),
    .I1(n881bar)
  );
  //OR U80
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U80 (
    .O(n881),
    .I0(in[118]),
    .I1(in[109])
  );
  //AND U80bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U80bar (
    .O(n881bar),
    .I0(inbar[118]),
    .I1(inbar[109])
  );
  //OR U81
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U81 (
    .O(n882),
    .I0(in[139]),
    .I1(in[120])
  );
  //AND U81bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U81bar (
    .O(n882bar),
    .I0(inbar[139]),
    .I1(inbar[120])
  );
  //OR U82
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U82 (
    .O(n884),
    .I0(n880),
    .I1(n879)
  );
  //AND U82bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U82bar (
    .O(n884bar),
    .I0(n880bar),
    .I1(n879bar)
  );
  //OR U83
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U83 (
    .O(n879),
    .I0(in[198]),
    .I1(in[154])
  );
  //AND U83bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U83bar (
    .O(n879bar),
    .I0(inbar[198]),
    .I1(inbar[154])
  );
  //OR U84
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U84 (
    .O(n880),
    .I0(in[210]),
    .I1(in[205])
  );
  //AND U84bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U84bar (
    .O(n880bar),
    .I0(inbar[210]),
    .I1(inbar[205])
  );
  //OR U85
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U85 (
    .O(n886),
    .I0(n878),
    .I1(n877)
  );
  //AND U85bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U85bar (
    .O(n886bar),
    .I0(n878bar),
    .I1(n877bar)
  );
  //OR U86
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U86 (
    .O(n877),
    .I0(n876),
    .I1(n875)
  );
  //AND U86bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U86bar (
    .O(n877bar),
    .I0(n876bar),
    .I1(n875bar)
  );
  //OR U87
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U87 (
    .O(n875),
    .I0(in[219]),
    .I1(in[217])
  );
  //AND U87bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U87bar (
    .O(n875bar),
    .I0(inbar[219]),
    .I1(inbar[217])
  );
  //OR U88
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U88 (
    .O(n876),
    .I0(in[86]),
    .I1(in[252])
  );
  //AND U88bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U88bar (
    .O(n876bar),
    .I0(inbar[86]),
    .I1(inbar[252])
  );
  //OR U89
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U89 (
    .O(n878),
    .I0(n874),
    .I1(n873)
  );
  //AND U89bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U89bar (
    .O(n878bar),
    .I0(n874bar),
    .I1(n873bar)
  );
  //OR U90
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U90 (
    .O(n873),
    .I0(in_40),
    .I1(in[91])
  );
  //AND U90bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U90bar (
    .O(n873bar),
    .I0(in_40bar),
    .I1(inbar[91])
  );
  //OR U91
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U91 (
    .O(n874),
    .I0(in_8),
    .I1(in_46)
  );
  //AND U91bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U91bar (
    .O(n874bar),
    .I0(in_8bar),
    .I1(in_46bar)
  );
  //OR U92
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U92 (
    .O(n889),
    .I0(n872),
    .I1(n871)
  );
  //AND U92bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U92bar (
    .O(n889bar),
    .I0(n872bar),
    .I1(n871bar)
  );
  //OR U93
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U93 (
    .O(n871),
    .I0(in[117]),
    .I1(n943)
  );
  //AND U93bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U93bar (
    .O(n871bar),
    .I0(inbar[117]),
    .I1(n943bar)
  );
  //OR U94
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U94 (
    .O(n943),
    .I0(n870),
    .I1(n869)
  );
  //AND U94bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U94bar (
    .O(n943bar),
    .I0(n870bar),
    .I1(n869bar)
  );
  //OR U95
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U95 (
    .O(n869),
    .I0(n868),
    .I1(n867)
  );
  //AND U95bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U95bar (
    .O(n869bar),
    .I0(n868bar),
    .I1(n867bar)
  );
  //OR U96
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U96 (
    .O(n867),
    .I0(n866),
    .I1(n865)
  );
  //AND U96bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U96bar (
    .O(n867bar),
    .I0(n866bar),
    .I1(n865bar)
  );
  //OR U97
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U97 (
    .O(n865),
    .I0(n864),
    .I1(n863)
  );
  //AND U97bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U97bar (
    .O(n865bar),
    .I0(n864bar),
    .I1(n863bar)
  );
  //OR U98
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U98 (
    .O(n866),
    .I0(in[108]),
    .I1(n919)
  );
  //AND U98bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U98bar (
    .O(n866bar),
    .I0(inbar[108]),
    .I1(n919bar)
  );
  //OR U99
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U99 (
    .O(n919),
    .I0(n862),
    .I1(n861)
  );
  //AND U99bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U99bar (
    .O(n919bar),
    .I0(n862bar),
    .I1(n861bar)
  );
  //OR U100
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U100 (
    .O(n861),
    .I0(n860),
    .I1(n859)
  );
  //AND U100bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U100bar (
    .O(n861bar),
    .I0(n860bar),
    .I1(n859bar)
  );
  //OR U101
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U101 (
    .O(n859),
    .I0(n858),
    .I1(n857)
  );
  //AND U101bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U101bar (
    .O(n859bar),
    .I0(n858bar),
    .I1(n857bar)
  );
  //OR U102
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U102 (
    .O(n857),
    .I0(in[119]),
    .I1(in[105])
  );
  //AND U102bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U102bar (
    .O(n857bar),
    .I0(inbar[119]),
    .I1(inbar[105])
  );
  //OR U103
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U103 (
    .O(n858),
    .I0(in[186]),
    .I1(in[175])
  );
  //AND U103bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U103bar (
    .O(n858bar),
    .I0(inbar[186]),
    .I1(inbar[175])
  );
  //OR U104
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U104 (
    .O(n860),
    .I0(n856),
    .I1(n855)
  );
  //AND U104bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U104bar (
    .O(n860bar),
    .I0(n856bar),
    .I1(n855bar)
  );
  //OR U105
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U105 (
    .O(n855),
    .I0(in[202]),
    .I1(in[193])
  );
  //AND U105bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U105bar (
    .O(n855bar),
    .I0(inbar[202]),
    .I1(inbar[193])
  );
  //OR U106
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U106 (
    .O(n856),
    .I0(in[225]),
    .I1(in[208])
  );
  //AND U106bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U106bar (
    .O(n856bar),
    .I0(inbar[225]),
    .I1(inbar[208])
  );
  //OR U107
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U107 (
    .O(n862),
    .I0(n854),
    .I1(n853)
  );
  //AND U107bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U107bar (
    .O(n862bar),
    .I0(n854bar),
    .I1(n853bar)
  );
  //OR U108
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U108 (
    .O(n853),
    .I0(n852),
    .I1(n851)
  );
  //AND U108bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U108bar (
    .O(n853bar),
    .I0(n852bar),
    .I1(n851bar)
  );
  //OR U109
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U109 (
    .O(n851),
    .I0(in_1),
    .I1(in[85])
  );
  //AND U109bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U109bar (
    .O(n851bar),
    .I0(in_1bar),
    .I1(inbar[85])
  );
  //OR U110
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U110 (
    .O(n852),
    .I0(in_23),
    .I1(in_19)
  );
  //AND U110bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U110bar (
    .O(n852bar),
    .I0(in_23bar),
    .I1(in_19bar)
  );
  //OR U111
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U111 (
    .O(n854),
    .I0(n850),
    .I1(n849)
  );
  //AND U111bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U111bar (
    .O(n854bar),
    .I0(n850bar),
    .I1(n849bar)
  );
  //OR U112
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U112 (
    .O(n849),
    .I0(in_43),
    .I1(in_33)
  );
  //AND U112bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U112bar (
    .O(n849bar),
    .I0(in_43bar),
    .I1(in_33bar)
  );
  //OR U113
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U113 (
    .O(n850),
    .I0(in_63),
    .I1(in_44)
  );
  //AND U113bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U113bar (
    .O(n850bar),
    .I0(in_63bar),
    .I1(in_44bar)
  );
  //OR U114
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U114 (
    .O(n868),
    .I0(n848),
    .I1(n847)
  );
  //AND U114bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U114bar (
    .O(n868bar),
    .I0(n848bar),
    .I1(n847bar)
  );
  //OR U115
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U115 (
    .O(n847),
    .I0(in[141]),
    .I1(in[112])
  );
  //AND U115bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U115bar (
    .O(n847bar),
    .I0(inbar[141]),
    .I1(inbar[112])
  );
  //OR U116
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U116 (
    .O(n848),
    .I0(in[147]),
    .I1(n846)
  );
  //AND U116bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U116bar (
    .O(n848bar),
    .I0(inbar[147]),
    .I1(n846bar)
  );
  //OR U117
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U117 (
    .O(n846),
    .I0(in[181]),
    .I1(in[167])
  );
  //AND U117bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U117bar (
    .O(n846bar),
    .I0(inbar[181]),
    .I1(inbar[167])
  );
  //OR U118
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U118 (
    .O(n870),
    .I0(n845),
    .I1(n844)
  );
  //AND U118bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U118bar (
    .O(n870bar),
    .I0(n845bar),
    .I1(n844bar)
  );
  //OR U119
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U119 (
    .O(n844),
    .I0(n843),
    .I1(n842)
  );
  //AND U119bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U119bar (
    .O(n844bar),
    .I0(n843bar),
    .I1(n842bar)
  );
  //OR U120
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U120 (
    .O(n842),
    .I0(in[229]),
    .I1(in[201])
  );
  //AND U120bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U120bar (
    .O(n842bar),
    .I0(inbar[229]),
    .I1(inbar[201])
  );
  //OR U121
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U121 (
    .O(n843),
    .I0(in[237]),
    .I1(n841)
  );
  //AND U121bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U121bar (
    .O(n843bar),
    .I0(inbar[237]),
    .I1(n841bar)
  );
  //OR U122
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U122 (
    .O(n841),
    .I0(in[94]),
    .I1(in[253])
  );
  //AND U122bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U122bar (
    .O(n841bar),
    .I0(inbar[94]),
    .I1(inbar[253])
  );
  //OR U123
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U123 (
    .O(n845),
    .I0(n840),
    .I1(n839)
  );
  //AND U123bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U123bar (
    .O(n845bar),
    .I0(n840bar),
    .I1(n839bar)
  );
  //OR U124
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U124 (
    .O(n839),
    .I0(in_21),
    .I1(in[96])
  );
  //AND U124bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U124bar (
    .O(n839bar),
    .I0(in_21bar),
    .I1(inbar[96])
  );
  //OR U125
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U125 (
    .O(n840),
    .I0(in_25),
    .I1(n838)
  );
  //AND U125bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U125bar (
    .O(n840bar),
    .I0(in_25bar),
    .I1(n838bar)
  );
  //OR U126
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U126 (
    .O(n838),
    .I0(in_81),
    .I1(in_45)
  );
  //AND U126bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U126bar (
    .O(n838bar),
    .I0(in_81bar),
    .I1(in_45bar)
  );
  //OR U127
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U127 (
    .O(n891),
    .I0(n837),
    .I1(n836)
  );
  //AND U127bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U127bar (
    .O(n891bar),
    .I0(n837bar),
    .I1(n836bar)
  );
  //OR U128
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U128 (
    .O(n836),
    .I0(in[142]),
    .I1(in[124])
  );
  //AND U128bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U128bar (
    .O(n836bar),
    .I0(inbar[142]),
    .I1(inbar[124])
  );
  //OR U129
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U129 (
    .O(n837),
    .I0(in[150]),
    .I1(n835)
  );
  //AND U129bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U129bar (
    .O(n837bar),
    .I0(inbar[150]),
    .I1(n835bar)
  );
  //OR U130
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U130 (
    .O(n835),
    .I0(in[172]),
    .I1(in[155])
  );
  //AND U130bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U130bar (
    .O(n835bar),
    .I0(inbar[172]),
    .I1(inbar[155])
  );
  //OR U131
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U131 (
    .O(n893),
    .I0(n834),
    .I1(n833)
  );
  //AND U131bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U131bar (
    .O(n893bar),
    .I0(n834bar),
    .I1(n833bar)
  );
  //OR U132
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U132 (
    .O(n833),
    .I0(n832),
    .I1(n831)
  );
  //AND U132bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U132bar (
    .O(n833bar),
    .I0(n832bar),
    .I1(n831bar)
  );
  //OR U133
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U133 (
    .O(n831),
    .I0(in[196]),
    .I1(in[173])
  );
  //AND U133bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U133bar (
    .O(n831bar),
    .I0(inbar[196]),
    .I1(inbar[173])
  );
  //OR U134
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U134 (
    .O(n832),
    .I0(in[222]),
    .I1(n830)
  );
  //AND U134bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U134bar (
    .O(n832bar),
    .I0(inbar[222]),
    .I1(n830bar)
  );
  //OR U135
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U135 (
    .O(n830),
    .I0(in[227]),
    .I1(in[226])
  );
  //AND U135bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U135bar (
    .O(n830bar),
    .I0(inbar[227]),
    .I1(inbar[226])
  );
  //OR U136
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U136 (
    .O(n834),
    .I0(n829),
    .I1(n828)
  );
  //AND U136bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U136bar (
    .O(n834bar),
    .I0(n829bar),
    .I1(n828bar)
  );
  //OR U137
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U137 (
    .O(n828),
    .I0(in[249]),
    .I1(in[231])
  );
  //AND U137bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U137bar (
    .O(n828bar),
    .I0(inbar[249]),
    .I1(inbar[231])
  );
  //OR U138
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U138 (
    .O(n829),
    .I0(in_28),
    .I1(n827)
  );
  //AND U138bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U138bar (
    .O(n829bar),
    .I0(in_28bar),
    .I1(n827bar)
  );
  //OR U139
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U139 (
    .O(n827),
    .I0(in_52),
    .I1(in_47)
  );
  //AND U139bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U139bar (
    .O(n827bar),
    .I0(in_52bar),
    .I1(in_47bar)
  );
  //OR U140
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U140 (
    .O(out[3]),
    .I0(n826),
    .I1(n825)
  );
  //AND U140bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U140bar (
    .O(outbar[3]),
    .I0(n826bar),
    .I1(n825bar)
  );
  //OR U141
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U141 (
    .O(n825),
    .I0(n824),
    .I1(n823)
  );
  //AND U141bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U141bar (
    .O(n825bar),
    .I0(n824bar),
    .I1(n823bar)
  );
  //OR U142
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U142 (
    .O(n823),
    .I0(n822),
    .I1(n821)
  );
  //AND U142bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U142bar (
    .O(n823bar),
    .I0(n822bar),
    .I1(n821bar)
  );
  //OR U143
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U143 (
    .O(n821),
    .I0(n820),
    .I1(n819)
  );
  //AND U143bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U143bar (
    .O(n821bar),
    .I0(n820bar),
    .I1(n819bar)
  );
  //OR U144
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U144 (
    .O(n822),
    .I0(n964),
    .I1(n818)
  );
  //AND U144bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U144bar (
    .O(n822bar),
    .I0(n964bar),
    .I1(n818bar)
  );
  //OR U145
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U145 (
    .O(n818),
    .I0(in[118]),
    .I1(n817)
  );
  //AND U145bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U145bar (
    .O(n818bar),
    .I0(inbar[118]),
    .I1(n817bar)
  );
  //OR U146
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U146 (
    .O(n964),
    .I0(n816),
    .I1(n815)
  );
  //AND U146bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U146bar (
    .O(n964bar),
    .I0(n816bar),
    .I1(n815bar)
  );
  //OR U147
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U147 (
    .O(n815),
    .I0(n814),
    .I1(n813)
  );
  //AND U147bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U147bar (
    .O(n815bar),
    .I0(n814bar),
    .I1(n813bar)
  );
  //OR U148
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U148 (
    .O(n813),
    .I0(n812),
    .I1(n811)
  );
  //AND U148bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U148bar (
    .O(n813bar),
    .I0(n812bar),
    .I1(n811bar)
  );
  //OR U149
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U149 (
    .O(n811),
    .I0(in[122]),
    .I1(in[111])
  );
  //AND U149bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U149bar (
    .O(n811bar),
    .I0(inbar[122]),
    .I1(inbar[111])
  );
  //OR U150
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U150 (
    .O(n812),
    .I0(in[154]),
    .I1(in[151])
  );
  //AND U150bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U150bar (
    .O(n812bar),
    .I0(inbar[154]),
    .I1(inbar[151])
  );
  //OR U151
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U151 (
    .O(n814),
    .I0(n810),
    .I1(n809)
  );
  //AND U151bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U151bar (
    .O(n814bar),
    .I0(n810bar),
    .I1(n809bar)
  );
  //OR U152
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U152 (
    .O(n809),
    .I0(in[187]),
    .I1(in[177])
  );
  //AND U152bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U152bar (
    .O(n809bar),
    .I0(inbar[187]),
    .I1(inbar[177])
  );
  //OR U153
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U153 (
    .O(n810),
    .I0(in[200]),
    .I1(in[192])
  );
  //AND U153bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U153bar (
    .O(n810bar),
    .I0(inbar[200]),
    .I1(inbar[192])
  );
  //OR U154
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U154 (
    .O(n816),
    .I0(n808),
    .I1(n807)
  );
  //AND U154bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U154bar (
    .O(n816bar),
    .I0(n808bar),
    .I1(n807bar)
  );
  //OR U155
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U155 (
    .O(n807),
    .I0(n806),
    .I1(n805)
  );
  //AND U155bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U155bar (
    .O(n807bar),
    .I0(n806bar),
    .I1(n805bar)
  );
  //OR U156
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U156 (
    .O(n805),
    .I0(in[225]),
    .I1(in[207])
  );
  //AND U156bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U156bar (
    .O(n805bar),
    .I0(inbar[225]),
    .I1(inbar[207])
  );
  //OR U157
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U157 (
    .O(n806),
    .I0(in[98]),
    .I1(in[226])
  );
  //AND U157bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U157bar (
    .O(n806bar),
    .I0(inbar[98]),
    .I1(inbar[226])
  );
  //OR U158
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U158 (
    .O(n808),
    .I0(n804),
    .I1(n803)
  );
  //AND U158bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U158bar (
    .O(n808bar),
    .I0(n804bar),
    .I1(n803bar)
  );
  //OR U159
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U159 (
    .O(n803),
    .I0(in_20),
    .I1(in_16)
  );
  //AND U159bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U159bar (
    .O(n803bar),
    .I0(in_20bar),
    .I1(in_16bar)
  );
  //OR U160
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U160 (
    .O(n804),
    .I0(in_55),
    .I1(in_45)
  );
  //AND U160bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U160bar (
    .O(n804bar),
    .I0(in_55bar),
    .I1(in_45bar)
  );
  //OR U161
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U161 (
    .O(n824),
    .I0(n802),
    .I1(n801)
  );
  //AND U161bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U161bar (
    .O(n824bar),
    .I0(n802bar),
    .I1(n801bar)
  );
  //OR U162
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U162 (
    .O(n801),
    .I0(in[162]),
    .I1(in[149])
  );
  //AND U162bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U162bar (
    .O(n801bar),
    .I0(inbar[162]),
    .I1(inbar[149])
  );
  //OR U163
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U163 (
    .O(n802),
    .I0(in[163]),
    .I1(n800)
  );
  //AND U163bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U163bar (
    .O(n802bar),
    .I0(inbar[163]),
    .I1(n800bar)
  );
  //OR U164
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U164 (
    .O(n800),
    .I0(in[191]),
    .I1(in[189])
  );
  //AND U164bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U164bar (
    .O(n800bar),
    .I0(inbar[191]),
    .I1(inbar[189])
  );
  //OR U165
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U165 (
    .O(n826),
    .I0(n799),
    .I1(n798)
  );
  //AND U165bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U165bar (
    .O(n826bar),
    .I0(n799bar),
    .I1(n798bar)
  );
  //OR U166
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U166 (
    .O(n798),
    .I0(n797),
    .I1(n796)
  );
  //AND U166bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U166bar (
    .O(n798bar),
    .I0(n797bar),
    .I1(n796bar)
  );
  //OR U167
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U167 (
    .O(n796),
    .I0(in[212]),
    .I1(in[193])
  );
  //AND U167bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U167bar (
    .O(n796bar),
    .I0(inbar[212]),
    .I1(inbar[193])
  );
  //OR U168
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U168 (
    .O(n797),
    .I0(in[238]),
    .I1(n795)
  );
  //AND U168bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U168bar (
    .O(n797bar),
    .I0(inbar[238]),
    .I1(n795bar)
  );
  //OR U169
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U169 (
    .O(n795),
    .I0(in[88]),
    .I1(in[247])
  );
  //AND U169bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U169bar (
    .O(n795bar),
    .I0(inbar[88]),
    .I1(inbar[247])
  );
  //OR U170
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U170 (
    .O(n799),
    .I0(n794),
    .I1(n793)
  );
  //AND U170bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U170bar (
    .O(n799bar),
    .I0(n794bar),
    .I1(n793bar)
  );
  //OR U171
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U171 (
    .O(n793),
    .I0(in[94]),
    .I1(in[92])
  );
  //AND U171bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U171bar (
    .O(n793bar),
    .I0(inbar[94]),
    .I1(inbar[92])
  );
  //OR U172
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U172 (
    .O(n794),
    .I0(in_52),
    .I1(n792)
  );
  //AND U172bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U172bar (
    .O(n794bar),
    .I0(in_52bar),
    .I1(n792bar)
  );
  //OR U173
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U173 (
    .O(n792),
    .I0(in_70),
    .I1(in_67)
  );
  //AND U173bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U173bar (
    .O(n792bar),
    .I0(in_70bar),
    .I1(in_67bar)
  );
  //OR U174
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U174 (
    .O(out[2]),
    .I0(n791),
    .I1(n790)
  );
  //AND U174bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U174bar (
    .O(outbar[2]),
    .I0(n791bar),
    .I1(n790bar)
  );
  //OR U175
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U175 (
    .O(n790),
    .I0(n789),
    .I1(n788)
  );
  //AND U175bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U175bar (
    .O(n790bar),
    .I0(n789bar),
    .I1(n788bar)
  );
  //OR U176
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U176 (
    .O(n788),
    .I0(n787),
    .I1(n786)
  );
  //AND U176bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U176bar (
    .O(n788bar),
    .I0(n787bar),
    .I1(n786bar)
  );
  //OR U177
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U177 (
    .O(n786),
    .I0(n819),
    .I1(n785)
  );
  //AND U177bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U177bar (
    .O(n786bar),
    .I0(n819bar),
    .I1(n785bar)
  );
  //OR U178
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U178 (
    .O(n819),
    .I0(n784),
    .I1(n783)
  );
  //AND U178bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U178bar (
    .O(n819bar),
    .I0(n784bar),
    .I1(n783bar)
  );
  //OR U179
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U179 (
    .O(n783),
    .I0(n782),
    .I1(n781)
  );
  //AND U179bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U179bar (
    .O(n783bar),
    .I0(n782bar),
    .I1(n781bar)
  );
  //OR U180
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U180 (
    .O(n781),
    .I0(n780),
    .I1(n779)
  );
  //AND U180bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U180bar (
    .O(n781bar),
    .I0(n780bar),
    .I1(n779bar)
  );
  //OR U181
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U181 (
    .O(n779),
    .I0(n962),
    .I1(n778)
  );
  //AND U181bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U181bar (
    .O(n779bar),
    .I0(n962bar),
    .I1(n778bar)
  );
  //OR U182
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U182 (
    .O(n962),
    .I0(n777),
    .I1(n776)
  );
  //AND U182bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U182bar (
    .O(n962bar),
    .I0(n777bar),
    .I1(n776bar)
  );
  //OR U183
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U183 (
    .O(n776),
    .I0(n775),
    .I1(n774)
  );
  //AND U183bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U183bar (
    .O(n776bar),
    .I0(n775bar),
    .I1(n774bar)
  );
  //OR U184
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U184 (
    .O(n774),
    .I0(n773),
    .I1(n772)
  );
  //AND U184bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U184bar (
    .O(n774bar),
    .I0(n773bar),
    .I1(n772bar)
  );
  //OR U185
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U185 (
    .O(n772),
    .I0(in[131]),
    .I1(in[120])
  );
  //AND U185bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U185bar (
    .O(n772bar),
    .I0(inbar[131]),
    .I1(inbar[120])
  );
  //OR U186
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U186 (
    .O(n773),
    .I0(in[153]),
    .I1(in[147])
  );
  //AND U186bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U186bar (
    .O(n773bar),
    .I0(inbar[153]),
    .I1(inbar[147])
  );
  //OR U187
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U187 (
    .O(n775),
    .I0(n771),
    .I1(n770)
  );
  //AND U187bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U187bar (
    .O(n775bar),
    .I0(n771bar),
    .I1(n770bar)
  );
  //OR U188
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U188 (
    .O(n770),
    .I0(in[170]),
    .I1(in[156])
  );
  //AND U188bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U188bar (
    .O(n770bar),
    .I0(inbar[170]),
    .I1(inbar[156])
  );
  //OR U189
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U189 (
    .O(n771),
    .I0(in[223]),
    .I1(in[190])
  );
  //AND U189bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U189bar (
    .O(n771bar),
    .I0(inbar[223]),
    .I1(inbar[190])
  );
  //OR U190
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U190 (
    .O(n777),
    .I0(n769),
    .I1(n768)
  );
  //AND U190bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U190bar (
    .O(n777bar),
    .I0(n769bar),
    .I1(n768bar)
  );
  //OR U191
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U191 (
    .O(n768),
    .I0(n767),
    .I1(n766)
  );
  //AND U191bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U191bar (
    .O(n768bar),
    .I0(n767bar),
    .I1(n766bar)
  );
  //OR U192
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U192 (
    .O(n766),
    .I0(in[236]),
    .I1(in[230])
  );
  //AND U192bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U192bar (
    .O(n766bar),
    .I0(inbar[236]),
    .I1(inbar[230])
  );
  //OR U193
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U193 (
    .O(n767),
    .I0(in[85]),
    .I1(in[240])
  );
  //AND U193bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U193bar (
    .O(n767bar),
    .I0(inbar[85]),
    .I1(inbar[240])
  );
  //OR U194
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U194 (
    .O(n769),
    .I0(n765),
    .I1(n764)
  );
  //AND U194bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U194bar (
    .O(n769bar),
    .I0(n765bar),
    .I1(n764bar)
  );
  //OR U195
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U195 (
    .O(n764),
    .I0(in_12),
    .I1(in[90])
  );
  //AND U195bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U195bar (
    .O(n764bar),
    .I0(in_12bar),
    .I1(inbar[90])
  );
  //OR U196
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U196 (
    .O(n765),
    .I0(in_39),
    .I1(in_28)
  );
  //AND U196bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U196bar (
    .O(n765bar),
    .I0(in_39bar),
    .I1(in_28bar)
  );
  //OR U197
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U197 (
    .O(n780),
    .I0(in[109]),
    .I1(n763)
  );
  //AND U197bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U197bar (
    .O(n780bar),
    .I0(inbar[109]),
    .I1(n763bar)
  );
  //OR U198
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U198 (
    .O(n782),
    .I0(n762),
    .I1(n761)
  );
  //AND U198bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U198bar (
    .O(n782bar),
    .I0(n762bar),
    .I1(n761bar)
  );
  //OR U199
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U199 (
    .O(n761),
    .I0(in[138]),
    .I1(in[129])
  );
  //AND U199bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U199bar (
    .O(n761bar),
    .I0(inbar[138]),
    .I1(inbar[129])
  );
  //OR U200
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U200 (
    .O(n762),
    .I0(in[157]),
    .I1(n760)
  );
  //AND U200bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U200bar (
    .O(n762bar),
    .I0(inbar[157]),
    .I1(n760bar)
  );
  //OR U201
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U201 (
    .O(n760),
    .I0(in[182]),
    .I1(in[167])
  );
  //AND U201bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U201bar (
    .O(n760bar),
    .I0(inbar[182]),
    .I1(inbar[167])
  );
  //OR U202
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U202 (
    .O(n784),
    .I0(n759),
    .I1(n758)
  );
  //AND U202bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U202bar (
    .O(n784bar),
    .I0(n759bar),
    .I1(n758bar)
  );
  //OR U203
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U203 (
    .O(n758),
    .I0(n757),
    .I1(n756)
  );
  //AND U203bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U203bar (
    .O(n758bar),
    .I0(n757bar),
    .I1(n756bar)
  );
  //OR U204
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U204 (
    .O(n756),
    .I0(in[195]),
    .I1(in[184])
  );
  //AND U204bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U204bar (
    .O(n756bar),
    .I0(inbar[195]),
    .I1(inbar[184])
  );
  //OR U205
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U205 (
    .O(n757),
    .I0(in[196]),
    .I1(n755)
  );
  //AND U205bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U205bar (
    .O(n757bar),
    .I0(inbar[196]),
    .I1(n755bar)
  );
  //OR U206
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U206 (
    .O(n755),
    .I0(in[215]),
    .I1(in[209])
  );
  //AND U206bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U206bar (
    .O(n755bar),
    .I0(inbar[215]),
    .I1(inbar[209])
  );
  //OR U207
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U207 (
    .O(n759),
    .I0(n754),
    .I1(n753)
  );
  //AND U207bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U207bar (
    .O(n759bar),
    .I0(n754bar),
    .I1(n753bar)
  );
  //OR U208
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U208 (
    .O(n753),
    .I0(in[93]),
    .I1(in[233])
  );
  //AND U208bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U208bar (
    .O(n753bar),
    .I0(inbar[93]),
    .I1(inbar[233])
  );
  //OR U209
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U209 (
    .O(n754),
    .I0(in_1),
    .I1(n752)
  );
  //AND U209bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U209bar (
    .O(n754bar),
    .I0(in_1bar),
    .I1(n752bar)
  );
  //OR U210
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U210 (
    .O(n752),
    .I0(in_69),
    .I1(in_66)
  );
  //AND U210bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U210bar (
    .O(n752bar),
    .I0(in_69bar),
    .I1(in_66bar)
  );
  //OR U211
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U211 (
    .O(n787),
    .I0(n966),
    .I1(n751)
  );
  //AND U211bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U211bar (
    .O(n787bar),
    .I0(n966bar),
    .I1(n751bar)
  );
  //OR U212
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U212 (
    .O(n751),
    .I0(in[134]),
    .I1(n750)
  );
  //AND U212bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U212bar (
    .O(n751bar),
    .I0(inbar[134]),
    .I1(n750bar)
  );
  //OR U213
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U213 (
    .O(n966),
    .I0(n749),
    .I1(n748)
  );
  //AND U213bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U213bar (
    .O(n966bar),
    .I0(n749bar),
    .I1(n748bar)
  );
  //OR U214
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U214 (
    .O(n748),
    .I0(n747),
    .I1(n746)
  );
  //AND U214bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U214bar (
    .O(n748bar),
    .I0(n747bar),
    .I1(n746bar)
  );
  //OR U215
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U215 (
    .O(n746),
    .I0(n745),
    .I1(n744)
  );
  //AND U215bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U215bar (
    .O(n746bar),
    .I0(n745bar),
    .I1(n744bar)
  );
  //OR U216
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U216 (
    .O(n744),
    .I0(in[136]),
    .I1(in[121])
  );
  //AND U216bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U216bar (
    .O(n744bar),
    .I0(inbar[136]),
    .I1(inbar[121])
  );
  //OR U217
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U217 (
    .O(n745),
    .I0(in[186]),
    .I1(in[174])
  );
  //AND U217bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U217bar (
    .O(n745bar),
    .I0(inbar[186]),
    .I1(inbar[174])
  );
  //OR U218
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U218 (
    .O(n747),
    .I0(n743),
    .I1(n742)
  );
  //AND U218bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U218bar (
    .O(n747bar),
    .I0(n743bar),
    .I1(n742bar)
  );
  //OR U219
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U219 (
    .O(n742),
    .I0(in[198]),
    .I1(in[197])
  );
  //AND U219bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U219bar (
    .O(n742bar),
    .I0(inbar[198]),
    .I1(inbar[197])
  );
  //OR U220
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U220 (
    .O(n743),
    .I0(in[214]),
    .I1(in[199])
  );
  //AND U220bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U220bar (
    .O(n743bar),
    .I0(inbar[214]),
    .I1(inbar[199])
  );
  //OR U221
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U221 (
    .O(n749),
    .I0(n741),
    .I1(n740)
  );
  //AND U221bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U221bar (
    .O(n749bar),
    .I0(n741bar),
    .I1(n740bar)
  );
  //OR U222
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U222 (
    .O(n740),
    .I0(n739),
    .I1(n738)
  );
  //AND U222bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U222bar (
    .O(n740bar),
    .I0(n739bar),
    .I1(n738bar)
  );
  //OR U223
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U223 (
    .O(n738),
    .I0(in[231]),
    .I1(in[220])
  );
  //AND U223bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U223bar (
    .O(n738bar),
    .I0(inbar[231]),
    .I1(inbar[220])
  );
  //OR U224
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U224 (
    .O(n739),
    .I0(in_25),
    .I1(in[245])
  );
  //AND U224bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U224bar (
    .O(n739bar),
    .I0(in_25bar),
    .I1(inbar[245])
  );
  //OR U225
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U225 (
    .O(n741),
    .I0(n737),
    .I1(n736)
  );
  //AND U225bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U225bar (
    .O(n741bar),
    .I0(n737bar),
    .I1(n736bar)
  );
  //OR U226
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U226 (
    .O(n736),
    .I0(in_53),
    .I1(in_29)
  );
  //AND U226bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U226bar (
    .O(n736bar),
    .I0(in_53bar),
    .I1(in_29bar)
  );
  //OR U227
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U227 (
    .O(n737),
    .I0(in_79),
    .I1(in_74)
  );
  //AND U227bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U227bar (
    .O(n737bar),
    .I0(in_79bar),
    .I1(in_74bar)
  );
  //OR U228
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U228 (
    .O(n789),
    .I0(n735),
    .I1(n734)
  );
  //AND U228bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U228bar (
    .O(n789bar),
    .I0(n735bar),
    .I1(n734bar)
  );
  //OR U229
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U229 (
    .O(n734),
    .I0(in[152]),
    .I1(in[140])
  );
  //AND U229bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U229bar (
    .O(n734bar),
    .I0(inbar[152]),
    .I1(inbar[140])
  );
  //OR U230
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U230 (
    .O(n735),
    .I0(in[155]),
    .I1(n733)
  );
  //AND U230bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U230bar (
    .O(n735bar),
    .I0(inbar[155]),
    .I1(n733bar)
  );
  //OR U231
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U231 (
    .O(n733),
    .I0(in[166]),
    .I1(in[165])
  );
  //AND U231bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U231bar (
    .O(n733bar),
    .I0(inbar[166]),
    .I1(inbar[165])
  );
  //OR U232
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U232 (
    .O(n791),
    .I0(n732),
    .I1(n731)
  );
  //AND U232bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U232bar (
    .O(n791bar),
    .I0(n732bar),
    .I1(n731bar)
  );
  //OR U233
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U233 (
    .O(n731),
    .I0(n730),
    .I1(n729)
  );
  //AND U233bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U233bar (
    .O(n731bar),
    .I0(n730bar),
    .I1(n729bar)
  );
  //OR U234
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U234 (
    .O(n729),
    .I0(in[202]),
    .I1(in[185])
  );
  //AND U234bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U234bar (
    .O(n729bar),
    .I0(inbar[202]),
    .I1(inbar[185])
  );
  //OR U235
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U235 (
    .O(n730),
    .I0(in[211]),
    .I1(n728)
  );
  //AND U235bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U235bar (
    .O(n730bar),
    .I0(inbar[211]),
    .I1(n728bar)
  );
  //OR U236
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U236 (
    .O(n728),
    .I0(in[255]),
    .I1(in[253])
  );
  //AND U236bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U236bar (
    .O(n728bar),
    .I0(inbar[255]),
    .I1(inbar[253])
  );
  //OR U237
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U237 (
    .O(n732),
    .I0(n727),
    .I1(n726)
  );
  //AND U237bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U237bar (
    .O(n732bar),
    .I0(n727bar),
    .I1(n726bar)
  );
  //OR U238
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U238 (
    .O(n726),
    .I0(in_35),
    .I1(in_15)
  );
  //AND U238bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U238bar (
    .O(n726bar),
    .I0(in_35bar),
    .I1(in_15bar)
  );
  //OR U239
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U239 (
    .O(n727),
    .I0(in_36),
    .I1(n725)
  );
  //AND U239bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U239bar (
    .O(n727bar),
    .I0(in_36bar),
    .I1(n725bar)
  );
  //OR U240
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U240 (
    .O(n725),
    .I0(in_48),
    .I1(in_40)
  );
  //AND U240bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U240bar (
    .O(n725bar),
    .I0(in_48bar),
    .I1(in_40bar)
  );
  //OR U241
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U241 (
    .O(out[1]),
    .I0(n724),
    .I1(n723)
  );
  //AND U241bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U241bar (
    .O(outbar[1]),
    .I0(n724bar),
    .I1(n723bar)
  );
  //OR U242
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U242 (
    .O(n723),
    .I0(n722),
    .I1(n721)
  );
  //AND U242bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U242bar (
    .O(n723bar),
    .I0(n722bar),
    .I1(n721bar)
  );
  //OR U243
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U243 (
    .O(n721),
    .I0(n720),
    .I1(n719)
  );
  //AND U243bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U243bar (
    .O(n721bar),
    .I0(n720bar),
    .I1(n719bar)
  );
  //OR U244
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U244 (
    .O(n719),
    .I0(n921),
    .I1(n887)
  );
  //AND U244bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U244bar (
    .O(n719bar),
    .I0(n921bar),
    .I1(n887bar)
  );
  //OR U245
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U245 (
    .O(n887),
    .I0(n718),
    .I1(n717)
  );
  //AND U245bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U245bar (
    .O(n887bar),
    .I0(n718bar),
    .I1(n717bar)
  );
  //OR U246
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U246 (
    .O(n717),
    .I0(n716),
    .I1(n715)
  );
  //AND U246bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U246bar (
    .O(n717bar),
    .I0(n716bar),
    .I1(n715bar)
  );
  //OR U247
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U247 (
    .O(n715),
    .I0(n714),
    .I1(n713)
  );
  //AND U247bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U247bar (
    .O(n715bar),
    .I0(n714bar),
    .I1(n713bar)
  );
  //OR U248
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U248 (
    .O(n713),
    .I0(in[116]),
    .I1(in[110])
  );
  //AND U248bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U248bar (
    .O(n713bar),
    .I0(inbar[116]),
    .I1(inbar[110])
  );
  //OR U249
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U249 (
    .O(n714),
    .I0(in[133]),
    .I1(in[130])
  );
  //AND U249bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U249bar (
    .O(n714bar),
    .I0(inbar[133]),
    .I1(inbar[130])
  );
  //OR U250
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U250 (
    .O(n716),
    .I0(n712),
    .I1(n711)
  );
  //AND U250bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U250bar (
    .O(n716bar),
    .I0(n712bar),
    .I1(n711bar)
  );
  //OR U251
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U251 (
    .O(n711),
    .I0(in[203]),
    .I1(in[135])
  );
  //AND U251bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U251bar (
    .O(n711bar),
    .I0(inbar[203]),
    .I1(inbar[135])
  );
  //OR U252
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U252 (
    .O(n712),
    .I0(in[232]),
    .I1(in[223])
  );
  //AND U252bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U252bar (
    .O(n712bar),
    .I0(inbar[232]),
    .I1(inbar[223])
  );
  //OR U253
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U253 (
    .O(n718),
    .I0(n710),
    .I1(n709)
  );
  //AND U253bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U253bar (
    .O(n718bar),
    .I0(n710bar),
    .I1(n709bar)
  );
  //OR U254
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U254 (
    .O(n709),
    .I0(n708),
    .I1(n707)
  );
  //AND U254bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U254bar (
    .O(n709bar),
    .I0(n708bar),
    .I1(n707bar)
  );
  //OR U255
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U255 (
    .O(n707),
    .I0(in[255]),
    .I1(in[233])
  );
  //AND U255bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U255bar (
    .O(n707bar),
    .I0(inbar[255]),
    .I1(inbar[233])
  );
  //OR U256
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U256 (
    .O(n708),
    .I0(in_53),
    .I1(in_34)
  );
  //AND U256bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U256bar (
    .O(n708bar),
    .I0(in_53bar),
    .I1(in_34bar)
  );
  //OR U257
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U257 (
    .O(n710),
    .I0(n706),
    .I1(n705)
  );
  //AND U257bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U257bar (
    .O(n710bar),
    .I0(n706bar),
    .I1(n705bar)
  );
  //OR U258
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U258 (
    .O(n705),
    .I0(in_57),
    .I1(in_55)
  );
  //AND U258bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U258bar (
    .O(n705bar),
    .I0(in_57bar),
    .I1(in_55bar)
  );
  //OR U259
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U259 (
    .O(n706),
    .I0(in_68),
    .I1(in_67)
  );
  //AND U259bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U259bar (
    .O(n706bar),
    .I0(in_68bar),
    .I1(in_67bar)
  );
  //OR U260
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U260 (
    .O(n921),
    .I0(n704),
    .I1(n703)
  );
  //AND U260bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U260bar (
    .O(n921bar),
    .I0(n704bar),
    .I1(n703bar)
  );
  //OR U261
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U261 (
    .O(n703),
    .I0(n702),
    .I1(n701)
  );
  //AND U261bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U261bar (
    .O(n703bar),
    .I0(n702bar),
    .I1(n701bar)
  );
  //OR U262
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U262 (
    .O(n701),
    .I0(n700),
    .I1(n699)
  );
  //AND U262bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U262bar (
    .O(n701bar),
    .I0(n700bar),
    .I1(n699bar)
  );
  //OR U263
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U263 (
    .O(n699),
    .I0(n944),
    .I1(n872)
  );
  //AND U263bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U263bar (
    .O(n699bar),
    .I0(n944bar),
    .I1(n872bar)
  );
  //OR U264
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U264 (
    .O(n872),
    .I0(n698),
    .I1(n697)
  );
  //AND U264bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U264bar (
    .O(n872bar),
    .I0(n698bar),
    .I1(n697bar)
  );
  //OR U265
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U265 (
    .O(n697),
    .I0(n696),
    .I1(n695)
  );
  //AND U265bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U265bar (
    .O(n697bar),
    .I0(n696bar),
    .I1(n695bar)
  );
  //OR U266
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U266 (
    .O(n695),
    .I0(n694),
    .I1(n693)
  );
  //AND U266bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U266bar (
    .O(n695bar),
    .I0(n694bar),
    .I1(n693bar)
  );
  //OR U267
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U267 (
    .O(n693),
    .I0(in[121]),
    .I1(in[102])
  );
  //AND U267bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U267bar (
    .O(n693bar),
    .I0(inbar[121]),
    .I1(inbar[102])
  );
  //OR U268
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U268 (
    .O(n694),
    .I0(in[162]),
    .I1(in[161])
  );
  //AND U268bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U268bar (
    .O(n694bar),
    .I0(inbar[162]),
    .I1(inbar[161])
  );
  //OR U269
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U269 (
    .O(n696),
    .I0(n692),
    .I1(n691)
  );
  //AND U269bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U269bar (
    .O(n696bar),
    .I0(n692bar),
    .I1(n691bar)
  );
  //OR U270
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U270 (
    .O(n691),
    .I0(in[192]),
    .I1(in[178])
  );
  //AND U270bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U270bar (
    .O(n691bar),
    .I0(inbar[192]),
    .I1(inbar[178])
  );
  //OR U271
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U271 (
    .O(n692),
    .I0(in[244]),
    .I1(in[209])
  );
  //AND U271bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U271bar (
    .O(n692bar),
    .I0(inbar[244]),
    .I1(inbar[209])
  );
  //OR U272
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U272 (
    .O(n698),
    .I0(n690),
    .I1(n689)
  );
  //AND U272bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U272bar (
    .O(n698bar),
    .I0(n690bar),
    .I1(n689bar)
  );
  //OR U273
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U273 (
    .O(n689),
    .I0(n688),
    .I1(n687)
  );
  //AND U273bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U273bar (
    .O(n689bar),
    .I0(n688bar),
    .I1(n687bar)
  );
  //OR U274
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U274 (
    .O(n687),
    .I0(in[90]),
    .I1(in[254])
  );
  //AND U274bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U274bar (
    .O(n687bar),
    .I0(inbar[90]),
    .I1(inbar[254])
  );
  //OR U275
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U275 (
    .O(n688),
    .I0(in_36),
    .I1(in_32)
  );
  //AND U275bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U275bar (
    .O(n688bar),
    .I0(in_36bar),
    .I1(in_32bar)
  );
  //OR U276
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U276 (
    .O(n690),
    .I0(n686),
    .I1(n685)
  );
  //AND U276bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U276bar (
    .O(n690bar),
    .I0(n686bar),
    .I1(n685bar)
  );
  //OR U277
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U277 (
    .O(n685),
    .I0(in_62),
    .I1(in_37)
  );
  //AND U277bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U277bar (
    .O(n685bar),
    .I0(in_62bar),
    .I1(in_37bar)
  );
  //OR U278
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U278 (
    .O(n686),
    .I0(in_75),
    .I1(in_73)
  );
  //AND U278bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U278bar (
    .O(n686bar),
    .I0(in_75bar),
    .I1(in_73bar)
  );
  //OR U279
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U279 (
    .O(n944),
    .I0(n684),
    .I1(n683)
  );
  //AND U279bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U279bar (
    .O(n944bar),
    .I0(n684bar),
    .I1(n683bar)
  );
  //OR U280
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U280 (
    .O(n683),
    .I0(n682),
    .I1(n681)
  );
  //AND U280bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U280bar (
    .O(n683bar),
    .I0(n682bar),
    .I1(n681bar)
  );
  //OR U281
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U281 (
    .O(n681),
    .I0(n680),
    .I1(n679)
  );
  //AND U281bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U281bar (
    .O(n681bar),
    .I0(n680bar),
    .I1(n679bar)
  );
  //OR U282
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U282 (
    .O(n679),
    .I0(in[171]),
    .I1(in[153])
  );
  //AND U282bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U282bar (
    .O(n679bar),
    .I0(inbar[171]),
    .I1(inbar[153])
  );
  //OR U283
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U283 (
    .O(n680),
    .I0(in[187]),
    .I1(in[176])
  );
  //AND U283bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U283bar (
    .O(n680bar),
    .I0(inbar[187]),
    .I1(inbar[176])
  );
  //OR U284
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U284 (
    .O(n682),
    .I0(n678),
    .I1(n677)
  );
  //AND U284bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U284bar (
    .O(n682bar),
    .I0(n678bar),
    .I1(n677bar)
  );
  //OR U285
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U285 (
    .O(n677),
    .I0(in[245]),
    .I1(in[211])
  );
  //AND U285bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U285bar (
    .O(n677bar),
    .I0(inbar[245]),
    .I1(inbar[211])
  );
  //OR U286
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U286 (
    .O(n678),
    .I0(in[97]),
    .I1(in[88])
  );
  //AND U286bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U286bar (
    .O(n678bar),
    .I0(inbar[97]),
    .I1(inbar[88])
  );
  //OR U287
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U287 (
    .O(n684),
    .I0(n676),
    .I1(n675)
  );
  //AND U287bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U287bar (
    .O(n684bar),
    .I0(n676bar),
    .I1(n675bar)
  );
  //OR U288
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U288 (
    .O(n675),
    .I0(n674),
    .I1(n673)
  );
  //AND U288bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U288bar (
    .O(n675bar),
    .I0(n674bar),
    .I1(n673bar)
  );
  //OR U289
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U289 (
    .O(n673),
    .I0(in_10),
    .I1(in_0)
  );
  //AND U289bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U289bar (
    .O(n673bar),
    .I0(in_10bar),
    .I1(in_0bar)
  );
  //OR U290
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U290 (
    .O(n674),
    .I0(in_59),
    .I1(in_5)
  );
  //AND U290bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U290bar (
    .O(n674bar),
    .I0(in_59bar),
    .I1(in_5bar)
  );
  //OR U291
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U291 (
    .O(n676),
    .I0(n672),
    .I1(n671)
  );
  //AND U291bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U291bar (
    .O(n676bar),
    .I0(n672bar),
    .I1(n671bar)
  );
  //OR U292
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U292 (
    .O(n671),
    .I0(in_60),
    .I1(in_6)
  );
  //AND U292bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U292bar (
    .O(n671bar),
    .I0(in_60bar),
    .I1(in_6bar)
  );
  //OR U293
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U293 (
    .O(n672),
    .I0(in_77),
    .I1(in_69)
  );
  //AND U293bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U293bar (
    .O(n672bar),
    .I0(in_77bar),
    .I1(in_69bar)
  );
  //OR U294
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U294 (
    .O(n700),
    .I0(in[113]),
    .I1(n864)
  );
  //AND U294bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U294bar (
    .O(n700bar),
    .I0(inbar[113]),
    .I1(n864bar)
  );
  //OR U295
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U295 (
    .O(n864),
    .I0(n670),
    .I1(n669)
  );
  //AND U295bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U295bar (
    .O(n864bar),
    .I0(n670bar),
    .I1(n669bar)
  );
  //OR U296
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U296 (
    .O(n669),
    .I0(n668),
    .I1(n667)
  );
  //AND U296bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U296bar (
    .O(n669bar),
    .I0(n668bar),
    .I1(n667bar)
  );
  //OR U297
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U297 (
    .O(n667),
    .I0(n666),
    .I1(n665)
  );
  //AND U297bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U297bar (
    .O(n667bar),
    .I0(n666bar),
    .I1(n665bar)
  );
  //OR U298
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U298 (
    .O(n665),
    .I0(in[125]),
    .I1(in[107])
  );
  //AND U298bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U298bar (
    .O(n665bar),
    .I0(inbar[125]),
    .I1(inbar[107])
  );
  //OR U299
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U299 (
    .O(n666),
    .I0(in[138]),
    .I1(in[126])
  );
  //AND U299bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U299bar (
    .O(n666bar),
    .I0(inbar[138]),
    .I1(inbar[126])
  );
  //OR U300
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U300 (
    .O(n668),
    .I0(n664),
    .I1(n663)
  );
  //AND U300bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U300bar (
    .O(n668bar),
    .I0(n664bar),
    .I1(n663bar)
  );
  //OR U301
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U301 (
    .O(n663),
    .I0(in[189]),
    .I1(in[143])
  );
  //AND U301bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U301bar (
    .O(n663bar),
    .I0(inbar[189]),
    .I1(inbar[143])
  );
  //OR U302
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U302 (
    .O(n664),
    .I0(in[99]),
    .I1(in[214])
  );
  //AND U302bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U302bar (
    .O(n664bar),
    .I0(inbar[99]),
    .I1(inbar[214])
  );
  //OR U303
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U303 (
    .O(n670),
    .I0(n662),
    .I1(n661)
  );
  //AND U303bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U303bar (
    .O(n670bar),
    .I0(n662bar),
    .I1(n661bar)
  );
  //OR U304
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U304 (
    .O(n661),
    .I0(n660),
    .I1(n659)
  );
  //AND U304bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U304bar (
    .O(n661bar),
    .I0(n660bar),
    .I1(n659bar)
  );
  //OR U305
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U305 (
    .O(n659),
    .I0(in_15),
    .I1(in_12)
  );
  //AND U305bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U305bar (
    .O(n659bar),
    .I0(in_15bar),
    .I1(in_12bar)
  );
  //OR U306
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U306 (
    .O(n660),
    .I0(in_20),
    .I1(in_2)
  );
  //AND U306bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U306bar (
    .O(n660bar),
    .I0(in_20bar),
    .I1(in_2bar)
  );
  //OR U307
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U307 (
    .O(n662),
    .I0(n658),
    .I1(n657)
  );
  //AND U307bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U307bar (
    .O(n662bar),
    .I0(n658bar),
    .I1(n657bar)
  );
  //OR U308
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U308 (
    .O(n657),
    .I0(in_30),
    .I1(in_3)
  );
  //AND U308bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U308bar (
    .O(n657bar),
    .I0(in_30bar),
    .I1(in_3bar)
  );
  //OR U309
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U309 (
    .O(n658),
    .I0(in_4),
    .I1(in_38)
  );
  //AND U309bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U309bar (
    .O(n658bar),
    .I0(in_4bar),
    .I1(in_38bar)
  );
  //OR U310
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U310 (
    .O(n702),
    .I0(n656),
    .I1(n655)
  );
  //AND U310bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U310bar (
    .O(n702bar),
    .I0(n656bar),
    .I1(n655bar)
  );
  //OR U311
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U311 (
    .O(n655),
    .I0(in[148]),
    .I1(in[137])
  );
  //AND U311bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U311bar (
    .O(n655bar),
    .I0(inbar[148]),
    .I1(inbar[137])
  );
  //OR U312
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U312 (
    .O(n656),
    .I0(in[149]),
    .I1(n654)
  );
  //AND U312bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U312bar (
    .O(n656bar),
    .I0(inbar[149]),
    .I1(n654bar)
  );
  //OR U313
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U313 (
    .O(n654),
    .I0(in[195]),
    .I1(in[190])
  );
  //AND U313bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U313bar (
    .O(n654bar),
    .I0(inbar[195]),
    .I1(inbar[190])
  );
  //OR U314
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U314 (
    .O(n704),
    .I0(n653),
    .I1(n652)
  );
  //AND U314bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U314bar (
    .O(n704bar),
    .I0(n653bar),
    .I1(n652bar)
  );
  //OR U315
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U315 (
    .O(n652),
    .I0(n651),
    .I1(n650)
  );
  //AND U315bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U315bar (
    .O(n652bar),
    .I0(n651bar),
    .I1(n650bar)
  );
  //OR U316
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U316 (
    .O(n650),
    .I0(in[98]),
    .I1(in[197])
  );
  //AND U316bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U316bar (
    .O(n650bar),
    .I0(inbar[98]),
    .I1(inbar[197])
  );
  //OR U317
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U317 (
    .O(n651),
    .I0(in_11),
    .I1(n649)
  );
  //AND U317bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U317bar (
    .O(n651bar),
    .I0(in_11bar),
    .I1(n649bar)
  );
  //OR U318
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U318 (
    .O(n649),
    .I0(in_26),
    .I1(in_14)
  );
  //AND U318bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U318bar (
    .O(n649bar),
    .I0(in_26bar),
    .I1(in_14bar)
  );
  //OR U319
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U319 (
    .O(n653),
    .I0(n648),
    .I1(n647)
  );
  //AND U319bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U319bar (
    .O(n653bar),
    .I0(n648bar),
    .I1(n647bar)
  );
  //OR U320
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U320 (
    .O(n647),
    .I0(in_35),
    .I1(in_27)
  );
  //AND U320bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U320bar (
    .O(n647bar),
    .I0(in_35bar),
    .I1(in_27bar)
  );
  //OR U321
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U321 (
    .O(n648),
    .I0(in_50),
    .I1(n646)
  );
  //AND U321bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U321bar (
    .O(n648bar),
    .I0(in_50bar),
    .I1(n646bar)
  );
  //OR U322
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U322 (
    .O(n646),
    .I0(in_78),
    .I1(in_61)
  );
  //AND U322bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U322bar (
    .O(n646bar),
    .I0(in_78bar),
    .I1(in_61bar)
  );
  //OR U323
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U323 (
    .O(n720),
    .I0(n942),
    .I1(n645)
  );
  //AND U323bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U323bar (
    .O(n720bar),
    .I0(n942bar),
    .I1(n645bar)
  );
  //OR U324
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U324 (
    .O(n645),
    .I0(in[106]),
    .I1(n863)
  );
  //AND U324bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U324bar (
    .O(n645bar),
    .I0(inbar[106]),
    .I1(n863bar)
  );
  //OR U325
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U325 (
    .O(n863),
    .I0(n644),
    .I1(n643)
  );
  //AND U325bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U325bar (
    .O(n863bar),
    .I0(n644bar),
    .I1(n643bar)
  );
  //OR U326
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U326 (
    .O(n643),
    .I0(n642),
    .I1(n641)
  );
  //AND U326bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U326bar (
    .O(n643bar),
    .I0(n642bar),
    .I1(n641bar)
  );
  //OR U327
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U327 (
    .O(n641),
    .I0(n640),
    .I1(n639)
  );
  //AND U327bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U327bar (
    .O(n641bar),
    .I0(n640bar),
    .I1(n639bar)
  );
  //OR U328
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U328 (
    .O(n639),
    .I0(in[127]),
    .I1(in[122])
  );
  //AND U328bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U328bar (
    .O(n639bar),
    .I0(inbar[127]),
    .I1(inbar[122])
  );
  //OR U329
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U329 (
    .O(n640),
    .I0(in[156]),
    .I1(in[132])
  );
  //AND U329bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U329bar (
    .O(n640bar),
    .I0(inbar[156]),
    .I1(inbar[132])
  );
  //OR U330
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U330 (
    .O(n642),
    .I0(n638),
    .I1(n637)
  );
  //AND U330bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U330bar (
    .O(n642bar),
    .I0(n638bar),
    .I1(n637bar)
  );
  //OR U331
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U331 (
    .O(n637),
    .I0(in[159]),
    .I1(in[157])
  );
  //AND U331bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U331bar (
    .O(n637bar),
    .I0(inbar[159]),
    .I1(inbar[157])
  );
  //OR U332
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U332 (
    .O(n638),
    .I0(in[185]),
    .I1(in[169])
  );
  //AND U332bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U332bar (
    .O(n638bar),
    .I0(inbar[185]),
    .I1(inbar[169])
  );
  //OR U333
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U333 (
    .O(n644),
    .I0(n636),
    .I1(n635)
  );
  //AND U333bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U333bar (
    .O(n644bar),
    .I0(n636bar),
    .I1(n635bar)
  );
  //OR U334
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U334 (
    .O(n635),
    .I0(n634),
    .I1(n633)
  );
  //AND U334bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U334bar (
    .O(n635bar),
    .I0(n634bar),
    .I1(n633bar)
  );
  //OR U335
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U335 (
    .O(n633),
    .I0(in[239]),
    .I1(in[218])
  );
  //AND U335bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U335bar (
    .O(n633bar),
    .I0(inbar[239]),
    .I1(inbar[218])
  );
  //OR U336
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U336 (
    .O(n634),
    .I0(in_13),
    .I1(in[87])
  );
  //AND U336bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U336bar (
    .O(n634bar),
    .I0(in_13bar),
    .I1(inbar[87])
  );
  //OR U337
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U337 (
    .O(n636),
    .I0(n632),
    .I1(n631)
  );
  //AND U337bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U337bar (
    .O(n636bar),
    .I0(n632bar),
    .I1(n631bar)
  );
  //OR U338
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U338 (
    .O(n631),
    .I0(in_72),
    .I1(in_70)
  );
  //AND U338bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U338bar (
    .O(n631bar),
    .I0(in_72bar),
    .I1(in_70bar)
  );
  //OR U339
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U339 (
    .O(n632),
    .I0(in_80),
    .I1(in_74)
  );
  //AND U339bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U339bar (
    .O(n632bar),
    .I0(in_80bar),
    .I1(in_74bar)
  );
  //OR U340
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U340 (
    .O(n942),
    .I0(n630),
    .I1(n629)
  );
  //AND U340bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U340bar (
    .O(n942bar),
    .I0(n630bar),
    .I1(n629bar)
  );
  //OR U341
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U341 (
    .O(n629),
    .I0(n628),
    .I1(n627)
  );
  //AND U341bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U341bar (
    .O(n629bar),
    .I0(n628bar),
    .I1(n627bar)
  );
  //OR U342
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U342 (
    .O(n627),
    .I0(n626),
    .I1(n625)
  );
  //AND U342bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U342bar (
    .O(n627bar),
    .I0(n626bar),
    .I1(n625bar)
  );
  //OR U343
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U343 (
    .O(n625),
    .I0(in[146]),
    .I1(in[100])
  );
  //AND U343bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U343bar (
    .O(n625bar),
    .I0(inbar[146]),
    .I1(inbar[100])
  );
  //OR U344
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U344 (
    .O(n626),
    .I0(in[168]),
    .I1(in[152])
  );
  //AND U344bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U344bar (
    .O(n626bar),
    .I0(inbar[168]),
    .I1(inbar[152])
  );
  //OR U345
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U345 (
    .O(n628),
    .I0(n624),
    .I1(n623)
  );
  //AND U345bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U345bar (
    .O(n628bar),
    .I0(n624bar),
    .I1(n623bar)
  );
  //OR U346
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U346 (
    .O(n623),
    .I0(in[199]),
    .I1(in[182])
  );
  //AND U346bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U346bar (
    .O(n623bar),
    .I0(inbar[199]),
    .I1(inbar[182])
  );
  //OR U347
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U347 (
    .O(n624),
    .I0(in[236]),
    .I1(in[204])
  );
  //AND U347bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U347bar (
    .O(n624bar),
    .I0(inbar[236]),
    .I1(inbar[204])
  );
  //OR U348
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U348 (
    .O(n630),
    .I0(n622),
    .I1(n621)
  );
  //AND U348bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U348bar (
    .O(n630bar),
    .I0(n622bar),
    .I1(n621bar)
  );
  //OR U349
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U349 (
    .O(n621),
    .I0(n620),
    .I1(n619)
  );
  //AND U349bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U349bar (
    .O(n621bar),
    .I0(n620bar),
    .I1(n619bar)
  );
  //OR U350
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U350 (
    .O(n619),
    .I0(in[89]),
    .I1(in[246])
  );
  //AND U350bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U350bar (
    .O(n619bar),
    .I0(inbar[89]),
    .I1(inbar[246])
  );
  //OR U351
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U351 (
    .O(n620),
    .I0(in[95]),
    .I1(in[92])
  );
  //AND U351bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U351bar (
    .O(n620bar),
    .I0(inbar[95]),
    .I1(inbar[92])
  );
  //OR U352
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U352 (
    .O(n622),
    .I0(n618),
    .I1(n617)
  );
  //AND U352bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U352bar (
    .O(n622bar),
    .I0(n618bar),
    .I1(n617bar)
  );
  //OR U353
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U353 (
    .O(n617),
    .I0(in_22),
    .I1(in_16)
  );
  //AND U353bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U353bar (
    .O(n617bar),
    .I0(in_22bar),
    .I1(in_16bar)
  );
  //OR U354
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U354 (
    .O(n618),
    .I0(in_51),
    .I1(in_49)
  );
  //AND U354bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U354bar (
    .O(n618bar),
    .I0(in_51bar),
    .I1(in_49bar)
  );
  //OR U355
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U355 (
    .O(n722),
    .I0(n616),
    .I1(n615)
  );
  //AND U355bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U355bar (
    .O(n722bar),
    .I0(n616bar),
    .I1(n615bar)
  );
  //OR U356
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U356 (
    .O(n615),
    .I0(in[158]),
    .I1(in[115])
  );
  //AND U356bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U356bar (
    .O(n615bar),
    .I0(inbar[158]),
    .I1(inbar[115])
  );
  //OR U357
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U357 (
    .O(n616),
    .I0(in[163]),
    .I1(n614)
  );
  //AND U357bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U357bar (
    .O(n616bar),
    .I0(inbar[163]),
    .I1(n614bar)
  );
  //OR U358
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U358 (
    .O(n614),
    .I0(in[206]),
    .I1(in[165])
  );
  //AND U358bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U358bar (
    .O(n614bar),
    .I0(inbar[206]),
    .I1(inbar[165])
  );
  //OR U359
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U359 (
    .O(n724),
    .I0(n613),
    .I1(n612)
  );
  //AND U359bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U359bar (
    .O(n724bar),
    .I0(n613bar),
    .I1(n612bar)
  );
  //OR U360
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U360 (
    .O(n612),
    .I0(n611),
    .I1(n610)
  );
  //AND U360bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U360bar (
    .O(n612bar),
    .I0(n611bar),
    .I1(n610bar)
  );
  //OR U361
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U361 (
    .O(n610),
    .I0(in[213]),
    .I1(in[207])
  );
  //AND U361bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U361bar (
    .O(n610bar),
    .I0(inbar[213]),
    .I1(inbar[207])
  );
  //OR U362
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U362 (
    .O(n611),
    .I0(in[215]),
    .I1(n609)
  );
  //AND U362bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U362bar (
    .O(n611bar),
    .I0(inbar[215]),
    .I1(n609bar)
  );
  //OR U363
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U363 (
    .O(n609),
    .I0(in[230]),
    .I1(in[220])
  );
  //AND U363bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U363bar (
    .O(n609bar),
    .I0(inbar[230]),
    .I1(inbar[220])
  );
  //OR U364
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U364 (
    .O(n613),
    .I0(n608),
    .I1(n607)
  );
  //AND U364bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U364bar (
    .O(n613bar),
    .I0(n608bar),
    .I1(n607bar)
  );
  //OR U365
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U365 (
    .O(n607),
    .I0(in[251]),
    .I1(in[234])
  );
  //AND U365bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U365bar (
    .O(n607bar),
    .I0(inbar[251]),
    .I1(inbar[234])
  );
  //OR U366
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U366 (
    .O(n608),
    .I0(in_17),
    .I1(n606)
  );
  //AND U366bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U366bar (
    .O(n608bar),
    .I0(in_17bar),
    .I1(n606bar)
  );
  //OR U367
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U367 (
    .O(n606),
    .I0(in_65),
    .I1(in_56)
  );
  //AND U367bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U367bar (
    .O(n606bar),
    .I0(in_65bar),
    .I1(in_56bar)
  );
  //OR U368
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U368 (
    .O(out[0]),
    .I0(n605),
    .I1(n604)
  );
  //AND U368bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U368bar (
    .O(outbar[0]),
    .I0(n605bar),
    .I1(n604bar)
  );
  //OR U369
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U369 (
    .O(n604),
    .I0(n603),
    .I1(n602)
  );
  //AND U369bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U369bar (
    .O(n604bar),
    .I0(n603bar),
    .I1(n602bar)
  );
  //OR U370
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U370 (
    .O(n602),
    .I0(n601),
    .I1(n600)
  );
  //AND U370bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U370bar (
    .O(n602bar),
    .I0(n601bar),
    .I1(n600bar)
  );
  //OR U371
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U371 (
    .O(n600),
    .I0(n820),
    .I1(n785)
  );
  //AND U371bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U371bar (
    .O(n600bar),
    .I0(n820bar),
    .I1(n785bar)
  );
  //OR U372
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U372 (
    .O(n785),
    .I0(n599),
    .I1(n598)
  );
  //AND U372bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U372bar (
    .O(n785bar),
    .I0(n599bar),
    .I1(n598bar)
  );
  //OR U373
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U373 (
    .O(n598),
    .I0(n597),
    .I1(n596)
  );
  //AND U373bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U373bar (
    .O(n598bar),
    .I0(n597bar),
    .I1(n596bar)
  );
  //OR U374
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U374 (
    .O(n596),
    .I0(n595),
    .I1(n594)
  );
  //AND U374bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U374bar (
    .O(n596bar),
    .I0(n595bar),
    .I1(n594bar)
  );
  //OR U375
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U375 (
    .O(n594),
    .I0(in[135]),
    .I1(in[104])
  );
  //AND U375bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U375bar (
    .O(n594bar),
    .I0(inbar[135]),
    .I1(inbar[104])
  );
  //OR U376
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U376 (
    .O(n595),
    .I0(in[188]),
    .I1(in[178])
  );
  //AND U376bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U376bar (
    .O(n595bar),
    .I0(inbar[188]),
    .I1(inbar[178])
  );
  //OR U377
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U377 (
    .O(n597),
    .I0(n593),
    .I1(n592)
  );
  //AND U377bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U377bar (
    .O(n597bar),
    .I0(n593bar),
    .I1(n592bar)
  );
  //OR U378
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U378 (
    .O(n592),
    .I0(in[217]),
    .I1(in[194])
  );
  //AND U378bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U378bar (
    .O(n592bar),
    .I0(inbar[217]),
    .I1(inbar[194])
  );
  //OR U379
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U379 (
    .O(n593),
    .I0(in[237]),
    .I1(in[218])
  );
  //AND U379bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U379bar (
    .O(n593bar),
    .I0(inbar[237]),
    .I1(inbar[218])
  );
  //OR U380
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U380 (
    .O(n599),
    .I0(n591),
    .I1(n590)
  );
  //AND U380bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U380bar (
    .O(n599bar),
    .I0(n591bar),
    .I1(n590bar)
  );
  //OR U381
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U381 (
    .O(n590),
    .I0(n589),
    .I1(n588)
  );
  //AND U381bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U381bar (
    .O(n590bar),
    .I0(n589bar),
    .I1(n588bar)
  );
  //OR U382
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U382 (
    .O(n588),
    .I0(in_2),
    .I1(in_10)
  );
  //AND U382bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U382bar (
    .O(n588bar),
    .I0(in_2bar),
    .I1(in_10bar)
  );
  //OR U383
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U383 (
    .O(n589),
    .I0(in_47),
    .I1(in_22)
  );
  //AND U383bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U383bar (
    .O(n589bar),
    .I0(in_47bar),
    .I1(in_22bar)
  );
  //OR U384
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U384 (
    .O(n591),
    .I0(n587),
    .I1(n586)
  );
  //AND U384bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U384bar (
    .O(n591bar),
    .I0(n587bar),
    .I1(n586bar)
  );
  //OR U385
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U385 (
    .O(n586),
    .I0(in_56),
    .I1(in_54)
  );
  //AND U385bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U385bar (
    .O(n586bar),
    .I0(in_56bar),
    .I1(in_54bar)
  );
  //OR U386
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U386 (
    .O(n587),
    .I0(in_63),
    .I1(in_61)
  );
  //AND U386bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U386bar (
    .O(n587bar),
    .I0(in_63bar),
    .I1(in_61bar)
  );
  //OR U387
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U387 (
    .O(n820),
    .I0(n585),
    .I1(n584)
  );
  //AND U387bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U387bar (
    .O(n820bar),
    .I0(n585bar),
    .I1(n584bar)
  );
  //OR U388
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U388 (
    .O(n584),
    .I0(n583),
    .I1(n582)
  );
  //AND U388bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U388bar (
    .O(n584bar),
    .I0(n583bar),
    .I1(n582bar)
  );
  //OR U389
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U389 (
    .O(n582),
    .I0(n581),
    .I1(n580)
  );
  //AND U389bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U389bar (
    .O(n582bar),
    .I0(n581bar),
    .I1(n580bar)
  );
  //OR U390
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U390 (
    .O(n580),
    .I0(in[158]),
    .I1(in[142])
  );
  //AND U390bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U390bar (
    .O(n580bar),
    .I0(inbar[158]),
    .I1(inbar[142])
  );
  //OR U391
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U391 (
    .O(n581),
    .I0(in[175]),
    .I1(in[164])
  );
  //AND U391bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U391bar (
    .O(n581bar),
    .I0(inbar[175]),
    .I1(inbar[164])
  );
  //OR U392
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U392 (
    .O(n583),
    .I0(n579),
    .I1(n578)
  );
  //AND U392bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U392bar (
    .O(n583bar),
    .I0(n579bar),
    .I1(n578bar)
  );
  //OR U393
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U393 (
    .O(n578),
    .I0(in[228]),
    .I1(in[204])
  );
  //AND U393bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U393bar (
    .O(n578bar),
    .I0(inbar[228]),
    .I1(inbar[204])
  );
  //OR U394
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U394 (
    .O(n579),
    .I0(in[91]),
    .I1(in[87])
  );
  //AND U394bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U394bar (
    .O(n579bar),
    .I0(inbar[91]),
    .I1(inbar[87])
  );
  //OR U395
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U395 (
    .O(n585),
    .I0(n577),
    .I1(n576)
  );
  //AND U395bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U395bar (
    .O(n585bar),
    .I0(n577bar),
    .I1(n576bar)
  );
  //OR U396
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U396 (
    .O(n576),
    .I0(n575),
    .I1(n574)
  );
  //AND U396bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U396bar (
    .O(n576bar),
    .I0(n575bar),
    .I1(n574bar)
  );
  //OR U397
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U397 (
    .O(n574),
    .I0(in_21),
    .I1(in_11)
  );
  //AND U397bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U397bar (
    .O(n574bar),
    .I0(in_21bar),
    .I1(in_11bar)
  );
  //OR U398
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U398 (
    .O(n575),
    .I0(in_5),
    .I1(in_3)
  );
  //AND U398bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U398bar (
    .O(n575bar),
    .I0(in_5bar),
    .I1(in_3bar)
  );
  //OR U399
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U399 (
    .O(n577),
    .I0(n573),
    .I1(n572)
  );
  //AND U399bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U399bar (
    .O(n577bar),
    .I0(n573bar),
    .I1(n572bar)
  );
  //OR U400
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U400 (
    .O(n572),
    .I0(in_68),
    .I1(in_64)
  );
  //AND U400bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U400bar (
    .O(n572bar),
    .I0(in_68bar),
    .I1(in_64bar)
  );
  //OR U401
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U401 (
    .O(n573),
    .I0(in_76),
    .I1(in_73)
  );
  //AND U401bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U401bar (
    .O(n573bar),
    .I0(in_76bar),
    .I1(in_73bar)
  );
  //OR U402
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U402 (
    .O(n601),
    .I0(n778),
    .I1(n571)
  );
  //AND U402bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U402bar (
    .O(n601bar),
    .I0(n778bar),
    .I1(n571bar)
  );
  //OR U403
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U403 (
    .O(n571),
    .I0(in[100]),
    .I1(n965)
  );
  //AND U403bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U403bar (
    .O(n571bar),
    .I0(inbar[100]),
    .I1(n965bar)
  );
  //OR U404
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U404 (
    .O(n965),
    .I0(n570),
    .I1(n569)
  );
  //AND U404bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U404bar (
    .O(n965bar),
    .I0(n570bar),
    .I1(n569bar)
  );
  //OR U405
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U405 (
    .O(n569),
    .I0(n568),
    .I1(n567)
  );
  //AND U405bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U405bar (
    .O(n569bar),
    .I0(n568bar),
    .I1(n567bar)
  );
  //OR U406
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U406 (
    .O(n567),
    .I0(n566),
    .I1(n565)
  );
  //AND U406bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U406bar (
    .O(n567bar),
    .I0(n566bar),
    .I1(n565bar)
  );
  //OR U407
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U407 (
    .O(n565),
    .I0(n817),
    .I1(n750)
  );
  //AND U407bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U407bar (
    .O(n565bar),
    .I0(n817bar),
    .I1(n750bar)
  );
  //OR U408
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U408 (
    .O(n750),
    .I0(n564),
    .I1(n563)
  );
  //AND U408bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U408bar (
    .O(n750bar),
    .I0(n564bar),
    .I1(n563bar)
  );
  //OR U409
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U409 (
    .O(n563),
    .I0(n562),
    .I1(n561)
  );
  //AND U409bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U409bar (
    .O(n563bar),
    .I0(n562bar),
    .I1(n561bar)
  );
  //OR U410
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U410 (
    .O(n561),
    .I0(n560),
    .I1(n559)
  );
  //AND U410bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U410bar (
    .O(n561bar),
    .I0(n560bar),
    .I1(n559bar)
  );
  //OR U411
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U411 (
    .O(n559),
    .I0(in[119]),
    .I1(in[103])
  );
  //AND U411bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U411bar (
    .O(n559bar),
    .I0(inbar[119]),
    .I1(inbar[103])
  );
  //OR U412
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U412 (
    .O(n560),
    .I0(in[137]),
    .I1(in[133])
  );
  //AND U412bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U412bar (
    .O(n560bar),
    .I0(inbar[137]),
    .I1(inbar[133])
  );
  //OR U413
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U413 (
    .O(n562),
    .I0(n558),
    .I1(n557)
  );
  //AND U413bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U413bar (
    .O(n562bar),
    .I0(n558bar),
    .I1(n557bar)
  );
  //OR U414
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U414 (
    .O(n557),
    .I0(in[176]),
    .I1(in[173])
  );
  //AND U414bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U414bar (
    .O(n557bar),
    .I0(inbar[176]),
    .I1(inbar[173])
  );
  //OR U415
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U415 (
    .O(n558),
    .I0(in[210]),
    .I1(in[181])
  );
  //AND U415bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U415bar (
    .O(n558bar),
    .I0(inbar[210]),
    .I1(inbar[181])
  );
  //OR U416
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U416 (
    .O(n564),
    .I0(n556),
    .I1(n555)
  );
  //AND U416bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U416bar (
    .O(n564bar),
    .I0(n556bar),
    .I1(n555bar)
  );
  //OR U417
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U417 (
    .O(n555),
    .I0(n554),
    .I1(n553)
  );
  //AND U417bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U417bar (
    .O(n555bar),
    .I0(n554bar),
    .I1(n553bar)
  );
  //OR U418
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U418 (
    .O(n553),
    .I0(in_13),
    .I1(in[234])
  );
  //AND U418bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U418bar (
    .O(n553bar),
    .I0(in_13bar),
    .I1(inbar[234])
  );
  //OR U419
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U419 (
    .O(n554),
    .I0(in_38),
    .I1(in_32)
  );
  //AND U419bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U419bar (
    .O(n554bar),
    .I0(in_38bar),
    .I1(in_32bar)
  );
  //OR U420
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U420 (
    .O(n556),
    .I0(n552),
    .I1(n551)
  );
  //AND U420bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U420bar (
    .O(n556bar),
    .I0(n552bar),
    .I1(n551bar)
  );
  //OR U421
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U421 (
    .O(n551),
    .I0(in_42),
    .I1(in_41)
  );
  //AND U421bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U421bar (
    .O(n551bar),
    .I0(in_42bar),
    .I1(in_41bar)
  );
  //OR U422
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U422 (
    .O(n552),
    .I0(in_7),
    .I1(in_49)
  );
  //AND U422bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U422bar (
    .O(n552bar),
    .I0(in_7bar),
    .I1(in_49bar)
  );
  //OR U423
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U423 (
    .O(n817),
    .I0(n550),
    .I1(n549)
  );
  //AND U423bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U423bar (
    .O(n817bar),
    .I0(n550bar),
    .I1(n549bar)
  );
  //OR U424
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U424 (
    .O(n549),
    .I0(n548),
    .I1(n547)
  );
  //AND U424bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U424bar (
    .O(n549bar),
    .I0(n548bar),
    .I1(n547bar)
  );
  //OR U425
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U425 (
    .O(n547),
    .I0(n546),
    .I1(n545)
  );
  //AND U425bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U425bar (
    .O(n547bar),
    .I0(n546bar),
    .I1(n545bar)
  );
  //OR U426
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U426 (
    .O(n545),
    .I0(in[159]),
    .I1(in[105])
  );
  //AND U426bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U426bar (
    .O(n545bar),
    .I0(inbar[159]),
    .I1(inbar[105])
  );
  //OR U427
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U427 (
    .O(n546),
    .I0(in[206]),
    .I1(in[183])
  );
  //AND U427bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U427bar (
    .O(n546bar),
    .I0(inbar[206]),
    .I1(inbar[183])
  );
  //OR U428
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U428 (
    .O(n548),
    .I0(n544),
    .I1(n543)
  );
  //AND U428bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U428bar (
    .O(n548bar),
    .I0(n544bar),
    .I1(n543bar)
  );
  //OR U429
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U429 (
    .O(n543),
    .I0(in[229]),
    .I1(in[219])
  );
  //AND U429bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U429bar (
    .O(n543bar),
    .I0(inbar[229]),
    .I1(inbar[219])
  );
  //OR U430
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U430 (
    .O(n544),
    .I0(in[235]),
    .I1(in[232])
  );
  //AND U430bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U430bar (
    .O(n544bar),
    .I0(inbar[235]),
    .I1(inbar[232])
  );
  //OR U431
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U431 (
    .O(n550),
    .I0(n542),
    .I1(n541)
  );
  //AND U431bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U431bar (
    .O(n550bar),
    .I0(n542bar),
    .I1(n541bar)
  );
  //OR U432
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U432 (
    .O(n541),
    .I0(n540),
    .I1(n539)
  );
  //AND U432bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U432bar (
    .O(n541bar),
    .I0(n540bar),
    .I1(n539bar)
  );
  //OR U433
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U433 (
    .O(n539),
    .I0(in[249]),
    .I1(in[242])
  );
  //AND U433bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U433bar (
    .O(n539bar),
    .I0(inbar[249]),
    .I1(inbar[242])
  );
  //OR U434
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U434 (
    .O(n540),
    .I0(in[89]),
    .I1(in[254])
  );
  //AND U434bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U434bar (
    .O(n540bar),
    .I0(inbar[89]),
    .I1(inbar[254])
  );
  //OR U435
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U435 (
    .O(n542),
    .I0(n538),
    .I1(n537)
  );
  //AND U435bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U435bar (
    .O(n542bar),
    .I0(n538bar),
    .I1(n537bar)
  );
  //OR U436
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U436 (
    .O(n537),
    .I0(in_14),
    .I1(in[99])
  );
  //AND U436bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U436bar (
    .O(n537bar),
    .I0(in_14bar),
    .I1(inbar[99])
  );
  //OR U437
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U437 (
    .O(n538),
    .I0(in_60),
    .I1(in_18)
  );
  //AND U437bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U437bar (
    .O(n538bar),
    .I0(in_60bar),
    .I1(in_18bar)
  );
  //OR U438
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U438 (
    .O(n566),
    .I0(in[113]),
    .I1(n763)
  );
  //AND U438bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U438bar (
    .O(n566bar),
    .I0(inbar[113]),
    .I1(n763bar)
  );
  //OR U439
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U439 (
    .O(n763),
    .I0(n536),
    .I1(n535)
  );
  //AND U439bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U439bar (
    .O(n763bar),
    .I0(n536bar),
    .I1(n535bar)
  );
  //OR U440
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U440 (
    .O(n535),
    .I0(n534),
    .I1(n533)
  );
  //AND U440bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U440bar (
    .O(n535bar),
    .I0(n534bar),
    .I1(n533bar)
  );
  //OR U441
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U441 (
    .O(n533),
    .I0(n532),
    .I1(n531)
  );
  //AND U441bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U441bar (
    .O(n533bar),
    .I0(n532bar),
    .I1(n531bar)
  );
  //OR U442
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U442 (
    .O(n531),
    .I0(in[115]),
    .I1(in[110])
  );
  //AND U442bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U442bar (
    .O(n531bar),
    .I0(inbar[115]),
    .I1(inbar[110])
  );
  //OR U443
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U443 (
    .O(n532),
    .I0(in[125]),
    .I1(in[117])
  );
  //AND U443bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U443bar (
    .O(n532bar),
    .I0(inbar[125]),
    .I1(inbar[117])
  );
  //OR U444
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U444 (
    .O(n534),
    .I0(n530),
    .I1(n529)
  );
  //AND U444bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U444bar (
    .O(n534bar),
    .I0(n530bar),
    .I1(n529bar)
  );
  //OR U445
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U445 (
    .O(n529),
    .I0(in[180]),
    .I1(in[128])
  );
  //AND U445bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U445bar (
    .O(n529bar),
    .I0(inbar[180]),
    .I1(inbar[128])
  );
  //OR U446
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U446 (
    .O(n530),
    .I0(in[205]),
    .I1(in[201])
  );
  //AND U446bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U446bar (
    .O(n530bar),
    .I0(inbar[205]),
    .I1(inbar[201])
  );
  //OR U447
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U447 (
    .O(n536),
    .I0(n528),
    .I1(n527)
  );
  //AND U447bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U447bar (
    .O(n536bar),
    .I0(n528bar),
    .I1(n527bar)
  );
  //OR U448
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U448 (
    .O(n527),
    .I0(n526),
    .I1(n525)
  );
  //AND U448bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U448bar (
    .O(n527bar),
    .I0(n526bar),
    .I1(n525bar)
  );
  //OR U449
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U449 (
    .O(n525),
    .I0(in[244]),
    .I1(in[239])
  );
  //AND U449bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U449bar (
    .O(n525bar),
    .I0(inbar[244]),
    .I1(inbar[239])
  );
  //OR U450
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U450 (
    .O(n526),
    .I0(in[95]),
    .I1(in[83])
  );
  //AND U450bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U450bar (
    .O(n526bar),
    .I0(inbar[95]),
    .I1(inbar[83])
  );
  //OR U451
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U451 (
    .O(n528),
    .I0(n524),
    .I1(n523)
  );
  //AND U451bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U451bar (
    .O(n528bar),
    .I0(n524bar),
    .I1(n523bar)
  );
  //OR U452
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U452 (
    .O(n523),
    .I0(in_24),
    .I1(in[97])
  );
  //AND U452bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U452bar (
    .O(n523bar),
    .I0(in_24bar),
    .I1(inbar[97])
  );
  //OR U453
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U453 (
    .O(n524),
    .I0(in_33),
    .I1(in_27)
  );
  //AND U453bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U453bar (
    .O(n524bar),
    .I0(in_33bar),
    .I1(in_27bar)
  );
  //OR U454
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U454 (
    .O(n568),
    .I0(n522),
    .I1(n521)
  );
  //AND U454bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U454bar (
    .O(n568bar),
    .I0(n522bar),
    .I1(n521bar)
  );
  //OR U455
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U455 (
    .O(n521),
    .I0(in[145]),
    .I1(in[126])
  );
  //AND U455bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U455bar (
    .O(n521bar),
    .I0(inbar[145]),
    .I1(inbar[126])
  );
  //OR U456
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U456 (
    .O(n522),
    .I0(in[169]),
    .I1(n520)
  );
  //AND U456bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U456bar (
    .O(n522bar),
    .I0(inbar[169]),
    .I1(n520bar)
  );
  //OR U457
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U457 (
    .O(n520),
    .I0(in[221]),
    .I1(in[172])
  );
  //AND U457bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U457bar (
    .O(n520bar),
    .I0(inbar[221]),
    .I1(inbar[172])
  );
  //OR U458
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U458 (
    .O(n570),
    .I0(n519),
    .I1(n518)
  );
  //AND U458bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U458bar (
    .O(n570bar),
    .I0(n519bar),
    .I1(n518bar)
  );
  //OR U459
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U459 (
    .O(n518),
    .I0(n517),
    .I1(n516)
  );
  //AND U459bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U459bar (
    .O(n518bar),
    .I0(n517bar),
    .I1(n516bar)
  );
  //OR U460
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U460 (
    .O(n516),
    .I0(in[241]),
    .I1(in[224])
  );
  //AND U460bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U460bar (
    .O(n516bar),
    .I0(inbar[241]),
    .I1(inbar[224])
  );
  //OR U461
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U461 (
    .O(n517),
    .I0(in[86]),
    .I1(n515)
  );
  //AND U461bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U461bar (
    .O(n517bar),
    .I0(inbar[86]),
    .I1(n515bar)
  );
  //OR U462
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U462 (
    .O(n515),
    .I0(in_43),
    .I1(in_34)
  );
  //AND U462bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U462bar (
    .O(n515bar),
    .I0(in_43bar),
    .I1(in_34bar)
  );
  //OR U463
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U463 (
    .O(n519),
    .I0(n514),
    .I1(n513)
  );
  //AND U463bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U463bar (
    .O(n519bar),
    .I0(n514bar),
    .I1(n513bar)
  );
  //OR U464
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U464 (
    .O(n513),
    .I0(in_65),
    .I1(in_51)
  );
  //AND U464bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U464bar (
    .O(n513bar),
    .I0(in_65bar),
    .I1(in_51bar)
  );
  //OR U465
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U465 (
    .O(n514),
    .I0(in_75),
    .I1(n512)
  );
  //AND U465bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U465bar (
    .O(n514bar),
    .I0(in_75bar),
    .I1(n512bar)
  );
  //OR U466
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U466 (
    .O(n512),
    .I0(in_81),
    .I1(in_77)
  );
  //AND U466bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U466bar (
    .O(n512bar),
    .I0(in_81bar),
    .I1(in_77bar)
  );
  //OR U467
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U467 (
    .O(n778),
    .I0(n511),
    .I1(n510)
  );
  //AND U467bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U467bar (
    .O(n778bar),
    .I0(n511bar),
    .I1(n510bar)
  );
  //OR U468
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U468 (
    .O(n510),
    .I0(n509),
    .I1(n508)
  );
  //AND U468bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U468bar (
    .O(n510bar),
    .I0(n509bar),
    .I1(n508bar)
  );
  //OR U469
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U469 (
    .O(n508),
    .I0(n507),
    .I1(n506)
  );
  //AND U469bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U469bar (
    .O(n508bar),
    .I0(n507bar),
    .I1(n506bar)
  );
  //OR U470
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U470 (
    .O(n506),
    .I0(in[107]),
    .I1(in[101])
  );
  //AND U470bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U470bar (
    .O(n506bar),
    .I0(inbar[107]),
    .I1(inbar[101])
  );
  //OR U471
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U471 (
    .O(n507),
    .I0(in[139]),
    .I1(in[132])
  );
  //AND U471bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U471bar (
    .O(n507bar),
    .I0(inbar[139]),
    .I1(inbar[132])
  );
  //OR U472
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U472 (
    .O(n509),
    .I0(n505),
    .I1(n504)
  );
  //AND U472bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U472bar (
    .O(n509bar),
    .I0(n505bar),
    .I1(n504bar)
  );
  //OR U473
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U473 (
    .O(n504),
    .I0(in[146]),
    .I1(in[141])
  );
  //AND U473bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U473bar (
    .O(n504bar),
    .I0(inbar[146]),
    .I1(inbar[141])
  );
  //OR U474
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U474 (
    .O(n505),
    .I0(in[203]),
    .I1(in[179])
  );
  //AND U474bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U474bar (
    .O(n505bar),
    .I0(inbar[203]),
    .I1(inbar[179])
  );
  //OR U475
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U475 (
    .O(n511),
    .I0(n503),
    .I1(n502)
  );
  //AND U475bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U475bar (
    .O(n511bar),
    .I0(n503bar),
    .I1(n502bar)
  );
  //OR U476
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U476 (
    .O(n502),
    .I0(n501),
    .I1(n500)
  );
  //AND U476bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U476bar (
    .O(n502bar),
    .I0(n501bar),
    .I1(n500bar)
  );
  //OR U477
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U477 (
    .O(n500),
    .I0(in[243]),
    .I1(in[222])
  );
  //AND U477bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U477bar (
    .O(n500bar),
    .I0(inbar[243]),
    .I1(inbar[222])
  );
  //OR U478
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U478 (
    .O(n501),
    .I0(in[251]),
    .I1(in[250])
  );
  //AND U478bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U478bar (
    .O(n501bar),
    .I0(inbar[251]),
    .I1(inbar[250])
  );
  //OR U479
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U479 (
    .O(n503),
    .I0(n499),
    .I1(n498)
  );
  //AND U479bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U479bar (
    .O(n503bar),
    .I0(n499bar),
    .I1(n498bar)
  );
  //OR U480
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U480 (
    .O(n498),
    .I0(in_37),
    .I1(in_19)
  );
  //AND U480bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U480bar (
    .O(n498bar),
    .I0(in_37bar),
    .I1(in_19bar)
  );
  //OR U481
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U481 (
    .O(n499),
    .I0(in_78),
    .I1(in_6)
  );
  //AND U481bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U481bar (
    .O(n499bar),
    .I0(in_78bar),
    .I1(in_6bar)
  );
  //OR U482
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U482 (
    .O(n603),
    .I0(n497),
    .I1(n496)
  );
  //AND U482bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U482bar (
    .O(n603bar),
    .I0(n497bar),
    .I1(n496bar)
  );
  //OR U483
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U483 (
    .O(n496),
    .I0(in[112]),
    .I1(in[102])
  );
  //AND U483bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U483bar (
    .O(n496bar),
    .I0(inbar[112]),
    .I1(inbar[102])
  );
  //OR U484
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U484 (
    .O(n497),
    .I0(in[123]),
    .I1(n495)
  );
  //AND U484bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U484bar (
    .O(n497bar),
    .I0(inbar[123]),
    .I1(n495bar)
  );
  //OR U485
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U485 (
    .O(n495),
    .I0(in[143]),
    .I1(in[130])
  );
  //AND U485bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U485bar (
    .O(n495bar),
    .I0(inbar[143]),
    .I1(inbar[130])
  );
  //OR U486
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U486 (
    .O(n605),
    .I0(n494),
    .I1(n493)
  );
  //AND U486bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U486bar (
    .O(n605bar),
    .I0(n494bar),
    .I1(n493bar)
  );
  //OR U487
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U487 (
    .O(n493),
    .I0(n492),
    .I1(n491)
  );
  //AND U487bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U487bar (
    .O(n493bar),
    .I0(n492bar),
    .I1(n491bar)
  );
  //OR U488
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U488 (
    .O(n491),
    .I0(in[216]),
    .I1(in[213])
  );
  //AND U488bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U488bar (
    .O(n491bar),
    .I0(inbar[216]),
    .I1(inbar[213])
  );
  //OR U489
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U489 (
    .O(n492),
    .I0(in[227]),
    .I1(n490)
  );
  //AND U489bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U489bar (
    .O(n492bar),
    .I0(inbar[227]),
    .I1(n490bar)
  );
  //OR U490
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U490 (
    .O(n490),
    .I0(in_0),
    .I1(in[248])
  );
  //AND U490bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U490bar (
    .O(n490bar),
    .I0(in_0bar),
    .I1(inbar[248])
  );
  //OR U491
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U491 (
    .O(n494),
    .I0(n489),
    .I1(n488)
  );
  //AND U491bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U491bar (
    .O(n494bar),
    .I0(n489bar),
    .I1(n488bar)
  );
  //OR U492
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U492 (
    .O(n488),
    .I0(in_46),
    .I1(in_44)
  );
  //AND U492bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U492bar (
    .O(n488bar),
    .I0(in_46bar),
    .I1(in_44bar)
  );
  //OR U493
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U493 (
    .O(n489),
    .I0(in_50),
    .I1(n487)
  );
  //AND U493bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U493bar (
    .O(n489bar),
    .I0(in_50bar),
    .I1(n487bar)
  );
  //OR U494
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U494 (
    .O(n487),
    .I0(in_9),
    .I1(in_80)
  );
  //AND U494bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U494bar (
    .O(n487bar),
    .I0(in_9bar),
    .I1(in_80bar)
  );
endmodule

module sBox_1 ( in, out );

  input wire [7:0] in;
//input_done

  output wire [7:0] out;
//output_done

  wire [255:0] decodeOut;
//wire_done

  decode_1 dec ( .in(in), .out(decodeOut) );
  encode_1 enc ( .in(decodeOut), .out(out) );
endmodule

module CD2_5 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD2_6 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD2_7 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD2_8 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD4_3 ( a, b, y );

  input wire [3:0] a;
  input wire [3:0] b;
  wire [3:0] abar;
  wire [3:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
//input_done

  output wire [15:0] y;
  wire [15:0] ybar;
//output_done

//wire_done

  //AND U1
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1 (
    .O(y[9]),
    .I0(b[1]),
    .I1(a[2])
  );
  //OR U1bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1bar (
    .O(ybar[9]),
    .I0(bbar[1]),
    .I1(abar[2])
  );
  //AND U2
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2 (
    .O(y[8]),
    .I0(b[0]),
    .I1(a[2])
  );
  //OR U2bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2bar (
    .O(ybar[8]),
    .I0(bbar[0]),
    .I1(abar[2])
  );
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[7]),
    .I0(b[3]),
    .I1(a[1])
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[7]),
    .I0(bbar[3]),
    .I1(abar[1])
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[6]),
    .I0(b[2]),
    .I1(a[1])
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[6]),
    .I0(bbar[2]),
    .I1(abar[1])
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[5]),
    .I0(a[1]),
    .I1(b[1])
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[5]),
    .I0(abar[1]),
    .I1(bbar[1])
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[4]),
    .I0(a[1]),
    .I1(b[0])
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[4]),
    .I0(abar[1]),
    .I1(bbar[0])
  );
  //AND U7
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7 (
    .O(y[3]),
    .I0(a[0]),
    .I1(b[3])
  );
  //OR U7bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7bar (
    .O(ybar[3]),
    .I0(abar[0]),
    .I1(bbar[3])
  );
  //AND U8
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8 (
    .O(y[2]),
    .I0(a[0]),
    .I1(b[2])
  );
  //OR U8bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8bar (
    .O(ybar[2]),
    .I0(abar[0]),
    .I1(bbar[2])
  );
  //AND U9
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9 (
    .O(y[1]),
    .I0(a[0]),
    .I1(b[1])
  );
  //OR U9bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9bar (
    .O(ybar[1]),
    .I0(abar[0]),
    .I1(bbar[1])
  );
  //AND U10
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10 (
    .O(y[15]),
    .I0(a[3]),
    .I1(b[3])
  );
  //OR U10bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10bar (
    .O(ybar[15]),
    .I0(abar[3]),
    .I1(bbar[3])
  );
  //AND U11
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11 (
    .O(y[14]),
    .I0(a[3]),
    .I1(b[2])
  );
  //OR U11bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11bar (
    .O(ybar[14]),
    .I0(abar[3]),
    .I1(bbar[2])
  );
  //AND U12
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12 (
    .O(y[13]),
    .I0(a[3]),
    .I1(b[1])
  );
  //OR U12bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12bar (
    .O(ybar[13]),
    .I0(abar[3]),
    .I1(bbar[1])
  );
  //AND U13
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13 (
    .O(y[12]),
    .I0(a[3]),
    .I1(b[0])
  );
  //OR U13bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13bar (
    .O(ybar[12]),
    .I0(abar[3]),
    .I1(bbar[0])
  );
  //AND U14
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14 (
    .O(y[11]),
    .I0(b[3]),
    .I1(a[2])
  );
  //OR U14bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14bar (
    .O(ybar[11]),
    .I0(bbar[3]),
    .I1(abar[2])
  );
  //AND U15
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15 (
    .O(y[10]),
    .I0(b[2]),
    .I1(a[2])
  );
  //OR U15bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15bar (
    .O(ybar[10]),
    .I0(bbar[2]),
    .I1(abar[2])
  );
  //AND U16
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16 (
    .O(y[0]),
    .I0(a[0]),
    .I1(b[0])
  );
  //OR U16bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16bar (
    .O(ybar[0]),
    .I0(abar[0]),
    .I1(bbar[0])
  );
endmodule

module CD4_4 ( a, b, y );

  input wire [3:0] a;
  input wire [3:0] b;
  wire [3:0] abar;
  wire [3:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
//input_done

  output wire [15:0] y;
  wire [15:0] ybar;
//output_done

//wire_done

  //AND U1
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1 (
    .O(y[9]),
    .I0(b[1]),
    .I1(a[2])
  );
  //OR U1bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1bar (
    .O(ybar[9]),
    .I0(bbar[1]),
    .I1(abar[2])
  );
  //AND U2
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2 (
    .O(y[8]),
    .I0(b[0]),
    .I1(a[2])
  );
  //OR U2bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2bar (
    .O(ybar[8]),
    .I0(bbar[0]),
    .I1(abar[2])
  );
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[7]),
    .I0(b[3]),
    .I1(a[1])
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[7]),
    .I0(bbar[3]),
    .I1(abar[1])
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[6]),
    .I0(b[2]),
    .I1(a[1])
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[6]),
    .I0(bbar[2]),
    .I1(abar[1])
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[5]),
    .I0(a[1]),
    .I1(b[1])
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[5]),
    .I0(abar[1]),
    .I1(bbar[1])
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[4]),
    .I0(a[1]),
    .I1(b[0])
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[4]),
    .I0(abar[1]),
    .I1(bbar[0])
  );
  //AND U7
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7 (
    .O(y[3]),
    .I0(a[0]),
    .I1(b[3])
  );
  //OR U7bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7bar (
    .O(ybar[3]),
    .I0(abar[0]),
    .I1(bbar[3])
  );
  //AND U8
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8 (
    .O(y[2]),
    .I0(a[0]),
    .I1(b[2])
  );
  //OR U8bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8bar (
    .O(ybar[2]),
    .I0(abar[0]),
    .I1(bbar[2])
  );
  //AND U9
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9 (
    .O(y[1]),
    .I0(a[0]),
    .I1(b[1])
  );
  //OR U9bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9bar (
    .O(ybar[1]),
    .I0(abar[0]),
    .I1(bbar[1])
  );
  //AND U10
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10 (
    .O(y[15]),
    .I0(a[3]),
    .I1(b[3])
  );
  //OR U10bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10bar (
    .O(ybar[15]),
    .I0(abar[3]),
    .I1(bbar[3])
  );
  //AND U11
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11 (
    .O(y[14]),
    .I0(a[3]),
    .I1(b[2])
  );
  //OR U11bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11bar (
    .O(ybar[14]),
    .I0(abar[3]),
    .I1(bbar[2])
  );
  //AND U12
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12 (
    .O(y[13]),
    .I0(a[3]),
    .I1(b[1])
  );
  //OR U12bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12bar (
    .O(ybar[13]),
    .I0(abar[3]),
    .I1(bbar[1])
  );
  //AND U13
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13 (
    .O(y[12]),
    .I0(a[3]),
    .I1(b[0])
  );
  //OR U13bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13bar (
    .O(ybar[12]),
    .I0(abar[3]),
    .I1(bbar[0])
  );
  //AND U14
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14 (
    .O(y[11]),
    .I0(b[3]),
    .I1(a[2])
  );
  //OR U14bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14bar (
    .O(ybar[11]),
    .I0(bbar[3]),
    .I1(abar[2])
  );
  //AND U15
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15 (
    .O(y[10]),
    .I0(b[2]),
    .I1(a[2])
  );
  //OR U15bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15bar (
    .O(ybar[10]),
    .I0(bbar[2]),
    .I1(abar[2])
  );
  //AND U16
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16 (
    .O(y[0]),
    .I0(a[0]),
    .I1(b[0])
  );
  //OR U16bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16bar (
    .O(ybar[0]),
    .I0(abar[0]),
    .I1(bbar[0])
  );
endmodule

module CD16_2 ( a, b, y );

  input wire [15:0] a;
  input wire [15:0] b;
  wire [15:0] abar;
  wire [15:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign abar[8] = ~a[8];
  assign abar[9] = ~a[9];
  assign abar[10] = ~a[10];
  assign abar[11] = ~a[11];
  assign abar[12] = ~a[12];
  assign abar[13] = ~a[13];
  assign abar[14] = ~a[14];
  assign abar[15] = ~a[15];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign bbar[8] = ~b[8];
  assign bbar[9] = ~b[9];
  assign bbar[10] = ~b[10];
  assign bbar[11] = ~b[11];
  assign bbar[12] = ~b[12];
  assign bbar[13] = ~b[13];
  assign bbar[14] = ~b[14];
  assign bbar[15] = ~b[15];
//input_done

  output wire [255:0] y;
  wire [255:0] ybar;
//output_done

//wire_done

  //AND U1
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1 (
    .O(y[9]),
    .I0(b[9]),
    .I1(a[0])
  );
  //OR U1bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1bar (
    .O(ybar[9]),
    .I0(bbar[9]),
    .I1(abar[0])
  );
  //AND U2
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2 (
    .O(y[99]),
    .I0(b[3]),
    .I1(a[6])
  );
  //OR U2bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2bar (
    .O(ybar[99]),
    .I0(bbar[3]),
    .I1(abar[6])
  );
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[98]),
    .I0(b[2]),
    .I1(a[6])
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[98]),
    .I0(bbar[2]),
    .I1(abar[6])
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[97]),
    .I0(b[1]),
    .I1(a[6])
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[97]),
    .I0(bbar[1]),
    .I1(abar[6])
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[96]),
    .I0(b[0]),
    .I1(a[6])
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[96]),
    .I0(bbar[0]),
    .I1(abar[6])
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[95]),
    .I0(b[15]),
    .I1(a[5])
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[95]),
    .I0(bbar[15]),
    .I1(abar[5])
  );
  //AND U7
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7 (
    .O(y[94]),
    .I0(b[14]),
    .I1(a[5])
  );
  //OR U7bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7bar (
    .O(ybar[94]),
    .I0(bbar[14]),
    .I1(abar[5])
  );
  //AND U8
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8 (
    .O(y[93]),
    .I0(b[13]),
    .I1(a[5])
  );
  //OR U8bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8bar (
    .O(ybar[93]),
    .I0(bbar[13]),
    .I1(abar[5])
  );
  //AND U9
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9 (
    .O(y[92]),
    .I0(b[12]),
    .I1(a[5])
  );
  //OR U9bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9bar (
    .O(ybar[92]),
    .I0(bbar[12]),
    .I1(abar[5])
  );
  //AND U10
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10 (
    .O(y[91]),
    .I0(b[11]),
    .I1(a[5])
  );
  //OR U10bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10bar (
    .O(ybar[91]),
    .I0(bbar[11]),
    .I1(abar[5])
  );
  //AND U11
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11 (
    .O(y[90]),
    .I0(b[10]),
    .I1(a[5])
  );
  //OR U11bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11bar (
    .O(ybar[90]),
    .I0(bbar[10]),
    .I1(abar[5])
  );
  //AND U12
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12 (
    .O(y[8]),
    .I0(b[8]),
    .I1(a[0])
  );
  //OR U12bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12bar (
    .O(ybar[8]),
    .I0(bbar[8]),
    .I1(abar[0])
  );
  //AND U13
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13 (
    .O(y[89]),
    .I0(a[5]),
    .I1(b[9])
  );
  //OR U13bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13bar (
    .O(ybar[89]),
    .I0(abar[5]),
    .I1(bbar[9])
  );
  //AND U14
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14 (
    .O(y[88]),
    .I0(b[8]),
    .I1(a[5])
  );
  //OR U14bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14bar (
    .O(ybar[88]),
    .I0(bbar[8]),
    .I1(abar[5])
  );
  //AND U15
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15 (
    .O(y[87]),
    .I0(b[7]),
    .I1(a[5])
  );
  //OR U15bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15bar (
    .O(ybar[87]),
    .I0(bbar[7]),
    .I1(abar[5])
  );
  //AND U16
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16 (
    .O(y[86]),
    .I0(b[6]),
    .I1(a[5])
  );
  //OR U16bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16bar (
    .O(ybar[86]),
    .I0(bbar[6]),
    .I1(abar[5])
  );
  //AND U17
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U17 (
    .O(y[85]),
    .I0(b[5]),
    .I1(a[5])
  );
  //OR U17bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U17bar (
    .O(ybar[85]),
    .I0(bbar[5]),
    .I1(abar[5])
  );
  //AND U18
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U18 (
    .O(y[84]),
    .I0(b[4]),
    .I1(a[5])
  );
  //OR U18bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U18bar (
    .O(ybar[84]),
    .I0(bbar[4]),
    .I1(abar[5])
  );
  //AND U19
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U19 (
    .O(y[83]),
    .I0(a[5]),
    .I1(b[3])
  );
  //OR U19bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U19bar (
    .O(ybar[83]),
    .I0(abar[5]),
    .I1(bbar[3])
  );
  //AND U20
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U20 (
    .O(y[82]),
    .I0(a[5]),
    .I1(b[2])
  );
  //OR U20bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U20bar (
    .O(ybar[82]),
    .I0(abar[5]),
    .I1(bbar[2])
  );
  //AND U21
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U21 (
    .O(y[81]),
    .I0(a[5]),
    .I1(b[1])
  );
  //OR U21bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U21bar (
    .O(ybar[81]),
    .I0(abar[5]),
    .I1(bbar[1])
  );
  //AND U22
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U22 (
    .O(y[80]),
    .I0(a[5]),
    .I1(b[0])
  );
  //OR U22bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U22bar (
    .O(ybar[80]),
    .I0(abar[5]),
    .I1(bbar[0])
  );
  //AND U23
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U23 (
    .O(y[7]),
    .I0(b[7]),
    .I1(a[0])
  );
  //OR U23bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U23bar (
    .O(ybar[7]),
    .I0(bbar[7]),
    .I1(abar[0])
  );
  //AND U24
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U24 (
    .O(y[79]),
    .I0(a[4]),
    .I1(b[15])
  );
  //OR U24bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U24bar (
    .O(ybar[79]),
    .I0(abar[4]),
    .I1(bbar[15])
  );
  //AND U25
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U25 (
    .O(y[78]),
    .I0(a[4]),
    .I1(b[14])
  );
  //OR U25bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U25bar (
    .O(ybar[78]),
    .I0(abar[4]),
    .I1(bbar[14])
  );
  //AND U26
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U26 (
    .O(y[77]),
    .I0(a[4]),
    .I1(b[13])
  );
  //OR U26bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U26bar (
    .O(ybar[77]),
    .I0(abar[4]),
    .I1(bbar[13])
  );
  //AND U27
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U27 (
    .O(y[76]),
    .I0(a[4]),
    .I1(b[12])
  );
  //OR U27bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U27bar (
    .O(ybar[76]),
    .I0(abar[4]),
    .I1(bbar[12])
  );
  //AND U28
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U28 (
    .O(y[75]),
    .I0(a[4]),
    .I1(b[11])
  );
  //OR U28bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U28bar (
    .O(ybar[75]),
    .I0(abar[4]),
    .I1(bbar[11])
  );
  //AND U29
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U29 (
    .O(y[74]),
    .I0(a[4]),
    .I1(b[10])
  );
  //OR U29bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U29bar (
    .O(ybar[74]),
    .I0(abar[4]),
    .I1(bbar[10])
  );
  //AND U30
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U30 (
    .O(y[73]),
    .I0(a[4]),
    .I1(b[9])
  );
  //OR U30bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U30bar (
    .O(ybar[73]),
    .I0(abar[4]),
    .I1(bbar[9])
  );
  //AND U31
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U31 (
    .O(y[72]),
    .I0(a[4]),
    .I1(b[8])
  );
  //OR U31bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U31bar (
    .O(ybar[72]),
    .I0(abar[4]),
    .I1(bbar[8])
  );
  //AND U32
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U32 (
    .O(y[71]),
    .I0(a[4]),
    .I1(b[7])
  );
  //OR U32bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U32bar (
    .O(ybar[71]),
    .I0(abar[4]),
    .I1(bbar[7])
  );
  //AND U33
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U33 (
    .O(y[70]),
    .I0(a[4]),
    .I1(b[6])
  );
  //OR U33bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U33bar (
    .O(ybar[70]),
    .I0(abar[4]),
    .I1(bbar[6])
  );
  //AND U34
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U34 (
    .O(y[6]),
    .I0(b[6]),
    .I1(a[0])
  );
  //OR U34bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U34bar (
    .O(ybar[6]),
    .I0(bbar[6]),
    .I1(abar[0])
  );
  //AND U35
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U35 (
    .O(y[69]),
    .I0(a[4]),
    .I1(b[5])
  );
  //OR U35bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U35bar (
    .O(ybar[69]),
    .I0(abar[4]),
    .I1(bbar[5])
  );
  //AND U36
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U36 (
    .O(y[68]),
    .I0(a[4]),
    .I1(b[4])
  );
  //OR U36bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U36bar (
    .O(ybar[68]),
    .I0(abar[4]),
    .I1(bbar[4])
  );
  //AND U37
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U37 (
    .O(y[67]),
    .I0(a[4]),
    .I1(b[3])
  );
  //OR U37bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U37bar (
    .O(ybar[67]),
    .I0(abar[4]),
    .I1(bbar[3])
  );
  //AND U38
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U38 (
    .O(y[66]),
    .I0(a[4]),
    .I1(b[2])
  );
  //OR U38bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U38bar (
    .O(ybar[66]),
    .I0(abar[4]),
    .I1(bbar[2])
  );
  //AND U39
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U39 (
    .O(y[65]),
    .I0(a[4]),
    .I1(b[1])
  );
  //OR U39bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U39bar (
    .O(ybar[65]),
    .I0(abar[4]),
    .I1(bbar[1])
  );
  //AND U40
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U40 (
    .O(y[64]),
    .I0(a[4]),
    .I1(b[0])
  );
  //OR U40bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U40bar (
    .O(ybar[64]),
    .I0(abar[4]),
    .I1(bbar[0])
  );
  //AND U41
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U41 (
    .O(y[63]),
    .I0(a[3]),
    .I1(b[15])
  );
  //OR U41bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U41bar (
    .O(ybar[63]),
    .I0(abar[3]),
    .I1(bbar[15])
  );
  //AND U42
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U42 (
    .O(y[62]),
    .I0(a[3]),
    .I1(b[14])
  );
  //OR U42bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U42bar (
    .O(ybar[62]),
    .I0(abar[3]),
    .I1(bbar[14])
  );
  //AND U43
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U43 (
    .O(y[61]),
    .I0(a[3]),
    .I1(b[13])
  );
  //OR U43bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U43bar (
    .O(ybar[61]),
    .I0(abar[3]),
    .I1(bbar[13])
  );
  //AND U44
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U44 (
    .O(y[60]),
    .I0(a[3]),
    .I1(b[12])
  );
  //OR U44bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U44bar (
    .O(ybar[60]),
    .I0(abar[3]),
    .I1(bbar[12])
  );
  //AND U45
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U45 (
    .O(y[5]),
    .I0(b[5]),
    .I1(a[0])
  );
  //OR U45bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U45bar (
    .O(ybar[5]),
    .I0(bbar[5]),
    .I1(abar[0])
  );
  //AND U46
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U46 (
    .O(y[59]),
    .I0(a[3]),
    .I1(b[11])
  );
  //OR U46bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U46bar (
    .O(ybar[59]),
    .I0(abar[3]),
    .I1(bbar[11])
  );
  //AND U47
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U47 (
    .O(y[58]),
    .I0(a[3]),
    .I1(b[10])
  );
  //OR U47bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U47bar (
    .O(ybar[58]),
    .I0(abar[3]),
    .I1(bbar[10])
  );
  //AND U48
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U48 (
    .O(y[57]),
    .I0(a[3]),
    .I1(b[9])
  );
  //OR U48bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U48bar (
    .O(ybar[57]),
    .I0(abar[3]),
    .I1(bbar[9])
  );
  //AND U49
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U49 (
    .O(y[56]),
    .I0(a[3]),
    .I1(b[8])
  );
  //OR U49bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U49bar (
    .O(ybar[56]),
    .I0(abar[3]),
    .I1(bbar[8])
  );
  //AND U50
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U50 (
    .O(y[55]),
    .I0(a[3]),
    .I1(b[7])
  );
  //OR U50bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U50bar (
    .O(ybar[55]),
    .I0(abar[3]),
    .I1(bbar[7])
  );
  //AND U51
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U51 (
    .O(y[54]),
    .I0(a[3]),
    .I1(b[6])
  );
  //OR U51bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U51bar (
    .O(ybar[54]),
    .I0(abar[3]),
    .I1(bbar[6])
  );
  //AND U52
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U52 (
    .O(y[53]),
    .I0(a[3]),
    .I1(b[5])
  );
  //OR U52bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U52bar (
    .O(ybar[53]),
    .I0(abar[3]),
    .I1(bbar[5])
  );
  //AND U53
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U53 (
    .O(y[52]),
    .I0(a[3]),
    .I1(b[4])
  );
  //OR U53bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U53bar (
    .O(ybar[52]),
    .I0(abar[3]),
    .I1(bbar[4])
  );
  //AND U54
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U54 (
    .O(y[51]),
    .I0(a[3]),
    .I1(b[3])
  );
  //OR U54bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U54bar (
    .O(ybar[51]),
    .I0(abar[3]),
    .I1(bbar[3])
  );
  //AND U55
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U55 (
    .O(y[50]),
    .I0(a[3]),
    .I1(b[2])
  );
  //OR U55bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U55bar (
    .O(ybar[50]),
    .I0(abar[3]),
    .I1(bbar[2])
  );
  //AND U56
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U56 (
    .O(y[4]),
    .I0(b[4]),
    .I1(a[0])
  );
  //OR U56bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U56bar (
    .O(ybar[4]),
    .I0(bbar[4]),
    .I1(abar[0])
  );
  //AND U57
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U57 (
    .O(y[49]),
    .I0(a[3]),
    .I1(b[1])
  );
  //OR U57bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U57bar (
    .O(ybar[49]),
    .I0(abar[3]),
    .I1(bbar[1])
  );
  //AND U58
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U58 (
    .O(y[48]),
    .I0(a[3]),
    .I1(b[0])
  );
  //OR U58bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U58bar (
    .O(ybar[48]),
    .I0(abar[3]),
    .I1(bbar[0])
  );
  //AND U59
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U59 (
    .O(y[47]),
    .I0(a[2]),
    .I1(b[15])
  );
  //OR U59bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U59bar (
    .O(ybar[47]),
    .I0(abar[2]),
    .I1(bbar[15])
  );
  //AND U60
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U60 (
    .O(y[46]),
    .I0(a[2]),
    .I1(b[14])
  );
  //OR U60bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U60bar (
    .O(ybar[46]),
    .I0(abar[2]),
    .I1(bbar[14])
  );
  //AND U61
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U61 (
    .O(y[45]),
    .I0(a[2]),
    .I1(b[13])
  );
  //OR U61bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U61bar (
    .O(ybar[45]),
    .I0(abar[2]),
    .I1(bbar[13])
  );
  //AND U62
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U62 (
    .O(y[44]),
    .I0(a[2]),
    .I1(b[12])
  );
  //OR U62bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U62bar (
    .O(ybar[44]),
    .I0(abar[2]),
    .I1(bbar[12])
  );
  //AND U63
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U63 (
    .O(y[43]),
    .I0(a[2]),
    .I1(b[11])
  );
  //OR U63bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U63bar (
    .O(ybar[43]),
    .I0(abar[2]),
    .I1(bbar[11])
  );
  //AND U64
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U64 (
    .O(y[42]),
    .I0(a[2]),
    .I1(b[10])
  );
  //OR U64bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U64bar (
    .O(ybar[42]),
    .I0(abar[2]),
    .I1(bbar[10])
  );
  //AND U65
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U65 (
    .O(y[41]),
    .I0(a[2]),
    .I1(b[9])
  );
  //OR U65bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U65bar (
    .O(ybar[41]),
    .I0(abar[2]),
    .I1(bbar[9])
  );
  //AND U66
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U66 (
    .O(y[40]),
    .I0(a[2]),
    .I1(b[8])
  );
  //OR U66bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U66bar (
    .O(ybar[40]),
    .I0(abar[2]),
    .I1(bbar[8])
  );
  //AND U67
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U67 (
    .O(y[3]),
    .I0(b[3]),
    .I1(a[0])
  );
  //OR U67bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U67bar (
    .O(ybar[3]),
    .I0(bbar[3]),
    .I1(abar[0])
  );
  //AND U68
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U68 (
    .O(y[39]),
    .I0(a[2]),
    .I1(b[7])
  );
  //OR U68bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U68bar (
    .O(ybar[39]),
    .I0(abar[2]),
    .I1(bbar[7])
  );
  //AND U69
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U69 (
    .O(y[38]),
    .I0(a[2]),
    .I1(b[6])
  );
  //OR U69bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U69bar (
    .O(ybar[38]),
    .I0(abar[2]),
    .I1(bbar[6])
  );
  //AND U70
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U70 (
    .O(y[37]),
    .I0(a[2]),
    .I1(b[5])
  );
  //OR U70bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U70bar (
    .O(ybar[37]),
    .I0(abar[2]),
    .I1(bbar[5])
  );
  //AND U71
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U71 (
    .O(y[36]),
    .I0(a[2]),
    .I1(b[4])
  );
  //OR U71bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U71bar (
    .O(ybar[36]),
    .I0(abar[2]),
    .I1(bbar[4])
  );
  //AND U72
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U72 (
    .O(y[35]),
    .I0(a[2]),
    .I1(b[3])
  );
  //OR U72bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U72bar (
    .O(ybar[35]),
    .I0(abar[2]),
    .I1(bbar[3])
  );
  //AND U73
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U73 (
    .O(y[34]),
    .I0(a[2]),
    .I1(b[2])
  );
  //OR U73bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U73bar (
    .O(ybar[34]),
    .I0(abar[2]),
    .I1(bbar[2])
  );
  //AND U74
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U74 (
    .O(y[33]),
    .I0(a[2]),
    .I1(b[1])
  );
  //OR U74bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U74bar (
    .O(ybar[33]),
    .I0(abar[2]),
    .I1(bbar[1])
  );
  //AND U75
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U75 (
    .O(y[32]),
    .I0(a[2]),
    .I1(b[0])
  );
  //OR U75bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U75bar (
    .O(ybar[32]),
    .I0(abar[2]),
    .I1(bbar[0])
  );
  //AND U76
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U76 (
    .O(y[31]),
    .I0(a[1]),
    .I1(b[15])
  );
  //OR U76bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U76bar (
    .O(ybar[31]),
    .I0(abar[1]),
    .I1(bbar[15])
  );
  //AND U77
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U77 (
    .O(y[30]),
    .I0(a[1]),
    .I1(b[14])
  );
  //OR U77bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U77bar (
    .O(ybar[30]),
    .I0(abar[1]),
    .I1(bbar[14])
  );
  //AND U78
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U78 (
    .O(y[2]),
    .I0(b[2]),
    .I1(a[0])
  );
  //OR U78bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U78bar (
    .O(ybar[2]),
    .I0(bbar[2]),
    .I1(abar[0])
  );
  //AND U79
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U79 (
    .O(y[29]),
    .I0(a[1]),
    .I1(b[13])
  );
  //OR U79bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U79bar (
    .O(ybar[29]),
    .I0(abar[1]),
    .I1(bbar[13])
  );
  //AND U80
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U80 (
    .O(y[28]),
    .I0(a[1]),
    .I1(b[12])
  );
  //OR U80bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U80bar (
    .O(ybar[28]),
    .I0(abar[1]),
    .I1(bbar[12])
  );
  //AND U81
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U81 (
    .O(y[27]),
    .I0(a[1]),
    .I1(b[11])
  );
  //OR U81bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U81bar (
    .O(ybar[27]),
    .I0(abar[1]),
    .I1(bbar[11])
  );
  //AND U82
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U82 (
    .O(y[26]),
    .I0(a[1]),
    .I1(b[10])
  );
  //OR U82bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U82bar (
    .O(ybar[26]),
    .I0(abar[1]),
    .I1(bbar[10])
  );
  //AND U83
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U83 (
    .O(y[25]),
    .I0(a[1]),
    .I1(b[9])
  );
  //OR U83bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U83bar (
    .O(ybar[25]),
    .I0(abar[1]),
    .I1(bbar[9])
  );
  //AND U84
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U84 (
    .O(y[255]),
    .I0(a[15]),
    .I1(b[15])
  );
  //OR U84bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U84bar (
    .O(ybar[255]),
    .I0(abar[15]),
    .I1(bbar[15])
  );
  //AND U85
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U85 (
    .O(y[254]),
    .I0(a[15]),
    .I1(b[14])
  );
  //OR U85bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U85bar (
    .O(ybar[254]),
    .I0(abar[15]),
    .I1(bbar[14])
  );
  //AND U86
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U86 (
    .O(y[253]),
    .I0(a[15]),
    .I1(b[13])
  );
  //OR U86bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U86bar (
    .O(ybar[253]),
    .I0(abar[15]),
    .I1(bbar[13])
  );
  //AND U87
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U87 (
    .O(y[252]),
    .I0(a[15]),
    .I1(b[12])
  );
  //OR U87bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U87bar (
    .O(ybar[252]),
    .I0(abar[15]),
    .I1(bbar[12])
  );
  //AND U88
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U88 (
    .O(y[251]),
    .I0(a[15]),
    .I1(b[11])
  );
  //OR U88bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U88bar (
    .O(ybar[251]),
    .I0(abar[15]),
    .I1(bbar[11])
  );
  //AND U89
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U89 (
    .O(y[250]),
    .I0(a[15]),
    .I1(b[10])
  );
  //OR U89bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U89bar (
    .O(ybar[250]),
    .I0(abar[15]),
    .I1(bbar[10])
  );
  //AND U90
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U90 (
    .O(y[24]),
    .I0(a[1]),
    .I1(b[8])
  );
  //OR U90bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U90bar (
    .O(ybar[24]),
    .I0(abar[1]),
    .I1(bbar[8])
  );
  //AND U91
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U91 (
    .O(y[249]),
    .I0(a[15]),
    .I1(b[9])
  );
  //OR U91bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U91bar (
    .O(ybar[249]),
    .I0(abar[15]),
    .I1(bbar[9])
  );
  //AND U92
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U92 (
    .O(y[248]),
    .I0(a[15]),
    .I1(b[8])
  );
  //OR U92bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U92bar (
    .O(ybar[248]),
    .I0(abar[15]),
    .I1(bbar[8])
  );
  //AND U93
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U93 (
    .O(y[247]),
    .I0(a[15]),
    .I1(b[7])
  );
  //OR U93bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U93bar (
    .O(ybar[247]),
    .I0(abar[15]),
    .I1(bbar[7])
  );
  //AND U94
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U94 (
    .O(y[246]),
    .I0(a[15]),
    .I1(b[6])
  );
  //OR U94bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U94bar (
    .O(ybar[246]),
    .I0(abar[15]),
    .I1(bbar[6])
  );
  //AND U95
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U95 (
    .O(y[245]),
    .I0(a[15]),
    .I1(b[5])
  );
  //OR U95bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U95bar (
    .O(ybar[245]),
    .I0(abar[15]),
    .I1(bbar[5])
  );
  //AND U96
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U96 (
    .O(y[244]),
    .I0(a[15]),
    .I1(b[4])
  );
  //OR U96bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U96bar (
    .O(ybar[244]),
    .I0(abar[15]),
    .I1(bbar[4])
  );
  //AND U97
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U97 (
    .O(y[243]),
    .I0(a[15]),
    .I1(b[3])
  );
  //OR U97bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U97bar (
    .O(ybar[243]),
    .I0(abar[15]),
    .I1(bbar[3])
  );
  //AND U98
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U98 (
    .O(y[242]),
    .I0(a[15]),
    .I1(b[2])
  );
  //OR U98bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U98bar (
    .O(ybar[242]),
    .I0(abar[15]),
    .I1(bbar[2])
  );
  //AND U99
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U99 (
    .O(y[241]),
    .I0(a[15]),
    .I1(b[1])
  );
  //OR U99bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U99bar (
    .O(ybar[241]),
    .I0(abar[15]),
    .I1(bbar[1])
  );
  //AND U100
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U100 (
    .O(y[240]),
    .I0(a[15]),
    .I1(b[0])
  );
  //OR U100bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U100bar (
    .O(ybar[240]),
    .I0(abar[15]),
    .I1(bbar[0])
  );
  //AND U101
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U101 (
    .O(y[23]),
    .I0(a[1]),
    .I1(b[7])
  );
  //OR U101bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U101bar (
    .O(ybar[23]),
    .I0(abar[1]),
    .I1(bbar[7])
  );
  //AND U102
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U102 (
    .O(y[239]),
    .I0(a[14]),
    .I1(b[15])
  );
  //OR U102bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U102bar (
    .O(ybar[239]),
    .I0(abar[14]),
    .I1(bbar[15])
  );
  //AND U103
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U103 (
    .O(y[238]),
    .I0(a[14]),
    .I1(b[14])
  );
  //OR U103bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U103bar (
    .O(ybar[238]),
    .I0(abar[14]),
    .I1(bbar[14])
  );
  //AND U104
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U104 (
    .O(y[237]),
    .I0(a[14]),
    .I1(b[13])
  );
  //OR U104bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U104bar (
    .O(ybar[237]),
    .I0(abar[14]),
    .I1(bbar[13])
  );
  //AND U105
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U105 (
    .O(y[236]),
    .I0(a[14]),
    .I1(b[12])
  );
  //OR U105bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U105bar (
    .O(ybar[236]),
    .I0(abar[14]),
    .I1(bbar[12])
  );
  //AND U106
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U106 (
    .O(y[235]),
    .I0(a[14]),
    .I1(b[11])
  );
  //OR U106bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U106bar (
    .O(ybar[235]),
    .I0(abar[14]),
    .I1(bbar[11])
  );
  //AND U107
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U107 (
    .O(y[234]),
    .I0(a[14]),
    .I1(b[10])
  );
  //OR U107bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U107bar (
    .O(ybar[234]),
    .I0(abar[14]),
    .I1(bbar[10])
  );
  //AND U108
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U108 (
    .O(y[233]),
    .I0(a[14]),
    .I1(b[9])
  );
  //OR U108bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U108bar (
    .O(ybar[233]),
    .I0(abar[14]),
    .I1(bbar[9])
  );
  //AND U109
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U109 (
    .O(y[232]),
    .I0(a[14]),
    .I1(b[8])
  );
  //OR U109bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U109bar (
    .O(ybar[232]),
    .I0(abar[14]),
    .I1(bbar[8])
  );
  //AND U110
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U110 (
    .O(y[231]),
    .I0(a[14]),
    .I1(b[7])
  );
  //OR U110bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U110bar (
    .O(ybar[231]),
    .I0(abar[14]),
    .I1(bbar[7])
  );
  //AND U111
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U111 (
    .O(y[230]),
    .I0(a[14]),
    .I1(b[6])
  );
  //OR U111bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U111bar (
    .O(ybar[230]),
    .I0(abar[14]),
    .I1(bbar[6])
  );
  //AND U112
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U112 (
    .O(y[22]),
    .I0(a[1]),
    .I1(b[6])
  );
  //OR U112bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U112bar (
    .O(ybar[22]),
    .I0(abar[1]),
    .I1(bbar[6])
  );
  //AND U113
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U113 (
    .O(y[229]),
    .I0(a[14]),
    .I1(b[5])
  );
  //OR U113bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U113bar (
    .O(ybar[229]),
    .I0(abar[14]),
    .I1(bbar[5])
  );
  //AND U114
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U114 (
    .O(y[228]),
    .I0(a[14]),
    .I1(b[4])
  );
  //OR U114bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U114bar (
    .O(ybar[228]),
    .I0(abar[14]),
    .I1(bbar[4])
  );
  //AND U115
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U115 (
    .O(y[227]),
    .I0(a[14]),
    .I1(b[3])
  );
  //OR U115bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U115bar (
    .O(ybar[227]),
    .I0(abar[14]),
    .I1(bbar[3])
  );
  //AND U116
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U116 (
    .O(y[226]),
    .I0(a[14]),
    .I1(b[2])
  );
  //OR U116bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U116bar (
    .O(ybar[226]),
    .I0(abar[14]),
    .I1(bbar[2])
  );
  //AND U117
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U117 (
    .O(y[225]),
    .I0(a[14]),
    .I1(b[1])
  );
  //OR U117bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U117bar (
    .O(ybar[225]),
    .I0(abar[14]),
    .I1(bbar[1])
  );
  //AND U118
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U118 (
    .O(y[224]),
    .I0(a[14]),
    .I1(b[0])
  );
  //OR U118bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U118bar (
    .O(ybar[224]),
    .I0(abar[14]),
    .I1(bbar[0])
  );
  //AND U119
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U119 (
    .O(y[223]),
    .I0(a[13]),
    .I1(b[15])
  );
  //OR U119bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U119bar (
    .O(ybar[223]),
    .I0(abar[13]),
    .I1(bbar[15])
  );
  //AND U120
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U120 (
    .O(y[222]),
    .I0(a[13]),
    .I1(b[14])
  );
  //OR U120bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U120bar (
    .O(ybar[222]),
    .I0(abar[13]),
    .I1(bbar[14])
  );
  //AND U121
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U121 (
    .O(y[221]),
    .I0(a[13]),
    .I1(b[13])
  );
  //OR U121bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U121bar (
    .O(ybar[221]),
    .I0(abar[13]),
    .I1(bbar[13])
  );
  //AND U122
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U122 (
    .O(y[220]),
    .I0(a[13]),
    .I1(b[12])
  );
  //OR U122bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U122bar (
    .O(ybar[220]),
    .I0(abar[13]),
    .I1(bbar[12])
  );
  //AND U123
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U123 (
    .O(y[21]),
    .I0(a[1]),
    .I1(b[5])
  );
  //OR U123bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U123bar (
    .O(ybar[21]),
    .I0(abar[1]),
    .I1(bbar[5])
  );
  //AND U124
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U124 (
    .O(y[219]),
    .I0(a[13]),
    .I1(b[11])
  );
  //OR U124bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U124bar (
    .O(ybar[219]),
    .I0(abar[13]),
    .I1(bbar[11])
  );
  //AND U125
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U125 (
    .O(y[218]),
    .I0(a[13]),
    .I1(b[10])
  );
  //OR U125bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U125bar (
    .O(ybar[218]),
    .I0(abar[13]),
    .I1(bbar[10])
  );
  //AND U126
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U126 (
    .O(y[217]),
    .I0(a[13]),
    .I1(b[9])
  );
  //OR U126bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U126bar (
    .O(ybar[217]),
    .I0(abar[13]),
    .I1(bbar[9])
  );
  //AND U127
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U127 (
    .O(y[216]),
    .I0(a[13]),
    .I1(b[8])
  );
  //OR U127bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U127bar (
    .O(ybar[216]),
    .I0(abar[13]),
    .I1(bbar[8])
  );
  //AND U128
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U128 (
    .O(y[215]),
    .I0(a[13]),
    .I1(b[7])
  );
  //OR U128bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U128bar (
    .O(ybar[215]),
    .I0(abar[13]),
    .I1(bbar[7])
  );
  //AND U129
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U129 (
    .O(y[214]),
    .I0(a[13]),
    .I1(b[6])
  );
  //OR U129bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U129bar (
    .O(ybar[214]),
    .I0(abar[13]),
    .I1(bbar[6])
  );
  //AND U130
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U130 (
    .O(y[213]),
    .I0(a[13]),
    .I1(b[5])
  );
  //OR U130bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U130bar (
    .O(ybar[213]),
    .I0(abar[13]),
    .I1(bbar[5])
  );
  //AND U131
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U131 (
    .O(y[212]),
    .I0(a[13]),
    .I1(b[4])
  );
  //OR U131bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U131bar (
    .O(ybar[212]),
    .I0(abar[13]),
    .I1(bbar[4])
  );
  //AND U132
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U132 (
    .O(y[211]),
    .I0(a[13]),
    .I1(b[3])
  );
  //OR U132bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U132bar (
    .O(ybar[211]),
    .I0(abar[13]),
    .I1(bbar[3])
  );
  //AND U133
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U133 (
    .O(y[210]),
    .I0(a[13]),
    .I1(b[2])
  );
  //OR U133bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U133bar (
    .O(ybar[210]),
    .I0(abar[13]),
    .I1(bbar[2])
  );
  //AND U134
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U134 (
    .O(y[20]),
    .I0(a[1]),
    .I1(b[4])
  );
  //OR U134bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U134bar (
    .O(ybar[20]),
    .I0(abar[1]),
    .I1(bbar[4])
  );
  //AND U135
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U135 (
    .O(y[209]),
    .I0(a[13]),
    .I1(b[1])
  );
  //OR U135bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U135bar (
    .O(ybar[209]),
    .I0(abar[13]),
    .I1(bbar[1])
  );
  //AND U136
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U136 (
    .O(y[208]),
    .I0(a[13]),
    .I1(b[0])
  );
  //OR U136bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U136bar (
    .O(ybar[208]),
    .I0(abar[13]),
    .I1(bbar[0])
  );
  //AND U137
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U137 (
    .O(y[207]),
    .I0(a[12]),
    .I1(b[15])
  );
  //OR U137bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U137bar (
    .O(ybar[207]),
    .I0(abar[12]),
    .I1(bbar[15])
  );
  //AND U138
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U138 (
    .O(y[206]),
    .I0(a[12]),
    .I1(b[14])
  );
  //OR U138bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U138bar (
    .O(ybar[206]),
    .I0(abar[12]),
    .I1(bbar[14])
  );
  //AND U139
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U139 (
    .O(y[205]),
    .I0(a[12]),
    .I1(b[13])
  );
  //OR U139bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U139bar (
    .O(ybar[205]),
    .I0(abar[12]),
    .I1(bbar[13])
  );
  //AND U140
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U140 (
    .O(y[204]),
    .I0(a[12]),
    .I1(b[12])
  );
  //OR U140bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U140bar (
    .O(ybar[204]),
    .I0(abar[12]),
    .I1(bbar[12])
  );
  //AND U141
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U141 (
    .O(y[203]),
    .I0(a[12]),
    .I1(b[11])
  );
  //OR U141bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U141bar (
    .O(ybar[203]),
    .I0(abar[12]),
    .I1(bbar[11])
  );
  //AND U142
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U142 (
    .O(y[202]),
    .I0(a[12]),
    .I1(b[10])
  );
  //OR U142bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U142bar (
    .O(ybar[202]),
    .I0(abar[12]),
    .I1(bbar[10])
  );
  //AND U143
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U143 (
    .O(y[201]),
    .I0(a[12]),
    .I1(b[9])
  );
  //OR U143bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U143bar (
    .O(ybar[201]),
    .I0(abar[12]),
    .I1(bbar[9])
  );
  //AND U144
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U144 (
    .O(y[200]),
    .I0(a[12]),
    .I1(b[8])
  );
  //OR U144bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U144bar (
    .O(ybar[200]),
    .I0(abar[12]),
    .I1(bbar[8])
  );
  //AND U145
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U145 (
    .O(y[1]),
    .I0(b[1]),
    .I1(a[0])
  );
  //OR U145bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U145bar (
    .O(ybar[1]),
    .I0(bbar[1]),
    .I1(abar[0])
  );
  //AND U146
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U146 (
    .O(y[19]),
    .I0(a[1]),
    .I1(b[3])
  );
  //OR U146bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U146bar (
    .O(ybar[19]),
    .I0(abar[1]),
    .I1(bbar[3])
  );
  //AND U147
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U147 (
    .O(y[199]),
    .I0(a[12]),
    .I1(b[7])
  );
  //OR U147bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U147bar (
    .O(ybar[199]),
    .I0(abar[12]),
    .I1(bbar[7])
  );
  //AND U148
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U148 (
    .O(y[198]),
    .I0(a[12]),
    .I1(b[6])
  );
  //OR U148bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U148bar (
    .O(ybar[198]),
    .I0(abar[12]),
    .I1(bbar[6])
  );
  //AND U149
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U149 (
    .O(y[197]),
    .I0(a[12]),
    .I1(b[5])
  );
  //OR U149bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U149bar (
    .O(ybar[197]),
    .I0(abar[12]),
    .I1(bbar[5])
  );
  //AND U150
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U150 (
    .O(y[196]),
    .I0(a[12]),
    .I1(b[4])
  );
  //OR U150bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U150bar (
    .O(ybar[196]),
    .I0(abar[12]),
    .I1(bbar[4])
  );
  //AND U151
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U151 (
    .O(y[195]),
    .I0(a[12]),
    .I1(b[3])
  );
  //OR U151bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U151bar (
    .O(ybar[195]),
    .I0(abar[12]),
    .I1(bbar[3])
  );
  //AND U152
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U152 (
    .O(y[194]),
    .I0(a[12]),
    .I1(b[2])
  );
  //OR U152bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U152bar (
    .O(ybar[194]),
    .I0(abar[12]),
    .I1(bbar[2])
  );
  //AND U153
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U153 (
    .O(y[193]),
    .I0(a[12]),
    .I1(b[1])
  );
  //OR U153bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U153bar (
    .O(ybar[193]),
    .I0(abar[12]),
    .I1(bbar[1])
  );
  //AND U154
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U154 (
    .O(y[192]),
    .I0(a[12]),
    .I1(b[0])
  );
  //OR U154bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U154bar (
    .O(ybar[192]),
    .I0(abar[12]),
    .I1(bbar[0])
  );
  //AND U155
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U155 (
    .O(y[191]),
    .I0(a[11]),
    .I1(b[15])
  );
  //OR U155bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U155bar (
    .O(ybar[191]),
    .I0(abar[11]),
    .I1(bbar[15])
  );
  //AND U156
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U156 (
    .O(y[190]),
    .I0(a[11]),
    .I1(b[14])
  );
  //OR U156bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U156bar (
    .O(ybar[190]),
    .I0(abar[11]),
    .I1(bbar[14])
  );
  //AND U157
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U157 (
    .O(y[18]),
    .I0(a[1]),
    .I1(b[2])
  );
  //OR U157bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U157bar (
    .O(ybar[18]),
    .I0(abar[1]),
    .I1(bbar[2])
  );
  //AND U158
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U158 (
    .O(y[189]),
    .I0(a[11]),
    .I1(b[13])
  );
  //OR U158bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U158bar (
    .O(ybar[189]),
    .I0(abar[11]),
    .I1(bbar[13])
  );
  //AND U159
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U159 (
    .O(y[188]),
    .I0(a[11]),
    .I1(b[12])
  );
  //OR U159bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U159bar (
    .O(ybar[188]),
    .I0(abar[11]),
    .I1(bbar[12])
  );
  //AND U160
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U160 (
    .O(y[187]),
    .I0(a[11]),
    .I1(b[11])
  );
  //OR U160bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U160bar (
    .O(ybar[187]),
    .I0(abar[11]),
    .I1(bbar[11])
  );
  //AND U161
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U161 (
    .O(y[186]),
    .I0(a[11]),
    .I1(b[10])
  );
  //OR U161bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U161bar (
    .O(ybar[186]),
    .I0(abar[11]),
    .I1(bbar[10])
  );
  //AND U162
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U162 (
    .O(y[185]),
    .I0(a[11]),
    .I1(b[9])
  );
  //OR U162bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U162bar (
    .O(ybar[185]),
    .I0(abar[11]),
    .I1(bbar[9])
  );
  //AND U163
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U163 (
    .O(y[184]),
    .I0(a[11]),
    .I1(b[8])
  );
  //OR U163bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U163bar (
    .O(ybar[184]),
    .I0(abar[11]),
    .I1(bbar[8])
  );
  //AND U164
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U164 (
    .O(y[183]),
    .I0(a[11]),
    .I1(b[7])
  );
  //OR U164bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U164bar (
    .O(ybar[183]),
    .I0(abar[11]),
    .I1(bbar[7])
  );
  //AND U165
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U165 (
    .O(y[182]),
    .I0(a[11]),
    .I1(b[6])
  );
  //OR U165bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U165bar (
    .O(ybar[182]),
    .I0(abar[11]),
    .I1(bbar[6])
  );
  //AND U166
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U166 (
    .O(y[181]),
    .I0(a[11]),
    .I1(b[5])
  );
  //OR U166bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U166bar (
    .O(ybar[181]),
    .I0(abar[11]),
    .I1(bbar[5])
  );
  //AND U167
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U167 (
    .O(y[180]),
    .I0(a[11]),
    .I1(b[4])
  );
  //OR U167bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U167bar (
    .O(ybar[180]),
    .I0(abar[11]),
    .I1(bbar[4])
  );
  //AND U168
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U168 (
    .O(y[17]),
    .I0(a[1]),
    .I1(b[1])
  );
  //OR U168bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U168bar (
    .O(ybar[17]),
    .I0(abar[1]),
    .I1(bbar[1])
  );
  //AND U169
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U169 (
    .O(y[179]),
    .I0(a[11]),
    .I1(b[3])
  );
  //OR U169bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U169bar (
    .O(ybar[179]),
    .I0(abar[11]),
    .I1(bbar[3])
  );
  //AND U170
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U170 (
    .O(y[178]),
    .I0(a[11]),
    .I1(b[2])
  );
  //OR U170bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U170bar (
    .O(ybar[178]),
    .I0(abar[11]),
    .I1(bbar[2])
  );
  //AND U171
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U171 (
    .O(y[177]),
    .I0(a[11]),
    .I1(b[1])
  );
  //OR U171bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U171bar (
    .O(ybar[177]),
    .I0(abar[11]),
    .I1(bbar[1])
  );
  //AND U172
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U172 (
    .O(y[176]),
    .I0(a[11]),
    .I1(b[0])
  );
  //OR U172bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U172bar (
    .O(ybar[176]),
    .I0(abar[11]),
    .I1(bbar[0])
  );
  //AND U173
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U173 (
    .O(y[175]),
    .I0(a[10]),
    .I1(b[15])
  );
  //OR U173bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U173bar (
    .O(ybar[175]),
    .I0(abar[10]),
    .I1(bbar[15])
  );
  //AND U174
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U174 (
    .O(y[174]),
    .I0(a[10]),
    .I1(b[14])
  );
  //OR U174bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U174bar (
    .O(ybar[174]),
    .I0(abar[10]),
    .I1(bbar[14])
  );
  //AND U175
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U175 (
    .O(y[173]),
    .I0(a[10]),
    .I1(b[13])
  );
  //OR U175bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U175bar (
    .O(ybar[173]),
    .I0(abar[10]),
    .I1(bbar[13])
  );
  //AND U176
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U176 (
    .O(y[172]),
    .I0(a[10]),
    .I1(b[12])
  );
  //OR U176bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U176bar (
    .O(ybar[172]),
    .I0(abar[10]),
    .I1(bbar[12])
  );
  //AND U177
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U177 (
    .O(y[171]),
    .I0(a[10]),
    .I1(b[11])
  );
  //OR U177bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U177bar (
    .O(ybar[171]),
    .I0(abar[10]),
    .I1(bbar[11])
  );
  //AND U178
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U178 (
    .O(y[170]),
    .I0(a[10]),
    .I1(b[10])
  );
  //OR U178bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U178bar (
    .O(ybar[170]),
    .I0(abar[10]),
    .I1(bbar[10])
  );
  //AND U179
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U179 (
    .O(y[16]),
    .I0(a[1]),
    .I1(b[0])
  );
  //OR U179bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U179bar (
    .O(ybar[16]),
    .I0(abar[1]),
    .I1(bbar[0])
  );
  //AND U180
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U180 (
    .O(y[169]),
    .I0(a[10]),
    .I1(b[9])
  );
  //OR U180bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U180bar (
    .O(ybar[169]),
    .I0(abar[10]),
    .I1(bbar[9])
  );
  //AND U181
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U181 (
    .O(y[168]),
    .I0(a[10]),
    .I1(b[8])
  );
  //OR U181bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U181bar (
    .O(ybar[168]),
    .I0(abar[10]),
    .I1(bbar[8])
  );
  //AND U182
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U182 (
    .O(y[167]),
    .I0(a[10]),
    .I1(b[7])
  );
  //OR U182bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U182bar (
    .O(ybar[167]),
    .I0(abar[10]),
    .I1(bbar[7])
  );
  //AND U183
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U183 (
    .O(y[166]),
    .I0(a[10]),
    .I1(b[6])
  );
  //OR U183bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U183bar (
    .O(ybar[166]),
    .I0(abar[10]),
    .I1(bbar[6])
  );
  //AND U184
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U184 (
    .O(y[165]),
    .I0(a[10]),
    .I1(b[5])
  );
  //OR U184bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U184bar (
    .O(ybar[165]),
    .I0(abar[10]),
    .I1(bbar[5])
  );
  //AND U185
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U185 (
    .O(y[164]),
    .I0(a[10]),
    .I1(b[4])
  );
  //OR U185bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U185bar (
    .O(ybar[164]),
    .I0(abar[10]),
    .I1(bbar[4])
  );
  //AND U186
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U186 (
    .O(y[163]),
    .I0(a[10]),
    .I1(b[3])
  );
  //OR U186bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U186bar (
    .O(ybar[163]),
    .I0(abar[10]),
    .I1(bbar[3])
  );
  //AND U187
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U187 (
    .O(y[162]),
    .I0(a[10]),
    .I1(b[2])
  );
  //OR U187bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U187bar (
    .O(ybar[162]),
    .I0(abar[10]),
    .I1(bbar[2])
  );
  //AND U188
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U188 (
    .O(y[161]),
    .I0(a[10]),
    .I1(b[1])
  );
  //OR U188bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U188bar (
    .O(ybar[161]),
    .I0(abar[10]),
    .I1(bbar[1])
  );
  //AND U189
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U189 (
    .O(y[160]),
    .I0(a[10]),
    .I1(b[0])
  );
  //OR U189bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U189bar (
    .O(ybar[160]),
    .I0(abar[10]),
    .I1(bbar[0])
  );
  //AND U190
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U190 (
    .O(y[15]),
    .I0(b[15]),
    .I1(a[0])
  );
  //OR U190bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U190bar (
    .O(ybar[15]),
    .I0(bbar[15]),
    .I1(abar[0])
  );
  //AND U191
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U191 (
    .O(y[159]),
    .I0(a[9]),
    .I1(b[15])
  );
  //OR U191bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U191bar (
    .O(ybar[159]),
    .I0(abar[9]),
    .I1(bbar[15])
  );
  //AND U192
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U192 (
    .O(y[158]),
    .I0(a[9]),
    .I1(b[14])
  );
  //OR U192bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U192bar (
    .O(ybar[158]),
    .I0(abar[9]),
    .I1(bbar[14])
  );
  //AND U193
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U193 (
    .O(y[157]),
    .I0(a[9]),
    .I1(b[13])
  );
  //OR U193bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U193bar (
    .O(ybar[157]),
    .I0(abar[9]),
    .I1(bbar[13])
  );
  //AND U194
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U194 (
    .O(y[156]),
    .I0(a[9]),
    .I1(b[12])
  );
  //OR U194bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U194bar (
    .O(ybar[156]),
    .I0(abar[9]),
    .I1(bbar[12])
  );
  //AND U195
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U195 (
    .O(y[155]),
    .I0(a[9]),
    .I1(b[11])
  );
  //OR U195bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U195bar (
    .O(ybar[155]),
    .I0(abar[9]),
    .I1(bbar[11])
  );
  //AND U196
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U196 (
    .O(y[154]),
    .I0(a[9]),
    .I1(b[10])
  );
  //OR U196bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U196bar (
    .O(ybar[154]),
    .I0(abar[9]),
    .I1(bbar[10])
  );
  //AND U197
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U197 (
    .O(y[153]),
    .I0(a[9]),
    .I1(b[9])
  );
  //OR U197bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U197bar (
    .O(ybar[153]),
    .I0(abar[9]),
    .I1(bbar[9])
  );
  //AND U198
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U198 (
    .O(y[152]),
    .I0(a[9]),
    .I1(b[8])
  );
  //OR U198bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U198bar (
    .O(ybar[152]),
    .I0(abar[9]),
    .I1(bbar[8])
  );
  //AND U199
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U199 (
    .O(y[151]),
    .I0(a[9]),
    .I1(b[7])
  );
  //OR U199bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U199bar (
    .O(ybar[151]),
    .I0(abar[9]),
    .I1(bbar[7])
  );
  //AND U200
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U200 (
    .O(y[150]),
    .I0(a[9]),
    .I1(b[6])
  );
  //OR U200bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U200bar (
    .O(ybar[150]),
    .I0(abar[9]),
    .I1(bbar[6])
  );
  //AND U201
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U201 (
    .O(y[14]),
    .I0(b[14]),
    .I1(a[0])
  );
  //OR U201bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U201bar (
    .O(ybar[14]),
    .I0(bbar[14]),
    .I1(abar[0])
  );
  //AND U202
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U202 (
    .O(y[149]),
    .I0(a[9]),
    .I1(b[5])
  );
  //OR U202bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U202bar (
    .O(ybar[149]),
    .I0(abar[9]),
    .I1(bbar[5])
  );
  //AND U203
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U203 (
    .O(y[148]),
    .I0(a[9]),
    .I1(b[4])
  );
  //OR U203bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U203bar (
    .O(ybar[148]),
    .I0(abar[9]),
    .I1(bbar[4])
  );
  //AND U204
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U204 (
    .O(y[147]),
    .I0(a[9]),
    .I1(b[3])
  );
  //OR U204bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U204bar (
    .O(ybar[147]),
    .I0(abar[9]),
    .I1(bbar[3])
  );
  //AND U205
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U205 (
    .O(y[146]),
    .I0(a[9]),
    .I1(b[2])
  );
  //OR U205bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U205bar (
    .O(ybar[146]),
    .I0(abar[9]),
    .I1(bbar[2])
  );
  //AND U206
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U206 (
    .O(y[145]),
    .I0(a[9]),
    .I1(b[1])
  );
  //OR U206bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U206bar (
    .O(ybar[145]),
    .I0(abar[9]),
    .I1(bbar[1])
  );
  //AND U207
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U207 (
    .O(y[144]),
    .I0(a[9]),
    .I1(b[0])
  );
  //OR U207bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U207bar (
    .O(ybar[144]),
    .I0(abar[9]),
    .I1(bbar[0])
  );
  //AND U208
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U208 (
    .O(y[143]),
    .I0(a[8]),
    .I1(b[15])
  );
  //OR U208bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U208bar (
    .O(ybar[143]),
    .I0(abar[8]),
    .I1(bbar[15])
  );
  //AND U209
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U209 (
    .O(y[142]),
    .I0(a[8]),
    .I1(b[14])
  );
  //OR U209bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U209bar (
    .O(ybar[142]),
    .I0(abar[8]),
    .I1(bbar[14])
  );
  //AND U210
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U210 (
    .O(y[141]),
    .I0(a[8]),
    .I1(b[13])
  );
  //OR U210bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U210bar (
    .O(ybar[141]),
    .I0(abar[8]),
    .I1(bbar[13])
  );
  //AND U211
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U211 (
    .O(y[140]),
    .I0(a[8]),
    .I1(b[12])
  );
  //OR U211bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U211bar (
    .O(ybar[140]),
    .I0(abar[8]),
    .I1(bbar[12])
  );
  //AND U212
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U212 (
    .O(y[13]),
    .I0(b[13]),
    .I1(a[0])
  );
  //OR U212bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U212bar (
    .O(ybar[13]),
    .I0(bbar[13]),
    .I1(abar[0])
  );
  //AND U213
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U213 (
    .O(y[139]),
    .I0(a[8]),
    .I1(b[11])
  );
  //OR U213bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U213bar (
    .O(ybar[139]),
    .I0(abar[8]),
    .I1(bbar[11])
  );
  //AND U214
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U214 (
    .O(y[138]),
    .I0(a[8]),
    .I1(b[10])
  );
  //OR U214bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U214bar (
    .O(ybar[138]),
    .I0(abar[8]),
    .I1(bbar[10])
  );
  //AND U215
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U215 (
    .O(y[137]),
    .I0(a[8]),
    .I1(b[9])
  );
  //OR U215bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U215bar (
    .O(ybar[137]),
    .I0(abar[8]),
    .I1(bbar[9])
  );
  //AND U216
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U216 (
    .O(y[136]),
    .I0(a[8]),
    .I1(b[8])
  );
  //OR U216bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U216bar (
    .O(ybar[136]),
    .I0(abar[8]),
    .I1(bbar[8])
  );
  //AND U217
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U217 (
    .O(y[135]),
    .I0(a[8]),
    .I1(b[7])
  );
  //OR U217bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U217bar (
    .O(ybar[135]),
    .I0(abar[8]),
    .I1(bbar[7])
  );
  //AND U218
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U218 (
    .O(y[134]),
    .I0(a[8]),
    .I1(b[6])
  );
  //OR U218bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U218bar (
    .O(ybar[134]),
    .I0(abar[8]),
    .I1(bbar[6])
  );
  //AND U219
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U219 (
    .O(y[133]),
    .I0(a[8]),
    .I1(b[5])
  );
  //OR U219bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U219bar (
    .O(ybar[133]),
    .I0(abar[8]),
    .I1(bbar[5])
  );
  //AND U220
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U220 (
    .O(y[132]),
    .I0(a[8]),
    .I1(b[4])
  );
  //OR U220bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U220bar (
    .O(ybar[132]),
    .I0(abar[8]),
    .I1(bbar[4])
  );
  //AND U221
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U221 (
    .O(y[131]),
    .I0(a[8]),
    .I1(b[3])
  );
  //OR U221bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U221bar (
    .O(ybar[131]),
    .I0(abar[8]),
    .I1(bbar[3])
  );
  //AND U222
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U222 (
    .O(y[130]),
    .I0(a[8]),
    .I1(b[2])
  );
  //OR U222bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U222bar (
    .O(ybar[130]),
    .I0(abar[8]),
    .I1(bbar[2])
  );
  //AND U223
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U223 (
    .O(y[12]),
    .I0(b[12]),
    .I1(a[0])
  );
  //OR U223bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U223bar (
    .O(ybar[12]),
    .I0(bbar[12]),
    .I1(abar[0])
  );
  //AND U224
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U224 (
    .O(y[129]),
    .I0(a[8]),
    .I1(b[1])
  );
  //OR U224bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U224bar (
    .O(ybar[129]),
    .I0(abar[8]),
    .I1(bbar[1])
  );
  //AND U225
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U225 (
    .O(y[128]),
    .I0(a[8]),
    .I1(b[0])
  );
  //OR U225bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U225bar (
    .O(ybar[128]),
    .I0(abar[8]),
    .I1(bbar[0])
  );
  //AND U226
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U226 (
    .O(y[127]),
    .I0(a[7]),
    .I1(b[15])
  );
  //OR U226bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U226bar (
    .O(ybar[127]),
    .I0(abar[7]),
    .I1(bbar[15])
  );
  //AND U227
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U227 (
    .O(y[126]),
    .I0(a[7]),
    .I1(b[14])
  );
  //OR U227bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U227bar (
    .O(ybar[126]),
    .I0(abar[7]),
    .I1(bbar[14])
  );
  //AND U228
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U228 (
    .O(y[125]),
    .I0(a[7]),
    .I1(b[13])
  );
  //OR U228bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U228bar (
    .O(ybar[125]),
    .I0(abar[7]),
    .I1(bbar[13])
  );
  //AND U229
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U229 (
    .O(y[124]),
    .I0(a[7]),
    .I1(b[12])
  );
  //OR U229bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U229bar (
    .O(ybar[124]),
    .I0(abar[7]),
    .I1(bbar[12])
  );
  //AND U230
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U230 (
    .O(y[123]),
    .I0(a[7]),
    .I1(b[11])
  );
  //OR U230bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U230bar (
    .O(ybar[123]),
    .I0(abar[7]),
    .I1(bbar[11])
  );
  //AND U231
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U231 (
    .O(y[122]),
    .I0(a[7]),
    .I1(b[10])
  );
  //OR U231bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U231bar (
    .O(ybar[122]),
    .I0(abar[7]),
    .I1(bbar[10])
  );
  //AND U232
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U232 (
    .O(y[121]),
    .I0(a[7]),
    .I1(b[9])
  );
  //OR U232bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U232bar (
    .O(ybar[121]),
    .I0(abar[7]),
    .I1(bbar[9])
  );
  //AND U233
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U233 (
    .O(y[120]),
    .I0(a[7]),
    .I1(b[8])
  );
  //OR U233bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U233bar (
    .O(ybar[120]),
    .I0(abar[7]),
    .I1(bbar[8])
  );
  //AND U234
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U234 (
    .O(y[11]),
    .I0(b[11]),
    .I1(a[0])
  );
  //OR U234bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U234bar (
    .O(ybar[11]),
    .I0(bbar[11]),
    .I1(abar[0])
  );
  //AND U235
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U235 (
    .O(y[119]),
    .I0(a[7]),
    .I1(b[7])
  );
  //OR U235bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U235bar (
    .O(ybar[119]),
    .I0(abar[7]),
    .I1(bbar[7])
  );
  //AND U236
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U236 (
    .O(y[118]),
    .I0(a[7]),
    .I1(b[6])
  );
  //OR U236bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U236bar (
    .O(ybar[118]),
    .I0(abar[7]),
    .I1(bbar[6])
  );
  //AND U237
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U237 (
    .O(y[117]),
    .I0(a[7]),
    .I1(b[5])
  );
  //OR U237bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U237bar (
    .O(ybar[117]),
    .I0(abar[7]),
    .I1(bbar[5])
  );
  //AND U238
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U238 (
    .O(y[116]),
    .I0(a[7]),
    .I1(b[4])
  );
  //OR U238bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U238bar (
    .O(ybar[116]),
    .I0(abar[7]),
    .I1(bbar[4])
  );
  //AND U239
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U239 (
    .O(y[115]),
    .I0(a[7]),
    .I1(b[3])
  );
  //OR U239bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U239bar (
    .O(ybar[115]),
    .I0(abar[7]),
    .I1(bbar[3])
  );
  //AND U240
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U240 (
    .O(y[114]),
    .I0(a[7]),
    .I1(b[2])
  );
  //OR U240bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U240bar (
    .O(ybar[114]),
    .I0(abar[7]),
    .I1(bbar[2])
  );
  //AND U241
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U241 (
    .O(y[113]),
    .I0(a[7]),
    .I1(b[1])
  );
  //OR U241bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U241bar (
    .O(ybar[113]),
    .I0(abar[7]),
    .I1(bbar[1])
  );
  //AND U242
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U242 (
    .O(y[112]),
    .I0(a[7]),
    .I1(b[0])
  );
  //OR U242bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U242bar (
    .O(ybar[112]),
    .I0(abar[7]),
    .I1(bbar[0])
  );
  //AND U243
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U243 (
    .O(y[111]),
    .I0(b[15]),
    .I1(a[6])
  );
  //OR U243bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U243bar (
    .O(ybar[111]),
    .I0(bbar[15]),
    .I1(abar[6])
  );
  //AND U244
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U244 (
    .O(y[110]),
    .I0(b[14]),
    .I1(a[6])
  );
  //OR U244bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U244bar (
    .O(ybar[110]),
    .I0(bbar[14]),
    .I1(abar[6])
  );
  //AND U245
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U245 (
    .O(y[10]),
    .I0(b[10]),
    .I1(a[0])
  );
  //OR U245bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U245bar (
    .O(ybar[10]),
    .I0(bbar[10]),
    .I1(abar[0])
  );
  //AND U246
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U246 (
    .O(y[109]),
    .I0(b[13]),
    .I1(a[6])
  );
  //OR U246bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U246bar (
    .O(ybar[109]),
    .I0(bbar[13]),
    .I1(abar[6])
  );
  //AND U247
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U247 (
    .O(y[108]),
    .I0(b[12]),
    .I1(a[6])
  );
  //OR U247bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U247bar (
    .O(ybar[108]),
    .I0(bbar[12]),
    .I1(abar[6])
  );
  //AND U248
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U248 (
    .O(y[107]),
    .I0(b[11]),
    .I1(a[6])
  );
  //OR U248bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U248bar (
    .O(ybar[107]),
    .I0(bbar[11]),
    .I1(abar[6])
  );
  //AND U249
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U249 (
    .O(y[106]),
    .I0(b[10]),
    .I1(a[6])
  );
  //OR U249bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U249bar (
    .O(ybar[106]),
    .I0(bbar[10]),
    .I1(abar[6])
  );
  //AND U250
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U250 (
    .O(y[105]),
    .I0(a[6]),
    .I1(b[9])
  );
  //OR U250bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U250bar (
    .O(ybar[105]),
    .I0(abar[6]),
    .I1(bbar[9])
  );
  //AND U251
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U251 (
    .O(y[104]),
    .I0(b[8]),
    .I1(a[6])
  );
  //OR U251bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U251bar (
    .O(ybar[104]),
    .I0(bbar[8]),
    .I1(abar[6])
  );
  //AND U252
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U252 (
    .O(y[103]),
    .I0(b[7]),
    .I1(a[6])
  );
  //OR U252bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U252bar (
    .O(ybar[103]),
    .I0(bbar[7]),
    .I1(abar[6])
  );
  //AND U253
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U253 (
    .O(y[102]),
    .I0(b[6]),
    .I1(a[6])
  );
  //OR U253bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U253bar (
    .O(ybar[102]),
    .I0(bbar[6]),
    .I1(abar[6])
  );
  //AND U254
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U254 (
    .O(y[101]),
    .I0(b[5]),
    .I1(a[6])
  );
  //OR U254bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U254bar (
    .O(ybar[101]),
    .I0(bbar[5]),
    .I1(abar[6])
  );
  //AND U255
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U255 (
    .O(y[100]),
    .I0(b[4]),
    .I1(a[6])
  );
  //OR U255bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U255bar (
    .O(ybar[100]),
    .I0(bbar[4]),
    .I1(abar[6])
  );
  //AND U256
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U256 (
    .O(y[0]),
    .I0(b[0]),
    .I1(a[0])
  );
  //OR U256bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U256bar (
    .O(ybar[0]),
    .I0(bbar[0]),
    .I1(abar[0])
  );
endmodule

module decode_2 ( in, out );

  input wire [7:0] in;
//input_done

  output wire [255:0] out;
//output_done

  wire [15:0] level1;
  wire [31:0] level2;
//wire_done

  CD2_8 cd_l1_1 ( .a(in[1]), .b(in[0]), .y(level1[3:0]) );
  CD2_7 cd_l1_2 ( .a(in[3]), .b(in[2]), .y(level1[7:4]) );
  CD2_6 cd_l1_3 ( .a(in[5]), .b(in[4]), .y(level1[11:8]) );
  CD2_5 cd_l1_4 ( .a(in[7]), .b(in[6]), .y(level1[15:12]) );
  CD4_4 cd_l2_1 ( .a(level1[7:4]), .b(level1[3:0]), .y(level2[15:0]) );
  CD4_3 cd_l2_2 ( .a(level1[15:12]), .b(level1[11:8]), .y(level2[31:16]) );
  CD16_2 cd_l3 ( .a(level2[31:16]), .b(level2[15:0]), .y(out) );
endmodule

module encode_2 ( in, out );

  input wire [255:0] in;
  wire [255:0] inbar;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
  assign inbar[8] = ~in[8];
  assign inbar[9] = ~in[9];
  assign inbar[10] = ~in[10];
  assign inbar[11] = ~in[11];
  assign inbar[12] = ~in[12];
  assign inbar[13] = ~in[13];
  assign inbar[14] = ~in[14];
  assign inbar[15] = ~in[15];
  assign inbar[16] = ~in[16];
  assign inbar[17] = ~in[17];
  assign inbar[18] = ~in[18];
  assign inbar[19] = ~in[19];
  assign inbar[20] = ~in[20];
  assign inbar[21] = ~in[21];
  assign inbar[22] = ~in[22];
  assign inbar[23] = ~in[23];
  assign inbar[24] = ~in[24];
  assign inbar[25] = ~in[25];
  assign inbar[26] = ~in[26];
  assign inbar[27] = ~in[27];
  assign inbar[28] = ~in[28];
  assign inbar[29] = ~in[29];
  assign inbar[30] = ~in[30];
  assign inbar[31] = ~in[31];
  assign inbar[32] = ~in[32];
  assign inbar[33] = ~in[33];
  assign inbar[34] = ~in[34];
  assign inbar[35] = ~in[35];
  assign inbar[36] = ~in[36];
  assign inbar[37] = ~in[37];
  assign inbar[38] = ~in[38];
  assign inbar[39] = ~in[39];
  assign inbar[40] = ~in[40];
  assign inbar[41] = ~in[41];
  assign inbar[42] = ~in[42];
  assign inbar[43] = ~in[43];
  assign inbar[44] = ~in[44];
  assign inbar[45] = ~in[45];
  assign inbar[46] = ~in[46];
  assign inbar[47] = ~in[47];
  assign inbar[48] = ~in[48];
  assign inbar[49] = ~in[49];
  assign inbar[50] = ~in[50];
  assign inbar[51] = ~in[51];
  assign inbar[52] = ~in[52];
  assign inbar[53] = ~in[53];
  assign inbar[54] = ~in[54];
  assign inbar[55] = ~in[55];
  assign inbar[56] = ~in[56];
  assign inbar[57] = ~in[57];
  assign inbar[58] = ~in[58];
  assign inbar[59] = ~in[59];
  assign inbar[60] = ~in[60];
  assign inbar[61] = ~in[61];
  assign inbar[62] = ~in[62];
  assign inbar[63] = ~in[63];
  assign inbar[64] = ~in[64];
  assign inbar[65] = ~in[65];
  assign inbar[66] = ~in[66];
  assign inbar[67] = ~in[67];
  assign inbar[68] = ~in[68];
  assign inbar[69] = ~in[69];
  assign inbar[70] = ~in[70];
  assign inbar[71] = ~in[71];
  assign inbar[72] = ~in[72];
  assign inbar[73] = ~in[73];
  assign inbar[74] = ~in[74];
  assign inbar[75] = ~in[75];
  assign inbar[76] = ~in[76];
  assign inbar[77] = ~in[77];
  assign inbar[78] = ~in[78];
  assign inbar[79] = ~in[79];
  assign inbar[80] = ~in[80];
  assign inbar[81] = ~in[81];
  assign inbar[82] = ~in[82];
  assign inbar[83] = ~in[83];
  assign inbar[84] = ~in[84];
  assign inbar[85] = ~in[85];
  assign inbar[86] = ~in[86];
  assign inbar[87] = ~in[87];
  assign inbar[88] = ~in[88];
  assign inbar[89] = ~in[89];
  assign inbar[90] = ~in[90];
  assign inbar[91] = ~in[91];
  assign inbar[92] = ~in[92];
  assign inbar[93] = ~in[93];
  assign inbar[94] = ~in[94];
  assign inbar[95] = ~in[95];
  assign inbar[96] = ~in[96];
  assign inbar[97] = ~in[97];
  assign inbar[98] = ~in[98];
  assign inbar[99] = ~in[99];
  assign inbar[100] = ~in[100];
  assign inbar[101] = ~in[101];
  assign inbar[102] = ~in[102];
  assign inbar[103] = ~in[103];
  assign inbar[104] = ~in[104];
  assign inbar[105] = ~in[105];
  assign inbar[106] = ~in[106];
  assign inbar[107] = ~in[107];
  assign inbar[108] = ~in[108];
  assign inbar[109] = ~in[109];
  assign inbar[110] = ~in[110];
  assign inbar[111] = ~in[111];
  assign inbar[112] = ~in[112];
  assign inbar[113] = ~in[113];
  assign inbar[114] = ~in[114];
  assign inbar[115] = ~in[115];
  assign inbar[116] = ~in[116];
  assign inbar[117] = ~in[117];
  assign inbar[118] = ~in[118];
  assign inbar[119] = ~in[119];
  assign inbar[120] = ~in[120];
  assign inbar[121] = ~in[121];
  assign inbar[122] = ~in[122];
  assign inbar[123] = ~in[123];
  assign inbar[124] = ~in[124];
  assign inbar[125] = ~in[125];
  assign inbar[126] = ~in[126];
  assign inbar[127] = ~in[127];
  assign inbar[128] = ~in[128];
  assign inbar[129] = ~in[129];
  assign inbar[130] = ~in[130];
  assign inbar[131] = ~in[131];
  assign inbar[132] = ~in[132];
  assign inbar[133] = ~in[133];
  assign inbar[134] = ~in[134];
  assign inbar[135] = ~in[135];
  assign inbar[136] = ~in[136];
  assign inbar[137] = ~in[137];
  assign inbar[138] = ~in[138];
  assign inbar[139] = ~in[139];
  assign inbar[140] = ~in[140];
  assign inbar[141] = ~in[141];
  assign inbar[142] = ~in[142];
  assign inbar[143] = ~in[143];
  assign inbar[144] = ~in[144];
  assign inbar[145] = ~in[145];
  assign inbar[146] = ~in[146];
  assign inbar[147] = ~in[147];
  assign inbar[148] = ~in[148];
  assign inbar[149] = ~in[149];
  assign inbar[150] = ~in[150];
  assign inbar[151] = ~in[151];
  assign inbar[152] = ~in[152];
  assign inbar[153] = ~in[153];
  assign inbar[154] = ~in[154];
  assign inbar[155] = ~in[155];
  assign inbar[156] = ~in[156];
  assign inbar[157] = ~in[157];
  assign inbar[158] = ~in[158];
  assign inbar[159] = ~in[159];
  assign inbar[160] = ~in[160];
  assign inbar[161] = ~in[161];
  assign inbar[162] = ~in[162];
  assign inbar[163] = ~in[163];
  assign inbar[164] = ~in[164];
  assign inbar[165] = ~in[165];
  assign inbar[166] = ~in[166];
  assign inbar[167] = ~in[167];
  assign inbar[168] = ~in[168];
  assign inbar[169] = ~in[169];
  assign inbar[170] = ~in[170];
  assign inbar[171] = ~in[171];
  assign inbar[172] = ~in[172];
  assign inbar[173] = ~in[173];
  assign inbar[174] = ~in[174];
  assign inbar[175] = ~in[175];
  assign inbar[176] = ~in[176];
  assign inbar[177] = ~in[177];
  assign inbar[178] = ~in[178];
  assign inbar[179] = ~in[179];
  assign inbar[180] = ~in[180];
  assign inbar[181] = ~in[181];
  assign inbar[182] = ~in[182];
  assign inbar[183] = ~in[183];
  assign inbar[184] = ~in[184];
  assign inbar[185] = ~in[185];
  assign inbar[186] = ~in[186];
  assign inbar[187] = ~in[187];
  assign inbar[188] = ~in[188];
  assign inbar[189] = ~in[189];
  assign inbar[190] = ~in[190];
  assign inbar[191] = ~in[191];
  assign inbar[192] = ~in[192];
  assign inbar[193] = ~in[193];
  assign inbar[194] = ~in[194];
  assign inbar[195] = ~in[195];
  assign inbar[196] = ~in[196];
  assign inbar[197] = ~in[197];
  assign inbar[198] = ~in[198];
  assign inbar[199] = ~in[199];
  assign inbar[200] = ~in[200];
  assign inbar[201] = ~in[201];
  assign inbar[202] = ~in[202];
  assign inbar[203] = ~in[203];
  assign inbar[204] = ~in[204];
  assign inbar[205] = ~in[205];
  assign inbar[206] = ~in[206];
  assign inbar[207] = ~in[207];
  assign inbar[208] = ~in[208];
  assign inbar[209] = ~in[209];
  assign inbar[210] = ~in[210];
  assign inbar[211] = ~in[211];
  assign inbar[212] = ~in[212];
  assign inbar[213] = ~in[213];
  assign inbar[214] = ~in[214];
  assign inbar[215] = ~in[215];
  assign inbar[216] = ~in[216];
  assign inbar[217] = ~in[217];
  assign inbar[218] = ~in[218];
  assign inbar[219] = ~in[219];
  assign inbar[220] = ~in[220];
  assign inbar[221] = ~in[221];
  assign inbar[222] = ~in[222];
  assign inbar[223] = ~in[223];
  assign inbar[224] = ~in[224];
  assign inbar[225] = ~in[225];
  assign inbar[226] = ~in[226];
  assign inbar[227] = ~in[227];
  assign inbar[228] = ~in[228];
  assign inbar[229] = ~in[229];
  assign inbar[230] = ~in[230];
  assign inbar[231] = ~in[231];
  assign inbar[232] = ~in[232];
  assign inbar[233] = ~in[233];
  assign inbar[234] = ~in[234];
  assign inbar[235] = ~in[235];
  assign inbar[236] = ~in[236];
  assign inbar[237] = ~in[237];
  assign inbar[238] = ~in[238];
  assign inbar[239] = ~in[239];
  assign inbar[240] = ~in[240];
  assign inbar[241] = ~in[241];
  assign inbar[242] = ~in[242];
  assign inbar[243] = ~in[243];
  assign inbar[244] = ~in[244];
  assign inbar[245] = ~in[245];
  assign inbar[246] = ~in[246];
  assign inbar[247] = ~in[247];
  assign inbar[248] = ~in[248];
  assign inbar[249] = ~in[249];
  assign inbar[250] = ~in[250];
  assign inbar[251] = ~in[251];
  assign inbar[252] = ~in[252];
  assign inbar[253] = ~in[253];
  assign inbar[254] = ~in[254];
  assign inbar[255] = ~in[255];
//input_done

  output wire [7:0] out;
  wire [7:0] outbar;
//output_done

  wire in_81;
  wire in_80;
  wire in_79;
  wire in_78;
  wire in_77;
  wire in_76;
  wire in_75;
  wire in_74;
  wire in_73;
  wire in_72;
  wire in_71;
  wire in_70;
  wire in_69;
  wire in_68;
  wire in_67;
  wire in_66;
  wire in_65;
  wire in_64;
  wire in_63;
  wire in_62;
  wire in_61;
  wire in_60;
  wire in_59;
  wire in_58;
  wire in_57;
  wire in_56;
  wire in_55;
  wire in_54;
  wire in_53;
  wire in_52;
  wire in_51;
  wire in_50;
  wire in_49;
  wire in_48;
  wire in_47;
  wire in_46;
  wire in_45;
  wire in_44;
  wire in_43;
  wire in_42;
  wire in_41;
  wire in_40;
  wire in_39;
  wire in_38;
  wire in_37;
  wire in_36;
  wire in_35;
  wire in_34;
  wire in_33;
  wire in_32;
  wire in_31;
  wire in_30;
  wire in_29;
  wire in_28;
  wire in_27;
  wire in_26;
  wire in_25;
  wire in_24;
  wire in_23;
  wire in_22;
  wire in_21;
  wire in_20;
  wire in_19;
  wire in_18;
  wire in_17;
  wire in_16;
  wire in_15;
  wire in_14;
  wire in_13;
  wire in_12;
  wire in_11;
  wire in_10;
  wire in_9;
  wire in_8;
  wire in_7;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_3;
  wire in_2;
  wire in_1;
  wire in_0;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire in_81bar;
  wire in_80bar;
  wire in_79bar;
  wire in_78bar;
  wire in_77bar;
  wire in_76bar;
  wire in_75bar;
  wire in_74bar;
  wire in_73bar;
  wire in_72bar;
  wire in_71bar;
  wire in_70bar;
  wire in_69bar;
  wire in_68bar;
  wire in_67bar;
  wire in_66bar;
  wire in_65bar;
  wire in_64bar;
  wire in_63bar;
  wire in_62bar;
  wire in_61bar;
  wire in_60bar;
  wire in_59bar;
  wire in_58bar;
  wire in_57bar;
  wire in_56bar;
  wire in_55bar;
  wire in_54bar;
  wire in_53bar;
  wire in_52bar;
  wire in_51bar;
  wire in_50bar;
  wire in_49bar;
  wire in_48bar;
  wire in_47bar;
  wire in_46bar;
  wire in_45bar;
  wire in_44bar;
  wire in_43bar;
  wire in_42bar;
  wire in_41bar;
  wire in_40bar;
  wire in_39bar;
  wire in_38bar;
  wire in_37bar;
  wire in_36bar;
  wire in_35bar;
  wire in_34bar;
  wire in_33bar;
  wire in_32bar;
  wire in_31bar;
  wire in_30bar;
  wire in_29bar;
  wire in_28bar;
  wire in_27bar;
  wire in_26bar;
  wire in_25bar;
  wire in_24bar;
  wire in_23bar;
  wire in_22bar;
  wire in_21bar;
  wire in_20bar;
  wire in_19bar;
  wire in_18bar;
  wire in_17bar;
  wire in_16bar;
  wire in_15bar;
  wire in_14bar;
  wire in_13bar;
  wire in_12bar;
  wire in_11bar;
  wire in_10bar;
  wire in_9bar;
  wire in_8bar;
  wire in_7bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_3bar;
  wire in_2bar;
  wire in_1bar;
  wire in_0bar;
  wire n487bar;
  wire n488bar;
  wire n489bar;
  wire n490bar;
  wire n491bar;
  wire n492bar;
  wire n493bar;
  wire n494bar;
  wire n495bar;
  wire n496bar;
  wire n497bar;
  wire n498bar;
  wire n499bar;
  wire n500bar;
  wire n501bar;
  wire n502bar;
  wire n503bar;
  wire n504bar;
  wire n505bar;
  wire n506bar;
  wire n507bar;
  wire n508bar;
  wire n509bar;
  wire n510bar;
  wire n511bar;
  wire n512bar;
  wire n513bar;
  wire n514bar;
  wire n515bar;
  wire n516bar;
  wire n517bar;
  wire n518bar;
  wire n519bar;
  wire n520bar;
  wire n521bar;
  wire n522bar;
  wire n523bar;
  wire n524bar;
  wire n525bar;
  wire n526bar;
  wire n527bar;
  wire n528bar;
  wire n529bar;
  wire n530bar;
  wire n531bar;
  wire n532bar;
  wire n533bar;
  wire n534bar;
  wire n535bar;
  wire n536bar;
  wire n537bar;
  wire n538bar;
  wire n539bar;
  wire n540bar;
  wire n541bar;
  wire n542bar;
  wire n543bar;
  wire n544bar;
  wire n545bar;
  wire n546bar;
  wire n547bar;
  wire n548bar;
  wire n549bar;
  wire n550bar;
  wire n551bar;
  wire n552bar;
  wire n553bar;
  wire n554bar;
  wire n555bar;
  wire n556bar;
  wire n557bar;
  wire n558bar;
  wire n559bar;
  wire n560bar;
  wire n561bar;
  wire n562bar;
  wire n563bar;
  wire n564bar;
  wire n565bar;
  wire n566bar;
  wire n567bar;
  wire n568bar;
  wire n569bar;
  wire n570bar;
  wire n571bar;
  wire n572bar;
  wire n573bar;
  wire n574bar;
  wire n575bar;
  wire n576bar;
  wire n577bar;
  wire n578bar;
  wire n579bar;
  wire n580bar;
  wire n581bar;
  wire n582bar;
  wire n583bar;
  wire n584bar;
  wire n585bar;
  wire n586bar;
  wire n587bar;
  wire n588bar;
  wire n589bar;
  wire n590bar;
  wire n591bar;
  wire n592bar;
  wire n593bar;
  wire n594bar;
  wire n595bar;
  wire n596bar;
  wire n597bar;
  wire n598bar;
  wire n599bar;
  wire n600bar;
  wire n601bar;
  wire n602bar;
  wire n603bar;
  wire n604bar;
  wire n605bar;
  wire n606bar;
  wire n607bar;
  wire n608bar;
  wire n609bar;
  wire n610bar;
  wire n611bar;
  wire n612bar;
  wire n613bar;
  wire n614bar;
  wire n615bar;
  wire n616bar;
  wire n617bar;
  wire n618bar;
  wire n619bar;
  wire n620bar;
  wire n621bar;
  wire n622bar;
  wire n623bar;
  wire n624bar;
  wire n625bar;
  wire n626bar;
  wire n627bar;
  wire n628bar;
  wire n629bar;
  wire n630bar;
  wire n631bar;
  wire n632bar;
  wire n633bar;
  wire n634bar;
  wire n635bar;
  wire n636bar;
  wire n637bar;
  wire n638bar;
  wire n639bar;
  wire n640bar;
  wire n641bar;
  wire n642bar;
  wire n643bar;
  wire n644bar;
  wire n645bar;
  wire n646bar;
  wire n647bar;
  wire n648bar;
  wire n649bar;
  wire n650bar;
  wire n651bar;
  wire n652bar;
  wire n653bar;
  wire n654bar;
  wire n655bar;
  wire n656bar;
  wire n657bar;
  wire n658bar;
  wire n659bar;
  wire n660bar;
  wire n661bar;
  wire n662bar;
  wire n663bar;
  wire n664bar;
  wire n665bar;
  wire n666bar;
  wire n667bar;
  wire n668bar;
  wire n669bar;
  wire n670bar;
  wire n671bar;
  wire n672bar;
  wire n673bar;
  wire n674bar;
  wire n675bar;
  wire n676bar;
  wire n677bar;
  wire n678bar;
  wire n679bar;
  wire n680bar;
  wire n681bar;
  wire n682bar;
  wire n683bar;
  wire n684bar;
  wire n685bar;
  wire n686bar;
  wire n687bar;
  wire n688bar;
  wire n689bar;
  wire n690bar;
  wire n691bar;
  wire n692bar;
  wire n693bar;
  wire n694bar;
  wire n695bar;
  wire n696bar;
  wire n697bar;
  wire n698bar;
  wire n699bar;
  wire n700bar;
  wire n701bar;
  wire n702bar;
  wire n703bar;
  wire n704bar;
  wire n705bar;
  wire n706bar;
  wire n707bar;
  wire n708bar;
  wire n709bar;
  wire n710bar;
  wire n711bar;
  wire n712bar;
  wire n713bar;
  wire n714bar;
  wire n715bar;
  wire n716bar;
  wire n717bar;
  wire n718bar;
  wire n719bar;
  wire n720bar;
  wire n721bar;
  wire n722bar;
  wire n723bar;
  wire n724bar;
  wire n725bar;
  wire n726bar;
  wire n727bar;
  wire n728bar;
  wire n729bar;
  wire n730bar;
  wire n731bar;
  wire n732bar;
  wire n733bar;
  wire n734bar;
  wire n735bar;
  wire n736bar;
  wire n737bar;
  wire n738bar;
  wire n739bar;
  wire n740bar;
  wire n741bar;
  wire n742bar;
  wire n743bar;
  wire n744bar;
  wire n745bar;
  wire n746bar;
  wire n747bar;
  wire n748bar;
  wire n749bar;
  wire n750bar;
  wire n751bar;
  wire n752bar;
  wire n753bar;
  wire n754bar;
  wire n755bar;
  wire n756bar;
  wire n757bar;
  wire n758bar;
  wire n759bar;
  wire n760bar;
  wire n761bar;
  wire n762bar;
  wire n763bar;
  wire n764bar;
  wire n765bar;
  wire n766bar;
  wire n767bar;
  wire n768bar;
  wire n769bar;
  wire n770bar;
  wire n771bar;
  wire n772bar;
  wire n773bar;
  wire n774bar;
  wire n775bar;
  wire n776bar;
  wire n777bar;
  wire n778bar;
  wire n779bar;
  wire n780bar;
  wire n781bar;
  wire n782bar;
  wire n783bar;
  wire n784bar;
  wire n785bar;
  wire n786bar;
  wire n787bar;
  wire n788bar;
  wire n789bar;
  wire n790bar;
  wire n791bar;
  wire n792bar;
  wire n793bar;
  wire n794bar;
  wire n795bar;
  wire n796bar;
  wire n797bar;
  wire n798bar;
  wire n799bar;
  wire n800bar;
  wire n801bar;
  wire n802bar;
  wire n803bar;
  wire n804bar;
  wire n805bar;
  wire n806bar;
  wire n807bar;
  wire n808bar;
  wire n809bar;
  wire n810bar;
  wire n811bar;
  wire n812bar;
  wire n813bar;
  wire n814bar;
  wire n815bar;
  wire n816bar;
  wire n817bar;
  wire n818bar;
  wire n819bar;
  wire n820bar;
  wire n821bar;
  wire n822bar;
  wire n823bar;
  wire n824bar;
  wire n825bar;
  wire n826bar;
  wire n827bar;
  wire n828bar;
  wire n829bar;
  wire n830bar;
  wire n831bar;
  wire n832bar;
  wire n833bar;
  wire n834bar;
  wire n835bar;
  wire n836bar;
  wire n837bar;
  wire n838bar;
  wire n839bar;
  wire n840bar;
  wire n841bar;
  wire n842bar;
  wire n843bar;
  wire n844bar;
  wire n845bar;
  wire n846bar;
  wire n847bar;
  wire n848bar;
  wire n849bar;
  wire n850bar;
  wire n851bar;
  wire n852bar;
  wire n853bar;
  wire n854bar;
  wire n855bar;
  wire n856bar;
  wire n857bar;
  wire n858bar;
  wire n859bar;
  wire n860bar;
  wire n861bar;
  wire n862bar;
  wire n863bar;
  wire n864bar;
  wire n865bar;
  wire n866bar;
  wire n867bar;
  wire n868bar;
  wire n869bar;
  wire n870bar;
  wire n871bar;
  wire n872bar;
  wire n873bar;
  wire n874bar;
  wire n875bar;
  wire n876bar;
  wire n877bar;
  wire n878bar;
  wire n879bar;
  wire n880bar;
  wire n881bar;
  wire n882bar;
  wire n883bar;
  wire n884bar;
  wire n885bar;
  wire n886bar;
  wire n887bar;
  wire n888bar;
  wire n889bar;
  wire n890bar;
  wire n891bar;
  wire n892bar;
  wire n893bar;
  wire n894bar;
  wire n895bar;
  wire n896bar;
  wire n897bar;
  wire n898bar;
  wire n899bar;
  wire n900bar;
  wire n901bar;
  wire n902bar;
  wire n903bar;
  wire n904bar;
  wire n905bar;
  wire n906bar;
  wire n907bar;
  wire n908bar;
  wire n909bar;
  wire n910bar;
  wire n911bar;
  wire n912bar;
  wire n913bar;
  wire n914bar;
  wire n915bar;
  wire n916bar;
  wire n917bar;
  wire n918bar;
  wire n919bar;
  wire n920bar;
  wire n921bar;
  wire n922bar;
  wire n923bar;
  wire n924bar;
  wire n925bar;
  wire n926bar;
  wire n927bar;
  wire n928bar;
  wire n929bar;
  wire n930bar;
  wire n931bar;
  wire n932bar;
  wire n933bar;
  wire n934bar;
  wire n935bar;
  wire n936bar;
  wire n937bar;
  wire n938bar;
  wire n939bar;
  wire n940bar;
  wire n941bar;
  wire n942bar;
  wire n943bar;
  wire n944bar;
  wire n945bar;
  wire n946bar;
  wire n947bar;
  wire n948bar;
  wire n949bar;
  wire n950bar;
  wire n951bar;
  wire n952bar;
  wire n953bar;
  wire n954bar;
  wire n955bar;
  wire n956bar;
  wire n957bar;
  wire n958bar;
  wire n959bar;
  wire n960bar;
  wire n961bar;
  wire n962bar;
  wire n963bar;
  wire n964bar;
  wire n965bar;
  wire n966bar;
  wire n967bar;
  wire n968bar;
  wire n969bar;
  wire n970bar;
  wire n971bar;
  wire n972bar;
//wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];
  //OR U1
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1 (
    .O(out[7]),
    .I0(n972),
    .I1(n971)
  );
  //AND U1bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1bar (
    .O(outbar[7]),
    .I0(n972bar),
    .I1(n971bar)
  );
  //OR U2
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2 (
    .O(n971),
    .I0(n970),
    .I1(n969)
  );
  //AND U2bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2bar (
    .O(n971bar),
    .I0(n970bar),
    .I1(n969bar)
  );
  //OR U3
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3 (
    .O(n969),
    .I0(n968),
    .I1(n967)
  );
  //AND U3bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3bar (
    .O(n969bar),
    .I0(n968bar),
    .I1(n967bar)
  );
  //OR U4
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4 (
    .O(n967),
    .I0(n966),
    .I1(n965)
  );
  //AND U4bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4bar (
    .O(n967bar),
    .I0(n966bar),
    .I1(n965bar)
  );
  //OR U5
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5 (
    .O(n968),
    .I0(n964),
    .I1(n963)
  );
  //AND U5bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5bar (
    .O(n968bar),
    .I0(n964bar),
    .I1(n963bar)
  );
  //OR U6
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6 (
    .O(n963),
    .I0(in[116]),
    .I1(n962)
  );
  //AND U6bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6bar (
    .O(n963bar),
    .I0(inbar[116]),
    .I1(n962bar)
  );
  //OR U7
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7 (
    .O(n970),
    .I0(n961),
    .I1(n960)
  );
  //AND U7bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7bar (
    .O(n970bar),
    .I0(n961bar),
    .I1(n960bar)
  );
  //OR U8
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8 (
    .O(n960),
    .I0(in[150]),
    .I1(in[127])
  );
  //AND U8bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8bar (
    .O(n960bar),
    .I0(inbar[150]),
    .I1(inbar[127])
  );
  //OR U9
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9 (
    .O(n961),
    .I0(in[160]),
    .I1(n959)
  );
  //AND U9bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9bar (
    .O(n961bar),
    .I0(inbar[160]),
    .I1(n959bar)
  );
  //OR U10
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10 (
    .O(n959),
    .I0(in[252]),
    .I1(in[168])
  );
  //AND U10bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10bar (
    .O(n959bar),
    .I0(inbar[252]),
    .I1(inbar[168])
  );
  //OR U11
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11 (
    .O(n972),
    .I0(n958),
    .I1(n957)
  );
  //AND U11bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11bar (
    .O(n972bar),
    .I0(n958bar),
    .I1(n957bar)
  );
  //OR U12
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12 (
    .O(n957),
    .I0(n956),
    .I1(n955)
  );
  //AND U12bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12bar (
    .O(n957bar),
    .I0(n956bar),
    .I1(n955bar)
  );
  //OR U13
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13 (
    .O(n955),
    .I0(in_17),
    .I1(in[96])
  );
  //AND U13bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13bar (
    .O(n955bar),
    .I0(in_17bar),
    .I1(inbar[96])
  );
  //OR U14
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14 (
    .O(n956),
    .I0(in_23),
    .I1(n954)
  );
  //AND U14bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14bar (
    .O(n956bar),
    .I0(in_23bar),
    .I1(n954bar)
  );
  //OR U15
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15 (
    .O(n954),
    .I0(in_31),
    .I1(in_26)
  );
  //AND U15bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15bar (
    .O(n954bar),
    .I0(in_31bar),
    .I1(in_26bar)
  );
  //OR U16
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16 (
    .O(n958),
    .I0(n953),
    .I1(n952)
  );
  //AND U16bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16bar (
    .O(n958bar),
    .I0(n953bar),
    .I1(n952bar)
  );
  //OR U17
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U17 (
    .O(n952),
    .I0(in_58),
    .I1(in_4)
  );
  //AND U17bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U17bar (
    .O(n952bar),
    .I0(in_58bar),
    .I1(in_4bar)
  );
  //OR U18
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U18 (
    .O(n953),
    .I0(in_59),
    .I1(n951)
  );
  //AND U18bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U18bar (
    .O(n953bar),
    .I0(in_59bar),
    .I1(n951bar)
  );
  //OR U19
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U19 (
    .O(n951),
    .I0(in_71),
    .I1(in_62)
  );
  //AND U19bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U19bar (
    .O(n951bar),
    .I0(in_71bar),
    .I1(in_62bar)
  );
  //OR U20
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U20 (
    .O(out[6]),
    .I0(n950),
    .I1(n949)
  );
  //AND U20bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U20bar (
    .O(outbar[6]),
    .I0(n950bar),
    .I1(n949bar)
  );
  //OR U21
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U21 (
    .O(n949),
    .I0(n948),
    .I1(n947)
  );
  //AND U21bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U21bar (
    .O(n949bar),
    .I0(n948bar),
    .I1(n947bar)
  );
  //OR U22
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U22 (
    .O(n947),
    .I0(n946),
    .I1(n945)
  );
  //AND U22bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U22bar (
    .O(n947bar),
    .I0(n946bar),
    .I1(n945bar)
  );
  //OR U23
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U23 (
    .O(n945),
    .I0(n944),
    .I1(n943)
  );
  //AND U23bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U23bar (
    .O(n945bar),
    .I0(n944bar),
    .I1(n943bar)
  );
  //OR U24
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U24 (
    .O(n946),
    .I0(n942),
    .I1(n941)
  );
  //AND U24bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U24bar (
    .O(n946bar),
    .I0(n942bar),
    .I1(n941bar)
  );
  //OR U25
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U25 (
    .O(n941),
    .I0(in[101]),
    .I1(n940)
  );
  //AND U25bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U25bar (
    .O(n941bar),
    .I0(inbar[101]),
    .I1(n940bar)
  );
  //OR U26
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U26 (
    .O(n948),
    .I0(n939),
    .I1(n938)
  );
  //AND U26bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U26bar (
    .O(n948bar),
    .I0(n939bar),
    .I1(n938bar)
  );
  //OR U27
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U27 (
    .O(n938),
    .I0(in[114]),
    .I1(in[104])
  );
  //AND U27bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U27bar (
    .O(n938bar),
    .I0(inbar[114]),
    .I1(inbar[104])
  );
  //OR U28
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U28 (
    .O(n939),
    .I0(in[128]),
    .I1(n937)
  );
  //AND U28bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U28bar (
    .O(n939bar),
    .I0(inbar[128]),
    .I1(n937bar)
  );
  //OR U29
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U29 (
    .O(n937),
    .I0(in[136]),
    .I1(in[134])
  );
  //AND U29bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U29bar (
    .O(n937bar),
    .I0(inbar[136]),
    .I1(inbar[134])
  );
  //OR U30
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U30 (
    .O(n950),
    .I0(n936),
    .I1(n935)
  );
  //AND U30bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U30bar (
    .O(n950bar),
    .I0(n936bar),
    .I1(n935bar)
  );
  //OR U31
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U31 (
    .O(n935),
    .I0(n934),
    .I1(n933)
  );
  //AND U31bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U31bar (
    .O(n935bar),
    .I0(n934bar),
    .I1(n933bar)
  );
  //OR U32
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U32 (
    .O(n933),
    .I0(in[177]),
    .I1(in[164])
  );
  //AND U32bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U32bar (
    .O(n933bar),
    .I0(inbar[177]),
    .I1(inbar[164])
  );
  //OR U33
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U33 (
    .O(n934),
    .I0(in[212]),
    .I1(n932)
  );
  //AND U33bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U33bar (
    .O(n934bar),
    .I0(inbar[212]),
    .I1(n932bar)
  );
  //OR U34
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U34 (
    .O(n932),
    .I0(in[248]),
    .I1(in[221])
  );
  //AND U34bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U34bar (
    .O(n932bar),
    .I0(inbar[248]),
    .I1(inbar[221])
  );
  //OR U35
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U35 (
    .O(n936),
    .I0(n931),
    .I1(n930)
  );
  //AND U35bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U35bar (
    .O(n936bar),
    .I0(n931bar),
    .I1(n930bar)
  );
  //OR U36
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U36 (
    .O(n930),
    .I0(in_18),
    .I1(in[93])
  );
  //AND U36bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U36bar (
    .O(n930bar),
    .I0(in_18bar),
    .I1(inbar[93])
  );
  //OR U37
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U37 (
    .O(n931),
    .I0(in_31),
    .I1(n929)
  );
  //AND U37bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U37bar (
    .O(n931bar),
    .I0(in_31bar),
    .I1(n929bar)
  );
  //OR U38
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U38 (
    .O(n929),
    .I0(in_7),
    .I1(in_39)
  );
  //AND U38bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U38bar (
    .O(n929bar),
    .I0(in_7bar),
    .I1(in_39bar)
  );
  //OR U39
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U39 (
    .O(out[5]),
    .I0(n928),
    .I1(n927)
  );
  //AND U39bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U39bar (
    .O(outbar[5]),
    .I0(n928bar),
    .I1(n927bar)
  );
  //OR U40
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U40 (
    .O(n927),
    .I0(n926),
    .I1(n925)
  );
  //AND U40bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U40bar (
    .O(n927bar),
    .I0(n926bar),
    .I1(n925bar)
  );
  //OR U41
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U41 (
    .O(n925),
    .I0(n924),
    .I1(n923)
  );
  //AND U41bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U41bar (
    .O(n925bar),
    .I0(n924bar),
    .I1(n923bar)
  );
  //OR U42
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U42 (
    .O(n923),
    .I0(n922),
    .I1(n921)
  );
  //AND U42bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U42bar (
    .O(n923bar),
    .I0(n922bar),
    .I1(n921bar)
  );
  //OR U43
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U43 (
    .O(n924),
    .I0(n940),
    .I1(n920)
  );
  //AND U43bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U43bar (
    .O(n924bar),
    .I0(n940bar),
    .I1(n920bar)
  );
  //OR U44
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U44 (
    .O(n920),
    .I0(in[111]),
    .I1(n919)
  );
  //AND U44bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U44bar (
    .O(n920bar),
    .I0(inbar[111]),
    .I1(n919bar)
  );
  //OR U45
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U45 (
    .O(n940),
    .I0(n918),
    .I1(n917)
  );
  //AND U45bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U45bar (
    .O(n940bar),
    .I0(n918bar),
    .I1(n917bar)
  );
  //OR U46
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U46 (
    .O(n917),
    .I0(n916),
    .I1(n915)
  );
  //AND U46bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U46bar (
    .O(n917bar),
    .I0(n916bar),
    .I1(n915bar)
  );
  //OR U47
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U47 (
    .O(n915),
    .I0(n914),
    .I1(n913)
  );
  //AND U47bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U47bar (
    .O(n915bar),
    .I0(n914bar),
    .I1(n913bar)
  );
  //OR U48
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U48 (
    .O(n913),
    .I0(in[140]),
    .I1(in[131])
  );
  //AND U48bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U48bar (
    .O(n913bar),
    .I0(inbar[140]),
    .I1(inbar[131])
  );
  //OR U49
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U49 (
    .O(n914),
    .I0(in[160]),
    .I1(in[144])
  );
  //AND U49bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U49bar (
    .O(n914bar),
    .I0(inbar[160]),
    .I1(inbar[144])
  );
  //OR U50
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U50 (
    .O(n916),
    .I0(n912),
    .I1(n911)
  );
  //AND U50bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U50bar (
    .O(n916bar),
    .I0(n912bar),
    .I1(n911bar)
  );
  //OR U51
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U51 (
    .O(n911),
    .I0(in[179]),
    .I1(in[174])
  );
  //AND U51bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U51bar (
    .O(n911bar),
    .I0(inbar[179]),
    .I1(inbar[174])
  );
  //OR U52
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U52 (
    .O(n912),
    .I0(in[188]),
    .I1(in[184])
  );
  //AND U52bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U52bar (
    .O(n912bar),
    .I0(inbar[188]),
    .I1(inbar[184])
  );
  //OR U53
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U53 (
    .O(n918),
    .I0(n910),
    .I1(n909)
  );
  //AND U53bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U53bar (
    .O(n918bar),
    .I0(n910bar),
    .I1(n909bar)
  );
  //OR U54
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U54 (
    .O(n909),
    .I0(n908),
    .I1(n907)
  );
  //AND U54bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U54bar (
    .O(n909bar),
    .I0(n908bar),
    .I1(n907bar)
  );
  //OR U55
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U55 (
    .O(n907),
    .I0(in[216]),
    .I1(in[200])
  );
  //AND U55bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U55bar (
    .O(n907bar),
    .I0(inbar[216]),
    .I1(inbar[200])
  );
  //OR U56
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U56 (
    .O(n908),
    .I0(in[228]),
    .I1(in[224])
  );
  //AND U56bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U56bar (
    .O(n908bar),
    .I0(inbar[228]),
    .I1(inbar[224])
  );
  //OR U57
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U57 (
    .O(n910),
    .I0(n906),
    .I1(n905)
  );
  //AND U57bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U57bar (
    .O(n910bar),
    .I0(n906bar),
    .I1(n905bar)
  );
  //OR U58
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U58 (
    .O(n905),
    .I0(in[247]),
    .I1(in[235])
  );
  //AND U58bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U58bar (
    .O(n905bar),
    .I0(inbar[247]),
    .I1(inbar[235])
  );
  //OR U59
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U59 (
    .O(n906),
    .I0(in_42),
    .I1(in[83])
  );
  //AND U59bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U59bar (
    .O(n906bar),
    .I0(in_42bar),
    .I1(inbar[83])
  );
  //OR U60
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U60 (
    .O(n926),
    .I0(n904),
    .I1(n903)
  );
  //AND U60bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U60bar (
    .O(n926bar),
    .I0(n904bar),
    .I1(n903bar)
  );
  //OR U61
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U61 (
    .O(n903),
    .I0(in[166]),
    .I1(in[123])
  );
  //AND U61bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U61bar (
    .O(n903bar),
    .I0(inbar[166]),
    .I1(inbar[123])
  );
  //OR U62
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U62 (
    .O(n904),
    .I0(in[170]),
    .I1(n902)
  );
  //AND U62bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U62bar (
    .O(n904bar),
    .I0(inbar[170]),
    .I1(n902bar)
  );
  //OR U63
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U63 (
    .O(n902),
    .I0(in[194]),
    .I1(in[183])
  );
  //AND U63bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U63bar (
    .O(n902bar),
    .I0(inbar[194]),
    .I1(inbar[183])
  );
  //OR U64
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U64 (
    .O(n928),
    .I0(n901),
    .I1(n900)
  );
  //AND U64bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U64bar (
    .O(n928bar),
    .I0(n901bar),
    .I1(n900bar)
  );
  //OR U65
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U65 (
    .O(n900),
    .I0(n899),
    .I1(n898)
  );
  //AND U65bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U65bar (
    .O(n900bar),
    .I0(n899bar),
    .I1(n898bar)
  );
  //OR U66
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U66 (
    .O(n898),
    .I0(in[241]),
    .I1(in[238])
  );
  //AND U66bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U66bar (
    .O(n898bar),
    .I0(inbar[241]),
    .I1(inbar[238])
  );
  //OR U67
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U67 (
    .O(n899),
    .I0(in[250]),
    .I1(n897)
  );
  //AND U67bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U67bar (
    .O(n899bar),
    .I0(inbar[250]),
    .I1(n897bar)
  );
  //OR U68
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U68 (
    .O(n897),
    .I0(in_24),
    .I1(in[84])
  );
  //AND U68bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U68bar (
    .O(n897bar),
    .I0(in_24bar),
    .I1(inbar[84])
  );
  //OR U69
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U69 (
    .O(n901),
    .I0(n896),
    .I1(n895)
  );
  //AND U69bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U69bar (
    .O(n901bar),
    .I0(n896bar),
    .I1(n895bar)
  );
  //OR U70
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U70 (
    .O(n895),
    .I0(in_41),
    .I1(in_29)
  );
  //AND U70bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U70bar (
    .O(n895bar),
    .I0(in_41bar),
    .I1(in_29bar)
  );
  //OR U71
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U71 (
    .O(n896),
    .I0(in_66),
    .I1(n894)
  );
  //AND U71bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U71bar (
    .O(n896bar),
    .I0(in_66bar),
    .I1(n894bar)
  );
  //OR U72
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U72 (
    .O(n894),
    .I0(in_76),
    .I1(in_71)
  );
  //AND U72bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U72bar (
    .O(n894bar),
    .I0(in_76bar),
    .I1(in_71bar)
  );
  //OR U73
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U73 (
    .O(out[4]),
    .I0(n893),
    .I1(n892)
  );
  //AND U73bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U73bar (
    .O(outbar[4]),
    .I0(n893bar),
    .I1(n892bar)
  );
  //OR U74
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U74 (
    .O(n892),
    .I0(n891),
    .I1(n890)
  );
  //AND U74bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U74bar (
    .O(n892bar),
    .I0(n891bar),
    .I1(n890bar)
  );
  //OR U75
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U75 (
    .O(n890),
    .I0(n889),
    .I1(n888)
  );
  //AND U75bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U75bar (
    .O(n890bar),
    .I0(n889bar),
    .I1(n888bar)
  );
  //OR U76
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U76 (
    .O(n888),
    .I0(n922),
    .I1(n887)
  );
  //AND U76bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U76bar (
    .O(n888bar),
    .I0(n922bar),
    .I1(n887bar)
  );
  //OR U77
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U77 (
    .O(n922),
    .I0(n886),
    .I1(n885)
  );
  //AND U77bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U77bar (
    .O(n922bar),
    .I0(n886bar),
    .I1(n885bar)
  );
  //OR U78
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U78 (
    .O(n885),
    .I0(n884),
    .I1(n883)
  );
  //AND U78bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U78bar (
    .O(n885bar),
    .I0(n884bar),
    .I1(n883bar)
  );
  //OR U79
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U79 (
    .O(n883),
    .I0(n882),
    .I1(n881)
  );
  //AND U79bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U79bar (
    .O(n883bar),
    .I0(n882bar),
    .I1(n881bar)
  );
  //OR U80
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U80 (
    .O(n881),
    .I0(in[118]),
    .I1(in[109])
  );
  //AND U80bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U80bar (
    .O(n881bar),
    .I0(inbar[118]),
    .I1(inbar[109])
  );
  //OR U81
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U81 (
    .O(n882),
    .I0(in[139]),
    .I1(in[120])
  );
  //AND U81bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U81bar (
    .O(n882bar),
    .I0(inbar[139]),
    .I1(inbar[120])
  );
  //OR U82
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U82 (
    .O(n884),
    .I0(n880),
    .I1(n879)
  );
  //AND U82bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U82bar (
    .O(n884bar),
    .I0(n880bar),
    .I1(n879bar)
  );
  //OR U83
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U83 (
    .O(n879),
    .I0(in[198]),
    .I1(in[154])
  );
  //AND U83bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U83bar (
    .O(n879bar),
    .I0(inbar[198]),
    .I1(inbar[154])
  );
  //OR U84
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U84 (
    .O(n880),
    .I0(in[210]),
    .I1(in[205])
  );
  //AND U84bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U84bar (
    .O(n880bar),
    .I0(inbar[210]),
    .I1(inbar[205])
  );
  //OR U85
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U85 (
    .O(n886),
    .I0(n878),
    .I1(n877)
  );
  //AND U85bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U85bar (
    .O(n886bar),
    .I0(n878bar),
    .I1(n877bar)
  );
  //OR U86
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U86 (
    .O(n877),
    .I0(n876),
    .I1(n875)
  );
  //AND U86bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U86bar (
    .O(n877bar),
    .I0(n876bar),
    .I1(n875bar)
  );
  //OR U87
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U87 (
    .O(n875),
    .I0(in[219]),
    .I1(in[217])
  );
  //AND U87bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U87bar (
    .O(n875bar),
    .I0(inbar[219]),
    .I1(inbar[217])
  );
  //OR U88
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U88 (
    .O(n876),
    .I0(in[86]),
    .I1(in[252])
  );
  //AND U88bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U88bar (
    .O(n876bar),
    .I0(inbar[86]),
    .I1(inbar[252])
  );
  //OR U89
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U89 (
    .O(n878),
    .I0(n874),
    .I1(n873)
  );
  //AND U89bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U89bar (
    .O(n878bar),
    .I0(n874bar),
    .I1(n873bar)
  );
  //OR U90
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U90 (
    .O(n873),
    .I0(in_40),
    .I1(in[91])
  );
  //AND U90bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U90bar (
    .O(n873bar),
    .I0(in_40bar),
    .I1(inbar[91])
  );
  //OR U91
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U91 (
    .O(n874),
    .I0(in_8),
    .I1(in_46)
  );
  //AND U91bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U91bar (
    .O(n874bar),
    .I0(in_8bar),
    .I1(in_46bar)
  );
  //OR U92
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U92 (
    .O(n889),
    .I0(n872),
    .I1(n871)
  );
  //AND U92bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U92bar (
    .O(n889bar),
    .I0(n872bar),
    .I1(n871bar)
  );
  //OR U93
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U93 (
    .O(n871),
    .I0(in[117]),
    .I1(n943)
  );
  //AND U93bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U93bar (
    .O(n871bar),
    .I0(inbar[117]),
    .I1(n943bar)
  );
  //OR U94
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U94 (
    .O(n943),
    .I0(n870),
    .I1(n869)
  );
  //AND U94bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U94bar (
    .O(n943bar),
    .I0(n870bar),
    .I1(n869bar)
  );
  //OR U95
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U95 (
    .O(n869),
    .I0(n868),
    .I1(n867)
  );
  //AND U95bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U95bar (
    .O(n869bar),
    .I0(n868bar),
    .I1(n867bar)
  );
  //OR U96
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U96 (
    .O(n867),
    .I0(n866),
    .I1(n865)
  );
  //AND U96bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U96bar (
    .O(n867bar),
    .I0(n866bar),
    .I1(n865bar)
  );
  //OR U97
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U97 (
    .O(n865),
    .I0(n864),
    .I1(n863)
  );
  //AND U97bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U97bar (
    .O(n865bar),
    .I0(n864bar),
    .I1(n863bar)
  );
  //OR U98
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U98 (
    .O(n866),
    .I0(in[108]),
    .I1(n919)
  );
  //AND U98bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U98bar (
    .O(n866bar),
    .I0(inbar[108]),
    .I1(n919bar)
  );
  //OR U99
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U99 (
    .O(n919),
    .I0(n862),
    .I1(n861)
  );
  //AND U99bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U99bar (
    .O(n919bar),
    .I0(n862bar),
    .I1(n861bar)
  );
  //OR U100
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U100 (
    .O(n861),
    .I0(n860),
    .I1(n859)
  );
  //AND U100bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U100bar (
    .O(n861bar),
    .I0(n860bar),
    .I1(n859bar)
  );
  //OR U101
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U101 (
    .O(n859),
    .I0(n858),
    .I1(n857)
  );
  //AND U101bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U101bar (
    .O(n859bar),
    .I0(n858bar),
    .I1(n857bar)
  );
  //OR U102
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U102 (
    .O(n857),
    .I0(in[119]),
    .I1(in[105])
  );
  //AND U102bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U102bar (
    .O(n857bar),
    .I0(inbar[119]),
    .I1(inbar[105])
  );
  //OR U103
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U103 (
    .O(n858),
    .I0(in[186]),
    .I1(in[175])
  );
  //AND U103bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U103bar (
    .O(n858bar),
    .I0(inbar[186]),
    .I1(inbar[175])
  );
  //OR U104
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U104 (
    .O(n860),
    .I0(n856),
    .I1(n855)
  );
  //AND U104bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U104bar (
    .O(n860bar),
    .I0(n856bar),
    .I1(n855bar)
  );
  //OR U105
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U105 (
    .O(n855),
    .I0(in[202]),
    .I1(in[193])
  );
  //AND U105bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U105bar (
    .O(n855bar),
    .I0(inbar[202]),
    .I1(inbar[193])
  );
  //OR U106
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U106 (
    .O(n856),
    .I0(in[225]),
    .I1(in[208])
  );
  //AND U106bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U106bar (
    .O(n856bar),
    .I0(inbar[225]),
    .I1(inbar[208])
  );
  //OR U107
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U107 (
    .O(n862),
    .I0(n854),
    .I1(n853)
  );
  //AND U107bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U107bar (
    .O(n862bar),
    .I0(n854bar),
    .I1(n853bar)
  );
  //OR U108
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U108 (
    .O(n853),
    .I0(n852),
    .I1(n851)
  );
  //AND U108bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U108bar (
    .O(n853bar),
    .I0(n852bar),
    .I1(n851bar)
  );
  //OR U109
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U109 (
    .O(n851),
    .I0(in_1),
    .I1(in[85])
  );
  //AND U109bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U109bar (
    .O(n851bar),
    .I0(in_1bar),
    .I1(inbar[85])
  );
  //OR U110
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U110 (
    .O(n852),
    .I0(in_23),
    .I1(in_19)
  );
  //AND U110bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U110bar (
    .O(n852bar),
    .I0(in_23bar),
    .I1(in_19bar)
  );
  //OR U111
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U111 (
    .O(n854),
    .I0(n850),
    .I1(n849)
  );
  //AND U111bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U111bar (
    .O(n854bar),
    .I0(n850bar),
    .I1(n849bar)
  );
  //OR U112
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U112 (
    .O(n849),
    .I0(in_43),
    .I1(in_33)
  );
  //AND U112bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U112bar (
    .O(n849bar),
    .I0(in_43bar),
    .I1(in_33bar)
  );
  //OR U113
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U113 (
    .O(n850),
    .I0(in_63),
    .I1(in_44)
  );
  //AND U113bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U113bar (
    .O(n850bar),
    .I0(in_63bar),
    .I1(in_44bar)
  );
  //OR U114
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U114 (
    .O(n868),
    .I0(n848),
    .I1(n847)
  );
  //AND U114bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U114bar (
    .O(n868bar),
    .I0(n848bar),
    .I1(n847bar)
  );
  //OR U115
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U115 (
    .O(n847),
    .I0(in[141]),
    .I1(in[112])
  );
  //AND U115bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U115bar (
    .O(n847bar),
    .I0(inbar[141]),
    .I1(inbar[112])
  );
  //OR U116
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U116 (
    .O(n848),
    .I0(in[147]),
    .I1(n846)
  );
  //AND U116bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U116bar (
    .O(n848bar),
    .I0(inbar[147]),
    .I1(n846bar)
  );
  //OR U117
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U117 (
    .O(n846),
    .I0(in[181]),
    .I1(in[167])
  );
  //AND U117bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U117bar (
    .O(n846bar),
    .I0(inbar[181]),
    .I1(inbar[167])
  );
  //OR U118
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U118 (
    .O(n870),
    .I0(n845),
    .I1(n844)
  );
  //AND U118bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U118bar (
    .O(n870bar),
    .I0(n845bar),
    .I1(n844bar)
  );
  //OR U119
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U119 (
    .O(n844),
    .I0(n843),
    .I1(n842)
  );
  //AND U119bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U119bar (
    .O(n844bar),
    .I0(n843bar),
    .I1(n842bar)
  );
  //OR U120
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U120 (
    .O(n842),
    .I0(in[229]),
    .I1(in[201])
  );
  //AND U120bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U120bar (
    .O(n842bar),
    .I0(inbar[229]),
    .I1(inbar[201])
  );
  //OR U121
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U121 (
    .O(n843),
    .I0(in[237]),
    .I1(n841)
  );
  //AND U121bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U121bar (
    .O(n843bar),
    .I0(inbar[237]),
    .I1(n841bar)
  );
  //OR U122
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U122 (
    .O(n841),
    .I0(in[94]),
    .I1(in[253])
  );
  //AND U122bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U122bar (
    .O(n841bar),
    .I0(inbar[94]),
    .I1(inbar[253])
  );
  //OR U123
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U123 (
    .O(n845),
    .I0(n840),
    .I1(n839)
  );
  //AND U123bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U123bar (
    .O(n845bar),
    .I0(n840bar),
    .I1(n839bar)
  );
  //OR U124
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U124 (
    .O(n839),
    .I0(in_21),
    .I1(in[96])
  );
  //AND U124bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U124bar (
    .O(n839bar),
    .I0(in_21bar),
    .I1(inbar[96])
  );
  //OR U125
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U125 (
    .O(n840),
    .I0(in_25),
    .I1(n838)
  );
  //AND U125bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U125bar (
    .O(n840bar),
    .I0(in_25bar),
    .I1(n838bar)
  );
  //OR U126
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U126 (
    .O(n838),
    .I0(in_81),
    .I1(in_45)
  );
  //AND U126bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U126bar (
    .O(n838bar),
    .I0(in_81bar),
    .I1(in_45bar)
  );
  //OR U127
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U127 (
    .O(n891),
    .I0(n837),
    .I1(n836)
  );
  //AND U127bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U127bar (
    .O(n891bar),
    .I0(n837bar),
    .I1(n836bar)
  );
  //OR U128
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U128 (
    .O(n836),
    .I0(in[142]),
    .I1(in[124])
  );
  //AND U128bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U128bar (
    .O(n836bar),
    .I0(inbar[142]),
    .I1(inbar[124])
  );
  //OR U129
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U129 (
    .O(n837),
    .I0(in[150]),
    .I1(n835)
  );
  //AND U129bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U129bar (
    .O(n837bar),
    .I0(inbar[150]),
    .I1(n835bar)
  );
  //OR U130
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U130 (
    .O(n835),
    .I0(in[172]),
    .I1(in[155])
  );
  //AND U130bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U130bar (
    .O(n835bar),
    .I0(inbar[172]),
    .I1(inbar[155])
  );
  //OR U131
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U131 (
    .O(n893),
    .I0(n834),
    .I1(n833)
  );
  //AND U131bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U131bar (
    .O(n893bar),
    .I0(n834bar),
    .I1(n833bar)
  );
  //OR U132
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U132 (
    .O(n833),
    .I0(n832),
    .I1(n831)
  );
  //AND U132bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U132bar (
    .O(n833bar),
    .I0(n832bar),
    .I1(n831bar)
  );
  //OR U133
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U133 (
    .O(n831),
    .I0(in[196]),
    .I1(in[173])
  );
  //AND U133bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U133bar (
    .O(n831bar),
    .I0(inbar[196]),
    .I1(inbar[173])
  );
  //OR U134
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U134 (
    .O(n832),
    .I0(in[222]),
    .I1(n830)
  );
  //AND U134bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U134bar (
    .O(n832bar),
    .I0(inbar[222]),
    .I1(n830bar)
  );
  //OR U135
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U135 (
    .O(n830),
    .I0(in[227]),
    .I1(in[226])
  );
  //AND U135bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U135bar (
    .O(n830bar),
    .I0(inbar[227]),
    .I1(inbar[226])
  );
  //OR U136
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U136 (
    .O(n834),
    .I0(n829),
    .I1(n828)
  );
  //AND U136bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U136bar (
    .O(n834bar),
    .I0(n829bar),
    .I1(n828bar)
  );
  //OR U137
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U137 (
    .O(n828),
    .I0(in[249]),
    .I1(in[231])
  );
  //AND U137bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U137bar (
    .O(n828bar),
    .I0(inbar[249]),
    .I1(inbar[231])
  );
  //OR U138
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U138 (
    .O(n829),
    .I0(in_28),
    .I1(n827)
  );
  //AND U138bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U138bar (
    .O(n829bar),
    .I0(in_28bar),
    .I1(n827bar)
  );
  //OR U139
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U139 (
    .O(n827),
    .I0(in_52),
    .I1(in_47)
  );
  //AND U139bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U139bar (
    .O(n827bar),
    .I0(in_52bar),
    .I1(in_47bar)
  );
  //OR U140
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U140 (
    .O(out[3]),
    .I0(n826),
    .I1(n825)
  );
  //AND U140bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U140bar (
    .O(outbar[3]),
    .I0(n826bar),
    .I1(n825bar)
  );
  //OR U141
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U141 (
    .O(n825),
    .I0(n824),
    .I1(n823)
  );
  //AND U141bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U141bar (
    .O(n825bar),
    .I0(n824bar),
    .I1(n823bar)
  );
  //OR U142
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U142 (
    .O(n823),
    .I0(n822),
    .I1(n821)
  );
  //AND U142bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U142bar (
    .O(n823bar),
    .I0(n822bar),
    .I1(n821bar)
  );
  //OR U143
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U143 (
    .O(n821),
    .I0(n820),
    .I1(n819)
  );
  //AND U143bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U143bar (
    .O(n821bar),
    .I0(n820bar),
    .I1(n819bar)
  );
  //OR U144
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U144 (
    .O(n822),
    .I0(n964),
    .I1(n818)
  );
  //AND U144bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U144bar (
    .O(n822bar),
    .I0(n964bar),
    .I1(n818bar)
  );
  //OR U145
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U145 (
    .O(n818),
    .I0(in[118]),
    .I1(n817)
  );
  //AND U145bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U145bar (
    .O(n818bar),
    .I0(inbar[118]),
    .I1(n817bar)
  );
  //OR U146
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U146 (
    .O(n964),
    .I0(n816),
    .I1(n815)
  );
  //AND U146bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U146bar (
    .O(n964bar),
    .I0(n816bar),
    .I1(n815bar)
  );
  //OR U147
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U147 (
    .O(n815),
    .I0(n814),
    .I1(n813)
  );
  //AND U147bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U147bar (
    .O(n815bar),
    .I0(n814bar),
    .I1(n813bar)
  );
  //OR U148
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U148 (
    .O(n813),
    .I0(n812),
    .I1(n811)
  );
  //AND U148bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U148bar (
    .O(n813bar),
    .I0(n812bar),
    .I1(n811bar)
  );
  //OR U149
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U149 (
    .O(n811),
    .I0(in[122]),
    .I1(in[111])
  );
  //AND U149bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U149bar (
    .O(n811bar),
    .I0(inbar[122]),
    .I1(inbar[111])
  );
  //OR U150
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U150 (
    .O(n812),
    .I0(in[154]),
    .I1(in[151])
  );
  //AND U150bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U150bar (
    .O(n812bar),
    .I0(inbar[154]),
    .I1(inbar[151])
  );
  //OR U151
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U151 (
    .O(n814),
    .I0(n810),
    .I1(n809)
  );
  //AND U151bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U151bar (
    .O(n814bar),
    .I0(n810bar),
    .I1(n809bar)
  );
  //OR U152
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U152 (
    .O(n809),
    .I0(in[187]),
    .I1(in[177])
  );
  //AND U152bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U152bar (
    .O(n809bar),
    .I0(inbar[187]),
    .I1(inbar[177])
  );
  //OR U153
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U153 (
    .O(n810),
    .I0(in[200]),
    .I1(in[192])
  );
  //AND U153bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U153bar (
    .O(n810bar),
    .I0(inbar[200]),
    .I1(inbar[192])
  );
  //OR U154
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U154 (
    .O(n816),
    .I0(n808),
    .I1(n807)
  );
  //AND U154bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U154bar (
    .O(n816bar),
    .I0(n808bar),
    .I1(n807bar)
  );
  //OR U155
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U155 (
    .O(n807),
    .I0(n806),
    .I1(n805)
  );
  //AND U155bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U155bar (
    .O(n807bar),
    .I0(n806bar),
    .I1(n805bar)
  );
  //OR U156
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U156 (
    .O(n805),
    .I0(in[225]),
    .I1(in[207])
  );
  //AND U156bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U156bar (
    .O(n805bar),
    .I0(inbar[225]),
    .I1(inbar[207])
  );
  //OR U157
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U157 (
    .O(n806),
    .I0(in[98]),
    .I1(in[226])
  );
  //AND U157bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U157bar (
    .O(n806bar),
    .I0(inbar[98]),
    .I1(inbar[226])
  );
  //OR U158
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U158 (
    .O(n808),
    .I0(n804),
    .I1(n803)
  );
  //AND U158bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U158bar (
    .O(n808bar),
    .I0(n804bar),
    .I1(n803bar)
  );
  //OR U159
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U159 (
    .O(n803),
    .I0(in_20),
    .I1(in_16)
  );
  //AND U159bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U159bar (
    .O(n803bar),
    .I0(in_20bar),
    .I1(in_16bar)
  );
  //OR U160
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U160 (
    .O(n804),
    .I0(in_55),
    .I1(in_45)
  );
  //AND U160bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U160bar (
    .O(n804bar),
    .I0(in_55bar),
    .I1(in_45bar)
  );
  //OR U161
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U161 (
    .O(n824),
    .I0(n802),
    .I1(n801)
  );
  //AND U161bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U161bar (
    .O(n824bar),
    .I0(n802bar),
    .I1(n801bar)
  );
  //OR U162
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U162 (
    .O(n801),
    .I0(in[162]),
    .I1(in[149])
  );
  //AND U162bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U162bar (
    .O(n801bar),
    .I0(inbar[162]),
    .I1(inbar[149])
  );
  //OR U163
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U163 (
    .O(n802),
    .I0(in[163]),
    .I1(n800)
  );
  //AND U163bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U163bar (
    .O(n802bar),
    .I0(inbar[163]),
    .I1(n800bar)
  );
  //OR U164
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U164 (
    .O(n800),
    .I0(in[191]),
    .I1(in[189])
  );
  //AND U164bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U164bar (
    .O(n800bar),
    .I0(inbar[191]),
    .I1(inbar[189])
  );
  //OR U165
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U165 (
    .O(n826),
    .I0(n799),
    .I1(n798)
  );
  //AND U165bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U165bar (
    .O(n826bar),
    .I0(n799bar),
    .I1(n798bar)
  );
  //OR U166
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U166 (
    .O(n798),
    .I0(n797),
    .I1(n796)
  );
  //AND U166bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U166bar (
    .O(n798bar),
    .I0(n797bar),
    .I1(n796bar)
  );
  //OR U167
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U167 (
    .O(n796),
    .I0(in[212]),
    .I1(in[193])
  );
  //AND U167bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U167bar (
    .O(n796bar),
    .I0(inbar[212]),
    .I1(inbar[193])
  );
  //OR U168
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U168 (
    .O(n797),
    .I0(in[238]),
    .I1(n795)
  );
  //AND U168bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U168bar (
    .O(n797bar),
    .I0(inbar[238]),
    .I1(n795bar)
  );
  //OR U169
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U169 (
    .O(n795),
    .I0(in[88]),
    .I1(in[247])
  );
  //AND U169bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U169bar (
    .O(n795bar),
    .I0(inbar[88]),
    .I1(inbar[247])
  );
  //OR U170
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U170 (
    .O(n799),
    .I0(n794),
    .I1(n793)
  );
  //AND U170bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U170bar (
    .O(n799bar),
    .I0(n794bar),
    .I1(n793bar)
  );
  //OR U171
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U171 (
    .O(n793),
    .I0(in[94]),
    .I1(in[92])
  );
  //AND U171bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U171bar (
    .O(n793bar),
    .I0(inbar[94]),
    .I1(inbar[92])
  );
  //OR U172
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U172 (
    .O(n794),
    .I0(in_52),
    .I1(n792)
  );
  //AND U172bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U172bar (
    .O(n794bar),
    .I0(in_52bar),
    .I1(n792bar)
  );
  //OR U173
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U173 (
    .O(n792),
    .I0(in_70),
    .I1(in_67)
  );
  //AND U173bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U173bar (
    .O(n792bar),
    .I0(in_70bar),
    .I1(in_67bar)
  );
  //OR U174
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U174 (
    .O(out[2]),
    .I0(n791),
    .I1(n790)
  );
  //AND U174bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U174bar (
    .O(outbar[2]),
    .I0(n791bar),
    .I1(n790bar)
  );
  //OR U175
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U175 (
    .O(n790),
    .I0(n789),
    .I1(n788)
  );
  //AND U175bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U175bar (
    .O(n790bar),
    .I0(n789bar),
    .I1(n788bar)
  );
  //OR U176
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U176 (
    .O(n788),
    .I0(n787),
    .I1(n786)
  );
  //AND U176bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U176bar (
    .O(n788bar),
    .I0(n787bar),
    .I1(n786bar)
  );
  //OR U177
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U177 (
    .O(n786),
    .I0(n819),
    .I1(n785)
  );
  //AND U177bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U177bar (
    .O(n786bar),
    .I0(n819bar),
    .I1(n785bar)
  );
  //OR U178
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U178 (
    .O(n819),
    .I0(n784),
    .I1(n783)
  );
  //AND U178bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U178bar (
    .O(n819bar),
    .I0(n784bar),
    .I1(n783bar)
  );
  //OR U179
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U179 (
    .O(n783),
    .I0(n782),
    .I1(n781)
  );
  //AND U179bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U179bar (
    .O(n783bar),
    .I0(n782bar),
    .I1(n781bar)
  );
  //OR U180
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U180 (
    .O(n781),
    .I0(n780),
    .I1(n779)
  );
  //AND U180bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U180bar (
    .O(n781bar),
    .I0(n780bar),
    .I1(n779bar)
  );
  //OR U181
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U181 (
    .O(n779),
    .I0(n962),
    .I1(n778)
  );
  //AND U181bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U181bar (
    .O(n779bar),
    .I0(n962bar),
    .I1(n778bar)
  );
  //OR U182
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U182 (
    .O(n962),
    .I0(n777),
    .I1(n776)
  );
  //AND U182bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U182bar (
    .O(n962bar),
    .I0(n777bar),
    .I1(n776bar)
  );
  //OR U183
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U183 (
    .O(n776),
    .I0(n775),
    .I1(n774)
  );
  //AND U183bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U183bar (
    .O(n776bar),
    .I0(n775bar),
    .I1(n774bar)
  );
  //OR U184
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U184 (
    .O(n774),
    .I0(n773),
    .I1(n772)
  );
  //AND U184bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U184bar (
    .O(n774bar),
    .I0(n773bar),
    .I1(n772bar)
  );
  //OR U185
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U185 (
    .O(n772),
    .I0(in[131]),
    .I1(in[120])
  );
  //AND U185bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U185bar (
    .O(n772bar),
    .I0(inbar[131]),
    .I1(inbar[120])
  );
  //OR U186
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U186 (
    .O(n773),
    .I0(in[153]),
    .I1(in[147])
  );
  //AND U186bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U186bar (
    .O(n773bar),
    .I0(inbar[153]),
    .I1(inbar[147])
  );
  //OR U187
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U187 (
    .O(n775),
    .I0(n771),
    .I1(n770)
  );
  //AND U187bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U187bar (
    .O(n775bar),
    .I0(n771bar),
    .I1(n770bar)
  );
  //OR U188
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U188 (
    .O(n770),
    .I0(in[170]),
    .I1(in[156])
  );
  //AND U188bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U188bar (
    .O(n770bar),
    .I0(inbar[170]),
    .I1(inbar[156])
  );
  //OR U189
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U189 (
    .O(n771),
    .I0(in[223]),
    .I1(in[190])
  );
  //AND U189bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U189bar (
    .O(n771bar),
    .I0(inbar[223]),
    .I1(inbar[190])
  );
  //OR U190
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U190 (
    .O(n777),
    .I0(n769),
    .I1(n768)
  );
  //AND U190bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U190bar (
    .O(n777bar),
    .I0(n769bar),
    .I1(n768bar)
  );
  //OR U191
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U191 (
    .O(n768),
    .I0(n767),
    .I1(n766)
  );
  //AND U191bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U191bar (
    .O(n768bar),
    .I0(n767bar),
    .I1(n766bar)
  );
  //OR U192
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U192 (
    .O(n766),
    .I0(in[236]),
    .I1(in[230])
  );
  //AND U192bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U192bar (
    .O(n766bar),
    .I0(inbar[236]),
    .I1(inbar[230])
  );
  //OR U193
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U193 (
    .O(n767),
    .I0(in[85]),
    .I1(in[240])
  );
  //AND U193bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U193bar (
    .O(n767bar),
    .I0(inbar[85]),
    .I1(inbar[240])
  );
  //OR U194
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U194 (
    .O(n769),
    .I0(n765),
    .I1(n764)
  );
  //AND U194bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U194bar (
    .O(n769bar),
    .I0(n765bar),
    .I1(n764bar)
  );
  //OR U195
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U195 (
    .O(n764),
    .I0(in_12),
    .I1(in[90])
  );
  //AND U195bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U195bar (
    .O(n764bar),
    .I0(in_12bar),
    .I1(inbar[90])
  );
  //OR U196
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U196 (
    .O(n765),
    .I0(in_39),
    .I1(in_28)
  );
  //AND U196bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U196bar (
    .O(n765bar),
    .I0(in_39bar),
    .I1(in_28bar)
  );
  //OR U197
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U197 (
    .O(n780),
    .I0(in[109]),
    .I1(n763)
  );
  //AND U197bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U197bar (
    .O(n780bar),
    .I0(inbar[109]),
    .I1(n763bar)
  );
  //OR U198
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U198 (
    .O(n782),
    .I0(n762),
    .I1(n761)
  );
  //AND U198bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U198bar (
    .O(n782bar),
    .I0(n762bar),
    .I1(n761bar)
  );
  //OR U199
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U199 (
    .O(n761),
    .I0(in[138]),
    .I1(in[129])
  );
  //AND U199bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U199bar (
    .O(n761bar),
    .I0(inbar[138]),
    .I1(inbar[129])
  );
  //OR U200
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U200 (
    .O(n762),
    .I0(in[157]),
    .I1(n760)
  );
  //AND U200bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U200bar (
    .O(n762bar),
    .I0(inbar[157]),
    .I1(n760bar)
  );
  //OR U201
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U201 (
    .O(n760),
    .I0(in[182]),
    .I1(in[167])
  );
  //AND U201bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U201bar (
    .O(n760bar),
    .I0(inbar[182]),
    .I1(inbar[167])
  );
  //OR U202
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U202 (
    .O(n784),
    .I0(n759),
    .I1(n758)
  );
  //AND U202bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U202bar (
    .O(n784bar),
    .I0(n759bar),
    .I1(n758bar)
  );
  //OR U203
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U203 (
    .O(n758),
    .I0(n757),
    .I1(n756)
  );
  //AND U203bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U203bar (
    .O(n758bar),
    .I0(n757bar),
    .I1(n756bar)
  );
  //OR U204
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U204 (
    .O(n756),
    .I0(in[195]),
    .I1(in[184])
  );
  //AND U204bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U204bar (
    .O(n756bar),
    .I0(inbar[195]),
    .I1(inbar[184])
  );
  //OR U205
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U205 (
    .O(n757),
    .I0(in[196]),
    .I1(n755)
  );
  //AND U205bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U205bar (
    .O(n757bar),
    .I0(inbar[196]),
    .I1(n755bar)
  );
  //OR U206
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U206 (
    .O(n755),
    .I0(in[215]),
    .I1(in[209])
  );
  //AND U206bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U206bar (
    .O(n755bar),
    .I0(inbar[215]),
    .I1(inbar[209])
  );
  //OR U207
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U207 (
    .O(n759),
    .I0(n754),
    .I1(n753)
  );
  //AND U207bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U207bar (
    .O(n759bar),
    .I0(n754bar),
    .I1(n753bar)
  );
  //OR U208
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U208 (
    .O(n753),
    .I0(in[93]),
    .I1(in[233])
  );
  //AND U208bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U208bar (
    .O(n753bar),
    .I0(inbar[93]),
    .I1(inbar[233])
  );
  //OR U209
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U209 (
    .O(n754),
    .I0(in_1),
    .I1(n752)
  );
  //AND U209bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U209bar (
    .O(n754bar),
    .I0(in_1bar),
    .I1(n752bar)
  );
  //OR U210
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U210 (
    .O(n752),
    .I0(in_69),
    .I1(in_66)
  );
  //AND U210bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U210bar (
    .O(n752bar),
    .I0(in_69bar),
    .I1(in_66bar)
  );
  //OR U211
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U211 (
    .O(n787),
    .I0(n966),
    .I1(n751)
  );
  //AND U211bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U211bar (
    .O(n787bar),
    .I0(n966bar),
    .I1(n751bar)
  );
  //OR U212
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U212 (
    .O(n751),
    .I0(in[134]),
    .I1(n750)
  );
  //AND U212bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U212bar (
    .O(n751bar),
    .I0(inbar[134]),
    .I1(n750bar)
  );
  //OR U213
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U213 (
    .O(n966),
    .I0(n749),
    .I1(n748)
  );
  //AND U213bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U213bar (
    .O(n966bar),
    .I0(n749bar),
    .I1(n748bar)
  );
  //OR U214
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U214 (
    .O(n748),
    .I0(n747),
    .I1(n746)
  );
  //AND U214bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U214bar (
    .O(n748bar),
    .I0(n747bar),
    .I1(n746bar)
  );
  //OR U215
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U215 (
    .O(n746),
    .I0(n745),
    .I1(n744)
  );
  //AND U215bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U215bar (
    .O(n746bar),
    .I0(n745bar),
    .I1(n744bar)
  );
  //OR U216
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U216 (
    .O(n744),
    .I0(in[136]),
    .I1(in[121])
  );
  //AND U216bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U216bar (
    .O(n744bar),
    .I0(inbar[136]),
    .I1(inbar[121])
  );
  //OR U217
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U217 (
    .O(n745),
    .I0(in[186]),
    .I1(in[174])
  );
  //AND U217bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U217bar (
    .O(n745bar),
    .I0(inbar[186]),
    .I1(inbar[174])
  );
  //OR U218
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U218 (
    .O(n747),
    .I0(n743),
    .I1(n742)
  );
  //AND U218bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U218bar (
    .O(n747bar),
    .I0(n743bar),
    .I1(n742bar)
  );
  //OR U219
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U219 (
    .O(n742),
    .I0(in[198]),
    .I1(in[197])
  );
  //AND U219bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U219bar (
    .O(n742bar),
    .I0(inbar[198]),
    .I1(inbar[197])
  );
  //OR U220
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U220 (
    .O(n743),
    .I0(in[214]),
    .I1(in[199])
  );
  //AND U220bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U220bar (
    .O(n743bar),
    .I0(inbar[214]),
    .I1(inbar[199])
  );
  //OR U221
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U221 (
    .O(n749),
    .I0(n741),
    .I1(n740)
  );
  //AND U221bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U221bar (
    .O(n749bar),
    .I0(n741bar),
    .I1(n740bar)
  );
  //OR U222
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U222 (
    .O(n740),
    .I0(n739),
    .I1(n738)
  );
  //AND U222bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U222bar (
    .O(n740bar),
    .I0(n739bar),
    .I1(n738bar)
  );
  //OR U223
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U223 (
    .O(n738),
    .I0(in[231]),
    .I1(in[220])
  );
  //AND U223bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U223bar (
    .O(n738bar),
    .I0(inbar[231]),
    .I1(inbar[220])
  );
  //OR U224
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U224 (
    .O(n739),
    .I0(in_25),
    .I1(in[245])
  );
  //AND U224bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U224bar (
    .O(n739bar),
    .I0(in_25bar),
    .I1(inbar[245])
  );
  //OR U225
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U225 (
    .O(n741),
    .I0(n737),
    .I1(n736)
  );
  //AND U225bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U225bar (
    .O(n741bar),
    .I0(n737bar),
    .I1(n736bar)
  );
  //OR U226
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U226 (
    .O(n736),
    .I0(in_53),
    .I1(in_29)
  );
  //AND U226bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U226bar (
    .O(n736bar),
    .I0(in_53bar),
    .I1(in_29bar)
  );
  //OR U227
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U227 (
    .O(n737),
    .I0(in_79),
    .I1(in_74)
  );
  //AND U227bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U227bar (
    .O(n737bar),
    .I0(in_79bar),
    .I1(in_74bar)
  );
  //OR U228
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U228 (
    .O(n789),
    .I0(n735),
    .I1(n734)
  );
  //AND U228bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U228bar (
    .O(n789bar),
    .I0(n735bar),
    .I1(n734bar)
  );
  //OR U229
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U229 (
    .O(n734),
    .I0(in[152]),
    .I1(in[140])
  );
  //AND U229bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U229bar (
    .O(n734bar),
    .I0(inbar[152]),
    .I1(inbar[140])
  );
  //OR U230
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U230 (
    .O(n735),
    .I0(in[155]),
    .I1(n733)
  );
  //AND U230bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U230bar (
    .O(n735bar),
    .I0(inbar[155]),
    .I1(n733bar)
  );
  //OR U231
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U231 (
    .O(n733),
    .I0(in[166]),
    .I1(in[165])
  );
  //AND U231bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U231bar (
    .O(n733bar),
    .I0(inbar[166]),
    .I1(inbar[165])
  );
  //OR U232
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U232 (
    .O(n791),
    .I0(n732),
    .I1(n731)
  );
  //AND U232bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U232bar (
    .O(n791bar),
    .I0(n732bar),
    .I1(n731bar)
  );
  //OR U233
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U233 (
    .O(n731),
    .I0(n730),
    .I1(n729)
  );
  //AND U233bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U233bar (
    .O(n731bar),
    .I0(n730bar),
    .I1(n729bar)
  );
  //OR U234
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U234 (
    .O(n729),
    .I0(in[202]),
    .I1(in[185])
  );
  //AND U234bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U234bar (
    .O(n729bar),
    .I0(inbar[202]),
    .I1(inbar[185])
  );
  //OR U235
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U235 (
    .O(n730),
    .I0(in[211]),
    .I1(n728)
  );
  //AND U235bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U235bar (
    .O(n730bar),
    .I0(inbar[211]),
    .I1(n728bar)
  );
  //OR U236
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U236 (
    .O(n728),
    .I0(in[255]),
    .I1(in[253])
  );
  //AND U236bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U236bar (
    .O(n728bar),
    .I0(inbar[255]),
    .I1(inbar[253])
  );
  //OR U237
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U237 (
    .O(n732),
    .I0(n727),
    .I1(n726)
  );
  //AND U237bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U237bar (
    .O(n732bar),
    .I0(n727bar),
    .I1(n726bar)
  );
  //OR U238
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U238 (
    .O(n726),
    .I0(in_35),
    .I1(in_15)
  );
  //AND U238bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U238bar (
    .O(n726bar),
    .I0(in_35bar),
    .I1(in_15bar)
  );
  //OR U239
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U239 (
    .O(n727),
    .I0(in_36),
    .I1(n725)
  );
  //AND U239bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U239bar (
    .O(n727bar),
    .I0(in_36bar),
    .I1(n725bar)
  );
  //OR U240
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U240 (
    .O(n725),
    .I0(in_48),
    .I1(in_40)
  );
  //AND U240bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U240bar (
    .O(n725bar),
    .I0(in_48bar),
    .I1(in_40bar)
  );
  //OR U241
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U241 (
    .O(out[1]),
    .I0(n724),
    .I1(n723)
  );
  //AND U241bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U241bar (
    .O(outbar[1]),
    .I0(n724bar),
    .I1(n723bar)
  );
  //OR U242
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U242 (
    .O(n723),
    .I0(n722),
    .I1(n721)
  );
  //AND U242bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U242bar (
    .O(n723bar),
    .I0(n722bar),
    .I1(n721bar)
  );
  //OR U243
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U243 (
    .O(n721),
    .I0(n720),
    .I1(n719)
  );
  //AND U243bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U243bar (
    .O(n721bar),
    .I0(n720bar),
    .I1(n719bar)
  );
  //OR U244
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U244 (
    .O(n719),
    .I0(n921),
    .I1(n887)
  );
  //AND U244bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U244bar (
    .O(n719bar),
    .I0(n921bar),
    .I1(n887bar)
  );
  //OR U245
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U245 (
    .O(n887),
    .I0(n718),
    .I1(n717)
  );
  //AND U245bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U245bar (
    .O(n887bar),
    .I0(n718bar),
    .I1(n717bar)
  );
  //OR U246
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U246 (
    .O(n717),
    .I0(n716),
    .I1(n715)
  );
  //AND U246bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U246bar (
    .O(n717bar),
    .I0(n716bar),
    .I1(n715bar)
  );
  //OR U247
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U247 (
    .O(n715),
    .I0(n714),
    .I1(n713)
  );
  //AND U247bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U247bar (
    .O(n715bar),
    .I0(n714bar),
    .I1(n713bar)
  );
  //OR U248
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U248 (
    .O(n713),
    .I0(in[116]),
    .I1(in[110])
  );
  //AND U248bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U248bar (
    .O(n713bar),
    .I0(inbar[116]),
    .I1(inbar[110])
  );
  //OR U249
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U249 (
    .O(n714),
    .I0(in[133]),
    .I1(in[130])
  );
  //AND U249bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U249bar (
    .O(n714bar),
    .I0(inbar[133]),
    .I1(inbar[130])
  );
  //OR U250
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U250 (
    .O(n716),
    .I0(n712),
    .I1(n711)
  );
  //AND U250bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U250bar (
    .O(n716bar),
    .I0(n712bar),
    .I1(n711bar)
  );
  //OR U251
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U251 (
    .O(n711),
    .I0(in[203]),
    .I1(in[135])
  );
  //AND U251bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U251bar (
    .O(n711bar),
    .I0(inbar[203]),
    .I1(inbar[135])
  );
  //OR U252
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U252 (
    .O(n712),
    .I0(in[232]),
    .I1(in[223])
  );
  //AND U252bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U252bar (
    .O(n712bar),
    .I0(inbar[232]),
    .I1(inbar[223])
  );
  //OR U253
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U253 (
    .O(n718),
    .I0(n710),
    .I1(n709)
  );
  //AND U253bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U253bar (
    .O(n718bar),
    .I0(n710bar),
    .I1(n709bar)
  );
  //OR U254
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U254 (
    .O(n709),
    .I0(n708),
    .I1(n707)
  );
  //AND U254bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U254bar (
    .O(n709bar),
    .I0(n708bar),
    .I1(n707bar)
  );
  //OR U255
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U255 (
    .O(n707),
    .I0(in[255]),
    .I1(in[233])
  );
  //AND U255bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U255bar (
    .O(n707bar),
    .I0(inbar[255]),
    .I1(inbar[233])
  );
  //OR U256
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U256 (
    .O(n708),
    .I0(in_53),
    .I1(in_34)
  );
  //AND U256bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U256bar (
    .O(n708bar),
    .I0(in_53bar),
    .I1(in_34bar)
  );
  //OR U257
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U257 (
    .O(n710),
    .I0(n706),
    .I1(n705)
  );
  //AND U257bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U257bar (
    .O(n710bar),
    .I0(n706bar),
    .I1(n705bar)
  );
  //OR U258
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U258 (
    .O(n705),
    .I0(in_57),
    .I1(in_55)
  );
  //AND U258bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U258bar (
    .O(n705bar),
    .I0(in_57bar),
    .I1(in_55bar)
  );
  //OR U259
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U259 (
    .O(n706),
    .I0(in_68),
    .I1(in_67)
  );
  //AND U259bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U259bar (
    .O(n706bar),
    .I0(in_68bar),
    .I1(in_67bar)
  );
  //OR U260
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U260 (
    .O(n921),
    .I0(n704),
    .I1(n703)
  );
  //AND U260bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U260bar (
    .O(n921bar),
    .I0(n704bar),
    .I1(n703bar)
  );
  //OR U261
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U261 (
    .O(n703),
    .I0(n702),
    .I1(n701)
  );
  //AND U261bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U261bar (
    .O(n703bar),
    .I0(n702bar),
    .I1(n701bar)
  );
  //OR U262
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U262 (
    .O(n701),
    .I0(n700),
    .I1(n699)
  );
  //AND U262bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U262bar (
    .O(n701bar),
    .I0(n700bar),
    .I1(n699bar)
  );
  //OR U263
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U263 (
    .O(n699),
    .I0(n944),
    .I1(n872)
  );
  //AND U263bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U263bar (
    .O(n699bar),
    .I0(n944bar),
    .I1(n872bar)
  );
  //OR U264
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U264 (
    .O(n872),
    .I0(n698),
    .I1(n697)
  );
  //AND U264bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U264bar (
    .O(n872bar),
    .I0(n698bar),
    .I1(n697bar)
  );
  //OR U265
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U265 (
    .O(n697),
    .I0(n696),
    .I1(n695)
  );
  //AND U265bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U265bar (
    .O(n697bar),
    .I0(n696bar),
    .I1(n695bar)
  );
  //OR U266
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U266 (
    .O(n695),
    .I0(n694),
    .I1(n693)
  );
  //AND U266bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U266bar (
    .O(n695bar),
    .I0(n694bar),
    .I1(n693bar)
  );
  //OR U267
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U267 (
    .O(n693),
    .I0(in[121]),
    .I1(in[102])
  );
  //AND U267bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U267bar (
    .O(n693bar),
    .I0(inbar[121]),
    .I1(inbar[102])
  );
  //OR U268
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U268 (
    .O(n694),
    .I0(in[162]),
    .I1(in[161])
  );
  //AND U268bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U268bar (
    .O(n694bar),
    .I0(inbar[162]),
    .I1(inbar[161])
  );
  //OR U269
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U269 (
    .O(n696),
    .I0(n692),
    .I1(n691)
  );
  //AND U269bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U269bar (
    .O(n696bar),
    .I0(n692bar),
    .I1(n691bar)
  );
  //OR U270
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U270 (
    .O(n691),
    .I0(in[192]),
    .I1(in[178])
  );
  //AND U270bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U270bar (
    .O(n691bar),
    .I0(inbar[192]),
    .I1(inbar[178])
  );
  //OR U271
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U271 (
    .O(n692),
    .I0(in[244]),
    .I1(in[209])
  );
  //AND U271bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U271bar (
    .O(n692bar),
    .I0(inbar[244]),
    .I1(inbar[209])
  );
  //OR U272
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U272 (
    .O(n698),
    .I0(n690),
    .I1(n689)
  );
  //AND U272bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U272bar (
    .O(n698bar),
    .I0(n690bar),
    .I1(n689bar)
  );
  //OR U273
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U273 (
    .O(n689),
    .I0(n688),
    .I1(n687)
  );
  //AND U273bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U273bar (
    .O(n689bar),
    .I0(n688bar),
    .I1(n687bar)
  );
  //OR U274
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U274 (
    .O(n687),
    .I0(in[90]),
    .I1(in[254])
  );
  //AND U274bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U274bar (
    .O(n687bar),
    .I0(inbar[90]),
    .I1(inbar[254])
  );
  //OR U275
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U275 (
    .O(n688),
    .I0(in_36),
    .I1(in_32)
  );
  //AND U275bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U275bar (
    .O(n688bar),
    .I0(in_36bar),
    .I1(in_32bar)
  );
  //OR U276
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U276 (
    .O(n690),
    .I0(n686),
    .I1(n685)
  );
  //AND U276bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U276bar (
    .O(n690bar),
    .I0(n686bar),
    .I1(n685bar)
  );
  //OR U277
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U277 (
    .O(n685),
    .I0(in_62),
    .I1(in_37)
  );
  //AND U277bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U277bar (
    .O(n685bar),
    .I0(in_62bar),
    .I1(in_37bar)
  );
  //OR U278
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U278 (
    .O(n686),
    .I0(in_75),
    .I1(in_73)
  );
  //AND U278bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U278bar (
    .O(n686bar),
    .I0(in_75bar),
    .I1(in_73bar)
  );
  //OR U279
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U279 (
    .O(n944),
    .I0(n684),
    .I1(n683)
  );
  //AND U279bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U279bar (
    .O(n944bar),
    .I0(n684bar),
    .I1(n683bar)
  );
  //OR U280
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U280 (
    .O(n683),
    .I0(n682),
    .I1(n681)
  );
  //AND U280bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U280bar (
    .O(n683bar),
    .I0(n682bar),
    .I1(n681bar)
  );
  //OR U281
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U281 (
    .O(n681),
    .I0(n680),
    .I1(n679)
  );
  //AND U281bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U281bar (
    .O(n681bar),
    .I0(n680bar),
    .I1(n679bar)
  );
  //OR U282
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U282 (
    .O(n679),
    .I0(in[171]),
    .I1(in[153])
  );
  //AND U282bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U282bar (
    .O(n679bar),
    .I0(inbar[171]),
    .I1(inbar[153])
  );
  //OR U283
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U283 (
    .O(n680),
    .I0(in[187]),
    .I1(in[176])
  );
  //AND U283bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U283bar (
    .O(n680bar),
    .I0(inbar[187]),
    .I1(inbar[176])
  );
  //OR U284
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U284 (
    .O(n682),
    .I0(n678),
    .I1(n677)
  );
  //AND U284bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U284bar (
    .O(n682bar),
    .I0(n678bar),
    .I1(n677bar)
  );
  //OR U285
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U285 (
    .O(n677),
    .I0(in[245]),
    .I1(in[211])
  );
  //AND U285bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U285bar (
    .O(n677bar),
    .I0(inbar[245]),
    .I1(inbar[211])
  );
  //OR U286
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U286 (
    .O(n678),
    .I0(in[97]),
    .I1(in[88])
  );
  //AND U286bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U286bar (
    .O(n678bar),
    .I0(inbar[97]),
    .I1(inbar[88])
  );
  //OR U287
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U287 (
    .O(n684),
    .I0(n676),
    .I1(n675)
  );
  //AND U287bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U287bar (
    .O(n684bar),
    .I0(n676bar),
    .I1(n675bar)
  );
  //OR U288
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U288 (
    .O(n675),
    .I0(n674),
    .I1(n673)
  );
  //AND U288bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U288bar (
    .O(n675bar),
    .I0(n674bar),
    .I1(n673bar)
  );
  //OR U289
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U289 (
    .O(n673),
    .I0(in_10),
    .I1(in_0)
  );
  //AND U289bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U289bar (
    .O(n673bar),
    .I0(in_10bar),
    .I1(in_0bar)
  );
  //OR U290
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U290 (
    .O(n674),
    .I0(in_59),
    .I1(in_5)
  );
  //AND U290bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U290bar (
    .O(n674bar),
    .I0(in_59bar),
    .I1(in_5bar)
  );
  //OR U291
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U291 (
    .O(n676),
    .I0(n672),
    .I1(n671)
  );
  //AND U291bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U291bar (
    .O(n676bar),
    .I0(n672bar),
    .I1(n671bar)
  );
  //OR U292
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U292 (
    .O(n671),
    .I0(in_60),
    .I1(in_6)
  );
  //AND U292bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U292bar (
    .O(n671bar),
    .I0(in_60bar),
    .I1(in_6bar)
  );
  //OR U293
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U293 (
    .O(n672),
    .I0(in_77),
    .I1(in_69)
  );
  //AND U293bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U293bar (
    .O(n672bar),
    .I0(in_77bar),
    .I1(in_69bar)
  );
  //OR U294
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U294 (
    .O(n700),
    .I0(in[113]),
    .I1(n864)
  );
  //AND U294bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U294bar (
    .O(n700bar),
    .I0(inbar[113]),
    .I1(n864bar)
  );
  //OR U295
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U295 (
    .O(n864),
    .I0(n670),
    .I1(n669)
  );
  //AND U295bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U295bar (
    .O(n864bar),
    .I0(n670bar),
    .I1(n669bar)
  );
  //OR U296
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U296 (
    .O(n669),
    .I0(n668),
    .I1(n667)
  );
  //AND U296bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U296bar (
    .O(n669bar),
    .I0(n668bar),
    .I1(n667bar)
  );
  //OR U297
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U297 (
    .O(n667),
    .I0(n666),
    .I1(n665)
  );
  //AND U297bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U297bar (
    .O(n667bar),
    .I0(n666bar),
    .I1(n665bar)
  );
  //OR U298
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U298 (
    .O(n665),
    .I0(in[125]),
    .I1(in[107])
  );
  //AND U298bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U298bar (
    .O(n665bar),
    .I0(inbar[125]),
    .I1(inbar[107])
  );
  //OR U299
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U299 (
    .O(n666),
    .I0(in[138]),
    .I1(in[126])
  );
  //AND U299bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U299bar (
    .O(n666bar),
    .I0(inbar[138]),
    .I1(inbar[126])
  );
  //OR U300
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U300 (
    .O(n668),
    .I0(n664),
    .I1(n663)
  );
  //AND U300bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U300bar (
    .O(n668bar),
    .I0(n664bar),
    .I1(n663bar)
  );
  //OR U301
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U301 (
    .O(n663),
    .I0(in[189]),
    .I1(in[143])
  );
  //AND U301bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U301bar (
    .O(n663bar),
    .I0(inbar[189]),
    .I1(inbar[143])
  );
  //OR U302
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U302 (
    .O(n664),
    .I0(in[99]),
    .I1(in[214])
  );
  //AND U302bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U302bar (
    .O(n664bar),
    .I0(inbar[99]),
    .I1(inbar[214])
  );
  //OR U303
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U303 (
    .O(n670),
    .I0(n662),
    .I1(n661)
  );
  //AND U303bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U303bar (
    .O(n670bar),
    .I0(n662bar),
    .I1(n661bar)
  );
  //OR U304
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U304 (
    .O(n661),
    .I0(n660),
    .I1(n659)
  );
  //AND U304bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U304bar (
    .O(n661bar),
    .I0(n660bar),
    .I1(n659bar)
  );
  //OR U305
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U305 (
    .O(n659),
    .I0(in_15),
    .I1(in_12)
  );
  //AND U305bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U305bar (
    .O(n659bar),
    .I0(in_15bar),
    .I1(in_12bar)
  );
  //OR U306
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U306 (
    .O(n660),
    .I0(in_20),
    .I1(in_2)
  );
  //AND U306bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U306bar (
    .O(n660bar),
    .I0(in_20bar),
    .I1(in_2bar)
  );
  //OR U307
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U307 (
    .O(n662),
    .I0(n658),
    .I1(n657)
  );
  //AND U307bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U307bar (
    .O(n662bar),
    .I0(n658bar),
    .I1(n657bar)
  );
  //OR U308
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U308 (
    .O(n657),
    .I0(in_30),
    .I1(in_3)
  );
  //AND U308bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U308bar (
    .O(n657bar),
    .I0(in_30bar),
    .I1(in_3bar)
  );
  //OR U309
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U309 (
    .O(n658),
    .I0(in_4),
    .I1(in_38)
  );
  //AND U309bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U309bar (
    .O(n658bar),
    .I0(in_4bar),
    .I1(in_38bar)
  );
  //OR U310
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U310 (
    .O(n702),
    .I0(n656),
    .I1(n655)
  );
  //AND U310bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U310bar (
    .O(n702bar),
    .I0(n656bar),
    .I1(n655bar)
  );
  //OR U311
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U311 (
    .O(n655),
    .I0(in[148]),
    .I1(in[137])
  );
  //AND U311bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U311bar (
    .O(n655bar),
    .I0(inbar[148]),
    .I1(inbar[137])
  );
  //OR U312
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U312 (
    .O(n656),
    .I0(in[149]),
    .I1(n654)
  );
  //AND U312bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U312bar (
    .O(n656bar),
    .I0(inbar[149]),
    .I1(n654bar)
  );
  //OR U313
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U313 (
    .O(n654),
    .I0(in[195]),
    .I1(in[190])
  );
  //AND U313bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U313bar (
    .O(n654bar),
    .I0(inbar[195]),
    .I1(inbar[190])
  );
  //OR U314
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U314 (
    .O(n704),
    .I0(n653),
    .I1(n652)
  );
  //AND U314bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U314bar (
    .O(n704bar),
    .I0(n653bar),
    .I1(n652bar)
  );
  //OR U315
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U315 (
    .O(n652),
    .I0(n651),
    .I1(n650)
  );
  //AND U315bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U315bar (
    .O(n652bar),
    .I0(n651bar),
    .I1(n650bar)
  );
  //OR U316
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U316 (
    .O(n650),
    .I0(in[98]),
    .I1(in[197])
  );
  //AND U316bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U316bar (
    .O(n650bar),
    .I0(inbar[98]),
    .I1(inbar[197])
  );
  //OR U317
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U317 (
    .O(n651),
    .I0(in_11),
    .I1(n649)
  );
  //AND U317bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U317bar (
    .O(n651bar),
    .I0(in_11bar),
    .I1(n649bar)
  );
  //OR U318
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U318 (
    .O(n649),
    .I0(in_26),
    .I1(in_14)
  );
  //AND U318bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U318bar (
    .O(n649bar),
    .I0(in_26bar),
    .I1(in_14bar)
  );
  //OR U319
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U319 (
    .O(n653),
    .I0(n648),
    .I1(n647)
  );
  //AND U319bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U319bar (
    .O(n653bar),
    .I0(n648bar),
    .I1(n647bar)
  );
  //OR U320
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U320 (
    .O(n647),
    .I0(in_35),
    .I1(in_27)
  );
  //AND U320bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U320bar (
    .O(n647bar),
    .I0(in_35bar),
    .I1(in_27bar)
  );
  //OR U321
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U321 (
    .O(n648),
    .I0(in_50),
    .I1(n646)
  );
  //AND U321bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U321bar (
    .O(n648bar),
    .I0(in_50bar),
    .I1(n646bar)
  );
  //OR U322
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U322 (
    .O(n646),
    .I0(in_78),
    .I1(in_61)
  );
  //AND U322bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U322bar (
    .O(n646bar),
    .I0(in_78bar),
    .I1(in_61bar)
  );
  //OR U323
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U323 (
    .O(n720),
    .I0(n942),
    .I1(n645)
  );
  //AND U323bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U323bar (
    .O(n720bar),
    .I0(n942bar),
    .I1(n645bar)
  );
  //OR U324
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U324 (
    .O(n645),
    .I0(in[106]),
    .I1(n863)
  );
  //AND U324bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U324bar (
    .O(n645bar),
    .I0(inbar[106]),
    .I1(n863bar)
  );
  //OR U325
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U325 (
    .O(n863),
    .I0(n644),
    .I1(n643)
  );
  //AND U325bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U325bar (
    .O(n863bar),
    .I0(n644bar),
    .I1(n643bar)
  );
  //OR U326
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U326 (
    .O(n643),
    .I0(n642),
    .I1(n641)
  );
  //AND U326bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U326bar (
    .O(n643bar),
    .I0(n642bar),
    .I1(n641bar)
  );
  //OR U327
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U327 (
    .O(n641),
    .I0(n640),
    .I1(n639)
  );
  //AND U327bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U327bar (
    .O(n641bar),
    .I0(n640bar),
    .I1(n639bar)
  );
  //OR U328
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U328 (
    .O(n639),
    .I0(in[127]),
    .I1(in[122])
  );
  //AND U328bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U328bar (
    .O(n639bar),
    .I0(inbar[127]),
    .I1(inbar[122])
  );
  //OR U329
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U329 (
    .O(n640),
    .I0(in[156]),
    .I1(in[132])
  );
  //AND U329bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U329bar (
    .O(n640bar),
    .I0(inbar[156]),
    .I1(inbar[132])
  );
  //OR U330
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U330 (
    .O(n642),
    .I0(n638),
    .I1(n637)
  );
  //AND U330bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U330bar (
    .O(n642bar),
    .I0(n638bar),
    .I1(n637bar)
  );
  //OR U331
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U331 (
    .O(n637),
    .I0(in[159]),
    .I1(in[157])
  );
  //AND U331bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U331bar (
    .O(n637bar),
    .I0(inbar[159]),
    .I1(inbar[157])
  );
  //OR U332
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U332 (
    .O(n638),
    .I0(in[185]),
    .I1(in[169])
  );
  //AND U332bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U332bar (
    .O(n638bar),
    .I0(inbar[185]),
    .I1(inbar[169])
  );
  //OR U333
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U333 (
    .O(n644),
    .I0(n636),
    .I1(n635)
  );
  //AND U333bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U333bar (
    .O(n644bar),
    .I0(n636bar),
    .I1(n635bar)
  );
  //OR U334
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U334 (
    .O(n635),
    .I0(n634),
    .I1(n633)
  );
  //AND U334bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U334bar (
    .O(n635bar),
    .I0(n634bar),
    .I1(n633bar)
  );
  //OR U335
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U335 (
    .O(n633),
    .I0(in[239]),
    .I1(in[218])
  );
  //AND U335bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U335bar (
    .O(n633bar),
    .I0(inbar[239]),
    .I1(inbar[218])
  );
  //OR U336
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U336 (
    .O(n634),
    .I0(in_13),
    .I1(in[87])
  );
  //AND U336bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U336bar (
    .O(n634bar),
    .I0(in_13bar),
    .I1(inbar[87])
  );
  //OR U337
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U337 (
    .O(n636),
    .I0(n632),
    .I1(n631)
  );
  //AND U337bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U337bar (
    .O(n636bar),
    .I0(n632bar),
    .I1(n631bar)
  );
  //OR U338
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U338 (
    .O(n631),
    .I0(in_72),
    .I1(in_70)
  );
  //AND U338bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U338bar (
    .O(n631bar),
    .I0(in_72bar),
    .I1(in_70bar)
  );
  //OR U339
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U339 (
    .O(n632),
    .I0(in_80),
    .I1(in_74)
  );
  //AND U339bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U339bar (
    .O(n632bar),
    .I0(in_80bar),
    .I1(in_74bar)
  );
  //OR U340
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U340 (
    .O(n942),
    .I0(n630),
    .I1(n629)
  );
  //AND U340bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U340bar (
    .O(n942bar),
    .I0(n630bar),
    .I1(n629bar)
  );
  //OR U341
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U341 (
    .O(n629),
    .I0(n628),
    .I1(n627)
  );
  //AND U341bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U341bar (
    .O(n629bar),
    .I0(n628bar),
    .I1(n627bar)
  );
  //OR U342
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U342 (
    .O(n627),
    .I0(n626),
    .I1(n625)
  );
  //AND U342bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U342bar (
    .O(n627bar),
    .I0(n626bar),
    .I1(n625bar)
  );
  //OR U343
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U343 (
    .O(n625),
    .I0(in[146]),
    .I1(in[100])
  );
  //AND U343bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U343bar (
    .O(n625bar),
    .I0(inbar[146]),
    .I1(inbar[100])
  );
  //OR U344
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U344 (
    .O(n626),
    .I0(in[168]),
    .I1(in[152])
  );
  //AND U344bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U344bar (
    .O(n626bar),
    .I0(inbar[168]),
    .I1(inbar[152])
  );
  //OR U345
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U345 (
    .O(n628),
    .I0(n624),
    .I1(n623)
  );
  //AND U345bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U345bar (
    .O(n628bar),
    .I0(n624bar),
    .I1(n623bar)
  );
  //OR U346
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U346 (
    .O(n623),
    .I0(in[199]),
    .I1(in[182])
  );
  //AND U346bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U346bar (
    .O(n623bar),
    .I0(inbar[199]),
    .I1(inbar[182])
  );
  //OR U347
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U347 (
    .O(n624),
    .I0(in[236]),
    .I1(in[204])
  );
  //AND U347bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U347bar (
    .O(n624bar),
    .I0(inbar[236]),
    .I1(inbar[204])
  );
  //OR U348
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U348 (
    .O(n630),
    .I0(n622),
    .I1(n621)
  );
  //AND U348bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U348bar (
    .O(n630bar),
    .I0(n622bar),
    .I1(n621bar)
  );
  //OR U349
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U349 (
    .O(n621),
    .I0(n620),
    .I1(n619)
  );
  //AND U349bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U349bar (
    .O(n621bar),
    .I0(n620bar),
    .I1(n619bar)
  );
  //OR U350
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U350 (
    .O(n619),
    .I0(in[89]),
    .I1(in[246])
  );
  //AND U350bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U350bar (
    .O(n619bar),
    .I0(inbar[89]),
    .I1(inbar[246])
  );
  //OR U351
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U351 (
    .O(n620),
    .I0(in[95]),
    .I1(in[92])
  );
  //AND U351bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U351bar (
    .O(n620bar),
    .I0(inbar[95]),
    .I1(inbar[92])
  );
  //OR U352
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U352 (
    .O(n622),
    .I0(n618),
    .I1(n617)
  );
  //AND U352bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U352bar (
    .O(n622bar),
    .I0(n618bar),
    .I1(n617bar)
  );
  //OR U353
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U353 (
    .O(n617),
    .I0(in_22),
    .I1(in_16)
  );
  //AND U353bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U353bar (
    .O(n617bar),
    .I0(in_22bar),
    .I1(in_16bar)
  );
  //OR U354
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U354 (
    .O(n618),
    .I0(in_51),
    .I1(in_49)
  );
  //AND U354bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U354bar (
    .O(n618bar),
    .I0(in_51bar),
    .I1(in_49bar)
  );
  //OR U355
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U355 (
    .O(n722),
    .I0(n616),
    .I1(n615)
  );
  //AND U355bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U355bar (
    .O(n722bar),
    .I0(n616bar),
    .I1(n615bar)
  );
  //OR U356
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U356 (
    .O(n615),
    .I0(in[158]),
    .I1(in[115])
  );
  //AND U356bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U356bar (
    .O(n615bar),
    .I0(inbar[158]),
    .I1(inbar[115])
  );
  //OR U357
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U357 (
    .O(n616),
    .I0(in[163]),
    .I1(n614)
  );
  //AND U357bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U357bar (
    .O(n616bar),
    .I0(inbar[163]),
    .I1(n614bar)
  );
  //OR U358
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U358 (
    .O(n614),
    .I0(in[206]),
    .I1(in[165])
  );
  //AND U358bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U358bar (
    .O(n614bar),
    .I0(inbar[206]),
    .I1(inbar[165])
  );
  //OR U359
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U359 (
    .O(n724),
    .I0(n613),
    .I1(n612)
  );
  //AND U359bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U359bar (
    .O(n724bar),
    .I0(n613bar),
    .I1(n612bar)
  );
  //OR U360
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U360 (
    .O(n612),
    .I0(n611),
    .I1(n610)
  );
  //AND U360bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U360bar (
    .O(n612bar),
    .I0(n611bar),
    .I1(n610bar)
  );
  //OR U361
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U361 (
    .O(n610),
    .I0(in[213]),
    .I1(in[207])
  );
  //AND U361bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U361bar (
    .O(n610bar),
    .I0(inbar[213]),
    .I1(inbar[207])
  );
  //OR U362
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U362 (
    .O(n611),
    .I0(in[215]),
    .I1(n609)
  );
  //AND U362bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U362bar (
    .O(n611bar),
    .I0(inbar[215]),
    .I1(n609bar)
  );
  //OR U363
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U363 (
    .O(n609),
    .I0(in[230]),
    .I1(in[220])
  );
  //AND U363bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U363bar (
    .O(n609bar),
    .I0(inbar[230]),
    .I1(inbar[220])
  );
  //OR U364
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U364 (
    .O(n613),
    .I0(n608),
    .I1(n607)
  );
  //AND U364bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U364bar (
    .O(n613bar),
    .I0(n608bar),
    .I1(n607bar)
  );
  //OR U365
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U365 (
    .O(n607),
    .I0(in[251]),
    .I1(in[234])
  );
  //AND U365bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U365bar (
    .O(n607bar),
    .I0(inbar[251]),
    .I1(inbar[234])
  );
  //OR U366
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U366 (
    .O(n608),
    .I0(in_17),
    .I1(n606)
  );
  //AND U366bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U366bar (
    .O(n608bar),
    .I0(in_17bar),
    .I1(n606bar)
  );
  //OR U367
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U367 (
    .O(n606),
    .I0(in_65),
    .I1(in_56)
  );
  //AND U367bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U367bar (
    .O(n606bar),
    .I0(in_65bar),
    .I1(in_56bar)
  );
  //OR U368
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U368 (
    .O(out[0]),
    .I0(n605),
    .I1(n604)
  );
  //AND U368bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U368bar (
    .O(outbar[0]),
    .I0(n605bar),
    .I1(n604bar)
  );
  //OR U369
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U369 (
    .O(n604),
    .I0(n603),
    .I1(n602)
  );
  //AND U369bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U369bar (
    .O(n604bar),
    .I0(n603bar),
    .I1(n602bar)
  );
  //OR U370
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U370 (
    .O(n602),
    .I0(n601),
    .I1(n600)
  );
  //AND U370bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U370bar (
    .O(n602bar),
    .I0(n601bar),
    .I1(n600bar)
  );
  //OR U371
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U371 (
    .O(n600),
    .I0(n820),
    .I1(n785)
  );
  //AND U371bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U371bar (
    .O(n600bar),
    .I0(n820bar),
    .I1(n785bar)
  );
  //OR U372
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U372 (
    .O(n785),
    .I0(n599),
    .I1(n598)
  );
  //AND U372bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U372bar (
    .O(n785bar),
    .I0(n599bar),
    .I1(n598bar)
  );
  //OR U373
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U373 (
    .O(n598),
    .I0(n597),
    .I1(n596)
  );
  //AND U373bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U373bar (
    .O(n598bar),
    .I0(n597bar),
    .I1(n596bar)
  );
  //OR U374
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U374 (
    .O(n596),
    .I0(n595),
    .I1(n594)
  );
  //AND U374bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U374bar (
    .O(n596bar),
    .I0(n595bar),
    .I1(n594bar)
  );
  //OR U375
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U375 (
    .O(n594),
    .I0(in[135]),
    .I1(in[104])
  );
  //AND U375bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U375bar (
    .O(n594bar),
    .I0(inbar[135]),
    .I1(inbar[104])
  );
  //OR U376
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U376 (
    .O(n595),
    .I0(in[188]),
    .I1(in[178])
  );
  //AND U376bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U376bar (
    .O(n595bar),
    .I0(inbar[188]),
    .I1(inbar[178])
  );
  //OR U377
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U377 (
    .O(n597),
    .I0(n593),
    .I1(n592)
  );
  //AND U377bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U377bar (
    .O(n597bar),
    .I0(n593bar),
    .I1(n592bar)
  );
  //OR U378
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U378 (
    .O(n592),
    .I0(in[217]),
    .I1(in[194])
  );
  //AND U378bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U378bar (
    .O(n592bar),
    .I0(inbar[217]),
    .I1(inbar[194])
  );
  //OR U379
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U379 (
    .O(n593),
    .I0(in[237]),
    .I1(in[218])
  );
  //AND U379bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U379bar (
    .O(n593bar),
    .I0(inbar[237]),
    .I1(inbar[218])
  );
  //OR U380
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U380 (
    .O(n599),
    .I0(n591),
    .I1(n590)
  );
  //AND U380bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U380bar (
    .O(n599bar),
    .I0(n591bar),
    .I1(n590bar)
  );
  //OR U381
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U381 (
    .O(n590),
    .I0(n589),
    .I1(n588)
  );
  //AND U381bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U381bar (
    .O(n590bar),
    .I0(n589bar),
    .I1(n588bar)
  );
  //OR U382
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U382 (
    .O(n588),
    .I0(in_2),
    .I1(in_10)
  );
  //AND U382bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U382bar (
    .O(n588bar),
    .I0(in_2bar),
    .I1(in_10bar)
  );
  //OR U383
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U383 (
    .O(n589),
    .I0(in_47),
    .I1(in_22)
  );
  //AND U383bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U383bar (
    .O(n589bar),
    .I0(in_47bar),
    .I1(in_22bar)
  );
  //OR U384
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U384 (
    .O(n591),
    .I0(n587),
    .I1(n586)
  );
  //AND U384bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U384bar (
    .O(n591bar),
    .I0(n587bar),
    .I1(n586bar)
  );
  //OR U385
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U385 (
    .O(n586),
    .I0(in_56),
    .I1(in_54)
  );
  //AND U385bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U385bar (
    .O(n586bar),
    .I0(in_56bar),
    .I1(in_54bar)
  );
  //OR U386
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U386 (
    .O(n587),
    .I0(in_63),
    .I1(in_61)
  );
  //AND U386bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U386bar (
    .O(n587bar),
    .I0(in_63bar),
    .I1(in_61bar)
  );
  //OR U387
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U387 (
    .O(n820),
    .I0(n585),
    .I1(n584)
  );
  //AND U387bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U387bar (
    .O(n820bar),
    .I0(n585bar),
    .I1(n584bar)
  );
  //OR U388
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U388 (
    .O(n584),
    .I0(n583),
    .I1(n582)
  );
  //AND U388bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U388bar (
    .O(n584bar),
    .I0(n583bar),
    .I1(n582bar)
  );
  //OR U389
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U389 (
    .O(n582),
    .I0(n581),
    .I1(n580)
  );
  //AND U389bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U389bar (
    .O(n582bar),
    .I0(n581bar),
    .I1(n580bar)
  );
  //OR U390
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U390 (
    .O(n580),
    .I0(in[158]),
    .I1(in[142])
  );
  //AND U390bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U390bar (
    .O(n580bar),
    .I0(inbar[158]),
    .I1(inbar[142])
  );
  //OR U391
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U391 (
    .O(n581),
    .I0(in[175]),
    .I1(in[164])
  );
  //AND U391bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U391bar (
    .O(n581bar),
    .I0(inbar[175]),
    .I1(inbar[164])
  );
  //OR U392
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U392 (
    .O(n583),
    .I0(n579),
    .I1(n578)
  );
  //AND U392bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U392bar (
    .O(n583bar),
    .I0(n579bar),
    .I1(n578bar)
  );
  //OR U393
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U393 (
    .O(n578),
    .I0(in[228]),
    .I1(in[204])
  );
  //AND U393bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U393bar (
    .O(n578bar),
    .I0(inbar[228]),
    .I1(inbar[204])
  );
  //OR U394
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U394 (
    .O(n579),
    .I0(in[91]),
    .I1(in[87])
  );
  //AND U394bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U394bar (
    .O(n579bar),
    .I0(inbar[91]),
    .I1(inbar[87])
  );
  //OR U395
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U395 (
    .O(n585),
    .I0(n577),
    .I1(n576)
  );
  //AND U395bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U395bar (
    .O(n585bar),
    .I0(n577bar),
    .I1(n576bar)
  );
  //OR U396
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U396 (
    .O(n576),
    .I0(n575),
    .I1(n574)
  );
  //AND U396bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U396bar (
    .O(n576bar),
    .I0(n575bar),
    .I1(n574bar)
  );
  //OR U397
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U397 (
    .O(n574),
    .I0(in_21),
    .I1(in_11)
  );
  //AND U397bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U397bar (
    .O(n574bar),
    .I0(in_21bar),
    .I1(in_11bar)
  );
  //OR U398
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U398 (
    .O(n575),
    .I0(in_5),
    .I1(in_3)
  );
  //AND U398bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U398bar (
    .O(n575bar),
    .I0(in_5bar),
    .I1(in_3bar)
  );
  //OR U399
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U399 (
    .O(n577),
    .I0(n573),
    .I1(n572)
  );
  //AND U399bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U399bar (
    .O(n577bar),
    .I0(n573bar),
    .I1(n572bar)
  );
  //OR U400
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U400 (
    .O(n572),
    .I0(in_68),
    .I1(in_64)
  );
  //AND U400bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U400bar (
    .O(n572bar),
    .I0(in_68bar),
    .I1(in_64bar)
  );
  //OR U401
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U401 (
    .O(n573),
    .I0(in_76),
    .I1(in_73)
  );
  //AND U401bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U401bar (
    .O(n573bar),
    .I0(in_76bar),
    .I1(in_73bar)
  );
  //OR U402
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U402 (
    .O(n601),
    .I0(n778),
    .I1(n571)
  );
  //AND U402bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U402bar (
    .O(n601bar),
    .I0(n778bar),
    .I1(n571bar)
  );
  //OR U403
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U403 (
    .O(n571),
    .I0(in[100]),
    .I1(n965)
  );
  //AND U403bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U403bar (
    .O(n571bar),
    .I0(inbar[100]),
    .I1(n965bar)
  );
  //OR U404
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U404 (
    .O(n965),
    .I0(n570),
    .I1(n569)
  );
  //AND U404bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U404bar (
    .O(n965bar),
    .I0(n570bar),
    .I1(n569bar)
  );
  //OR U405
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U405 (
    .O(n569),
    .I0(n568),
    .I1(n567)
  );
  //AND U405bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U405bar (
    .O(n569bar),
    .I0(n568bar),
    .I1(n567bar)
  );
  //OR U406
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U406 (
    .O(n567),
    .I0(n566),
    .I1(n565)
  );
  //AND U406bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U406bar (
    .O(n567bar),
    .I0(n566bar),
    .I1(n565bar)
  );
  //OR U407
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U407 (
    .O(n565),
    .I0(n817),
    .I1(n750)
  );
  //AND U407bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U407bar (
    .O(n565bar),
    .I0(n817bar),
    .I1(n750bar)
  );
  //OR U408
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U408 (
    .O(n750),
    .I0(n564),
    .I1(n563)
  );
  //AND U408bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U408bar (
    .O(n750bar),
    .I0(n564bar),
    .I1(n563bar)
  );
  //OR U409
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U409 (
    .O(n563),
    .I0(n562),
    .I1(n561)
  );
  //AND U409bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U409bar (
    .O(n563bar),
    .I0(n562bar),
    .I1(n561bar)
  );
  //OR U410
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U410 (
    .O(n561),
    .I0(n560),
    .I1(n559)
  );
  //AND U410bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U410bar (
    .O(n561bar),
    .I0(n560bar),
    .I1(n559bar)
  );
  //OR U411
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U411 (
    .O(n559),
    .I0(in[119]),
    .I1(in[103])
  );
  //AND U411bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U411bar (
    .O(n559bar),
    .I0(inbar[119]),
    .I1(inbar[103])
  );
  //OR U412
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U412 (
    .O(n560),
    .I0(in[137]),
    .I1(in[133])
  );
  //AND U412bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U412bar (
    .O(n560bar),
    .I0(inbar[137]),
    .I1(inbar[133])
  );
  //OR U413
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U413 (
    .O(n562),
    .I0(n558),
    .I1(n557)
  );
  //AND U413bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U413bar (
    .O(n562bar),
    .I0(n558bar),
    .I1(n557bar)
  );
  //OR U414
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U414 (
    .O(n557),
    .I0(in[176]),
    .I1(in[173])
  );
  //AND U414bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U414bar (
    .O(n557bar),
    .I0(inbar[176]),
    .I1(inbar[173])
  );
  //OR U415
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U415 (
    .O(n558),
    .I0(in[210]),
    .I1(in[181])
  );
  //AND U415bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U415bar (
    .O(n558bar),
    .I0(inbar[210]),
    .I1(inbar[181])
  );
  //OR U416
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U416 (
    .O(n564),
    .I0(n556),
    .I1(n555)
  );
  //AND U416bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U416bar (
    .O(n564bar),
    .I0(n556bar),
    .I1(n555bar)
  );
  //OR U417
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U417 (
    .O(n555),
    .I0(n554),
    .I1(n553)
  );
  //AND U417bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U417bar (
    .O(n555bar),
    .I0(n554bar),
    .I1(n553bar)
  );
  //OR U418
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U418 (
    .O(n553),
    .I0(in_13),
    .I1(in[234])
  );
  //AND U418bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U418bar (
    .O(n553bar),
    .I0(in_13bar),
    .I1(inbar[234])
  );
  //OR U419
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U419 (
    .O(n554),
    .I0(in_38),
    .I1(in_32)
  );
  //AND U419bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U419bar (
    .O(n554bar),
    .I0(in_38bar),
    .I1(in_32bar)
  );
  //OR U420
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U420 (
    .O(n556),
    .I0(n552),
    .I1(n551)
  );
  //AND U420bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U420bar (
    .O(n556bar),
    .I0(n552bar),
    .I1(n551bar)
  );
  //OR U421
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U421 (
    .O(n551),
    .I0(in_42),
    .I1(in_41)
  );
  //AND U421bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U421bar (
    .O(n551bar),
    .I0(in_42bar),
    .I1(in_41bar)
  );
  //OR U422
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U422 (
    .O(n552),
    .I0(in_7),
    .I1(in_49)
  );
  //AND U422bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U422bar (
    .O(n552bar),
    .I0(in_7bar),
    .I1(in_49bar)
  );
  //OR U423
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U423 (
    .O(n817),
    .I0(n550),
    .I1(n549)
  );
  //AND U423bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U423bar (
    .O(n817bar),
    .I0(n550bar),
    .I1(n549bar)
  );
  //OR U424
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U424 (
    .O(n549),
    .I0(n548),
    .I1(n547)
  );
  //AND U424bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U424bar (
    .O(n549bar),
    .I0(n548bar),
    .I1(n547bar)
  );
  //OR U425
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U425 (
    .O(n547),
    .I0(n546),
    .I1(n545)
  );
  //AND U425bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U425bar (
    .O(n547bar),
    .I0(n546bar),
    .I1(n545bar)
  );
  //OR U426
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U426 (
    .O(n545),
    .I0(in[159]),
    .I1(in[105])
  );
  //AND U426bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U426bar (
    .O(n545bar),
    .I0(inbar[159]),
    .I1(inbar[105])
  );
  //OR U427
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U427 (
    .O(n546),
    .I0(in[206]),
    .I1(in[183])
  );
  //AND U427bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U427bar (
    .O(n546bar),
    .I0(inbar[206]),
    .I1(inbar[183])
  );
  //OR U428
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U428 (
    .O(n548),
    .I0(n544),
    .I1(n543)
  );
  //AND U428bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U428bar (
    .O(n548bar),
    .I0(n544bar),
    .I1(n543bar)
  );
  //OR U429
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U429 (
    .O(n543),
    .I0(in[229]),
    .I1(in[219])
  );
  //AND U429bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U429bar (
    .O(n543bar),
    .I0(inbar[229]),
    .I1(inbar[219])
  );
  //OR U430
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U430 (
    .O(n544),
    .I0(in[235]),
    .I1(in[232])
  );
  //AND U430bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U430bar (
    .O(n544bar),
    .I0(inbar[235]),
    .I1(inbar[232])
  );
  //OR U431
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U431 (
    .O(n550),
    .I0(n542),
    .I1(n541)
  );
  //AND U431bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U431bar (
    .O(n550bar),
    .I0(n542bar),
    .I1(n541bar)
  );
  //OR U432
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U432 (
    .O(n541),
    .I0(n540),
    .I1(n539)
  );
  //AND U432bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U432bar (
    .O(n541bar),
    .I0(n540bar),
    .I1(n539bar)
  );
  //OR U433
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U433 (
    .O(n539),
    .I0(in[249]),
    .I1(in[242])
  );
  //AND U433bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U433bar (
    .O(n539bar),
    .I0(inbar[249]),
    .I1(inbar[242])
  );
  //OR U434
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U434 (
    .O(n540),
    .I0(in[89]),
    .I1(in[254])
  );
  //AND U434bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U434bar (
    .O(n540bar),
    .I0(inbar[89]),
    .I1(inbar[254])
  );
  //OR U435
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U435 (
    .O(n542),
    .I0(n538),
    .I1(n537)
  );
  //AND U435bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U435bar (
    .O(n542bar),
    .I0(n538bar),
    .I1(n537bar)
  );
  //OR U436
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U436 (
    .O(n537),
    .I0(in_14),
    .I1(in[99])
  );
  //AND U436bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U436bar (
    .O(n537bar),
    .I0(in_14bar),
    .I1(inbar[99])
  );
  //OR U437
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U437 (
    .O(n538),
    .I0(in_60),
    .I1(in_18)
  );
  //AND U437bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U437bar (
    .O(n538bar),
    .I0(in_60bar),
    .I1(in_18bar)
  );
  //OR U438
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U438 (
    .O(n566),
    .I0(in[113]),
    .I1(n763)
  );
  //AND U438bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U438bar (
    .O(n566bar),
    .I0(inbar[113]),
    .I1(n763bar)
  );
  //OR U439
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U439 (
    .O(n763),
    .I0(n536),
    .I1(n535)
  );
  //AND U439bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U439bar (
    .O(n763bar),
    .I0(n536bar),
    .I1(n535bar)
  );
  //OR U440
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U440 (
    .O(n535),
    .I0(n534),
    .I1(n533)
  );
  //AND U440bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U440bar (
    .O(n535bar),
    .I0(n534bar),
    .I1(n533bar)
  );
  //OR U441
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U441 (
    .O(n533),
    .I0(n532),
    .I1(n531)
  );
  //AND U441bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U441bar (
    .O(n533bar),
    .I0(n532bar),
    .I1(n531bar)
  );
  //OR U442
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U442 (
    .O(n531),
    .I0(in[115]),
    .I1(in[110])
  );
  //AND U442bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U442bar (
    .O(n531bar),
    .I0(inbar[115]),
    .I1(inbar[110])
  );
  //OR U443
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U443 (
    .O(n532),
    .I0(in[125]),
    .I1(in[117])
  );
  //AND U443bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U443bar (
    .O(n532bar),
    .I0(inbar[125]),
    .I1(inbar[117])
  );
  //OR U444
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U444 (
    .O(n534),
    .I0(n530),
    .I1(n529)
  );
  //AND U444bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U444bar (
    .O(n534bar),
    .I0(n530bar),
    .I1(n529bar)
  );
  //OR U445
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U445 (
    .O(n529),
    .I0(in[180]),
    .I1(in[128])
  );
  //AND U445bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U445bar (
    .O(n529bar),
    .I0(inbar[180]),
    .I1(inbar[128])
  );
  //OR U446
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U446 (
    .O(n530),
    .I0(in[205]),
    .I1(in[201])
  );
  //AND U446bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U446bar (
    .O(n530bar),
    .I0(inbar[205]),
    .I1(inbar[201])
  );
  //OR U447
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U447 (
    .O(n536),
    .I0(n528),
    .I1(n527)
  );
  //AND U447bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U447bar (
    .O(n536bar),
    .I0(n528bar),
    .I1(n527bar)
  );
  //OR U448
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U448 (
    .O(n527),
    .I0(n526),
    .I1(n525)
  );
  //AND U448bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U448bar (
    .O(n527bar),
    .I0(n526bar),
    .I1(n525bar)
  );
  //OR U449
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U449 (
    .O(n525),
    .I0(in[244]),
    .I1(in[239])
  );
  //AND U449bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U449bar (
    .O(n525bar),
    .I0(inbar[244]),
    .I1(inbar[239])
  );
  //OR U450
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U450 (
    .O(n526),
    .I0(in[95]),
    .I1(in[83])
  );
  //AND U450bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U450bar (
    .O(n526bar),
    .I0(inbar[95]),
    .I1(inbar[83])
  );
  //OR U451
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U451 (
    .O(n528),
    .I0(n524),
    .I1(n523)
  );
  //AND U451bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U451bar (
    .O(n528bar),
    .I0(n524bar),
    .I1(n523bar)
  );
  //OR U452
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U452 (
    .O(n523),
    .I0(in_24),
    .I1(in[97])
  );
  //AND U452bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U452bar (
    .O(n523bar),
    .I0(in_24bar),
    .I1(inbar[97])
  );
  //OR U453
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U453 (
    .O(n524),
    .I0(in_33),
    .I1(in_27)
  );
  //AND U453bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U453bar (
    .O(n524bar),
    .I0(in_33bar),
    .I1(in_27bar)
  );
  //OR U454
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U454 (
    .O(n568),
    .I0(n522),
    .I1(n521)
  );
  //AND U454bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U454bar (
    .O(n568bar),
    .I0(n522bar),
    .I1(n521bar)
  );
  //OR U455
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U455 (
    .O(n521),
    .I0(in[145]),
    .I1(in[126])
  );
  //AND U455bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U455bar (
    .O(n521bar),
    .I0(inbar[145]),
    .I1(inbar[126])
  );
  //OR U456
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U456 (
    .O(n522),
    .I0(in[169]),
    .I1(n520)
  );
  //AND U456bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U456bar (
    .O(n522bar),
    .I0(inbar[169]),
    .I1(n520bar)
  );
  //OR U457
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U457 (
    .O(n520),
    .I0(in[221]),
    .I1(in[172])
  );
  //AND U457bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U457bar (
    .O(n520bar),
    .I0(inbar[221]),
    .I1(inbar[172])
  );
  //OR U458
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U458 (
    .O(n570),
    .I0(n519),
    .I1(n518)
  );
  //AND U458bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U458bar (
    .O(n570bar),
    .I0(n519bar),
    .I1(n518bar)
  );
  //OR U459
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U459 (
    .O(n518),
    .I0(n517),
    .I1(n516)
  );
  //AND U459bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U459bar (
    .O(n518bar),
    .I0(n517bar),
    .I1(n516bar)
  );
  //OR U460
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U460 (
    .O(n516),
    .I0(in[241]),
    .I1(in[224])
  );
  //AND U460bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U460bar (
    .O(n516bar),
    .I0(inbar[241]),
    .I1(inbar[224])
  );
  //OR U461
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U461 (
    .O(n517),
    .I0(in[86]),
    .I1(n515)
  );
  //AND U461bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U461bar (
    .O(n517bar),
    .I0(inbar[86]),
    .I1(n515bar)
  );
  //OR U462
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U462 (
    .O(n515),
    .I0(in_43),
    .I1(in_34)
  );
  //AND U462bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U462bar (
    .O(n515bar),
    .I0(in_43bar),
    .I1(in_34bar)
  );
  //OR U463
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U463 (
    .O(n519),
    .I0(n514),
    .I1(n513)
  );
  //AND U463bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U463bar (
    .O(n519bar),
    .I0(n514bar),
    .I1(n513bar)
  );
  //OR U464
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U464 (
    .O(n513),
    .I0(in_65),
    .I1(in_51)
  );
  //AND U464bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U464bar (
    .O(n513bar),
    .I0(in_65bar),
    .I1(in_51bar)
  );
  //OR U465
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U465 (
    .O(n514),
    .I0(in_75),
    .I1(n512)
  );
  //AND U465bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U465bar (
    .O(n514bar),
    .I0(in_75bar),
    .I1(n512bar)
  );
  //OR U466
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U466 (
    .O(n512),
    .I0(in_81),
    .I1(in_77)
  );
  //AND U466bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U466bar (
    .O(n512bar),
    .I0(in_81bar),
    .I1(in_77bar)
  );
  //OR U467
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U467 (
    .O(n778),
    .I0(n511),
    .I1(n510)
  );
  //AND U467bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U467bar (
    .O(n778bar),
    .I0(n511bar),
    .I1(n510bar)
  );
  //OR U468
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U468 (
    .O(n510),
    .I0(n509),
    .I1(n508)
  );
  //AND U468bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U468bar (
    .O(n510bar),
    .I0(n509bar),
    .I1(n508bar)
  );
  //OR U469
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U469 (
    .O(n508),
    .I0(n507),
    .I1(n506)
  );
  //AND U469bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U469bar (
    .O(n508bar),
    .I0(n507bar),
    .I1(n506bar)
  );
  //OR U470
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U470 (
    .O(n506),
    .I0(in[107]),
    .I1(in[101])
  );
  //AND U470bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U470bar (
    .O(n506bar),
    .I0(inbar[107]),
    .I1(inbar[101])
  );
  //OR U471
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U471 (
    .O(n507),
    .I0(in[139]),
    .I1(in[132])
  );
  //AND U471bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U471bar (
    .O(n507bar),
    .I0(inbar[139]),
    .I1(inbar[132])
  );
  //OR U472
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U472 (
    .O(n509),
    .I0(n505),
    .I1(n504)
  );
  //AND U472bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U472bar (
    .O(n509bar),
    .I0(n505bar),
    .I1(n504bar)
  );
  //OR U473
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U473 (
    .O(n504),
    .I0(in[146]),
    .I1(in[141])
  );
  //AND U473bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U473bar (
    .O(n504bar),
    .I0(inbar[146]),
    .I1(inbar[141])
  );
  //OR U474
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U474 (
    .O(n505),
    .I0(in[203]),
    .I1(in[179])
  );
  //AND U474bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U474bar (
    .O(n505bar),
    .I0(inbar[203]),
    .I1(inbar[179])
  );
  //OR U475
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U475 (
    .O(n511),
    .I0(n503),
    .I1(n502)
  );
  //AND U475bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U475bar (
    .O(n511bar),
    .I0(n503bar),
    .I1(n502bar)
  );
  //OR U476
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U476 (
    .O(n502),
    .I0(n501),
    .I1(n500)
  );
  //AND U476bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U476bar (
    .O(n502bar),
    .I0(n501bar),
    .I1(n500bar)
  );
  //OR U477
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U477 (
    .O(n500),
    .I0(in[243]),
    .I1(in[222])
  );
  //AND U477bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U477bar (
    .O(n500bar),
    .I0(inbar[243]),
    .I1(inbar[222])
  );
  //OR U478
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U478 (
    .O(n501),
    .I0(in[251]),
    .I1(in[250])
  );
  //AND U478bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U478bar (
    .O(n501bar),
    .I0(inbar[251]),
    .I1(inbar[250])
  );
  //OR U479
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U479 (
    .O(n503),
    .I0(n499),
    .I1(n498)
  );
  //AND U479bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U479bar (
    .O(n503bar),
    .I0(n499bar),
    .I1(n498bar)
  );
  //OR U480
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U480 (
    .O(n498),
    .I0(in_37),
    .I1(in_19)
  );
  //AND U480bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U480bar (
    .O(n498bar),
    .I0(in_37bar),
    .I1(in_19bar)
  );
  //OR U481
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U481 (
    .O(n499),
    .I0(in_78),
    .I1(in_6)
  );
  //AND U481bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U481bar (
    .O(n499bar),
    .I0(in_78bar),
    .I1(in_6bar)
  );
  //OR U482
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U482 (
    .O(n603),
    .I0(n497),
    .I1(n496)
  );
  //AND U482bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U482bar (
    .O(n603bar),
    .I0(n497bar),
    .I1(n496bar)
  );
  //OR U483
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U483 (
    .O(n496),
    .I0(in[112]),
    .I1(in[102])
  );
  //AND U483bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U483bar (
    .O(n496bar),
    .I0(inbar[112]),
    .I1(inbar[102])
  );
  //OR U484
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U484 (
    .O(n497),
    .I0(in[123]),
    .I1(n495)
  );
  //AND U484bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U484bar (
    .O(n497bar),
    .I0(inbar[123]),
    .I1(n495bar)
  );
  //OR U485
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U485 (
    .O(n495),
    .I0(in[143]),
    .I1(in[130])
  );
  //AND U485bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U485bar (
    .O(n495bar),
    .I0(inbar[143]),
    .I1(inbar[130])
  );
  //OR U486
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U486 (
    .O(n605),
    .I0(n494),
    .I1(n493)
  );
  //AND U486bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U486bar (
    .O(n605bar),
    .I0(n494bar),
    .I1(n493bar)
  );
  //OR U487
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U487 (
    .O(n493),
    .I0(n492),
    .I1(n491)
  );
  //AND U487bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U487bar (
    .O(n493bar),
    .I0(n492bar),
    .I1(n491bar)
  );
  //OR U488
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U488 (
    .O(n491),
    .I0(in[216]),
    .I1(in[213])
  );
  //AND U488bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U488bar (
    .O(n491bar),
    .I0(inbar[216]),
    .I1(inbar[213])
  );
  //OR U489
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U489 (
    .O(n492),
    .I0(in[227]),
    .I1(n490)
  );
  //AND U489bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U489bar (
    .O(n492bar),
    .I0(inbar[227]),
    .I1(n490bar)
  );
  //OR U490
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U490 (
    .O(n490),
    .I0(in_0),
    .I1(in[248])
  );
  //AND U490bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U490bar (
    .O(n490bar),
    .I0(in_0bar),
    .I1(inbar[248])
  );
  //OR U491
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U491 (
    .O(n494),
    .I0(n489),
    .I1(n488)
  );
  //AND U491bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U491bar (
    .O(n494bar),
    .I0(n489bar),
    .I1(n488bar)
  );
  //OR U492
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U492 (
    .O(n488),
    .I0(in_46),
    .I1(in_44)
  );
  //AND U492bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U492bar (
    .O(n488bar),
    .I0(in_46bar),
    .I1(in_44bar)
  );
  //OR U493
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U493 (
    .O(n489),
    .I0(in_50),
    .I1(n487)
  );
  //AND U493bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U493bar (
    .O(n489bar),
    .I0(in_50bar),
    .I1(n487bar)
  );
  //OR U494
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U494 (
    .O(n487),
    .I0(in_9),
    .I1(in_80)
  );
  //AND U494bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U494bar (
    .O(n487bar),
    .I0(in_9bar),
    .I1(in_80bar)
  );
endmodule

module sBox_2 ( in, out );

  input wire [7:0] in;
//input_done

  output wire [7:0] out;
//output_done

  wire [255:0] decodeOut;
//wire_done

  decode_2 dec ( .in(in), .out(decodeOut) );
  encode_2 enc ( .in(decodeOut), .out(out) );
endmodule

module CD2_9 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD2_10 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD2_11 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD2_12 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD4_5 ( a, b, y );

  input wire [3:0] a;
  input wire [3:0] b;
  wire [3:0] abar;
  wire [3:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
//input_done

  output wire [15:0] y;
  wire [15:0] ybar;
//output_done

//wire_done

  //AND U1
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1 (
    .O(y[9]),
    .I0(b[1]),
    .I1(a[2])
  );
  //OR U1bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1bar (
    .O(ybar[9]),
    .I0(bbar[1]),
    .I1(abar[2])
  );
  //AND U2
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2 (
    .O(y[8]),
    .I0(b[0]),
    .I1(a[2])
  );
  //OR U2bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2bar (
    .O(ybar[8]),
    .I0(bbar[0]),
    .I1(abar[2])
  );
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[7]),
    .I0(b[3]),
    .I1(a[1])
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[7]),
    .I0(bbar[3]),
    .I1(abar[1])
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[6]),
    .I0(b[2]),
    .I1(a[1])
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[6]),
    .I0(bbar[2]),
    .I1(abar[1])
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[5]),
    .I0(a[1]),
    .I1(b[1])
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[5]),
    .I0(abar[1]),
    .I1(bbar[1])
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[4]),
    .I0(a[1]),
    .I1(b[0])
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[4]),
    .I0(abar[1]),
    .I1(bbar[0])
  );
  //AND U7
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7 (
    .O(y[3]),
    .I0(a[0]),
    .I1(b[3])
  );
  //OR U7bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7bar (
    .O(ybar[3]),
    .I0(abar[0]),
    .I1(bbar[3])
  );
  //AND U8
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8 (
    .O(y[2]),
    .I0(a[0]),
    .I1(b[2])
  );
  //OR U8bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8bar (
    .O(ybar[2]),
    .I0(abar[0]),
    .I1(bbar[2])
  );
  //AND U9
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9 (
    .O(y[1]),
    .I0(a[0]),
    .I1(b[1])
  );
  //OR U9bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9bar (
    .O(ybar[1]),
    .I0(abar[0]),
    .I1(bbar[1])
  );
  //AND U10
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10 (
    .O(y[15]),
    .I0(a[3]),
    .I1(b[3])
  );
  //OR U10bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10bar (
    .O(ybar[15]),
    .I0(abar[3]),
    .I1(bbar[3])
  );
  //AND U11
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11 (
    .O(y[14]),
    .I0(a[3]),
    .I1(b[2])
  );
  //OR U11bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11bar (
    .O(ybar[14]),
    .I0(abar[3]),
    .I1(bbar[2])
  );
  //AND U12
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12 (
    .O(y[13]),
    .I0(a[3]),
    .I1(b[1])
  );
  //OR U12bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12bar (
    .O(ybar[13]),
    .I0(abar[3]),
    .I1(bbar[1])
  );
  //AND U13
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13 (
    .O(y[12]),
    .I0(a[3]),
    .I1(b[0])
  );
  //OR U13bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13bar (
    .O(ybar[12]),
    .I0(abar[3]),
    .I1(bbar[0])
  );
  //AND U14
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14 (
    .O(y[11]),
    .I0(b[3]),
    .I1(a[2])
  );
  //OR U14bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14bar (
    .O(ybar[11]),
    .I0(bbar[3]),
    .I1(abar[2])
  );
  //AND U15
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15 (
    .O(y[10]),
    .I0(b[2]),
    .I1(a[2])
  );
  //OR U15bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15bar (
    .O(ybar[10]),
    .I0(bbar[2]),
    .I1(abar[2])
  );
  //AND U16
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16 (
    .O(y[0]),
    .I0(a[0]),
    .I1(b[0])
  );
  //OR U16bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16bar (
    .O(ybar[0]),
    .I0(abar[0]),
    .I1(bbar[0])
  );
endmodule

module CD4_6 ( a, b, y );

  input wire [3:0] a;
  input wire [3:0] b;
  wire [3:0] abar;
  wire [3:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
//input_done

  output wire [15:0] y;
  wire [15:0] ybar;
//output_done

//wire_done

  //AND U1
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1 (
    .O(y[9]),
    .I0(b[1]),
    .I1(a[2])
  );
  //OR U1bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1bar (
    .O(ybar[9]),
    .I0(bbar[1]),
    .I1(abar[2])
  );
  //AND U2
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2 (
    .O(y[8]),
    .I0(b[0]),
    .I1(a[2])
  );
  //OR U2bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2bar (
    .O(ybar[8]),
    .I0(bbar[0]),
    .I1(abar[2])
  );
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[7]),
    .I0(b[3]),
    .I1(a[1])
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[7]),
    .I0(bbar[3]),
    .I1(abar[1])
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[6]),
    .I0(b[2]),
    .I1(a[1])
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[6]),
    .I0(bbar[2]),
    .I1(abar[1])
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[5]),
    .I0(a[1]),
    .I1(b[1])
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[5]),
    .I0(abar[1]),
    .I1(bbar[1])
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[4]),
    .I0(a[1]),
    .I1(b[0])
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[4]),
    .I0(abar[1]),
    .I1(bbar[0])
  );
  //AND U7
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7 (
    .O(y[3]),
    .I0(a[0]),
    .I1(b[3])
  );
  //OR U7bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7bar (
    .O(ybar[3]),
    .I0(abar[0]),
    .I1(bbar[3])
  );
  //AND U8
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8 (
    .O(y[2]),
    .I0(a[0]),
    .I1(b[2])
  );
  //OR U8bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8bar (
    .O(ybar[2]),
    .I0(abar[0]),
    .I1(bbar[2])
  );
  //AND U9
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9 (
    .O(y[1]),
    .I0(a[0]),
    .I1(b[1])
  );
  //OR U9bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9bar (
    .O(ybar[1]),
    .I0(abar[0]),
    .I1(bbar[1])
  );
  //AND U10
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10 (
    .O(y[15]),
    .I0(a[3]),
    .I1(b[3])
  );
  //OR U10bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10bar (
    .O(ybar[15]),
    .I0(abar[3]),
    .I1(bbar[3])
  );
  //AND U11
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11 (
    .O(y[14]),
    .I0(a[3]),
    .I1(b[2])
  );
  //OR U11bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11bar (
    .O(ybar[14]),
    .I0(abar[3]),
    .I1(bbar[2])
  );
  //AND U12
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12 (
    .O(y[13]),
    .I0(a[3]),
    .I1(b[1])
  );
  //OR U12bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12bar (
    .O(ybar[13]),
    .I0(abar[3]),
    .I1(bbar[1])
  );
  //AND U13
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13 (
    .O(y[12]),
    .I0(a[3]),
    .I1(b[0])
  );
  //OR U13bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13bar (
    .O(ybar[12]),
    .I0(abar[3]),
    .I1(bbar[0])
  );
  //AND U14
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14 (
    .O(y[11]),
    .I0(b[3]),
    .I1(a[2])
  );
  //OR U14bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14bar (
    .O(ybar[11]),
    .I0(bbar[3]),
    .I1(abar[2])
  );
  //AND U15
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15 (
    .O(y[10]),
    .I0(b[2]),
    .I1(a[2])
  );
  //OR U15bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15bar (
    .O(ybar[10]),
    .I0(bbar[2]),
    .I1(abar[2])
  );
  //AND U16
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16 (
    .O(y[0]),
    .I0(a[0]),
    .I1(b[0])
  );
  //OR U16bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16bar (
    .O(ybar[0]),
    .I0(abar[0]),
    .I1(bbar[0])
  );
endmodule

module CD16_3 ( a, b, y );

  input wire [15:0] a;
  input wire [15:0] b;
  wire [15:0] abar;
  wire [15:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign abar[8] = ~a[8];
  assign abar[9] = ~a[9];
  assign abar[10] = ~a[10];
  assign abar[11] = ~a[11];
  assign abar[12] = ~a[12];
  assign abar[13] = ~a[13];
  assign abar[14] = ~a[14];
  assign abar[15] = ~a[15];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign bbar[8] = ~b[8];
  assign bbar[9] = ~b[9];
  assign bbar[10] = ~b[10];
  assign bbar[11] = ~b[11];
  assign bbar[12] = ~b[12];
  assign bbar[13] = ~b[13];
  assign bbar[14] = ~b[14];
  assign bbar[15] = ~b[15];
//input_done

  output wire [255:0] y;
  wire [255:0] ybar;
//output_done

//wire_done

  //AND U1
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1 (
    .O(y[9]),
    .I0(b[9]),
    .I1(a[0])
  );
  //OR U1bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1bar (
    .O(ybar[9]),
    .I0(bbar[9]),
    .I1(abar[0])
  );
  //AND U2
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2 (
    .O(y[99]),
    .I0(b[3]),
    .I1(a[6])
  );
  //OR U2bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2bar (
    .O(ybar[99]),
    .I0(bbar[3]),
    .I1(abar[6])
  );
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[98]),
    .I0(b[2]),
    .I1(a[6])
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[98]),
    .I0(bbar[2]),
    .I1(abar[6])
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[97]),
    .I0(b[1]),
    .I1(a[6])
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[97]),
    .I0(bbar[1]),
    .I1(abar[6])
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[96]),
    .I0(b[0]),
    .I1(a[6])
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[96]),
    .I0(bbar[0]),
    .I1(abar[6])
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[95]),
    .I0(b[15]),
    .I1(a[5])
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[95]),
    .I0(bbar[15]),
    .I1(abar[5])
  );
  //AND U7
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7 (
    .O(y[94]),
    .I0(b[14]),
    .I1(a[5])
  );
  //OR U7bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7bar (
    .O(ybar[94]),
    .I0(bbar[14]),
    .I1(abar[5])
  );
  //AND U8
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8 (
    .O(y[93]),
    .I0(b[13]),
    .I1(a[5])
  );
  //OR U8bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8bar (
    .O(ybar[93]),
    .I0(bbar[13]),
    .I1(abar[5])
  );
  //AND U9
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9 (
    .O(y[92]),
    .I0(b[12]),
    .I1(a[5])
  );
  //OR U9bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9bar (
    .O(ybar[92]),
    .I0(bbar[12]),
    .I1(abar[5])
  );
  //AND U10
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10 (
    .O(y[91]),
    .I0(b[11]),
    .I1(a[5])
  );
  //OR U10bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10bar (
    .O(ybar[91]),
    .I0(bbar[11]),
    .I1(abar[5])
  );
  //AND U11
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11 (
    .O(y[90]),
    .I0(b[10]),
    .I1(a[5])
  );
  //OR U11bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11bar (
    .O(ybar[90]),
    .I0(bbar[10]),
    .I1(abar[5])
  );
  //AND U12
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12 (
    .O(y[8]),
    .I0(b[8]),
    .I1(a[0])
  );
  //OR U12bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12bar (
    .O(ybar[8]),
    .I0(bbar[8]),
    .I1(abar[0])
  );
  //AND U13
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13 (
    .O(y[89]),
    .I0(a[5]),
    .I1(b[9])
  );
  //OR U13bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13bar (
    .O(ybar[89]),
    .I0(abar[5]),
    .I1(bbar[9])
  );
  //AND U14
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14 (
    .O(y[88]),
    .I0(b[8]),
    .I1(a[5])
  );
  //OR U14bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14bar (
    .O(ybar[88]),
    .I0(bbar[8]),
    .I1(abar[5])
  );
  //AND U15
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15 (
    .O(y[87]),
    .I0(b[7]),
    .I1(a[5])
  );
  //OR U15bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15bar (
    .O(ybar[87]),
    .I0(bbar[7]),
    .I1(abar[5])
  );
  //AND U16
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16 (
    .O(y[86]),
    .I0(b[6]),
    .I1(a[5])
  );
  //OR U16bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16bar (
    .O(ybar[86]),
    .I0(bbar[6]),
    .I1(abar[5])
  );
  //AND U17
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U17 (
    .O(y[85]),
    .I0(b[5]),
    .I1(a[5])
  );
  //OR U17bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U17bar (
    .O(ybar[85]),
    .I0(bbar[5]),
    .I1(abar[5])
  );
  //AND U18
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U18 (
    .O(y[84]),
    .I0(b[4]),
    .I1(a[5])
  );
  //OR U18bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U18bar (
    .O(ybar[84]),
    .I0(bbar[4]),
    .I1(abar[5])
  );
  //AND U19
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U19 (
    .O(y[83]),
    .I0(a[5]),
    .I1(b[3])
  );
  //OR U19bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U19bar (
    .O(ybar[83]),
    .I0(abar[5]),
    .I1(bbar[3])
  );
  //AND U20
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U20 (
    .O(y[82]),
    .I0(a[5]),
    .I1(b[2])
  );
  //OR U20bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U20bar (
    .O(ybar[82]),
    .I0(abar[5]),
    .I1(bbar[2])
  );
  //AND U21
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U21 (
    .O(y[81]),
    .I0(a[5]),
    .I1(b[1])
  );
  //OR U21bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U21bar (
    .O(ybar[81]),
    .I0(abar[5]),
    .I1(bbar[1])
  );
  //AND U22
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U22 (
    .O(y[80]),
    .I0(a[5]),
    .I1(b[0])
  );
  //OR U22bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U22bar (
    .O(ybar[80]),
    .I0(abar[5]),
    .I1(bbar[0])
  );
  //AND U23
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U23 (
    .O(y[7]),
    .I0(b[7]),
    .I1(a[0])
  );
  //OR U23bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U23bar (
    .O(ybar[7]),
    .I0(bbar[7]),
    .I1(abar[0])
  );
  //AND U24
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U24 (
    .O(y[79]),
    .I0(a[4]),
    .I1(b[15])
  );
  //OR U24bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U24bar (
    .O(ybar[79]),
    .I0(abar[4]),
    .I1(bbar[15])
  );
  //AND U25
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U25 (
    .O(y[78]),
    .I0(a[4]),
    .I1(b[14])
  );
  //OR U25bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U25bar (
    .O(ybar[78]),
    .I0(abar[4]),
    .I1(bbar[14])
  );
  //AND U26
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U26 (
    .O(y[77]),
    .I0(a[4]),
    .I1(b[13])
  );
  //OR U26bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U26bar (
    .O(ybar[77]),
    .I0(abar[4]),
    .I1(bbar[13])
  );
  //AND U27
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U27 (
    .O(y[76]),
    .I0(a[4]),
    .I1(b[12])
  );
  //OR U27bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U27bar (
    .O(ybar[76]),
    .I0(abar[4]),
    .I1(bbar[12])
  );
  //AND U28
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U28 (
    .O(y[75]),
    .I0(a[4]),
    .I1(b[11])
  );
  //OR U28bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U28bar (
    .O(ybar[75]),
    .I0(abar[4]),
    .I1(bbar[11])
  );
  //AND U29
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U29 (
    .O(y[74]),
    .I0(a[4]),
    .I1(b[10])
  );
  //OR U29bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U29bar (
    .O(ybar[74]),
    .I0(abar[4]),
    .I1(bbar[10])
  );
  //AND U30
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U30 (
    .O(y[73]),
    .I0(a[4]),
    .I1(b[9])
  );
  //OR U30bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U30bar (
    .O(ybar[73]),
    .I0(abar[4]),
    .I1(bbar[9])
  );
  //AND U31
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U31 (
    .O(y[72]),
    .I0(a[4]),
    .I1(b[8])
  );
  //OR U31bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U31bar (
    .O(ybar[72]),
    .I0(abar[4]),
    .I1(bbar[8])
  );
  //AND U32
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U32 (
    .O(y[71]),
    .I0(a[4]),
    .I1(b[7])
  );
  //OR U32bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U32bar (
    .O(ybar[71]),
    .I0(abar[4]),
    .I1(bbar[7])
  );
  //AND U33
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U33 (
    .O(y[70]),
    .I0(a[4]),
    .I1(b[6])
  );
  //OR U33bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U33bar (
    .O(ybar[70]),
    .I0(abar[4]),
    .I1(bbar[6])
  );
  //AND U34
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U34 (
    .O(y[6]),
    .I0(b[6]),
    .I1(a[0])
  );
  //OR U34bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U34bar (
    .O(ybar[6]),
    .I0(bbar[6]),
    .I1(abar[0])
  );
  //AND U35
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U35 (
    .O(y[69]),
    .I0(a[4]),
    .I1(b[5])
  );
  //OR U35bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U35bar (
    .O(ybar[69]),
    .I0(abar[4]),
    .I1(bbar[5])
  );
  //AND U36
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U36 (
    .O(y[68]),
    .I0(a[4]),
    .I1(b[4])
  );
  //OR U36bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U36bar (
    .O(ybar[68]),
    .I0(abar[4]),
    .I1(bbar[4])
  );
  //AND U37
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U37 (
    .O(y[67]),
    .I0(a[4]),
    .I1(b[3])
  );
  //OR U37bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U37bar (
    .O(ybar[67]),
    .I0(abar[4]),
    .I1(bbar[3])
  );
  //AND U38
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U38 (
    .O(y[66]),
    .I0(a[4]),
    .I1(b[2])
  );
  //OR U38bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U38bar (
    .O(ybar[66]),
    .I0(abar[4]),
    .I1(bbar[2])
  );
  //AND U39
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U39 (
    .O(y[65]),
    .I0(a[4]),
    .I1(b[1])
  );
  //OR U39bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U39bar (
    .O(ybar[65]),
    .I0(abar[4]),
    .I1(bbar[1])
  );
  //AND U40
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U40 (
    .O(y[64]),
    .I0(a[4]),
    .I1(b[0])
  );
  //OR U40bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U40bar (
    .O(ybar[64]),
    .I0(abar[4]),
    .I1(bbar[0])
  );
  //AND U41
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U41 (
    .O(y[63]),
    .I0(a[3]),
    .I1(b[15])
  );
  //OR U41bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U41bar (
    .O(ybar[63]),
    .I0(abar[3]),
    .I1(bbar[15])
  );
  //AND U42
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U42 (
    .O(y[62]),
    .I0(a[3]),
    .I1(b[14])
  );
  //OR U42bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U42bar (
    .O(ybar[62]),
    .I0(abar[3]),
    .I1(bbar[14])
  );
  //AND U43
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U43 (
    .O(y[61]),
    .I0(a[3]),
    .I1(b[13])
  );
  //OR U43bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U43bar (
    .O(ybar[61]),
    .I0(abar[3]),
    .I1(bbar[13])
  );
  //AND U44
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U44 (
    .O(y[60]),
    .I0(a[3]),
    .I1(b[12])
  );
  //OR U44bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U44bar (
    .O(ybar[60]),
    .I0(abar[3]),
    .I1(bbar[12])
  );
  //AND U45
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U45 (
    .O(y[5]),
    .I0(b[5]),
    .I1(a[0])
  );
  //OR U45bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U45bar (
    .O(ybar[5]),
    .I0(bbar[5]),
    .I1(abar[0])
  );
  //AND U46
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U46 (
    .O(y[59]),
    .I0(a[3]),
    .I1(b[11])
  );
  //OR U46bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U46bar (
    .O(ybar[59]),
    .I0(abar[3]),
    .I1(bbar[11])
  );
  //AND U47
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U47 (
    .O(y[58]),
    .I0(a[3]),
    .I1(b[10])
  );
  //OR U47bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U47bar (
    .O(ybar[58]),
    .I0(abar[3]),
    .I1(bbar[10])
  );
  //AND U48
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U48 (
    .O(y[57]),
    .I0(a[3]),
    .I1(b[9])
  );
  //OR U48bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U48bar (
    .O(ybar[57]),
    .I0(abar[3]),
    .I1(bbar[9])
  );
  //AND U49
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U49 (
    .O(y[56]),
    .I0(a[3]),
    .I1(b[8])
  );
  //OR U49bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U49bar (
    .O(ybar[56]),
    .I0(abar[3]),
    .I1(bbar[8])
  );
  //AND U50
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U50 (
    .O(y[55]),
    .I0(a[3]),
    .I1(b[7])
  );
  //OR U50bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U50bar (
    .O(ybar[55]),
    .I0(abar[3]),
    .I1(bbar[7])
  );
  //AND U51
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U51 (
    .O(y[54]),
    .I0(a[3]),
    .I1(b[6])
  );
  //OR U51bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U51bar (
    .O(ybar[54]),
    .I0(abar[3]),
    .I1(bbar[6])
  );
  //AND U52
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U52 (
    .O(y[53]),
    .I0(a[3]),
    .I1(b[5])
  );
  //OR U52bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U52bar (
    .O(ybar[53]),
    .I0(abar[3]),
    .I1(bbar[5])
  );
  //AND U53
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U53 (
    .O(y[52]),
    .I0(a[3]),
    .I1(b[4])
  );
  //OR U53bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U53bar (
    .O(ybar[52]),
    .I0(abar[3]),
    .I1(bbar[4])
  );
  //AND U54
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U54 (
    .O(y[51]),
    .I0(a[3]),
    .I1(b[3])
  );
  //OR U54bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U54bar (
    .O(ybar[51]),
    .I0(abar[3]),
    .I1(bbar[3])
  );
  //AND U55
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U55 (
    .O(y[50]),
    .I0(a[3]),
    .I1(b[2])
  );
  //OR U55bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U55bar (
    .O(ybar[50]),
    .I0(abar[3]),
    .I1(bbar[2])
  );
  //AND U56
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U56 (
    .O(y[4]),
    .I0(b[4]),
    .I1(a[0])
  );
  //OR U56bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U56bar (
    .O(ybar[4]),
    .I0(bbar[4]),
    .I1(abar[0])
  );
  //AND U57
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U57 (
    .O(y[49]),
    .I0(a[3]),
    .I1(b[1])
  );
  //OR U57bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U57bar (
    .O(ybar[49]),
    .I0(abar[3]),
    .I1(bbar[1])
  );
  //AND U58
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U58 (
    .O(y[48]),
    .I0(a[3]),
    .I1(b[0])
  );
  //OR U58bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U58bar (
    .O(ybar[48]),
    .I0(abar[3]),
    .I1(bbar[0])
  );
  //AND U59
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U59 (
    .O(y[47]),
    .I0(a[2]),
    .I1(b[15])
  );
  //OR U59bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U59bar (
    .O(ybar[47]),
    .I0(abar[2]),
    .I1(bbar[15])
  );
  //AND U60
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U60 (
    .O(y[46]),
    .I0(a[2]),
    .I1(b[14])
  );
  //OR U60bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U60bar (
    .O(ybar[46]),
    .I0(abar[2]),
    .I1(bbar[14])
  );
  //AND U61
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U61 (
    .O(y[45]),
    .I0(a[2]),
    .I1(b[13])
  );
  //OR U61bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U61bar (
    .O(ybar[45]),
    .I0(abar[2]),
    .I1(bbar[13])
  );
  //AND U62
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U62 (
    .O(y[44]),
    .I0(a[2]),
    .I1(b[12])
  );
  //OR U62bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U62bar (
    .O(ybar[44]),
    .I0(abar[2]),
    .I1(bbar[12])
  );
  //AND U63
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U63 (
    .O(y[43]),
    .I0(a[2]),
    .I1(b[11])
  );
  //OR U63bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U63bar (
    .O(ybar[43]),
    .I0(abar[2]),
    .I1(bbar[11])
  );
  //AND U64
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U64 (
    .O(y[42]),
    .I0(a[2]),
    .I1(b[10])
  );
  //OR U64bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U64bar (
    .O(ybar[42]),
    .I0(abar[2]),
    .I1(bbar[10])
  );
  //AND U65
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U65 (
    .O(y[41]),
    .I0(a[2]),
    .I1(b[9])
  );
  //OR U65bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U65bar (
    .O(ybar[41]),
    .I0(abar[2]),
    .I1(bbar[9])
  );
  //AND U66
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U66 (
    .O(y[40]),
    .I0(a[2]),
    .I1(b[8])
  );
  //OR U66bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U66bar (
    .O(ybar[40]),
    .I0(abar[2]),
    .I1(bbar[8])
  );
  //AND U67
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U67 (
    .O(y[3]),
    .I0(b[3]),
    .I1(a[0])
  );
  //OR U67bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U67bar (
    .O(ybar[3]),
    .I0(bbar[3]),
    .I1(abar[0])
  );
  //AND U68
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U68 (
    .O(y[39]),
    .I0(a[2]),
    .I1(b[7])
  );
  //OR U68bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U68bar (
    .O(ybar[39]),
    .I0(abar[2]),
    .I1(bbar[7])
  );
  //AND U69
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U69 (
    .O(y[38]),
    .I0(a[2]),
    .I1(b[6])
  );
  //OR U69bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U69bar (
    .O(ybar[38]),
    .I0(abar[2]),
    .I1(bbar[6])
  );
  //AND U70
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U70 (
    .O(y[37]),
    .I0(a[2]),
    .I1(b[5])
  );
  //OR U70bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U70bar (
    .O(ybar[37]),
    .I0(abar[2]),
    .I1(bbar[5])
  );
  //AND U71
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U71 (
    .O(y[36]),
    .I0(a[2]),
    .I1(b[4])
  );
  //OR U71bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U71bar (
    .O(ybar[36]),
    .I0(abar[2]),
    .I1(bbar[4])
  );
  //AND U72
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U72 (
    .O(y[35]),
    .I0(a[2]),
    .I1(b[3])
  );
  //OR U72bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U72bar (
    .O(ybar[35]),
    .I0(abar[2]),
    .I1(bbar[3])
  );
  //AND U73
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U73 (
    .O(y[34]),
    .I0(a[2]),
    .I1(b[2])
  );
  //OR U73bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U73bar (
    .O(ybar[34]),
    .I0(abar[2]),
    .I1(bbar[2])
  );
  //AND U74
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U74 (
    .O(y[33]),
    .I0(a[2]),
    .I1(b[1])
  );
  //OR U74bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U74bar (
    .O(ybar[33]),
    .I0(abar[2]),
    .I1(bbar[1])
  );
  //AND U75
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U75 (
    .O(y[32]),
    .I0(a[2]),
    .I1(b[0])
  );
  //OR U75bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U75bar (
    .O(ybar[32]),
    .I0(abar[2]),
    .I1(bbar[0])
  );
  //AND U76
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U76 (
    .O(y[31]),
    .I0(a[1]),
    .I1(b[15])
  );
  //OR U76bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U76bar (
    .O(ybar[31]),
    .I0(abar[1]),
    .I1(bbar[15])
  );
  //AND U77
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U77 (
    .O(y[30]),
    .I0(a[1]),
    .I1(b[14])
  );
  //OR U77bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U77bar (
    .O(ybar[30]),
    .I0(abar[1]),
    .I1(bbar[14])
  );
  //AND U78
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U78 (
    .O(y[2]),
    .I0(b[2]),
    .I1(a[0])
  );
  //OR U78bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U78bar (
    .O(ybar[2]),
    .I0(bbar[2]),
    .I1(abar[0])
  );
  //AND U79
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U79 (
    .O(y[29]),
    .I0(a[1]),
    .I1(b[13])
  );
  //OR U79bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U79bar (
    .O(ybar[29]),
    .I0(abar[1]),
    .I1(bbar[13])
  );
  //AND U80
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U80 (
    .O(y[28]),
    .I0(a[1]),
    .I1(b[12])
  );
  //OR U80bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U80bar (
    .O(ybar[28]),
    .I0(abar[1]),
    .I1(bbar[12])
  );
  //AND U81
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U81 (
    .O(y[27]),
    .I0(a[1]),
    .I1(b[11])
  );
  //OR U81bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U81bar (
    .O(ybar[27]),
    .I0(abar[1]),
    .I1(bbar[11])
  );
  //AND U82
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U82 (
    .O(y[26]),
    .I0(a[1]),
    .I1(b[10])
  );
  //OR U82bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U82bar (
    .O(ybar[26]),
    .I0(abar[1]),
    .I1(bbar[10])
  );
  //AND U83
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U83 (
    .O(y[25]),
    .I0(a[1]),
    .I1(b[9])
  );
  //OR U83bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U83bar (
    .O(ybar[25]),
    .I0(abar[1]),
    .I1(bbar[9])
  );
  //AND U84
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U84 (
    .O(y[255]),
    .I0(a[15]),
    .I1(b[15])
  );
  //OR U84bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U84bar (
    .O(ybar[255]),
    .I0(abar[15]),
    .I1(bbar[15])
  );
  //AND U85
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U85 (
    .O(y[254]),
    .I0(a[15]),
    .I1(b[14])
  );
  //OR U85bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U85bar (
    .O(ybar[254]),
    .I0(abar[15]),
    .I1(bbar[14])
  );
  //AND U86
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U86 (
    .O(y[253]),
    .I0(a[15]),
    .I1(b[13])
  );
  //OR U86bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U86bar (
    .O(ybar[253]),
    .I0(abar[15]),
    .I1(bbar[13])
  );
  //AND U87
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U87 (
    .O(y[252]),
    .I0(a[15]),
    .I1(b[12])
  );
  //OR U87bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U87bar (
    .O(ybar[252]),
    .I0(abar[15]),
    .I1(bbar[12])
  );
  //AND U88
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U88 (
    .O(y[251]),
    .I0(a[15]),
    .I1(b[11])
  );
  //OR U88bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U88bar (
    .O(ybar[251]),
    .I0(abar[15]),
    .I1(bbar[11])
  );
  //AND U89
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U89 (
    .O(y[250]),
    .I0(a[15]),
    .I1(b[10])
  );
  //OR U89bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U89bar (
    .O(ybar[250]),
    .I0(abar[15]),
    .I1(bbar[10])
  );
  //AND U90
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U90 (
    .O(y[24]),
    .I0(a[1]),
    .I1(b[8])
  );
  //OR U90bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U90bar (
    .O(ybar[24]),
    .I0(abar[1]),
    .I1(bbar[8])
  );
  //AND U91
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U91 (
    .O(y[249]),
    .I0(a[15]),
    .I1(b[9])
  );
  //OR U91bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U91bar (
    .O(ybar[249]),
    .I0(abar[15]),
    .I1(bbar[9])
  );
  //AND U92
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U92 (
    .O(y[248]),
    .I0(a[15]),
    .I1(b[8])
  );
  //OR U92bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U92bar (
    .O(ybar[248]),
    .I0(abar[15]),
    .I1(bbar[8])
  );
  //AND U93
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U93 (
    .O(y[247]),
    .I0(a[15]),
    .I1(b[7])
  );
  //OR U93bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U93bar (
    .O(ybar[247]),
    .I0(abar[15]),
    .I1(bbar[7])
  );
  //AND U94
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U94 (
    .O(y[246]),
    .I0(a[15]),
    .I1(b[6])
  );
  //OR U94bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U94bar (
    .O(ybar[246]),
    .I0(abar[15]),
    .I1(bbar[6])
  );
  //AND U95
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U95 (
    .O(y[245]),
    .I0(a[15]),
    .I1(b[5])
  );
  //OR U95bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U95bar (
    .O(ybar[245]),
    .I0(abar[15]),
    .I1(bbar[5])
  );
  //AND U96
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U96 (
    .O(y[244]),
    .I0(a[15]),
    .I1(b[4])
  );
  //OR U96bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U96bar (
    .O(ybar[244]),
    .I0(abar[15]),
    .I1(bbar[4])
  );
  //AND U97
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U97 (
    .O(y[243]),
    .I0(a[15]),
    .I1(b[3])
  );
  //OR U97bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U97bar (
    .O(ybar[243]),
    .I0(abar[15]),
    .I1(bbar[3])
  );
  //AND U98
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U98 (
    .O(y[242]),
    .I0(a[15]),
    .I1(b[2])
  );
  //OR U98bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U98bar (
    .O(ybar[242]),
    .I0(abar[15]),
    .I1(bbar[2])
  );
  //AND U99
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U99 (
    .O(y[241]),
    .I0(a[15]),
    .I1(b[1])
  );
  //OR U99bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U99bar (
    .O(ybar[241]),
    .I0(abar[15]),
    .I1(bbar[1])
  );
  //AND U100
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U100 (
    .O(y[240]),
    .I0(a[15]),
    .I1(b[0])
  );
  //OR U100bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U100bar (
    .O(ybar[240]),
    .I0(abar[15]),
    .I1(bbar[0])
  );
  //AND U101
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U101 (
    .O(y[23]),
    .I0(a[1]),
    .I1(b[7])
  );
  //OR U101bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U101bar (
    .O(ybar[23]),
    .I0(abar[1]),
    .I1(bbar[7])
  );
  //AND U102
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U102 (
    .O(y[239]),
    .I0(a[14]),
    .I1(b[15])
  );
  //OR U102bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U102bar (
    .O(ybar[239]),
    .I0(abar[14]),
    .I1(bbar[15])
  );
  //AND U103
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U103 (
    .O(y[238]),
    .I0(a[14]),
    .I1(b[14])
  );
  //OR U103bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U103bar (
    .O(ybar[238]),
    .I0(abar[14]),
    .I1(bbar[14])
  );
  //AND U104
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U104 (
    .O(y[237]),
    .I0(a[14]),
    .I1(b[13])
  );
  //OR U104bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U104bar (
    .O(ybar[237]),
    .I0(abar[14]),
    .I1(bbar[13])
  );
  //AND U105
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U105 (
    .O(y[236]),
    .I0(a[14]),
    .I1(b[12])
  );
  //OR U105bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U105bar (
    .O(ybar[236]),
    .I0(abar[14]),
    .I1(bbar[12])
  );
  //AND U106
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U106 (
    .O(y[235]),
    .I0(a[14]),
    .I1(b[11])
  );
  //OR U106bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U106bar (
    .O(ybar[235]),
    .I0(abar[14]),
    .I1(bbar[11])
  );
  //AND U107
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U107 (
    .O(y[234]),
    .I0(a[14]),
    .I1(b[10])
  );
  //OR U107bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U107bar (
    .O(ybar[234]),
    .I0(abar[14]),
    .I1(bbar[10])
  );
  //AND U108
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U108 (
    .O(y[233]),
    .I0(a[14]),
    .I1(b[9])
  );
  //OR U108bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U108bar (
    .O(ybar[233]),
    .I0(abar[14]),
    .I1(bbar[9])
  );
  //AND U109
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U109 (
    .O(y[232]),
    .I0(a[14]),
    .I1(b[8])
  );
  //OR U109bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U109bar (
    .O(ybar[232]),
    .I0(abar[14]),
    .I1(bbar[8])
  );
  //AND U110
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U110 (
    .O(y[231]),
    .I0(a[14]),
    .I1(b[7])
  );
  //OR U110bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U110bar (
    .O(ybar[231]),
    .I0(abar[14]),
    .I1(bbar[7])
  );
  //AND U111
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U111 (
    .O(y[230]),
    .I0(a[14]),
    .I1(b[6])
  );
  //OR U111bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U111bar (
    .O(ybar[230]),
    .I0(abar[14]),
    .I1(bbar[6])
  );
  //AND U112
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U112 (
    .O(y[22]),
    .I0(a[1]),
    .I1(b[6])
  );
  //OR U112bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U112bar (
    .O(ybar[22]),
    .I0(abar[1]),
    .I1(bbar[6])
  );
  //AND U113
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U113 (
    .O(y[229]),
    .I0(a[14]),
    .I1(b[5])
  );
  //OR U113bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U113bar (
    .O(ybar[229]),
    .I0(abar[14]),
    .I1(bbar[5])
  );
  //AND U114
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U114 (
    .O(y[228]),
    .I0(a[14]),
    .I1(b[4])
  );
  //OR U114bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U114bar (
    .O(ybar[228]),
    .I0(abar[14]),
    .I1(bbar[4])
  );
  //AND U115
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U115 (
    .O(y[227]),
    .I0(a[14]),
    .I1(b[3])
  );
  //OR U115bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U115bar (
    .O(ybar[227]),
    .I0(abar[14]),
    .I1(bbar[3])
  );
  //AND U116
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U116 (
    .O(y[226]),
    .I0(a[14]),
    .I1(b[2])
  );
  //OR U116bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U116bar (
    .O(ybar[226]),
    .I0(abar[14]),
    .I1(bbar[2])
  );
  //AND U117
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U117 (
    .O(y[225]),
    .I0(a[14]),
    .I1(b[1])
  );
  //OR U117bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U117bar (
    .O(ybar[225]),
    .I0(abar[14]),
    .I1(bbar[1])
  );
  //AND U118
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U118 (
    .O(y[224]),
    .I0(a[14]),
    .I1(b[0])
  );
  //OR U118bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U118bar (
    .O(ybar[224]),
    .I0(abar[14]),
    .I1(bbar[0])
  );
  //AND U119
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U119 (
    .O(y[223]),
    .I0(a[13]),
    .I1(b[15])
  );
  //OR U119bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U119bar (
    .O(ybar[223]),
    .I0(abar[13]),
    .I1(bbar[15])
  );
  //AND U120
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U120 (
    .O(y[222]),
    .I0(a[13]),
    .I1(b[14])
  );
  //OR U120bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U120bar (
    .O(ybar[222]),
    .I0(abar[13]),
    .I1(bbar[14])
  );
  //AND U121
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U121 (
    .O(y[221]),
    .I0(a[13]),
    .I1(b[13])
  );
  //OR U121bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U121bar (
    .O(ybar[221]),
    .I0(abar[13]),
    .I1(bbar[13])
  );
  //AND U122
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U122 (
    .O(y[220]),
    .I0(a[13]),
    .I1(b[12])
  );
  //OR U122bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U122bar (
    .O(ybar[220]),
    .I0(abar[13]),
    .I1(bbar[12])
  );
  //AND U123
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U123 (
    .O(y[21]),
    .I0(a[1]),
    .I1(b[5])
  );
  //OR U123bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U123bar (
    .O(ybar[21]),
    .I0(abar[1]),
    .I1(bbar[5])
  );
  //AND U124
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U124 (
    .O(y[219]),
    .I0(a[13]),
    .I1(b[11])
  );
  //OR U124bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U124bar (
    .O(ybar[219]),
    .I0(abar[13]),
    .I1(bbar[11])
  );
  //AND U125
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U125 (
    .O(y[218]),
    .I0(a[13]),
    .I1(b[10])
  );
  //OR U125bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U125bar (
    .O(ybar[218]),
    .I0(abar[13]),
    .I1(bbar[10])
  );
  //AND U126
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U126 (
    .O(y[217]),
    .I0(a[13]),
    .I1(b[9])
  );
  //OR U126bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U126bar (
    .O(ybar[217]),
    .I0(abar[13]),
    .I1(bbar[9])
  );
  //AND U127
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U127 (
    .O(y[216]),
    .I0(a[13]),
    .I1(b[8])
  );
  //OR U127bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U127bar (
    .O(ybar[216]),
    .I0(abar[13]),
    .I1(bbar[8])
  );
  //AND U128
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U128 (
    .O(y[215]),
    .I0(a[13]),
    .I1(b[7])
  );
  //OR U128bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U128bar (
    .O(ybar[215]),
    .I0(abar[13]),
    .I1(bbar[7])
  );
  //AND U129
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U129 (
    .O(y[214]),
    .I0(a[13]),
    .I1(b[6])
  );
  //OR U129bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U129bar (
    .O(ybar[214]),
    .I0(abar[13]),
    .I1(bbar[6])
  );
  //AND U130
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U130 (
    .O(y[213]),
    .I0(a[13]),
    .I1(b[5])
  );
  //OR U130bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U130bar (
    .O(ybar[213]),
    .I0(abar[13]),
    .I1(bbar[5])
  );
  //AND U131
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U131 (
    .O(y[212]),
    .I0(a[13]),
    .I1(b[4])
  );
  //OR U131bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U131bar (
    .O(ybar[212]),
    .I0(abar[13]),
    .I1(bbar[4])
  );
  //AND U132
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U132 (
    .O(y[211]),
    .I0(a[13]),
    .I1(b[3])
  );
  //OR U132bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U132bar (
    .O(ybar[211]),
    .I0(abar[13]),
    .I1(bbar[3])
  );
  //AND U133
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U133 (
    .O(y[210]),
    .I0(a[13]),
    .I1(b[2])
  );
  //OR U133bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U133bar (
    .O(ybar[210]),
    .I0(abar[13]),
    .I1(bbar[2])
  );
  //AND U134
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U134 (
    .O(y[20]),
    .I0(a[1]),
    .I1(b[4])
  );
  //OR U134bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U134bar (
    .O(ybar[20]),
    .I0(abar[1]),
    .I1(bbar[4])
  );
  //AND U135
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U135 (
    .O(y[209]),
    .I0(a[13]),
    .I1(b[1])
  );
  //OR U135bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U135bar (
    .O(ybar[209]),
    .I0(abar[13]),
    .I1(bbar[1])
  );
  //AND U136
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U136 (
    .O(y[208]),
    .I0(a[13]),
    .I1(b[0])
  );
  //OR U136bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U136bar (
    .O(ybar[208]),
    .I0(abar[13]),
    .I1(bbar[0])
  );
  //AND U137
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U137 (
    .O(y[207]),
    .I0(a[12]),
    .I1(b[15])
  );
  //OR U137bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U137bar (
    .O(ybar[207]),
    .I0(abar[12]),
    .I1(bbar[15])
  );
  //AND U138
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U138 (
    .O(y[206]),
    .I0(a[12]),
    .I1(b[14])
  );
  //OR U138bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U138bar (
    .O(ybar[206]),
    .I0(abar[12]),
    .I1(bbar[14])
  );
  //AND U139
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U139 (
    .O(y[205]),
    .I0(a[12]),
    .I1(b[13])
  );
  //OR U139bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U139bar (
    .O(ybar[205]),
    .I0(abar[12]),
    .I1(bbar[13])
  );
  //AND U140
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U140 (
    .O(y[204]),
    .I0(a[12]),
    .I1(b[12])
  );
  //OR U140bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U140bar (
    .O(ybar[204]),
    .I0(abar[12]),
    .I1(bbar[12])
  );
  //AND U141
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U141 (
    .O(y[203]),
    .I0(a[12]),
    .I1(b[11])
  );
  //OR U141bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U141bar (
    .O(ybar[203]),
    .I0(abar[12]),
    .I1(bbar[11])
  );
  //AND U142
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U142 (
    .O(y[202]),
    .I0(a[12]),
    .I1(b[10])
  );
  //OR U142bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U142bar (
    .O(ybar[202]),
    .I0(abar[12]),
    .I1(bbar[10])
  );
  //AND U143
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U143 (
    .O(y[201]),
    .I0(a[12]),
    .I1(b[9])
  );
  //OR U143bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U143bar (
    .O(ybar[201]),
    .I0(abar[12]),
    .I1(bbar[9])
  );
  //AND U144
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U144 (
    .O(y[200]),
    .I0(a[12]),
    .I1(b[8])
  );
  //OR U144bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U144bar (
    .O(ybar[200]),
    .I0(abar[12]),
    .I1(bbar[8])
  );
  //AND U145
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U145 (
    .O(y[1]),
    .I0(b[1]),
    .I1(a[0])
  );
  //OR U145bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U145bar (
    .O(ybar[1]),
    .I0(bbar[1]),
    .I1(abar[0])
  );
  //AND U146
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U146 (
    .O(y[19]),
    .I0(a[1]),
    .I1(b[3])
  );
  //OR U146bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U146bar (
    .O(ybar[19]),
    .I0(abar[1]),
    .I1(bbar[3])
  );
  //AND U147
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U147 (
    .O(y[199]),
    .I0(a[12]),
    .I1(b[7])
  );
  //OR U147bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U147bar (
    .O(ybar[199]),
    .I0(abar[12]),
    .I1(bbar[7])
  );
  //AND U148
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U148 (
    .O(y[198]),
    .I0(a[12]),
    .I1(b[6])
  );
  //OR U148bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U148bar (
    .O(ybar[198]),
    .I0(abar[12]),
    .I1(bbar[6])
  );
  //AND U149
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U149 (
    .O(y[197]),
    .I0(a[12]),
    .I1(b[5])
  );
  //OR U149bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U149bar (
    .O(ybar[197]),
    .I0(abar[12]),
    .I1(bbar[5])
  );
  //AND U150
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U150 (
    .O(y[196]),
    .I0(a[12]),
    .I1(b[4])
  );
  //OR U150bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U150bar (
    .O(ybar[196]),
    .I0(abar[12]),
    .I1(bbar[4])
  );
  //AND U151
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U151 (
    .O(y[195]),
    .I0(a[12]),
    .I1(b[3])
  );
  //OR U151bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U151bar (
    .O(ybar[195]),
    .I0(abar[12]),
    .I1(bbar[3])
  );
  //AND U152
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U152 (
    .O(y[194]),
    .I0(a[12]),
    .I1(b[2])
  );
  //OR U152bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U152bar (
    .O(ybar[194]),
    .I0(abar[12]),
    .I1(bbar[2])
  );
  //AND U153
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U153 (
    .O(y[193]),
    .I0(a[12]),
    .I1(b[1])
  );
  //OR U153bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U153bar (
    .O(ybar[193]),
    .I0(abar[12]),
    .I1(bbar[1])
  );
  //AND U154
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U154 (
    .O(y[192]),
    .I0(a[12]),
    .I1(b[0])
  );
  //OR U154bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U154bar (
    .O(ybar[192]),
    .I0(abar[12]),
    .I1(bbar[0])
  );
  //AND U155
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U155 (
    .O(y[191]),
    .I0(a[11]),
    .I1(b[15])
  );
  //OR U155bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U155bar (
    .O(ybar[191]),
    .I0(abar[11]),
    .I1(bbar[15])
  );
  //AND U156
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U156 (
    .O(y[190]),
    .I0(a[11]),
    .I1(b[14])
  );
  //OR U156bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U156bar (
    .O(ybar[190]),
    .I0(abar[11]),
    .I1(bbar[14])
  );
  //AND U157
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U157 (
    .O(y[18]),
    .I0(a[1]),
    .I1(b[2])
  );
  //OR U157bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U157bar (
    .O(ybar[18]),
    .I0(abar[1]),
    .I1(bbar[2])
  );
  //AND U158
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U158 (
    .O(y[189]),
    .I0(a[11]),
    .I1(b[13])
  );
  //OR U158bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U158bar (
    .O(ybar[189]),
    .I0(abar[11]),
    .I1(bbar[13])
  );
  //AND U159
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U159 (
    .O(y[188]),
    .I0(a[11]),
    .I1(b[12])
  );
  //OR U159bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U159bar (
    .O(ybar[188]),
    .I0(abar[11]),
    .I1(bbar[12])
  );
  //AND U160
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U160 (
    .O(y[187]),
    .I0(a[11]),
    .I1(b[11])
  );
  //OR U160bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U160bar (
    .O(ybar[187]),
    .I0(abar[11]),
    .I1(bbar[11])
  );
  //AND U161
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U161 (
    .O(y[186]),
    .I0(a[11]),
    .I1(b[10])
  );
  //OR U161bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U161bar (
    .O(ybar[186]),
    .I0(abar[11]),
    .I1(bbar[10])
  );
  //AND U162
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U162 (
    .O(y[185]),
    .I0(a[11]),
    .I1(b[9])
  );
  //OR U162bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U162bar (
    .O(ybar[185]),
    .I0(abar[11]),
    .I1(bbar[9])
  );
  //AND U163
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U163 (
    .O(y[184]),
    .I0(a[11]),
    .I1(b[8])
  );
  //OR U163bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U163bar (
    .O(ybar[184]),
    .I0(abar[11]),
    .I1(bbar[8])
  );
  //AND U164
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U164 (
    .O(y[183]),
    .I0(a[11]),
    .I1(b[7])
  );
  //OR U164bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U164bar (
    .O(ybar[183]),
    .I0(abar[11]),
    .I1(bbar[7])
  );
  //AND U165
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U165 (
    .O(y[182]),
    .I0(a[11]),
    .I1(b[6])
  );
  //OR U165bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U165bar (
    .O(ybar[182]),
    .I0(abar[11]),
    .I1(bbar[6])
  );
  //AND U166
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U166 (
    .O(y[181]),
    .I0(a[11]),
    .I1(b[5])
  );
  //OR U166bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U166bar (
    .O(ybar[181]),
    .I0(abar[11]),
    .I1(bbar[5])
  );
  //AND U167
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U167 (
    .O(y[180]),
    .I0(a[11]),
    .I1(b[4])
  );
  //OR U167bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U167bar (
    .O(ybar[180]),
    .I0(abar[11]),
    .I1(bbar[4])
  );
  //AND U168
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U168 (
    .O(y[17]),
    .I0(a[1]),
    .I1(b[1])
  );
  //OR U168bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U168bar (
    .O(ybar[17]),
    .I0(abar[1]),
    .I1(bbar[1])
  );
  //AND U169
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U169 (
    .O(y[179]),
    .I0(a[11]),
    .I1(b[3])
  );
  //OR U169bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U169bar (
    .O(ybar[179]),
    .I0(abar[11]),
    .I1(bbar[3])
  );
  //AND U170
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U170 (
    .O(y[178]),
    .I0(a[11]),
    .I1(b[2])
  );
  //OR U170bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U170bar (
    .O(ybar[178]),
    .I0(abar[11]),
    .I1(bbar[2])
  );
  //AND U171
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U171 (
    .O(y[177]),
    .I0(a[11]),
    .I1(b[1])
  );
  //OR U171bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U171bar (
    .O(ybar[177]),
    .I0(abar[11]),
    .I1(bbar[1])
  );
  //AND U172
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U172 (
    .O(y[176]),
    .I0(a[11]),
    .I1(b[0])
  );
  //OR U172bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U172bar (
    .O(ybar[176]),
    .I0(abar[11]),
    .I1(bbar[0])
  );
  //AND U173
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U173 (
    .O(y[175]),
    .I0(a[10]),
    .I1(b[15])
  );
  //OR U173bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U173bar (
    .O(ybar[175]),
    .I0(abar[10]),
    .I1(bbar[15])
  );
  //AND U174
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U174 (
    .O(y[174]),
    .I0(a[10]),
    .I1(b[14])
  );
  //OR U174bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U174bar (
    .O(ybar[174]),
    .I0(abar[10]),
    .I1(bbar[14])
  );
  //AND U175
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U175 (
    .O(y[173]),
    .I0(a[10]),
    .I1(b[13])
  );
  //OR U175bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U175bar (
    .O(ybar[173]),
    .I0(abar[10]),
    .I1(bbar[13])
  );
  //AND U176
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U176 (
    .O(y[172]),
    .I0(a[10]),
    .I1(b[12])
  );
  //OR U176bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U176bar (
    .O(ybar[172]),
    .I0(abar[10]),
    .I1(bbar[12])
  );
  //AND U177
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U177 (
    .O(y[171]),
    .I0(a[10]),
    .I1(b[11])
  );
  //OR U177bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U177bar (
    .O(ybar[171]),
    .I0(abar[10]),
    .I1(bbar[11])
  );
  //AND U178
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U178 (
    .O(y[170]),
    .I0(a[10]),
    .I1(b[10])
  );
  //OR U178bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U178bar (
    .O(ybar[170]),
    .I0(abar[10]),
    .I1(bbar[10])
  );
  //AND U179
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U179 (
    .O(y[16]),
    .I0(a[1]),
    .I1(b[0])
  );
  //OR U179bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U179bar (
    .O(ybar[16]),
    .I0(abar[1]),
    .I1(bbar[0])
  );
  //AND U180
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U180 (
    .O(y[169]),
    .I0(a[10]),
    .I1(b[9])
  );
  //OR U180bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U180bar (
    .O(ybar[169]),
    .I0(abar[10]),
    .I1(bbar[9])
  );
  //AND U181
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U181 (
    .O(y[168]),
    .I0(a[10]),
    .I1(b[8])
  );
  //OR U181bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U181bar (
    .O(ybar[168]),
    .I0(abar[10]),
    .I1(bbar[8])
  );
  //AND U182
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U182 (
    .O(y[167]),
    .I0(a[10]),
    .I1(b[7])
  );
  //OR U182bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U182bar (
    .O(ybar[167]),
    .I0(abar[10]),
    .I1(bbar[7])
  );
  //AND U183
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U183 (
    .O(y[166]),
    .I0(a[10]),
    .I1(b[6])
  );
  //OR U183bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U183bar (
    .O(ybar[166]),
    .I0(abar[10]),
    .I1(bbar[6])
  );
  //AND U184
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U184 (
    .O(y[165]),
    .I0(a[10]),
    .I1(b[5])
  );
  //OR U184bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U184bar (
    .O(ybar[165]),
    .I0(abar[10]),
    .I1(bbar[5])
  );
  //AND U185
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U185 (
    .O(y[164]),
    .I0(a[10]),
    .I1(b[4])
  );
  //OR U185bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U185bar (
    .O(ybar[164]),
    .I0(abar[10]),
    .I1(bbar[4])
  );
  //AND U186
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U186 (
    .O(y[163]),
    .I0(a[10]),
    .I1(b[3])
  );
  //OR U186bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U186bar (
    .O(ybar[163]),
    .I0(abar[10]),
    .I1(bbar[3])
  );
  //AND U187
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U187 (
    .O(y[162]),
    .I0(a[10]),
    .I1(b[2])
  );
  //OR U187bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U187bar (
    .O(ybar[162]),
    .I0(abar[10]),
    .I1(bbar[2])
  );
  //AND U188
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U188 (
    .O(y[161]),
    .I0(a[10]),
    .I1(b[1])
  );
  //OR U188bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U188bar (
    .O(ybar[161]),
    .I0(abar[10]),
    .I1(bbar[1])
  );
  //AND U189
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U189 (
    .O(y[160]),
    .I0(a[10]),
    .I1(b[0])
  );
  //OR U189bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U189bar (
    .O(ybar[160]),
    .I0(abar[10]),
    .I1(bbar[0])
  );
  //AND U190
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U190 (
    .O(y[15]),
    .I0(b[15]),
    .I1(a[0])
  );
  //OR U190bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U190bar (
    .O(ybar[15]),
    .I0(bbar[15]),
    .I1(abar[0])
  );
  //AND U191
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U191 (
    .O(y[159]),
    .I0(a[9]),
    .I1(b[15])
  );
  //OR U191bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U191bar (
    .O(ybar[159]),
    .I0(abar[9]),
    .I1(bbar[15])
  );
  //AND U192
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U192 (
    .O(y[158]),
    .I0(a[9]),
    .I1(b[14])
  );
  //OR U192bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U192bar (
    .O(ybar[158]),
    .I0(abar[9]),
    .I1(bbar[14])
  );
  //AND U193
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U193 (
    .O(y[157]),
    .I0(a[9]),
    .I1(b[13])
  );
  //OR U193bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U193bar (
    .O(ybar[157]),
    .I0(abar[9]),
    .I1(bbar[13])
  );
  //AND U194
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U194 (
    .O(y[156]),
    .I0(a[9]),
    .I1(b[12])
  );
  //OR U194bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U194bar (
    .O(ybar[156]),
    .I0(abar[9]),
    .I1(bbar[12])
  );
  //AND U195
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U195 (
    .O(y[155]),
    .I0(a[9]),
    .I1(b[11])
  );
  //OR U195bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U195bar (
    .O(ybar[155]),
    .I0(abar[9]),
    .I1(bbar[11])
  );
  //AND U196
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U196 (
    .O(y[154]),
    .I0(a[9]),
    .I1(b[10])
  );
  //OR U196bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U196bar (
    .O(ybar[154]),
    .I0(abar[9]),
    .I1(bbar[10])
  );
  //AND U197
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U197 (
    .O(y[153]),
    .I0(a[9]),
    .I1(b[9])
  );
  //OR U197bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U197bar (
    .O(ybar[153]),
    .I0(abar[9]),
    .I1(bbar[9])
  );
  //AND U198
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U198 (
    .O(y[152]),
    .I0(a[9]),
    .I1(b[8])
  );
  //OR U198bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U198bar (
    .O(ybar[152]),
    .I0(abar[9]),
    .I1(bbar[8])
  );
  //AND U199
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U199 (
    .O(y[151]),
    .I0(a[9]),
    .I1(b[7])
  );
  //OR U199bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U199bar (
    .O(ybar[151]),
    .I0(abar[9]),
    .I1(bbar[7])
  );
  //AND U200
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U200 (
    .O(y[150]),
    .I0(a[9]),
    .I1(b[6])
  );
  //OR U200bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U200bar (
    .O(ybar[150]),
    .I0(abar[9]),
    .I1(bbar[6])
  );
  //AND U201
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U201 (
    .O(y[14]),
    .I0(b[14]),
    .I1(a[0])
  );
  //OR U201bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U201bar (
    .O(ybar[14]),
    .I0(bbar[14]),
    .I1(abar[0])
  );
  //AND U202
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U202 (
    .O(y[149]),
    .I0(a[9]),
    .I1(b[5])
  );
  //OR U202bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U202bar (
    .O(ybar[149]),
    .I0(abar[9]),
    .I1(bbar[5])
  );
  //AND U203
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U203 (
    .O(y[148]),
    .I0(a[9]),
    .I1(b[4])
  );
  //OR U203bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U203bar (
    .O(ybar[148]),
    .I0(abar[9]),
    .I1(bbar[4])
  );
  //AND U204
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U204 (
    .O(y[147]),
    .I0(a[9]),
    .I1(b[3])
  );
  //OR U204bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U204bar (
    .O(ybar[147]),
    .I0(abar[9]),
    .I1(bbar[3])
  );
  //AND U205
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U205 (
    .O(y[146]),
    .I0(a[9]),
    .I1(b[2])
  );
  //OR U205bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U205bar (
    .O(ybar[146]),
    .I0(abar[9]),
    .I1(bbar[2])
  );
  //AND U206
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U206 (
    .O(y[145]),
    .I0(a[9]),
    .I1(b[1])
  );
  //OR U206bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U206bar (
    .O(ybar[145]),
    .I0(abar[9]),
    .I1(bbar[1])
  );
  //AND U207
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U207 (
    .O(y[144]),
    .I0(a[9]),
    .I1(b[0])
  );
  //OR U207bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U207bar (
    .O(ybar[144]),
    .I0(abar[9]),
    .I1(bbar[0])
  );
  //AND U208
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U208 (
    .O(y[143]),
    .I0(a[8]),
    .I1(b[15])
  );
  //OR U208bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U208bar (
    .O(ybar[143]),
    .I0(abar[8]),
    .I1(bbar[15])
  );
  //AND U209
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U209 (
    .O(y[142]),
    .I0(a[8]),
    .I1(b[14])
  );
  //OR U209bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U209bar (
    .O(ybar[142]),
    .I0(abar[8]),
    .I1(bbar[14])
  );
  //AND U210
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U210 (
    .O(y[141]),
    .I0(a[8]),
    .I1(b[13])
  );
  //OR U210bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U210bar (
    .O(ybar[141]),
    .I0(abar[8]),
    .I1(bbar[13])
  );
  //AND U211
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U211 (
    .O(y[140]),
    .I0(a[8]),
    .I1(b[12])
  );
  //OR U211bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U211bar (
    .O(ybar[140]),
    .I0(abar[8]),
    .I1(bbar[12])
  );
  //AND U212
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U212 (
    .O(y[13]),
    .I0(b[13]),
    .I1(a[0])
  );
  //OR U212bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U212bar (
    .O(ybar[13]),
    .I0(bbar[13]),
    .I1(abar[0])
  );
  //AND U213
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U213 (
    .O(y[139]),
    .I0(a[8]),
    .I1(b[11])
  );
  //OR U213bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U213bar (
    .O(ybar[139]),
    .I0(abar[8]),
    .I1(bbar[11])
  );
  //AND U214
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U214 (
    .O(y[138]),
    .I0(a[8]),
    .I1(b[10])
  );
  //OR U214bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U214bar (
    .O(ybar[138]),
    .I0(abar[8]),
    .I1(bbar[10])
  );
  //AND U215
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U215 (
    .O(y[137]),
    .I0(a[8]),
    .I1(b[9])
  );
  //OR U215bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U215bar (
    .O(ybar[137]),
    .I0(abar[8]),
    .I1(bbar[9])
  );
  //AND U216
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U216 (
    .O(y[136]),
    .I0(a[8]),
    .I1(b[8])
  );
  //OR U216bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U216bar (
    .O(ybar[136]),
    .I0(abar[8]),
    .I1(bbar[8])
  );
  //AND U217
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U217 (
    .O(y[135]),
    .I0(a[8]),
    .I1(b[7])
  );
  //OR U217bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U217bar (
    .O(ybar[135]),
    .I0(abar[8]),
    .I1(bbar[7])
  );
  //AND U218
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U218 (
    .O(y[134]),
    .I0(a[8]),
    .I1(b[6])
  );
  //OR U218bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U218bar (
    .O(ybar[134]),
    .I0(abar[8]),
    .I1(bbar[6])
  );
  //AND U219
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U219 (
    .O(y[133]),
    .I0(a[8]),
    .I1(b[5])
  );
  //OR U219bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U219bar (
    .O(ybar[133]),
    .I0(abar[8]),
    .I1(bbar[5])
  );
  //AND U220
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U220 (
    .O(y[132]),
    .I0(a[8]),
    .I1(b[4])
  );
  //OR U220bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U220bar (
    .O(ybar[132]),
    .I0(abar[8]),
    .I1(bbar[4])
  );
  //AND U221
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U221 (
    .O(y[131]),
    .I0(a[8]),
    .I1(b[3])
  );
  //OR U221bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U221bar (
    .O(ybar[131]),
    .I0(abar[8]),
    .I1(bbar[3])
  );
  //AND U222
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U222 (
    .O(y[130]),
    .I0(a[8]),
    .I1(b[2])
  );
  //OR U222bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U222bar (
    .O(ybar[130]),
    .I0(abar[8]),
    .I1(bbar[2])
  );
  //AND U223
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U223 (
    .O(y[12]),
    .I0(b[12]),
    .I1(a[0])
  );
  //OR U223bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U223bar (
    .O(ybar[12]),
    .I0(bbar[12]),
    .I1(abar[0])
  );
  //AND U224
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U224 (
    .O(y[129]),
    .I0(a[8]),
    .I1(b[1])
  );
  //OR U224bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U224bar (
    .O(ybar[129]),
    .I0(abar[8]),
    .I1(bbar[1])
  );
  //AND U225
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U225 (
    .O(y[128]),
    .I0(a[8]),
    .I1(b[0])
  );
  //OR U225bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U225bar (
    .O(ybar[128]),
    .I0(abar[8]),
    .I1(bbar[0])
  );
  //AND U226
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U226 (
    .O(y[127]),
    .I0(a[7]),
    .I1(b[15])
  );
  //OR U226bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U226bar (
    .O(ybar[127]),
    .I0(abar[7]),
    .I1(bbar[15])
  );
  //AND U227
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U227 (
    .O(y[126]),
    .I0(a[7]),
    .I1(b[14])
  );
  //OR U227bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U227bar (
    .O(ybar[126]),
    .I0(abar[7]),
    .I1(bbar[14])
  );
  //AND U228
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U228 (
    .O(y[125]),
    .I0(a[7]),
    .I1(b[13])
  );
  //OR U228bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U228bar (
    .O(ybar[125]),
    .I0(abar[7]),
    .I1(bbar[13])
  );
  //AND U229
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U229 (
    .O(y[124]),
    .I0(a[7]),
    .I1(b[12])
  );
  //OR U229bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U229bar (
    .O(ybar[124]),
    .I0(abar[7]),
    .I1(bbar[12])
  );
  //AND U230
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U230 (
    .O(y[123]),
    .I0(a[7]),
    .I1(b[11])
  );
  //OR U230bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U230bar (
    .O(ybar[123]),
    .I0(abar[7]),
    .I1(bbar[11])
  );
  //AND U231
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U231 (
    .O(y[122]),
    .I0(a[7]),
    .I1(b[10])
  );
  //OR U231bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U231bar (
    .O(ybar[122]),
    .I0(abar[7]),
    .I1(bbar[10])
  );
  //AND U232
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U232 (
    .O(y[121]),
    .I0(a[7]),
    .I1(b[9])
  );
  //OR U232bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U232bar (
    .O(ybar[121]),
    .I0(abar[7]),
    .I1(bbar[9])
  );
  //AND U233
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U233 (
    .O(y[120]),
    .I0(a[7]),
    .I1(b[8])
  );
  //OR U233bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U233bar (
    .O(ybar[120]),
    .I0(abar[7]),
    .I1(bbar[8])
  );
  //AND U234
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U234 (
    .O(y[11]),
    .I0(b[11]),
    .I1(a[0])
  );
  //OR U234bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U234bar (
    .O(ybar[11]),
    .I0(bbar[11]),
    .I1(abar[0])
  );
  //AND U235
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U235 (
    .O(y[119]),
    .I0(a[7]),
    .I1(b[7])
  );
  //OR U235bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U235bar (
    .O(ybar[119]),
    .I0(abar[7]),
    .I1(bbar[7])
  );
  //AND U236
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U236 (
    .O(y[118]),
    .I0(a[7]),
    .I1(b[6])
  );
  //OR U236bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U236bar (
    .O(ybar[118]),
    .I0(abar[7]),
    .I1(bbar[6])
  );
  //AND U237
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U237 (
    .O(y[117]),
    .I0(a[7]),
    .I1(b[5])
  );
  //OR U237bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U237bar (
    .O(ybar[117]),
    .I0(abar[7]),
    .I1(bbar[5])
  );
  //AND U238
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U238 (
    .O(y[116]),
    .I0(a[7]),
    .I1(b[4])
  );
  //OR U238bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U238bar (
    .O(ybar[116]),
    .I0(abar[7]),
    .I1(bbar[4])
  );
  //AND U239
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U239 (
    .O(y[115]),
    .I0(a[7]),
    .I1(b[3])
  );
  //OR U239bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U239bar (
    .O(ybar[115]),
    .I0(abar[7]),
    .I1(bbar[3])
  );
  //AND U240
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U240 (
    .O(y[114]),
    .I0(a[7]),
    .I1(b[2])
  );
  //OR U240bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U240bar (
    .O(ybar[114]),
    .I0(abar[7]),
    .I1(bbar[2])
  );
  //AND U241
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U241 (
    .O(y[113]),
    .I0(a[7]),
    .I1(b[1])
  );
  //OR U241bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U241bar (
    .O(ybar[113]),
    .I0(abar[7]),
    .I1(bbar[1])
  );
  //AND U242
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U242 (
    .O(y[112]),
    .I0(a[7]),
    .I1(b[0])
  );
  //OR U242bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U242bar (
    .O(ybar[112]),
    .I0(abar[7]),
    .I1(bbar[0])
  );
  //AND U243
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U243 (
    .O(y[111]),
    .I0(b[15]),
    .I1(a[6])
  );
  //OR U243bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U243bar (
    .O(ybar[111]),
    .I0(bbar[15]),
    .I1(abar[6])
  );
  //AND U244
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U244 (
    .O(y[110]),
    .I0(b[14]),
    .I1(a[6])
  );
  //OR U244bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U244bar (
    .O(ybar[110]),
    .I0(bbar[14]),
    .I1(abar[6])
  );
  //AND U245
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U245 (
    .O(y[10]),
    .I0(b[10]),
    .I1(a[0])
  );
  //OR U245bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U245bar (
    .O(ybar[10]),
    .I0(bbar[10]),
    .I1(abar[0])
  );
  //AND U246
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U246 (
    .O(y[109]),
    .I0(b[13]),
    .I1(a[6])
  );
  //OR U246bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U246bar (
    .O(ybar[109]),
    .I0(bbar[13]),
    .I1(abar[6])
  );
  //AND U247
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U247 (
    .O(y[108]),
    .I0(b[12]),
    .I1(a[6])
  );
  //OR U247bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U247bar (
    .O(ybar[108]),
    .I0(bbar[12]),
    .I1(abar[6])
  );
  //AND U248
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U248 (
    .O(y[107]),
    .I0(b[11]),
    .I1(a[6])
  );
  //OR U248bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U248bar (
    .O(ybar[107]),
    .I0(bbar[11]),
    .I1(abar[6])
  );
  //AND U249
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U249 (
    .O(y[106]),
    .I0(b[10]),
    .I1(a[6])
  );
  //OR U249bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U249bar (
    .O(ybar[106]),
    .I0(bbar[10]),
    .I1(abar[6])
  );
  //AND U250
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U250 (
    .O(y[105]),
    .I0(a[6]),
    .I1(b[9])
  );
  //OR U250bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U250bar (
    .O(ybar[105]),
    .I0(abar[6]),
    .I1(bbar[9])
  );
  //AND U251
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U251 (
    .O(y[104]),
    .I0(b[8]),
    .I1(a[6])
  );
  //OR U251bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U251bar (
    .O(ybar[104]),
    .I0(bbar[8]),
    .I1(abar[6])
  );
  //AND U252
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U252 (
    .O(y[103]),
    .I0(b[7]),
    .I1(a[6])
  );
  //OR U252bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U252bar (
    .O(ybar[103]),
    .I0(bbar[7]),
    .I1(abar[6])
  );
  //AND U253
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U253 (
    .O(y[102]),
    .I0(b[6]),
    .I1(a[6])
  );
  //OR U253bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U253bar (
    .O(ybar[102]),
    .I0(bbar[6]),
    .I1(abar[6])
  );
  //AND U254
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U254 (
    .O(y[101]),
    .I0(b[5]),
    .I1(a[6])
  );
  //OR U254bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U254bar (
    .O(ybar[101]),
    .I0(bbar[5]),
    .I1(abar[6])
  );
  //AND U255
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U255 (
    .O(y[100]),
    .I0(b[4]),
    .I1(a[6])
  );
  //OR U255bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U255bar (
    .O(ybar[100]),
    .I0(bbar[4]),
    .I1(abar[6])
  );
  //AND U256
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U256 (
    .O(y[0]),
    .I0(b[0]),
    .I1(a[0])
  );
  //OR U256bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U256bar (
    .O(ybar[0]),
    .I0(bbar[0]),
    .I1(abar[0])
  );
endmodule

module decode_3 ( in, out );

  input wire [7:0] in;
//input_done

  output wire [255:0] out;
//output_done

  wire [15:0] level1;
  wire [31:0] level2;
//wire_done

  CD2_12 cd_l1_1 ( .a(in[1]), .b(in[0]), .y(level1[3:0]) );
  CD2_11 cd_l1_2 ( .a(in[3]), .b(in[2]), .y(level1[7:4]) );
  CD2_10 cd_l1_3 ( .a(in[5]), .b(in[4]), .y(level1[11:8]) );
  CD2_9 cd_l1_4 ( .a(in[7]), .b(in[6]), .y(level1[15:12]) );
  CD4_6 cd_l2_1 ( .a(level1[7:4]), .b(level1[3:0]), .y(level2[15:0]) );
  CD4_5 cd_l2_2 ( .a(level1[15:12]), .b(level1[11:8]), .y(level2[31:16]) );
  CD16_3 cd_l3 ( .a(level2[31:16]), .b(level2[15:0]), .y(out) );
endmodule

module encode_3 ( in, out );

  input wire [255:0] in;
  wire [255:0] inbar;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
  assign inbar[8] = ~in[8];
  assign inbar[9] = ~in[9];
  assign inbar[10] = ~in[10];
  assign inbar[11] = ~in[11];
  assign inbar[12] = ~in[12];
  assign inbar[13] = ~in[13];
  assign inbar[14] = ~in[14];
  assign inbar[15] = ~in[15];
  assign inbar[16] = ~in[16];
  assign inbar[17] = ~in[17];
  assign inbar[18] = ~in[18];
  assign inbar[19] = ~in[19];
  assign inbar[20] = ~in[20];
  assign inbar[21] = ~in[21];
  assign inbar[22] = ~in[22];
  assign inbar[23] = ~in[23];
  assign inbar[24] = ~in[24];
  assign inbar[25] = ~in[25];
  assign inbar[26] = ~in[26];
  assign inbar[27] = ~in[27];
  assign inbar[28] = ~in[28];
  assign inbar[29] = ~in[29];
  assign inbar[30] = ~in[30];
  assign inbar[31] = ~in[31];
  assign inbar[32] = ~in[32];
  assign inbar[33] = ~in[33];
  assign inbar[34] = ~in[34];
  assign inbar[35] = ~in[35];
  assign inbar[36] = ~in[36];
  assign inbar[37] = ~in[37];
  assign inbar[38] = ~in[38];
  assign inbar[39] = ~in[39];
  assign inbar[40] = ~in[40];
  assign inbar[41] = ~in[41];
  assign inbar[42] = ~in[42];
  assign inbar[43] = ~in[43];
  assign inbar[44] = ~in[44];
  assign inbar[45] = ~in[45];
  assign inbar[46] = ~in[46];
  assign inbar[47] = ~in[47];
  assign inbar[48] = ~in[48];
  assign inbar[49] = ~in[49];
  assign inbar[50] = ~in[50];
  assign inbar[51] = ~in[51];
  assign inbar[52] = ~in[52];
  assign inbar[53] = ~in[53];
  assign inbar[54] = ~in[54];
  assign inbar[55] = ~in[55];
  assign inbar[56] = ~in[56];
  assign inbar[57] = ~in[57];
  assign inbar[58] = ~in[58];
  assign inbar[59] = ~in[59];
  assign inbar[60] = ~in[60];
  assign inbar[61] = ~in[61];
  assign inbar[62] = ~in[62];
  assign inbar[63] = ~in[63];
  assign inbar[64] = ~in[64];
  assign inbar[65] = ~in[65];
  assign inbar[66] = ~in[66];
  assign inbar[67] = ~in[67];
  assign inbar[68] = ~in[68];
  assign inbar[69] = ~in[69];
  assign inbar[70] = ~in[70];
  assign inbar[71] = ~in[71];
  assign inbar[72] = ~in[72];
  assign inbar[73] = ~in[73];
  assign inbar[74] = ~in[74];
  assign inbar[75] = ~in[75];
  assign inbar[76] = ~in[76];
  assign inbar[77] = ~in[77];
  assign inbar[78] = ~in[78];
  assign inbar[79] = ~in[79];
  assign inbar[80] = ~in[80];
  assign inbar[81] = ~in[81];
  assign inbar[82] = ~in[82];
  assign inbar[83] = ~in[83];
  assign inbar[84] = ~in[84];
  assign inbar[85] = ~in[85];
  assign inbar[86] = ~in[86];
  assign inbar[87] = ~in[87];
  assign inbar[88] = ~in[88];
  assign inbar[89] = ~in[89];
  assign inbar[90] = ~in[90];
  assign inbar[91] = ~in[91];
  assign inbar[92] = ~in[92];
  assign inbar[93] = ~in[93];
  assign inbar[94] = ~in[94];
  assign inbar[95] = ~in[95];
  assign inbar[96] = ~in[96];
  assign inbar[97] = ~in[97];
  assign inbar[98] = ~in[98];
  assign inbar[99] = ~in[99];
  assign inbar[100] = ~in[100];
  assign inbar[101] = ~in[101];
  assign inbar[102] = ~in[102];
  assign inbar[103] = ~in[103];
  assign inbar[104] = ~in[104];
  assign inbar[105] = ~in[105];
  assign inbar[106] = ~in[106];
  assign inbar[107] = ~in[107];
  assign inbar[108] = ~in[108];
  assign inbar[109] = ~in[109];
  assign inbar[110] = ~in[110];
  assign inbar[111] = ~in[111];
  assign inbar[112] = ~in[112];
  assign inbar[113] = ~in[113];
  assign inbar[114] = ~in[114];
  assign inbar[115] = ~in[115];
  assign inbar[116] = ~in[116];
  assign inbar[117] = ~in[117];
  assign inbar[118] = ~in[118];
  assign inbar[119] = ~in[119];
  assign inbar[120] = ~in[120];
  assign inbar[121] = ~in[121];
  assign inbar[122] = ~in[122];
  assign inbar[123] = ~in[123];
  assign inbar[124] = ~in[124];
  assign inbar[125] = ~in[125];
  assign inbar[126] = ~in[126];
  assign inbar[127] = ~in[127];
  assign inbar[128] = ~in[128];
  assign inbar[129] = ~in[129];
  assign inbar[130] = ~in[130];
  assign inbar[131] = ~in[131];
  assign inbar[132] = ~in[132];
  assign inbar[133] = ~in[133];
  assign inbar[134] = ~in[134];
  assign inbar[135] = ~in[135];
  assign inbar[136] = ~in[136];
  assign inbar[137] = ~in[137];
  assign inbar[138] = ~in[138];
  assign inbar[139] = ~in[139];
  assign inbar[140] = ~in[140];
  assign inbar[141] = ~in[141];
  assign inbar[142] = ~in[142];
  assign inbar[143] = ~in[143];
  assign inbar[144] = ~in[144];
  assign inbar[145] = ~in[145];
  assign inbar[146] = ~in[146];
  assign inbar[147] = ~in[147];
  assign inbar[148] = ~in[148];
  assign inbar[149] = ~in[149];
  assign inbar[150] = ~in[150];
  assign inbar[151] = ~in[151];
  assign inbar[152] = ~in[152];
  assign inbar[153] = ~in[153];
  assign inbar[154] = ~in[154];
  assign inbar[155] = ~in[155];
  assign inbar[156] = ~in[156];
  assign inbar[157] = ~in[157];
  assign inbar[158] = ~in[158];
  assign inbar[159] = ~in[159];
  assign inbar[160] = ~in[160];
  assign inbar[161] = ~in[161];
  assign inbar[162] = ~in[162];
  assign inbar[163] = ~in[163];
  assign inbar[164] = ~in[164];
  assign inbar[165] = ~in[165];
  assign inbar[166] = ~in[166];
  assign inbar[167] = ~in[167];
  assign inbar[168] = ~in[168];
  assign inbar[169] = ~in[169];
  assign inbar[170] = ~in[170];
  assign inbar[171] = ~in[171];
  assign inbar[172] = ~in[172];
  assign inbar[173] = ~in[173];
  assign inbar[174] = ~in[174];
  assign inbar[175] = ~in[175];
  assign inbar[176] = ~in[176];
  assign inbar[177] = ~in[177];
  assign inbar[178] = ~in[178];
  assign inbar[179] = ~in[179];
  assign inbar[180] = ~in[180];
  assign inbar[181] = ~in[181];
  assign inbar[182] = ~in[182];
  assign inbar[183] = ~in[183];
  assign inbar[184] = ~in[184];
  assign inbar[185] = ~in[185];
  assign inbar[186] = ~in[186];
  assign inbar[187] = ~in[187];
  assign inbar[188] = ~in[188];
  assign inbar[189] = ~in[189];
  assign inbar[190] = ~in[190];
  assign inbar[191] = ~in[191];
  assign inbar[192] = ~in[192];
  assign inbar[193] = ~in[193];
  assign inbar[194] = ~in[194];
  assign inbar[195] = ~in[195];
  assign inbar[196] = ~in[196];
  assign inbar[197] = ~in[197];
  assign inbar[198] = ~in[198];
  assign inbar[199] = ~in[199];
  assign inbar[200] = ~in[200];
  assign inbar[201] = ~in[201];
  assign inbar[202] = ~in[202];
  assign inbar[203] = ~in[203];
  assign inbar[204] = ~in[204];
  assign inbar[205] = ~in[205];
  assign inbar[206] = ~in[206];
  assign inbar[207] = ~in[207];
  assign inbar[208] = ~in[208];
  assign inbar[209] = ~in[209];
  assign inbar[210] = ~in[210];
  assign inbar[211] = ~in[211];
  assign inbar[212] = ~in[212];
  assign inbar[213] = ~in[213];
  assign inbar[214] = ~in[214];
  assign inbar[215] = ~in[215];
  assign inbar[216] = ~in[216];
  assign inbar[217] = ~in[217];
  assign inbar[218] = ~in[218];
  assign inbar[219] = ~in[219];
  assign inbar[220] = ~in[220];
  assign inbar[221] = ~in[221];
  assign inbar[222] = ~in[222];
  assign inbar[223] = ~in[223];
  assign inbar[224] = ~in[224];
  assign inbar[225] = ~in[225];
  assign inbar[226] = ~in[226];
  assign inbar[227] = ~in[227];
  assign inbar[228] = ~in[228];
  assign inbar[229] = ~in[229];
  assign inbar[230] = ~in[230];
  assign inbar[231] = ~in[231];
  assign inbar[232] = ~in[232];
  assign inbar[233] = ~in[233];
  assign inbar[234] = ~in[234];
  assign inbar[235] = ~in[235];
  assign inbar[236] = ~in[236];
  assign inbar[237] = ~in[237];
  assign inbar[238] = ~in[238];
  assign inbar[239] = ~in[239];
  assign inbar[240] = ~in[240];
  assign inbar[241] = ~in[241];
  assign inbar[242] = ~in[242];
  assign inbar[243] = ~in[243];
  assign inbar[244] = ~in[244];
  assign inbar[245] = ~in[245];
  assign inbar[246] = ~in[246];
  assign inbar[247] = ~in[247];
  assign inbar[248] = ~in[248];
  assign inbar[249] = ~in[249];
  assign inbar[250] = ~in[250];
  assign inbar[251] = ~in[251];
  assign inbar[252] = ~in[252];
  assign inbar[253] = ~in[253];
  assign inbar[254] = ~in[254];
  assign inbar[255] = ~in[255];
//input_done

  output wire [7:0] out;
  wire [7:0] outbar;
//output_done

  wire in_81;
  wire in_80;
  wire in_79;
  wire in_78;
  wire in_77;
  wire in_76;
  wire in_75;
  wire in_74;
  wire in_73;
  wire in_72;
  wire in_71;
  wire in_70;
  wire in_69;
  wire in_68;
  wire in_67;
  wire in_66;
  wire in_65;
  wire in_64;
  wire in_63;
  wire in_62;
  wire in_61;
  wire in_60;
  wire in_59;
  wire in_58;
  wire in_57;
  wire in_56;
  wire in_55;
  wire in_54;
  wire in_53;
  wire in_52;
  wire in_51;
  wire in_50;
  wire in_49;
  wire in_48;
  wire in_47;
  wire in_46;
  wire in_45;
  wire in_44;
  wire in_43;
  wire in_42;
  wire in_41;
  wire in_40;
  wire in_39;
  wire in_38;
  wire in_37;
  wire in_36;
  wire in_35;
  wire in_34;
  wire in_33;
  wire in_32;
  wire in_31;
  wire in_30;
  wire in_29;
  wire in_28;
  wire in_27;
  wire in_26;
  wire in_25;
  wire in_24;
  wire in_23;
  wire in_22;
  wire in_21;
  wire in_20;
  wire in_19;
  wire in_18;
  wire in_17;
  wire in_16;
  wire in_15;
  wire in_14;
  wire in_13;
  wire in_12;
  wire in_11;
  wire in_10;
  wire in_9;
  wire in_8;
  wire in_7;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_3;
  wire in_2;
  wire in_1;
  wire in_0;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire in_81bar;
  wire in_80bar;
  wire in_79bar;
  wire in_78bar;
  wire in_77bar;
  wire in_76bar;
  wire in_75bar;
  wire in_74bar;
  wire in_73bar;
  wire in_72bar;
  wire in_71bar;
  wire in_70bar;
  wire in_69bar;
  wire in_68bar;
  wire in_67bar;
  wire in_66bar;
  wire in_65bar;
  wire in_64bar;
  wire in_63bar;
  wire in_62bar;
  wire in_61bar;
  wire in_60bar;
  wire in_59bar;
  wire in_58bar;
  wire in_57bar;
  wire in_56bar;
  wire in_55bar;
  wire in_54bar;
  wire in_53bar;
  wire in_52bar;
  wire in_51bar;
  wire in_50bar;
  wire in_49bar;
  wire in_48bar;
  wire in_47bar;
  wire in_46bar;
  wire in_45bar;
  wire in_44bar;
  wire in_43bar;
  wire in_42bar;
  wire in_41bar;
  wire in_40bar;
  wire in_39bar;
  wire in_38bar;
  wire in_37bar;
  wire in_36bar;
  wire in_35bar;
  wire in_34bar;
  wire in_33bar;
  wire in_32bar;
  wire in_31bar;
  wire in_30bar;
  wire in_29bar;
  wire in_28bar;
  wire in_27bar;
  wire in_26bar;
  wire in_25bar;
  wire in_24bar;
  wire in_23bar;
  wire in_22bar;
  wire in_21bar;
  wire in_20bar;
  wire in_19bar;
  wire in_18bar;
  wire in_17bar;
  wire in_16bar;
  wire in_15bar;
  wire in_14bar;
  wire in_13bar;
  wire in_12bar;
  wire in_11bar;
  wire in_10bar;
  wire in_9bar;
  wire in_8bar;
  wire in_7bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_3bar;
  wire in_2bar;
  wire in_1bar;
  wire in_0bar;
  wire n487bar;
  wire n488bar;
  wire n489bar;
  wire n490bar;
  wire n491bar;
  wire n492bar;
  wire n493bar;
  wire n494bar;
  wire n495bar;
  wire n496bar;
  wire n497bar;
  wire n498bar;
  wire n499bar;
  wire n500bar;
  wire n501bar;
  wire n502bar;
  wire n503bar;
  wire n504bar;
  wire n505bar;
  wire n506bar;
  wire n507bar;
  wire n508bar;
  wire n509bar;
  wire n510bar;
  wire n511bar;
  wire n512bar;
  wire n513bar;
  wire n514bar;
  wire n515bar;
  wire n516bar;
  wire n517bar;
  wire n518bar;
  wire n519bar;
  wire n520bar;
  wire n521bar;
  wire n522bar;
  wire n523bar;
  wire n524bar;
  wire n525bar;
  wire n526bar;
  wire n527bar;
  wire n528bar;
  wire n529bar;
  wire n530bar;
  wire n531bar;
  wire n532bar;
  wire n533bar;
  wire n534bar;
  wire n535bar;
  wire n536bar;
  wire n537bar;
  wire n538bar;
  wire n539bar;
  wire n540bar;
  wire n541bar;
  wire n542bar;
  wire n543bar;
  wire n544bar;
  wire n545bar;
  wire n546bar;
  wire n547bar;
  wire n548bar;
  wire n549bar;
  wire n550bar;
  wire n551bar;
  wire n552bar;
  wire n553bar;
  wire n554bar;
  wire n555bar;
  wire n556bar;
  wire n557bar;
  wire n558bar;
  wire n559bar;
  wire n560bar;
  wire n561bar;
  wire n562bar;
  wire n563bar;
  wire n564bar;
  wire n565bar;
  wire n566bar;
  wire n567bar;
  wire n568bar;
  wire n569bar;
  wire n570bar;
  wire n571bar;
  wire n572bar;
  wire n573bar;
  wire n574bar;
  wire n575bar;
  wire n576bar;
  wire n577bar;
  wire n578bar;
  wire n579bar;
  wire n580bar;
  wire n581bar;
  wire n582bar;
  wire n583bar;
  wire n584bar;
  wire n585bar;
  wire n586bar;
  wire n587bar;
  wire n588bar;
  wire n589bar;
  wire n590bar;
  wire n591bar;
  wire n592bar;
  wire n593bar;
  wire n594bar;
  wire n595bar;
  wire n596bar;
  wire n597bar;
  wire n598bar;
  wire n599bar;
  wire n600bar;
  wire n601bar;
  wire n602bar;
  wire n603bar;
  wire n604bar;
  wire n605bar;
  wire n606bar;
  wire n607bar;
  wire n608bar;
  wire n609bar;
  wire n610bar;
  wire n611bar;
  wire n612bar;
  wire n613bar;
  wire n614bar;
  wire n615bar;
  wire n616bar;
  wire n617bar;
  wire n618bar;
  wire n619bar;
  wire n620bar;
  wire n621bar;
  wire n622bar;
  wire n623bar;
  wire n624bar;
  wire n625bar;
  wire n626bar;
  wire n627bar;
  wire n628bar;
  wire n629bar;
  wire n630bar;
  wire n631bar;
  wire n632bar;
  wire n633bar;
  wire n634bar;
  wire n635bar;
  wire n636bar;
  wire n637bar;
  wire n638bar;
  wire n639bar;
  wire n640bar;
  wire n641bar;
  wire n642bar;
  wire n643bar;
  wire n644bar;
  wire n645bar;
  wire n646bar;
  wire n647bar;
  wire n648bar;
  wire n649bar;
  wire n650bar;
  wire n651bar;
  wire n652bar;
  wire n653bar;
  wire n654bar;
  wire n655bar;
  wire n656bar;
  wire n657bar;
  wire n658bar;
  wire n659bar;
  wire n660bar;
  wire n661bar;
  wire n662bar;
  wire n663bar;
  wire n664bar;
  wire n665bar;
  wire n666bar;
  wire n667bar;
  wire n668bar;
  wire n669bar;
  wire n670bar;
  wire n671bar;
  wire n672bar;
  wire n673bar;
  wire n674bar;
  wire n675bar;
  wire n676bar;
  wire n677bar;
  wire n678bar;
  wire n679bar;
  wire n680bar;
  wire n681bar;
  wire n682bar;
  wire n683bar;
  wire n684bar;
  wire n685bar;
  wire n686bar;
  wire n687bar;
  wire n688bar;
  wire n689bar;
  wire n690bar;
  wire n691bar;
  wire n692bar;
  wire n693bar;
  wire n694bar;
  wire n695bar;
  wire n696bar;
  wire n697bar;
  wire n698bar;
  wire n699bar;
  wire n700bar;
  wire n701bar;
  wire n702bar;
  wire n703bar;
  wire n704bar;
  wire n705bar;
  wire n706bar;
  wire n707bar;
  wire n708bar;
  wire n709bar;
  wire n710bar;
  wire n711bar;
  wire n712bar;
  wire n713bar;
  wire n714bar;
  wire n715bar;
  wire n716bar;
  wire n717bar;
  wire n718bar;
  wire n719bar;
  wire n720bar;
  wire n721bar;
  wire n722bar;
  wire n723bar;
  wire n724bar;
  wire n725bar;
  wire n726bar;
  wire n727bar;
  wire n728bar;
  wire n729bar;
  wire n730bar;
  wire n731bar;
  wire n732bar;
  wire n733bar;
  wire n734bar;
  wire n735bar;
  wire n736bar;
  wire n737bar;
  wire n738bar;
  wire n739bar;
  wire n740bar;
  wire n741bar;
  wire n742bar;
  wire n743bar;
  wire n744bar;
  wire n745bar;
  wire n746bar;
  wire n747bar;
  wire n748bar;
  wire n749bar;
  wire n750bar;
  wire n751bar;
  wire n752bar;
  wire n753bar;
  wire n754bar;
  wire n755bar;
  wire n756bar;
  wire n757bar;
  wire n758bar;
  wire n759bar;
  wire n760bar;
  wire n761bar;
  wire n762bar;
  wire n763bar;
  wire n764bar;
  wire n765bar;
  wire n766bar;
  wire n767bar;
  wire n768bar;
  wire n769bar;
  wire n770bar;
  wire n771bar;
  wire n772bar;
  wire n773bar;
  wire n774bar;
  wire n775bar;
  wire n776bar;
  wire n777bar;
  wire n778bar;
  wire n779bar;
  wire n780bar;
  wire n781bar;
  wire n782bar;
  wire n783bar;
  wire n784bar;
  wire n785bar;
  wire n786bar;
  wire n787bar;
  wire n788bar;
  wire n789bar;
  wire n790bar;
  wire n791bar;
  wire n792bar;
  wire n793bar;
  wire n794bar;
  wire n795bar;
  wire n796bar;
  wire n797bar;
  wire n798bar;
  wire n799bar;
  wire n800bar;
  wire n801bar;
  wire n802bar;
  wire n803bar;
  wire n804bar;
  wire n805bar;
  wire n806bar;
  wire n807bar;
  wire n808bar;
  wire n809bar;
  wire n810bar;
  wire n811bar;
  wire n812bar;
  wire n813bar;
  wire n814bar;
  wire n815bar;
  wire n816bar;
  wire n817bar;
  wire n818bar;
  wire n819bar;
  wire n820bar;
  wire n821bar;
  wire n822bar;
  wire n823bar;
  wire n824bar;
  wire n825bar;
  wire n826bar;
  wire n827bar;
  wire n828bar;
  wire n829bar;
  wire n830bar;
  wire n831bar;
  wire n832bar;
  wire n833bar;
  wire n834bar;
  wire n835bar;
  wire n836bar;
  wire n837bar;
  wire n838bar;
  wire n839bar;
  wire n840bar;
  wire n841bar;
  wire n842bar;
  wire n843bar;
  wire n844bar;
  wire n845bar;
  wire n846bar;
  wire n847bar;
  wire n848bar;
  wire n849bar;
  wire n850bar;
  wire n851bar;
  wire n852bar;
  wire n853bar;
  wire n854bar;
  wire n855bar;
  wire n856bar;
  wire n857bar;
  wire n858bar;
  wire n859bar;
  wire n860bar;
  wire n861bar;
  wire n862bar;
  wire n863bar;
  wire n864bar;
  wire n865bar;
  wire n866bar;
  wire n867bar;
  wire n868bar;
  wire n869bar;
  wire n870bar;
  wire n871bar;
  wire n872bar;
  wire n873bar;
  wire n874bar;
  wire n875bar;
  wire n876bar;
  wire n877bar;
  wire n878bar;
  wire n879bar;
  wire n880bar;
  wire n881bar;
  wire n882bar;
  wire n883bar;
  wire n884bar;
  wire n885bar;
  wire n886bar;
  wire n887bar;
  wire n888bar;
  wire n889bar;
  wire n890bar;
  wire n891bar;
  wire n892bar;
  wire n893bar;
  wire n894bar;
  wire n895bar;
  wire n896bar;
  wire n897bar;
  wire n898bar;
  wire n899bar;
  wire n900bar;
  wire n901bar;
  wire n902bar;
  wire n903bar;
  wire n904bar;
  wire n905bar;
  wire n906bar;
  wire n907bar;
  wire n908bar;
  wire n909bar;
  wire n910bar;
  wire n911bar;
  wire n912bar;
  wire n913bar;
  wire n914bar;
  wire n915bar;
  wire n916bar;
  wire n917bar;
  wire n918bar;
  wire n919bar;
  wire n920bar;
  wire n921bar;
  wire n922bar;
  wire n923bar;
  wire n924bar;
  wire n925bar;
  wire n926bar;
  wire n927bar;
  wire n928bar;
  wire n929bar;
  wire n930bar;
  wire n931bar;
  wire n932bar;
  wire n933bar;
  wire n934bar;
  wire n935bar;
  wire n936bar;
  wire n937bar;
  wire n938bar;
  wire n939bar;
  wire n940bar;
  wire n941bar;
  wire n942bar;
  wire n943bar;
  wire n944bar;
  wire n945bar;
  wire n946bar;
  wire n947bar;
  wire n948bar;
  wire n949bar;
  wire n950bar;
  wire n951bar;
  wire n952bar;
  wire n953bar;
  wire n954bar;
  wire n955bar;
  wire n956bar;
  wire n957bar;
  wire n958bar;
  wire n959bar;
  wire n960bar;
  wire n961bar;
  wire n962bar;
  wire n963bar;
  wire n964bar;
  wire n965bar;
  wire n966bar;
  wire n967bar;
  wire n968bar;
  wire n969bar;
  wire n970bar;
  wire n971bar;
  wire n972bar;
//wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];
  //OR U1
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1 (
    .O(out[7]),
    .I0(n972),
    .I1(n971)
  );
  //AND U1bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1bar (
    .O(outbar[7]),
    .I0(n972bar),
    .I1(n971bar)
  );
  //OR U2
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2 (
    .O(n971),
    .I0(n970),
    .I1(n969)
  );
  //AND U2bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2bar (
    .O(n971bar),
    .I0(n970bar),
    .I1(n969bar)
  );
  //OR U3
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3 (
    .O(n969),
    .I0(n968),
    .I1(n967)
  );
  //AND U3bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3bar (
    .O(n969bar),
    .I0(n968bar),
    .I1(n967bar)
  );
  //OR U4
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4 (
    .O(n967),
    .I0(n966),
    .I1(n965)
  );
  //AND U4bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4bar (
    .O(n967bar),
    .I0(n966bar),
    .I1(n965bar)
  );
  //OR U5
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5 (
    .O(n968),
    .I0(n964),
    .I1(n963)
  );
  //AND U5bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5bar (
    .O(n968bar),
    .I0(n964bar),
    .I1(n963bar)
  );
  //OR U6
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6 (
    .O(n963),
    .I0(in[116]),
    .I1(n962)
  );
  //AND U6bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6bar (
    .O(n963bar),
    .I0(inbar[116]),
    .I1(n962bar)
  );
  //OR U7
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7 (
    .O(n970),
    .I0(n961),
    .I1(n960)
  );
  //AND U7bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7bar (
    .O(n970bar),
    .I0(n961bar),
    .I1(n960bar)
  );
  //OR U8
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8 (
    .O(n960),
    .I0(in[150]),
    .I1(in[127])
  );
  //AND U8bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8bar (
    .O(n960bar),
    .I0(inbar[150]),
    .I1(inbar[127])
  );
  //OR U9
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9 (
    .O(n961),
    .I0(in[160]),
    .I1(n959)
  );
  //AND U9bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9bar (
    .O(n961bar),
    .I0(inbar[160]),
    .I1(n959bar)
  );
  //OR U10
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10 (
    .O(n959),
    .I0(in[252]),
    .I1(in[168])
  );
  //AND U10bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10bar (
    .O(n959bar),
    .I0(inbar[252]),
    .I1(inbar[168])
  );
  //OR U11
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11 (
    .O(n972),
    .I0(n958),
    .I1(n957)
  );
  //AND U11bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11bar (
    .O(n972bar),
    .I0(n958bar),
    .I1(n957bar)
  );
  //OR U12
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12 (
    .O(n957),
    .I0(n956),
    .I1(n955)
  );
  //AND U12bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12bar (
    .O(n957bar),
    .I0(n956bar),
    .I1(n955bar)
  );
  //OR U13
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13 (
    .O(n955),
    .I0(in_17),
    .I1(in[96])
  );
  //AND U13bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13bar (
    .O(n955bar),
    .I0(in_17bar),
    .I1(inbar[96])
  );
  //OR U14
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14 (
    .O(n956),
    .I0(in_23),
    .I1(n954)
  );
  //AND U14bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14bar (
    .O(n956bar),
    .I0(in_23bar),
    .I1(n954bar)
  );
  //OR U15
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15 (
    .O(n954),
    .I0(in_31),
    .I1(in_26)
  );
  //AND U15bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15bar (
    .O(n954bar),
    .I0(in_31bar),
    .I1(in_26bar)
  );
  //OR U16
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16 (
    .O(n958),
    .I0(n953),
    .I1(n952)
  );
  //AND U16bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16bar (
    .O(n958bar),
    .I0(n953bar),
    .I1(n952bar)
  );
  //OR U17
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U17 (
    .O(n952),
    .I0(in_58),
    .I1(in_4)
  );
  //AND U17bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U17bar (
    .O(n952bar),
    .I0(in_58bar),
    .I1(in_4bar)
  );
  //OR U18
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U18 (
    .O(n953),
    .I0(in_59),
    .I1(n951)
  );
  //AND U18bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U18bar (
    .O(n953bar),
    .I0(in_59bar),
    .I1(n951bar)
  );
  //OR U19
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U19 (
    .O(n951),
    .I0(in_71),
    .I1(in_62)
  );
  //AND U19bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U19bar (
    .O(n951bar),
    .I0(in_71bar),
    .I1(in_62bar)
  );
  //OR U20
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U20 (
    .O(out[6]),
    .I0(n950),
    .I1(n949)
  );
  //AND U20bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U20bar (
    .O(outbar[6]),
    .I0(n950bar),
    .I1(n949bar)
  );
  //OR U21
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U21 (
    .O(n949),
    .I0(n948),
    .I1(n947)
  );
  //AND U21bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U21bar (
    .O(n949bar),
    .I0(n948bar),
    .I1(n947bar)
  );
  //OR U22
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U22 (
    .O(n947),
    .I0(n946),
    .I1(n945)
  );
  //AND U22bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U22bar (
    .O(n947bar),
    .I0(n946bar),
    .I1(n945bar)
  );
  //OR U23
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U23 (
    .O(n945),
    .I0(n944),
    .I1(n943)
  );
  //AND U23bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U23bar (
    .O(n945bar),
    .I0(n944bar),
    .I1(n943bar)
  );
  //OR U24
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U24 (
    .O(n946),
    .I0(n942),
    .I1(n941)
  );
  //AND U24bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U24bar (
    .O(n946bar),
    .I0(n942bar),
    .I1(n941bar)
  );
  //OR U25
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U25 (
    .O(n941),
    .I0(in[101]),
    .I1(n940)
  );
  //AND U25bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U25bar (
    .O(n941bar),
    .I0(inbar[101]),
    .I1(n940bar)
  );
  //OR U26
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U26 (
    .O(n948),
    .I0(n939),
    .I1(n938)
  );
  //AND U26bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U26bar (
    .O(n948bar),
    .I0(n939bar),
    .I1(n938bar)
  );
  //OR U27
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U27 (
    .O(n938),
    .I0(in[114]),
    .I1(in[104])
  );
  //AND U27bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U27bar (
    .O(n938bar),
    .I0(inbar[114]),
    .I1(inbar[104])
  );
  //OR U28
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U28 (
    .O(n939),
    .I0(in[128]),
    .I1(n937)
  );
  //AND U28bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U28bar (
    .O(n939bar),
    .I0(inbar[128]),
    .I1(n937bar)
  );
  //OR U29
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U29 (
    .O(n937),
    .I0(in[136]),
    .I1(in[134])
  );
  //AND U29bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U29bar (
    .O(n937bar),
    .I0(inbar[136]),
    .I1(inbar[134])
  );
  //OR U30
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U30 (
    .O(n950),
    .I0(n936),
    .I1(n935)
  );
  //AND U30bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U30bar (
    .O(n950bar),
    .I0(n936bar),
    .I1(n935bar)
  );
  //OR U31
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U31 (
    .O(n935),
    .I0(n934),
    .I1(n933)
  );
  //AND U31bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U31bar (
    .O(n935bar),
    .I0(n934bar),
    .I1(n933bar)
  );
  //OR U32
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U32 (
    .O(n933),
    .I0(in[177]),
    .I1(in[164])
  );
  //AND U32bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U32bar (
    .O(n933bar),
    .I0(inbar[177]),
    .I1(inbar[164])
  );
  //OR U33
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U33 (
    .O(n934),
    .I0(in[212]),
    .I1(n932)
  );
  //AND U33bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U33bar (
    .O(n934bar),
    .I0(inbar[212]),
    .I1(n932bar)
  );
  //OR U34
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U34 (
    .O(n932),
    .I0(in[248]),
    .I1(in[221])
  );
  //AND U34bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U34bar (
    .O(n932bar),
    .I0(inbar[248]),
    .I1(inbar[221])
  );
  //OR U35
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U35 (
    .O(n936),
    .I0(n931),
    .I1(n930)
  );
  //AND U35bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U35bar (
    .O(n936bar),
    .I0(n931bar),
    .I1(n930bar)
  );
  //OR U36
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U36 (
    .O(n930),
    .I0(in_18),
    .I1(in[93])
  );
  //AND U36bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U36bar (
    .O(n930bar),
    .I0(in_18bar),
    .I1(inbar[93])
  );
  //OR U37
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U37 (
    .O(n931),
    .I0(in_31),
    .I1(n929)
  );
  //AND U37bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U37bar (
    .O(n931bar),
    .I0(in_31bar),
    .I1(n929bar)
  );
  //OR U38
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U38 (
    .O(n929),
    .I0(in_7),
    .I1(in_39)
  );
  //AND U38bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U38bar (
    .O(n929bar),
    .I0(in_7bar),
    .I1(in_39bar)
  );
  //OR U39
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U39 (
    .O(out[5]),
    .I0(n928),
    .I1(n927)
  );
  //AND U39bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U39bar (
    .O(outbar[5]),
    .I0(n928bar),
    .I1(n927bar)
  );
  //OR U40
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U40 (
    .O(n927),
    .I0(n926),
    .I1(n925)
  );
  //AND U40bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U40bar (
    .O(n927bar),
    .I0(n926bar),
    .I1(n925bar)
  );
  //OR U41
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U41 (
    .O(n925),
    .I0(n924),
    .I1(n923)
  );
  //AND U41bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U41bar (
    .O(n925bar),
    .I0(n924bar),
    .I1(n923bar)
  );
  //OR U42
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U42 (
    .O(n923),
    .I0(n922),
    .I1(n921)
  );
  //AND U42bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U42bar (
    .O(n923bar),
    .I0(n922bar),
    .I1(n921bar)
  );
  //OR U43
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U43 (
    .O(n924),
    .I0(n940),
    .I1(n920)
  );
  //AND U43bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U43bar (
    .O(n924bar),
    .I0(n940bar),
    .I1(n920bar)
  );
  //OR U44
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U44 (
    .O(n920),
    .I0(in[111]),
    .I1(n919)
  );
  //AND U44bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U44bar (
    .O(n920bar),
    .I0(inbar[111]),
    .I1(n919bar)
  );
  //OR U45
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U45 (
    .O(n940),
    .I0(n918),
    .I1(n917)
  );
  //AND U45bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U45bar (
    .O(n940bar),
    .I0(n918bar),
    .I1(n917bar)
  );
  //OR U46
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U46 (
    .O(n917),
    .I0(n916),
    .I1(n915)
  );
  //AND U46bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U46bar (
    .O(n917bar),
    .I0(n916bar),
    .I1(n915bar)
  );
  //OR U47
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U47 (
    .O(n915),
    .I0(n914),
    .I1(n913)
  );
  //AND U47bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U47bar (
    .O(n915bar),
    .I0(n914bar),
    .I1(n913bar)
  );
  //OR U48
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U48 (
    .O(n913),
    .I0(in[140]),
    .I1(in[131])
  );
  //AND U48bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U48bar (
    .O(n913bar),
    .I0(inbar[140]),
    .I1(inbar[131])
  );
  //OR U49
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U49 (
    .O(n914),
    .I0(in[160]),
    .I1(in[144])
  );
  //AND U49bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U49bar (
    .O(n914bar),
    .I0(inbar[160]),
    .I1(inbar[144])
  );
  //OR U50
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U50 (
    .O(n916),
    .I0(n912),
    .I1(n911)
  );
  //AND U50bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U50bar (
    .O(n916bar),
    .I0(n912bar),
    .I1(n911bar)
  );
  //OR U51
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U51 (
    .O(n911),
    .I0(in[179]),
    .I1(in[174])
  );
  //AND U51bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U51bar (
    .O(n911bar),
    .I0(inbar[179]),
    .I1(inbar[174])
  );
  //OR U52
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U52 (
    .O(n912),
    .I0(in[188]),
    .I1(in[184])
  );
  //AND U52bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U52bar (
    .O(n912bar),
    .I0(inbar[188]),
    .I1(inbar[184])
  );
  //OR U53
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U53 (
    .O(n918),
    .I0(n910),
    .I1(n909)
  );
  //AND U53bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U53bar (
    .O(n918bar),
    .I0(n910bar),
    .I1(n909bar)
  );
  //OR U54
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U54 (
    .O(n909),
    .I0(n908),
    .I1(n907)
  );
  //AND U54bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U54bar (
    .O(n909bar),
    .I0(n908bar),
    .I1(n907bar)
  );
  //OR U55
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U55 (
    .O(n907),
    .I0(in[216]),
    .I1(in[200])
  );
  //AND U55bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U55bar (
    .O(n907bar),
    .I0(inbar[216]),
    .I1(inbar[200])
  );
  //OR U56
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U56 (
    .O(n908),
    .I0(in[228]),
    .I1(in[224])
  );
  //AND U56bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U56bar (
    .O(n908bar),
    .I0(inbar[228]),
    .I1(inbar[224])
  );
  //OR U57
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U57 (
    .O(n910),
    .I0(n906),
    .I1(n905)
  );
  //AND U57bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U57bar (
    .O(n910bar),
    .I0(n906bar),
    .I1(n905bar)
  );
  //OR U58
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U58 (
    .O(n905),
    .I0(in[247]),
    .I1(in[235])
  );
  //AND U58bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U58bar (
    .O(n905bar),
    .I0(inbar[247]),
    .I1(inbar[235])
  );
  //OR U59
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U59 (
    .O(n906),
    .I0(in_42),
    .I1(in[83])
  );
  //AND U59bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U59bar (
    .O(n906bar),
    .I0(in_42bar),
    .I1(inbar[83])
  );
  //OR U60
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U60 (
    .O(n926),
    .I0(n904),
    .I1(n903)
  );
  //AND U60bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U60bar (
    .O(n926bar),
    .I0(n904bar),
    .I1(n903bar)
  );
  //OR U61
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U61 (
    .O(n903),
    .I0(in[166]),
    .I1(in[123])
  );
  //AND U61bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U61bar (
    .O(n903bar),
    .I0(inbar[166]),
    .I1(inbar[123])
  );
  //OR U62
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U62 (
    .O(n904),
    .I0(in[170]),
    .I1(n902)
  );
  //AND U62bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U62bar (
    .O(n904bar),
    .I0(inbar[170]),
    .I1(n902bar)
  );
  //OR U63
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U63 (
    .O(n902),
    .I0(in[194]),
    .I1(in[183])
  );
  //AND U63bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U63bar (
    .O(n902bar),
    .I0(inbar[194]),
    .I1(inbar[183])
  );
  //OR U64
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U64 (
    .O(n928),
    .I0(n901),
    .I1(n900)
  );
  //AND U64bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U64bar (
    .O(n928bar),
    .I0(n901bar),
    .I1(n900bar)
  );
  //OR U65
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U65 (
    .O(n900),
    .I0(n899),
    .I1(n898)
  );
  //AND U65bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U65bar (
    .O(n900bar),
    .I0(n899bar),
    .I1(n898bar)
  );
  //OR U66
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U66 (
    .O(n898),
    .I0(in[241]),
    .I1(in[238])
  );
  //AND U66bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U66bar (
    .O(n898bar),
    .I0(inbar[241]),
    .I1(inbar[238])
  );
  //OR U67
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U67 (
    .O(n899),
    .I0(in[250]),
    .I1(n897)
  );
  //AND U67bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U67bar (
    .O(n899bar),
    .I0(inbar[250]),
    .I1(n897bar)
  );
  //OR U68
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U68 (
    .O(n897),
    .I0(in_24),
    .I1(in[84])
  );
  //AND U68bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U68bar (
    .O(n897bar),
    .I0(in_24bar),
    .I1(inbar[84])
  );
  //OR U69
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U69 (
    .O(n901),
    .I0(n896),
    .I1(n895)
  );
  //AND U69bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U69bar (
    .O(n901bar),
    .I0(n896bar),
    .I1(n895bar)
  );
  //OR U70
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U70 (
    .O(n895),
    .I0(in_41),
    .I1(in_29)
  );
  //AND U70bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U70bar (
    .O(n895bar),
    .I0(in_41bar),
    .I1(in_29bar)
  );
  //OR U71
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U71 (
    .O(n896),
    .I0(in_66),
    .I1(n894)
  );
  //AND U71bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U71bar (
    .O(n896bar),
    .I0(in_66bar),
    .I1(n894bar)
  );
  //OR U72
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U72 (
    .O(n894),
    .I0(in_76),
    .I1(in_71)
  );
  //AND U72bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U72bar (
    .O(n894bar),
    .I0(in_76bar),
    .I1(in_71bar)
  );
  //OR U73
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U73 (
    .O(out[4]),
    .I0(n893),
    .I1(n892)
  );
  //AND U73bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U73bar (
    .O(outbar[4]),
    .I0(n893bar),
    .I1(n892bar)
  );
  //OR U74
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U74 (
    .O(n892),
    .I0(n891),
    .I1(n890)
  );
  //AND U74bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U74bar (
    .O(n892bar),
    .I0(n891bar),
    .I1(n890bar)
  );
  //OR U75
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U75 (
    .O(n890),
    .I0(n889),
    .I1(n888)
  );
  //AND U75bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U75bar (
    .O(n890bar),
    .I0(n889bar),
    .I1(n888bar)
  );
  //OR U76
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U76 (
    .O(n888),
    .I0(n922),
    .I1(n887)
  );
  //AND U76bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U76bar (
    .O(n888bar),
    .I0(n922bar),
    .I1(n887bar)
  );
  //OR U77
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U77 (
    .O(n922),
    .I0(n886),
    .I1(n885)
  );
  //AND U77bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U77bar (
    .O(n922bar),
    .I0(n886bar),
    .I1(n885bar)
  );
  //OR U78
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U78 (
    .O(n885),
    .I0(n884),
    .I1(n883)
  );
  //AND U78bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U78bar (
    .O(n885bar),
    .I0(n884bar),
    .I1(n883bar)
  );
  //OR U79
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U79 (
    .O(n883),
    .I0(n882),
    .I1(n881)
  );
  //AND U79bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U79bar (
    .O(n883bar),
    .I0(n882bar),
    .I1(n881bar)
  );
  //OR U80
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U80 (
    .O(n881),
    .I0(in[118]),
    .I1(in[109])
  );
  //AND U80bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U80bar (
    .O(n881bar),
    .I0(inbar[118]),
    .I1(inbar[109])
  );
  //OR U81
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U81 (
    .O(n882),
    .I0(in[139]),
    .I1(in[120])
  );
  //AND U81bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U81bar (
    .O(n882bar),
    .I0(inbar[139]),
    .I1(inbar[120])
  );
  //OR U82
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U82 (
    .O(n884),
    .I0(n880),
    .I1(n879)
  );
  //AND U82bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U82bar (
    .O(n884bar),
    .I0(n880bar),
    .I1(n879bar)
  );
  //OR U83
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U83 (
    .O(n879),
    .I0(in[198]),
    .I1(in[154])
  );
  //AND U83bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U83bar (
    .O(n879bar),
    .I0(inbar[198]),
    .I1(inbar[154])
  );
  //OR U84
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U84 (
    .O(n880),
    .I0(in[210]),
    .I1(in[205])
  );
  //AND U84bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U84bar (
    .O(n880bar),
    .I0(inbar[210]),
    .I1(inbar[205])
  );
  //OR U85
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U85 (
    .O(n886),
    .I0(n878),
    .I1(n877)
  );
  //AND U85bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U85bar (
    .O(n886bar),
    .I0(n878bar),
    .I1(n877bar)
  );
  //OR U86
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U86 (
    .O(n877),
    .I0(n876),
    .I1(n875)
  );
  //AND U86bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U86bar (
    .O(n877bar),
    .I0(n876bar),
    .I1(n875bar)
  );
  //OR U87
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U87 (
    .O(n875),
    .I0(in[219]),
    .I1(in[217])
  );
  //AND U87bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U87bar (
    .O(n875bar),
    .I0(inbar[219]),
    .I1(inbar[217])
  );
  //OR U88
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U88 (
    .O(n876),
    .I0(in[86]),
    .I1(in[252])
  );
  //AND U88bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U88bar (
    .O(n876bar),
    .I0(inbar[86]),
    .I1(inbar[252])
  );
  //OR U89
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U89 (
    .O(n878),
    .I0(n874),
    .I1(n873)
  );
  //AND U89bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U89bar (
    .O(n878bar),
    .I0(n874bar),
    .I1(n873bar)
  );
  //OR U90
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U90 (
    .O(n873),
    .I0(in_40),
    .I1(in[91])
  );
  //AND U90bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U90bar (
    .O(n873bar),
    .I0(in_40bar),
    .I1(inbar[91])
  );
  //OR U91
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U91 (
    .O(n874),
    .I0(in_8),
    .I1(in_46)
  );
  //AND U91bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U91bar (
    .O(n874bar),
    .I0(in_8bar),
    .I1(in_46bar)
  );
  //OR U92
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U92 (
    .O(n889),
    .I0(n872),
    .I1(n871)
  );
  //AND U92bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U92bar (
    .O(n889bar),
    .I0(n872bar),
    .I1(n871bar)
  );
  //OR U93
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U93 (
    .O(n871),
    .I0(in[117]),
    .I1(n943)
  );
  //AND U93bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U93bar (
    .O(n871bar),
    .I0(inbar[117]),
    .I1(n943bar)
  );
  //OR U94
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U94 (
    .O(n943),
    .I0(n870),
    .I1(n869)
  );
  //AND U94bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U94bar (
    .O(n943bar),
    .I0(n870bar),
    .I1(n869bar)
  );
  //OR U95
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U95 (
    .O(n869),
    .I0(n868),
    .I1(n867)
  );
  //AND U95bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U95bar (
    .O(n869bar),
    .I0(n868bar),
    .I1(n867bar)
  );
  //OR U96
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U96 (
    .O(n867),
    .I0(n866),
    .I1(n865)
  );
  //AND U96bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U96bar (
    .O(n867bar),
    .I0(n866bar),
    .I1(n865bar)
  );
  //OR U97
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U97 (
    .O(n865),
    .I0(n864),
    .I1(n863)
  );
  //AND U97bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U97bar (
    .O(n865bar),
    .I0(n864bar),
    .I1(n863bar)
  );
  //OR U98
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U98 (
    .O(n866),
    .I0(in[108]),
    .I1(n919)
  );
  //AND U98bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U98bar (
    .O(n866bar),
    .I0(inbar[108]),
    .I1(n919bar)
  );
  //OR U99
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U99 (
    .O(n919),
    .I0(n862),
    .I1(n861)
  );
  //AND U99bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U99bar (
    .O(n919bar),
    .I0(n862bar),
    .I1(n861bar)
  );
  //OR U100
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U100 (
    .O(n861),
    .I0(n860),
    .I1(n859)
  );
  //AND U100bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U100bar (
    .O(n861bar),
    .I0(n860bar),
    .I1(n859bar)
  );
  //OR U101
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U101 (
    .O(n859),
    .I0(n858),
    .I1(n857)
  );
  //AND U101bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U101bar (
    .O(n859bar),
    .I0(n858bar),
    .I1(n857bar)
  );
  //OR U102
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U102 (
    .O(n857),
    .I0(in[119]),
    .I1(in[105])
  );
  //AND U102bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U102bar (
    .O(n857bar),
    .I0(inbar[119]),
    .I1(inbar[105])
  );
  //OR U103
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U103 (
    .O(n858),
    .I0(in[186]),
    .I1(in[175])
  );
  //AND U103bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U103bar (
    .O(n858bar),
    .I0(inbar[186]),
    .I1(inbar[175])
  );
  //OR U104
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U104 (
    .O(n860),
    .I0(n856),
    .I1(n855)
  );
  //AND U104bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U104bar (
    .O(n860bar),
    .I0(n856bar),
    .I1(n855bar)
  );
  //OR U105
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U105 (
    .O(n855),
    .I0(in[202]),
    .I1(in[193])
  );
  //AND U105bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U105bar (
    .O(n855bar),
    .I0(inbar[202]),
    .I1(inbar[193])
  );
  //OR U106
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U106 (
    .O(n856),
    .I0(in[225]),
    .I1(in[208])
  );
  //AND U106bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U106bar (
    .O(n856bar),
    .I0(inbar[225]),
    .I1(inbar[208])
  );
  //OR U107
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U107 (
    .O(n862),
    .I0(n854),
    .I1(n853)
  );
  //AND U107bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U107bar (
    .O(n862bar),
    .I0(n854bar),
    .I1(n853bar)
  );
  //OR U108
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U108 (
    .O(n853),
    .I0(n852),
    .I1(n851)
  );
  //AND U108bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U108bar (
    .O(n853bar),
    .I0(n852bar),
    .I1(n851bar)
  );
  //OR U109
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U109 (
    .O(n851),
    .I0(in_1),
    .I1(in[85])
  );
  //AND U109bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U109bar (
    .O(n851bar),
    .I0(in_1bar),
    .I1(inbar[85])
  );
  //OR U110
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U110 (
    .O(n852),
    .I0(in_23),
    .I1(in_19)
  );
  //AND U110bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U110bar (
    .O(n852bar),
    .I0(in_23bar),
    .I1(in_19bar)
  );
  //OR U111
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U111 (
    .O(n854),
    .I0(n850),
    .I1(n849)
  );
  //AND U111bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U111bar (
    .O(n854bar),
    .I0(n850bar),
    .I1(n849bar)
  );
  //OR U112
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U112 (
    .O(n849),
    .I0(in_43),
    .I1(in_33)
  );
  //AND U112bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U112bar (
    .O(n849bar),
    .I0(in_43bar),
    .I1(in_33bar)
  );
  //OR U113
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U113 (
    .O(n850),
    .I0(in_63),
    .I1(in_44)
  );
  //AND U113bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U113bar (
    .O(n850bar),
    .I0(in_63bar),
    .I1(in_44bar)
  );
  //OR U114
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U114 (
    .O(n868),
    .I0(n848),
    .I1(n847)
  );
  //AND U114bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U114bar (
    .O(n868bar),
    .I0(n848bar),
    .I1(n847bar)
  );
  //OR U115
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U115 (
    .O(n847),
    .I0(in[141]),
    .I1(in[112])
  );
  //AND U115bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U115bar (
    .O(n847bar),
    .I0(inbar[141]),
    .I1(inbar[112])
  );
  //OR U116
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U116 (
    .O(n848),
    .I0(in[147]),
    .I1(n846)
  );
  //AND U116bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U116bar (
    .O(n848bar),
    .I0(inbar[147]),
    .I1(n846bar)
  );
  //OR U117
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U117 (
    .O(n846),
    .I0(in[181]),
    .I1(in[167])
  );
  //AND U117bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U117bar (
    .O(n846bar),
    .I0(inbar[181]),
    .I1(inbar[167])
  );
  //OR U118
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U118 (
    .O(n870),
    .I0(n845),
    .I1(n844)
  );
  //AND U118bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U118bar (
    .O(n870bar),
    .I0(n845bar),
    .I1(n844bar)
  );
  //OR U119
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U119 (
    .O(n844),
    .I0(n843),
    .I1(n842)
  );
  //AND U119bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U119bar (
    .O(n844bar),
    .I0(n843bar),
    .I1(n842bar)
  );
  //OR U120
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U120 (
    .O(n842),
    .I0(in[229]),
    .I1(in[201])
  );
  //AND U120bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U120bar (
    .O(n842bar),
    .I0(inbar[229]),
    .I1(inbar[201])
  );
  //OR U121
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U121 (
    .O(n843),
    .I0(in[237]),
    .I1(n841)
  );
  //AND U121bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U121bar (
    .O(n843bar),
    .I0(inbar[237]),
    .I1(n841bar)
  );
  //OR U122
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U122 (
    .O(n841),
    .I0(in[94]),
    .I1(in[253])
  );
  //AND U122bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U122bar (
    .O(n841bar),
    .I0(inbar[94]),
    .I1(inbar[253])
  );
  //OR U123
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U123 (
    .O(n845),
    .I0(n840),
    .I1(n839)
  );
  //AND U123bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U123bar (
    .O(n845bar),
    .I0(n840bar),
    .I1(n839bar)
  );
  //OR U124
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U124 (
    .O(n839),
    .I0(in_21),
    .I1(in[96])
  );
  //AND U124bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U124bar (
    .O(n839bar),
    .I0(in_21bar),
    .I1(inbar[96])
  );
  //OR U125
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U125 (
    .O(n840),
    .I0(in_25),
    .I1(n838)
  );
  //AND U125bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U125bar (
    .O(n840bar),
    .I0(in_25bar),
    .I1(n838bar)
  );
  //OR U126
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U126 (
    .O(n838),
    .I0(in_81),
    .I1(in_45)
  );
  //AND U126bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U126bar (
    .O(n838bar),
    .I0(in_81bar),
    .I1(in_45bar)
  );
  //OR U127
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U127 (
    .O(n891),
    .I0(n837),
    .I1(n836)
  );
  //AND U127bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U127bar (
    .O(n891bar),
    .I0(n837bar),
    .I1(n836bar)
  );
  //OR U128
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U128 (
    .O(n836),
    .I0(in[142]),
    .I1(in[124])
  );
  //AND U128bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U128bar (
    .O(n836bar),
    .I0(inbar[142]),
    .I1(inbar[124])
  );
  //OR U129
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U129 (
    .O(n837),
    .I0(in[150]),
    .I1(n835)
  );
  //AND U129bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U129bar (
    .O(n837bar),
    .I0(inbar[150]),
    .I1(n835bar)
  );
  //OR U130
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U130 (
    .O(n835),
    .I0(in[172]),
    .I1(in[155])
  );
  //AND U130bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U130bar (
    .O(n835bar),
    .I0(inbar[172]),
    .I1(inbar[155])
  );
  //OR U131
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U131 (
    .O(n893),
    .I0(n834),
    .I1(n833)
  );
  //AND U131bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U131bar (
    .O(n893bar),
    .I0(n834bar),
    .I1(n833bar)
  );
  //OR U132
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U132 (
    .O(n833),
    .I0(n832),
    .I1(n831)
  );
  //AND U132bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U132bar (
    .O(n833bar),
    .I0(n832bar),
    .I1(n831bar)
  );
  //OR U133
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U133 (
    .O(n831),
    .I0(in[196]),
    .I1(in[173])
  );
  //AND U133bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U133bar (
    .O(n831bar),
    .I0(inbar[196]),
    .I1(inbar[173])
  );
  //OR U134
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U134 (
    .O(n832),
    .I0(in[222]),
    .I1(n830)
  );
  //AND U134bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U134bar (
    .O(n832bar),
    .I0(inbar[222]),
    .I1(n830bar)
  );
  //OR U135
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U135 (
    .O(n830),
    .I0(in[227]),
    .I1(in[226])
  );
  //AND U135bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U135bar (
    .O(n830bar),
    .I0(inbar[227]),
    .I1(inbar[226])
  );
  //OR U136
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U136 (
    .O(n834),
    .I0(n829),
    .I1(n828)
  );
  //AND U136bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U136bar (
    .O(n834bar),
    .I0(n829bar),
    .I1(n828bar)
  );
  //OR U137
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U137 (
    .O(n828),
    .I0(in[249]),
    .I1(in[231])
  );
  //AND U137bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U137bar (
    .O(n828bar),
    .I0(inbar[249]),
    .I1(inbar[231])
  );
  //OR U138
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U138 (
    .O(n829),
    .I0(in_28),
    .I1(n827)
  );
  //AND U138bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U138bar (
    .O(n829bar),
    .I0(in_28bar),
    .I1(n827bar)
  );
  //OR U139
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U139 (
    .O(n827),
    .I0(in_52),
    .I1(in_47)
  );
  //AND U139bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U139bar (
    .O(n827bar),
    .I0(in_52bar),
    .I1(in_47bar)
  );
  //OR U140
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U140 (
    .O(out[3]),
    .I0(n826),
    .I1(n825)
  );
  //AND U140bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U140bar (
    .O(outbar[3]),
    .I0(n826bar),
    .I1(n825bar)
  );
  //OR U141
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U141 (
    .O(n825),
    .I0(n824),
    .I1(n823)
  );
  //AND U141bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U141bar (
    .O(n825bar),
    .I0(n824bar),
    .I1(n823bar)
  );
  //OR U142
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U142 (
    .O(n823),
    .I0(n822),
    .I1(n821)
  );
  //AND U142bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U142bar (
    .O(n823bar),
    .I0(n822bar),
    .I1(n821bar)
  );
  //OR U143
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U143 (
    .O(n821),
    .I0(n820),
    .I1(n819)
  );
  //AND U143bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U143bar (
    .O(n821bar),
    .I0(n820bar),
    .I1(n819bar)
  );
  //OR U144
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U144 (
    .O(n822),
    .I0(n964),
    .I1(n818)
  );
  //AND U144bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U144bar (
    .O(n822bar),
    .I0(n964bar),
    .I1(n818bar)
  );
  //OR U145
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U145 (
    .O(n818),
    .I0(in[118]),
    .I1(n817)
  );
  //AND U145bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U145bar (
    .O(n818bar),
    .I0(inbar[118]),
    .I1(n817bar)
  );
  //OR U146
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U146 (
    .O(n964),
    .I0(n816),
    .I1(n815)
  );
  //AND U146bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U146bar (
    .O(n964bar),
    .I0(n816bar),
    .I1(n815bar)
  );
  //OR U147
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U147 (
    .O(n815),
    .I0(n814),
    .I1(n813)
  );
  //AND U147bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U147bar (
    .O(n815bar),
    .I0(n814bar),
    .I1(n813bar)
  );
  //OR U148
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U148 (
    .O(n813),
    .I0(n812),
    .I1(n811)
  );
  //AND U148bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U148bar (
    .O(n813bar),
    .I0(n812bar),
    .I1(n811bar)
  );
  //OR U149
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U149 (
    .O(n811),
    .I0(in[122]),
    .I1(in[111])
  );
  //AND U149bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U149bar (
    .O(n811bar),
    .I0(inbar[122]),
    .I1(inbar[111])
  );
  //OR U150
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U150 (
    .O(n812),
    .I0(in[154]),
    .I1(in[151])
  );
  //AND U150bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U150bar (
    .O(n812bar),
    .I0(inbar[154]),
    .I1(inbar[151])
  );
  //OR U151
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U151 (
    .O(n814),
    .I0(n810),
    .I1(n809)
  );
  //AND U151bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U151bar (
    .O(n814bar),
    .I0(n810bar),
    .I1(n809bar)
  );
  //OR U152
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U152 (
    .O(n809),
    .I0(in[187]),
    .I1(in[177])
  );
  //AND U152bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U152bar (
    .O(n809bar),
    .I0(inbar[187]),
    .I1(inbar[177])
  );
  //OR U153
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U153 (
    .O(n810),
    .I0(in[200]),
    .I1(in[192])
  );
  //AND U153bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U153bar (
    .O(n810bar),
    .I0(inbar[200]),
    .I1(inbar[192])
  );
  //OR U154
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U154 (
    .O(n816),
    .I0(n808),
    .I1(n807)
  );
  //AND U154bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U154bar (
    .O(n816bar),
    .I0(n808bar),
    .I1(n807bar)
  );
  //OR U155
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U155 (
    .O(n807),
    .I0(n806),
    .I1(n805)
  );
  //AND U155bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U155bar (
    .O(n807bar),
    .I0(n806bar),
    .I1(n805bar)
  );
  //OR U156
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U156 (
    .O(n805),
    .I0(in[225]),
    .I1(in[207])
  );
  //AND U156bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U156bar (
    .O(n805bar),
    .I0(inbar[225]),
    .I1(inbar[207])
  );
  //OR U157
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U157 (
    .O(n806),
    .I0(in[98]),
    .I1(in[226])
  );
  //AND U157bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U157bar (
    .O(n806bar),
    .I0(inbar[98]),
    .I1(inbar[226])
  );
  //OR U158
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U158 (
    .O(n808),
    .I0(n804),
    .I1(n803)
  );
  //AND U158bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U158bar (
    .O(n808bar),
    .I0(n804bar),
    .I1(n803bar)
  );
  //OR U159
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U159 (
    .O(n803),
    .I0(in_20),
    .I1(in_16)
  );
  //AND U159bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U159bar (
    .O(n803bar),
    .I0(in_20bar),
    .I1(in_16bar)
  );
  //OR U160
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U160 (
    .O(n804),
    .I0(in_55),
    .I1(in_45)
  );
  //AND U160bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U160bar (
    .O(n804bar),
    .I0(in_55bar),
    .I1(in_45bar)
  );
  //OR U161
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U161 (
    .O(n824),
    .I0(n802),
    .I1(n801)
  );
  //AND U161bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U161bar (
    .O(n824bar),
    .I0(n802bar),
    .I1(n801bar)
  );
  //OR U162
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U162 (
    .O(n801),
    .I0(in[162]),
    .I1(in[149])
  );
  //AND U162bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U162bar (
    .O(n801bar),
    .I0(inbar[162]),
    .I1(inbar[149])
  );
  //OR U163
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U163 (
    .O(n802),
    .I0(in[163]),
    .I1(n800)
  );
  //AND U163bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U163bar (
    .O(n802bar),
    .I0(inbar[163]),
    .I1(n800bar)
  );
  //OR U164
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U164 (
    .O(n800),
    .I0(in[191]),
    .I1(in[189])
  );
  //AND U164bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U164bar (
    .O(n800bar),
    .I0(inbar[191]),
    .I1(inbar[189])
  );
  //OR U165
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U165 (
    .O(n826),
    .I0(n799),
    .I1(n798)
  );
  //AND U165bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U165bar (
    .O(n826bar),
    .I0(n799bar),
    .I1(n798bar)
  );
  //OR U166
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U166 (
    .O(n798),
    .I0(n797),
    .I1(n796)
  );
  //AND U166bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U166bar (
    .O(n798bar),
    .I0(n797bar),
    .I1(n796bar)
  );
  //OR U167
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U167 (
    .O(n796),
    .I0(in[212]),
    .I1(in[193])
  );
  //AND U167bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U167bar (
    .O(n796bar),
    .I0(inbar[212]),
    .I1(inbar[193])
  );
  //OR U168
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U168 (
    .O(n797),
    .I0(in[238]),
    .I1(n795)
  );
  //AND U168bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U168bar (
    .O(n797bar),
    .I0(inbar[238]),
    .I1(n795bar)
  );
  //OR U169
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U169 (
    .O(n795),
    .I0(in[88]),
    .I1(in[247])
  );
  //AND U169bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U169bar (
    .O(n795bar),
    .I0(inbar[88]),
    .I1(inbar[247])
  );
  //OR U170
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U170 (
    .O(n799),
    .I0(n794),
    .I1(n793)
  );
  //AND U170bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U170bar (
    .O(n799bar),
    .I0(n794bar),
    .I1(n793bar)
  );
  //OR U171
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U171 (
    .O(n793),
    .I0(in[94]),
    .I1(in[92])
  );
  //AND U171bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U171bar (
    .O(n793bar),
    .I0(inbar[94]),
    .I1(inbar[92])
  );
  //OR U172
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U172 (
    .O(n794),
    .I0(in_52),
    .I1(n792)
  );
  //AND U172bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U172bar (
    .O(n794bar),
    .I0(in_52bar),
    .I1(n792bar)
  );
  //OR U173
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U173 (
    .O(n792),
    .I0(in_70),
    .I1(in_67)
  );
  //AND U173bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U173bar (
    .O(n792bar),
    .I0(in_70bar),
    .I1(in_67bar)
  );
  //OR U174
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U174 (
    .O(out[2]),
    .I0(n791),
    .I1(n790)
  );
  //AND U174bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U174bar (
    .O(outbar[2]),
    .I0(n791bar),
    .I1(n790bar)
  );
  //OR U175
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U175 (
    .O(n790),
    .I0(n789),
    .I1(n788)
  );
  //AND U175bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U175bar (
    .O(n790bar),
    .I0(n789bar),
    .I1(n788bar)
  );
  //OR U176
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U176 (
    .O(n788),
    .I0(n787),
    .I1(n786)
  );
  //AND U176bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U176bar (
    .O(n788bar),
    .I0(n787bar),
    .I1(n786bar)
  );
  //OR U177
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U177 (
    .O(n786),
    .I0(n819),
    .I1(n785)
  );
  //AND U177bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U177bar (
    .O(n786bar),
    .I0(n819bar),
    .I1(n785bar)
  );
  //OR U178
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U178 (
    .O(n819),
    .I0(n784),
    .I1(n783)
  );
  //AND U178bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U178bar (
    .O(n819bar),
    .I0(n784bar),
    .I1(n783bar)
  );
  //OR U179
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U179 (
    .O(n783),
    .I0(n782),
    .I1(n781)
  );
  //AND U179bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U179bar (
    .O(n783bar),
    .I0(n782bar),
    .I1(n781bar)
  );
  //OR U180
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U180 (
    .O(n781),
    .I0(n780),
    .I1(n779)
  );
  //AND U180bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U180bar (
    .O(n781bar),
    .I0(n780bar),
    .I1(n779bar)
  );
  //OR U181
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U181 (
    .O(n779),
    .I0(n962),
    .I1(n778)
  );
  //AND U181bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U181bar (
    .O(n779bar),
    .I0(n962bar),
    .I1(n778bar)
  );
  //OR U182
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U182 (
    .O(n962),
    .I0(n777),
    .I1(n776)
  );
  //AND U182bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U182bar (
    .O(n962bar),
    .I0(n777bar),
    .I1(n776bar)
  );
  //OR U183
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U183 (
    .O(n776),
    .I0(n775),
    .I1(n774)
  );
  //AND U183bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U183bar (
    .O(n776bar),
    .I0(n775bar),
    .I1(n774bar)
  );
  //OR U184
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U184 (
    .O(n774),
    .I0(n773),
    .I1(n772)
  );
  //AND U184bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U184bar (
    .O(n774bar),
    .I0(n773bar),
    .I1(n772bar)
  );
  //OR U185
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U185 (
    .O(n772),
    .I0(in[131]),
    .I1(in[120])
  );
  //AND U185bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U185bar (
    .O(n772bar),
    .I0(inbar[131]),
    .I1(inbar[120])
  );
  //OR U186
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U186 (
    .O(n773),
    .I0(in[153]),
    .I1(in[147])
  );
  //AND U186bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U186bar (
    .O(n773bar),
    .I0(inbar[153]),
    .I1(inbar[147])
  );
  //OR U187
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U187 (
    .O(n775),
    .I0(n771),
    .I1(n770)
  );
  //AND U187bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U187bar (
    .O(n775bar),
    .I0(n771bar),
    .I1(n770bar)
  );
  //OR U188
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U188 (
    .O(n770),
    .I0(in[170]),
    .I1(in[156])
  );
  //AND U188bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U188bar (
    .O(n770bar),
    .I0(inbar[170]),
    .I1(inbar[156])
  );
  //OR U189
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U189 (
    .O(n771),
    .I0(in[223]),
    .I1(in[190])
  );
  //AND U189bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U189bar (
    .O(n771bar),
    .I0(inbar[223]),
    .I1(inbar[190])
  );
  //OR U190
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U190 (
    .O(n777),
    .I0(n769),
    .I1(n768)
  );
  //AND U190bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U190bar (
    .O(n777bar),
    .I0(n769bar),
    .I1(n768bar)
  );
  //OR U191
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U191 (
    .O(n768),
    .I0(n767),
    .I1(n766)
  );
  //AND U191bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U191bar (
    .O(n768bar),
    .I0(n767bar),
    .I1(n766bar)
  );
  //OR U192
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U192 (
    .O(n766),
    .I0(in[236]),
    .I1(in[230])
  );
  //AND U192bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U192bar (
    .O(n766bar),
    .I0(inbar[236]),
    .I1(inbar[230])
  );
  //OR U193
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U193 (
    .O(n767),
    .I0(in[85]),
    .I1(in[240])
  );
  //AND U193bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U193bar (
    .O(n767bar),
    .I0(inbar[85]),
    .I1(inbar[240])
  );
  //OR U194
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U194 (
    .O(n769),
    .I0(n765),
    .I1(n764)
  );
  //AND U194bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U194bar (
    .O(n769bar),
    .I0(n765bar),
    .I1(n764bar)
  );
  //OR U195
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U195 (
    .O(n764),
    .I0(in_12),
    .I1(in[90])
  );
  //AND U195bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U195bar (
    .O(n764bar),
    .I0(in_12bar),
    .I1(inbar[90])
  );
  //OR U196
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U196 (
    .O(n765),
    .I0(in_39),
    .I1(in_28)
  );
  //AND U196bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U196bar (
    .O(n765bar),
    .I0(in_39bar),
    .I1(in_28bar)
  );
  //OR U197
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U197 (
    .O(n780),
    .I0(in[109]),
    .I1(n763)
  );
  //AND U197bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U197bar (
    .O(n780bar),
    .I0(inbar[109]),
    .I1(n763bar)
  );
  //OR U198
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U198 (
    .O(n782),
    .I0(n762),
    .I1(n761)
  );
  //AND U198bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U198bar (
    .O(n782bar),
    .I0(n762bar),
    .I1(n761bar)
  );
  //OR U199
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U199 (
    .O(n761),
    .I0(in[138]),
    .I1(in[129])
  );
  //AND U199bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U199bar (
    .O(n761bar),
    .I0(inbar[138]),
    .I1(inbar[129])
  );
  //OR U200
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U200 (
    .O(n762),
    .I0(in[157]),
    .I1(n760)
  );
  //AND U200bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U200bar (
    .O(n762bar),
    .I0(inbar[157]),
    .I1(n760bar)
  );
  //OR U201
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U201 (
    .O(n760),
    .I0(in[182]),
    .I1(in[167])
  );
  //AND U201bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U201bar (
    .O(n760bar),
    .I0(inbar[182]),
    .I1(inbar[167])
  );
  //OR U202
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U202 (
    .O(n784),
    .I0(n759),
    .I1(n758)
  );
  //AND U202bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U202bar (
    .O(n784bar),
    .I0(n759bar),
    .I1(n758bar)
  );
  //OR U203
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U203 (
    .O(n758),
    .I0(n757),
    .I1(n756)
  );
  //AND U203bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U203bar (
    .O(n758bar),
    .I0(n757bar),
    .I1(n756bar)
  );
  //OR U204
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U204 (
    .O(n756),
    .I0(in[195]),
    .I1(in[184])
  );
  //AND U204bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U204bar (
    .O(n756bar),
    .I0(inbar[195]),
    .I1(inbar[184])
  );
  //OR U205
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U205 (
    .O(n757),
    .I0(in[196]),
    .I1(n755)
  );
  //AND U205bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U205bar (
    .O(n757bar),
    .I0(inbar[196]),
    .I1(n755bar)
  );
  //OR U206
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U206 (
    .O(n755),
    .I0(in[215]),
    .I1(in[209])
  );
  //AND U206bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U206bar (
    .O(n755bar),
    .I0(inbar[215]),
    .I1(inbar[209])
  );
  //OR U207
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U207 (
    .O(n759),
    .I0(n754),
    .I1(n753)
  );
  //AND U207bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U207bar (
    .O(n759bar),
    .I0(n754bar),
    .I1(n753bar)
  );
  //OR U208
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U208 (
    .O(n753),
    .I0(in[93]),
    .I1(in[233])
  );
  //AND U208bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U208bar (
    .O(n753bar),
    .I0(inbar[93]),
    .I1(inbar[233])
  );
  //OR U209
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U209 (
    .O(n754),
    .I0(in_1),
    .I1(n752)
  );
  //AND U209bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U209bar (
    .O(n754bar),
    .I0(in_1bar),
    .I1(n752bar)
  );
  //OR U210
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U210 (
    .O(n752),
    .I0(in_69),
    .I1(in_66)
  );
  //AND U210bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U210bar (
    .O(n752bar),
    .I0(in_69bar),
    .I1(in_66bar)
  );
  //OR U211
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U211 (
    .O(n787),
    .I0(n966),
    .I1(n751)
  );
  //AND U211bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U211bar (
    .O(n787bar),
    .I0(n966bar),
    .I1(n751bar)
  );
  //OR U212
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U212 (
    .O(n751),
    .I0(in[134]),
    .I1(n750)
  );
  //AND U212bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U212bar (
    .O(n751bar),
    .I0(inbar[134]),
    .I1(n750bar)
  );
  //OR U213
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U213 (
    .O(n966),
    .I0(n749),
    .I1(n748)
  );
  //AND U213bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U213bar (
    .O(n966bar),
    .I0(n749bar),
    .I1(n748bar)
  );
  //OR U214
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U214 (
    .O(n748),
    .I0(n747),
    .I1(n746)
  );
  //AND U214bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U214bar (
    .O(n748bar),
    .I0(n747bar),
    .I1(n746bar)
  );
  //OR U215
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U215 (
    .O(n746),
    .I0(n745),
    .I1(n744)
  );
  //AND U215bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U215bar (
    .O(n746bar),
    .I0(n745bar),
    .I1(n744bar)
  );
  //OR U216
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U216 (
    .O(n744),
    .I0(in[136]),
    .I1(in[121])
  );
  //AND U216bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U216bar (
    .O(n744bar),
    .I0(inbar[136]),
    .I1(inbar[121])
  );
  //OR U217
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U217 (
    .O(n745),
    .I0(in[186]),
    .I1(in[174])
  );
  //AND U217bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U217bar (
    .O(n745bar),
    .I0(inbar[186]),
    .I1(inbar[174])
  );
  //OR U218
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U218 (
    .O(n747),
    .I0(n743),
    .I1(n742)
  );
  //AND U218bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U218bar (
    .O(n747bar),
    .I0(n743bar),
    .I1(n742bar)
  );
  //OR U219
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U219 (
    .O(n742),
    .I0(in[198]),
    .I1(in[197])
  );
  //AND U219bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U219bar (
    .O(n742bar),
    .I0(inbar[198]),
    .I1(inbar[197])
  );
  //OR U220
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U220 (
    .O(n743),
    .I0(in[214]),
    .I1(in[199])
  );
  //AND U220bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U220bar (
    .O(n743bar),
    .I0(inbar[214]),
    .I1(inbar[199])
  );
  //OR U221
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U221 (
    .O(n749),
    .I0(n741),
    .I1(n740)
  );
  //AND U221bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U221bar (
    .O(n749bar),
    .I0(n741bar),
    .I1(n740bar)
  );
  //OR U222
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U222 (
    .O(n740),
    .I0(n739),
    .I1(n738)
  );
  //AND U222bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U222bar (
    .O(n740bar),
    .I0(n739bar),
    .I1(n738bar)
  );
  //OR U223
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U223 (
    .O(n738),
    .I0(in[231]),
    .I1(in[220])
  );
  //AND U223bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U223bar (
    .O(n738bar),
    .I0(inbar[231]),
    .I1(inbar[220])
  );
  //OR U224
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U224 (
    .O(n739),
    .I0(in_25),
    .I1(in[245])
  );
  //AND U224bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U224bar (
    .O(n739bar),
    .I0(in_25bar),
    .I1(inbar[245])
  );
  //OR U225
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U225 (
    .O(n741),
    .I0(n737),
    .I1(n736)
  );
  //AND U225bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U225bar (
    .O(n741bar),
    .I0(n737bar),
    .I1(n736bar)
  );
  //OR U226
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U226 (
    .O(n736),
    .I0(in_53),
    .I1(in_29)
  );
  //AND U226bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U226bar (
    .O(n736bar),
    .I0(in_53bar),
    .I1(in_29bar)
  );
  //OR U227
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U227 (
    .O(n737),
    .I0(in_79),
    .I1(in_74)
  );
  //AND U227bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U227bar (
    .O(n737bar),
    .I0(in_79bar),
    .I1(in_74bar)
  );
  //OR U228
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U228 (
    .O(n789),
    .I0(n735),
    .I1(n734)
  );
  //AND U228bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U228bar (
    .O(n789bar),
    .I0(n735bar),
    .I1(n734bar)
  );
  //OR U229
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U229 (
    .O(n734),
    .I0(in[152]),
    .I1(in[140])
  );
  //AND U229bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U229bar (
    .O(n734bar),
    .I0(inbar[152]),
    .I1(inbar[140])
  );
  //OR U230
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U230 (
    .O(n735),
    .I0(in[155]),
    .I1(n733)
  );
  //AND U230bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U230bar (
    .O(n735bar),
    .I0(inbar[155]),
    .I1(n733bar)
  );
  //OR U231
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U231 (
    .O(n733),
    .I0(in[166]),
    .I1(in[165])
  );
  //AND U231bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U231bar (
    .O(n733bar),
    .I0(inbar[166]),
    .I1(inbar[165])
  );
  //OR U232
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U232 (
    .O(n791),
    .I0(n732),
    .I1(n731)
  );
  //AND U232bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U232bar (
    .O(n791bar),
    .I0(n732bar),
    .I1(n731bar)
  );
  //OR U233
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U233 (
    .O(n731),
    .I0(n730),
    .I1(n729)
  );
  //AND U233bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U233bar (
    .O(n731bar),
    .I0(n730bar),
    .I1(n729bar)
  );
  //OR U234
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U234 (
    .O(n729),
    .I0(in[202]),
    .I1(in[185])
  );
  //AND U234bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U234bar (
    .O(n729bar),
    .I0(inbar[202]),
    .I1(inbar[185])
  );
  //OR U235
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U235 (
    .O(n730),
    .I0(in[211]),
    .I1(n728)
  );
  //AND U235bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U235bar (
    .O(n730bar),
    .I0(inbar[211]),
    .I1(n728bar)
  );
  //OR U236
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U236 (
    .O(n728),
    .I0(in[255]),
    .I1(in[253])
  );
  //AND U236bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U236bar (
    .O(n728bar),
    .I0(inbar[255]),
    .I1(inbar[253])
  );
  //OR U237
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U237 (
    .O(n732),
    .I0(n727),
    .I1(n726)
  );
  //AND U237bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U237bar (
    .O(n732bar),
    .I0(n727bar),
    .I1(n726bar)
  );
  //OR U238
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U238 (
    .O(n726),
    .I0(in_35),
    .I1(in_15)
  );
  //AND U238bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U238bar (
    .O(n726bar),
    .I0(in_35bar),
    .I1(in_15bar)
  );
  //OR U239
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U239 (
    .O(n727),
    .I0(in_36),
    .I1(n725)
  );
  //AND U239bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U239bar (
    .O(n727bar),
    .I0(in_36bar),
    .I1(n725bar)
  );
  //OR U240
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U240 (
    .O(n725),
    .I0(in_48),
    .I1(in_40)
  );
  //AND U240bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U240bar (
    .O(n725bar),
    .I0(in_48bar),
    .I1(in_40bar)
  );
  //OR U241
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U241 (
    .O(out[1]),
    .I0(n724),
    .I1(n723)
  );
  //AND U241bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U241bar (
    .O(outbar[1]),
    .I0(n724bar),
    .I1(n723bar)
  );
  //OR U242
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U242 (
    .O(n723),
    .I0(n722),
    .I1(n721)
  );
  //AND U242bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U242bar (
    .O(n723bar),
    .I0(n722bar),
    .I1(n721bar)
  );
  //OR U243
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U243 (
    .O(n721),
    .I0(n720),
    .I1(n719)
  );
  //AND U243bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U243bar (
    .O(n721bar),
    .I0(n720bar),
    .I1(n719bar)
  );
  //OR U244
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U244 (
    .O(n719),
    .I0(n921),
    .I1(n887)
  );
  //AND U244bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U244bar (
    .O(n719bar),
    .I0(n921bar),
    .I1(n887bar)
  );
  //OR U245
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U245 (
    .O(n887),
    .I0(n718),
    .I1(n717)
  );
  //AND U245bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U245bar (
    .O(n887bar),
    .I0(n718bar),
    .I1(n717bar)
  );
  //OR U246
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U246 (
    .O(n717),
    .I0(n716),
    .I1(n715)
  );
  //AND U246bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U246bar (
    .O(n717bar),
    .I0(n716bar),
    .I1(n715bar)
  );
  //OR U247
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U247 (
    .O(n715),
    .I0(n714),
    .I1(n713)
  );
  //AND U247bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U247bar (
    .O(n715bar),
    .I0(n714bar),
    .I1(n713bar)
  );
  //OR U248
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U248 (
    .O(n713),
    .I0(in[116]),
    .I1(in[110])
  );
  //AND U248bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U248bar (
    .O(n713bar),
    .I0(inbar[116]),
    .I1(inbar[110])
  );
  //OR U249
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U249 (
    .O(n714),
    .I0(in[133]),
    .I1(in[130])
  );
  //AND U249bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U249bar (
    .O(n714bar),
    .I0(inbar[133]),
    .I1(inbar[130])
  );
  //OR U250
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U250 (
    .O(n716),
    .I0(n712),
    .I1(n711)
  );
  //AND U250bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U250bar (
    .O(n716bar),
    .I0(n712bar),
    .I1(n711bar)
  );
  //OR U251
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U251 (
    .O(n711),
    .I0(in[203]),
    .I1(in[135])
  );
  //AND U251bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U251bar (
    .O(n711bar),
    .I0(inbar[203]),
    .I1(inbar[135])
  );
  //OR U252
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U252 (
    .O(n712),
    .I0(in[232]),
    .I1(in[223])
  );
  //AND U252bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U252bar (
    .O(n712bar),
    .I0(inbar[232]),
    .I1(inbar[223])
  );
  //OR U253
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U253 (
    .O(n718),
    .I0(n710),
    .I1(n709)
  );
  //AND U253bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U253bar (
    .O(n718bar),
    .I0(n710bar),
    .I1(n709bar)
  );
  //OR U254
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U254 (
    .O(n709),
    .I0(n708),
    .I1(n707)
  );
  //AND U254bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U254bar (
    .O(n709bar),
    .I0(n708bar),
    .I1(n707bar)
  );
  //OR U255
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U255 (
    .O(n707),
    .I0(in[255]),
    .I1(in[233])
  );
  //AND U255bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U255bar (
    .O(n707bar),
    .I0(inbar[255]),
    .I1(inbar[233])
  );
  //OR U256
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U256 (
    .O(n708),
    .I0(in_53),
    .I1(in_34)
  );
  //AND U256bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U256bar (
    .O(n708bar),
    .I0(in_53bar),
    .I1(in_34bar)
  );
  //OR U257
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U257 (
    .O(n710),
    .I0(n706),
    .I1(n705)
  );
  //AND U257bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U257bar (
    .O(n710bar),
    .I0(n706bar),
    .I1(n705bar)
  );
  //OR U258
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U258 (
    .O(n705),
    .I0(in_57),
    .I1(in_55)
  );
  //AND U258bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U258bar (
    .O(n705bar),
    .I0(in_57bar),
    .I1(in_55bar)
  );
  //OR U259
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U259 (
    .O(n706),
    .I0(in_68),
    .I1(in_67)
  );
  //AND U259bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U259bar (
    .O(n706bar),
    .I0(in_68bar),
    .I1(in_67bar)
  );
  //OR U260
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U260 (
    .O(n921),
    .I0(n704),
    .I1(n703)
  );
  //AND U260bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U260bar (
    .O(n921bar),
    .I0(n704bar),
    .I1(n703bar)
  );
  //OR U261
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U261 (
    .O(n703),
    .I0(n702),
    .I1(n701)
  );
  //AND U261bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U261bar (
    .O(n703bar),
    .I0(n702bar),
    .I1(n701bar)
  );
  //OR U262
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U262 (
    .O(n701),
    .I0(n700),
    .I1(n699)
  );
  //AND U262bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U262bar (
    .O(n701bar),
    .I0(n700bar),
    .I1(n699bar)
  );
  //OR U263
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U263 (
    .O(n699),
    .I0(n944),
    .I1(n872)
  );
  //AND U263bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U263bar (
    .O(n699bar),
    .I0(n944bar),
    .I1(n872bar)
  );
  //OR U264
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U264 (
    .O(n872),
    .I0(n698),
    .I1(n697)
  );
  //AND U264bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U264bar (
    .O(n872bar),
    .I0(n698bar),
    .I1(n697bar)
  );
  //OR U265
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U265 (
    .O(n697),
    .I0(n696),
    .I1(n695)
  );
  //AND U265bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U265bar (
    .O(n697bar),
    .I0(n696bar),
    .I1(n695bar)
  );
  //OR U266
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U266 (
    .O(n695),
    .I0(n694),
    .I1(n693)
  );
  //AND U266bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U266bar (
    .O(n695bar),
    .I0(n694bar),
    .I1(n693bar)
  );
  //OR U267
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U267 (
    .O(n693),
    .I0(in[121]),
    .I1(in[102])
  );
  //AND U267bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U267bar (
    .O(n693bar),
    .I0(inbar[121]),
    .I1(inbar[102])
  );
  //OR U268
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U268 (
    .O(n694),
    .I0(in[162]),
    .I1(in[161])
  );
  //AND U268bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U268bar (
    .O(n694bar),
    .I0(inbar[162]),
    .I1(inbar[161])
  );
  //OR U269
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U269 (
    .O(n696),
    .I0(n692),
    .I1(n691)
  );
  //AND U269bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U269bar (
    .O(n696bar),
    .I0(n692bar),
    .I1(n691bar)
  );
  //OR U270
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U270 (
    .O(n691),
    .I0(in[192]),
    .I1(in[178])
  );
  //AND U270bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U270bar (
    .O(n691bar),
    .I0(inbar[192]),
    .I1(inbar[178])
  );
  //OR U271
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U271 (
    .O(n692),
    .I0(in[244]),
    .I1(in[209])
  );
  //AND U271bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U271bar (
    .O(n692bar),
    .I0(inbar[244]),
    .I1(inbar[209])
  );
  //OR U272
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U272 (
    .O(n698),
    .I0(n690),
    .I1(n689)
  );
  //AND U272bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U272bar (
    .O(n698bar),
    .I0(n690bar),
    .I1(n689bar)
  );
  //OR U273
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U273 (
    .O(n689),
    .I0(n688),
    .I1(n687)
  );
  //AND U273bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U273bar (
    .O(n689bar),
    .I0(n688bar),
    .I1(n687bar)
  );
  //OR U274
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U274 (
    .O(n687),
    .I0(in[90]),
    .I1(in[254])
  );
  //AND U274bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U274bar (
    .O(n687bar),
    .I0(inbar[90]),
    .I1(inbar[254])
  );
  //OR U275
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U275 (
    .O(n688),
    .I0(in_36),
    .I1(in_32)
  );
  //AND U275bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U275bar (
    .O(n688bar),
    .I0(in_36bar),
    .I1(in_32bar)
  );
  //OR U276
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U276 (
    .O(n690),
    .I0(n686),
    .I1(n685)
  );
  //AND U276bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U276bar (
    .O(n690bar),
    .I0(n686bar),
    .I1(n685bar)
  );
  //OR U277
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U277 (
    .O(n685),
    .I0(in_62),
    .I1(in_37)
  );
  //AND U277bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U277bar (
    .O(n685bar),
    .I0(in_62bar),
    .I1(in_37bar)
  );
  //OR U278
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U278 (
    .O(n686),
    .I0(in_75),
    .I1(in_73)
  );
  //AND U278bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U278bar (
    .O(n686bar),
    .I0(in_75bar),
    .I1(in_73bar)
  );
  //OR U279
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U279 (
    .O(n944),
    .I0(n684),
    .I1(n683)
  );
  //AND U279bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U279bar (
    .O(n944bar),
    .I0(n684bar),
    .I1(n683bar)
  );
  //OR U280
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U280 (
    .O(n683),
    .I0(n682),
    .I1(n681)
  );
  //AND U280bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U280bar (
    .O(n683bar),
    .I0(n682bar),
    .I1(n681bar)
  );
  //OR U281
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U281 (
    .O(n681),
    .I0(n680),
    .I1(n679)
  );
  //AND U281bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U281bar (
    .O(n681bar),
    .I0(n680bar),
    .I1(n679bar)
  );
  //OR U282
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U282 (
    .O(n679),
    .I0(in[171]),
    .I1(in[153])
  );
  //AND U282bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U282bar (
    .O(n679bar),
    .I0(inbar[171]),
    .I1(inbar[153])
  );
  //OR U283
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U283 (
    .O(n680),
    .I0(in[187]),
    .I1(in[176])
  );
  //AND U283bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U283bar (
    .O(n680bar),
    .I0(inbar[187]),
    .I1(inbar[176])
  );
  //OR U284
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U284 (
    .O(n682),
    .I0(n678),
    .I1(n677)
  );
  //AND U284bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U284bar (
    .O(n682bar),
    .I0(n678bar),
    .I1(n677bar)
  );
  //OR U285
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U285 (
    .O(n677),
    .I0(in[245]),
    .I1(in[211])
  );
  //AND U285bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U285bar (
    .O(n677bar),
    .I0(inbar[245]),
    .I1(inbar[211])
  );
  //OR U286
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U286 (
    .O(n678),
    .I0(in[97]),
    .I1(in[88])
  );
  //AND U286bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U286bar (
    .O(n678bar),
    .I0(inbar[97]),
    .I1(inbar[88])
  );
  //OR U287
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U287 (
    .O(n684),
    .I0(n676),
    .I1(n675)
  );
  //AND U287bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U287bar (
    .O(n684bar),
    .I0(n676bar),
    .I1(n675bar)
  );
  //OR U288
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U288 (
    .O(n675),
    .I0(n674),
    .I1(n673)
  );
  //AND U288bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U288bar (
    .O(n675bar),
    .I0(n674bar),
    .I1(n673bar)
  );
  //OR U289
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U289 (
    .O(n673),
    .I0(in_10),
    .I1(in_0)
  );
  //AND U289bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U289bar (
    .O(n673bar),
    .I0(in_10bar),
    .I1(in_0bar)
  );
  //OR U290
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U290 (
    .O(n674),
    .I0(in_59),
    .I1(in_5)
  );
  //AND U290bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U290bar (
    .O(n674bar),
    .I0(in_59bar),
    .I1(in_5bar)
  );
  //OR U291
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U291 (
    .O(n676),
    .I0(n672),
    .I1(n671)
  );
  //AND U291bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U291bar (
    .O(n676bar),
    .I0(n672bar),
    .I1(n671bar)
  );
  //OR U292
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U292 (
    .O(n671),
    .I0(in_60),
    .I1(in_6)
  );
  //AND U292bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U292bar (
    .O(n671bar),
    .I0(in_60bar),
    .I1(in_6bar)
  );
  //OR U293
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U293 (
    .O(n672),
    .I0(in_77),
    .I1(in_69)
  );
  //AND U293bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U293bar (
    .O(n672bar),
    .I0(in_77bar),
    .I1(in_69bar)
  );
  //OR U294
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U294 (
    .O(n700),
    .I0(in[113]),
    .I1(n864)
  );
  //AND U294bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U294bar (
    .O(n700bar),
    .I0(inbar[113]),
    .I1(n864bar)
  );
  //OR U295
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U295 (
    .O(n864),
    .I0(n670),
    .I1(n669)
  );
  //AND U295bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U295bar (
    .O(n864bar),
    .I0(n670bar),
    .I1(n669bar)
  );
  //OR U296
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U296 (
    .O(n669),
    .I0(n668),
    .I1(n667)
  );
  //AND U296bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U296bar (
    .O(n669bar),
    .I0(n668bar),
    .I1(n667bar)
  );
  //OR U297
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U297 (
    .O(n667),
    .I0(n666),
    .I1(n665)
  );
  //AND U297bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U297bar (
    .O(n667bar),
    .I0(n666bar),
    .I1(n665bar)
  );
  //OR U298
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U298 (
    .O(n665),
    .I0(in[125]),
    .I1(in[107])
  );
  //AND U298bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U298bar (
    .O(n665bar),
    .I0(inbar[125]),
    .I1(inbar[107])
  );
  //OR U299
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U299 (
    .O(n666),
    .I0(in[138]),
    .I1(in[126])
  );
  //AND U299bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U299bar (
    .O(n666bar),
    .I0(inbar[138]),
    .I1(inbar[126])
  );
  //OR U300
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U300 (
    .O(n668),
    .I0(n664),
    .I1(n663)
  );
  //AND U300bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U300bar (
    .O(n668bar),
    .I0(n664bar),
    .I1(n663bar)
  );
  //OR U301
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U301 (
    .O(n663),
    .I0(in[189]),
    .I1(in[143])
  );
  //AND U301bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U301bar (
    .O(n663bar),
    .I0(inbar[189]),
    .I1(inbar[143])
  );
  //OR U302
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U302 (
    .O(n664),
    .I0(in[99]),
    .I1(in[214])
  );
  //AND U302bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U302bar (
    .O(n664bar),
    .I0(inbar[99]),
    .I1(inbar[214])
  );
  //OR U303
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U303 (
    .O(n670),
    .I0(n662),
    .I1(n661)
  );
  //AND U303bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U303bar (
    .O(n670bar),
    .I0(n662bar),
    .I1(n661bar)
  );
  //OR U304
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U304 (
    .O(n661),
    .I0(n660),
    .I1(n659)
  );
  //AND U304bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U304bar (
    .O(n661bar),
    .I0(n660bar),
    .I1(n659bar)
  );
  //OR U305
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U305 (
    .O(n659),
    .I0(in_15),
    .I1(in_12)
  );
  //AND U305bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U305bar (
    .O(n659bar),
    .I0(in_15bar),
    .I1(in_12bar)
  );
  //OR U306
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U306 (
    .O(n660),
    .I0(in_20),
    .I1(in_2)
  );
  //AND U306bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U306bar (
    .O(n660bar),
    .I0(in_20bar),
    .I1(in_2bar)
  );
  //OR U307
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U307 (
    .O(n662),
    .I0(n658),
    .I1(n657)
  );
  //AND U307bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U307bar (
    .O(n662bar),
    .I0(n658bar),
    .I1(n657bar)
  );
  //OR U308
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U308 (
    .O(n657),
    .I0(in_30),
    .I1(in_3)
  );
  //AND U308bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U308bar (
    .O(n657bar),
    .I0(in_30bar),
    .I1(in_3bar)
  );
  //OR U309
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U309 (
    .O(n658),
    .I0(in_4),
    .I1(in_38)
  );
  //AND U309bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U309bar (
    .O(n658bar),
    .I0(in_4bar),
    .I1(in_38bar)
  );
  //OR U310
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U310 (
    .O(n702),
    .I0(n656),
    .I1(n655)
  );
  //AND U310bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U310bar (
    .O(n702bar),
    .I0(n656bar),
    .I1(n655bar)
  );
  //OR U311
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U311 (
    .O(n655),
    .I0(in[148]),
    .I1(in[137])
  );
  //AND U311bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U311bar (
    .O(n655bar),
    .I0(inbar[148]),
    .I1(inbar[137])
  );
  //OR U312
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U312 (
    .O(n656),
    .I0(in[149]),
    .I1(n654)
  );
  //AND U312bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U312bar (
    .O(n656bar),
    .I0(inbar[149]),
    .I1(n654bar)
  );
  //OR U313
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U313 (
    .O(n654),
    .I0(in[195]),
    .I1(in[190])
  );
  //AND U313bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U313bar (
    .O(n654bar),
    .I0(inbar[195]),
    .I1(inbar[190])
  );
  //OR U314
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U314 (
    .O(n704),
    .I0(n653),
    .I1(n652)
  );
  //AND U314bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U314bar (
    .O(n704bar),
    .I0(n653bar),
    .I1(n652bar)
  );
  //OR U315
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U315 (
    .O(n652),
    .I0(n651),
    .I1(n650)
  );
  //AND U315bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U315bar (
    .O(n652bar),
    .I0(n651bar),
    .I1(n650bar)
  );
  //OR U316
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U316 (
    .O(n650),
    .I0(in[98]),
    .I1(in[197])
  );
  //AND U316bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U316bar (
    .O(n650bar),
    .I0(inbar[98]),
    .I1(inbar[197])
  );
  //OR U317
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U317 (
    .O(n651),
    .I0(in_11),
    .I1(n649)
  );
  //AND U317bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U317bar (
    .O(n651bar),
    .I0(in_11bar),
    .I1(n649bar)
  );
  //OR U318
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U318 (
    .O(n649),
    .I0(in_26),
    .I1(in_14)
  );
  //AND U318bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U318bar (
    .O(n649bar),
    .I0(in_26bar),
    .I1(in_14bar)
  );
  //OR U319
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U319 (
    .O(n653),
    .I0(n648),
    .I1(n647)
  );
  //AND U319bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U319bar (
    .O(n653bar),
    .I0(n648bar),
    .I1(n647bar)
  );
  //OR U320
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U320 (
    .O(n647),
    .I0(in_35),
    .I1(in_27)
  );
  //AND U320bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U320bar (
    .O(n647bar),
    .I0(in_35bar),
    .I1(in_27bar)
  );
  //OR U321
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U321 (
    .O(n648),
    .I0(in_50),
    .I1(n646)
  );
  //AND U321bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U321bar (
    .O(n648bar),
    .I0(in_50bar),
    .I1(n646bar)
  );
  //OR U322
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U322 (
    .O(n646),
    .I0(in_78),
    .I1(in_61)
  );
  //AND U322bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U322bar (
    .O(n646bar),
    .I0(in_78bar),
    .I1(in_61bar)
  );
  //OR U323
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U323 (
    .O(n720),
    .I0(n942),
    .I1(n645)
  );
  //AND U323bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U323bar (
    .O(n720bar),
    .I0(n942bar),
    .I1(n645bar)
  );
  //OR U324
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U324 (
    .O(n645),
    .I0(in[106]),
    .I1(n863)
  );
  //AND U324bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U324bar (
    .O(n645bar),
    .I0(inbar[106]),
    .I1(n863bar)
  );
  //OR U325
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U325 (
    .O(n863),
    .I0(n644),
    .I1(n643)
  );
  //AND U325bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U325bar (
    .O(n863bar),
    .I0(n644bar),
    .I1(n643bar)
  );
  //OR U326
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U326 (
    .O(n643),
    .I0(n642),
    .I1(n641)
  );
  //AND U326bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U326bar (
    .O(n643bar),
    .I0(n642bar),
    .I1(n641bar)
  );
  //OR U327
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U327 (
    .O(n641),
    .I0(n640),
    .I1(n639)
  );
  //AND U327bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U327bar (
    .O(n641bar),
    .I0(n640bar),
    .I1(n639bar)
  );
  //OR U328
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U328 (
    .O(n639),
    .I0(in[127]),
    .I1(in[122])
  );
  //AND U328bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U328bar (
    .O(n639bar),
    .I0(inbar[127]),
    .I1(inbar[122])
  );
  //OR U329
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U329 (
    .O(n640),
    .I0(in[156]),
    .I1(in[132])
  );
  //AND U329bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U329bar (
    .O(n640bar),
    .I0(inbar[156]),
    .I1(inbar[132])
  );
  //OR U330
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U330 (
    .O(n642),
    .I0(n638),
    .I1(n637)
  );
  //AND U330bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U330bar (
    .O(n642bar),
    .I0(n638bar),
    .I1(n637bar)
  );
  //OR U331
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U331 (
    .O(n637),
    .I0(in[159]),
    .I1(in[157])
  );
  //AND U331bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U331bar (
    .O(n637bar),
    .I0(inbar[159]),
    .I1(inbar[157])
  );
  //OR U332
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U332 (
    .O(n638),
    .I0(in[185]),
    .I1(in[169])
  );
  //AND U332bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U332bar (
    .O(n638bar),
    .I0(inbar[185]),
    .I1(inbar[169])
  );
  //OR U333
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U333 (
    .O(n644),
    .I0(n636),
    .I1(n635)
  );
  //AND U333bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U333bar (
    .O(n644bar),
    .I0(n636bar),
    .I1(n635bar)
  );
  //OR U334
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U334 (
    .O(n635),
    .I0(n634),
    .I1(n633)
  );
  //AND U334bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U334bar (
    .O(n635bar),
    .I0(n634bar),
    .I1(n633bar)
  );
  //OR U335
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U335 (
    .O(n633),
    .I0(in[239]),
    .I1(in[218])
  );
  //AND U335bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U335bar (
    .O(n633bar),
    .I0(inbar[239]),
    .I1(inbar[218])
  );
  //OR U336
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U336 (
    .O(n634),
    .I0(in_13),
    .I1(in[87])
  );
  //AND U336bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U336bar (
    .O(n634bar),
    .I0(in_13bar),
    .I1(inbar[87])
  );
  //OR U337
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U337 (
    .O(n636),
    .I0(n632),
    .I1(n631)
  );
  //AND U337bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U337bar (
    .O(n636bar),
    .I0(n632bar),
    .I1(n631bar)
  );
  //OR U338
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U338 (
    .O(n631),
    .I0(in_72),
    .I1(in_70)
  );
  //AND U338bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U338bar (
    .O(n631bar),
    .I0(in_72bar),
    .I1(in_70bar)
  );
  //OR U339
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U339 (
    .O(n632),
    .I0(in_80),
    .I1(in_74)
  );
  //AND U339bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U339bar (
    .O(n632bar),
    .I0(in_80bar),
    .I1(in_74bar)
  );
  //OR U340
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U340 (
    .O(n942),
    .I0(n630),
    .I1(n629)
  );
  //AND U340bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U340bar (
    .O(n942bar),
    .I0(n630bar),
    .I1(n629bar)
  );
  //OR U341
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U341 (
    .O(n629),
    .I0(n628),
    .I1(n627)
  );
  //AND U341bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U341bar (
    .O(n629bar),
    .I0(n628bar),
    .I1(n627bar)
  );
  //OR U342
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U342 (
    .O(n627),
    .I0(n626),
    .I1(n625)
  );
  //AND U342bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U342bar (
    .O(n627bar),
    .I0(n626bar),
    .I1(n625bar)
  );
  //OR U343
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U343 (
    .O(n625),
    .I0(in[146]),
    .I1(in[100])
  );
  //AND U343bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U343bar (
    .O(n625bar),
    .I0(inbar[146]),
    .I1(inbar[100])
  );
  //OR U344
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U344 (
    .O(n626),
    .I0(in[168]),
    .I1(in[152])
  );
  //AND U344bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U344bar (
    .O(n626bar),
    .I0(inbar[168]),
    .I1(inbar[152])
  );
  //OR U345
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U345 (
    .O(n628),
    .I0(n624),
    .I1(n623)
  );
  //AND U345bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U345bar (
    .O(n628bar),
    .I0(n624bar),
    .I1(n623bar)
  );
  //OR U346
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U346 (
    .O(n623),
    .I0(in[199]),
    .I1(in[182])
  );
  //AND U346bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U346bar (
    .O(n623bar),
    .I0(inbar[199]),
    .I1(inbar[182])
  );
  //OR U347
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U347 (
    .O(n624),
    .I0(in[236]),
    .I1(in[204])
  );
  //AND U347bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U347bar (
    .O(n624bar),
    .I0(inbar[236]),
    .I1(inbar[204])
  );
  //OR U348
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U348 (
    .O(n630),
    .I0(n622),
    .I1(n621)
  );
  //AND U348bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U348bar (
    .O(n630bar),
    .I0(n622bar),
    .I1(n621bar)
  );
  //OR U349
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U349 (
    .O(n621),
    .I0(n620),
    .I1(n619)
  );
  //AND U349bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U349bar (
    .O(n621bar),
    .I0(n620bar),
    .I1(n619bar)
  );
  //OR U350
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U350 (
    .O(n619),
    .I0(in[89]),
    .I1(in[246])
  );
  //AND U350bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U350bar (
    .O(n619bar),
    .I0(inbar[89]),
    .I1(inbar[246])
  );
  //OR U351
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U351 (
    .O(n620),
    .I0(in[95]),
    .I1(in[92])
  );
  //AND U351bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U351bar (
    .O(n620bar),
    .I0(inbar[95]),
    .I1(inbar[92])
  );
  //OR U352
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U352 (
    .O(n622),
    .I0(n618),
    .I1(n617)
  );
  //AND U352bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U352bar (
    .O(n622bar),
    .I0(n618bar),
    .I1(n617bar)
  );
  //OR U353
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U353 (
    .O(n617),
    .I0(in_22),
    .I1(in_16)
  );
  //AND U353bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U353bar (
    .O(n617bar),
    .I0(in_22bar),
    .I1(in_16bar)
  );
  //OR U354
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U354 (
    .O(n618),
    .I0(in_51),
    .I1(in_49)
  );
  //AND U354bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U354bar (
    .O(n618bar),
    .I0(in_51bar),
    .I1(in_49bar)
  );
  //OR U355
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U355 (
    .O(n722),
    .I0(n616),
    .I1(n615)
  );
  //AND U355bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U355bar (
    .O(n722bar),
    .I0(n616bar),
    .I1(n615bar)
  );
  //OR U356
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U356 (
    .O(n615),
    .I0(in[158]),
    .I1(in[115])
  );
  //AND U356bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U356bar (
    .O(n615bar),
    .I0(inbar[158]),
    .I1(inbar[115])
  );
  //OR U357
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U357 (
    .O(n616),
    .I0(in[163]),
    .I1(n614)
  );
  //AND U357bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U357bar (
    .O(n616bar),
    .I0(inbar[163]),
    .I1(n614bar)
  );
  //OR U358
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U358 (
    .O(n614),
    .I0(in[206]),
    .I1(in[165])
  );
  //AND U358bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U358bar (
    .O(n614bar),
    .I0(inbar[206]),
    .I1(inbar[165])
  );
  //OR U359
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U359 (
    .O(n724),
    .I0(n613),
    .I1(n612)
  );
  //AND U359bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U359bar (
    .O(n724bar),
    .I0(n613bar),
    .I1(n612bar)
  );
  //OR U360
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U360 (
    .O(n612),
    .I0(n611),
    .I1(n610)
  );
  //AND U360bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U360bar (
    .O(n612bar),
    .I0(n611bar),
    .I1(n610bar)
  );
  //OR U361
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U361 (
    .O(n610),
    .I0(in[213]),
    .I1(in[207])
  );
  //AND U361bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U361bar (
    .O(n610bar),
    .I0(inbar[213]),
    .I1(inbar[207])
  );
  //OR U362
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U362 (
    .O(n611),
    .I0(in[215]),
    .I1(n609)
  );
  //AND U362bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U362bar (
    .O(n611bar),
    .I0(inbar[215]),
    .I1(n609bar)
  );
  //OR U363
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U363 (
    .O(n609),
    .I0(in[230]),
    .I1(in[220])
  );
  //AND U363bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U363bar (
    .O(n609bar),
    .I0(inbar[230]),
    .I1(inbar[220])
  );
  //OR U364
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U364 (
    .O(n613),
    .I0(n608),
    .I1(n607)
  );
  //AND U364bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U364bar (
    .O(n613bar),
    .I0(n608bar),
    .I1(n607bar)
  );
  //OR U365
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U365 (
    .O(n607),
    .I0(in[251]),
    .I1(in[234])
  );
  //AND U365bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U365bar (
    .O(n607bar),
    .I0(inbar[251]),
    .I1(inbar[234])
  );
  //OR U366
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U366 (
    .O(n608),
    .I0(in_17),
    .I1(n606)
  );
  //AND U366bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U366bar (
    .O(n608bar),
    .I0(in_17bar),
    .I1(n606bar)
  );
  //OR U367
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U367 (
    .O(n606),
    .I0(in_65),
    .I1(in_56)
  );
  //AND U367bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U367bar (
    .O(n606bar),
    .I0(in_65bar),
    .I1(in_56bar)
  );
  //OR U368
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U368 (
    .O(out[0]),
    .I0(n605),
    .I1(n604)
  );
  //AND U368bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U368bar (
    .O(outbar[0]),
    .I0(n605bar),
    .I1(n604bar)
  );
  //OR U369
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U369 (
    .O(n604),
    .I0(n603),
    .I1(n602)
  );
  //AND U369bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U369bar (
    .O(n604bar),
    .I0(n603bar),
    .I1(n602bar)
  );
  //OR U370
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U370 (
    .O(n602),
    .I0(n601),
    .I1(n600)
  );
  //AND U370bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U370bar (
    .O(n602bar),
    .I0(n601bar),
    .I1(n600bar)
  );
  //OR U371
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U371 (
    .O(n600),
    .I0(n820),
    .I1(n785)
  );
  //AND U371bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U371bar (
    .O(n600bar),
    .I0(n820bar),
    .I1(n785bar)
  );
  //OR U372
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U372 (
    .O(n785),
    .I0(n599),
    .I1(n598)
  );
  //AND U372bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U372bar (
    .O(n785bar),
    .I0(n599bar),
    .I1(n598bar)
  );
  //OR U373
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U373 (
    .O(n598),
    .I0(n597),
    .I1(n596)
  );
  //AND U373bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U373bar (
    .O(n598bar),
    .I0(n597bar),
    .I1(n596bar)
  );
  //OR U374
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U374 (
    .O(n596),
    .I0(n595),
    .I1(n594)
  );
  //AND U374bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U374bar (
    .O(n596bar),
    .I0(n595bar),
    .I1(n594bar)
  );
  //OR U375
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U375 (
    .O(n594),
    .I0(in[135]),
    .I1(in[104])
  );
  //AND U375bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U375bar (
    .O(n594bar),
    .I0(inbar[135]),
    .I1(inbar[104])
  );
  //OR U376
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U376 (
    .O(n595),
    .I0(in[188]),
    .I1(in[178])
  );
  //AND U376bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U376bar (
    .O(n595bar),
    .I0(inbar[188]),
    .I1(inbar[178])
  );
  //OR U377
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U377 (
    .O(n597),
    .I0(n593),
    .I1(n592)
  );
  //AND U377bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U377bar (
    .O(n597bar),
    .I0(n593bar),
    .I1(n592bar)
  );
  //OR U378
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U378 (
    .O(n592),
    .I0(in[217]),
    .I1(in[194])
  );
  //AND U378bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U378bar (
    .O(n592bar),
    .I0(inbar[217]),
    .I1(inbar[194])
  );
  //OR U379
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U379 (
    .O(n593),
    .I0(in[237]),
    .I1(in[218])
  );
  //AND U379bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U379bar (
    .O(n593bar),
    .I0(inbar[237]),
    .I1(inbar[218])
  );
  //OR U380
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U380 (
    .O(n599),
    .I0(n591),
    .I1(n590)
  );
  //AND U380bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U380bar (
    .O(n599bar),
    .I0(n591bar),
    .I1(n590bar)
  );
  //OR U381
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U381 (
    .O(n590),
    .I0(n589),
    .I1(n588)
  );
  //AND U381bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U381bar (
    .O(n590bar),
    .I0(n589bar),
    .I1(n588bar)
  );
  //OR U382
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U382 (
    .O(n588),
    .I0(in_2),
    .I1(in_10)
  );
  //AND U382bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U382bar (
    .O(n588bar),
    .I0(in_2bar),
    .I1(in_10bar)
  );
  //OR U383
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U383 (
    .O(n589),
    .I0(in_47),
    .I1(in_22)
  );
  //AND U383bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U383bar (
    .O(n589bar),
    .I0(in_47bar),
    .I1(in_22bar)
  );
  //OR U384
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U384 (
    .O(n591),
    .I0(n587),
    .I1(n586)
  );
  //AND U384bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U384bar (
    .O(n591bar),
    .I0(n587bar),
    .I1(n586bar)
  );
  //OR U385
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U385 (
    .O(n586),
    .I0(in_56),
    .I1(in_54)
  );
  //AND U385bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U385bar (
    .O(n586bar),
    .I0(in_56bar),
    .I1(in_54bar)
  );
  //OR U386
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U386 (
    .O(n587),
    .I0(in_63),
    .I1(in_61)
  );
  //AND U386bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U386bar (
    .O(n587bar),
    .I0(in_63bar),
    .I1(in_61bar)
  );
  //OR U387
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U387 (
    .O(n820),
    .I0(n585),
    .I1(n584)
  );
  //AND U387bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U387bar (
    .O(n820bar),
    .I0(n585bar),
    .I1(n584bar)
  );
  //OR U388
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U388 (
    .O(n584),
    .I0(n583),
    .I1(n582)
  );
  //AND U388bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U388bar (
    .O(n584bar),
    .I0(n583bar),
    .I1(n582bar)
  );
  //OR U389
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U389 (
    .O(n582),
    .I0(n581),
    .I1(n580)
  );
  //AND U389bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U389bar (
    .O(n582bar),
    .I0(n581bar),
    .I1(n580bar)
  );
  //OR U390
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U390 (
    .O(n580),
    .I0(in[158]),
    .I1(in[142])
  );
  //AND U390bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U390bar (
    .O(n580bar),
    .I0(inbar[158]),
    .I1(inbar[142])
  );
  //OR U391
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U391 (
    .O(n581),
    .I0(in[175]),
    .I1(in[164])
  );
  //AND U391bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U391bar (
    .O(n581bar),
    .I0(inbar[175]),
    .I1(inbar[164])
  );
  //OR U392
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U392 (
    .O(n583),
    .I0(n579),
    .I1(n578)
  );
  //AND U392bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U392bar (
    .O(n583bar),
    .I0(n579bar),
    .I1(n578bar)
  );
  //OR U393
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U393 (
    .O(n578),
    .I0(in[228]),
    .I1(in[204])
  );
  //AND U393bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U393bar (
    .O(n578bar),
    .I0(inbar[228]),
    .I1(inbar[204])
  );
  //OR U394
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U394 (
    .O(n579),
    .I0(in[91]),
    .I1(in[87])
  );
  //AND U394bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U394bar (
    .O(n579bar),
    .I0(inbar[91]),
    .I1(inbar[87])
  );
  //OR U395
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U395 (
    .O(n585),
    .I0(n577),
    .I1(n576)
  );
  //AND U395bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U395bar (
    .O(n585bar),
    .I0(n577bar),
    .I1(n576bar)
  );
  //OR U396
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U396 (
    .O(n576),
    .I0(n575),
    .I1(n574)
  );
  //AND U396bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U396bar (
    .O(n576bar),
    .I0(n575bar),
    .I1(n574bar)
  );
  //OR U397
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U397 (
    .O(n574),
    .I0(in_21),
    .I1(in_11)
  );
  //AND U397bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U397bar (
    .O(n574bar),
    .I0(in_21bar),
    .I1(in_11bar)
  );
  //OR U398
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U398 (
    .O(n575),
    .I0(in_5),
    .I1(in_3)
  );
  //AND U398bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U398bar (
    .O(n575bar),
    .I0(in_5bar),
    .I1(in_3bar)
  );
  //OR U399
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U399 (
    .O(n577),
    .I0(n573),
    .I1(n572)
  );
  //AND U399bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U399bar (
    .O(n577bar),
    .I0(n573bar),
    .I1(n572bar)
  );
  //OR U400
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U400 (
    .O(n572),
    .I0(in_68),
    .I1(in_64)
  );
  //AND U400bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U400bar (
    .O(n572bar),
    .I0(in_68bar),
    .I1(in_64bar)
  );
  //OR U401
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U401 (
    .O(n573),
    .I0(in_76),
    .I1(in_73)
  );
  //AND U401bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U401bar (
    .O(n573bar),
    .I0(in_76bar),
    .I1(in_73bar)
  );
  //OR U402
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U402 (
    .O(n601),
    .I0(n778),
    .I1(n571)
  );
  //AND U402bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U402bar (
    .O(n601bar),
    .I0(n778bar),
    .I1(n571bar)
  );
  //OR U403
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U403 (
    .O(n571),
    .I0(in[100]),
    .I1(n965)
  );
  //AND U403bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U403bar (
    .O(n571bar),
    .I0(inbar[100]),
    .I1(n965bar)
  );
  //OR U404
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U404 (
    .O(n965),
    .I0(n570),
    .I1(n569)
  );
  //AND U404bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U404bar (
    .O(n965bar),
    .I0(n570bar),
    .I1(n569bar)
  );
  //OR U405
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U405 (
    .O(n569),
    .I0(n568),
    .I1(n567)
  );
  //AND U405bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U405bar (
    .O(n569bar),
    .I0(n568bar),
    .I1(n567bar)
  );
  //OR U406
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U406 (
    .O(n567),
    .I0(n566),
    .I1(n565)
  );
  //AND U406bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U406bar (
    .O(n567bar),
    .I0(n566bar),
    .I1(n565bar)
  );
  //OR U407
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U407 (
    .O(n565),
    .I0(n817),
    .I1(n750)
  );
  //AND U407bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U407bar (
    .O(n565bar),
    .I0(n817bar),
    .I1(n750bar)
  );
  //OR U408
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U408 (
    .O(n750),
    .I0(n564),
    .I1(n563)
  );
  //AND U408bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U408bar (
    .O(n750bar),
    .I0(n564bar),
    .I1(n563bar)
  );
  //OR U409
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U409 (
    .O(n563),
    .I0(n562),
    .I1(n561)
  );
  //AND U409bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U409bar (
    .O(n563bar),
    .I0(n562bar),
    .I1(n561bar)
  );
  //OR U410
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U410 (
    .O(n561),
    .I0(n560),
    .I1(n559)
  );
  //AND U410bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U410bar (
    .O(n561bar),
    .I0(n560bar),
    .I1(n559bar)
  );
  //OR U411
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U411 (
    .O(n559),
    .I0(in[119]),
    .I1(in[103])
  );
  //AND U411bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U411bar (
    .O(n559bar),
    .I0(inbar[119]),
    .I1(inbar[103])
  );
  //OR U412
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U412 (
    .O(n560),
    .I0(in[137]),
    .I1(in[133])
  );
  //AND U412bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U412bar (
    .O(n560bar),
    .I0(inbar[137]),
    .I1(inbar[133])
  );
  //OR U413
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U413 (
    .O(n562),
    .I0(n558),
    .I1(n557)
  );
  //AND U413bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U413bar (
    .O(n562bar),
    .I0(n558bar),
    .I1(n557bar)
  );
  //OR U414
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U414 (
    .O(n557),
    .I0(in[176]),
    .I1(in[173])
  );
  //AND U414bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U414bar (
    .O(n557bar),
    .I0(inbar[176]),
    .I1(inbar[173])
  );
  //OR U415
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U415 (
    .O(n558),
    .I0(in[210]),
    .I1(in[181])
  );
  //AND U415bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U415bar (
    .O(n558bar),
    .I0(inbar[210]),
    .I1(inbar[181])
  );
  //OR U416
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U416 (
    .O(n564),
    .I0(n556),
    .I1(n555)
  );
  //AND U416bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U416bar (
    .O(n564bar),
    .I0(n556bar),
    .I1(n555bar)
  );
  //OR U417
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U417 (
    .O(n555),
    .I0(n554),
    .I1(n553)
  );
  //AND U417bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U417bar (
    .O(n555bar),
    .I0(n554bar),
    .I1(n553bar)
  );
  //OR U418
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U418 (
    .O(n553),
    .I0(in_13),
    .I1(in[234])
  );
  //AND U418bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U418bar (
    .O(n553bar),
    .I0(in_13bar),
    .I1(inbar[234])
  );
  //OR U419
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U419 (
    .O(n554),
    .I0(in_38),
    .I1(in_32)
  );
  //AND U419bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U419bar (
    .O(n554bar),
    .I0(in_38bar),
    .I1(in_32bar)
  );
  //OR U420
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U420 (
    .O(n556),
    .I0(n552),
    .I1(n551)
  );
  //AND U420bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U420bar (
    .O(n556bar),
    .I0(n552bar),
    .I1(n551bar)
  );
  //OR U421
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U421 (
    .O(n551),
    .I0(in_42),
    .I1(in_41)
  );
  //AND U421bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U421bar (
    .O(n551bar),
    .I0(in_42bar),
    .I1(in_41bar)
  );
  //OR U422
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U422 (
    .O(n552),
    .I0(in_7),
    .I1(in_49)
  );
  //AND U422bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U422bar (
    .O(n552bar),
    .I0(in_7bar),
    .I1(in_49bar)
  );
  //OR U423
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U423 (
    .O(n817),
    .I0(n550),
    .I1(n549)
  );
  //AND U423bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U423bar (
    .O(n817bar),
    .I0(n550bar),
    .I1(n549bar)
  );
  //OR U424
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U424 (
    .O(n549),
    .I0(n548),
    .I1(n547)
  );
  //AND U424bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U424bar (
    .O(n549bar),
    .I0(n548bar),
    .I1(n547bar)
  );
  //OR U425
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U425 (
    .O(n547),
    .I0(n546),
    .I1(n545)
  );
  //AND U425bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U425bar (
    .O(n547bar),
    .I0(n546bar),
    .I1(n545bar)
  );
  //OR U426
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U426 (
    .O(n545),
    .I0(in[159]),
    .I1(in[105])
  );
  //AND U426bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U426bar (
    .O(n545bar),
    .I0(inbar[159]),
    .I1(inbar[105])
  );
  //OR U427
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U427 (
    .O(n546),
    .I0(in[206]),
    .I1(in[183])
  );
  //AND U427bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U427bar (
    .O(n546bar),
    .I0(inbar[206]),
    .I1(inbar[183])
  );
  //OR U428
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U428 (
    .O(n548),
    .I0(n544),
    .I1(n543)
  );
  //AND U428bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U428bar (
    .O(n548bar),
    .I0(n544bar),
    .I1(n543bar)
  );
  //OR U429
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U429 (
    .O(n543),
    .I0(in[229]),
    .I1(in[219])
  );
  //AND U429bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U429bar (
    .O(n543bar),
    .I0(inbar[229]),
    .I1(inbar[219])
  );
  //OR U430
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U430 (
    .O(n544),
    .I0(in[235]),
    .I1(in[232])
  );
  //AND U430bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U430bar (
    .O(n544bar),
    .I0(inbar[235]),
    .I1(inbar[232])
  );
  //OR U431
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U431 (
    .O(n550),
    .I0(n542),
    .I1(n541)
  );
  //AND U431bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U431bar (
    .O(n550bar),
    .I0(n542bar),
    .I1(n541bar)
  );
  //OR U432
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U432 (
    .O(n541),
    .I0(n540),
    .I1(n539)
  );
  //AND U432bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U432bar (
    .O(n541bar),
    .I0(n540bar),
    .I1(n539bar)
  );
  //OR U433
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U433 (
    .O(n539),
    .I0(in[249]),
    .I1(in[242])
  );
  //AND U433bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U433bar (
    .O(n539bar),
    .I0(inbar[249]),
    .I1(inbar[242])
  );
  //OR U434
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U434 (
    .O(n540),
    .I0(in[89]),
    .I1(in[254])
  );
  //AND U434bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U434bar (
    .O(n540bar),
    .I0(inbar[89]),
    .I1(inbar[254])
  );
  //OR U435
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U435 (
    .O(n542),
    .I0(n538),
    .I1(n537)
  );
  //AND U435bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U435bar (
    .O(n542bar),
    .I0(n538bar),
    .I1(n537bar)
  );
  //OR U436
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U436 (
    .O(n537),
    .I0(in_14),
    .I1(in[99])
  );
  //AND U436bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U436bar (
    .O(n537bar),
    .I0(in_14bar),
    .I1(inbar[99])
  );
  //OR U437
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U437 (
    .O(n538),
    .I0(in_60),
    .I1(in_18)
  );
  //AND U437bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U437bar (
    .O(n538bar),
    .I0(in_60bar),
    .I1(in_18bar)
  );
  //OR U438
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U438 (
    .O(n566),
    .I0(in[113]),
    .I1(n763)
  );
  //AND U438bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U438bar (
    .O(n566bar),
    .I0(inbar[113]),
    .I1(n763bar)
  );
  //OR U439
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U439 (
    .O(n763),
    .I0(n536),
    .I1(n535)
  );
  //AND U439bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U439bar (
    .O(n763bar),
    .I0(n536bar),
    .I1(n535bar)
  );
  //OR U440
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U440 (
    .O(n535),
    .I0(n534),
    .I1(n533)
  );
  //AND U440bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U440bar (
    .O(n535bar),
    .I0(n534bar),
    .I1(n533bar)
  );
  //OR U441
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U441 (
    .O(n533),
    .I0(n532),
    .I1(n531)
  );
  //AND U441bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U441bar (
    .O(n533bar),
    .I0(n532bar),
    .I1(n531bar)
  );
  //OR U442
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U442 (
    .O(n531),
    .I0(in[115]),
    .I1(in[110])
  );
  //AND U442bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U442bar (
    .O(n531bar),
    .I0(inbar[115]),
    .I1(inbar[110])
  );
  //OR U443
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U443 (
    .O(n532),
    .I0(in[125]),
    .I1(in[117])
  );
  //AND U443bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U443bar (
    .O(n532bar),
    .I0(inbar[125]),
    .I1(inbar[117])
  );
  //OR U444
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U444 (
    .O(n534),
    .I0(n530),
    .I1(n529)
  );
  //AND U444bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U444bar (
    .O(n534bar),
    .I0(n530bar),
    .I1(n529bar)
  );
  //OR U445
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U445 (
    .O(n529),
    .I0(in[180]),
    .I1(in[128])
  );
  //AND U445bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U445bar (
    .O(n529bar),
    .I0(inbar[180]),
    .I1(inbar[128])
  );
  //OR U446
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U446 (
    .O(n530),
    .I0(in[205]),
    .I1(in[201])
  );
  //AND U446bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U446bar (
    .O(n530bar),
    .I0(inbar[205]),
    .I1(inbar[201])
  );
  //OR U447
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U447 (
    .O(n536),
    .I0(n528),
    .I1(n527)
  );
  //AND U447bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U447bar (
    .O(n536bar),
    .I0(n528bar),
    .I1(n527bar)
  );
  //OR U448
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U448 (
    .O(n527),
    .I0(n526),
    .I1(n525)
  );
  //AND U448bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U448bar (
    .O(n527bar),
    .I0(n526bar),
    .I1(n525bar)
  );
  //OR U449
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U449 (
    .O(n525),
    .I0(in[244]),
    .I1(in[239])
  );
  //AND U449bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U449bar (
    .O(n525bar),
    .I0(inbar[244]),
    .I1(inbar[239])
  );
  //OR U450
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U450 (
    .O(n526),
    .I0(in[95]),
    .I1(in[83])
  );
  //AND U450bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U450bar (
    .O(n526bar),
    .I0(inbar[95]),
    .I1(inbar[83])
  );
  //OR U451
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U451 (
    .O(n528),
    .I0(n524),
    .I1(n523)
  );
  //AND U451bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U451bar (
    .O(n528bar),
    .I0(n524bar),
    .I1(n523bar)
  );
  //OR U452
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U452 (
    .O(n523),
    .I0(in_24),
    .I1(in[97])
  );
  //AND U452bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U452bar (
    .O(n523bar),
    .I0(in_24bar),
    .I1(inbar[97])
  );
  //OR U453
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U453 (
    .O(n524),
    .I0(in_33),
    .I1(in_27)
  );
  //AND U453bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U453bar (
    .O(n524bar),
    .I0(in_33bar),
    .I1(in_27bar)
  );
  //OR U454
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U454 (
    .O(n568),
    .I0(n522),
    .I1(n521)
  );
  //AND U454bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U454bar (
    .O(n568bar),
    .I0(n522bar),
    .I1(n521bar)
  );
  //OR U455
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U455 (
    .O(n521),
    .I0(in[145]),
    .I1(in[126])
  );
  //AND U455bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U455bar (
    .O(n521bar),
    .I0(inbar[145]),
    .I1(inbar[126])
  );
  //OR U456
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U456 (
    .O(n522),
    .I0(in[169]),
    .I1(n520)
  );
  //AND U456bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U456bar (
    .O(n522bar),
    .I0(inbar[169]),
    .I1(n520bar)
  );
  //OR U457
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U457 (
    .O(n520),
    .I0(in[221]),
    .I1(in[172])
  );
  //AND U457bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U457bar (
    .O(n520bar),
    .I0(inbar[221]),
    .I1(inbar[172])
  );
  //OR U458
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U458 (
    .O(n570),
    .I0(n519),
    .I1(n518)
  );
  //AND U458bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U458bar (
    .O(n570bar),
    .I0(n519bar),
    .I1(n518bar)
  );
  //OR U459
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U459 (
    .O(n518),
    .I0(n517),
    .I1(n516)
  );
  //AND U459bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U459bar (
    .O(n518bar),
    .I0(n517bar),
    .I1(n516bar)
  );
  //OR U460
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U460 (
    .O(n516),
    .I0(in[241]),
    .I1(in[224])
  );
  //AND U460bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U460bar (
    .O(n516bar),
    .I0(inbar[241]),
    .I1(inbar[224])
  );
  //OR U461
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U461 (
    .O(n517),
    .I0(in[86]),
    .I1(n515)
  );
  //AND U461bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U461bar (
    .O(n517bar),
    .I0(inbar[86]),
    .I1(n515bar)
  );
  //OR U462
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U462 (
    .O(n515),
    .I0(in_43),
    .I1(in_34)
  );
  //AND U462bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U462bar (
    .O(n515bar),
    .I0(in_43bar),
    .I1(in_34bar)
  );
  //OR U463
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U463 (
    .O(n519),
    .I0(n514),
    .I1(n513)
  );
  //AND U463bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U463bar (
    .O(n519bar),
    .I0(n514bar),
    .I1(n513bar)
  );
  //OR U464
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U464 (
    .O(n513),
    .I0(in_65),
    .I1(in_51)
  );
  //AND U464bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U464bar (
    .O(n513bar),
    .I0(in_65bar),
    .I1(in_51bar)
  );
  //OR U465
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U465 (
    .O(n514),
    .I0(in_75),
    .I1(n512)
  );
  //AND U465bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U465bar (
    .O(n514bar),
    .I0(in_75bar),
    .I1(n512bar)
  );
  //OR U466
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U466 (
    .O(n512),
    .I0(in_81),
    .I1(in_77)
  );
  //AND U466bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U466bar (
    .O(n512bar),
    .I0(in_81bar),
    .I1(in_77bar)
  );
  //OR U467
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U467 (
    .O(n778),
    .I0(n511),
    .I1(n510)
  );
  //AND U467bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U467bar (
    .O(n778bar),
    .I0(n511bar),
    .I1(n510bar)
  );
  //OR U468
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U468 (
    .O(n510),
    .I0(n509),
    .I1(n508)
  );
  //AND U468bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U468bar (
    .O(n510bar),
    .I0(n509bar),
    .I1(n508bar)
  );
  //OR U469
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U469 (
    .O(n508),
    .I0(n507),
    .I1(n506)
  );
  //AND U469bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U469bar (
    .O(n508bar),
    .I0(n507bar),
    .I1(n506bar)
  );
  //OR U470
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U470 (
    .O(n506),
    .I0(in[107]),
    .I1(in[101])
  );
  //AND U470bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U470bar (
    .O(n506bar),
    .I0(inbar[107]),
    .I1(inbar[101])
  );
  //OR U471
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U471 (
    .O(n507),
    .I0(in[139]),
    .I1(in[132])
  );
  //AND U471bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U471bar (
    .O(n507bar),
    .I0(inbar[139]),
    .I1(inbar[132])
  );
  //OR U472
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U472 (
    .O(n509),
    .I0(n505),
    .I1(n504)
  );
  //AND U472bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U472bar (
    .O(n509bar),
    .I0(n505bar),
    .I1(n504bar)
  );
  //OR U473
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U473 (
    .O(n504),
    .I0(in[146]),
    .I1(in[141])
  );
  //AND U473bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U473bar (
    .O(n504bar),
    .I0(inbar[146]),
    .I1(inbar[141])
  );
  //OR U474
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U474 (
    .O(n505),
    .I0(in[203]),
    .I1(in[179])
  );
  //AND U474bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U474bar (
    .O(n505bar),
    .I0(inbar[203]),
    .I1(inbar[179])
  );
  //OR U475
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U475 (
    .O(n511),
    .I0(n503),
    .I1(n502)
  );
  //AND U475bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U475bar (
    .O(n511bar),
    .I0(n503bar),
    .I1(n502bar)
  );
  //OR U476
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U476 (
    .O(n502),
    .I0(n501),
    .I1(n500)
  );
  //AND U476bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U476bar (
    .O(n502bar),
    .I0(n501bar),
    .I1(n500bar)
  );
  //OR U477
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U477 (
    .O(n500),
    .I0(in[243]),
    .I1(in[222])
  );
  //AND U477bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U477bar (
    .O(n500bar),
    .I0(inbar[243]),
    .I1(inbar[222])
  );
  //OR U478
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U478 (
    .O(n501),
    .I0(in[251]),
    .I1(in[250])
  );
  //AND U478bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U478bar (
    .O(n501bar),
    .I0(inbar[251]),
    .I1(inbar[250])
  );
  //OR U479
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U479 (
    .O(n503),
    .I0(n499),
    .I1(n498)
  );
  //AND U479bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U479bar (
    .O(n503bar),
    .I0(n499bar),
    .I1(n498bar)
  );
  //OR U480
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U480 (
    .O(n498),
    .I0(in_37),
    .I1(in_19)
  );
  //AND U480bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U480bar (
    .O(n498bar),
    .I0(in_37bar),
    .I1(in_19bar)
  );
  //OR U481
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U481 (
    .O(n499),
    .I0(in_78),
    .I1(in_6)
  );
  //AND U481bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U481bar (
    .O(n499bar),
    .I0(in_78bar),
    .I1(in_6bar)
  );
  //OR U482
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U482 (
    .O(n603),
    .I0(n497),
    .I1(n496)
  );
  //AND U482bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U482bar (
    .O(n603bar),
    .I0(n497bar),
    .I1(n496bar)
  );
  //OR U483
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U483 (
    .O(n496),
    .I0(in[112]),
    .I1(in[102])
  );
  //AND U483bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U483bar (
    .O(n496bar),
    .I0(inbar[112]),
    .I1(inbar[102])
  );
  //OR U484
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U484 (
    .O(n497),
    .I0(in[123]),
    .I1(n495)
  );
  //AND U484bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U484bar (
    .O(n497bar),
    .I0(inbar[123]),
    .I1(n495bar)
  );
  //OR U485
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U485 (
    .O(n495),
    .I0(in[143]),
    .I1(in[130])
  );
  //AND U485bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U485bar (
    .O(n495bar),
    .I0(inbar[143]),
    .I1(inbar[130])
  );
  //OR U486
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U486 (
    .O(n605),
    .I0(n494),
    .I1(n493)
  );
  //AND U486bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U486bar (
    .O(n605bar),
    .I0(n494bar),
    .I1(n493bar)
  );
  //OR U487
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U487 (
    .O(n493),
    .I0(n492),
    .I1(n491)
  );
  //AND U487bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U487bar (
    .O(n493bar),
    .I0(n492bar),
    .I1(n491bar)
  );
  //OR U488
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U488 (
    .O(n491),
    .I0(in[216]),
    .I1(in[213])
  );
  //AND U488bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U488bar (
    .O(n491bar),
    .I0(inbar[216]),
    .I1(inbar[213])
  );
  //OR U489
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U489 (
    .O(n492),
    .I0(in[227]),
    .I1(n490)
  );
  //AND U489bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U489bar (
    .O(n492bar),
    .I0(inbar[227]),
    .I1(n490bar)
  );
  //OR U490
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U490 (
    .O(n490),
    .I0(in_0),
    .I1(in[248])
  );
  //AND U490bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U490bar (
    .O(n490bar),
    .I0(in_0bar),
    .I1(inbar[248])
  );
  //OR U491
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U491 (
    .O(n494),
    .I0(n489),
    .I1(n488)
  );
  //AND U491bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U491bar (
    .O(n494bar),
    .I0(n489bar),
    .I1(n488bar)
  );
  //OR U492
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U492 (
    .O(n488),
    .I0(in_46),
    .I1(in_44)
  );
  //AND U492bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U492bar (
    .O(n488bar),
    .I0(in_46bar),
    .I1(in_44bar)
  );
  //OR U493
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U493 (
    .O(n489),
    .I0(in_50),
    .I1(n487)
  );
  //AND U493bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U493bar (
    .O(n489bar),
    .I0(in_50bar),
    .I1(n487bar)
  );
  //OR U494
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U494 (
    .O(n487),
    .I0(in_9),
    .I1(in_80)
  );
  //AND U494bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U494bar (
    .O(n487bar),
    .I0(in_9bar),
    .I1(in_80bar)
  );
endmodule

module sBox_3 ( in, out );

  input wire [7:0] in;
//input_done

  output wire [7:0] out;
//output_done

  wire [255:0] decodeOut;
//wire_done

  decode_3 dec ( .in(in), .out(decodeOut) );
  encode_3 enc ( .in(decodeOut), .out(out) );
endmodule

module CD2_13 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD2_14 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD2_15 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD2_16 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD4_7 ( a, b, y );

  input wire [3:0] a;
  input wire [3:0] b;
  wire [3:0] abar;
  wire [3:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
//input_done

  output wire [15:0] y;
  wire [15:0] ybar;
//output_done

//wire_done

  //AND U1
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1 (
    .O(y[9]),
    .I0(b[1]),
    .I1(a[2])
  );
  //OR U1bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1bar (
    .O(ybar[9]),
    .I0(bbar[1]),
    .I1(abar[2])
  );
  //AND U2
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2 (
    .O(y[8]),
    .I0(b[0]),
    .I1(a[2])
  );
  //OR U2bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2bar (
    .O(ybar[8]),
    .I0(bbar[0]),
    .I1(abar[2])
  );
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[7]),
    .I0(b[3]),
    .I1(a[1])
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[7]),
    .I0(bbar[3]),
    .I1(abar[1])
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[6]),
    .I0(b[2]),
    .I1(a[1])
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[6]),
    .I0(bbar[2]),
    .I1(abar[1])
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[5]),
    .I0(a[1]),
    .I1(b[1])
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[5]),
    .I0(abar[1]),
    .I1(bbar[1])
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[4]),
    .I0(a[1]),
    .I1(b[0])
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[4]),
    .I0(abar[1]),
    .I1(bbar[0])
  );
  //AND U7
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7 (
    .O(y[3]),
    .I0(a[0]),
    .I1(b[3])
  );
  //OR U7bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7bar (
    .O(ybar[3]),
    .I0(abar[0]),
    .I1(bbar[3])
  );
  //AND U8
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8 (
    .O(y[2]),
    .I0(a[0]),
    .I1(b[2])
  );
  //OR U8bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8bar (
    .O(ybar[2]),
    .I0(abar[0]),
    .I1(bbar[2])
  );
  //AND U9
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9 (
    .O(y[1]),
    .I0(a[0]),
    .I1(b[1])
  );
  //OR U9bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9bar (
    .O(ybar[1]),
    .I0(abar[0]),
    .I1(bbar[1])
  );
  //AND U10
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10 (
    .O(y[15]),
    .I0(a[3]),
    .I1(b[3])
  );
  //OR U10bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10bar (
    .O(ybar[15]),
    .I0(abar[3]),
    .I1(bbar[3])
  );
  //AND U11
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11 (
    .O(y[14]),
    .I0(a[3]),
    .I1(b[2])
  );
  //OR U11bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11bar (
    .O(ybar[14]),
    .I0(abar[3]),
    .I1(bbar[2])
  );
  //AND U12
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12 (
    .O(y[13]),
    .I0(a[3]),
    .I1(b[1])
  );
  //OR U12bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12bar (
    .O(ybar[13]),
    .I0(abar[3]),
    .I1(bbar[1])
  );
  //AND U13
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13 (
    .O(y[12]),
    .I0(a[3]),
    .I1(b[0])
  );
  //OR U13bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13bar (
    .O(ybar[12]),
    .I0(abar[3]),
    .I1(bbar[0])
  );
  //AND U14
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14 (
    .O(y[11]),
    .I0(b[3]),
    .I1(a[2])
  );
  //OR U14bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14bar (
    .O(ybar[11]),
    .I0(bbar[3]),
    .I1(abar[2])
  );
  //AND U15
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15 (
    .O(y[10]),
    .I0(b[2]),
    .I1(a[2])
  );
  //OR U15bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15bar (
    .O(ybar[10]),
    .I0(bbar[2]),
    .I1(abar[2])
  );
  //AND U16
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16 (
    .O(y[0]),
    .I0(a[0]),
    .I1(b[0])
  );
  //OR U16bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16bar (
    .O(ybar[0]),
    .I0(abar[0]),
    .I1(bbar[0])
  );
endmodule

module CD4_8 ( a, b, y );

  input wire [3:0] a;
  input wire [3:0] b;
  wire [3:0] abar;
  wire [3:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
//input_done

  output wire [15:0] y;
  wire [15:0] ybar;
//output_done

//wire_done

  //AND U1
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1 (
    .O(y[9]),
    .I0(b[1]),
    .I1(a[2])
  );
  //OR U1bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1bar (
    .O(ybar[9]),
    .I0(bbar[1]),
    .I1(abar[2])
  );
  //AND U2
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2 (
    .O(y[8]),
    .I0(b[0]),
    .I1(a[2])
  );
  //OR U2bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2bar (
    .O(ybar[8]),
    .I0(bbar[0]),
    .I1(abar[2])
  );
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[7]),
    .I0(b[3]),
    .I1(a[1])
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[7]),
    .I0(bbar[3]),
    .I1(abar[1])
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[6]),
    .I0(b[2]),
    .I1(a[1])
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[6]),
    .I0(bbar[2]),
    .I1(abar[1])
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[5]),
    .I0(a[1]),
    .I1(b[1])
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[5]),
    .I0(abar[1]),
    .I1(bbar[1])
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[4]),
    .I0(a[1]),
    .I1(b[0])
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[4]),
    .I0(abar[1]),
    .I1(bbar[0])
  );
  //AND U7
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7 (
    .O(y[3]),
    .I0(a[0]),
    .I1(b[3])
  );
  //OR U7bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7bar (
    .O(ybar[3]),
    .I0(abar[0]),
    .I1(bbar[3])
  );
  //AND U8
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8 (
    .O(y[2]),
    .I0(a[0]),
    .I1(b[2])
  );
  //OR U8bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8bar (
    .O(ybar[2]),
    .I0(abar[0]),
    .I1(bbar[2])
  );
  //AND U9
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9 (
    .O(y[1]),
    .I0(a[0]),
    .I1(b[1])
  );
  //OR U9bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9bar (
    .O(ybar[1]),
    .I0(abar[0]),
    .I1(bbar[1])
  );
  //AND U10
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10 (
    .O(y[15]),
    .I0(a[3]),
    .I1(b[3])
  );
  //OR U10bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10bar (
    .O(ybar[15]),
    .I0(abar[3]),
    .I1(bbar[3])
  );
  //AND U11
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11 (
    .O(y[14]),
    .I0(a[3]),
    .I1(b[2])
  );
  //OR U11bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11bar (
    .O(ybar[14]),
    .I0(abar[3]),
    .I1(bbar[2])
  );
  //AND U12
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12 (
    .O(y[13]),
    .I0(a[3]),
    .I1(b[1])
  );
  //OR U12bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12bar (
    .O(ybar[13]),
    .I0(abar[3]),
    .I1(bbar[1])
  );
  //AND U13
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13 (
    .O(y[12]),
    .I0(a[3]),
    .I1(b[0])
  );
  //OR U13bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13bar (
    .O(ybar[12]),
    .I0(abar[3]),
    .I1(bbar[0])
  );
  //AND U14
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14 (
    .O(y[11]),
    .I0(b[3]),
    .I1(a[2])
  );
  //OR U14bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14bar (
    .O(ybar[11]),
    .I0(bbar[3]),
    .I1(abar[2])
  );
  //AND U15
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15 (
    .O(y[10]),
    .I0(b[2]),
    .I1(a[2])
  );
  //OR U15bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15bar (
    .O(ybar[10]),
    .I0(bbar[2]),
    .I1(abar[2])
  );
  //AND U16
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16 (
    .O(y[0]),
    .I0(a[0]),
    .I1(b[0])
  );
  //OR U16bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16bar (
    .O(ybar[0]),
    .I0(abar[0]),
    .I1(bbar[0])
  );
endmodule

module CD16_4 ( a, b, y );

  input wire [15:0] a;
  input wire [15:0] b;
  wire [15:0] abar;
  wire [15:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign abar[8] = ~a[8];
  assign abar[9] = ~a[9];
  assign abar[10] = ~a[10];
  assign abar[11] = ~a[11];
  assign abar[12] = ~a[12];
  assign abar[13] = ~a[13];
  assign abar[14] = ~a[14];
  assign abar[15] = ~a[15];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign bbar[8] = ~b[8];
  assign bbar[9] = ~b[9];
  assign bbar[10] = ~b[10];
  assign bbar[11] = ~b[11];
  assign bbar[12] = ~b[12];
  assign bbar[13] = ~b[13];
  assign bbar[14] = ~b[14];
  assign bbar[15] = ~b[15];
//input_done

  output wire [255:0] y;
  wire [255:0] ybar;
//output_done

//wire_done

  //AND U1
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1 (
    .O(y[9]),
    .I0(b[9]),
    .I1(a[0])
  );
  //OR U1bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1bar (
    .O(ybar[9]),
    .I0(bbar[9]),
    .I1(abar[0])
  );
  //AND U2
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2 (
    .O(y[99]),
    .I0(b[3]),
    .I1(a[6])
  );
  //OR U2bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2bar (
    .O(ybar[99]),
    .I0(bbar[3]),
    .I1(abar[6])
  );
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[98]),
    .I0(b[2]),
    .I1(a[6])
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[98]),
    .I0(bbar[2]),
    .I1(abar[6])
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[97]),
    .I0(b[1]),
    .I1(a[6])
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[97]),
    .I0(bbar[1]),
    .I1(abar[6])
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[96]),
    .I0(b[0]),
    .I1(a[6])
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[96]),
    .I0(bbar[0]),
    .I1(abar[6])
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[95]),
    .I0(b[15]),
    .I1(a[5])
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[95]),
    .I0(bbar[15]),
    .I1(abar[5])
  );
  //AND U7
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7 (
    .O(y[94]),
    .I0(b[14]),
    .I1(a[5])
  );
  //OR U7bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7bar (
    .O(ybar[94]),
    .I0(bbar[14]),
    .I1(abar[5])
  );
  //AND U8
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8 (
    .O(y[93]),
    .I0(b[13]),
    .I1(a[5])
  );
  //OR U8bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8bar (
    .O(ybar[93]),
    .I0(bbar[13]),
    .I1(abar[5])
  );
  //AND U9
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9 (
    .O(y[92]),
    .I0(b[12]),
    .I1(a[5])
  );
  //OR U9bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9bar (
    .O(ybar[92]),
    .I0(bbar[12]),
    .I1(abar[5])
  );
  //AND U10
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10 (
    .O(y[91]),
    .I0(b[11]),
    .I1(a[5])
  );
  //OR U10bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10bar (
    .O(ybar[91]),
    .I0(bbar[11]),
    .I1(abar[5])
  );
  //AND U11
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11 (
    .O(y[90]),
    .I0(b[10]),
    .I1(a[5])
  );
  //OR U11bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11bar (
    .O(ybar[90]),
    .I0(bbar[10]),
    .I1(abar[5])
  );
  //AND U12
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12 (
    .O(y[8]),
    .I0(b[8]),
    .I1(a[0])
  );
  //OR U12bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12bar (
    .O(ybar[8]),
    .I0(bbar[8]),
    .I1(abar[0])
  );
  //AND U13
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13 (
    .O(y[89]),
    .I0(a[5]),
    .I1(b[9])
  );
  //OR U13bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13bar (
    .O(ybar[89]),
    .I0(abar[5]),
    .I1(bbar[9])
  );
  //AND U14
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14 (
    .O(y[88]),
    .I0(b[8]),
    .I1(a[5])
  );
  //OR U14bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14bar (
    .O(ybar[88]),
    .I0(bbar[8]),
    .I1(abar[5])
  );
  //AND U15
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15 (
    .O(y[87]),
    .I0(b[7]),
    .I1(a[5])
  );
  //OR U15bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15bar (
    .O(ybar[87]),
    .I0(bbar[7]),
    .I1(abar[5])
  );
  //AND U16
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16 (
    .O(y[86]),
    .I0(b[6]),
    .I1(a[5])
  );
  //OR U16bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16bar (
    .O(ybar[86]),
    .I0(bbar[6]),
    .I1(abar[5])
  );
  //AND U17
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U17 (
    .O(y[85]),
    .I0(b[5]),
    .I1(a[5])
  );
  //OR U17bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U17bar (
    .O(ybar[85]),
    .I0(bbar[5]),
    .I1(abar[5])
  );
  //AND U18
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U18 (
    .O(y[84]),
    .I0(b[4]),
    .I1(a[5])
  );
  //OR U18bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U18bar (
    .O(ybar[84]),
    .I0(bbar[4]),
    .I1(abar[5])
  );
  //AND U19
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U19 (
    .O(y[83]),
    .I0(a[5]),
    .I1(b[3])
  );
  //OR U19bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U19bar (
    .O(ybar[83]),
    .I0(abar[5]),
    .I1(bbar[3])
  );
  //AND U20
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U20 (
    .O(y[82]),
    .I0(a[5]),
    .I1(b[2])
  );
  //OR U20bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U20bar (
    .O(ybar[82]),
    .I0(abar[5]),
    .I1(bbar[2])
  );
  //AND U21
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U21 (
    .O(y[81]),
    .I0(a[5]),
    .I1(b[1])
  );
  //OR U21bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U21bar (
    .O(ybar[81]),
    .I0(abar[5]),
    .I1(bbar[1])
  );
  //AND U22
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U22 (
    .O(y[80]),
    .I0(a[5]),
    .I1(b[0])
  );
  //OR U22bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U22bar (
    .O(ybar[80]),
    .I0(abar[5]),
    .I1(bbar[0])
  );
  //AND U23
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U23 (
    .O(y[7]),
    .I0(b[7]),
    .I1(a[0])
  );
  //OR U23bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U23bar (
    .O(ybar[7]),
    .I0(bbar[7]),
    .I1(abar[0])
  );
  //AND U24
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U24 (
    .O(y[79]),
    .I0(a[4]),
    .I1(b[15])
  );
  //OR U24bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U24bar (
    .O(ybar[79]),
    .I0(abar[4]),
    .I1(bbar[15])
  );
  //AND U25
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U25 (
    .O(y[78]),
    .I0(a[4]),
    .I1(b[14])
  );
  //OR U25bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U25bar (
    .O(ybar[78]),
    .I0(abar[4]),
    .I1(bbar[14])
  );
  //AND U26
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U26 (
    .O(y[77]),
    .I0(a[4]),
    .I1(b[13])
  );
  //OR U26bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U26bar (
    .O(ybar[77]),
    .I0(abar[4]),
    .I1(bbar[13])
  );
  //AND U27
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U27 (
    .O(y[76]),
    .I0(a[4]),
    .I1(b[12])
  );
  //OR U27bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U27bar (
    .O(ybar[76]),
    .I0(abar[4]),
    .I1(bbar[12])
  );
  //AND U28
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U28 (
    .O(y[75]),
    .I0(a[4]),
    .I1(b[11])
  );
  //OR U28bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U28bar (
    .O(ybar[75]),
    .I0(abar[4]),
    .I1(bbar[11])
  );
  //AND U29
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U29 (
    .O(y[74]),
    .I0(a[4]),
    .I1(b[10])
  );
  //OR U29bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U29bar (
    .O(ybar[74]),
    .I0(abar[4]),
    .I1(bbar[10])
  );
  //AND U30
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U30 (
    .O(y[73]),
    .I0(a[4]),
    .I1(b[9])
  );
  //OR U30bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U30bar (
    .O(ybar[73]),
    .I0(abar[4]),
    .I1(bbar[9])
  );
  //AND U31
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U31 (
    .O(y[72]),
    .I0(a[4]),
    .I1(b[8])
  );
  //OR U31bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U31bar (
    .O(ybar[72]),
    .I0(abar[4]),
    .I1(bbar[8])
  );
  //AND U32
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U32 (
    .O(y[71]),
    .I0(a[4]),
    .I1(b[7])
  );
  //OR U32bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U32bar (
    .O(ybar[71]),
    .I0(abar[4]),
    .I1(bbar[7])
  );
  //AND U33
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U33 (
    .O(y[70]),
    .I0(a[4]),
    .I1(b[6])
  );
  //OR U33bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U33bar (
    .O(ybar[70]),
    .I0(abar[4]),
    .I1(bbar[6])
  );
  //AND U34
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U34 (
    .O(y[6]),
    .I0(b[6]),
    .I1(a[0])
  );
  //OR U34bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U34bar (
    .O(ybar[6]),
    .I0(bbar[6]),
    .I1(abar[0])
  );
  //AND U35
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U35 (
    .O(y[69]),
    .I0(a[4]),
    .I1(b[5])
  );
  //OR U35bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U35bar (
    .O(ybar[69]),
    .I0(abar[4]),
    .I1(bbar[5])
  );
  //AND U36
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U36 (
    .O(y[68]),
    .I0(a[4]),
    .I1(b[4])
  );
  //OR U36bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U36bar (
    .O(ybar[68]),
    .I0(abar[4]),
    .I1(bbar[4])
  );
  //AND U37
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U37 (
    .O(y[67]),
    .I0(a[4]),
    .I1(b[3])
  );
  //OR U37bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U37bar (
    .O(ybar[67]),
    .I0(abar[4]),
    .I1(bbar[3])
  );
  //AND U38
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U38 (
    .O(y[66]),
    .I0(a[4]),
    .I1(b[2])
  );
  //OR U38bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U38bar (
    .O(ybar[66]),
    .I0(abar[4]),
    .I1(bbar[2])
  );
  //AND U39
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U39 (
    .O(y[65]),
    .I0(a[4]),
    .I1(b[1])
  );
  //OR U39bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U39bar (
    .O(ybar[65]),
    .I0(abar[4]),
    .I1(bbar[1])
  );
  //AND U40
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U40 (
    .O(y[64]),
    .I0(a[4]),
    .I1(b[0])
  );
  //OR U40bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U40bar (
    .O(ybar[64]),
    .I0(abar[4]),
    .I1(bbar[0])
  );
  //AND U41
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U41 (
    .O(y[63]),
    .I0(a[3]),
    .I1(b[15])
  );
  //OR U41bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U41bar (
    .O(ybar[63]),
    .I0(abar[3]),
    .I1(bbar[15])
  );
  //AND U42
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U42 (
    .O(y[62]),
    .I0(a[3]),
    .I1(b[14])
  );
  //OR U42bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U42bar (
    .O(ybar[62]),
    .I0(abar[3]),
    .I1(bbar[14])
  );
  //AND U43
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U43 (
    .O(y[61]),
    .I0(a[3]),
    .I1(b[13])
  );
  //OR U43bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U43bar (
    .O(ybar[61]),
    .I0(abar[3]),
    .I1(bbar[13])
  );
  //AND U44
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U44 (
    .O(y[60]),
    .I0(a[3]),
    .I1(b[12])
  );
  //OR U44bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U44bar (
    .O(ybar[60]),
    .I0(abar[3]),
    .I1(bbar[12])
  );
  //AND U45
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U45 (
    .O(y[5]),
    .I0(b[5]),
    .I1(a[0])
  );
  //OR U45bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U45bar (
    .O(ybar[5]),
    .I0(bbar[5]),
    .I1(abar[0])
  );
  //AND U46
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U46 (
    .O(y[59]),
    .I0(a[3]),
    .I1(b[11])
  );
  //OR U46bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U46bar (
    .O(ybar[59]),
    .I0(abar[3]),
    .I1(bbar[11])
  );
  //AND U47
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U47 (
    .O(y[58]),
    .I0(a[3]),
    .I1(b[10])
  );
  //OR U47bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U47bar (
    .O(ybar[58]),
    .I0(abar[3]),
    .I1(bbar[10])
  );
  //AND U48
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U48 (
    .O(y[57]),
    .I0(a[3]),
    .I1(b[9])
  );
  //OR U48bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U48bar (
    .O(ybar[57]),
    .I0(abar[3]),
    .I1(bbar[9])
  );
  //AND U49
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U49 (
    .O(y[56]),
    .I0(a[3]),
    .I1(b[8])
  );
  //OR U49bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U49bar (
    .O(ybar[56]),
    .I0(abar[3]),
    .I1(bbar[8])
  );
  //AND U50
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U50 (
    .O(y[55]),
    .I0(a[3]),
    .I1(b[7])
  );
  //OR U50bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U50bar (
    .O(ybar[55]),
    .I0(abar[3]),
    .I1(bbar[7])
  );
  //AND U51
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U51 (
    .O(y[54]),
    .I0(a[3]),
    .I1(b[6])
  );
  //OR U51bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U51bar (
    .O(ybar[54]),
    .I0(abar[3]),
    .I1(bbar[6])
  );
  //AND U52
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U52 (
    .O(y[53]),
    .I0(a[3]),
    .I1(b[5])
  );
  //OR U52bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U52bar (
    .O(ybar[53]),
    .I0(abar[3]),
    .I1(bbar[5])
  );
  //AND U53
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U53 (
    .O(y[52]),
    .I0(a[3]),
    .I1(b[4])
  );
  //OR U53bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U53bar (
    .O(ybar[52]),
    .I0(abar[3]),
    .I1(bbar[4])
  );
  //AND U54
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U54 (
    .O(y[51]),
    .I0(a[3]),
    .I1(b[3])
  );
  //OR U54bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U54bar (
    .O(ybar[51]),
    .I0(abar[3]),
    .I1(bbar[3])
  );
  //AND U55
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U55 (
    .O(y[50]),
    .I0(a[3]),
    .I1(b[2])
  );
  //OR U55bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U55bar (
    .O(ybar[50]),
    .I0(abar[3]),
    .I1(bbar[2])
  );
  //AND U56
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U56 (
    .O(y[4]),
    .I0(b[4]),
    .I1(a[0])
  );
  //OR U56bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U56bar (
    .O(ybar[4]),
    .I0(bbar[4]),
    .I1(abar[0])
  );
  //AND U57
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U57 (
    .O(y[49]),
    .I0(a[3]),
    .I1(b[1])
  );
  //OR U57bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U57bar (
    .O(ybar[49]),
    .I0(abar[3]),
    .I1(bbar[1])
  );
  //AND U58
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U58 (
    .O(y[48]),
    .I0(a[3]),
    .I1(b[0])
  );
  //OR U58bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U58bar (
    .O(ybar[48]),
    .I0(abar[3]),
    .I1(bbar[0])
  );
  //AND U59
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U59 (
    .O(y[47]),
    .I0(a[2]),
    .I1(b[15])
  );
  //OR U59bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U59bar (
    .O(ybar[47]),
    .I0(abar[2]),
    .I1(bbar[15])
  );
  //AND U60
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U60 (
    .O(y[46]),
    .I0(a[2]),
    .I1(b[14])
  );
  //OR U60bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U60bar (
    .O(ybar[46]),
    .I0(abar[2]),
    .I1(bbar[14])
  );
  //AND U61
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U61 (
    .O(y[45]),
    .I0(a[2]),
    .I1(b[13])
  );
  //OR U61bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U61bar (
    .O(ybar[45]),
    .I0(abar[2]),
    .I1(bbar[13])
  );
  //AND U62
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U62 (
    .O(y[44]),
    .I0(a[2]),
    .I1(b[12])
  );
  //OR U62bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U62bar (
    .O(ybar[44]),
    .I0(abar[2]),
    .I1(bbar[12])
  );
  //AND U63
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U63 (
    .O(y[43]),
    .I0(a[2]),
    .I1(b[11])
  );
  //OR U63bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U63bar (
    .O(ybar[43]),
    .I0(abar[2]),
    .I1(bbar[11])
  );
  //AND U64
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U64 (
    .O(y[42]),
    .I0(a[2]),
    .I1(b[10])
  );
  //OR U64bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U64bar (
    .O(ybar[42]),
    .I0(abar[2]),
    .I1(bbar[10])
  );
  //AND U65
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U65 (
    .O(y[41]),
    .I0(a[2]),
    .I1(b[9])
  );
  //OR U65bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U65bar (
    .O(ybar[41]),
    .I0(abar[2]),
    .I1(bbar[9])
  );
  //AND U66
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U66 (
    .O(y[40]),
    .I0(a[2]),
    .I1(b[8])
  );
  //OR U66bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U66bar (
    .O(ybar[40]),
    .I0(abar[2]),
    .I1(bbar[8])
  );
  //AND U67
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U67 (
    .O(y[3]),
    .I0(b[3]),
    .I1(a[0])
  );
  //OR U67bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U67bar (
    .O(ybar[3]),
    .I0(bbar[3]),
    .I1(abar[0])
  );
  //AND U68
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U68 (
    .O(y[39]),
    .I0(a[2]),
    .I1(b[7])
  );
  //OR U68bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U68bar (
    .O(ybar[39]),
    .I0(abar[2]),
    .I1(bbar[7])
  );
  //AND U69
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U69 (
    .O(y[38]),
    .I0(a[2]),
    .I1(b[6])
  );
  //OR U69bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U69bar (
    .O(ybar[38]),
    .I0(abar[2]),
    .I1(bbar[6])
  );
  //AND U70
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U70 (
    .O(y[37]),
    .I0(a[2]),
    .I1(b[5])
  );
  //OR U70bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U70bar (
    .O(ybar[37]),
    .I0(abar[2]),
    .I1(bbar[5])
  );
  //AND U71
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U71 (
    .O(y[36]),
    .I0(a[2]),
    .I1(b[4])
  );
  //OR U71bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U71bar (
    .O(ybar[36]),
    .I0(abar[2]),
    .I1(bbar[4])
  );
  //AND U72
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U72 (
    .O(y[35]),
    .I0(a[2]),
    .I1(b[3])
  );
  //OR U72bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U72bar (
    .O(ybar[35]),
    .I0(abar[2]),
    .I1(bbar[3])
  );
  //AND U73
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U73 (
    .O(y[34]),
    .I0(a[2]),
    .I1(b[2])
  );
  //OR U73bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U73bar (
    .O(ybar[34]),
    .I0(abar[2]),
    .I1(bbar[2])
  );
  //AND U74
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U74 (
    .O(y[33]),
    .I0(a[2]),
    .I1(b[1])
  );
  //OR U74bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U74bar (
    .O(ybar[33]),
    .I0(abar[2]),
    .I1(bbar[1])
  );
  //AND U75
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U75 (
    .O(y[32]),
    .I0(a[2]),
    .I1(b[0])
  );
  //OR U75bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U75bar (
    .O(ybar[32]),
    .I0(abar[2]),
    .I1(bbar[0])
  );
  //AND U76
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U76 (
    .O(y[31]),
    .I0(a[1]),
    .I1(b[15])
  );
  //OR U76bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U76bar (
    .O(ybar[31]),
    .I0(abar[1]),
    .I1(bbar[15])
  );
  //AND U77
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U77 (
    .O(y[30]),
    .I0(a[1]),
    .I1(b[14])
  );
  //OR U77bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U77bar (
    .O(ybar[30]),
    .I0(abar[1]),
    .I1(bbar[14])
  );
  //AND U78
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U78 (
    .O(y[2]),
    .I0(b[2]),
    .I1(a[0])
  );
  //OR U78bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U78bar (
    .O(ybar[2]),
    .I0(bbar[2]),
    .I1(abar[0])
  );
  //AND U79
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U79 (
    .O(y[29]),
    .I0(a[1]),
    .I1(b[13])
  );
  //OR U79bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U79bar (
    .O(ybar[29]),
    .I0(abar[1]),
    .I1(bbar[13])
  );
  //AND U80
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U80 (
    .O(y[28]),
    .I0(a[1]),
    .I1(b[12])
  );
  //OR U80bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U80bar (
    .O(ybar[28]),
    .I0(abar[1]),
    .I1(bbar[12])
  );
  //AND U81
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U81 (
    .O(y[27]),
    .I0(a[1]),
    .I1(b[11])
  );
  //OR U81bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U81bar (
    .O(ybar[27]),
    .I0(abar[1]),
    .I1(bbar[11])
  );
  //AND U82
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U82 (
    .O(y[26]),
    .I0(a[1]),
    .I1(b[10])
  );
  //OR U82bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U82bar (
    .O(ybar[26]),
    .I0(abar[1]),
    .I1(bbar[10])
  );
  //AND U83
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U83 (
    .O(y[25]),
    .I0(a[1]),
    .I1(b[9])
  );
  //OR U83bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U83bar (
    .O(ybar[25]),
    .I0(abar[1]),
    .I1(bbar[9])
  );
  //AND U84
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U84 (
    .O(y[255]),
    .I0(a[15]),
    .I1(b[15])
  );
  //OR U84bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U84bar (
    .O(ybar[255]),
    .I0(abar[15]),
    .I1(bbar[15])
  );
  //AND U85
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U85 (
    .O(y[254]),
    .I0(a[15]),
    .I1(b[14])
  );
  //OR U85bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U85bar (
    .O(ybar[254]),
    .I0(abar[15]),
    .I1(bbar[14])
  );
  //AND U86
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U86 (
    .O(y[253]),
    .I0(a[15]),
    .I1(b[13])
  );
  //OR U86bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U86bar (
    .O(ybar[253]),
    .I0(abar[15]),
    .I1(bbar[13])
  );
  //AND U87
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U87 (
    .O(y[252]),
    .I0(a[15]),
    .I1(b[12])
  );
  //OR U87bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U87bar (
    .O(ybar[252]),
    .I0(abar[15]),
    .I1(bbar[12])
  );
  //AND U88
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U88 (
    .O(y[251]),
    .I0(a[15]),
    .I1(b[11])
  );
  //OR U88bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U88bar (
    .O(ybar[251]),
    .I0(abar[15]),
    .I1(bbar[11])
  );
  //AND U89
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U89 (
    .O(y[250]),
    .I0(a[15]),
    .I1(b[10])
  );
  //OR U89bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U89bar (
    .O(ybar[250]),
    .I0(abar[15]),
    .I1(bbar[10])
  );
  //AND U90
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U90 (
    .O(y[24]),
    .I0(a[1]),
    .I1(b[8])
  );
  //OR U90bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U90bar (
    .O(ybar[24]),
    .I0(abar[1]),
    .I1(bbar[8])
  );
  //AND U91
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U91 (
    .O(y[249]),
    .I0(a[15]),
    .I1(b[9])
  );
  //OR U91bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U91bar (
    .O(ybar[249]),
    .I0(abar[15]),
    .I1(bbar[9])
  );
  //AND U92
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U92 (
    .O(y[248]),
    .I0(a[15]),
    .I1(b[8])
  );
  //OR U92bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U92bar (
    .O(ybar[248]),
    .I0(abar[15]),
    .I1(bbar[8])
  );
  //AND U93
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U93 (
    .O(y[247]),
    .I0(a[15]),
    .I1(b[7])
  );
  //OR U93bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U93bar (
    .O(ybar[247]),
    .I0(abar[15]),
    .I1(bbar[7])
  );
  //AND U94
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U94 (
    .O(y[246]),
    .I0(a[15]),
    .I1(b[6])
  );
  //OR U94bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U94bar (
    .O(ybar[246]),
    .I0(abar[15]),
    .I1(bbar[6])
  );
  //AND U95
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U95 (
    .O(y[245]),
    .I0(a[15]),
    .I1(b[5])
  );
  //OR U95bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U95bar (
    .O(ybar[245]),
    .I0(abar[15]),
    .I1(bbar[5])
  );
  //AND U96
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U96 (
    .O(y[244]),
    .I0(a[15]),
    .I1(b[4])
  );
  //OR U96bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U96bar (
    .O(ybar[244]),
    .I0(abar[15]),
    .I1(bbar[4])
  );
  //AND U97
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U97 (
    .O(y[243]),
    .I0(a[15]),
    .I1(b[3])
  );
  //OR U97bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U97bar (
    .O(ybar[243]),
    .I0(abar[15]),
    .I1(bbar[3])
  );
  //AND U98
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U98 (
    .O(y[242]),
    .I0(a[15]),
    .I1(b[2])
  );
  //OR U98bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U98bar (
    .O(ybar[242]),
    .I0(abar[15]),
    .I1(bbar[2])
  );
  //AND U99
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U99 (
    .O(y[241]),
    .I0(a[15]),
    .I1(b[1])
  );
  //OR U99bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U99bar (
    .O(ybar[241]),
    .I0(abar[15]),
    .I1(bbar[1])
  );
  //AND U100
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U100 (
    .O(y[240]),
    .I0(a[15]),
    .I1(b[0])
  );
  //OR U100bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U100bar (
    .O(ybar[240]),
    .I0(abar[15]),
    .I1(bbar[0])
  );
  //AND U101
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U101 (
    .O(y[23]),
    .I0(a[1]),
    .I1(b[7])
  );
  //OR U101bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U101bar (
    .O(ybar[23]),
    .I0(abar[1]),
    .I1(bbar[7])
  );
  //AND U102
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U102 (
    .O(y[239]),
    .I0(a[14]),
    .I1(b[15])
  );
  //OR U102bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U102bar (
    .O(ybar[239]),
    .I0(abar[14]),
    .I1(bbar[15])
  );
  //AND U103
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U103 (
    .O(y[238]),
    .I0(a[14]),
    .I1(b[14])
  );
  //OR U103bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U103bar (
    .O(ybar[238]),
    .I0(abar[14]),
    .I1(bbar[14])
  );
  //AND U104
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U104 (
    .O(y[237]),
    .I0(a[14]),
    .I1(b[13])
  );
  //OR U104bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U104bar (
    .O(ybar[237]),
    .I0(abar[14]),
    .I1(bbar[13])
  );
  //AND U105
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U105 (
    .O(y[236]),
    .I0(a[14]),
    .I1(b[12])
  );
  //OR U105bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U105bar (
    .O(ybar[236]),
    .I0(abar[14]),
    .I1(bbar[12])
  );
  //AND U106
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U106 (
    .O(y[235]),
    .I0(a[14]),
    .I1(b[11])
  );
  //OR U106bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U106bar (
    .O(ybar[235]),
    .I0(abar[14]),
    .I1(bbar[11])
  );
  //AND U107
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U107 (
    .O(y[234]),
    .I0(a[14]),
    .I1(b[10])
  );
  //OR U107bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U107bar (
    .O(ybar[234]),
    .I0(abar[14]),
    .I1(bbar[10])
  );
  //AND U108
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U108 (
    .O(y[233]),
    .I0(a[14]),
    .I1(b[9])
  );
  //OR U108bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U108bar (
    .O(ybar[233]),
    .I0(abar[14]),
    .I1(bbar[9])
  );
  //AND U109
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U109 (
    .O(y[232]),
    .I0(a[14]),
    .I1(b[8])
  );
  //OR U109bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U109bar (
    .O(ybar[232]),
    .I0(abar[14]),
    .I1(bbar[8])
  );
  //AND U110
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U110 (
    .O(y[231]),
    .I0(a[14]),
    .I1(b[7])
  );
  //OR U110bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U110bar (
    .O(ybar[231]),
    .I0(abar[14]),
    .I1(bbar[7])
  );
  //AND U111
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U111 (
    .O(y[230]),
    .I0(a[14]),
    .I1(b[6])
  );
  //OR U111bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U111bar (
    .O(ybar[230]),
    .I0(abar[14]),
    .I1(bbar[6])
  );
  //AND U112
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U112 (
    .O(y[22]),
    .I0(a[1]),
    .I1(b[6])
  );
  //OR U112bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U112bar (
    .O(ybar[22]),
    .I0(abar[1]),
    .I1(bbar[6])
  );
  //AND U113
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U113 (
    .O(y[229]),
    .I0(a[14]),
    .I1(b[5])
  );
  //OR U113bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U113bar (
    .O(ybar[229]),
    .I0(abar[14]),
    .I1(bbar[5])
  );
  //AND U114
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U114 (
    .O(y[228]),
    .I0(a[14]),
    .I1(b[4])
  );
  //OR U114bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U114bar (
    .O(ybar[228]),
    .I0(abar[14]),
    .I1(bbar[4])
  );
  //AND U115
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U115 (
    .O(y[227]),
    .I0(a[14]),
    .I1(b[3])
  );
  //OR U115bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U115bar (
    .O(ybar[227]),
    .I0(abar[14]),
    .I1(bbar[3])
  );
  //AND U116
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U116 (
    .O(y[226]),
    .I0(a[14]),
    .I1(b[2])
  );
  //OR U116bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U116bar (
    .O(ybar[226]),
    .I0(abar[14]),
    .I1(bbar[2])
  );
  //AND U117
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U117 (
    .O(y[225]),
    .I0(a[14]),
    .I1(b[1])
  );
  //OR U117bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U117bar (
    .O(ybar[225]),
    .I0(abar[14]),
    .I1(bbar[1])
  );
  //AND U118
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U118 (
    .O(y[224]),
    .I0(a[14]),
    .I1(b[0])
  );
  //OR U118bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U118bar (
    .O(ybar[224]),
    .I0(abar[14]),
    .I1(bbar[0])
  );
  //AND U119
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U119 (
    .O(y[223]),
    .I0(a[13]),
    .I1(b[15])
  );
  //OR U119bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U119bar (
    .O(ybar[223]),
    .I0(abar[13]),
    .I1(bbar[15])
  );
  //AND U120
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U120 (
    .O(y[222]),
    .I0(a[13]),
    .I1(b[14])
  );
  //OR U120bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U120bar (
    .O(ybar[222]),
    .I0(abar[13]),
    .I1(bbar[14])
  );
  //AND U121
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U121 (
    .O(y[221]),
    .I0(a[13]),
    .I1(b[13])
  );
  //OR U121bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U121bar (
    .O(ybar[221]),
    .I0(abar[13]),
    .I1(bbar[13])
  );
  //AND U122
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U122 (
    .O(y[220]),
    .I0(a[13]),
    .I1(b[12])
  );
  //OR U122bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U122bar (
    .O(ybar[220]),
    .I0(abar[13]),
    .I1(bbar[12])
  );
  //AND U123
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U123 (
    .O(y[21]),
    .I0(a[1]),
    .I1(b[5])
  );
  //OR U123bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U123bar (
    .O(ybar[21]),
    .I0(abar[1]),
    .I1(bbar[5])
  );
  //AND U124
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U124 (
    .O(y[219]),
    .I0(a[13]),
    .I1(b[11])
  );
  //OR U124bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U124bar (
    .O(ybar[219]),
    .I0(abar[13]),
    .I1(bbar[11])
  );
  //AND U125
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U125 (
    .O(y[218]),
    .I0(a[13]),
    .I1(b[10])
  );
  //OR U125bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U125bar (
    .O(ybar[218]),
    .I0(abar[13]),
    .I1(bbar[10])
  );
  //AND U126
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U126 (
    .O(y[217]),
    .I0(a[13]),
    .I1(b[9])
  );
  //OR U126bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U126bar (
    .O(ybar[217]),
    .I0(abar[13]),
    .I1(bbar[9])
  );
  //AND U127
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U127 (
    .O(y[216]),
    .I0(a[13]),
    .I1(b[8])
  );
  //OR U127bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U127bar (
    .O(ybar[216]),
    .I0(abar[13]),
    .I1(bbar[8])
  );
  //AND U128
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U128 (
    .O(y[215]),
    .I0(a[13]),
    .I1(b[7])
  );
  //OR U128bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U128bar (
    .O(ybar[215]),
    .I0(abar[13]),
    .I1(bbar[7])
  );
  //AND U129
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U129 (
    .O(y[214]),
    .I0(a[13]),
    .I1(b[6])
  );
  //OR U129bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U129bar (
    .O(ybar[214]),
    .I0(abar[13]),
    .I1(bbar[6])
  );
  //AND U130
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U130 (
    .O(y[213]),
    .I0(a[13]),
    .I1(b[5])
  );
  //OR U130bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U130bar (
    .O(ybar[213]),
    .I0(abar[13]),
    .I1(bbar[5])
  );
  //AND U131
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U131 (
    .O(y[212]),
    .I0(a[13]),
    .I1(b[4])
  );
  //OR U131bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U131bar (
    .O(ybar[212]),
    .I0(abar[13]),
    .I1(bbar[4])
  );
  //AND U132
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U132 (
    .O(y[211]),
    .I0(a[13]),
    .I1(b[3])
  );
  //OR U132bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U132bar (
    .O(ybar[211]),
    .I0(abar[13]),
    .I1(bbar[3])
  );
  //AND U133
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U133 (
    .O(y[210]),
    .I0(a[13]),
    .I1(b[2])
  );
  //OR U133bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U133bar (
    .O(ybar[210]),
    .I0(abar[13]),
    .I1(bbar[2])
  );
  //AND U134
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U134 (
    .O(y[20]),
    .I0(a[1]),
    .I1(b[4])
  );
  //OR U134bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U134bar (
    .O(ybar[20]),
    .I0(abar[1]),
    .I1(bbar[4])
  );
  //AND U135
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U135 (
    .O(y[209]),
    .I0(a[13]),
    .I1(b[1])
  );
  //OR U135bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U135bar (
    .O(ybar[209]),
    .I0(abar[13]),
    .I1(bbar[1])
  );
  //AND U136
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U136 (
    .O(y[208]),
    .I0(a[13]),
    .I1(b[0])
  );
  //OR U136bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U136bar (
    .O(ybar[208]),
    .I0(abar[13]),
    .I1(bbar[0])
  );
  //AND U137
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U137 (
    .O(y[207]),
    .I0(a[12]),
    .I1(b[15])
  );
  //OR U137bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U137bar (
    .O(ybar[207]),
    .I0(abar[12]),
    .I1(bbar[15])
  );
  //AND U138
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U138 (
    .O(y[206]),
    .I0(a[12]),
    .I1(b[14])
  );
  //OR U138bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U138bar (
    .O(ybar[206]),
    .I0(abar[12]),
    .I1(bbar[14])
  );
  //AND U139
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U139 (
    .O(y[205]),
    .I0(a[12]),
    .I1(b[13])
  );
  //OR U139bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U139bar (
    .O(ybar[205]),
    .I0(abar[12]),
    .I1(bbar[13])
  );
  //AND U140
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U140 (
    .O(y[204]),
    .I0(a[12]),
    .I1(b[12])
  );
  //OR U140bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U140bar (
    .O(ybar[204]),
    .I0(abar[12]),
    .I1(bbar[12])
  );
  //AND U141
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U141 (
    .O(y[203]),
    .I0(a[12]),
    .I1(b[11])
  );
  //OR U141bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U141bar (
    .O(ybar[203]),
    .I0(abar[12]),
    .I1(bbar[11])
  );
  //AND U142
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U142 (
    .O(y[202]),
    .I0(a[12]),
    .I1(b[10])
  );
  //OR U142bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U142bar (
    .O(ybar[202]),
    .I0(abar[12]),
    .I1(bbar[10])
  );
  //AND U143
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U143 (
    .O(y[201]),
    .I0(a[12]),
    .I1(b[9])
  );
  //OR U143bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U143bar (
    .O(ybar[201]),
    .I0(abar[12]),
    .I1(bbar[9])
  );
  //AND U144
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U144 (
    .O(y[200]),
    .I0(a[12]),
    .I1(b[8])
  );
  //OR U144bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U144bar (
    .O(ybar[200]),
    .I0(abar[12]),
    .I1(bbar[8])
  );
  //AND U145
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U145 (
    .O(y[1]),
    .I0(b[1]),
    .I1(a[0])
  );
  //OR U145bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U145bar (
    .O(ybar[1]),
    .I0(bbar[1]),
    .I1(abar[0])
  );
  //AND U146
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U146 (
    .O(y[19]),
    .I0(a[1]),
    .I1(b[3])
  );
  //OR U146bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U146bar (
    .O(ybar[19]),
    .I0(abar[1]),
    .I1(bbar[3])
  );
  //AND U147
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U147 (
    .O(y[199]),
    .I0(a[12]),
    .I1(b[7])
  );
  //OR U147bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U147bar (
    .O(ybar[199]),
    .I0(abar[12]),
    .I1(bbar[7])
  );
  //AND U148
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U148 (
    .O(y[198]),
    .I0(a[12]),
    .I1(b[6])
  );
  //OR U148bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U148bar (
    .O(ybar[198]),
    .I0(abar[12]),
    .I1(bbar[6])
  );
  //AND U149
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U149 (
    .O(y[197]),
    .I0(a[12]),
    .I1(b[5])
  );
  //OR U149bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U149bar (
    .O(ybar[197]),
    .I0(abar[12]),
    .I1(bbar[5])
  );
  //AND U150
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U150 (
    .O(y[196]),
    .I0(a[12]),
    .I1(b[4])
  );
  //OR U150bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U150bar (
    .O(ybar[196]),
    .I0(abar[12]),
    .I1(bbar[4])
  );
  //AND U151
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U151 (
    .O(y[195]),
    .I0(a[12]),
    .I1(b[3])
  );
  //OR U151bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U151bar (
    .O(ybar[195]),
    .I0(abar[12]),
    .I1(bbar[3])
  );
  //AND U152
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U152 (
    .O(y[194]),
    .I0(a[12]),
    .I1(b[2])
  );
  //OR U152bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U152bar (
    .O(ybar[194]),
    .I0(abar[12]),
    .I1(bbar[2])
  );
  //AND U153
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U153 (
    .O(y[193]),
    .I0(a[12]),
    .I1(b[1])
  );
  //OR U153bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U153bar (
    .O(ybar[193]),
    .I0(abar[12]),
    .I1(bbar[1])
  );
  //AND U154
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U154 (
    .O(y[192]),
    .I0(a[12]),
    .I1(b[0])
  );
  //OR U154bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U154bar (
    .O(ybar[192]),
    .I0(abar[12]),
    .I1(bbar[0])
  );
  //AND U155
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U155 (
    .O(y[191]),
    .I0(a[11]),
    .I1(b[15])
  );
  //OR U155bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U155bar (
    .O(ybar[191]),
    .I0(abar[11]),
    .I1(bbar[15])
  );
  //AND U156
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U156 (
    .O(y[190]),
    .I0(a[11]),
    .I1(b[14])
  );
  //OR U156bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U156bar (
    .O(ybar[190]),
    .I0(abar[11]),
    .I1(bbar[14])
  );
  //AND U157
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U157 (
    .O(y[18]),
    .I0(a[1]),
    .I1(b[2])
  );
  //OR U157bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U157bar (
    .O(ybar[18]),
    .I0(abar[1]),
    .I1(bbar[2])
  );
  //AND U158
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U158 (
    .O(y[189]),
    .I0(a[11]),
    .I1(b[13])
  );
  //OR U158bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U158bar (
    .O(ybar[189]),
    .I0(abar[11]),
    .I1(bbar[13])
  );
  //AND U159
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U159 (
    .O(y[188]),
    .I0(a[11]),
    .I1(b[12])
  );
  //OR U159bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U159bar (
    .O(ybar[188]),
    .I0(abar[11]),
    .I1(bbar[12])
  );
  //AND U160
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U160 (
    .O(y[187]),
    .I0(a[11]),
    .I1(b[11])
  );
  //OR U160bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U160bar (
    .O(ybar[187]),
    .I0(abar[11]),
    .I1(bbar[11])
  );
  //AND U161
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U161 (
    .O(y[186]),
    .I0(a[11]),
    .I1(b[10])
  );
  //OR U161bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U161bar (
    .O(ybar[186]),
    .I0(abar[11]),
    .I1(bbar[10])
  );
  //AND U162
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U162 (
    .O(y[185]),
    .I0(a[11]),
    .I1(b[9])
  );
  //OR U162bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U162bar (
    .O(ybar[185]),
    .I0(abar[11]),
    .I1(bbar[9])
  );
  //AND U163
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U163 (
    .O(y[184]),
    .I0(a[11]),
    .I1(b[8])
  );
  //OR U163bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U163bar (
    .O(ybar[184]),
    .I0(abar[11]),
    .I1(bbar[8])
  );
  //AND U164
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U164 (
    .O(y[183]),
    .I0(a[11]),
    .I1(b[7])
  );
  //OR U164bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U164bar (
    .O(ybar[183]),
    .I0(abar[11]),
    .I1(bbar[7])
  );
  //AND U165
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U165 (
    .O(y[182]),
    .I0(a[11]),
    .I1(b[6])
  );
  //OR U165bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U165bar (
    .O(ybar[182]),
    .I0(abar[11]),
    .I1(bbar[6])
  );
  //AND U166
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U166 (
    .O(y[181]),
    .I0(a[11]),
    .I1(b[5])
  );
  //OR U166bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U166bar (
    .O(ybar[181]),
    .I0(abar[11]),
    .I1(bbar[5])
  );
  //AND U167
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U167 (
    .O(y[180]),
    .I0(a[11]),
    .I1(b[4])
  );
  //OR U167bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U167bar (
    .O(ybar[180]),
    .I0(abar[11]),
    .I1(bbar[4])
  );
  //AND U168
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U168 (
    .O(y[17]),
    .I0(a[1]),
    .I1(b[1])
  );
  //OR U168bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U168bar (
    .O(ybar[17]),
    .I0(abar[1]),
    .I1(bbar[1])
  );
  //AND U169
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U169 (
    .O(y[179]),
    .I0(a[11]),
    .I1(b[3])
  );
  //OR U169bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U169bar (
    .O(ybar[179]),
    .I0(abar[11]),
    .I1(bbar[3])
  );
  //AND U170
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U170 (
    .O(y[178]),
    .I0(a[11]),
    .I1(b[2])
  );
  //OR U170bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U170bar (
    .O(ybar[178]),
    .I0(abar[11]),
    .I1(bbar[2])
  );
  //AND U171
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U171 (
    .O(y[177]),
    .I0(a[11]),
    .I1(b[1])
  );
  //OR U171bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U171bar (
    .O(ybar[177]),
    .I0(abar[11]),
    .I1(bbar[1])
  );
  //AND U172
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U172 (
    .O(y[176]),
    .I0(a[11]),
    .I1(b[0])
  );
  //OR U172bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U172bar (
    .O(ybar[176]),
    .I0(abar[11]),
    .I1(bbar[0])
  );
  //AND U173
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U173 (
    .O(y[175]),
    .I0(a[10]),
    .I1(b[15])
  );
  //OR U173bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U173bar (
    .O(ybar[175]),
    .I0(abar[10]),
    .I1(bbar[15])
  );
  //AND U174
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U174 (
    .O(y[174]),
    .I0(a[10]),
    .I1(b[14])
  );
  //OR U174bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U174bar (
    .O(ybar[174]),
    .I0(abar[10]),
    .I1(bbar[14])
  );
  //AND U175
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U175 (
    .O(y[173]),
    .I0(a[10]),
    .I1(b[13])
  );
  //OR U175bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U175bar (
    .O(ybar[173]),
    .I0(abar[10]),
    .I1(bbar[13])
  );
  //AND U176
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U176 (
    .O(y[172]),
    .I0(a[10]),
    .I1(b[12])
  );
  //OR U176bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U176bar (
    .O(ybar[172]),
    .I0(abar[10]),
    .I1(bbar[12])
  );
  //AND U177
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U177 (
    .O(y[171]),
    .I0(a[10]),
    .I1(b[11])
  );
  //OR U177bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U177bar (
    .O(ybar[171]),
    .I0(abar[10]),
    .I1(bbar[11])
  );
  //AND U178
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U178 (
    .O(y[170]),
    .I0(a[10]),
    .I1(b[10])
  );
  //OR U178bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U178bar (
    .O(ybar[170]),
    .I0(abar[10]),
    .I1(bbar[10])
  );
  //AND U179
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U179 (
    .O(y[16]),
    .I0(a[1]),
    .I1(b[0])
  );
  //OR U179bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U179bar (
    .O(ybar[16]),
    .I0(abar[1]),
    .I1(bbar[0])
  );
  //AND U180
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U180 (
    .O(y[169]),
    .I0(a[10]),
    .I1(b[9])
  );
  //OR U180bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U180bar (
    .O(ybar[169]),
    .I0(abar[10]),
    .I1(bbar[9])
  );
  //AND U181
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U181 (
    .O(y[168]),
    .I0(a[10]),
    .I1(b[8])
  );
  //OR U181bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U181bar (
    .O(ybar[168]),
    .I0(abar[10]),
    .I1(bbar[8])
  );
  //AND U182
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U182 (
    .O(y[167]),
    .I0(a[10]),
    .I1(b[7])
  );
  //OR U182bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U182bar (
    .O(ybar[167]),
    .I0(abar[10]),
    .I1(bbar[7])
  );
  //AND U183
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U183 (
    .O(y[166]),
    .I0(a[10]),
    .I1(b[6])
  );
  //OR U183bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U183bar (
    .O(ybar[166]),
    .I0(abar[10]),
    .I1(bbar[6])
  );
  //AND U184
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U184 (
    .O(y[165]),
    .I0(a[10]),
    .I1(b[5])
  );
  //OR U184bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U184bar (
    .O(ybar[165]),
    .I0(abar[10]),
    .I1(bbar[5])
  );
  //AND U185
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U185 (
    .O(y[164]),
    .I0(a[10]),
    .I1(b[4])
  );
  //OR U185bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U185bar (
    .O(ybar[164]),
    .I0(abar[10]),
    .I1(bbar[4])
  );
  //AND U186
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U186 (
    .O(y[163]),
    .I0(a[10]),
    .I1(b[3])
  );
  //OR U186bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U186bar (
    .O(ybar[163]),
    .I0(abar[10]),
    .I1(bbar[3])
  );
  //AND U187
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U187 (
    .O(y[162]),
    .I0(a[10]),
    .I1(b[2])
  );
  //OR U187bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U187bar (
    .O(ybar[162]),
    .I0(abar[10]),
    .I1(bbar[2])
  );
  //AND U188
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U188 (
    .O(y[161]),
    .I0(a[10]),
    .I1(b[1])
  );
  //OR U188bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U188bar (
    .O(ybar[161]),
    .I0(abar[10]),
    .I1(bbar[1])
  );
  //AND U189
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U189 (
    .O(y[160]),
    .I0(a[10]),
    .I1(b[0])
  );
  //OR U189bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U189bar (
    .O(ybar[160]),
    .I0(abar[10]),
    .I1(bbar[0])
  );
  //AND U190
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U190 (
    .O(y[15]),
    .I0(b[15]),
    .I1(a[0])
  );
  //OR U190bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U190bar (
    .O(ybar[15]),
    .I0(bbar[15]),
    .I1(abar[0])
  );
  //AND U191
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U191 (
    .O(y[159]),
    .I0(a[9]),
    .I1(b[15])
  );
  //OR U191bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U191bar (
    .O(ybar[159]),
    .I0(abar[9]),
    .I1(bbar[15])
  );
  //AND U192
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U192 (
    .O(y[158]),
    .I0(a[9]),
    .I1(b[14])
  );
  //OR U192bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U192bar (
    .O(ybar[158]),
    .I0(abar[9]),
    .I1(bbar[14])
  );
  //AND U193
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U193 (
    .O(y[157]),
    .I0(a[9]),
    .I1(b[13])
  );
  //OR U193bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U193bar (
    .O(ybar[157]),
    .I0(abar[9]),
    .I1(bbar[13])
  );
  //AND U194
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U194 (
    .O(y[156]),
    .I0(a[9]),
    .I1(b[12])
  );
  //OR U194bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U194bar (
    .O(ybar[156]),
    .I0(abar[9]),
    .I1(bbar[12])
  );
  //AND U195
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U195 (
    .O(y[155]),
    .I0(a[9]),
    .I1(b[11])
  );
  //OR U195bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U195bar (
    .O(ybar[155]),
    .I0(abar[9]),
    .I1(bbar[11])
  );
  //AND U196
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U196 (
    .O(y[154]),
    .I0(a[9]),
    .I1(b[10])
  );
  //OR U196bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U196bar (
    .O(ybar[154]),
    .I0(abar[9]),
    .I1(bbar[10])
  );
  //AND U197
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U197 (
    .O(y[153]),
    .I0(a[9]),
    .I1(b[9])
  );
  //OR U197bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U197bar (
    .O(ybar[153]),
    .I0(abar[9]),
    .I1(bbar[9])
  );
  //AND U198
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U198 (
    .O(y[152]),
    .I0(a[9]),
    .I1(b[8])
  );
  //OR U198bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U198bar (
    .O(ybar[152]),
    .I0(abar[9]),
    .I1(bbar[8])
  );
  //AND U199
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U199 (
    .O(y[151]),
    .I0(a[9]),
    .I1(b[7])
  );
  //OR U199bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U199bar (
    .O(ybar[151]),
    .I0(abar[9]),
    .I1(bbar[7])
  );
  //AND U200
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U200 (
    .O(y[150]),
    .I0(a[9]),
    .I1(b[6])
  );
  //OR U200bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U200bar (
    .O(ybar[150]),
    .I0(abar[9]),
    .I1(bbar[6])
  );
  //AND U201
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U201 (
    .O(y[14]),
    .I0(b[14]),
    .I1(a[0])
  );
  //OR U201bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U201bar (
    .O(ybar[14]),
    .I0(bbar[14]),
    .I1(abar[0])
  );
  //AND U202
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U202 (
    .O(y[149]),
    .I0(a[9]),
    .I1(b[5])
  );
  //OR U202bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U202bar (
    .O(ybar[149]),
    .I0(abar[9]),
    .I1(bbar[5])
  );
  //AND U203
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U203 (
    .O(y[148]),
    .I0(a[9]),
    .I1(b[4])
  );
  //OR U203bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U203bar (
    .O(ybar[148]),
    .I0(abar[9]),
    .I1(bbar[4])
  );
  //AND U204
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U204 (
    .O(y[147]),
    .I0(a[9]),
    .I1(b[3])
  );
  //OR U204bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U204bar (
    .O(ybar[147]),
    .I0(abar[9]),
    .I1(bbar[3])
  );
  //AND U205
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U205 (
    .O(y[146]),
    .I0(a[9]),
    .I1(b[2])
  );
  //OR U205bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U205bar (
    .O(ybar[146]),
    .I0(abar[9]),
    .I1(bbar[2])
  );
  //AND U206
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U206 (
    .O(y[145]),
    .I0(a[9]),
    .I1(b[1])
  );
  //OR U206bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U206bar (
    .O(ybar[145]),
    .I0(abar[9]),
    .I1(bbar[1])
  );
  //AND U207
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U207 (
    .O(y[144]),
    .I0(a[9]),
    .I1(b[0])
  );
  //OR U207bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U207bar (
    .O(ybar[144]),
    .I0(abar[9]),
    .I1(bbar[0])
  );
  //AND U208
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U208 (
    .O(y[143]),
    .I0(a[8]),
    .I1(b[15])
  );
  //OR U208bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U208bar (
    .O(ybar[143]),
    .I0(abar[8]),
    .I1(bbar[15])
  );
  //AND U209
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U209 (
    .O(y[142]),
    .I0(a[8]),
    .I1(b[14])
  );
  //OR U209bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U209bar (
    .O(ybar[142]),
    .I0(abar[8]),
    .I1(bbar[14])
  );
  //AND U210
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U210 (
    .O(y[141]),
    .I0(a[8]),
    .I1(b[13])
  );
  //OR U210bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U210bar (
    .O(ybar[141]),
    .I0(abar[8]),
    .I1(bbar[13])
  );
  //AND U211
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U211 (
    .O(y[140]),
    .I0(a[8]),
    .I1(b[12])
  );
  //OR U211bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U211bar (
    .O(ybar[140]),
    .I0(abar[8]),
    .I1(bbar[12])
  );
  //AND U212
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U212 (
    .O(y[13]),
    .I0(b[13]),
    .I1(a[0])
  );
  //OR U212bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U212bar (
    .O(ybar[13]),
    .I0(bbar[13]),
    .I1(abar[0])
  );
  //AND U213
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U213 (
    .O(y[139]),
    .I0(a[8]),
    .I1(b[11])
  );
  //OR U213bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U213bar (
    .O(ybar[139]),
    .I0(abar[8]),
    .I1(bbar[11])
  );
  //AND U214
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U214 (
    .O(y[138]),
    .I0(a[8]),
    .I1(b[10])
  );
  //OR U214bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U214bar (
    .O(ybar[138]),
    .I0(abar[8]),
    .I1(bbar[10])
  );
  //AND U215
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U215 (
    .O(y[137]),
    .I0(a[8]),
    .I1(b[9])
  );
  //OR U215bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U215bar (
    .O(ybar[137]),
    .I0(abar[8]),
    .I1(bbar[9])
  );
  //AND U216
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U216 (
    .O(y[136]),
    .I0(a[8]),
    .I1(b[8])
  );
  //OR U216bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U216bar (
    .O(ybar[136]),
    .I0(abar[8]),
    .I1(bbar[8])
  );
  //AND U217
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U217 (
    .O(y[135]),
    .I0(a[8]),
    .I1(b[7])
  );
  //OR U217bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U217bar (
    .O(ybar[135]),
    .I0(abar[8]),
    .I1(bbar[7])
  );
  //AND U218
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U218 (
    .O(y[134]),
    .I0(a[8]),
    .I1(b[6])
  );
  //OR U218bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U218bar (
    .O(ybar[134]),
    .I0(abar[8]),
    .I1(bbar[6])
  );
  //AND U219
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U219 (
    .O(y[133]),
    .I0(a[8]),
    .I1(b[5])
  );
  //OR U219bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U219bar (
    .O(ybar[133]),
    .I0(abar[8]),
    .I1(bbar[5])
  );
  //AND U220
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U220 (
    .O(y[132]),
    .I0(a[8]),
    .I1(b[4])
  );
  //OR U220bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U220bar (
    .O(ybar[132]),
    .I0(abar[8]),
    .I1(bbar[4])
  );
  //AND U221
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U221 (
    .O(y[131]),
    .I0(a[8]),
    .I1(b[3])
  );
  //OR U221bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U221bar (
    .O(ybar[131]),
    .I0(abar[8]),
    .I1(bbar[3])
  );
  //AND U222
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U222 (
    .O(y[130]),
    .I0(a[8]),
    .I1(b[2])
  );
  //OR U222bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U222bar (
    .O(ybar[130]),
    .I0(abar[8]),
    .I1(bbar[2])
  );
  //AND U223
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U223 (
    .O(y[12]),
    .I0(b[12]),
    .I1(a[0])
  );
  //OR U223bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U223bar (
    .O(ybar[12]),
    .I0(bbar[12]),
    .I1(abar[0])
  );
  //AND U224
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U224 (
    .O(y[129]),
    .I0(a[8]),
    .I1(b[1])
  );
  //OR U224bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U224bar (
    .O(ybar[129]),
    .I0(abar[8]),
    .I1(bbar[1])
  );
  //AND U225
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U225 (
    .O(y[128]),
    .I0(a[8]),
    .I1(b[0])
  );
  //OR U225bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U225bar (
    .O(ybar[128]),
    .I0(abar[8]),
    .I1(bbar[0])
  );
  //AND U226
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U226 (
    .O(y[127]),
    .I0(a[7]),
    .I1(b[15])
  );
  //OR U226bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U226bar (
    .O(ybar[127]),
    .I0(abar[7]),
    .I1(bbar[15])
  );
  //AND U227
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U227 (
    .O(y[126]),
    .I0(a[7]),
    .I1(b[14])
  );
  //OR U227bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U227bar (
    .O(ybar[126]),
    .I0(abar[7]),
    .I1(bbar[14])
  );
  //AND U228
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U228 (
    .O(y[125]),
    .I0(a[7]),
    .I1(b[13])
  );
  //OR U228bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U228bar (
    .O(ybar[125]),
    .I0(abar[7]),
    .I1(bbar[13])
  );
  //AND U229
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U229 (
    .O(y[124]),
    .I0(a[7]),
    .I1(b[12])
  );
  //OR U229bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U229bar (
    .O(ybar[124]),
    .I0(abar[7]),
    .I1(bbar[12])
  );
  //AND U230
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U230 (
    .O(y[123]),
    .I0(a[7]),
    .I1(b[11])
  );
  //OR U230bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U230bar (
    .O(ybar[123]),
    .I0(abar[7]),
    .I1(bbar[11])
  );
  //AND U231
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U231 (
    .O(y[122]),
    .I0(a[7]),
    .I1(b[10])
  );
  //OR U231bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U231bar (
    .O(ybar[122]),
    .I0(abar[7]),
    .I1(bbar[10])
  );
  //AND U232
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U232 (
    .O(y[121]),
    .I0(a[7]),
    .I1(b[9])
  );
  //OR U232bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U232bar (
    .O(ybar[121]),
    .I0(abar[7]),
    .I1(bbar[9])
  );
  //AND U233
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U233 (
    .O(y[120]),
    .I0(a[7]),
    .I1(b[8])
  );
  //OR U233bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U233bar (
    .O(ybar[120]),
    .I0(abar[7]),
    .I1(bbar[8])
  );
  //AND U234
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U234 (
    .O(y[11]),
    .I0(b[11]),
    .I1(a[0])
  );
  //OR U234bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U234bar (
    .O(ybar[11]),
    .I0(bbar[11]),
    .I1(abar[0])
  );
  //AND U235
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U235 (
    .O(y[119]),
    .I0(a[7]),
    .I1(b[7])
  );
  //OR U235bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U235bar (
    .O(ybar[119]),
    .I0(abar[7]),
    .I1(bbar[7])
  );
  //AND U236
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U236 (
    .O(y[118]),
    .I0(a[7]),
    .I1(b[6])
  );
  //OR U236bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U236bar (
    .O(ybar[118]),
    .I0(abar[7]),
    .I1(bbar[6])
  );
  //AND U237
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U237 (
    .O(y[117]),
    .I0(a[7]),
    .I1(b[5])
  );
  //OR U237bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U237bar (
    .O(ybar[117]),
    .I0(abar[7]),
    .I1(bbar[5])
  );
  //AND U238
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U238 (
    .O(y[116]),
    .I0(a[7]),
    .I1(b[4])
  );
  //OR U238bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U238bar (
    .O(ybar[116]),
    .I0(abar[7]),
    .I1(bbar[4])
  );
  //AND U239
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U239 (
    .O(y[115]),
    .I0(a[7]),
    .I1(b[3])
  );
  //OR U239bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U239bar (
    .O(ybar[115]),
    .I0(abar[7]),
    .I1(bbar[3])
  );
  //AND U240
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U240 (
    .O(y[114]),
    .I0(a[7]),
    .I1(b[2])
  );
  //OR U240bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U240bar (
    .O(ybar[114]),
    .I0(abar[7]),
    .I1(bbar[2])
  );
  //AND U241
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U241 (
    .O(y[113]),
    .I0(a[7]),
    .I1(b[1])
  );
  //OR U241bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U241bar (
    .O(ybar[113]),
    .I0(abar[7]),
    .I1(bbar[1])
  );
  //AND U242
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U242 (
    .O(y[112]),
    .I0(a[7]),
    .I1(b[0])
  );
  //OR U242bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U242bar (
    .O(ybar[112]),
    .I0(abar[7]),
    .I1(bbar[0])
  );
  //AND U243
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U243 (
    .O(y[111]),
    .I0(b[15]),
    .I1(a[6])
  );
  //OR U243bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U243bar (
    .O(ybar[111]),
    .I0(bbar[15]),
    .I1(abar[6])
  );
  //AND U244
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U244 (
    .O(y[110]),
    .I0(b[14]),
    .I1(a[6])
  );
  //OR U244bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U244bar (
    .O(ybar[110]),
    .I0(bbar[14]),
    .I1(abar[6])
  );
  //AND U245
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U245 (
    .O(y[10]),
    .I0(b[10]),
    .I1(a[0])
  );
  //OR U245bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U245bar (
    .O(ybar[10]),
    .I0(bbar[10]),
    .I1(abar[0])
  );
  //AND U246
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U246 (
    .O(y[109]),
    .I0(b[13]),
    .I1(a[6])
  );
  //OR U246bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U246bar (
    .O(ybar[109]),
    .I0(bbar[13]),
    .I1(abar[6])
  );
  //AND U247
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U247 (
    .O(y[108]),
    .I0(b[12]),
    .I1(a[6])
  );
  //OR U247bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U247bar (
    .O(ybar[108]),
    .I0(bbar[12]),
    .I1(abar[6])
  );
  //AND U248
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U248 (
    .O(y[107]),
    .I0(b[11]),
    .I1(a[6])
  );
  //OR U248bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U248bar (
    .O(ybar[107]),
    .I0(bbar[11]),
    .I1(abar[6])
  );
  //AND U249
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U249 (
    .O(y[106]),
    .I0(b[10]),
    .I1(a[6])
  );
  //OR U249bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U249bar (
    .O(ybar[106]),
    .I0(bbar[10]),
    .I1(abar[6])
  );
  //AND U250
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U250 (
    .O(y[105]),
    .I0(a[6]),
    .I1(b[9])
  );
  //OR U250bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U250bar (
    .O(ybar[105]),
    .I0(abar[6]),
    .I1(bbar[9])
  );
  //AND U251
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U251 (
    .O(y[104]),
    .I0(b[8]),
    .I1(a[6])
  );
  //OR U251bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U251bar (
    .O(ybar[104]),
    .I0(bbar[8]),
    .I1(abar[6])
  );
  //AND U252
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U252 (
    .O(y[103]),
    .I0(b[7]),
    .I1(a[6])
  );
  //OR U252bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U252bar (
    .O(ybar[103]),
    .I0(bbar[7]),
    .I1(abar[6])
  );
  //AND U253
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U253 (
    .O(y[102]),
    .I0(b[6]),
    .I1(a[6])
  );
  //OR U253bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U253bar (
    .O(ybar[102]),
    .I0(bbar[6]),
    .I1(abar[6])
  );
  //AND U254
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U254 (
    .O(y[101]),
    .I0(b[5]),
    .I1(a[6])
  );
  //OR U254bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U254bar (
    .O(ybar[101]),
    .I0(bbar[5]),
    .I1(abar[6])
  );
  //AND U255
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U255 (
    .O(y[100]),
    .I0(b[4]),
    .I1(a[6])
  );
  //OR U255bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U255bar (
    .O(ybar[100]),
    .I0(bbar[4]),
    .I1(abar[6])
  );
  //AND U256
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U256 (
    .O(y[0]),
    .I0(b[0]),
    .I1(a[0])
  );
  //OR U256bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U256bar (
    .O(ybar[0]),
    .I0(bbar[0]),
    .I1(abar[0])
  );
endmodule

module decode_4 ( in, out );

  input wire [7:0] in;
//input_done

  output wire [255:0] out;
//output_done

  wire [15:0] level1;
  wire [31:0] level2;
//wire_done

  CD2_16 cd_l1_1 ( .a(in[1]), .b(in[0]), .y(level1[3:0]) );
  CD2_15 cd_l1_2 ( .a(in[3]), .b(in[2]), .y(level1[7:4]) );
  CD2_14 cd_l1_3 ( .a(in[5]), .b(in[4]), .y(level1[11:8]) );
  CD2_13 cd_l1_4 ( .a(in[7]), .b(in[6]), .y(level1[15:12]) );
  CD4_8 cd_l2_1 ( .a(level1[7:4]), .b(level1[3:0]), .y(level2[15:0]) );
  CD4_7 cd_l2_2 ( .a(level1[15:12]), .b(level1[11:8]), .y(level2[31:16]) );
  CD16_4 cd_l3 ( .a(level2[31:16]), .b(level2[15:0]), .y(out) );
endmodule

module encode_4 ( in, out );

  input wire [255:0] in;
  wire [255:0] inbar;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
  assign inbar[8] = ~in[8];
  assign inbar[9] = ~in[9];
  assign inbar[10] = ~in[10];
  assign inbar[11] = ~in[11];
  assign inbar[12] = ~in[12];
  assign inbar[13] = ~in[13];
  assign inbar[14] = ~in[14];
  assign inbar[15] = ~in[15];
  assign inbar[16] = ~in[16];
  assign inbar[17] = ~in[17];
  assign inbar[18] = ~in[18];
  assign inbar[19] = ~in[19];
  assign inbar[20] = ~in[20];
  assign inbar[21] = ~in[21];
  assign inbar[22] = ~in[22];
  assign inbar[23] = ~in[23];
  assign inbar[24] = ~in[24];
  assign inbar[25] = ~in[25];
  assign inbar[26] = ~in[26];
  assign inbar[27] = ~in[27];
  assign inbar[28] = ~in[28];
  assign inbar[29] = ~in[29];
  assign inbar[30] = ~in[30];
  assign inbar[31] = ~in[31];
  assign inbar[32] = ~in[32];
  assign inbar[33] = ~in[33];
  assign inbar[34] = ~in[34];
  assign inbar[35] = ~in[35];
  assign inbar[36] = ~in[36];
  assign inbar[37] = ~in[37];
  assign inbar[38] = ~in[38];
  assign inbar[39] = ~in[39];
  assign inbar[40] = ~in[40];
  assign inbar[41] = ~in[41];
  assign inbar[42] = ~in[42];
  assign inbar[43] = ~in[43];
  assign inbar[44] = ~in[44];
  assign inbar[45] = ~in[45];
  assign inbar[46] = ~in[46];
  assign inbar[47] = ~in[47];
  assign inbar[48] = ~in[48];
  assign inbar[49] = ~in[49];
  assign inbar[50] = ~in[50];
  assign inbar[51] = ~in[51];
  assign inbar[52] = ~in[52];
  assign inbar[53] = ~in[53];
  assign inbar[54] = ~in[54];
  assign inbar[55] = ~in[55];
  assign inbar[56] = ~in[56];
  assign inbar[57] = ~in[57];
  assign inbar[58] = ~in[58];
  assign inbar[59] = ~in[59];
  assign inbar[60] = ~in[60];
  assign inbar[61] = ~in[61];
  assign inbar[62] = ~in[62];
  assign inbar[63] = ~in[63];
  assign inbar[64] = ~in[64];
  assign inbar[65] = ~in[65];
  assign inbar[66] = ~in[66];
  assign inbar[67] = ~in[67];
  assign inbar[68] = ~in[68];
  assign inbar[69] = ~in[69];
  assign inbar[70] = ~in[70];
  assign inbar[71] = ~in[71];
  assign inbar[72] = ~in[72];
  assign inbar[73] = ~in[73];
  assign inbar[74] = ~in[74];
  assign inbar[75] = ~in[75];
  assign inbar[76] = ~in[76];
  assign inbar[77] = ~in[77];
  assign inbar[78] = ~in[78];
  assign inbar[79] = ~in[79];
  assign inbar[80] = ~in[80];
  assign inbar[81] = ~in[81];
  assign inbar[82] = ~in[82];
  assign inbar[83] = ~in[83];
  assign inbar[84] = ~in[84];
  assign inbar[85] = ~in[85];
  assign inbar[86] = ~in[86];
  assign inbar[87] = ~in[87];
  assign inbar[88] = ~in[88];
  assign inbar[89] = ~in[89];
  assign inbar[90] = ~in[90];
  assign inbar[91] = ~in[91];
  assign inbar[92] = ~in[92];
  assign inbar[93] = ~in[93];
  assign inbar[94] = ~in[94];
  assign inbar[95] = ~in[95];
  assign inbar[96] = ~in[96];
  assign inbar[97] = ~in[97];
  assign inbar[98] = ~in[98];
  assign inbar[99] = ~in[99];
  assign inbar[100] = ~in[100];
  assign inbar[101] = ~in[101];
  assign inbar[102] = ~in[102];
  assign inbar[103] = ~in[103];
  assign inbar[104] = ~in[104];
  assign inbar[105] = ~in[105];
  assign inbar[106] = ~in[106];
  assign inbar[107] = ~in[107];
  assign inbar[108] = ~in[108];
  assign inbar[109] = ~in[109];
  assign inbar[110] = ~in[110];
  assign inbar[111] = ~in[111];
  assign inbar[112] = ~in[112];
  assign inbar[113] = ~in[113];
  assign inbar[114] = ~in[114];
  assign inbar[115] = ~in[115];
  assign inbar[116] = ~in[116];
  assign inbar[117] = ~in[117];
  assign inbar[118] = ~in[118];
  assign inbar[119] = ~in[119];
  assign inbar[120] = ~in[120];
  assign inbar[121] = ~in[121];
  assign inbar[122] = ~in[122];
  assign inbar[123] = ~in[123];
  assign inbar[124] = ~in[124];
  assign inbar[125] = ~in[125];
  assign inbar[126] = ~in[126];
  assign inbar[127] = ~in[127];
  assign inbar[128] = ~in[128];
  assign inbar[129] = ~in[129];
  assign inbar[130] = ~in[130];
  assign inbar[131] = ~in[131];
  assign inbar[132] = ~in[132];
  assign inbar[133] = ~in[133];
  assign inbar[134] = ~in[134];
  assign inbar[135] = ~in[135];
  assign inbar[136] = ~in[136];
  assign inbar[137] = ~in[137];
  assign inbar[138] = ~in[138];
  assign inbar[139] = ~in[139];
  assign inbar[140] = ~in[140];
  assign inbar[141] = ~in[141];
  assign inbar[142] = ~in[142];
  assign inbar[143] = ~in[143];
  assign inbar[144] = ~in[144];
  assign inbar[145] = ~in[145];
  assign inbar[146] = ~in[146];
  assign inbar[147] = ~in[147];
  assign inbar[148] = ~in[148];
  assign inbar[149] = ~in[149];
  assign inbar[150] = ~in[150];
  assign inbar[151] = ~in[151];
  assign inbar[152] = ~in[152];
  assign inbar[153] = ~in[153];
  assign inbar[154] = ~in[154];
  assign inbar[155] = ~in[155];
  assign inbar[156] = ~in[156];
  assign inbar[157] = ~in[157];
  assign inbar[158] = ~in[158];
  assign inbar[159] = ~in[159];
  assign inbar[160] = ~in[160];
  assign inbar[161] = ~in[161];
  assign inbar[162] = ~in[162];
  assign inbar[163] = ~in[163];
  assign inbar[164] = ~in[164];
  assign inbar[165] = ~in[165];
  assign inbar[166] = ~in[166];
  assign inbar[167] = ~in[167];
  assign inbar[168] = ~in[168];
  assign inbar[169] = ~in[169];
  assign inbar[170] = ~in[170];
  assign inbar[171] = ~in[171];
  assign inbar[172] = ~in[172];
  assign inbar[173] = ~in[173];
  assign inbar[174] = ~in[174];
  assign inbar[175] = ~in[175];
  assign inbar[176] = ~in[176];
  assign inbar[177] = ~in[177];
  assign inbar[178] = ~in[178];
  assign inbar[179] = ~in[179];
  assign inbar[180] = ~in[180];
  assign inbar[181] = ~in[181];
  assign inbar[182] = ~in[182];
  assign inbar[183] = ~in[183];
  assign inbar[184] = ~in[184];
  assign inbar[185] = ~in[185];
  assign inbar[186] = ~in[186];
  assign inbar[187] = ~in[187];
  assign inbar[188] = ~in[188];
  assign inbar[189] = ~in[189];
  assign inbar[190] = ~in[190];
  assign inbar[191] = ~in[191];
  assign inbar[192] = ~in[192];
  assign inbar[193] = ~in[193];
  assign inbar[194] = ~in[194];
  assign inbar[195] = ~in[195];
  assign inbar[196] = ~in[196];
  assign inbar[197] = ~in[197];
  assign inbar[198] = ~in[198];
  assign inbar[199] = ~in[199];
  assign inbar[200] = ~in[200];
  assign inbar[201] = ~in[201];
  assign inbar[202] = ~in[202];
  assign inbar[203] = ~in[203];
  assign inbar[204] = ~in[204];
  assign inbar[205] = ~in[205];
  assign inbar[206] = ~in[206];
  assign inbar[207] = ~in[207];
  assign inbar[208] = ~in[208];
  assign inbar[209] = ~in[209];
  assign inbar[210] = ~in[210];
  assign inbar[211] = ~in[211];
  assign inbar[212] = ~in[212];
  assign inbar[213] = ~in[213];
  assign inbar[214] = ~in[214];
  assign inbar[215] = ~in[215];
  assign inbar[216] = ~in[216];
  assign inbar[217] = ~in[217];
  assign inbar[218] = ~in[218];
  assign inbar[219] = ~in[219];
  assign inbar[220] = ~in[220];
  assign inbar[221] = ~in[221];
  assign inbar[222] = ~in[222];
  assign inbar[223] = ~in[223];
  assign inbar[224] = ~in[224];
  assign inbar[225] = ~in[225];
  assign inbar[226] = ~in[226];
  assign inbar[227] = ~in[227];
  assign inbar[228] = ~in[228];
  assign inbar[229] = ~in[229];
  assign inbar[230] = ~in[230];
  assign inbar[231] = ~in[231];
  assign inbar[232] = ~in[232];
  assign inbar[233] = ~in[233];
  assign inbar[234] = ~in[234];
  assign inbar[235] = ~in[235];
  assign inbar[236] = ~in[236];
  assign inbar[237] = ~in[237];
  assign inbar[238] = ~in[238];
  assign inbar[239] = ~in[239];
  assign inbar[240] = ~in[240];
  assign inbar[241] = ~in[241];
  assign inbar[242] = ~in[242];
  assign inbar[243] = ~in[243];
  assign inbar[244] = ~in[244];
  assign inbar[245] = ~in[245];
  assign inbar[246] = ~in[246];
  assign inbar[247] = ~in[247];
  assign inbar[248] = ~in[248];
  assign inbar[249] = ~in[249];
  assign inbar[250] = ~in[250];
  assign inbar[251] = ~in[251];
  assign inbar[252] = ~in[252];
  assign inbar[253] = ~in[253];
  assign inbar[254] = ~in[254];
  assign inbar[255] = ~in[255];
//input_done

  output wire [7:0] out;
  wire [7:0] outbar;
//output_done

  wire in_81;
  wire in_80;
  wire in_79;
  wire in_78;
  wire in_77;
  wire in_76;
  wire in_75;
  wire in_74;
  wire in_73;
  wire in_72;
  wire in_71;
  wire in_70;
  wire in_69;
  wire in_68;
  wire in_67;
  wire in_66;
  wire in_65;
  wire in_64;
  wire in_63;
  wire in_62;
  wire in_61;
  wire in_60;
  wire in_59;
  wire in_58;
  wire in_57;
  wire in_56;
  wire in_55;
  wire in_54;
  wire in_53;
  wire in_52;
  wire in_51;
  wire in_50;
  wire in_49;
  wire in_48;
  wire in_47;
  wire in_46;
  wire in_45;
  wire in_44;
  wire in_43;
  wire in_42;
  wire in_41;
  wire in_40;
  wire in_39;
  wire in_38;
  wire in_37;
  wire in_36;
  wire in_35;
  wire in_34;
  wire in_33;
  wire in_32;
  wire in_31;
  wire in_30;
  wire in_29;
  wire in_28;
  wire in_27;
  wire in_26;
  wire in_25;
  wire in_24;
  wire in_23;
  wire in_22;
  wire in_21;
  wire in_20;
  wire in_19;
  wire in_18;
  wire in_17;
  wire in_16;
  wire in_15;
  wire in_14;
  wire in_13;
  wire in_12;
  wire in_11;
  wire in_10;
  wire in_9;
  wire in_8;
  wire in_7;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_3;
  wire in_2;
  wire in_1;
  wire in_0;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire in_81bar;
  wire in_80bar;
  wire in_79bar;
  wire in_78bar;
  wire in_77bar;
  wire in_76bar;
  wire in_75bar;
  wire in_74bar;
  wire in_73bar;
  wire in_72bar;
  wire in_71bar;
  wire in_70bar;
  wire in_69bar;
  wire in_68bar;
  wire in_67bar;
  wire in_66bar;
  wire in_65bar;
  wire in_64bar;
  wire in_63bar;
  wire in_62bar;
  wire in_61bar;
  wire in_60bar;
  wire in_59bar;
  wire in_58bar;
  wire in_57bar;
  wire in_56bar;
  wire in_55bar;
  wire in_54bar;
  wire in_53bar;
  wire in_52bar;
  wire in_51bar;
  wire in_50bar;
  wire in_49bar;
  wire in_48bar;
  wire in_47bar;
  wire in_46bar;
  wire in_45bar;
  wire in_44bar;
  wire in_43bar;
  wire in_42bar;
  wire in_41bar;
  wire in_40bar;
  wire in_39bar;
  wire in_38bar;
  wire in_37bar;
  wire in_36bar;
  wire in_35bar;
  wire in_34bar;
  wire in_33bar;
  wire in_32bar;
  wire in_31bar;
  wire in_30bar;
  wire in_29bar;
  wire in_28bar;
  wire in_27bar;
  wire in_26bar;
  wire in_25bar;
  wire in_24bar;
  wire in_23bar;
  wire in_22bar;
  wire in_21bar;
  wire in_20bar;
  wire in_19bar;
  wire in_18bar;
  wire in_17bar;
  wire in_16bar;
  wire in_15bar;
  wire in_14bar;
  wire in_13bar;
  wire in_12bar;
  wire in_11bar;
  wire in_10bar;
  wire in_9bar;
  wire in_8bar;
  wire in_7bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_3bar;
  wire in_2bar;
  wire in_1bar;
  wire in_0bar;
  wire n487bar;
  wire n488bar;
  wire n489bar;
  wire n490bar;
  wire n491bar;
  wire n492bar;
  wire n493bar;
  wire n494bar;
  wire n495bar;
  wire n496bar;
  wire n497bar;
  wire n498bar;
  wire n499bar;
  wire n500bar;
  wire n501bar;
  wire n502bar;
  wire n503bar;
  wire n504bar;
  wire n505bar;
  wire n506bar;
  wire n507bar;
  wire n508bar;
  wire n509bar;
  wire n510bar;
  wire n511bar;
  wire n512bar;
  wire n513bar;
  wire n514bar;
  wire n515bar;
  wire n516bar;
  wire n517bar;
  wire n518bar;
  wire n519bar;
  wire n520bar;
  wire n521bar;
  wire n522bar;
  wire n523bar;
  wire n524bar;
  wire n525bar;
  wire n526bar;
  wire n527bar;
  wire n528bar;
  wire n529bar;
  wire n530bar;
  wire n531bar;
  wire n532bar;
  wire n533bar;
  wire n534bar;
  wire n535bar;
  wire n536bar;
  wire n537bar;
  wire n538bar;
  wire n539bar;
  wire n540bar;
  wire n541bar;
  wire n542bar;
  wire n543bar;
  wire n544bar;
  wire n545bar;
  wire n546bar;
  wire n547bar;
  wire n548bar;
  wire n549bar;
  wire n550bar;
  wire n551bar;
  wire n552bar;
  wire n553bar;
  wire n554bar;
  wire n555bar;
  wire n556bar;
  wire n557bar;
  wire n558bar;
  wire n559bar;
  wire n560bar;
  wire n561bar;
  wire n562bar;
  wire n563bar;
  wire n564bar;
  wire n565bar;
  wire n566bar;
  wire n567bar;
  wire n568bar;
  wire n569bar;
  wire n570bar;
  wire n571bar;
  wire n572bar;
  wire n573bar;
  wire n574bar;
  wire n575bar;
  wire n576bar;
  wire n577bar;
  wire n578bar;
  wire n579bar;
  wire n580bar;
  wire n581bar;
  wire n582bar;
  wire n583bar;
  wire n584bar;
  wire n585bar;
  wire n586bar;
  wire n587bar;
  wire n588bar;
  wire n589bar;
  wire n590bar;
  wire n591bar;
  wire n592bar;
  wire n593bar;
  wire n594bar;
  wire n595bar;
  wire n596bar;
  wire n597bar;
  wire n598bar;
  wire n599bar;
  wire n600bar;
  wire n601bar;
  wire n602bar;
  wire n603bar;
  wire n604bar;
  wire n605bar;
  wire n606bar;
  wire n607bar;
  wire n608bar;
  wire n609bar;
  wire n610bar;
  wire n611bar;
  wire n612bar;
  wire n613bar;
  wire n614bar;
  wire n615bar;
  wire n616bar;
  wire n617bar;
  wire n618bar;
  wire n619bar;
  wire n620bar;
  wire n621bar;
  wire n622bar;
  wire n623bar;
  wire n624bar;
  wire n625bar;
  wire n626bar;
  wire n627bar;
  wire n628bar;
  wire n629bar;
  wire n630bar;
  wire n631bar;
  wire n632bar;
  wire n633bar;
  wire n634bar;
  wire n635bar;
  wire n636bar;
  wire n637bar;
  wire n638bar;
  wire n639bar;
  wire n640bar;
  wire n641bar;
  wire n642bar;
  wire n643bar;
  wire n644bar;
  wire n645bar;
  wire n646bar;
  wire n647bar;
  wire n648bar;
  wire n649bar;
  wire n650bar;
  wire n651bar;
  wire n652bar;
  wire n653bar;
  wire n654bar;
  wire n655bar;
  wire n656bar;
  wire n657bar;
  wire n658bar;
  wire n659bar;
  wire n660bar;
  wire n661bar;
  wire n662bar;
  wire n663bar;
  wire n664bar;
  wire n665bar;
  wire n666bar;
  wire n667bar;
  wire n668bar;
  wire n669bar;
  wire n670bar;
  wire n671bar;
  wire n672bar;
  wire n673bar;
  wire n674bar;
  wire n675bar;
  wire n676bar;
  wire n677bar;
  wire n678bar;
  wire n679bar;
  wire n680bar;
  wire n681bar;
  wire n682bar;
  wire n683bar;
  wire n684bar;
  wire n685bar;
  wire n686bar;
  wire n687bar;
  wire n688bar;
  wire n689bar;
  wire n690bar;
  wire n691bar;
  wire n692bar;
  wire n693bar;
  wire n694bar;
  wire n695bar;
  wire n696bar;
  wire n697bar;
  wire n698bar;
  wire n699bar;
  wire n700bar;
  wire n701bar;
  wire n702bar;
  wire n703bar;
  wire n704bar;
  wire n705bar;
  wire n706bar;
  wire n707bar;
  wire n708bar;
  wire n709bar;
  wire n710bar;
  wire n711bar;
  wire n712bar;
  wire n713bar;
  wire n714bar;
  wire n715bar;
  wire n716bar;
  wire n717bar;
  wire n718bar;
  wire n719bar;
  wire n720bar;
  wire n721bar;
  wire n722bar;
  wire n723bar;
  wire n724bar;
  wire n725bar;
  wire n726bar;
  wire n727bar;
  wire n728bar;
  wire n729bar;
  wire n730bar;
  wire n731bar;
  wire n732bar;
  wire n733bar;
  wire n734bar;
  wire n735bar;
  wire n736bar;
  wire n737bar;
  wire n738bar;
  wire n739bar;
  wire n740bar;
  wire n741bar;
  wire n742bar;
  wire n743bar;
  wire n744bar;
  wire n745bar;
  wire n746bar;
  wire n747bar;
  wire n748bar;
  wire n749bar;
  wire n750bar;
  wire n751bar;
  wire n752bar;
  wire n753bar;
  wire n754bar;
  wire n755bar;
  wire n756bar;
  wire n757bar;
  wire n758bar;
  wire n759bar;
  wire n760bar;
  wire n761bar;
  wire n762bar;
  wire n763bar;
  wire n764bar;
  wire n765bar;
  wire n766bar;
  wire n767bar;
  wire n768bar;
  wire n769bar;
  wire n770bar;
  wire n771bar;
  wire n772bar;
  wire n773bar;
  wire n774bar;
  wire n775bar;
  wire n776bar;
  wire n777bar;
  wire n778bar;
  wire n779bar;
  wire n780bar;
  wire n781bar;
  wire n782bar;
  wire n783bar;
  wire n784bar;
  wire n785bar;
  wire n786bar;
  wire n787bar;
  wire n788bar;
  wire n789bar;
  wire n790bar;
  wire n791bar;
  wire n792bar;
  wire n793bar;
  wire n794bar;
  wire n795bar;
  wire n796bar;
  wire n797bar;
  wire n798bar;
  wire n799bar;
  wire n800bar;
  wire n801bar;
  wire n802bar;
  wire n803bar;
  wire n804bar;
  wire n805bar;
  wire n806bar;
  wire n807bar;
  wire n808bar;
  wire n809bar;
  wire n810bar;
  wire n811bar;
  wire n812bar;
  wire n813bar;
  wire n814bar;
  wire n815bar;
  wire n816bar;
  wire n817bar;
  wire n818bar;
  wire n819bar;
  wire n820bar;
  wire n821bar;
  wire n822bar;
  wire n823bar;
  wire n824bar;
  wire n825bar;
  wire n826bar;
  wire n827bar;
  wire n828bar;
  wire n829bar;
  wire n830bar;
  wire n831bar;
  wire n832bar;
  wire n833bar;
  wire n834bar;
  wire n835bar;
  wire n836bar;
  wire n837bar;
  wire n838bar;
  wire n839bar;
  wire n840bar;
  wire n841bar;
  wire n842bar;
  wire n843bar;
  wire n844bar;
  wire n845bar;
  wire n846bar;
  wire n847bar;
  wire n848bar;
  wire n849bar;
  wire n850bar;
  wire n851bar;
  wire n852bar;
  wire n853bar;
  wire n854bar;
  wire n855bar;
  wire n856bar;
  wire n857bar;
  wire n858bar;
  wire n859bar;
  wire n860bar;
  wire n861bar;
  wire n862bar;
  wire n863bar;
  wire n864bar;
  wire n865bar;
  wire n866bar;
  wire n867bar;
  wire n868bar;
  wire n869bar;
  wire n870bar;
  wire n871bar;
  wire n872bar;
  wire n873bar;
  wire n874bar;
  wire n875bar;
  wire n876bar;
  wire n877bar;
  wire n878bar;
  wire n879bar;
  wire n880bar;
  wire n881bar;
  wire n882bar;
  wire n883bar;
  wire n884bar;
  wire n885bar;
  wire n886bar;
  wire n887bar;
  wire n888bar;
  wire n889bar;
  wire n890bar;
  wire n891bar;
  wire n892bar;
  wire n893bar;
  wire n894bar;
  wire n895bar;
  wire n896bar;
  wire n897bar;
  wire n898bar;
  wire n899bar;
  wire n900bar;
  wire n901bar;
  wire n902bar;
  wire n903bar;
  wire n904bar;
  wire n905bar;
  wire n906bar;
  wire n907bar;
  wire n908bar;
  wire n909bar;
  wire n910bar;
  wire n911bar;
  wire n912bar;
  wire n913bar;
  wire n914bar;
  wire n915bar;
  wire n916bar;
  wire n917bar;
  wire n918bar;
  wire n919bar;
  wire n920bar;
  wire n921bar;
  wire n922bar;
  wire n923bar;
  wire n924bar;
  wire n925bar;
  wire n926bar;
  wire n927bar;
  wire n928bar;
  wire n929bar;
  wire n930bar;
  wire n931bar;
  wire n932bar;
  wire n933bar;
  wire n934bar;
  wire n935bar;
  wire n936bar;
  wire n937bar;
  wire n938bar;
  wire n939bar;
  wire n940bar;
  wire n941bar;
  wire n942bar;
  wire n943bar;
  wire n944bar;
  wire n945bar;
  wire n946bar;
  wire n947bar;
  wire n948bar;
  wire n949bar;
  wire n950bar;
  wire n951bar;
  wire n952bar;
  wire n953bar;
  wire n954bar;
  wire n955bar;
  wire n956bar;
  wire n957bar;
  wire n958bar;
  wire n959bar;
  wire n960bar;
  wire n961bar;
  wire n962bar;
  wire n963bar;
  wire n964bar;
  wire n965bar;
  wire n966bar;
  wire n967bar;
  wire n968bar;
  wire n969bar;
  wire n970bar;
  wire n971bar;
  wire n972bar;
//wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];
  //OR U1
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1 (
    .O(out[7]),
    .I0(n972),
    .I1(n971)
  );
  //AND U1bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1bar (
    .O(outbar[7]),
    .I0(n972bar),
    .I1(n971bar)
  );
  //OR U2
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2 (
    .O(n971),
    .I0(n970),
    .I1(n969)
  );
  //AND U2bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2bar (
    .O(n971bar),
    .I0(n970bar),
    .I1(n969bar)
  );
  //OR U3
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3 (
    .O(n969),
    .I0(n968),
    .I1(n967)
  );
  //AND U3bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3bar (
    .O(n969bar),
    .I0(n968bar),
    .I1(n967bar)
  );
  //OR U4
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4 (
    .O(n967),
    .I0(n966),
    .I1(n965)
  );
  //AND U4bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4bar (
    .O(n967bar),
    .I0(n966bar),
    .I1(n965bar)
  );
  //OR U5
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5 (
    .O(n968),
    .I0(n964),
    .I1(n963)
  );
  //AND U5bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5bar (
    .O(n968bar),
    .I0(n964bar),
    .I1(n963bar)
  );
  //OR U6
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6 (
    .O(n963),
    .I0(in[116]),
    .I1(n962)
  );
  //AND U6bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6bar (
    .O(n963bar),
    .I0(inbar[116]),
    .I1(n962bar)
  );
  //OR U7
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7 (
    .O(n970),
    .I0(n961),
    .I1(n960)
  );
  //AND U7bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7bar (
    .O(n970bar),
    .I0(n961bar),
    .I1(n960bar)
  );
  //OR U8
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8 (
    .O(n960),
    .I0(in[150]),
    .I1(in[127])
  );
  //AND U8bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8bar (
    .O(n960bar),
    .I0(inbar[150]),
    .I1(inbar[127])
  );
  //OR U9
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9 (
    .O(n961),
    .I0(in[160]),
    .I1(n959)
  );
  //AND U9bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9bar (
    .O(n961bar),
    .I0(inbar[160]),
    .I1(n959bar)
  );
  //OR U10
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10 (
    .O(n959),
    .I0(in[252]),
    .I1(in[168])
  );
  //AND U10bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10bar (
    .O(n959bar),
    .I0(inbar[252]),
    .I1(inbar[168])
  );
  //OR U11
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11 (
    .O(n972),
    .I0(n958),
    .I1(n957)
  );
  //AND U11bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11bar (
    .O(n972bar),
    .I0(n958bar),
    .I1(n957bar)
  );
  //OR U12
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12 (
    .O(n957),
    .I0(n956),
    .I1(n955)
  );
  //AND U12bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12bar (
    .O(n957bar),
    .I0(n956bar),
    .I1(n955bar)
  );
  //OR U13
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13 (
    .O(n955),
    .I0(in_17),
    .I1(in[96])
  );
  //AND U13bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13bar (
    .O(n955bar),
    .I0(in_17bar),
    .I1(inbar[96])
  );
  //OR U14
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14 (
    .O(n956),
    .I0(in_23),
    .I1(n954)
  );
  //AND U14bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14bar (
    .O(n956bar),
    .I0(in_23bar),
    .I1(n954bar)
  );
  //OR U15
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15 (
    .O(n954),
    .I0(in_31),
    .I1(in_26)
  );
  //AND U15bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15bar (
    .O(n954bar),
    .I0(in_31bar),
    .I1(in_26bar)
  );
  //OR U16
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16 (
    .O(n958),
    .I0(n953),
    .I1(n952)
  );
  //AND U16bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16bar (
    .O(n958bar),
    .I0(n953bar),
    .I1(n952bar)
  );
  //OR U17
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U17 (
    .O(n952),
    .I0(in_58),
    .I1(in_4)
  );
  //AND U17bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U17bar (
    .O(n952bar),
    .I0(in_58bar),
    .I1(in_4bar)
  );
  //OR U18
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U18 (
    .O(n953),
    .I0(in_59),
    .I1(n951)
  );
  //AND U18bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U18bar (
    .O(n953bar),
    .I0(in_59bar),
    .I1(n951bar)
  );
  //OR U19
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U19 (
    .O(n951),
    .I0(in_71),
    .I1(in_62)
  );
  //AND U19bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U19bar (
    .O(n951bar),
    .I0(in_71bar),
    .I1(in_62bar)
  );
  //OR U20
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U20 (
    .O(out[6]),
    .I0(n950),
    .I1(n949)
  );
  //AND U20bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U20bar (
    .O(outbar[6]),
    .I0(n950bar),
    .I1(n949bar)
  );
  //OR U21
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U21 (
    .O(n949),
    .I0(n948),
    .I1(n947)
  );
  //AND U21bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U21bar (
    .O(n949bar),
    .I0(n948bar),
    .I1(n947bar)
  );
  //OR U22
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U22 (
    .O(n947),
    .I0(n946),
    .I1(n945)
  );
  //AND U22bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U22bar (
    .O(n947bar),
    .I0(n946bar),
    .I1(n945bar)
  );
  //OR U23
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U23 (
    .O(n945),
    .I0(n944),
    .I1(n943)
  );
  //AND U23bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U23bar (
    .O(n945bar),
    .I0(n944bar),
    .I1(n943bar)
  );
  //OR U24
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U24 (
    .O(n946),
    .I0(n942),
    .I1(n941)
  );
  //AND U24bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U24bar (
    .O(n946bar),
    .I0(n942bar),
    .I1(n941bar)
  );
  //OR U25
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U25 (
    .O(n941),
    .I0(in[101]),
    .I1(n940)
  );
  //AND U25bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U25bar (
    .O(n941bar),
    .I0(inbar[101]),
    .I1(n940bar)
  );
  //OR U26
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U26 (
    .O(n948),
    .I0(n939),
    .I1(n938)
  );
  //AND U26bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U26bar (
    .O(n948bar),
    .I0(n939bar),
    .I1(n938bar)
  );
  //OR U27
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U27 (
    .O(n938),
    .I0(in[114]),
    .I1(in[104])
  );
  //AND U27bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U27bar (
    .O(n938bar),
    .I0(inbar[114]),
    .I1(inbar[104])
  );
  //OR U28
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U28 (
    .O(n939),
    .I0(in[128]),
    .I1(n937)
  );
  //AND U28bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U28bar (
    .O(n939bar),
    .I0(inbar[128]),
    .I1(n937bar)
  );
  //OR U29
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U29 (
    .O(n937),
    .I0(in[136]),
    .I1(in[134])
  );
  //AND U29bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U29bar (
    .O(n937bar),
    .I0(inbar[136]),
    .I1(inbar[134])
  );
  //OR U30
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U30 (
    .O(n950),
    .I0(n936),
    .I1(n935)
  );
  //AND U30bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U30bar (
    .O(n950bar),
    .I0(n936bar),
    .I1(n935bar)
  );
  //OR U31
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U31 (
    .O(n935),
    .I0(n934),
    .I1(n933)
  );
  //AND U31bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U31bar (
    .O(n935bar),
    .I0(n934bar),
    .I1(n933bar)
  );
  //OR U32
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U32 (
    .O(n933),
    .I0(in[177]),
    .I1(in[164])
  );
  //AND U32bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U32bar (
    .O(n933bar),
    .I0(inbar[177]),
    .I1(inbar[164])
  );
  //OR U33
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U33 (
    .O(n934),
    .I0(in[212]),
    .I1(n932)
  );
  //AND U33bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U33bar (
    .O(n934bar),
    .I0(inbar[212]),
    .I1(n932bar)
  );
  //OR U34
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U34 (
    .O(n932),
    .I0(in[248]),
    .I1(in[221])
  );
  //AND U34bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U34bar (
    .O(n932bar),
    .I0(inbar[248]),
    .I1(inbar[221])
  );
  //OR U35
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U35 (
    .O(n936),
    .I0(n931),
    .I1(n930)
  );
  //AND U35bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U35bar (
    .O(n936bar),
    .I0(n931bar),
    .I1(n930bar)
  );
  //OR U36
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U36 (
    .O(n930),
    .I0(in_18),
    .I1(in[93])
  );
  //AND U36bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U36bar (
    .O(n930bar),
    .I0(in_18bar),
    .I1(inbar[93])
  );
  //OR U37
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U37 (
    .O(n931),
    .I0(in_31),
    .I1(n929)
  );
  //AND U37bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U37bar (
    .O(n931bar),
    .I0(in_31bar),
    .I1(n929bar)
  );
  //OR U38
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U38 (
    .O(n929),
    .I0(in_7),
    .I1(in_39)
  );
  //AND U38bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U38bar (
    .O(n929bar),
    .I0(in_7bar),
    .I1(in_39bar)
  );
  //OR U39
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U39 (
    .O(out[5]),
    .I0(n928),
    .I1(n927)
  );
  //AND U39bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U39bar (
    .O(outbar[5]),
    .I0(n928bar),
    .I1(n927bar)
  );
  //OR U40
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U40 (
    .O(n927),
    .I0(n926),
    .I1(n925)
  );
  //AND U40bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U40bar (
    .O(n927bar),
    .I0(n926bar),
    .I1(n925bar)
  );
  //OR U41
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U41 (
    .O(n925),
    .I0(n924),
    .I1(n923)
  );
  //AND U41bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U41bar (
    .O(n925bar),
    .I0(n924bar),
    .I1(n923bar)
  );
  //OR U42
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U42 (
    .O(n923),
    .I0(n922),
    .I1(n921)
  );
  //AND U42bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U42bar (
    .O(n923bar),
    .I0(n922bar),
    .I1(n921bar)
  );
  //OR U43
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U43 (
    .O(n924),
    .I0(n940),
    .I1(n920)
  );
  //AND U43bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U43bar (
    .O(n924bar),
    .I0(n940bar),
    .I1(n920bar)
  );
  //OR U44
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U44 (
    .O(n920),
    .I0(in[111]),
    .I1(n919)
  );
  //AND U44bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U44bar (
    .O(n920bar),
    .I0(inbar[111]),
    .I1(n919bar)
  );
  //OR U45
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U45 (
    .O(n940),
    .I0(n918),
    .I1(n917)
  );
  //AND U45bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U45bar (
    .O(n940bar),
    .I0(n918bar),
    .I1(n917bar)
  );
  //OR U46
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U46 (
    .O(n917),
    .I0(n916),
    .I1(n915)
  );
  //AND U46bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U46bar (
    .O(n917bar),
    .I0(n916bar),
    .I1(n915bar)
  );
  //OR U47
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U47 (
    .O(n915),
    .I0(n914),
    .I1(n913)
  );
  //AND U47bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U47bar (
    .O(n915bar),
    .I0(n914bar),
    .I1(n913bar)
  );
  //OR U48
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U48 (
    .O(n913),
    .I0(in[140]),
    .I1(in[131])
  );
  //AND U48bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U48bar (
    .O(n913bar),
    .I0(inbar[140]),
    .I1(inbar[131])
  );
  //OR U49
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U49 (
    .O(n914),
    .I0(in[160]),
    .I1(in[144])
  );
  //AND U49bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U49bar (
    .O(n914bar),
    .I0(inbar[160]),
    .I1(inbar[144])
  );
  //OR U50
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U50 (
    .O(n916),
    .I0(n912),
    .I1(n911)
  );
  //AND U50bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U50bar (
    .O(n916bar),
    .I0(n912bar),
    .I1(n911bar)
  );
  //OR U51
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U51 (
    .O(n911),
    .I0(in[179]),
    .I1(in[174])
  );
  //AND U51bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U51bar (
    .O(n911bar),
    .I0(inbar[179]),
    .I1(inbar[174])
  );
  //OR U52
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U52 (
    .O(n912),
    .I0(in[188]),
    .I1(in[184])
  );
  //AND U52bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U52bar (
    .O(n912bar),
    .I0(inbar[188]),
    .I1(inbar[184])
  );
  //OR U53
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U53 (
    .O(n918),
    .I0(n910),
    .I1(n909)
  );
  //AND U53bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U53bar (
    .O(n918bar),
    .I0(n910bar),
    .I1(n909bar)
  );
  //OR U54
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U54 (
    .O(n909),
    .I0(n908),
    .I1(n907)
  );
  //AND U54bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U54bar (
    .O(n909bar),
    .I0(n908bar),
    .I1(n907bar)
  );
  //OR U55
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U55 (
    .O(n907),
    .I0(in[216]),
    .I1(in[200])
  );
  //AND U55bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U55bar (
    .O(n907bar),
    .I0(inbar[216]),
    .I1(inbar[200])
  );
  //OR U56
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U56 (
    .O(n908),
    .I0(in[228]),
    .I1(in[224])
  );
  //AND U56bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U56bar (
    .O(n908bar),
    .I0(inbar[228]),
    .I1(inbar[224])
  );
  //OR U57
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U57 (
    .O(n910),
    .I0(n906),
    .I1(n905)
  );
  //AND U57bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U57bar (
    .O(n910bar),
    .I0(n906bar),
    .I1(n905bar)
  );
  //OR U58
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U58 (
    .O(n905),
    .I0(in[247]),
    .I1(in[235])
  );
  //AND U58bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U58bar (
    .O(n905bar),
    .I0(inbar[247]),
    .I1(inbar[235])
  );
  //OR U59
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U59 (
    .O(n906),
    .I0(in_42),
    .I1(in[83])
  );
  //AND U59bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U59bar (
    .O(n906bar),
    .I0(in_42bar),
    .I1(inbar[83])
  );
  //OR U60
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U60 (
    .O(n926),
    .I0(n904),
    .I1(n903)
  );
  //AND U60bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U60bar (
    .O(n926bar),
    .I0(n904bar),
    .I1(n903bar)
  );
  //OR U61
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U61 (
    .O(n903),
    .I0(in[166]),
    .I1(in[123])
  );
  //AND U61bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U61bar (
    .O(n903bar),
    .I0(inbar[166]),
    .I1(inbar[123])
  );
  //OR U62
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U62 (
    .O(n904),
    .I0(in[170]),
    .I1(n902)
  );
  //AND U62bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U62bar (
    .O(n904bar),
    .I0(inbar[170]),
    .I1(n902bar)
  );
  //OR U63
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U63 (
    .O(n902),
    .I0(in[194]),
    .I1(in[183])
  );
  //AND U63bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U63bar (
    .O(n902bar),
    .I0(inbar[194]),
    .I1(inbar[183])
  );
  //OR U64
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U64 (
    .O(n928),
    .I0(n901),
    .I1(n900)
  );
  //AND U64bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U64bar (
    .O(n928bar),
    .I0(n901bar),
    .I1(n900bar)
  );
  //OR U65
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U65 (
    .O(n900),
    .I0(n899),
    .I1(n898)
  );
  //AND U65bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U65bar (
    .O(n900bar),
    .I0(n899bar),
    .I1(n898bar)
  );
  //OR U66
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U66 (
    .O(n898),
    .I0(in[241]),
    .I1(in[238])
  );
  //AND U66bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U66bar (
    .O(n898bar),
    .I0(inbar[241]),
    .I1(inbar[238])
  );
  //OR U67
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U67 (
    .O(n899),
    .I0(in[250]),
    .I1(n897)
  );
  //AND U67bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U67bar (
    .O(n899bar),
    .I0(inbar[250]),
    .I1(n897bar)
  );
  //OR U68
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U68 (
    .O(n897),
    .I0(in_24),
    .I1(in[84])
  );
  //AND U68bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U68bar (
    .O(n897bar),
    .I0(in_24bar),
    .I1(inbar[84])
  );
  //OR U69
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U69 (
    .O(n901),
    .I0(n896),
    .I1(n895)
  );
  //AND U69bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U69bar (
    .O(n901bar),
    .I0(n896bar),
    .I1(n895bar)
  );
  //OR U70
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U70 (
    .O(n895),
    .I0(in_41),
    .I1(in_29)
  );
  //AND U70bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U70bar (
    .O(n895bar),
    .I0(in_41bar),
    .I1(in_29bar)
  );
  //OR U71
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U71 (
    .O(n896),
    .I0(in_66),
    .I1(n894)
  );
  //AND U71bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U71bar (
    .O(n896bar),
    .I0(in_66bar),
    .I1(n894bar)
  );
  //OR U72
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U72 (
    .O(n894),
    .I0(in_76),
    .I1(in_71)
  );
  //AND U72bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U72bar (
    .O(n894bar),
    .I0(in_76bar),
    .I1(in_71bar)
  );
  //OR U73
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U73 (
    .O(out[4]),
    .I0(n893),
    .I1(n892)
  );
  //AND U73bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U73bar (
    .O(outbar[4]),
    .I0(n893bar),
    .I1(n892bar)
  );
  //OR U74
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U74 (
    .O(n892),
    .I0(n891),
    .I1(n890)
  );
  //AND U74bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U74bar (
    .O(n892bar),
    .I0(n891bar),
    .I1(n890bar)
  );
  //OR U75
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U75 (
    .O(n890),
    .I0(n889),
    .I1(n888)
  );
  //AND U75bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U75bar (
    .O(n890bar),
    .I0(n889bar),
    .I1(n888bar)
  );
  //OR U76
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U76 (
    .O(n888),
    .I0(n922),
    .I1(n887)
  );
  //AND U76bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U76bar (
    .O(n888bar),
    .I0(n922bar),
    .I1(n887bar)
  );
  //OR U77
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U77 (
    .O(n922),
    .I0(n886),
    .I1(n885)
  );
  //AND U77bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U77bar (
    .O(n922bar),
    .I0(n886bar),
    .I1(n885bar)
  );
  //OR U78
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U78 (
    .O(n885),
    .I0(n884),
    .I1(n883)
  );
  //AND U78bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U78bar (
    .O(n885bar),
    .I0(n884bar),
    .I1(n883bar)
  );
  //OR U79
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U79 (
    .O(n883),
    .I0(n882),
    .I1(n881)
  );
  //AND U79bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U79bar (
    .O(n883bar),
    .I0(n882bar),
    .I1(n881bar)
  );
  //OR U80
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U80 (
    .O(n881),
    .I0(in[118]),
    .I1(in[109])
  );
  //AND U80bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U80bar (
    .O(n881bar),
    .I0(inbar[118]),
    .I1(inbar[109])
  );
  //OR U81
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U81 (
    .O(n882),
    .I0(in[139]),
    .I1(in[120])
  );
  //AND U81bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U81bar (
    .O(n882bar),
    .I0(inbar[139]),
    .I1(inbar[120])
  );
  //OR U82
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U82 (
    .O(n884),
    .I0(n880),
    .I1(n879)
  );
  //AND U82bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U82bar (
    .O(n884bar),
    .I0(n880bar),
    .I1(n879bar)
  );
  //OR U83
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U83 (
    .O(n879),
    .I0(in[198]),
    .I1(in[154])
  );
  //AND U83bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U83bar (
    .O(n879bar),
    .I0(inbar[198]),
    .I1(inbar[154])
  );
  //OR U84
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U84 (
    .O(n880),
    .I0(in[210]),
    .I1(in[205])
  );
  //AND U84bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U84bar (
    .O(n880bar),
    .I0(inbar[210]),
    .I1(inbar[205])
  );
  //OR U85
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U85 (
    .O(n886),
    .I0(n878),
    .I1(n877)
  );
  //AND U85bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U85bar (
    .O(n886bar),
    .I0(n878bar),
    .I1(n877bar)
  );
  //OR U86
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U86 (
    .O(n877),
    .I0(n876),
    .I1(n875)
  );
  //AND U86bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U86bar (
    .O(n877bar),
    .I0(n876bar),
    .I1(n875bar)
  );
  //OR U87
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U87 (
    .O(n875),
    .I0(in[219]),
    .I1(in[217])
  );
  //AND U87bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U87bar (
    .O(n875bar),
    .I0(inbar[219]),
    .I1(inbar[217])
  );
  //OR U88
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U88 (
    .O(n876),
    .I0(in[86]),
    .I1(in[252])
  );
  //AND U88bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U88bar (
    .O(n876bar),
    .I0(inbar[86]),
    .I1(inbar[252])
  );
  //OR U89
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U89 (
    .O(n878),
    .I0(n874),
    .I1(n873)
  );
  //AND U89bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U89bar (
    .O(n878bar),
    .I0(n874bar),
    .I1(n873bar)
  );
  //OR U90
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U90 (
    .O(n873),
    .I0(in_40),
    .I1(in[91])
  );
  //AND U90bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U90bar (
    .O(n873bar),
    .I0(in_40bar),
    .I1(inbar[91])
  );
  //OR U91
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U91 (
    .O(n874),
    .I0(in_8),
    .I1(in_46)
  );
  //AND U91bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U91bar (
    .O(n874bar),
    .I0(in_8bar),
    .I1(in_46bar)
  );
  //OR U92
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U92 (
    .O(n889),
    .I0(n872),
    .I1(n871)
  );
  //AND U92bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U92bar (
    .O(n889bar),
    .I0(n872bar),
    .I1(n871bar)
  );
  //OR U93
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U93 (
    .O(n871),
    .I0(in[117]),
    .I1(n943)
  );
  //AND U93bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U93bar (
    .O(n871bar),
    .I0(inbar[117]),
    .I1(n943bar)
  );
  //OR U94
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U94 (
    .O(n943),
    .I0(n870),
    .I1(n869)
  );
  //AND U94bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U94bar (
    .O(n943bar),
    .I0(n870bar),
    .I1(n869bar)
  );
  //OR U95
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U95 (
    .O(n869),
    .I0(n868),
    .I1(n867)
  );
  //AND U95bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U95bar (
    .O(n869bar),
    .I0(n868bar),
    .I1(n867bar)
  );
  //OR U96
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U96 (
    .O(n867),
    .I0(n866),
    .I1(n865)
  );
  //AND U96bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U96bar (
    .O(n867bar),
    .I0(n866bar),
    .I1(n865bar)
  );
  //OR U97
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U97 (
    .O(n865),
    .I0(n864),
    .I1(n863)
  );
  //AND U97bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U97bar (
    .O(n865bar),
    .I0(n864bar),
    .I1(n863bar)
  );
  //OR U98
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U98 (
    .O(n866),
    .I0(in[108]),
    .I1(n919)
  );
  //AND U98bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U98bar (
    .O(n866bar),
    .I0(inbar[108]),
    .I1(n919bar)
  );
  //OR U99
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U99 (
    .O(n919),
    .I0(n862),
    .I1(n861)
  );
  //AND U99bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U99bar (
    .O(n919bar),
    .I0(n862bar),
    .I1(n861bar)
  );
  //OR U100
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U100 (
    .O(n861),
    .I0(n860),
    .I1(n859)
  );
  //AND U100bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U100bar (
    .O(n861bar),
    .I0(n860bar),
    .I1(n859bar)
  );
  //OR U101
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U101 (
    .O(n859),
    .I0(n858),
    .I1(n857)
  );
  //AND U101bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U101bar (
    .O(n859bar),
    .I0(n858bar),
    .I1(n857bar)
  );
  //OR U102
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U102 (
    .O(n857),
    .I0(in[119]),
    .I1(in[105])
  );
  //AND U102bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U102bar (
    .O(n857bar),
    .I0(inbar[119]),
    .I1(inbar[105])
  );
  //OR U103
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U103 (
    .O(n858),
    .I0(in[186]),
    .I1(in[175])
  );
  //AND U103bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U103bar (
    .O(n858bar),
    .I0(inbar[186]),
    .I1(inbar[175])
  );
  //OR U104
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U104 (
    .O(n860),
    .I0(n856),
    .I1(n855)
  );
  //AND U104bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U104bar (
    .O(n860bar),
    .I0(n856bar),
    .I1(n855bar)
  );
  //OR U105
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U105 (
    .O(n855),
    .I0(in[202]),
    .I1(in[193])
  );
  //AND U105bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U105bar (
    .O(n855bar),
    .I0(inbar[202]),
    .I1(inbar[193])
  );
  //OR U106
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U106 (
    .O(n856),
    .I0(in[225]),
    .I1(in[208])
  );
  //AND U106bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U106bar (
    .O(n856bar),
    .I0(inbar[225]),
    .I1(inbar[208])
  );
  //OR U107
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U107 (
    .O(n862),
    .I0(n854),
    .I1(n853)
  );
  //AND U107bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U107bar (
    .O(n862bar),
    .I0(n854bar),
    .I1(n853bar)
  );
  //OR U108
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U108 (
    .O(n853),
    .I0(n852),
    .I1(n851)
  );
  //AND U108bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U108bar (
    .O(n853bar),
    .I0(n852bar),
    .I1(n851bar)
  );
  //OR U109
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U109 (
    .O(n851),
    .I0(in_1),
    .I1(in[85])
  );
  //AND U109bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U109bar (
    .O(n851bar),
    .I0(in_1bar),
    .I1(inbar[85])
  );
  //OR U110
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U110 (
    .O(n852),
    .I0(in_23),
    .I1(in_19)
  );
  //AND U110bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U110bar (
    .O(n852bar),
    .I0(in_23bar),
    .I1(in_19bar)
  );
  //OR U111
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U111 (
    .O(n854),
    .I0(n850),
    .I1(n849)
  );
  //AND U111bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U111bar (
    .O(n854bar),
    .I0(n850bar),
    .I1(n849bar)
  );
  //OR U112
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U112 (
    .O(n849),
    .I0(in_43),
    .I1(in_33)
  );
  //AND U112bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U112bar (
    .O(n849bar),
    .I0(in_43bar),
    .I1(in_33bar)
  );
  //OR U113
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U113 (
    .O(n850),
    .I0(in_63),
    .I1(in_44)
  );
  //AND U113bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U113bar (
    .O(n850bar),
    .I0(in_63bar),
    .I1(in_44bar)
  );
  //OR U114
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U114 (
    .O(n868),
    .I0(n848),
    .I1(n847)
  );
  //AND U114bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U114bar (
    .O(n868bar),
    .I0(n848bar),
    .I1(n847bar)
  );
  //OR U115
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U115 (
    .O(n847),
    .I0(in[141]),
    .I1(in[112])
  );
  //AND U115bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U115bar (
    .O(n847bar),
    .I0(inbar[141]),
    .I1(inbar[112])
  );
  //OR U116
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U116 (
    .O(n848),
    .I0(in[147]),
    .I1(n846)
  );
  //AND U116bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U116bar (
    .O(n848bar),
    .I0(inbar[147]),
    .I1(n846bar)
  );
  //OR U117
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U117 (
    .O(n846),
    .I0(in[181]),
    .I1(in[167])
  );
  //AND U117bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U117bar (
    .O(n846bar),
    .I0(inbar[181]),
    .I1(inbar[167])
  );
  //OR U118
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U118 (
    .O(n870),
    .I0(n845),
    .I1(n844)
  );
  //AND U118bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U118bar (
    .O(n870bar),
    .I0(n845bar),
    .I1(n844bar)
  );
  //OR U119
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U119 (
    .O(n844),
    .I0(n843),
    .I1(n842)
  );
  //AND U119bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U119bar (
    .O(n844bar),
    .I0(n843bar),
    .I1(n842bar)
  );
  //OR U120
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U120 (
    .O(n842),
    .I0(in[229]),
    .I1(in[201])
  );
  //AND U120bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U120bar (
    .O(n842bar),
    .I0(inbar[229]),
    .I1(inbar[201])
  );
  //OR U121
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U121 (
    .O(n843),
    .I0(in[237]),
    .I1(n841)
  );
  //AND U121bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U121bar (
    .O(n843bar),
    .I0(inbar[237]),
    .I1(n841bar)
  );
  //OR U122
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U122 (
    .O(n841),
    .I0(in[94]),
    .I1(in[253])
  );
  //AND U122bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U122bar (
    .O(n841bar),
    .I0(inbar[94]),
    .I1(inbar[253])
  );
  //OR U123
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U123 (
    .O(n845),
    .I0(n840),
    .I1(n839)
  );
  //AND U123bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U123bar (
    .O(n845bar),
    .I0(n840bar),
    .I1(n839bar)
  );
  //OR U124
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U124 (
    .O(n839),
    .I0(in_21),
    .I1(in[96])
  );
  //AND U124bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U124bar (
    .O(n839bar),
    .I0(in_21bar),
    .I1(inbar[96])
  );
  //OR U125
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U125 (
    .O(n840),
    .I0(in_25),
    .I1(n838)
  );
  //AND U125bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U125bar (
    .O(n840bar),
    .I0(in_25bar),
    .I1(n838bar)
  );
  //OR U126
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U126 (
    .O(n838),
    .I0(in_81),
    .I1(in_45)
  );
  //AND U126bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U126bar (
    .O(n838bar),
    .I0(in_81bar),
    .I1(in_45bar)
  );
  //OR U127
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U127 (
    .O(n891),
    .I0(n837),
    .I1(n836)
  );
  //AND U127bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U127bar (
    .O(n891bar),
    .I0(n837bar),
    .I1(n836bar)
  );
  //OR U128
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U128 (
    .O(n836),
    .I0(in[142]),
    .I1(in[124])
  );
  //AND U128bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U128bar (
    .O(n836bar),
    .I0(inbar[142]),
    .I1(inbar[124])
  );
  //OR U129
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U129 (
    .O(n837),
    .I0(in[150]),
    .I1(n835)
  );
  //AND U129bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U129bar (
    .O(n837bar),
    .I0(inbar[150]),
    .I1(n835bar)
  );
  //OR U130
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U130 (
    .O(n835),
    .I0(in[172]),
    .I1(in[155])
  );
  //AND U130bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U130bar (
    .O(n835bar),
    .I0(inbar[172]),
    .I1(inbar[155])
  );
  //OR U131
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U131 (
    .O(n893),
    .I0(n834),
    .I1(n833)
  );
  //AND U131bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U131bar (
    .O(n893bar),
    .I0(n834bar),
    .I1(n833bar)
  );
  //OR U132
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U132 (
    .O(n833),
    .I0(n832),
    .I1(n831)
  );
  //AND U132bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U132bar (
    .O(n833bar),
    .I0(n832bar),
    .I1(n831bar)
  );
  //OR U133
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U133 (
    .O(n831),
    .I0(in[196]),
    .I1(in[173])
  );
  //AND U133bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U133bar (
    .O(n831bar),
    .I0(inbar[196]),
    .I1(inbar[173])
  );
  //OR U134
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U134 (
    .O(n832),
    .I0(in[222]),
    .I1(n830)
  );
  //AND U134bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U134bar (
    .O(n832bar),
    .I0(inbar[222]),
    .I1(n830bar)
  );
  //OR U135
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U135 (
    .O(n830),
    .I0(in[227]),
    .I1(in[226])
  );
  //AND U135bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U135bar (
    .O(n830bar),
    .I0(inbar[227]),
    .I1(inbar[226])
  );
  //OR U136
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U136 (
    .O(n834),
    .I0(n829),
    .I1(n828)
  );
  //AND U136bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U136bar (
    .O(n834bar),
    .I0(n829bar),
    .I1(n828bar)
  );
  //OR U137
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U137 (
    .O(n828),
    .I0(in[249]),
    .I1(in[231])
  );
  //AND U137bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U137bar (
    .O(n828bar),
    .I0(inbar[249]),
    .I1(inbar[231])
  );
  //OR U138
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U138 (
    .O(n829),
    .I0(in_28),
    .I1(n827)
  );
  //AND U138bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U138bar (
    .O(n829bar),
    .I0(in_28bar),
    .I1(n827bar)
  );
  //OR U139
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U139 (
    .O(n827),
    .I0(in_52),
    .I1(in_47)
  );
  //AND U139bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U139bar (
    .O(n827bar),
    .I0(in_52bar),
    .I1(in_47bar)
  );
  //OR U140
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U140 (
    .O(out[3]),
    .I0(n826),
    .I1(n825)
  );
  //AND U140bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U140bar (
    .O(outbar[3]),
    .I0(n826bar),
    .I1(n825bar)
  );
  //OR U141
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U141 (
    .O(n825),
    .I0(n824),
    .I1(n823)
  );
  //AND U141bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U141bar (
    .O(n825bar),
    .I0(n824bar),
    .I1(n823bar)
  );
  //OR U142
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U142 (
    .O(n823),
    .I0(n822),
    .I1(n821)
  );
  //AND U142bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U142bar (
    .O(n823bar),
    .I0(n822bar),
    .I1(n821bar)
  );
  //OR U143
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U143 (
    .O(n821),
    .I0(n820),
    .I1(n819)
  );
  //AND U143bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U143bar (
    .O(n821bar),
    .I0(n820bar),
    .I1(n819bar)
  );
  //OR U144
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U144 (
    .O(n822),
    .I0(n964),
    .I1(n818)
  );
  //AND U144bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U144bar (
    .O(n822bar),
    .I0(n964bar),
    .I1(n818bar)
  );
  //OR U145
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U145 (
    .O(n818),
    .I0(in[118]),
    .I1(n817)
  );
  //AND U145bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U145bar (
    .O(n818bar),
    .I0(inbar[118]),
    .I1(n817bar)
  );
  //OR U146
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U146 (
    .O(n964),
    .I0(n816),
    .I1(n815)
  );
  //AND U146bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U146bar (
    .O(n964bar),
    .I0(n816bar),
    .I1(n815bar)
  );
  //OR U147
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U147 (
    .O(n815),
    .I0(n814),
    .I1(n813)
  );
  //AND U147bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U147bar (
    .O(n815bar),
    .I0(n814bar),
    .I1(n813bar)
  );
  //OR U148
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U148 (
    .O(n813),
    .I0(n812),
    .I1(n811)
  );
  //AND U148bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U148bar (
    .O(n813bar),
    .I0(n812bar),
    .I1(n811bar)
  );
  //OR U149
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U149 (
    .O(n811),
    .I0(in[122]),
    .I1(in[111])
  );
  //AND U149bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U149bar (
    .O(n811bar),
    .I0(inbar[122]),
    .I1(inbar[111])
  );
  //OR U150
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U150 (
    .O(n812),
    .I0(in[154]),
    .I1(in[151])
  );
  //AND U150bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U150bar (
    .O(n812bar),
    .I0(inbar[154]),
    .I1(inbar[151])
  );
  //OR U151
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U151 (
    .O(n814),
    .I0(n810),
    .I1(n809)
  );
  //AND U151bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U151bar (
    .O(n814bar),
    .I0(n810bar),
    .I1(n809bar)
  );
  //OR U152
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U152 (
    .O(n809),
    .I0(in[187]),
    .I1(in[177])
  );
  //AND U152bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U152bar (
    .O(n809bar),
    .I0(inbar[187]),
    .I1(inbar[177])
  );
  //OR U153
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U153 (
    .O(n810),
    .I0(in[200]),
    .I1(in[192])
  );
  //AND U153bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U153bar (
    .O(n810bar),
    .I0(inbar[200]),
    .I1(inbar[192])
  );
  //OR U154
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U154 (
    .O(n816),
    .I0(n808),
    .I1(n807)
  );
  //AND U154bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U154bar (
    .O(n816bar),
    .I0(n808bar),
    .I1(n807bar)
  );
  //OR U155
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U155 (
    .O(n807),
    .I0(n806),
    .I1(n805)
  );
  //AND U155bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U155bar (
    .O(n807bar),
    .I0(n806bar),
    .I1(n805bar)
  );
  //OR U156
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U156 (
    .O(n805),
    .I0(in[225]),
    .I1(in[207])
  );
  //AND U156bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U156bar (
    .O(n805bar),
    .I0(inbar[225]),
    .I1(inbar[207])
  );
  //OR U157
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U157 (
    .O(n806),
    .I0(in[98]),
    .I1(in[226])
  );
  //AND U157bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U157bar (
    .O(n806bar),
    .I0(inbar[98]),
    .I1(inbar[226])
  );
  //OR U158
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U158 (
    .O(n808),
    .I0(n804),
    .I1(n803)
  );
  //AND U158bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U158bar (
    .O(n808bar),
    .I0(n804bar),
    .I1(n803bar)
  );
  //OR U159
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U159 (
    .O(n803),
    .I0(in_20),
    .I1(in_16)
  );
  //AND U159bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U159bar (
    .O(n803bar),
    .I0(in_20bar),
    .I1(in_16bar)
  );
  //OR U160
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U160 (
    .O(n804),
    .I0(in_55),
    .I1(in_45)
  );
  //AND U160bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U160bar (
    .O(n804bar),
    .I0(in_55bar),
    .I1(in_45bar)
  );
  //OR U161
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U161 (
    .O(n824),
    .I0(n802),
    .I1(n801)
  );
  //AND U161bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U161bar (
    .O(n824bar),
    .I0(n802bar),
    .I1(n801bar)
  );
  //OR U162
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U162 (
    .O(n801),
    .I0(in[162]),
    .I1(in[149])
  );
  //AND U162bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U162bar (
    .O(n801bar),
    .I0(inbar[162]),
    .I1(inbar[149])
  );
  //OR U163
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U163 (
    .O(n802),
    .I0(in[163]),
    .I1(n800)
  );
  //AND U163bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U163bar (
    .O(n802bar),
    .I0(inbar[163]),
    .I1(n800bar)
  );
  //OR U164
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U164 (
    .O(n800),
    .I0(in[191]),
    .I1(in[189])
  );
  //AND U164bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U164bar (
    .O(n800bar),
    .I0(inbar[191]),
    .I1(inbar[189])
  );
  //OR U165
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U165 (
    .O(n826),
    .I0(n799),
    .I1(n798)
  );
  //AND U165bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U165bar (
    .O(n826bar),
    .I0(n799bar),
    .I1(n798bar)
  );
  //OR U166
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U166 (
    .O(n798),
    .I0(n797),
    .I1(n796)
  );
  //AND U166bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U166bar (
    .O(n798bar),
    .I0(n797bar),
    .I1(n796bar)
  );
  //OR U167
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U167 (
    .O(n796),
    .I0(in[212]),
    .I1(in[193])
  );
  //AND U167bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U167bar (
    .O(n796bar),
    .I0(inbar[212]),
    .I1(inbar[193])
  );
  //OR U168
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U168 (
    .O(n797),
    .I0(in[238]),
    .I1(n795)
  );
  //AND U168bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U168bar (
    .O(n797bar),
    .I0(inbar[238]),
    .I1(n795bar)
  );
  //OR U169
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U169 (
    .O(n795),
    .I0(in[88]),
    .I1(in[247])
  );
  //AND U169bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U169bar (
    .O(n795bar),
    .I0(inbar[88]),
    .I1(inbar[247])
  );
  //OR U170
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U170 (
    .O(n799),
    .I0(n794),
    .I1(n793)
  );
  //AND U170bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U170bar (
    .O(n799bar),
    .I0(n794bar),
    .I1(n793bar)
  );
  //OR U171
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U171 (
    .O(n793),
    .I0(in[94]),
    .I1(in[92])
  );
  //AND U171bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U171bar (
    .O(n793bar),
    .I0(inbar[94]),
    .I1(inbar[92])
  );
  //OR U172
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U172 (
    .O(n794),
    .I0(in_52),
    .I1(n792)
  );
  //AND U172bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U172bar (
    .O(n794bar),
    .I0(in_52bar),
    .I1(n792bar)
  );
  //OR U173
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U173 (
    .O(n792),
    .I0(in_70),
    .I1(in_67)
  );
  //AND U173bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U173bar (
    .O(n792bar),
    .I0(in_70bar),
    .I1(in_67bar)
  );
  //OR U174
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U174 (
    .O(out[2]),
    .I0(n791),
    .I1(n790)
  );
  //AND U174bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U174bar (
    .O(outbar[2]),
    .I0(n791bar),
    .I1(n790bar)
  );
  //OR U175
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U175 (
    .O(n790),
    .I0(n789),
    .I1(n788)
  );
  //AND U175bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U175bar (
    .O(n790bar),
    .I0(n789bar),
    .I1(n788bar)
  );
  //OR U176
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U176 (
    .O(n788),
    .I0(n787),
    .I1(n786)
  );
  //AND U176bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U176bar (
    .O(n788bar),
    .I0(n787bar),
    .I1(n786bar)
  );
  //OR U177
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U177 (
    .O(n786),
    .I0(n819),
    .I1(n785)
  );
  //AND U177bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U177bar (
    .O(n786bar),
    .I0(n819bar),
    .I1(n785bar)
  );
  //OR U178
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U178 (
    .O(n819),
    .I0(n784),
    .I1(n783)
  );
  //AND U178bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U178bar (
    .O(n819bar),
    .I0(n784bar),
    .I1(n783bar)
  );
  //OR U179
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U179 (
    .O(n783),
    .I0(n782),
    .I1(n781)
  );
  //AND U179bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U179bar (
    .O(n783bar),
    .I0(n782bar),
    .I1(n781bar)
  );
  //OR U180
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U180 (
    .O(n781),
    .I0(n780),
    .I1(n779)
  );
  //AND U180bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U180bar (
    .O(n781bar),
    .I0(n780bar),
    .I1(n779bar)
  );
  //OR U181
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U181 (
    .O(n779),
    .I0(n962),
    .I1(n778)
  );
  //AND U181bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U181bar (
    .O(n779bar),
    .I0(n962bar),
    .I1(n778bar)
  );
  //OR U182
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U182 (
    .O(n962),
    .I0(n777),
    .I1(n776)
  );
  //AND U182bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U182bar (
    .O(n962bar),
    .I0(n777bar),
    .I1(n776bar)
  );
  //OR U183
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U183 (
    .O(n776),
    .I0(n775),
    .I1(n774)
  );
  //AND U183bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U183bar (
    .O(n776bar),
    .I0(n775bar),
    .I1(n774bar)
  );
  //OR U184
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U184 (
    .O(n774),
    .I0(n773),
    .I1(n772)
  );
  //AND U184bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U184bar (
    .O(n774bar),
    .I0(n773bar),
    .I1(n772bar)
  );
  //OR U185
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U185 (
    .O(n772),
    .I0(in[131]),
    .I1(in[120])
  );
  //AND U185bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U185bar (
    .O(n772bar),
    .I0(inbar[131]),
    .I1(inbar[120])
  );
  //OR U186
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U186 (
    .O(n773),
    .I0(in[153]),
    .I1(in[147])
  );
  //AND U186bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U186bar (
    .O(n773bar),
    .I0(inbar[153]),
    .I1(inbar[147])
  );
  //OR U187
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U187 (
    .O(n775),
    .I0(n771),
    .I1(n770)
  );
  //AND U187bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U187bar (
    .O(n775bar),
    .I0(n771bar),
    .I1(n770bar)
  );
  //OR U188
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U188 (
    .O(n770),
    .I0(in[170]),
    .I1(in[156])
  );
  //AND U188bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U188bar (
    .O(n770bar),
    .I0(inbar[170]),
    .I1(inbar[156])
  );
  //OR U189
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U189 (
    .O(n771),
    .I0(in[223]),
    .I1(in[190])
  );
  //AND U189bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U189bar (
    .O(n771bar),
    .I0(inbar[223]),
    .I1(inbar[190])
  );
  //OR U190
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U190 (
    .O(n777),
    .I0(n769),
    .I1(n768)
  );
  //AND U190bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U190bar (
    .O(n777bar),
    .I0(n769bar),
    .I1(n768bar)
  );
  //OR U191
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U191 (
    .O(n768),
    .I0(n767),
    .I1(n766)
  );
  //AND U191bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U191bar (
    .O(n768bar),
    .I0(n767bar),
    .I1(n766bar)
  );
  //OR U192
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U192 (
    .O(n766),
    .I0(in[236]),
    .I1(in[230])
  );
  //AND U192bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U192bar (
    .O(n766bar),
    .I0(inbar[236]),
    .I1(inbar[230])
  );
  //OR U193
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U193 (
    .O(n767),
    .I0(in[85]),
    .I1(in[240])
  );
  //AND U193bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U193bar (
    .O(n767bar),
    .I0(inbar[85]),
    .I1(inbar[240])
  );
  //OR U194
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U194 (
    .O(n769),
    .I0(n765),
    .I1(n764)
  );
  //AND U194bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U194bar (
    .O(n769bar),
    .I0(n765bar),
    .I1(n764bar)
  );
  //OR U195
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U195 (
    .O(n764),
    .I0(in_12),
    .I1(in[90])
  );
  //AND U195bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U195bar (
    .O(n764bar),
    .I0(in_12bar),
    .I1(inbar[90])
  );
  //OR U196
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U196 (
    .O(n765),
    .I0(in_39),
    .I1(in_28)
  );
  //AND U196bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U196bar (
    .O(n765bar),
    .I0(in_39bar),
    .I1(in_28bar)
  );
  //OR U197
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U197 (
    .O(n780),
    .I0(in[109]),
    .I1(n763)
  );
  //AND U197bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U197bar (
    .O(n780bar),
    .I0(inbar[109]),
    .I1(n763bar)
  );
  //OR U198
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U198 (
    .O(n782),
    .I0(n762),
    .I1(n761)
  );
  //AND U198bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U198bar (
    .O(n782bar),
    .I0(n762bar),
    .I1(n761bar)
  );
  //OR U199
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U199 (
    .O(n761),
    .I0(in[138]),
    .I1(in[129])
  );
  //AND U199bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U199bar (
    .O(n761bar),
    .I0(inbar[138]),
    .I1(inbar[129])
  );
  //OR U200
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U200 (
    .O(n762),
    .I0(in[157]),
    .I1(n760)
  );
  //AND U200bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U200bar (
    .O(n762bar),
    .I0(inbar[157]),
    .I1(n760bar)
  );
  //OR U201
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U201 (
    .O(n760),
    .I0(in[182]),
    .I1(in[167])
  );
  //AND U201bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U201bar (
    .O(n760bar),
    .I0(inbar[182]),
    .I1(inbar[167])
  );
  //OR U202
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U202 (
    .O(n784),
    .I0(n759),
    .I1(n758)
  );
  //AND U202bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U202bar (
    .O(n784bar),
    .I0(n759bar),
    .I1(n758bar)
  );
  //OR U203
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U203 (
    .O(n758),
    .I0(n757),
    .I1(n756)
  );
  //AND U203bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U203bar (
    .O(n758bar),
    .I0(n757bar),
    .I1(n756bar)
  );
  //OR U204
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U204 (
    .O(n756),
    .I0(in[195]),
    .I1(in[184])
  );
  //AND U204bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U204bar (
    .O(n756bar),
    .I0(inbar[195]),
    .I1(inbar[184])
  );
  //OR U205
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U205 (
    .O(n757),
    .I0(in[196]),
    .I1(n755)
  );
  //AND U205bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U205bar (
    .O(n757bar),
    .I0(inbar[196]),
    .I1(n755bar)
  );
  //OR U206
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U206 (
    .O(n755),
    .I0(in[215]),
    .I1(in[209])
  );
  //AND U206bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U206bar (
    .O(n755bar),
    .I0(inbar[215]),
    .I1(inbar[209])
  );
  //OR U207
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U207 (
    .O(n759),
    .I0(n754),
    .I1(n753)
  );
  //AND U207bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U207bar (
    .O(n759bar),
    .I0(n754bar),
    .I1(n753bar)
  );
  //OR U208
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U208 (
    .O(n753),
    .I0(in[93]),
    .I1(in[233])
  );
  //AND U208bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U208bar (
    .O(n753bar),
    .I0(inbar[93]),
    .I1(inbar[233])
  );
  //OR U209
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U209 (
    .O(n754),
    .I0(in_1),
    .I1(n752)
  );
  //AND U209bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U209bar (
    .O(n754bar),
    .I0(in_1bar),
    .I1(n752bar)
  );
  //OR U210
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U210 (
    .O(n752),
    .I0(in_69),
    .I1(in_66)
  );
  //AND U210bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U210bar (
    .O(n752bar),
    .I0(in_69bar),
    .I1(in_66bar)
  );
  //OR U211
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U211 (
    .O(n787),
    .I0(n966),
    .I1(n751)
  );
  //AND U211bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U211bar (
    .O(n787bar),
    .I0(n966bar),
    .I1(n751bar)
  );
  //OR U212
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U212 (
    .O(n751),
    .I0(in[134]),
    .I1(n750)
  );
  //AND U212bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U212bar (
    .O(n751bar),
    .I0(inbar[134]),
    .I1(n750bar)
  );
  //OR U213
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U213 (
    .O(n966),
    .I0(n749),
    .I1(n748)
  );
  //AND U213bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U213bar (
    .O(n966bar),
    .I0(n749bar),
    .I1(n748bar)
  );
  //OR U214
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U214 (
    .O(n748),
    .I0(n747),
    .I1(n746)
  );
  //AND U214bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U214bar (
    .O(n748bar),
    .I0(n747bar),
    .I1(n746bar)
  );
  //OR U215
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U215 (
    .O(n746),
    .I0(n745),
    .I1(n744)
  );
  //AND U215bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U215bar (
    .O(n746bar),
    .I0(n745bar),
    .I1(n744bar)
  );
  //OR U216
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U216 (
    .O(n744),
    .I0(in[136]),
    .I1(in[121])
  );
  //AND U216bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U216bar (
    .O(n744bar),
    .I0(inbar[136]),
    .I1(inbar[121])
  );
  //OR U217
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U217 (
    .O(n745),
    .I0(in[186]),
    .I1(in[174])
  );
  //AND U217bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U217bar (
    .O(n745bar),
    .I0(inbar[186]),
    .I1(inbar[174])
  );
  //OR U218
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U218 (
    .O(n747),
    .I0(n743),
    .I1(n742)
  );
  //AND U218bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U218bar (
    .O(n747bar),
    .I0(n743bar),
    .I1(n742bar)
  );
  //OR U219
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U219 (
    .O(n742),
    .I0(in[198]),
    .I1(in[197])
  );
  //AND U219bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U219bar (
    .O(n742bar),
    .I0(inbar[198]),
    .I1(inbar[197])
  );
  //OR U220
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U220 (
    .O(n743),
    .I0(in[214]),
    .I1(in[199])
  );
  //AND U220bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U220bar (
    .O(n743bar),
    .I0(inbar[214]),
    .I1(inbar[199])
  );
  //OR U221
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U221 (
    .O(n749),
    .I0(n741),
    .I1(n740)
  );
  //AND U221bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U221bar (
    .O(n749bar),
    .I0(n741bar),
    .I1(n740bar)
  );
  //OR U222
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U222 (
    .O(n740),
    .I0(n739),
    .I1(n738)
  );
  //AND U222bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U222bar (
    .O(n740bar),
    .I0(n739bar),
    .I1(n738bar)
  );
  //OR U223
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U223 (
    .O(n738),
    .I0(in[231]),
    .I1(in[220])
  );
  //AND U223bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U223bar (
    .O(n738bar),
    .I0(inbar[231]),
    .I1(inbar[220])
  );
  //OR U224
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U224 (
    .O(n739),
    .I0(in_25),
    .I1(in[245])
  );
  //AND U224bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U224bar (
    .O(n739bar),
    .I0(in_25bar),
    .I1(inbar[245])
  );
  //OR U225
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U225 (
    .O(n741),
    .I0(n737),
    .I1(n736)
  );
  //AND U225bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U225bar (
    .O(n741bar),
    .I0(n737bar),
    .I1(n736bar)
  );
  //OR U226
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U226 (
    .O(n736),
    .I0(in_53),
    .I1(in_29)
  );
  //AND U226bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U226bar (
    .O(n736bar),
    .I0(in_53bar),
    .I1(in_29bar)
  );
  //OR U227
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U227 (
    .O(n737),
    .I0(in_79),
    .I1(in_74)
  );
  //AND U227bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U227bar (
    .O(n737bar),
    .I0(in_79bar),
    .I1(in_74bar)
  );
  //OR U228
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U228 (
    .O(n789),
    .I0(n735),
    .I1(n734)
  );
  //AND U228bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U228bar (
    .O(n789bar),
    .I0(n735bar),
    .I1(n734bar)
  );
  //OR U229
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U229 (
    .O(n734),
    .I0(in[152]),
    .I1(in[140])
  );
  //AND U229bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U229bar (
    .O(n734bar),
    .I0(inbar[152]),
    .I1(inbar[140])
  );
  //OR U230
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U230 (
    .O(n735),
    .I0(in[155]),
    .I1(n733)
  );
  //AND U230bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U230bar (
    .O(n735bar),
    .I0(inbar[155]),
    .I1(n733bar)
  );
  //OR U231
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U231 (
    .O(n733),
    .I0(in[166]),
    .I1(in[165])
  );
  //AND U231bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U231bar (
    .O(n733bar),
    .I0(inbar[166]),
    .I1(inbar[165])
  );
  //OR U232
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U232 (
    .O(n791),
    .I0(n732),
    .I1(n731)
  );
  //AND U232bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U232bar (
    .O(n791bar),
    .I0(n732bar),
    .I1(n731bar)
  );
  //OR U233
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U233 (
    .O(n731),
    .I0(n730),
    .I1(n729)
  );
  //AND U233bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U233bar (
    .O(n731bar),
    .I0(n730bar),
    .I1(n729bar)
  );
  //OR U234
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U234 (
    .O(n729),
    .I0(in[202]),
    .I1(in[185])
  );
  //AND U234bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U234bar (
    .O(n729bar),
    .I0(inbar[202]),
    .I1(inbar[185])
  );
  //OR U235
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U235 (
    .O(n730),
    .I0(in[211]),
    .I1(n728)
  );
  //AND U235bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U235bar (
    .O(n730bar),
    .I0(inbar[211]),
    .I1(n728bar)
  );
  //OR U236
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U236 (
    .O(n728),
    .I0(in[255]),
    .I1(in[253])
  );
  //AND U236bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U236bar (
    .O(n728bar),
    .I0(inbar[255]),
    .I1(inbar[253])
  );
  //OR U237
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U237 (
    .O(n732),
    .I0(n727),
    .I1(n726)
  );
  //AND U237bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U237bar (
    .O(n732bar),
    .I0(n727bar),
    .I1(n726bar)
  );
  //OR U238
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U238 (
    .O(n726),
    .I0(in_35),
    .I1(in_15)
  );
  //AND U238bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U238bar (
    .O(n726bar),
    .I0(in_35bar),
    .I1(in_15bar)
  );
  //OR U239
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U239 (
    .O(n727),
    .I0(in_36),
    .I1(n725)
  );
  //AND U239bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U239bar (
    .O(n727bar),
    .I0(in_36bar),
    .I1(n725bar)
  );
  //OR U240
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U240 (
    .O(n725),
    .I0(in_48),
    .I1(in_40)
  );
  //AND U240bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U240bar (
    .O(n725bar),
    .I0(in_48bar),
    .I1(in_40bar)
  );
  //OR U241
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U241 (
    .O(out[1]),
    .I0(n724),
    .I1(n723)
  );
  //AND U241bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U241bar (
    .O(outbar[1]),
    .I0(n724bar),
    .I1(n723bar)
  );
  //OR U242
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U242 (
    .O(n723),
    .I0(n722),
    .I1(n721)
  );
  //AND U242bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U242bar (
    .O(n723bar),
    .I0(n722bar),
    .I1(n721bar)
  );
  //OR U243
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U243 (
    .O(n721),
    .I0(n720),
    .I1(n719)
  );
  //AND U243bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U243bar (
    .O(n721bar),
    .I0(n720bar),
    .I1(n719bar)
  );
  //OR U244
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U244 (
    .O(n719),
    .I0(n921),
    .I1(n887)
  );
  //AND U244bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U244bar (
    .O(n719bar),
    .I0(n921bar),
    .I1(n887bar)
  );
  //OR U245
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U245 (
    .O(n887),
    .I0(n718),
    .I1(n717)
  );
  //AND U245bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U245bar (
    .O(n887bar),
    .I0(n718bar),
    .I1(n717bar)
  );
  //OR U246
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U246 (
    .O(n717),
    .I0(n716),
    .I1(n715)
  );
  //AND U246bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U246bar (
    .O(n717bar),
    .I0(n716bar),
    .I1(n715bar)
  );
  //OR U247
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U247 (
    .O(n715),
    .I0(n714),
    .I1(n713)
  );
  //AND U247bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U247bar (
    .O(n715bar),
    .I0(n714bar),
    .I1(n713bar)
  );
  //OR U248
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U248 (
    .O(n713),
    .I0(in[116]),
    .I1(in[110])
  );
  //AND U248bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U248bar (
    .O(n713bar),
    .I0(inbar[116]),
    .I1(inbar[110])
  );
  //OR U249
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U249 (
    .O(n714),
    .I0(in[133]),
    .I1(in[130])
  );
  //AND U249bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U249bar (
    .O(n714bar),
    .I0(inbar[133]),
    .I1(inbar[130])
  );
  //OR U250
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U250 (
    .O(n716),
    .I0(n712),
    .I1(n711)
  );
  //AND U250bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U250bar (
    .O(n716bar),
    .I0(n712bar),
    .I1(n711bar)
  );
  //OR U251
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U251 (
    .O(n711),
    .I0(in[203]),
    .I1(in[135])
  );
  //AND U251bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U251bar (
    .O(n711bar),
    .I0(inbar[203]),
    .I1(inbar[135])
  );
  //OR U252
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U252 (
    .O(n712),
    .I0(in[232]),
    .I1(in[223])
  );
  //AND U252bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U252bar (
    .O(n712bar),
    .I0(inbar[232]),
    .I1(inbar[223])
  );
  //OR U253
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U253 (
    .O(n718),
    .I0(n710),
    .I1(n709)
  );
  //AND U253bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U253bar (
    .O(n718bar),
    .I0(n710bar),
    .I1(n709bar)
  );
  //OR U254
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U254 (
    .O(n709),
    .I0(n708),
    .I1(n707)
  );
  //AND U254bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U254bar (
    .O(n709bar),
    .I0(n708bar),
    .I1(n707bar)
  );
  //OR U255
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U255 (
    .O(n707),
    .I0(in[255]),
    .I1(in[233])
  );
  //AND U255bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U255bar (
    .O(n707bar),
    .I0(inbar[255]),
    .I1(inbar[233])
  );
  //OR U256
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U256 (
    .O(n708),
    .I0(in_53),
    .I1(in_34)
  );
  //AND U256bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U256bar (
    .O(n708bar),
    .I0(in_53bar),
    .I1(in_34bar)
  );
  //OR U257
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U257 (
    .O(n710),
    .I0(n706),
    .I1(n705)
  );
  //AND U257bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U257bar (
    .O(n710bar),
    .I0(n706bar),
    .I1(n705bar)
  );
  //OR U258
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U258 (
    .O(n705),
    .I0(in_57),
    .I1(in_55)
  );
  //AND U258bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U258bar (
    .O(n705bar),
    .I0(in_57bar),
    .I1(in_55bar)
  );
  //OR U259
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U259 (
    .O(n706),
    .I0(in_68),
    .I1(in_67)
  );
  //AND U259bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U259bar (
    .O(n706bar),
    .I0(in_68bar),
    .I1(in_67bar)
  );
  //OR U260
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U260 (
    .O(n921),
    .I0(n704),
    .I1(n703)
  );
  //AND U260bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U260bar (
    .O(n921bar),
    .I0(n704bar),
    .I1(n703bar)
  );
  //OR U261
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U261 (
    .O(n703),
    .I0(n702),
    .I1(n701)
  );
  //AND U261bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U261bar (
    .O(n703bar),
    .I0(n702bar),
    .I1(n701bar)
  );
  //OR U262
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U262 (
    .O(n701),
    .I0(n700),
    .I1(n699)
  );
  //AND U262bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U262bar (
    .O(n701bar),
    .I0(n700bar),
    .I1(n699bar)
  );
  //OR U263
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U263 (
    .O(n699),
    .I0(n944),
    .I1(n872)
  );
  //AND U263bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U263bar (
    .O(n699bar),
    .I0(n944bar),
    .I1(n872bar)
  );
  //OR U264
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U264 (
    .O(n872),
    .I0(n698),
    .I1(n697)
  );
  //AND U264bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U264bar (
    .O(n872bar),
    .I0(n698bar),
    .I1(n697bar)
  );
  //OR U265
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U265 (
    .O(n697),
    .I0(n696),
    .I1(n695)
  );
  //AND U265bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U265bar (
    .O(n697bar),
    .I0(n696bar),
    .I1(n695bar)
  );
  //OR U266
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U266 (
    .O(n695),
    .I0(n694),
    .I1(n693)
  );
  //AND U266bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U266bar (
    .O(n695bar),
    .I0(n694bar),
    .I1(n693bar)
  );
  //OR U267
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U267 (
    .O(n693),
    .I0(in[121]),
    .I1(in[102])
  );
  //AND U267bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U267bar (
    .O(n693bar),
    .I0(inbar[121]),
    .I1(inbar[102])
  );
  //OR U268
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U268 (
    .O(n694),
    .I0(in[162]),
    .I1(in[161])
  );
  //AND U268bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U268bar (
    .O(n694bar),
    .I0(inbar[162]),
    .I1(inbar[161])
  );
  //OR U269
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U269 (
    .O(n696),
    .I0(n692),
    .I1(n691)
  );
  //AND U269bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U269bar (
    .O(n696bar),
    .I0(n692bar),
    .I1(n691bar)
  );
  //OR U270
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U270 (
    .O(n691),
    .I0(in[192]),
    .I1(in[178])
  );
  //AND U270bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U270bar (
    .O(n691bar),
    .I0(inbar[192]),
    .I1(inbar[178])
  );
  //OR U271
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U271 (
    .O(n692),
    .I0(in[244]),
    .I1(in[209])
  );
  //AND U271bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U271bar (
    .O(n692bar),
    .I0(inbar[244]),
    .I1(inbar[209])
  );
  //OR U272
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U272 (
    .O(n698),
    .I0(n690),
    .I1(n689)
  );
  //AND U272bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U272bar (
    .O(n698bar),
    .I0(n690bar),
    .I1(n689bar)
  );
  //OR U273
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U273 (
    .O(n689),
    .I0(n688),
    .I1(n687)
  );
  //AND U273bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U273bar (
    .O(n689bar),
    .I0(n688bar),
    .I1(n687bar)
  );
  //OR U274
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U274 (
    .O(n687),
    .I0(in[90]),
    .I1(in[254])
  );
  //AND U274bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U274bar (
    .O(n687bar),
    .I0(inbar[90]),
    .I1(inbar[254])
  );
  //OR U275
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U275 (
    .O(n688),
    .I0(in_36),
    .I1(in_32)
  );
  //AND U275bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U275bar (
    .O(n688bar),
    .I0(in_36bar),
    .I1(in_32bar)
  );
  //OR U276
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U276 (
    .O(n690),
    .I0(n686),
    .I1(n685)
  );
  //AND U276bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U276bar (
    .O(n690bar),
    .I0(n686bar),
    .I1(n685bar)
  );
  //OR U277
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U277 (
    .O(n685),
    .I0(in_62),
    .I1(in_37)
  );
  //AND U277bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U277bar (
    .O(n685bar),
    .I0(in_62bar),
    .I1(in_37bar)
  );
  //OR U278
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U278 (
    .O(n686),
    .I0(in_75),
    .I1(in_73)
  );
  //AND U278bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U278bar (
    .O(n686bar),
    .I0(in_75bar),
    .I1(in_73bar)
  );
  //OR U279
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U279 (
    .O(n944),
    .I0(n684),
    .I1(n683)
  );
  //AND U279bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U279bar (
    .O(n944bar),
    .I0(n684bar),
    .I1(n683bar)
  );
  //OR U280
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U280 (
    .O(n683),
    .I0(n682),
    .I1(n681)
  );
  //AND U280bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U280bar (
    .O(n683bar),
    .I0(n682bar),
    .I1(n681bar)
  );
  //OR U281
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U281 (
    .O(n681),
    .I0(n680),
    .I1(n679)
  );
  //AND U281bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U281bar (
    .O(n681bar),
    .I0(n680bar),
    .I1(n679bar)
  );
  //OR U282
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U282 (
    .O(n679),
    .I0(in[171]),
    .I1(in[153])
  );
  //AND U282bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U282bar (
    .O(n679bar),
    .I0(inbar[171]),
    .I1(inbar[153])
  );
  //OR U283
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U283 (
    .O(n680),
    .I0(in[187]),
    .I1(in[176])
  );
  //AND U283bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U283bar (
    .O(n680bar),
    .I0(inbar[187]),
    .I1(inbar[176])
  );
  //OR U284
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U284 (
    .O(n682),
    .I0(n678),
    .I1(n677)
  );
  //AND U284bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U284bar (
    .O(n682bar),
    .I0(n678bar),
    .I1(n677bar)
  );
  //OR U285
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U285 (
    .O(n677),
    .I0(in[245]),
    .I1(in[211])
  );
  //AND U285bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U285bar (
    .O(n677bar),
    .I0(inbar[245]),
    .I1(inbar[211])
  );
  //OR U286
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U286 (
    .O(n678),
    .I0(in[97]),
    .I1(in[88])
  );
  //AND U286bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U286bar (
    .O(n678bar),
    .I0(inbar[97]),
    .I1(inbar[88])
  );
  //OR U287
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U287 (
    .O(n684),
    .I0(n676),
    .I1(n675)
  );
  //AND U287bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U287bar (
    .O(n684bar),
    .I0(n676bar),
    .I1(n675bar)
  );
  //OR U288
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U288 (
    .O(n675),
    .I0(n674),
    .I1(n673)
  );
  //AND U288bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U288bar (
    .O(n675bar),
    .I0(n674bar),
    .I1(n673bar)
  );
  //OR U289
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U289 (
    .O(n673),
    .I0(in_10),
    .I1(in_0)
  );
  //AND U289bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U289bar (
    .O(n673bar),
    .I0(in_10bar),
    .I1(in_0bar)
  );
  //OR U290
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U290 (
    .O(n674),
    .I0(in_59),
    .I1(in_5)
  );
  //AND U290bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U290bar (
    .O(n674bar),
    .I0(in_59bar),
    .I1(in_5bar)
  );
  //OR U291
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U291 (
    .O(n676),
    .I0(n672),
    .I1(n671)
  );
  //AND U291bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U291bar (
    .O(n676bar),
    .I0(n672bar),
    .I1(n671bar)
  );
  //OR U292
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U292 (
    .O(n671),
    .I0(in_60),
    .I1(in_6)
  );
  //AND U292bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U292bar (
    .O(n671bar),
    .I0(in_60bar),
    .I1(in_6bar)
  );
  //OR U293
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U293 (
    .O(n672),
    .I0(in_77),
    .I1(in_69)
  );
  //AND U293bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U293bar (
    .O(n672bar),
    .I0(in_77bar),
    .I1(in_69bar)
  );
  //OR U294
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U294 (
    .O(n700),
    .I0(in[113]),
    .I1(n864)
  );
  //AND U294bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U294bar (
    .O(n700bar),
    .I0(inbar[113]),
    .I1(n864bar)
  );
  //OR U295
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U295 (
    .O(n864),
    .I0(n670),
    .I1(n669)
  );
  //AND U295bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U295bar (
    .O(n864bar),
    .I0(n670bar),
    .I1(n669bar)
  );
  //OR U296
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U296 (
    .O(n669),
    .I0(n668),
    .I1(n667)
  );
  //AND U296bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U296bar (
    .O(n669bar),
    .I0(n668bar),
    .I1(n667bar)
  );
  //OR U297
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U297 (
    .O(n667),
    .I0(n666),
    .I1(n665)
  );
  //AND U297bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U297bar (
    .O(n667bar),
    .I0(n666bar),
    .I1(n665bar)
  );
  //OR U298
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U298 (
    .O(n665),
    .I0(in[125]),
    .I1(in[107])
  );
  //AND U298bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U298bar (
    .O(n665bar),
    .I0(inbar[125]),
    .I1(inbar[107])
  );
  //OR U299
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U299 (
    .O(n666),
    .I0(in[138]),
    .I1(in[126])
  );
  //AND U299bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U299bar (
    .O(n666bar),
    .I0(inbar[138]),
    .I1(inbar[126])
  );
  //OR U300
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U300 (
    .O(n668),
    .I0(n664),
    .I1(n663)
  );
  //AND U300bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U300bar (
    .O(n668bar),
    .I0(n664bar),
    .I1(n663bar)
  );
  //OR U301
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U301 (
    .O(n663),
    .I0(in[189]),
    .I1(in[143])
  );
  //AND U301bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U301bar (
    .O(n663bar),
    .I0(inbar[189]),
    .I1(inbar[143])
  );
  //OR U302
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U302 (
    .O(n664),
    .I0(in[99]),
    .I1(in[214])
  );
  //AND U302bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U302bar (
    .O(n664bar),
    .I0(inbar[99]),
    .I1(inbar[214])
  );
  //OR U303
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U303 (
    .O(n670),
    .I0(n662),
    .I1(n661)
  );
  //AND U303bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U303bar (
    .O(n670bar),
    .I0(n662bar),
    .I1(n661bar)
  );
  //OR U304
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U304 (
    .O(n661),
    .I0(n660),
    .I1(n659)
  );
  //AND U304bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U304bar (
    .O(n661bar),
    .I0(n660bar),
    .I1(n659bar)
  );
  //OR U305
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U305 (
    .O(n659),
    .I0(in_15),
    .I1(in_12)
  );
  //AND U305bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U305bar (
    .O(n659bar),
    .I0(in_15bar),
    .I1(in_12bar)
  );
  //OR U306
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U306 (
    .O(n660),
    .I0(in_20),
    .I1(in_2)
  );
  //AND U306bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U306bar (
    .O(n660bar),
    .I0(in_20bar),
    .I1(in_2bar)
  );
  //OR U307
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U307 (
    .O(n662),
    .I0(n658),
    .I1(n657)
  );
  //AND U307bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U307bar (
    .O(n662bar),
    .I0(n658bar),
    .I1(n657bar)
  );
  //OR U308
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U308 (
    .O(n657),
    .I0(in_30),
    .I1(in_3)
  );
  //AND U308bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U308bar (
    .O(n657bar),
    .I0(in_30bar),
    .I1(in_3bar)
  );
  //OR U309
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U309 (
    .O(n658),
    .I0(in_4),
    .I1(in_38)
  );
  //AND U309bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U309bar (
    .O(n658bar),
    .I0(in_4bar),
    .I1(in_38bar)
  );
  //OR U310
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U310 (
    .O(n702),
    .I0(n656),
    .I1(n655)
  );
  //AND U310bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U310bar (
    .O(n702bar),
    .I0(n656bar),
    .I1(n655bar)
  );
  //OR U311
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U311 (
    .O(n655),
    .I0(in[148]),
    .I1(in[137])
  );
  //AND U311bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U311bar (
    .O(n655bar),
    .I0(inbar[148]),
    .I1(inbar[137])
  );
  //OR U312
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U312 (
    .O(n656),
    .I0(in[149]),
    .I1(n654)
  );
  //AND U312bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U312bar (
    .O(n656bar),
    .I0(inbar[149]),
    .I1(n654bar)
  );
  //OR U313
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U313 (
    .O(n654),
    .I0(in[195]),
    .I1(in[190])
  );
  //AND U313bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U313bar (
    .O(n654bar),
    .I0(inbar[195]),
    .I1(inbar[190])
  );
  //OR U314
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U314 (
    .O(n704),
    .I0(n653),
    .I1(n652)
  );
  //AND U314bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U314bar (
    .O(n704bar),
    .I0(n653bar),
    .I1(n652bar)
  );
  //OR U315
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U315 (
    .O(n652),
    .I0(n651),
    .I1(n650)
  );
  //AND U315bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U315bar (
    .O(n652bar),
    .I0(n651bar),
    .I1(n650bar)
  );
  //OR U316
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U316 (
    .O(n650),
    .I0(in[98]),
    .I1(in[197])
  );
  //AND U316bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U316bar (
    .O(n650bar),
    .I0(inbar[98]),
    .I1(inbar[197])
  );
  //OR U317
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U317 (
    .O(n651),
    .I0(in_11),
    .I1(n649)
  );
  //AND U317bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U317bar (
    .O(n651bar),
    .I0(in_11bar),
    .I1(n649bar)
  );
  //OR U318
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U318 (
    .O(n649),
    .I0(in_26),
    .I1(in_14)
  );
  //AND U318bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U318bar (
    .O(n649bar),
    .I0(in_26bar),
    .I1(in_14bar)
  );
  //OR U319
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U319 (
    .O(n653),
    .I0(n648),
    .I1(n647)
  );
  //AND U319bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U319bar (
    .O(n653bar),
    .I0(n648bar),
    .I1(n647bar)
  );
  //OR U320
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U320 (
    .O(n647),
    .I0(in_35),
    .I1(in_27)
  );
  //AND U320bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U320bar (
    .O(n647bar),
    .I0(in_35bar),
    .I1(in_27bar)
  );
  //OR U321
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U321 (
    .O(n648),
    .I0(in_50),
    .I1(n646)
  );
  //AND U321bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U321bar (
    .O(n648bar),
    .I0(in_50bar),
    .I1(n646bar)
  );
  //OR U322
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U322 (
    .O(n646),
    .I0(in_78),
    .I1(in_61)
  );
  //AND U322bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U322bar (
    .O(n646bar),
    .I0(in_78bar),
    .I1(in_61bar)
  );
  //OR U323
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U323 (
    .O(n720),
    .I0(n942),
    .I1(n645)
  );
  //AND U323bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U323bar (
    .O(n720bar),
    .I0(n942bar),
    .I1(n645bar)
  );
  //OR U324
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U324 (
    .O(n645),
    .I0(in[106]),
    .I1(n863)
  );
  //AND U324bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U324bar (
    .O(n645bar),
    .I0(inbar[106]),
    .I1(n863bar)
  );
  //OR U325
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U325 (
    .O(n863),
    .I0(n644),
    .I1(n643)
  );
  //AND U325bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U325bar (
    .O(n863bar),
    .I0(n644bar),
    .I1(n643bar)
  );
  //OR U326
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U326 (
    .O(n643),
    .I0(n642),
    .I1(n641)
  );
  //AND U326bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U326bar (
    .O(n643bar),
    .I0(n642bar),
    .I1(n641bar)
  );
  //OR U327
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U327 (
    .O(n641),
    .I0(n640),
    .I1(n639)
  );
  //AND U327bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U327bar (
    .O(n641bar),
    .I0(n640bar),
    .I1(n639bar)
  );
  //OR U328
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U328 (
    .O(n639),
    .I0(in[127]),
    .I1(in[122])
  );
  //AND U328bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U328bar (
    .O(n639bar),
    .I0(inbar[127]),
    .I1(inbar[122])
  );
  //OR U329
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U329 (
    .O(n640),
    .I0(in[156]),
    .I1(in[132])
  );
  //AND U329bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U329bar (
    .O(n640bar),
    .I0(inbar[156]),
    .I1(inbar[132])
  );
  //OR U330
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U330 (
    .O(n642),
    .I0(n638),
    .I1(n637)
  );
  //AND U330bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U330bar (
    .O(n642bar),
    .I0(n638bar),
    .I1(n637bar)
  );
  //OR U331
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U331 (
    .O(n637),
    .I0(in[159]),
    .I1(in[157])
  );
  //AND U331bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U331bar (
    .O(n637bar),
    .I0(inbar[159]),
    .I1(inbar[157])
  );
  //OR U332
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U332 (
    .O(n638),
    .I0(in[185]),
    .I1(in[169])
  );
  //AND U332bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U332bar (
    .O(n638bar),
    .I0(inbar[185]),
    .I1(inbar[169])
  );
  //OR U333
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U333 (
    .O(n644),
    .I0(n636),
    .I1(n635)
  );
  //AND U333bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U333bar (
    .O(n644bar),
    .I0(n636bar),
    .I1(n635bar)
  );
  //OR U334
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U334 (
    .O(n635),
    .I0(n634),
    .I1(n633)
  );
  //AND U334bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U334bar (
    .O(n635bar),
    .I0(n634bar),
    .I1(n633bar)
  );
  //OR U335
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U335 (
    .O(n633),
    .I0(in[239]),
    .I1(in[218])
  );
  //AND U335bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U335bar (
    .O(n633bar),
    .I0(inbar[239]),
    .I1(inbar[218])
  );
  //OR U336
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U336 (
    .O(n634),
    .I0(in_13),
    .I1(in[87])
  );
  //AND U336bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U336bar (
    .O(n634bar),
    .I0(in_13bar),
    .I1(inbar[87])
  );
  //OR U337
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U337 (
    .O(n636),
    .I0(n632),
    .I1(n631)
  );
  //AND U337bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U337bar (
    .O(n636bar),
    .I0(n632bar),
    .I1(n631bar)
  );
  //OR U338
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U338 (
    .O(n631),
    .I0(in_72),
    .I1(in_70)
  );
  //AND U338bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U338bar (
    .O(n631bar),
    .I0(in_72bar),
    .I1(in_70bar)
  );
  //OR U339
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U339 (
    .O(n632),
    .I0(in_80),
    .I1(in_74)
  );
  //AND U339bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U339bar (
    .O(n632bar),
    .I0(in_80bar),
    .I1(in_74bar)
  );
  //OR U340
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U340 (
    .O(n942),
    .I0(n630),
    .I1(n629)
  );
  //AND U340bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U340bar (
    .O(n942bar),
    .I0(n630bar),
    .I1(n629bar)
  );
  //OR U341
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U341 (
    .O(n629),
    .I0(n628),
    .I1(n627)
  );
  //AND U341bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U341bar (
    .O(n629bar),
    .I0(n628bar),
    .I1(n627bar)
  );
  //OR U342
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U342 (
    .O(n627),
    .I0(n626),
    .I1(n625)
  );
  //AND U342bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U342bar (
    .O(n627bar),
    .I0(n626bar),
    .I1(n625bar)
  );
  //OR U343
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U343 (
    .O(n625),
    .I0(in[146]),
    .I1(in[100])
  );
  //AND U343bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U343bar (
    .O(n625bar),
    .I0(inbar[146]),
    .I1(inbar[100])
  );
  //OR U344
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U344 (
    .O(n626),
    .I0(in[168]),
    .I1(in[152])
  );
  //AND U344bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U344bar (
    .O(n626bar),
    .I0(inbar[168]),
    .I1(inbar[152])
  );
  //OR U345
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U345 (
    .O(n628),
    .I0(n624),
    .I1(n623)
  );
  //AND U345bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U345bar (
    .O(n628bar),
    .I0(n624bar),
    .I1(n623bar)
  );
  //OR U346
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U346 (
    .O(n623),
    .I0(in[199]),
    .I1(in[182])
  );
  //AND U346bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U346bar (
    .O(n623bar),
    .I0(inbar[199]),
    .I1(inbar[182])
  );
  //OR U347
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U347 (
    .O(n624),
    .I0(in[236]),
    .I1(in[204])
  );
  //AND U347bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U347bar (
    .O(n624bar),
    .I0(inbar[236]),
    .I1(inbar[204])
  );
  //OR U348
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U348 (
    .O(n630),
    .I0(n622),
    .I1(n621)
  );
  //AND U348bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U348bar (
    .O(n630bar),
    .I0(n622bar),
    .I1(n621bar)
  );
  //OR U349
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U349 (
    .O(n621),
    .I0(n620),
    .I1(n619)
  );
  //AND U349bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U349bar (
    .O(n621bar),
    .I0(n620bar),
    .I1(n619bar)
  );
  //OR U350
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U350 (
    .O(n619),
    .I0(in[89]),
    .I1(in[246])
  );
  //AND U350bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U350bar (
    .O(n619bar),
    .I0(inbar[89]),
    .I1(inbar[246])
  );
  //OR U351
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U351 (
    .O(n620),
    .I0(in[95]),
    .I1(in[92])
  );
  //AND U351bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U351bar (
    .O(n620bar),
    .I0(inbar[95]),
    .I1(inbar[92])
  );
  //OR U352
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U352 (
    .O(n622),
    .I0(n618),
    .I1(n617)
  );
  //AND U352bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U352bar (
    .O(n622bar),
    .I0(n618bar),
    .I1(n617bar)
  );
  //OR U353
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U353 (
    .O(n617),
    .I0(in_22),
    .I1(in_16)
  );
  //AND U353bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U353bar (
    .O(n617bar),
    .I0(in_22bar),
    .I1(in_16bar)
  );
  //OR U354
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U354 (
    .O(n618),
    .I0(in_51),
    .I1(in_49)
  );
  //AND U354bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U354bar (
    .O(n618bar),
    .I0(in_51bar),
    .I1(in_49bar)
  );
  //OR U355
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U355 (
    .O(n722),
    .I0(n616),
    .I1(n615)
  );
  //AND U355bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U355bar (
    .O(n722bar),
    .I0(n616bar),
    .I1(n615bar)
  );
  //OR U356
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U356 (
    .O(n615),
    .I0(in[158]),
    .I1(in[115])
  );
  //AND U356bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U356bar (
    .O(n615bar),
    .I0(inbar[158]),
    .I1(inbar[115])
  );
  //OR U357
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U357 (
    .O(n616),
    .I0(in[163]),
    .I1(n614)
  );
  //AND U357bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U357bar (
    .O(n616bar),
    .I0(inbar[163]),
    .I1(n614bar)
  );
  //OR U358
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U358 (
    .O(n614),
    .I0(in[206]),
    .I1(in[165])
  );
  //AND U358bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U358bar (
    .O(n614bar),
    .I0(inbar[206]),
    .I1(inbar[165])
  );
  //OR U359
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U359 (
    .O(n724),
    .I0(n613),
    .I1(n612)
  );
  //AND U359bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U359bar (
    .O(n724bar),
    .I0(n613bar),
    .I1(n612bar)
  );
  //OR U360
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U360 (
    .O(n612),
    .I0(n611),
    .I1(n610)
  );
  //AND U360bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U360bar (
    .O(n612bar),
    .I0(n611bar),
    .I1(n610bar)
  );
  //OR U361
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U361 (
    .O(n610),
    .I0(in[213]),
    .I1(in[207])
  );
  //AND U361bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U361bar (
    .O(n610bar),
    .I0(inbar[213]),
    .I1(inbar[207])
  );
  //OR U362
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U362 (
    .O(n611),
    .I0(in[215]),
    .I1(n609)
  );
  //AND U362bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U362bar (
    .O(n611bar),
    .I0(inbar[215]),
    .I1(n609bar)
  );
  //OR U363
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U363 (
    .O(n609),
    .I0(in[230]),
    .I1(in[220])
  );
  //AND U363bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U363bar (
    .O(n609bar),
    .I0(inbar[230]),
    .I1(inbar[220])
  );
  //OR U364
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U364 (
    .O(n613),
    .I0(n608),
    .I1(n607)
  );
  //AND U364bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U364bar (
    .O(n613bar),
    .I0(n608bar),
    .I1(n607bar)
  );
  //OR U365
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U365 (
    .O(n607),
    .I0(in[251]),
    .I1(in[234])
  );
  //AND U365bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U365bar (
    .O(n607bar),
    .I0(inbar[251]),
    .I1(inbar[234])
  );
  //OR U366
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U366 (
    .O(n608),
    .I0(in_17),
    .I1(n606)
  );
  //AND U366bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U366bar (
    .O(n608bar),
    .I0(in_17bar),
    .I1(n606bar)
  );
  //OR U367
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U367 (
    .O(n606),
    .I0(in_65),
    .I1(in_56)
  );
  //AND U367bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U367bar (
    .O(n606bar),
    .I0(in_65bar),
    .I1(in_56bar)
  );
  //OR U368
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U368 (
    .O(out[0]),
    .I0(n605),
    .I1(n604)
  );
  //AND U368bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U368bar (
    .O(outbar[0]),
    .I0(n605bar),
    .I1(n604bar)
  );
  //OR U369
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U369 (
    .O(n604),
    .I0(n603),
    .I1(n602)
  );
  //AND U369bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U369bar (
    .O(n604bar),
    .I0(n603bar),
    .I1(n602bar)
  );
  //OR U370
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U370 (
    .O(n602),
    .I0(n601),
    .I1(n600)
  );
  //AND U370bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U370bar (
    .O(n602bar),
    .I0(n601bar),
    .I1(n600bar)
  );
  //OR U371
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U371 (
    .O(n600),
    .I0(n820),
    .I1(n785)
  );
  //AND U371bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U371bar (
    .O(n600bar),
    .I0(n820bar),
    .I1(n785bar)
  );
  //OR U372
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U372 (
    .O(n785),
    .I0(n599),
    .I1(n598)
  );
  //AND U372bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U372bar (
    .O(n785bar),
    .I0(n599bar),
    .I1(n598bar)
  );
  //OR U373
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U373 (
    .O(n598),
    .I0(n597),
    .I1(n596)
  );
  //AND U373bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U373bar (
    .O(n598bar),
    .I0(n597bar),
    .I1(n596bar)
  );
  //OR U374
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U374 (
    .O(n596),
    .I0(n595),
    .I1(n594)
  );
  //AND U374bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U374bar (
    .O(n596bar),
    .I0(n595bar),
    .I1(n594bar)
  );
  //OR U375
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U375 (
    .O(n594),
    .I0(in[135]),
    .I1(in[104])
  );
  //AND U375bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U375bar (
    .O(n594bar),
    .I0(inbar[135]),
    .I1(inbar[104])
  );
  //OR U376
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U376 (
    .O(n595),
    .I0(in[188]),
    .I1(in[178])
  );
  //AND U376bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U376bar (
    .O(n595bar),
    .I0(inbar[188]),
    .I1(inbar[178])
  );
  //OR U377
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U377 (
    .O(n597),
    .I0(n593),
    .I1(n592)
  );
  //AND U377bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U377bar (
    .O(n597bar),
    .I0(n593bar),
    .I1(n592bar)
  );
  //OR U378
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U378 (
    .O(n592),
    .I0(in[217]),
    .I1(in[194])
  );
  //AND U378bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U378bar (
    .O(n592bar),
    .I0(inbar[217]),
    .I1(inbar[194])
  );
  //OR U379
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U379 (
    .O(n593),
    .I0(in[237]),
    .I1(in[218])
  );
  //AND U379bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U379bar (
    .O(n593bar),
    .I0(inbar[237]),
    .I1(inbar[218])
  );
  //OR U380
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U380 (
    .O(n599),
    .I0(n591),
    .I1(n590)
  );
  //AND U380bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U380bar (
    .O(n599bar),
    .I0(n591bar),
    .I1(n590bar)
  );
  //OR U381
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U381 (
    .O(n590),
    .I0(n589),
    .I1(n588)
  );
  //AND U381bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U381bar (
    .O(n590bar),
    .I0(n589bar),
    .I1(n588bar)
  );
  //OR U382
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U382 (
    .O(n588),
    .I0(in_2),
    .I1(in_10)
  );
  //AND U382bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U382bar (
    .O(n588bar),
    .I0(in_2bar),
    .I1(in_10bar)
  );
  //OR U383
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U383 (
    .O(n589),
    .I0(in_47),
    .I1(in_22)
  );
  //AND U383bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U383bar (
    .O(n589bar),
    .I0(in_47bar),
    .I1(in_22bar)
  );
  //OR U384
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U384 (
    .O(n591),
    .I0(n587),
    .I1(n586)
  );
  //AND U384bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U384bar (
    .O(n591bar),
    .I0(n587bar),
    .I1(n586bar)
  );
  //OR U385
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U385 (
    .O(n586),
    .I0(in_56),
    .I1(in_54)
  );
  //AND U385bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U385bar (
    .O(n586bar),
    .I0(in_56bar),
    .I1(in_54bar)
  );
  //OR U386
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U386 (
    .O(n587),
    .I0(in_63),
    .I1(in_61)
  );
  //AND U386bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U386bar (
    .O(n587bar),
    .I0(in_63bar),
    .I1(in_61bar)
  );
  //OR U387
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U387 (
    .O(n820),
    .I0(n585),
    .I1(n584)
  );
  //AND U387bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U387bar (
    .O(n820bar),
    .I0(n585bar),
    .I1(n584bar)
  );
  //OR U388
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U388 (
    .O(n584),
    .I0(n583),
    .I1(n582)
  );
  //AND U388bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U388bar (
    .O(n584bar),
    .I0(n583bar),
    .I1(n582bar)
  );
  //OR U389
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U389 (
    .O(n582),
    .I0(n581),
    .I1(n580)
  );
  //AND U389bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U389bar (
    .O(n582bar),
    .I0(n581bar),
    .I1(n580bar)
  );
  //OR U390
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U390 (
    .O(n580),
    .I0(in[158]),
    .I1(in[142])
  );
  //AND U390bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U390bar (
    .O(n580bar),
    .I0(inbar[158]),
    .I1(inbar[142])
  );
  //OR U391
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U391 (
    .O(n581),
    .I0(in[175]),
    .I1(in[164])
  );
  //AND U391bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U391bar (
    .O(n581bar),
    .I0(inbar[175]),
    .I1(inbar[164])
  );
  //OR U392
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U392 (
    .O(n583),
    .I0(n579),
    .I1(n578)
  );
  //AND U392bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U392bar (
    .O(n583bar),
    .I0(n579bar),
    .I1(n578bar)
  );
  //OR U393
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U393 (
    .O(n578),
    .I0(in[228]),
    .I1(in[204])
  );
  //AND U393bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U393bar (
    .O(n578bar),
    .I0(inbar[228]),
    .I1(inbar[204])
  );
  //OR U394
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U394 (
    .O(n579),
    .I0(in[91]),
    .I1(in[87])
  );
  //AND U394bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U394bar (
    .O(n579bar),
    .I0(inbar[91]),
    .I1(inbar[87])
  );
  //OR U395
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U395 (
    .O(n585),
    .I0(n577),
    .I1(n576)
  );
  //AND U395bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U395bar (
    .O(n585bar),
    .I0(n577bar),
    .I1(n576bar)
  );
  //OR U396
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U396 (
    .O(n576),
    .I0(n575),
    .I1(n574)
  );
  //AND U396bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U396bar (
    .O(n576bar),
    .I0(n575bar),
    .I1(n574bar)
  );
  //OR U397
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U397 (
    .O(n574),
    .I0(in_21),
    .I1(in_11)
  );
  //AND U397bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U397bar (
    .O(n574bar),
    .I0(in_21bar),
    .I1(in_11bar)
  );
  //OR U398
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U398 (
    .O(n575),
    .I0(in_5),
    .I1(in_3)
  );
  //AND U398bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U398bar (
    .O(n575bar),
    .I0(in_5bar),
    .I1(in_3bar)
  );
  //OR U399
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U399 (
    .O(n577),
    .I0(n573),
    .I1(n572)
  );
  //AND U399bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U399bar (
    .O(n577bar),
    .I0(n573bar),
    .I1(n572bar)
  );
  //OR U400
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U400 (
    .O(n572),
    .I0(in_68),
    .I1(in_64)
  );
  //AND U400bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U400bar (
    .O(n572bar),
    .I0(in_68bar),
    .I1(in_64bar)
  );
  //OR U401
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U401 (
    .O(n573),
    .I0(in_76),
    .I1(in_73)
  );
  //AND U401bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U401bar (
    .O(n573bar),
    .I0(in_76bar),
    .I1(in_73bar)
  );
  //OR U402
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U402 (
    .O(n601),
    .I0(n778),
    .I1(n571)
  );
  //AND U402bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U402bar (
    .O(n601bar),
    .I0(n778bar),
    .I1(n571bar)
  );
  //OR U403
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U403 (
    .O(n571),
    .I0(in[100]),
    .I1(n965)
  );
  //AND U403bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U403bar (
    .O(n571bar),
    .I0(inbar[100]),
    .I1(n965bar)
  );
  //OR U404
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U404 (
    .O(n965),
    .I0(n570),
    .I1(n569)
  );
  //AND U404bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U404bar (
    .O(n965bar),
    .I0(n570bar),
    .I1(n569bar)
  );
  //OR U405
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U405 (
    .O(n569),
    .I0(n568),
    .I1(n567)
  );
  //AND U405bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U405bar (
    .O(n569bar),
    .I0(n568bar),
    .I1(n567bar)
  );
  //OR U406
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U406 (
    .O(n567),
    .I0(n566),
    .I1(n565)
  );
  //AND U406bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U406bar (
    .O(n567bar),
    .I0(n566bar),
    .I1(n565bar)
  );
  //OR U407
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U407 (
    .O(n565),
    .I0(n817),
    .I1(n750)
  );
  //AND U407bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U407bar (
    .O(n565bar),
    .I0(n817bar),
    .I1(n750bar)
  );
  //OR U408
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U408 (
    .O(n750),
    .I0(n564),
    .I1(n563)
  );
  //AND U408bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U408bar (
    .O(n750bar),
    .I0(n564bar),
    .I1(n563bar)
  );
  //OR U409
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U409 (
    .O(n563),
    .I0(n562),
    .I1(n561)
  );
  //AND U409bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U409bar (
    .O(n563bar),
    .I0(n562bar),
    .I1(n561bar)
  );
  //OR U410
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U410 (
    .O(n561),
    .I0(n560),
    .I1(n559)
  );
  //AND U410bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U410bar (
    .O(n561bar),
    .I0(n560bar),
    .I1(n559bar)
  );
  //OR U411
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U411 (
    .O(n559),
    .I0(in[119]),
    .I1(in[103])
  );
  //AND U411bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U411bar (
    .O(n559bar),
    .I0(inbar[119]),
    .I1(inbar[103])
  );
  //OR U412
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U412 (
    .O(n560),
    .I0(in[137]),
    .I1(in[133])
  );
  //AND U412bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U412bar (
    .O(n560bar),
    .I0(inbar[137]),
    .I1(inbar[133])
  );
  //OR U413
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U413 (
    .O(n562),
    .I0(n558),
    .I1(n557)
  );
  //AND U413bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U413bar (
    .O(n562bar),
    .I0(n558bar),
    .I1(n557bar)
  );
  //OR U414
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U414 (
    .O(n557),
    .I0(in[176]),
    .I1(in[173])
  );
  //AND U414bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U414bar (
    .O(n557bar),
    .I0(inbar[176]),
    .I1(inbar[173])
  );
  //OR U415
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U415 (
    .O(n558),
    .I0(in[210]),
    .I1(in[181])
  );
  //AND U415bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U415bar (
    .O(n558bar),
    .I0(inbar[210]),
    .I1(inbar[181])
  );
  //OR U416
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U416 (
    .O(n564),
    .I0(n556),
    .I1(n555)
  );
  //AND U416bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U416bar (
    .O(n564bar),
    .I0(n556bar),
    .I1(n555bar)
  );
  //OR U417
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U417 (
    .O(n555),
    .I0(n554),
    .I1(n553)
  );
  //AND U417bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U417bar (
    .O(n555bar),
    .I0(n554bar),
    .I1(n553bar)
  );
  //OR U418
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U418 (
    .O(n553),
    .I0(in_13),
    .I1(in[234])
  );
  //AND U418bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U418bar (
    .O(n553bar),
    .I0(in_13bar),
    .I1(inbar[234])
  );
  //OR U419
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U419 (
    .O(n554),
    .I0(in_38),
    .I1(in_32)
  );
  //AND U419bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U419bar (
    .O(n554bar),
    .I0(in_38bar),
    .I1(in_32bar)
  );
  //OR U420
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U420 (
    .O(n556),
    .I0(n552),
    .I1(n551)
  );
  //AND U420bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U420bar (
    .O(n556bar),
    .I0(n552bar),
    .I1(n551bar)
  );
  //OR U421
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U421 (
    .O(n551),
    .I0(in_42),
    .I1(in_41)
  );
  //AND U421bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U421bar (
    .O(n551bar),
    .I0(in_42bar),
    .I1(in_41bar)
  );
  //OR U422
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U422 (
    .O(n552),
    .I0(in_7),
    .I1(in_49)
  );
  //AND U422bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U422bar (
    .O(n552bar),
    .I0(in_7bar),
    .I1(in_49bar)
  );
  //OR U423
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U423 (
    .O(n817),
    .I0(n550),
    .I1(n549)
  );
  //AND U423bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U423bar (
    .O(n817bar),
    .I0(n550bar),
    .I1(n549bar)
  );
  //OR U424
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U424 (
    .O(n549),
    .I0(n548),
    .I1(n547)
  );
  //AND U424bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U424bar (
    .O(n549bar),
    .I0(n548bar),
    .I1(n547bar)
  );
  //OR U425
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U425 (
    .O(n547),
    .I0(n546),
    .I1(n545)
  );
  //AND U425bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U425bar (
    .O(n547bar),
    .I0(n546bar),
    .I1(n545bar)
  );
  //OR U426
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U426 (
    .O(n545),
    .I0(in[159]),
    .I1(in[105])
  );
  //AND U426bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U426bar (
    .O(n545bar),
    .I0(inbar[159]),
    .I1(inbar[105])
  );
  //OR U427
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U427 (
    .O(n546),
    .I0(in[206]),
    .I1(in[183])
  );
  //AND U427bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U427bar (
    .O(n546bar),
    .I0(inbar[206]),
    .I1(inbar[183])
  );
  //OR U428
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U428 (
    .O(n548),
    .I0(n544),
    .I1(n543)
  );
  //AND U428bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U428bar (
    .O(n548bar),
    .I0(n544bar),
    .I1(n543bar)
  );
  //OR U429
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U429 (
    .O(n543),
    .I0(in[229]),
    .I1(in[219])
  );
  //AND U429bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U429bar (
    .O(n543bar),
    .I0(inbar[229]),
    .I1(inbar[219])
  );
  //OR U430
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U430 (
    .O(n544),
    .I0(in[235]),
    .I1(in[232])
  );
  //AND U430bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U430bar (
    .O(n544bar),
    .I0(inbar[235]),
    .I1(inbar[232])
  );
  //OR U431
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U431 (
    .O(n550),
    .I0(n542),
    .I1(n541)
  );
  //AND U431bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U431bar (
    .O(n550bar),
    .I0(n542bar),
    .I1(n541bar)
  );
  //OR U432
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U432 (
    .O(n541),
    .I0(n540),
    .I1(n539)
  );
  //AND U432bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U432bar (
    .O(n541bar),
    .I0(n540bar),
    .I1(n539bar)
  );
  //OR U433
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U433 (
    .O(n539),
    .I0(in[249]),
    .I1(in[242])
  );
  //AND U433bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U433bar (
    .O(n539bar),
    .I0(inbar[249]),
    .I1(inbar[242])
  );
  //OR U434
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U434 (
    .O(n540),
    .I0(in[89]),
    .I1(in[254])
  );
  //AND U434bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U434bar (
    .O(n540bar),
    .I0(inbar[89]),
    .I1(inbar[254])
  );
  //OR U435
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U435 (
    .O(n542),
    .I0(n538),
    .I1(n537)
  );
  //AND U435bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U435bar (
    .O(n542bar),
    .I0(n538bar),
    .I1(n537bar)
  );
  //OR U436
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U436 (
    .O(n537),
    .I0(in_14),
    .I1(in[99])
  );
  //AND U436bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U436bar (
    .O(n537bar),
    .I0(in_14bar),
    .I1(inbar[99])
  );
  //OR U437
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U437 (
    .O(n538),
    .I0(in_60),
    .I1(in_18)
  );
  //AND U437bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U437bar (
    .O(n538bar),
    .I0(in_60bar),
    .I1(in_18bar)
  );
  //OR U438
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U438 (
    .O(n566),
    .I0(in[113]),
    .I1(n763)
  );
  //AND U438bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U438bar (
    .O(n566bar),
    .I0(inbar[113]),
    .I1(n763bar)
  );
  //OR U439
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U439 (
    .O(n763),
    .I0(n536),
    .I1(n535)
  );
  //AND U439bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U439bar (
    .O(n763bar),
    .I0(n536bar),
    .I1(n535bar)
  );
  //OR U440
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U440 (
    .O(n535),
    .I0(n534),
    .I1(n533)
  );
  //AND U440bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U440bar (
    .O(n535bar),
    .I0(n534bar),
    .I1(n533bar)
  );
  //OR U441
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U441 (
    .O(n533),
    .I0(n532),
    .I1(n531)
  );
  //AND U441bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U441bar (
    .O(n533bar),
    .I0(n532bar),
    .I1(n531bar)
  );
  //OR U442
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U442 (
    .O(n531),
    .I0(in[115]),
    .I1(in[110])
  );
  //AND U442bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U442bar (
    .O(n531bar),
    .I0(inbar[115]),
    .I1(inbar[110])
  );
  //OR U443
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U443 (
    .O(n532),
    .I0(in[125]),
    .I1(in[117])
  );
  //AND U443bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U443bar (
    .O(n532bar),
    .I0(inbar[125]),
    .I1(inbar[117])
  );
  //OR U444
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U444 (
    .O(n534),
    .I0(n530),
    .I1(n529)
  );
  //AND U444bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U444bar (
    .O(n534bar),
    .I0(n530bar),
    .I1(n529bar)
  );
  //OR U445
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U445 (
    .O(n529),
    .I0(in[180]),
    .I1(in[128])
  );
  //AND U445bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U445bar (
    .O(n529bar),
    .I0(inbar[180]),
    .I1(inbar[128])
  );
  //OR U446
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U446 (
    .O(n530),
    .I0(in[205]),
    .I1(in[201])
  );
  //AND U446bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U446bar (
    .O(n530bar),
    .I0(inbar[205]),
    .I1(inbar[201])
  );
  //OR U447
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U447 (
    .O(n536),
    .I0(n528),
    .I1(n527)
  );
  //AND U447bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U447bar (
    .O(n536bar),
    .I0(n528bar),
    .I1(n527bar)
  );
  //OR U448
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U448 (
    .O(n527),
    .I0(n526),
    .I1(n525)
  );
  //AND U448bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U448bar (
    .O(n527bar),
    .I0(n526bar),
    .I1(n525bar)
  );
  //OR U449
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U449 (
    .O(n525),
    .I0(in[244]),
    .I1(in[239])
  );
  //AND U449bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U449bar (
    .O(n525bar),
    .I0(inbar[244]),
    .I1(inbar[239])
  );
  //OR U450
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U450 (
    .O(n526),
    .I0(in[95]),
    .I1(in[83])
  );
  //AND U450bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U450bar (
    .O(n526bar),
    .I0(inbar[95]),
    .I1(inbar[83])
  );
  //OR U451
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U451 (
    .O(n528),
    .I0(n524),
    .I1(n523)
  );
  //AND U451bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U451bar (
    .O(n528bar),
    .I0(n524bar),
    .I1(n523bar)
  );
  //OR U452
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U452 (
    .O(n523),
    .I0(in_24),
    .I1(in[97])
  );
  //AND U452bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U452bar (
    .O(n523bar),
    .I0(in_24bar),
    .I1(inbar[97])
  );
  //OR U453
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U453 (
    .O(n524),
    .I0(in_33),
    .I1(in_27)
  );
  //AND U453bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U453bar (
    .O(n524bar),
    .I0(in_33bar),
    .I1(in_27bar)
  );
  //OR U454
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U454 (
    .O(n568),
    .I0(n522),
    .I1(n521)
  );
  //AND U454bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U454bar (
    .O(n568bar),
    .I0(n522bar),
    .I1(n521bar)
  );
  //OR U455
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U455 (
    .O(n521),
    .I0(in[145]),
    .I1(in[126])
  );
  //AND U455bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U455bar (
    .O(n521bar),
    .I0(inbar[145]),
    .I1(inbar[126])
  );
  //OR U456
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U456 (
    .O(n522),
    .I0(in[169]),
    .I1(n520)
  );
  //AND U456bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U456bar (
    .O(n522bar),
    .I0(inbar[169]),
    .I1(n520bar)
  );
  //OR U457
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U457 (
    .O(n520),
    .I0(in[221]),
    .I1(in[172])
  );
  //AND U457bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U457bar (
    .O(n520bar),
    .I0(inbar[221]),
    .I1(inbar[172])
  );
  //OR U458
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U458 (
    .O(n570),
    .I0(n519),
    .I1(n518)
  );
  //AND U458bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U458bar (
    .O(n570bar),
    .I0(n519bar),
    .I1(n518bar)
  );
  //OR U459
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U459 (
    .O(n518),
    .I0(n517),
    .I1(n516)
  );
  //AND U459bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U459bar (
    .O(n518bar),
    .I0(n517bar),
    .I1(n516bar)
  );
  //OR U460
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U460 (
    .O(n516),
    .I0(in[241]),
    .I1(in[224])
  );
  //AND U460bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U460bar (
    .O(n516bar),
    .I0(inbar[241]),
    .I1(inbar[224])
  );
  //OR U461
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U461 (
    .O(n517),
    .I0(in[86]),
    .I1(n515)
  );
  //AND U461bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U461bar (
    .O(n517bar),
    .I0(inbar[86]),
    .I1(n515bar)
  );
  //OR U462
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U462 (
    .O(n515),
    .I0(in_43),
    .I1(in_34)
  );
  //AND U462bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U462bar (
    .O(n515bar),
    .I0(in_43bar),
    .I1(in_34bar)
  );
  //OR U463
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U463 (
    .O(n519),
    .I0(n514),
    .I1(n513)
  );
  //AND U463bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U463bar (
    .O(n519bar),
    .I0(n514bar),
    .I1(n513bar)
  );
  //OR U464
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U464 (
    .O(n513),
    .I0(in_65),
    .I1(in_51)
  );
  //AND U464bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U464bar (
    .O(n513bar),
    .I0(in_65bar),
    .I1(in_51bar)
  );
  //OR U465
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U465 (
    .O(n514),
    .I0(in_75),
    .I1(n512)
  );
  //AND U465bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U465bar (
    .O(n514bar),
    .I0(in_75bar),
    .I1(n512bar)
  );
  //OR U466
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U466 (
    .O(n512),
    .I0(in_81),
    .I1(in_77)
  );
  //AND U466bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U466bar (
    .O(n512bar),
    .I0(in_81bar),
    .I1(in_77bar)
  );
  //OR U467
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U467 (
    .O(n778),
    .I0(n511),
    .I1(n510)
  );
  //AND U467bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U467bar (
    .O(n778bar),
    .I0(n511bar),
    .I1(n510bar)
  );
  //OR U468
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U468 (
    .O(n510),
    .I0(n509),
    .I1(n508)
  );
  //AND U468bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U468bar (
    .O(n510bar),
    .I0(n509bar),
    .I1(n508bar)
  );
  //OR U469
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U469 (
    .O(n508),
    .I0(n507),
    .I1(n506)
  );
  //AND U469bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U469bar (
    .O(n508bar),
    .I0(n507bar),
    .I1(n506bar)
  );
  //OR U470
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U470 (
    .O(n506),
    .I0(in[107]),
    .I1(in[101])
  );
  //AND U470bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U470bar (
    .O(n506bar),
    .I0(inbar[107]),
    .I1(inbar[101])
  );
  //OR U471
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U471 (
    .O(n507),
    .I0(in[139]),
    .I1(in[132])
  );
  //AND U471bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U471bar (
    .O(n507bar),
    .I0(inbar[139]),
    .I1(inbar[132])
  );
  //OR U472
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U472 (
    .O(n509),
    .I0(n505),
    .I1(n504)
  );
  //AND U472bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U472bar (
    .O(n509bar),
    .I0(n505bar),
    .I1(n504bar)
  );
  //OR U473
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U473 (
    .O(n504),
    .I0(in[146]),
    .I1(in[141])
  );
  //AND U473bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U473bar (
    .O(n504bar),
    .I0(inbar[146]),
    .I1(inbar[141])
  );
  //OR U474
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U474 (
    .O(n505),
    .I0(in[203]),
    .I1(in[179])
  );
  //AND U474bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U474bar (
    .O(n505bar),
    .I0(inbar[203]),
    .I1(inbar[179])
  );
  //OR U475
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U475 (
    .O(n511),
    .I0(n503),
    .I1(n502)
  );
  //AND U475bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U475bar (
    .O(n511bar),
    .I0(n503bar),
    .I1(n502bar)
  );
  //OR U476
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U476 (
    .O(n502),
    .I0(n501),
    .I1(n500)
  );
  //AND U476bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U476bar (
    .O(n502bar),
    .I0(n501bar),
    .I1(n500bar)
  );
  //OR U477
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U477 (
    .O(n500),
    .I0(in[243]),
    .I1(in[222])
  );
  //AND U477bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U477bar (
    .O(n500bar),
    .I0(inbar[243]),
    .I1(inbar[222])
  );
  //OR U478
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U478 (
    .O(n501),
    .I0(in[251]),
    .I1(in[250])
  );
  //AND U478bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U478bar (
    .O(n501bar),
    .I0(inbar[251]),
    .I1(inbar[250])
  );
  //OR U479
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U479 (
    .O(n503),
    .I0(n499),
    .I1(n498)
  );
  //AND U479bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U479bar (
    .O(n503bar),
    .I0(n499bar),
    .I1(n498bar)
  );
  //OR U480
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U480 (
    .O(n498),
    .I0(in_37),
    .I1(in_19)
  );
  //AND U480bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U480bar (
    .O(n498bar),
    .I0(in_37bar),
    .I1(in_19bar)
  );
  //OR U481
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U481 (
    .O(n499),
    .I0(in_78),
    .I1(in_6)
  );
  //AND U481bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U481bar (
    .O(n499bar),
    .I0(in_78bar),
    .I1(in_6bar)
  );
  //OR U482
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U482 (
    .O(n603),
    .I0(n497),
    .I1(n496)
  );
  //AND U482bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U482bar (
    .O(n603bar),
    .I0(n497bar),
    .I1(n496bar)
  );
  //OR U483
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U483 (
    .O(n496),
    .I0(in[112]),
    .I1(in[102])
  );
  //AND U483bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U483bar (
    .O(n496bar),
    .I0(inbar[112]),
    .I1(inbar[102])
  );
  //OR U484
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U484 (
    .O(n497),
    .I0(in[123]),
    .I1(n495)
  );
  //AND U484bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U484bar (
    .O(n497bar),
    .I0(inbar[123]),
    .I1(n495bar)
  );
  //OR U485
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U485 (
    .O(n495),
    .I0(in[143]),
    .I1(in[130])
  );
  //AND U485bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U485bar (
    .O(n495bar),
    .I0(inbar[143]),
    .I1(inbar[130])
  );
  //OR U486
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U486 (
    .O(n605),
    .I0(n494),
    .I1(n493)
  );
  //AND U486bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U486bar (
    .O(n605bar),
    .I0(n494bar),
    .I1(n493bar)
  );
  //OR U487
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U487 (
    .O(n493),
    .I0(n492),
    .I1(n491)
  );
  //AND U487bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U487bar (
    .O(n493bar),
    .I0(n492bar),
    .I1(n491bar)
  );
  //OR U488
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U488 (
    .O(n491),
    .I0(in[216]),
    .I1(in[213])
  );
  //AND U488bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U488bar (
    .O(n491bar),
    .I0(inbar[216]),
    .I1(inbar[213])
  );
  //OR U489
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U489 (
    .O(n492),
    .I0(in[227]),
    .I1(n490)
  );
  //AND U489bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U489bar (
    .O(n492bar),
    .I0(inbar[227]),
    .I1(n490bar)
  );
  //OR U490
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U490 (
    .O(n490),
    .I0(in_0),
    .I1(in[248])
  );
  //AND U490bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U490bar (
    .O(n490bar),
    .I0(in_0bar),
    .I1(inbar[248])
  );
  //OR U491
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U491 (
    .O(n494),
    .I0(n489),
    .I1(n488)
  );
  //AND U491bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U491bar (
    .O(n494bar),
    .I0(n489bar),
    .I1(n488bar)
  );
  //OR U492
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U492 (
    .O(n488),
    .I0(in_46),
    .I1(in_44)
  );
  //AND U492bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U492bar (
    .O(n488bar),
    .I0(in_46bar),
    .I1(in_44bar)
  );
  //OR U493
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U493 (
    .O(n489),
    .I0(in_50),
    .I1(n487)
  );
  //AND U493bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U493bar (
    .O(n489bar),
    .I0(in_50bar),
    .I1(n487bar)
  );
  //OR U494
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U494 (
    .O(n487),
    .I0(in_9),
    .I1(in_80)
  );
  //AND U494bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U494bar (
    .O(n487bar),
    .I0(in_9bar),
    .I1(in_80bar)
  );
endmodule

module sBox_4 ( in, out );

  input wire [7:0] in;
//input_done

  output wire [7:0] out;
//output_done

  wire [255:0] decodeOut;
//wire_done

  decode_4 dec ( .in(in), .out(decodeOut) );
  encode_4 enc ( .in(decodeOut), .out(out) );
endmodule

module CD2_17 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD2_18 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD2_19 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD2_20 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD4_9 ( a, b, y );

  input wire [3:0] a;
  input wire [3:0] b;
  wire [3:0] abar;
  wire [3:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
//input_done

  output wire [15:0] y;
  wire [15:0] ybar;
//output_done

//wire_done

  //AND U1
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1 (
    .O(y[9]),
    .I0(b[1]),
    .I1(a[2])
  );
  //OR U1bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1bar (
    .O(ybar[9]),
    .I0(bbar[1]),
    .I1(abar[2])
  );
  //AND U2
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2 (
    .O(y[8]),
    .I0(b[0]),
    .I1(a[2])
  );
  //OR U2bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2bar (
    .O(ybar[8]),
    .I0(bbar[0]),
    .I1(abar[2])
  );
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[7]),
    .I0(b[3]),
    .I1(a[1])
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[7]),
    .I0(bbar[3]),
    .I1(abar[1])
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[6]),
    .I0(b[2]),
    .I1(a[1])
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[6]),
    .I0(bbar[2]),
    .I1(abar[1])
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[5]),
    .I0(a[1]),
    .I1(b[1])
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[5]),
    .I0(abar[1]),
    .I1(bbar[1])
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[4]),
    .I0(a[1]),
    .I1(b[0])
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[4]),
    .I0(abar[1]),
    .I1(bbar[0])
  );
  //AND U7
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7 (
    .O(y[3]),
    .I0(a[0]),
    .I1(b[3])
  );
  //OR U7bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7bar (
    .O(ybar[3]),
    .I0(abar[0]),
    .I1(bbar[3])
  );
  //AND U8
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8 (
    .O(y[2]),
    .I0(a[0]),
    .I1(b[2])
  );
  //OR U8bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8bar (
    .O(ybar[2]),
    .I0(abar[0]),
    .I1(bbar[2])
  );
  //AND U9
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9 (
    .O(y[1]),
    .I0(a[0]),
    .I1(b[1])
  );
  //OR U9bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9bar (
    .O(ybar[1]),
    .I0(abar[0]),
    .I1(bbar[1])
  );
  //AND U10
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10 (
    .O(y[15]),
    .I0(a[3]),
    .I1(b[3])
  );
  //OR U10bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10bar (
    .O(ybar[15]),
    .I0(abar[3]),
    .I1(bbar[3])
  );
  //AND U11
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11 (
    .O(y[14]),
    .I0(a[3]),
    .I1(b[2])
  );
  //OR U11bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11bar (
    .O(ybar[14]),
    .I0(abar[3]),
    .I1(bbar[2])
  );
  //AND U12
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12 (
    .O(y[13]),
    .I0(a[3]),
    .I1(b[1])
  );
  //OR U12bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12bar (
    .O(ybar[13]),
    .I0(abar[3]),
    .I1(bbar[1])
  );
  //AND U13
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13 (
    .O(y[12]),
    .I0(a[3]),
    .I1(b[0])
  );
  //OR U13bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13bar (
    .O(ybar[12]),
    .I0(abar[3]),
    .I1(bbar[0])
  );
  //AND U14
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14 (
    .O(y[11]),
    .I0(b[3]),
    .I1(a[2])
  );
  //OR U14bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14bar (
    .O(ybar[11]),
    .I0(bbar[3]),
    .I1(abar[2])
  );
  //AND U15
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15 (
    .O(y[10]),
    .I0(b[2]),
    .I1(a[2])
  );
  //OR U15bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15bar (
    .O(ybar[10]),
    .I0(bbar[2]),
    .I1(abar[2])
  );
  //AND U16
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16 (
    .O(y[0]),
    .I0(a[0]),
    .I1(b[0])
  );
  //OR U16bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16bar (
    .O(ybar[0]),
    .I0(abar[0]),
    .I1(bbar[0])
  );
endmodule

module CD4_10 ( a, b, y );

  input wire [3:0] a;
  input wire [3:0] b;
  wire [3:0] abar;
  wire [3:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
//input_done

  output wire [15:0] y;
  wire [15:0] ybar;
//output_done

//wire_done

  //AND U1
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1 (
    .O(y[9]),
    .I0(b[1]),
    .I1(a[2])
  );
  //OR U1bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1bar (
    .O(ybar[9]),
    .I0(bbar[1]),
    .I1(abar[2])
  );
  //AND U2
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2 (
    .O(y[8]),
    .I0(b[0]),
    .I1(a[2])
  );
  //OR U2bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2bar (
    .O(ybar[8]),
    .I0(bbar[0]),
    .I1(abar[2])
  );
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[7]),
    .I0(b[3]),
    .I1(a[1])
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[7]),
    .I0(bbar[3]),
    .I1(abar[1])
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[6]),
    .I0(b[2]),
    .I1(a[1])
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[6]),
    .I0(bbar[2]),
    .I1(abar[1])
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[5]),
    .I0(a[1]),
    .I1(b[1])
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[5]),
    .I0(abar[1]),
    .I1(bbar[1])
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[4]),
    .I0(a[1]),
    .I1(b[0])
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[4]),
    .I0(abar[1]),
    .I1(bbar[0])
  );
  //AND U7
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7 (
    .O(y[3]),
    .I0(a[0]),
    .I1(b[3])
  );
  //OR U7bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7bar (
    .O(ybar[3]),
    .I0(abar[0]),
    .I1(bbar[3])
  );
  //AND U8
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8 (
    .O(y[2]),
    .I0(a[0]),
    .I1(b[2])
  );
  //OR U8bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8bar (
    .O(ybar[2]),
    .I0(abar[0]),
    .I1(bbar[2])
  );
  //AND U9
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9 (
    .O(y[1]),
    .I0(a[0]),
    .I1(b[1])
  );
  //OR U9bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9bar (
    .O(ybar[1]),
    .I0(abar[0]),
    .I1(bbar[1])
  );
  //AND U10
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10 (
    .O(y[15]),
    .I0(a[3]),
    .I1(b[3])
  );
  //OR U10bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10bar (
    .O(ybar[15]),
    .I0(abar[3]),
    .I1(bbar[3])
  );
  //AND U11
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11 (
    .O(y[14]),
    .I0(a[3]),
    .I1(b[2])
  );
  //OR U11bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11bar (
    .O(ybar[14]),
    .I0(abar[3]),
    .I1(bbar[2])
  );
  //AND U12
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12 (
    .O(y[13]),
    .I0(a[3]),
    .I1(b[1])
  );
  //OR U12bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12bar (
    .O(ybar[13]),
    .I0(abar[3]),
    .I1(bbar[1])
  );
  //AND U13
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13 (
    .O(y[12]),
    .I0(a[3]),
    .I1(b[0])
  );
  //OR U13bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13bar (
    .O(ybar[12]),
    .I0(abar[3]),
    .I1(bbar[0])
  );
  //AND U14
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14 (
    .O(y[11]),
    .I0(b[3]),
    .I1(a[2])
  );
  //OR U14bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14bar (
    .O(ybar[11]),
    .I0(bbar[3]),
    .I1(abar[2])
  );
  //AND U15
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15 (
    .O(y[10]),
    .I0(b[2]),
    .I1(a[2])
  );
  //OR U15bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15bar (
    .O(ybar[10]),
    .I0(bbar[2]),
    .I1(abar[2])
  );
  //AND U16
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16 (
    .O(y[0]),
    .I0(a[0]),
    .I1(b[0])
  );
  //OR U16bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16bar (
    .O(ybar[0]),
    .I0(abar[0]),
    .I1(bbar[0])
  );
endmodule

module CD16_5 ( a, b, y );

  input wire [15:0] a;
  input wire [15:0] b;
  wire [15:0] abar;
  wire [15:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign abar[8] = ~a[8];
  assign abar[9] = ~a[9];
  assign abar[10] = ~a[10];
  assign abar[11] = ~a[11];
  assign abar[12] = ~a[12];
  assign abar[13] = ~a[13];
  assign abar[14] = ~a[14];
  assign abar[15] = ~a[15];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign bbar[8] = ~b[8];
  assign bbar[9] = ~b[9];
  assign bbar[10] = ~b[10];
  assign bbar[11] = ~b[11];
  assign bbar[12] = ~b[12];
  assign bbar[13] = ~b[13];
  assign bbar[14] = ~b[14];
  assign bbar[15] = ~b[15];
//input_done

  output wire [255:0] y;
  wire [255:0] ybar;
//output_done

//wire_done

  //AND U1
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1 (
    .O(y[9]),
    .I0(b[9]),
    .I1(a[0])
  );
  //OR U1bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1bar (
    .O(ybar[9]),
    .I0(bbar[9]),
    .I1(abar[0])
  );
  //AND U2
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2 (
    .O(y[99]),
    .I0(b[3]),
    .I1(a[6])
  );
  //OR U2bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2bar (
    .O(ybar[99]),
    .I0(bbar[3]),
    .I1(abar[6])
  );
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[98]),
    .I0(b[2]),
    .I1(a[6])
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[98]),
    .I0(bbar[2]),
    .I1(abar[6])
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[97]),
    .I0(b[1]),
    .I1(a[6])
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[97]),
    .I0(bbar[1]),
    .I1(abar[6])
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[96]),
    .I0(b[0]),
    .I1(a[6])
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[96]),
    .I0(bbar[0]),
    .I1(abar[6])
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[95]),
    .I0(b[15]),
    .I1(a[5])
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[95]),
    .I0(bbar[15]),
    .I1(abar[5])
  );
  //AND U7
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7 (
    .O(y[94]),
    .I0(b[14]),
    .I1(a[5])
  );
  //OR U7bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7bar (
    .O(ybar[94]),
    .I0(bbar[14]),
    .I1(abar[5])
  );
  //AND U8
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8 (
    .O(y[93]),
    .I0(b[13]),
    .I1(a[5])
  );
  //OR U8bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8bar (
    .O(ybar[93]),
    .I0(bbar[13]),
    .I1(abar[5])
  );
  //AND U9
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9 (
    .O(y[92]),
    .I0(b[12]),
    .I1(a[5])
  );
  //OR U9bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9bar (
    .O(ybar[92]),
    .I0(bbar[12]),
    .I1(abar[5])
  );
  //AND U10
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10 (
    .O(y[91]),
    .I0(b[11]),
    .I1(a[5])
  );
  //OR U10bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10bar (
    .O(ybar[91]),
    .I0(bbar[11]),
    .I1(abar[5])
  );
  //AND U11
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11 (
    .O(y[90]),
    .I0(b[10]),
    .I1(a[5])
  );
  //OR U11bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11bar (
    .O(ybar[90]),
    .I0(bbar[10]),
    .I1(abar[5])
  );
  //AND U12
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12 (
    .O(y[8]),
    .I0(b[8]),
    .I1(a[0])
  );
  //OR U12bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12bar (
    .O(ybar[8]),
    .I0(bbar[8]),
    .I1(abar[0])
  );
  //AND U13
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13 (
    .O(y[89]),
    .I0(a[5]),
    .I1(b[9])
  );
  //OR U13bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13bar (
    .O(ybar[89]),
    .I0(abar[5]),
    .I1(bbar[9])
  );
  //AND U14
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14 (
    .O(y[88]),
    .I0(b[8]),
    .I1(a[5])
  );
  //OR U14bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14bar (
    .O(ybar[88]),
    .I0(bbar[8]),
    .I1(abar[5])
  );
  //AND U15
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15 (
    .O(y[87]),
    .I0(b[7]),
    .I1(a[5])
  );
  //OR U15bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15bar (
    .O(ybar[87]),
    .I0(bbar[7]),
    .I1(abar[5])
  );
  //AND U16
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16 (
    .O(y[86]),
    .I0(b[6]),
    .I1(a[5])
  );
  //OR U16bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16bar (
    .O(ybar[86]),
    .I0(bbar[6]),
    .I1(abar[5])
  );
  //AND U17
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U17 (
    .O(y[85]),
    .I0(b[5]),
    .I1(a[5])
  );
  //OR U17bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U17bar (
    .O(ybar[85]),
    .I0(bbar[5]),
    .I1(abar[5])
  );
  //AND U18
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U18 (
    .O(y[84]),
    .I0(b[4]),
    .I1(a[5])
  );
  //OR U18bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U18bar (
    .O(ybar[84]),
    .I0(bbar[4]),
    .I1(abar[5])
  );
  //AND U19
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U19 (
    .O(y[83]),
    .I0(a[5]),
    .I1(b[3])
  );
  //OR U19bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U19bar (
    .O(ybar[83]),
    .I0(abar[5]),
    .I1(bbar[3])
  );
  //AND U20
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U20 (
    .O(y[82]),
    .I0(a[5]),
    .I1(b[2])
  );
  //OR U20bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U20bar (
    .O(ybar[82]),
    .I0(abar[5]),
    .I1(bbar[2])
  );
  //AND U21
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U21 (
    .O(y[81]),
    .I0(a[5]),
    .I1(b[1])
  );
  //OR U21bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U21bar (
    .O(ybar[81]),
    .I0(abar[5]),
    .I1(bbar[1])
  );
  //AND U22
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U22 (
    .O(y[80]),
    .I0(a[5]),
    .I1(b[0])
  );
  //OR U22bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U22bar (
    .O(ybar[80]),
    .I0(abar[5]),
    .I1(bbar[0])
  );
  //AND U23
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U23 (
    .O(y[7]),
    .I0(b[7]),
    .I1(a[0])
  );
  //OR U23bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U23bar (
    .O(ybar[7]),
    .I0(bbar[7]),
    .I1(abar[0])
  );
  //AND U24
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U24 (
    .O(y[79]),
    .I0(a[4]),
    .I1(b[15])
  );
  //OR U24bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U24bar (
    .O(ybar[79]),
    .I0(abar[4]),
    .I1(bbar[15])
  );
  //AND U25
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U25 (
    .O(y[78]),
    .I0(a[4]),
    .I1(b[14])
  );
  //OR U25bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U25bar (
    .O(ybar[78]),
    .I0(abar[4]),
    .I1(bbar[14])
  );
  //AND U26
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U26 (
    .O(y[77]),
    .I0(a[4]),
    .I1(b[13])
  );
  //OR U26bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U26bar (
    .O(ybar[77]),
    .I0(abar[4]),
    .I1(bbar[13])
  );
  //AND U27
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U27 (
    .O(y[76]),
    .I0(a[4]),
    .I1(b[12])
  );
  //OR U27bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U27bar (
    .O(ybar[76]),
    .I0(abar[4]),
    .I1(bbar[12])
  );
  //AND U28
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U28 (
    .O(y[75]),
    .I0(a[4]),
    .I1(b[11])
  );
  //OR U28bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U28bar (
    .O(ybar[75]),
    .I0(abar[4]),
    .I1(bbar[11])
  );
  //AND U29
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U29 (
    .O(y[74]),
    .I0(a[4]),
    .I1(b[10])
  );
  //OR U29bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U29bar (
    .O(ybar[74]),
    .I0(abar[4]),
    .I1(bbar[10])
  );
  //AND U30
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U30 (
    .O(y[73]),
    .I0(a[4]),
    .I1(b[9])
  );
  //OR U30bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U30bar (
    .O(ybar[73]),
    .I0(abar[4]),
    .I1(bbar[9])
  );
  //AND U31
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U31 (
    .O(y[72]),
    .I0(a[4]),
    .I1(b[8])
  );
  //OR U31bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U31bar (
    .O(ybar[72]),
    .I0(abar[4]),
    .I1(bbar[8])
  );
  //AND U32
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U32 (
    .O(y[71]),
    .I0(a[4]),
    .I1(b[7])
  );
  //OR U32bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U32bar (
    .O(ybar[71]),
    .I0(abar[4]),
    .I1(bbar[7])
  );
  //AND U33
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U33 (
    .O(y[70]),
    .I0(a[4]),
    .I1(b[6])
  );
  //OR U33bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U33bar (
    .O(ybar[70]),
    .I0(abar[4]),
    .I1(bbar[6])
  );
  //AND U34
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U34 (
    .O(y[6]),
    .I0(b[6]),
    .I1(a[0])
  );
  //OR U34bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U34bar (
    .O(ybar[6]),
    .I0(bbar[6]),
    .I1(abar[0])
  );
  //AND U35
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U35 (
    .O(y[69]),
    .I0(a[4]),
    .I1(b[5])
  );
  //OR U35bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U35bar (
    .O(ybar[69]),
    .I0(abar[4]),
    .I1(bbar[5])
  );
  //AND U36
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U36 (
    .O(y[68]),
    .I0(a[4]),
    .I1(b[4])
  );
  //OR U36bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U36bar (
    .O(ybar[68]),
    .I0(abar[4]),
    .I1(bbar[4])
  );
  //AND U37
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U37 (
    .O(y[67]),
    .I0(a[4]),
    .I1(b[3])
  );
  //OR U37bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U37bar (
    .O(ybar[67]),
    .I0(abar[4]),
    .I1(bbar[3])
  );
  //AND U38
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U38 (
    .O(y[66]),
    .I0(a[4]),
    .I1(b[2])
  );
  //OR U38bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U38bar (
    .O(ybar[66]),
    .I0(abar[4]),
    .I1(bbar[2])
  );
  //AND U39
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U39 (
    .O(y[65]),
    .I0(a[4]),
    .I1(b[1])
  );
  //OR U39bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U39bar (
    .O(ybar[65]),
    .I0(abar[4]),
    .I1(bbar[1])
  );
  //AND U40
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U40 (
    .O(y[64]),
    .I0(a[4]),
    .I1(b[0])
  );
  //OR U40bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U40bar (
    .O(ybar[64]),
    .I0(abar[4]),
    .I1(bbar[0])
  );
  //AND U41
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U41 (
    .O(y[63]),
    .I0(a[3]),
    .I1(b[15])
  );
  //OR U41bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U41bar (
    .O(ybar[63]),
    .I0(abar[3]),
    .I1(bbar[15])
  );
  //AND U42
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U42 (
    .O(y[62]),
    .I0(a[3]),
    .I1(b[14])
  );
  //OR U42bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U42bar (
    .O(ybar[62]),
    .I0(abar[3]),
    .I1(bbar[14])
  );
  //AND U43
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U43 (
    .O(y[61]),
    .I0(a[3]),
    .I1(b[13])
  );
  //OR U43bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U43bar (
    .O(ybar[61]),
    .I0(abar[3]),
    .I1(bbar[13])
  );
  //AND U44
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U44 (
    .O(y[60]),
    .I0(a[3]),
    .I1(b[12])
  );
  //OR U44bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U44bar (
    .O(ybar[60]),
    .I0(abar[3]),
    .I1(bbar[12])
  );
  //AND U45
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U45 (
    .O(y[5]),
    .I0(b[5]),
    .I1(a[0])
  );
  //OR U45bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U45bar (
    .O(ybar[5]),
    .I0(bbar[5]),
    .I1(abar[0])
  );
  //AND U46
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U46 (
    .O(y[59]),
    .I0(a[3]),
    .I1(b[11])
  );
  //OR U46bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U46bar (
    .O(ybar[59]),
    .I0(abar[3]),
    .I1(bbar[11])
  );
  //AND U47
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U47 (
    .O(y[58]),
    .I0(a[3]),
    .I1(b[10])
  );
  //OR U47bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U47bar (
    .O(ybar[58]),
    .I0(abar[3]),
    .I1(bbar[10])
  );
  //AND U48
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U48 (
    .O(y[57]),
    .I0(a[3]),
    .I1(b[9])
  );
  //OR U48bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U48bar (
    .O(ybar[57]),
    .I0(abar[3]),
    .I1(bbar[9])
  );
  //AND U49
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U49 (
    .O(y[56]),
    .I0(a[3]),
    .I1(b[8])
  );
  //OR U49bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U49bar (
    .O(ybar[56]),
    .I0(abar[3]),
    .I1(bbar[8])
  );
  //AND U50
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U50 (
    .O(y[55]),
    .I0(a[3]),
    .I1(b[7])
  );
  //OR U50bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U50bar (
    .O(ybar[55]),
    .I0(abar[3]),
    .I1(bbar[7])
  );
  //AND U51
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U51 (
    .O(y[54]),
    .I0(a[3]),
    .I1(b[6])
  );
  //OR U51bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U51bar (
    .O(ybar[54]),
    .I0(abar[3]),
    .I1(bbar[6])
  );
  //AND U52
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U52 (
    .O(y[53]),
    .I0(a[3]),
    .I1(b[5])
  );
  //OR U52bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U52bar (
    .O(ybar[53]),
    .I0(abar[3]),
    .I1(bbar[5])
  );
  //AND U53
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U53 (
    .O(y[52]),
    .I0(a[3]),
    .I1(b[4])
  );
  //OR U53bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U53bar (
    .O(ybar[52]),
    .I0(abar[3]),
    .I1(bbar[4])
  );
  //AND U54
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U54 (
    .O(y[51]),
    .I0(a[3]),
    .I1(b[3])
  );
  //OR U54bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U54bar (
    .O(ybar[51]),
    .I0(abar[3]),
    .I1(bbar[3])
  );
  //AND U55
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U55 (
    .O(y[50]),
    .I0(a[3]),
    .I1(b[2])
  );
  //OR U55bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U55bar (
    .O(ybar[50]),
    .I0(abar[3]),
    .I1(bbar[2])
  );
  //AND U56
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U56 (
    .O(y[4]),
    .I0(b[4]),
    .I1(a[0])
  );
  //OR U56bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U56bar (
    .O(ybar[4]),
    .I0(bbar[4]),
    .I1(abar[0])
  );
  //AND U57
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U57 (
    .O(y[49]),
    .I0(a[3]),
    .I1(b[1])
  );
  //OR U57bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U57bar (
    .O(ybar[49]),
    .I0(abar[3]),
    .I1(bbar[1])
  );
  //AND U58
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U58 (
    .O(y[48]),
    .I0(a[3]),
    .I1(b[0])
  );
  //OR U58bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U58bar (
    .O(ybar[48]),
    .I0(abar[3]),
    .I1(bbar[0])
  );
  //AND U59
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U59 (
    .O(y[47]),
    .I0(a[2]),
    .I1(b[15])
  );
  //OR U59bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U59bar (
    .O(ybar[47]),
    .I0(abar[2]),
    .I1(bbar[15])
  );
  //AND U60
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U60 (
    .O(y[46]),
    .I0(a[2]),
    .I1(b[14])
  );
  //OR U60bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U60bar (
    .O(ybar[46]),
    .I0(abar[2]),
    .I1(bbar[14])
  );
  //AND U61
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U61 (
    .O(y[45]),
    .I0(a[2]),
    .I1(b[13])
  );
  //OR U61bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U61bar (
    .O(ybar[45]),
    .I0(abar[2]),
    .I1(bbar[13])
  );
  //AND U62
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U62 (
    .O(y[44]),
    .I0(a[2]),
    .I1(b[12])
  );
  //OR U62bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U62bar (
    .O(ybar[44]),
    .I0(abar[2]),
    .I1(bbar[12])
  );
  //AND U63
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U63 (
    .O(y[43]),
    .I0(a[2]),
    .I1(b[11])
  );
  //OR U63bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U63bar (
    .O(ybar[43]),
    .I0(abar[2]),
    .I1(bbar[11])
  );
  //AND U64
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U64 (
    .O(y[42]),
    .I0(a[2]),
    .I1(b[10])
  );
  //OR U64bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U64bar (
    .O(ybar[42]),
    .I0(abar[2]),
    .I1(bbar[10])
  );
  //AND U65
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U65 (
    .O(y[41]),
    .I0(a[2]),
    .I1(b[9])
  );
  //OR U65bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U65bar (
    .O(ybar[41]),
    .I0(abar[2]),
    .I1(bbar[9])
  );
  //AND U66
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U66 (
    .O(y[40]),
    .I0(a[2]),
    .I1(b[8])
  );
  //OR U66bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U66bar (
    .O(ybar[40]),
    .I0(abar[2]),
    .I1(bbar[8])
  );
  //AND U67
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U67 (
    .O(y[3]),
    .I0(b[3]),
    .I1(a[0])
  );
  //OR U67bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U67bar (
    .O(ybar[3]),
    .I0(bbar[3]),
    .I1(abar[0])
  );
  //AND U68
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U68 (
    .O(y[39]),
    .I0(a[2]),
    .I1(b[7])
  );
  //OR U68bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U68bar (
    .O(ybar[39]),
    .I0(abar[2]),
    .I1(bbar[7])
  );
  //AND U69
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U69 (
    .O(y[38]),
    .I0(a[2]),
    .I1(b[6])
  );
  //OR U69bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U69bar (
    .O(ybar[38]),
    .I0(abar[2]),
    .I1(bbar[6])
  );
  //AND U70
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U70 (
    .O(y[37]),
    .I0(a[2]),
    .I1(b[5])
  );
  //OR U70bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U70bar (
    .O(ybar[37]),
    .I0(abar[2]),
    .I1(bbar[5])
  );
  //AND U71
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U71 (
    .O(y[36]),
    .I0(a[2]),
    .I1(b[4])
  );
  //OR U71bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U71bar (
    .O(ybar[36]),
    .I0(abar[2]),
    .I1(bbar[4])
  );
  //AND U72
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U72 (
    .O(y[35]),
    .I0(a[2]),
    .I1(b[3])
  );
  //OR U72bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U72bar (
    .O(ybar[35]),
    .I0(abar[2]),
    .I1(bbar[3])
  );
  //AND U73
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U73 (
    .O(y[34]),
    .I0(a[2]),
    .I1(b[2])
  );
  //OR U73bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U73bar (
    .O(ybar[34]),
    .I0(abar[2]),
    .I1(bbar[2])
  );
  //AND U74
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U74 (
    .O(y[33]),
    .I0(a[2]),
    .I1(b[1])
  );
  //OR U74bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U74bar (
    .O(ybar[33]),
    .I0(abar[2]),
    .I1(bbar[1])
  );
  //AND U75
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U75 (
    .O(y[32]),
    .I0(a[2]),
    .I1(b[0])
  );
  //OR U75bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U75bar (
    .O(ybar[32]),
    .I0(abar[2]),
    .I1(bbar[0])
  );
  //AND U76
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U76 (
    .O(y[31]),
    .I0(a[1]),
    .I1(b[15])
  );
  //OR U76bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U76bar (
    .O(ybar[31]),
    .I0(abar[1]),
    .I1(bbar[15])
  );
  //AND U77
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U77 (
    .O(y[30]),
    .I0(a[1]),
    .I1(b[14])
  );
  //OR U77bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U77bar (
    .O(ybar[30]),
    .I0(abar[1]),
    .I1(bbar[14])
  );
  //AND U78
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U78 (
    .O(y[2]),
    .I0(b[2]),
    .I1(a[0])
  );
  //OR U78bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U78bar (
    .O(ybar[2]),
    .I0(bbar[2]),
    .I1(abar[0])
  );
  //AND U79
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U79 (
    .O(y[29]),
    .I0(a[1]),
    .I1(b[13])
  );
  //OR U79bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U79bar (
    .O(ybar[29]),
    .I0(abar[1]),
    .I1(bbar[13])
  );
  //AND U80
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U80 (
    .O(y[28]),
    .I0(a[1]),
    .I1(b[12])
  );
  //OR U80bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U80bar (
    .O(ybar[28]),
    .I0(abar[1]),
    .I1(bbar[12])
  );
  //AND U81
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U81 (
    .O(y[27]),
    .I0(a[1]),
    .I1(b[11])
  );
  //OR U81bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U81bar (
    .O(ybar[27]),
    .I0(abar[1]),
    .I1(bbar[11])
  );
  //AND U82
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U82 (
    .O(y[26]),
    .I0(a[1]),
    .I1(b[10])
  );
  //OR U82bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U82bar (
    .O(ybar[26]),
    .I0(abar[1]),
    .I1(bbar[10])
  );
  //AND U83
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U83 (
    .O(y[25]),
    .I0(a[1]),
    .I1(b[9])
  );
  //OR U83bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U83bar (
    .O(ybar[25]),
    .I0(abar[1]),
    .I1(bbar[9])
  );
  //AND U84
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U84 (
    .O(y[255]),
    .I0(a[15]),
    .I1(b[15])
  );
  //OR U84bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U84bar (
    .O(ybar[255]),
    .I0(abar[15]),
    .I1(bbar[15])
  );
  //AND U85
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U85 (
    .O(y[254]),
    .I0(a[15]),
    .I1(b[14])
  );
  //OR U85bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U85bar (
    .O(ybar[254]),
    .I0(abar[15]),
    .I1(bbar[14])
  );
  //AND U86
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U86 (
    .O(y[253]),
    .I0(a[15]),
    .I1(b[13])
  );
  //OR U86bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U86bar (
    .O(ybar[253]),
    .I0(abar[15]),
    .I1(bbar[13])
  );
  //AND U87
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U87 (
    .O(y[252]),
    .I0(a[15]),
    .I1(b[12])
  );
  //OR U87bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U87bar (
    .O(ybar[252]),
    .I0(abar[15]),
    .I1(bbar[12])
  );
  //AND U88
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U88 (
    .O(y[251]),
    .I0(a[15]),
    .I1(b[11])
  );
  //OR U88bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U88bar (
    .O(ybar[251]),
    .I0(abar[15]),
    .I1(bbar[11])
  );
  //AND U89
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U89 (
    .O(y[250]),
    .I0(a[15]),
    .I1(b[10])
  );
  //OR U89bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U89bar (
    .O(ybar[250]),
    .I0(abar[15]),
    .I1(bbar[10])
  );
  //AND U90
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U90 (
    .O(y[24]),
    .I0(a[1]),
    .I1(b[8])
  );
  //OR U90bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U90bar (
    .O(ybar[24]),
    .I0(abar[1]),
    .I1(bbar[8])
  );
  //AND U91
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U91 (
    .O(y[249]),
    .I0(a[15]),
    .I1(b[9])
  );
  //OR U91bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U91bar (
    .O(ybar[249]),
    .I0(abar[15]),
    .I1(bbar[9])
  );
  //AND U92
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U92 (
    .O(y[248]),
    .I0(a[15]),
    .I1(b[8])
  );
  //OR U92bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U92bar (
    .O(ybar[248]),
    .I0(abar[15]),
    .I1(bbar[8])
  );
  //AND U93
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U93 (
    .O(y[247]),
    .I0(a[15]),
    .I1(b[7])
  );
  //OR U93bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U93bar (
    .O(ybar[247]),
    .I0(abar[15]),
    .I1(bbar[7])
  );
  //AND U94
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U94 (
    .O(y[246]),
    .I0(a[15]),
    .I1(b[6])
  );
  //OR U94bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U94bar (
    .O(ybar[246]),
    .I0(abar[15]),
    .I1(bbar[6])
  );
  //AND U95
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U95 (
    .O(y[245]),
    .I0(a[15]),
    .I1(b[5])
  );
  //OR U95bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U95bar (
    .O(ybar[245]),
    .I0(abar[15]),
    .I1(bbar[5])
  );
  //AND U96
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U96 (
    .O(y[244]),
    .I0(a[15]),
    .I1(b[4])
  );
  //OR U96bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U96bar (
    .O(ybar[244]),
    .I0(abar[15]),
    .I1(bbar[4])
  );
  //AND U97
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U97 (
    .O(y[243]),
    .I0(a[15]),
    .I1(b[3])
  );
  //OR U97bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U97bar (
    .O(ybar[243]),
    .I0(abar[15]),
    .I1(bbar[3])
  );
  //AND U98
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U98 (
    .O(y[242]),
    .I0(a[15]),
    .I1(b[2])
  );
  //OR U98bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U98bar (
    .O(ybar[242]),
    .I0(abar[15]),
    .I1(bbar[2])
  );
  //AND U99
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U99 (
    .O(y[241]),
    .I0(a[15]),
    .I1(b[1])
  );
  //OR U99bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U99bar (
    .O(ybar[241]),
    .I0(abar[15]),
    .I1(bbar[1])
  );
  //AND U100
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U100 (
    .O(y[240]),
    .I0(a[15]),
    .I1(b[0])
  );
  //OR U100bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U100bar (
    .O(ybar[240]),
    .I0(abar[15]),
    .I1(bbar[0])
  );
  //AND U101
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U101 (
    .O(y[23]),
    .I0(a[1]),
    .I1(b[7])
  );
  //OR U101bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U101bar (
    .O(ybar[23]),
    .I0(abar[1]),
    .I1(bbar[7])
  );
  //AND U102
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U102 (
    .O(y[239]),
    .I0(a[14]),
    .I1(b[15])
  );
  //OR U102bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U102bar (
    .O(ybar[239]),
    .I0(abar[14]),
    .I1(bbar[15])
  );
  //AND U103
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U103 (
    .O(y[238]),
    .I0(a[14]),
    .I1(b[14])
  );
  //OR U103bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U103bar (
    .O(ybar[238]),
    .I0(abar[14]),
    .I1(bbar[14])
  );
  //AND U104
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U104 (
    .O(y[237]),
    .I0(a[14]),
    .I1(b[13])
  );
  //OR U104bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U104bar (
    .O(ybar[237]),
    .I0(abar[14]),
    .I1(bbar[13])
  );
  //AND U105
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U105 (
    .O(y[236]),
    .I0(a[14]),
    .I1(b[12])
  );
  //OR U105bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U105bar (
    .O(ybar[236]),
    .I0(abar[14]),
    .I1(bbar[12])
  );
  //AND U106
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U106 (
    .O(y[235]),
    .I0(a[14]),
    .I1(b[11])
  );
  //OR U106bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U106bar (
    .O(ybar[235]),
    .I0(abar[14]),
    .I1(bbar[11])
  );
  //AND U107
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U107 (
    .O(y[234]),
    .I0(a[14]),
    .I1(b[10])
  );
  //OR U107bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U107bar (
    .O(ybar[234]),
    .I0(abar[14]),
    .I1(bbar[10])
  );
  //AND U108
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U108 (
    .O(y[233]),
    .I0(a[14]),
    .I1(b[9])
  );
  //OR U108bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U108bar (
    .O(ybar[233]),
    .I0(abar[14]),
    .I1(bbar[9])
  );
  //AND U109
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U109 (
    .O(y[232]),
    .I0(a[14]),
    .I1(b[8])
  );
  //OR U109bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U109bar (
    .O(ybar[232]),
    .I0(abar[14]),
    .I1(bbar[8])
  );
  //AND U110
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U110 (
    .O(y[231]),
    .I0(a[14]),
    .I1(b[7])
  );
  //OR U110bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U110bar (
    .O(ybar[231]),
    .I0(abar[14]),
    .I1(bbar[7])
  );
  //AND U111
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U111 (
    .O(y[230]),
    .I0(a[14]),
    .I1(b[6])
  );
  //OR U111bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U111bar (
    .O(ybar[230]),
    .I0(abar[14]),
    .I1(bbar[6])
  );
  //AND U112
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U112 (
    .O(y[22]),
    .I0(a[1]),
    .I1(b[6])
  );
  //OR U112bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U112bar (
    .O(ybar[22]),
    .I0(abar[1]),
    .I1(bbar[6])
  );
  //AND U113
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U113 (
    .O(y[229]),
    .I0(a[14]),
    .I1(b[5])
  );
  //OR U113bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U113bar (
    .O(ybar[229]),
    .I0(abar[14]),
    .I1(bbar[5])
  );
  //AND U114
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U114 (
    .O(y[228]),
    .I0(a[14]),
    .I1(b[4])
  );
  //OR U114bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U114bar (
    .O(ybar[228]),
    .I0(abar[14]),
    .I1(bbar[4])
  );
  //AND U115
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U115 (
    .O(y[227]),
    .I0(a[14]),
    .I1(b[3])
  );
  //OR U115bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U115bar (
    .O(ybar[227]),
    .I0(abar[14]),
    .I1(bbar[3])
  );
  //AND U116
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U116 (
    .O(y[226]),
    .I0(a[14]),
    .I1(b[2])
  );
  //OR U116bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U116bar (
    .O(ybar[226]),
    .I0(abar[14]),
    .I1(bbar[2])
  );
  //AND U117
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U117 (
    .O(y[225]),
    .I0(a[14]),
    .I1(b[1])
  );
  //OR U117bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U117bar (
    .O(ybar[225]),
    .I0(abar[14]),
    .I1(bbar[1])
  );
  //AND U118
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U118 (
    .O(y[224]),
    .I0(a[14]),
    .I1(b[0])
  );
  //OR U118bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U118bar (
    .O(ybar[224]),
    .I0(abar[14]),
    .I1(bbar[0])
  );
  //AND U119
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U119 (
    .O(y[223]),
    .I0(a[13]),
    .I1(b[15])
  );
  //OR U119bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U119bar (
    .O(ybar[223]),
    .I0(abar[13]),
    .I1(bbar[15])
  );
  //AND U120
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U120 (
    .O(y[222]),
    .I0(a[13]),
    .I1(b[14])
  );
  //OR U120bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U120bar (
    .O(ybar[222]),
    .I0(abar[13]),
    .I1(bbar[14])
  );
  //AND U121
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U121 (
    .O(y[221]),
    .I0(a[13]),
    .I1(b[13])
  );
  //OR U121bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U121bar (
    .O(ybar[221]),
    .I0(abar[13]),
    .I1(bbar[13])
  );
  //AND U122
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U122 (
    .O(y[220]),
    .I0(a[13]),
    .I1(b[12])
  );
  //OR U122bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U122bar (
    .O(ybar[220]),
    .I0(abar[13]),
    .I1(bbar[12])
  );
  //AND U123
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U123 (
    .O(y[21]),
    .I0(a[1]),
    .I1(b[5])
  );
  //OR U123bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U123bar (
    .O(ybar[21]),
    .I0(abar[1]),
    .I1(bbar[5])
  );
  //AND U124
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U124 (
    .O(y[219]),
    .I0(a[13]),
    .I1(b[11])
  );
  //OR U124bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U124bar (
    .O(ybar[219]),
    .I0(abar[13]),
    .I1(bbar[11])
  );
  //AND U125
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U125 (
    .O(y[218]),
    .I0(a[13]),
    .I1(b[10])
  );
  //OR U125bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U125bar (
    .O(ybar[218]),
    .I0(abar[13]),
    .I1(bbar[10])
  );
  //AND U126
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U126 (
    .O(y[217]),
    .I0(a[13]),
    .I1(b[9])
  );
  //OR U126bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U126bar (
    .O(ybar[217]),
    .I0(abar[13]),
    .I1(bbar[9])
  );
  //AND U127
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U127 (
    .O(y[216]),
    .I0(a[13]),
    .I1(b[8])
  );
  //OR U127bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U127bar (
    .O(ybar[216]),
    .I0(abar[13]),
    .I1(bbar[8])
  );
  //AND U128
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U128 (
    .O(y[215]),
    .I0(a[13]),
    .I1(b[7])
  );
  //OR U128bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U128bar (
    .O(ybar[215]),
    .I0(abar[13]),
    .I1(bbar[7])
  );
  //AND U129
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U129 (
    .O(y[214]),
    .I0(a[13]),
    .I1(b[6])
  );
  //OR U129bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U129bar (
    .O(ybar[214]),
    .I0(abar[13]),
    .I1(bbar[6])
  );
  //AND U130
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U130 (
    .O(y[213]),
    .I0(a[13]),
    .I1(b[5])
  );
  //OR U130bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U130bar (
    .O(ybar[213]),
    .I0(abar[13]),
    .I1(bbar[5])
  );
  //AND U131
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U131 (
    .O(y[212]),
    .I0(a[13]),
    .I1(b[4])
  );
  //OR U131bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U131bar (
    .O(ybar[212]),
    .I0(abar[13]),
    .I1(bbar[4])
  );
  //AND U132
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U132 (
    .O(y[211]),
    .I0(a[13]),
    .I1(b[3])
  );
  //OR U132bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U132bar (
    .O(ybar[211]),
    .I0(abar[13]),
    .I1(bbar[3])
  );
  //AND U133
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U133 (
    .O(y[210]),
    .I0(a[13]),
    .I1(b[2])
  );
  //OR U133bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U133bar (
    .O(ybar[210]),
    .I0(abar[13]),
    .I1(bbar[2])
  );
  //AND U134
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U134 (
    .O(y[20]),
    .I0(a[1]),
    .I1(b[4])
  );
  //OR U134bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U134bar (
    .O(ybar[20]),
    .I0(abar[1]),
    .I1(bbar[4])
  );
  //AND U135
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U135 (
    .O(y[209]),
    .I0(a[13]),
    .I1(b[1])
  );
  //OR U135bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U135bar (
    .O(ybar[209]),
    .I0(abar[13]),
    .I1(bbar[1])
  );
  //AND U136
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U136 (
    .O(y[208]),
    .I0(a[13]),
    .I1(b[0])
  );
  //OR U136bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U136bar (
    .O(ybar[208]),
    .I0(abar[13]),
    .I1(bbar[0])
  );
  //AND U137
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U137 (
    .O(y[207]),
    .I0(a[12]),
    .I1(b[15])
  );
  //OR U137bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U137bar (
    .O(ybar[207]),
    .I0(abar[12]),
    .I1(bbar[15])
  );
  //AND U138
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U138 (
    .O(y[206]),
    .I0(a[12]),
    .I1(b[14])
  );
  //OR U138bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U138bar (
    .O(ybar[206]),
    .I0(abar[12]),
    .I1(bbar[14])
  );
  //AND U139
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U139 (
    .O(y[205]),
    .I0(a[12]),
    .I1(b[13])
  );
  //OR U139bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U139bar (
    .O(ybar[205]),
    .I0(abar[12]),
    .I1(bbar[13])
  );
  //AND U140
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U140 (
    .O(y[204]),
    .I0(a[12]),
    .I1(b[12])
  );
  //OR U140bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U140bar (
    .O(ybar[204]),
    .I0(abar[12]),
    .I1(bbar[12])
  );
  //AND U141
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U141 (
    .O(y[203]),
    .I0(a[12]),
    .I1(b[11])
  );
  //OR U141bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U141bar (
    .O(ybar[203]),
    .I0(abar[12]),
    .I1(bbar[11])
  );
  //AND U142
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U142 (
    .O(y[202]),
    .I0(a[12]),
    .I1(b[10])
  );
  //OR U142bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U142bar (
    .O(ybar[202]),
    .I0(abar[12]),
    .I1(bbar[10])
  );
  //AND U143
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U143 (
    .O(y[201]),
    .I0(a[12]),
    .I1(b[9])
  );
  //OR U143bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U143bar (
    .O(ybar[201]),
    .I0(abar[12]),
    .I1(bbar[9])
  );
  //AND U144
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U144 (
    .O(y[200]),
    .I0(a[12]),
    .I1(b[8])
  );
  //OR U144bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U144bar (
    .O(ybar[200]),
    .I0(abar[12]),
    .I1(bbar[8])
  );
  //AND U145
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U145 (
    .O(y[1]),
    .I0(b[1]),
    .I1(a[0])
  );
  //OR U145bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U145bar (
    .O(ybar[1]),
    .I0(bbar[1]),
    .I1(abar[0])
  );
  //AND U146
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U146 (
    .O(y[19]),
    .I0(a[1]),
    .I1(b[3])
  );
  //OR U146bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U146bar (
    .O(ybar[19]),
    .I0(abar[1]),
    .I1(bbar[3])
  );
  //AND U147
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U147 (
    .O(y[199]),
    .I0(a[12]),
    .I1(b[7])
  );
  //OR U147bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U147bar (
    .O(ybar[199]),
    .I0(abar[12]),
    .I1(bbar[7])
  );
  //AND U148
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U148 (
    .O(y[198]),
    .I0(a[12]),
    .I1(b[6])
  );
  //OR U148bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U148bar (
    .O(ybar[198]),
    .I0(abar[12]),
    .I1(bbar[6])
  );
  //AND U149
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U149 (
    .O(y[197]),
    .I0(a[12]),
    .I1(b[5])
  );
  //OR U149bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U149bar (
    .O(ybar[197]),
    .I0(abar[12]),
    .I1(bbar[5])
  );
  //AND U150
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U150 (
    .O(y[196]),
    .I0(a[12]),
    .I1(b[4])
  );
  //OR U150bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U150bar (
    .O(ybar[196]),
    .I0(abar[12]),
    .I1(bbar[4])
  );
  //AND U151
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U151 (
    .O(y[195]),
    .I0(a[12]),
    .I1(b[3])
  );
  //OR U151bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U151bar (
    .O(ybar[195]),
    .I0(abar[12]),
    .I1(bbar[3])
  );
  //AND U152
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U152 (
    .O(y[194]),
    .I0(a[12]),
    .I1(b[2])
  );
  //OR U152bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U152bar (
    .O(ybar[194]),
    .I0(abar[12]),
    .I1(bbar[2])
  );
  //AND U153
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U153 (
    .O(y[193]),
    .I0(a[12]),
    .I1(b[1])
  );
  //OR U153bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U153bar (
    .O(ybar[193]),
    .I0(abar[12]),
    .I1(bbar[1])
  );
  //AND U154
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U154 (
    .O(y[192]),
    .I0(a[12]),
    .I1(b[0])
  );
  //OR U154bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U154bar (
    .O(ybar[192]),
    .I0(abar[12]),
    .I1(bbar[0])
  );
  //AND U155
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U155 (
    .O(y[191]),
    .I0(a[11]),
    .I1(b[15])
  );
  //OR U155bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U155bar (
    .O(ybar[191]),
    .I0(abar[11]),
    .I1(bbar[15])
  );
  //AND U156
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U156 (
    .O(y[190]),
    .I0(a[11]),
    .I1(b[14])
  );
  //OR U156bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U156bar (
    .O(ybar[190]),
    .I0(abar[11]),
    .I1(bbar[14])
  );
  //AND U157
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U157 (
    .O(y[18]),
    .I0(a[1]),
    .I1(b[2])
  );
  //OR U157bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U157bar (
    .O(ybar[18]),
    .I0(abar[1]),
    .I1(bbar[2])
  );
  //AND U158
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U158 (
    .O(y[189]),
    .I0(a[11]),
    .I1(b[13])
  );
  //OR U158bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U158bar (
    .O(ybar[189]),
    .I0(abar[11]),
    .I1(bbar[13])
  );
  //AND U159
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U159 (
    .O(y[188]),
    .I0(a[11]),
    .I1(b[12])
  );
  //OR U159bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U159bar (
    .O(ybar[188]),
    .I0(abar[11]),
    .I1(bbar[12])
  );
  //AND U160
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U160 (
    .O(y[187]),
    .I0(a[11]),
    .I1(b[11])
  );
  //OR U160bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U160bar (
    .O(ybar[187]),
    .I0(abar[11]),
    .I1(bbar[11])
  );
  //AND U161
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U161 (
    .O(y[186]),
    .I0(a[11]),
    .I1(b[10])
  );
  //OR U161bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U161bar (
    .O(ybar[186]),
    .I0(abar[11]),
    .I1(bbar[10])
  );
  //AND U162
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U162 (
    .O(y[185]),
    .I0(a[11]),
    .I1(b[9])
  );
  //OR U162bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U162bar (
    .O(ybar[185]),
    .I0(abar[11]),
    .I1(bbar[9])
  );
  //AND U163
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U163 (
    .O(y[184]),
    .I0(a[11]),
    .I1(b[8])
  );
  //OR U163bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U163bar (
    .O(ybar[184]),
    .I0(abar[11]),
    .I1(bbar[8])
  );
  //AND U164
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U164 (
    .O(y[183]),
    .I0(a[11]),
    .I1(b[7])
  );
  //OR U164bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U164bar (
    .O(ybar[183]),
    .I0(abar[11]),
    .I1(bbar[7])
  );
  //AND U165
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U165 (
    .O(y[182]),
    .I0(a[11]),
    .I1(b[6])
  );
  //OR U165bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U165bar (
    .O(ybar[182]),
    .I0(abar[11]),
    .I1(bbar[6])
  );
  //AND U166
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U166 (
    .O(y[181]),
    .I0(a[11]),
    .I1(b[5])
  );
  //OR U166bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U166bar (
    .O(ybar[181]),
    .I0(abar[11]),
    .I1(bbar[5])
  );
  //AND U167
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U167 (
    .O(y[180]),
    .I0(a[11]),
    .I1(b[4])
  );
  //OR U167bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U167bar (
    .O(ybar[180]),
    .I0(abar[11]),
    .I1(bbar[4])
  );
  //AND U168
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U168 (
    .O(y[17]),
    .I0(a[1]),
    .I1(b[1])
  );
  //OR U168bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U168bar (
    .O(ybar[17]),
    .I0(abar[1]),
    .I1(bbar[1])
  );
  //AND U169
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U169 (
    .O(y[179]),
    .I0(a[11]),
    .I1(b[3])
  );
  //OR U169bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U169bar (
    .O(ybar[179]),
    .I0(abar[11]),
    .I1(bbar[3])
  );
  //AND U170
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U170 (
    .O(y[178]),
    .I0(a[11]),
    .I1(b[2])
  );
  //OR U170bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U170bar (
    .O(ybar[178]),
    .I0(abar[11]),
    .I1(bbar[2])
  );
  //AND U171
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U171 (
    .O(y[177]),
    .I0(a[11]),
    .I1(b[1])
  );
  //OR U171bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U171bar (
    .O(ybar[177]),
    .I0(abar[11]),
    .I1(bbar[1])
  );
  //AND U172
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U172 (
    .O(y[176]),
    .I0(a[11]),
    .I1(b[0])
  );
  //OR U172bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U172bar (
    .O(ybar[176]),
    .I0(abar[11]),
    .I1(bbar[0])
  );
  //AND U173
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U173 (
    .O(y[175]),
    .I0(a[10]),
    .I1(b[15])
  );
  //OR U173bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U173bar (
    .O(ybar[175]),
    .I0(abar[10]),
    .I1(bbar[15])
  );
  //AND U174
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U174 (
    .O(y[174]),
    .I0(a[10]),
    .I1(b[14])
  );
  //OR U174bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U174bar (
    .O(ybar[174]),
    .I0(abar[10]),
    .I1(bbar[14])
  );
  //AND U175
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U175 (
    .O(y[173]),
    .I0(a[10]),
    .I1(b[13])
  );
  //OR U175bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U175bar (
    .O(ybar[173]),
    .I0(abar[10]),
    .I1(bbar[13])
  );
  //AND U176
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U176 (
    .O(y[172]),
    .I0(a[10]),
    .I1(b[12])
  );
  //OR U176bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U176bar (
    .O(ybar[172]),
    .I0(abar[10]),
    .I1(bbar[12])
  );
  //AND U177
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U177 (
    .O(y[171]),
    .I0(a[10]),
    .I1(b[11])
  );
  //OR U177bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U177bar (
    .O(ybar[171]),
    .I0(abar[10]),
    .I1(bbar[11])
  );
  //AND U178
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U178 (
    .O(y[170]),
    .I0(a[10]),
    .I1(b[10])
  );
  //OR U178bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U178bar (
    .O(ybar[170]),
    .I0(abar[10]),
    .I1(bbar[10])
  );
  //AND U179
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U179 (
    .O(y[16]),
    .I0(a[1]),
    .I1(b[0])
  );
  //OR U179bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U179bar (
    .O(ybar[16]),
    .I0(abar[1]),
    .I1(bbar[0])
  );
  //AND U180
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U180 (
    .O(y[169]),
    .I0(a[10]),
    .I1(b[9])
  );
  //OR U180bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U180bar (
    .O(ybar[169]),
    .I0(abar[10]),
    .I1(bbar[9])
  );
  //AND U181
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U181 (
    .O(y[168]),
    .I0(a[10]),
    .I1(b[8])
  );
  //OR U181bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U181bar (
    .O(ybar[168]),
    .I0(abar[10]),
    .I1(bbar[8])
  );
  //AND U182
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U182 (
    .O(y[167]),
    .I0(a[10]),
    .I1(b[7])
  );
  //OR U182bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U182bar (
    .O(ybar[167]),
    .I0(abar[10]),
    .I1(bbar[7])
  );
  //AND U183
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U183 (
    .O(y[166]),
    .I0(a[10]),
    .I1(b[6])
  );
  //OR U183bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U183bar (
    .O(ybar[166]),
    .I0(abar[10]),
    .I1(bbar[6])
  );
  //AND U184
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U184 (
    .O(y[165]),
    .I0(a[10]),
    .I1(b[5])
  );
  //OR U184bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U184bar (
    .O(ybar[165]),
    .I0(abar[10]),
    .I1(bbar[5])
  );
  //AND U185
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U185 (
    .O(y[164]),
    .I0(a[10]),
    .I1(b[4])
  );
  //OR U185bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U185bar (
    .O(ybar[164]),
    .I0(abar[10]),
    .I1(bbar[4])
  );
  //AND U186
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U186 (
    .O(y[163]),
    .I0(a[10]),
    .I1(b[3])
  );
  //OR U186bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U186bar (
    .O(ybar[163]),
    .I0(abar[10]),
    .I1(bbar[3])
  );
  //AND U187
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U187 (
    .O(y[162]),
    .I0(a[10]),
    .I1(b[2])
  );
  //OR U187bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U187bar (
    .O(ybar[162]),
    .I0(abar[10]),
    .I1(bbar[2])
  );
  //AND U188
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U188 (
    .O(y[161]),
    .I0(a[10]),
    .I1(b[1])
  );
  //OR U188bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U188bar (
    .O(ybar[161]),
    .I0(abar[10]),
    .I1(bbar[1])
  );
  //AND U189
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U189 (
    .O(y[160]),
    .I0(a[10]),
    .I1(b[0])
  );
  //OR U189bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U189bar (
    .O(ybar[160]),
    .I0(abar[10]),
    .I1(bbar[0])
  );
  //AND U190
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U190 (
    .O(y[15]),
    .I0(b[15]),
    .I1(a[0])
  );
  //OR U190bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U190bar (
    .O(ybar[15]),
    .I0(bbar[15]),
    .I1(abar[0])
  );
  //AND U191
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U191 (
    .O(y[159]),
    .I0(a[9]),
    .I1(b[15])
  );
  //OR U191bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U191bar (
    .O(ybar[159]),
    .I0(abar[9]),
    .I1(bbar[15])
  );
  //AND U192
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U192 (
    .O(y[158]),
    .I0(a[9]),
    .I1(b[14])
  );
  //OR U192bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U192bar (
    .O(ybar[158]),
    .I0(abar[9]),
    .I1(bbar[14])
  );
  //AND U193
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U193 (
    .O(y[157]),
    .I0(a[9]),
    .I1(b[13])
  );
  //OR U193bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U193bar (
    .O(ybar[157]),
    .I0(abar[9]),
    .I1(bbar[13])
  );
  //AND U194
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U194 (
    .O(y[156]),
    .I0(a[9]),
    .I1(b[12])
  );
  //OR U194bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U194bar (
    .O(ybar[156]),
    .I0(abar[9]),
    .I1(bbar[12])
  );
  //AND U195
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U195 (
    .O(y[155]),
    .I0(a[9]),
    .I1(b[11])
  );
  //OR U195bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U195bar (
    .O(ybar[155]),
    .I0(abar[9]),
    .I1(bbar[11])
  );
  //AND U196
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U196 (
    .O(y[154]),
    .I0(a[9]),
    .I1(b[10])
  );
  //OR U196bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U196bar (
    .O(ybar[154]),
    .I0(abar[9]),
    .I1(bbar[10])
  );
  //AND U197
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U197 (
    .O(y[153]),
    .I0(a[9]),
    .I1(b[9])
  );
  //OR U197bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U197bar (
    .O(ybar[153]),
    .I0(abar[9]),
    .I1(bbar[9])
  );
  //AND U198
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U198 (
    .O(y[152]),
    .I0(a[9]),
    .I1(b[8])
  );
  //OR U198bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U198bar (
    .O(ybar[152]),
    .I0(abar[9]),
    .I1(bbar[8])
  );
  //AND U199
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U199 (
    .O(y[151]),
    .I0(a[9]),
    .I1(b[7])
  );
  //OR U199bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U199bar (
    .O(ybar[151]),
    .I0(abar[9]),
    .I1(bbar[7])
  );
  //AND U200
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U200 (
    .O(y[150]),
    .I0(a[9]),
    .I1(b[6])
  );
  //OR U200bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U200bar (
    .O(ybar[150]),
    .I0(abar[9]),
    .I1(bbar[6])
  );
  //AND U201
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U201 (
    .O(y[14]),
    .I0(b[14]),
    .I1(a[0])
  );
  //OR U201bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U201bar (
    .O(ybar[14]),
    .I0(bbar[14]),
    .I1(abar[0])
  );
  //AND U202
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U202 (
    .O(y[149]),
    .I0(a[9]),
    .I1(b[5])
  );
  //OR U202bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U202bar (
    .O(ybar[149]),
    .I0(abar[9]),
    .I1(bbar[5])
  );
  //AND U203
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U203 (
    .O(y[148]),
    .I0(a[9]),
    .I1(b[4])
  );
  //OR U203bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U203bar (
    .O(ybar[148]),
    .I0(abar[9]),
    .I1(bbar[4])
  );
  //AND U204
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U204 (
    .O(y[147]),
    .I0(a[9]),
    .I1(b[3])
  );
  //OR U204bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U204bar (
    .O(ybar[147]),
    .I0(abar[9]),
    .I1(bbar[3])
  );
  //AND U205
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U205 (
    .O(y[146]),
    .I0(a[9]),
    .I1(b[2])
  );
  //OR U205bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U205bar (
    .O(ybar[146]),
    .I0(abar[9]),
    .I1(bbar[2])
  );
  //AND U206
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U206 (
    .O(y[145]),
    .I0(a[9]),
    .I1(b[1])
  );
  //OR U206bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U206bar (
    .O(ybar[145]),
    .I0(abar[9]),
    .I1(bbar[1])
  );
  //AND U207
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U207 (
    .O(y[144]),
    .I0(a[9]),
    .I1(b[0])
  );
  //OR U207bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U207bar (
    .O(ybar[144]),
    .I0(abar[9]),
    .I1(bbar[0])
  );
  //AND U208
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U208 (
    .O(y[143]),
    .I0(a[8]),
    .I1(b[15])
  );
  //OR U208bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U208bar (
    .O(ybar[143]),
    .I0(abar[8]),
    .I1(bbar[15])
  );
  //AND U209
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U209 (
    .O(y[142]),
    .I0(a[8]),
    .I1(b[14])
  );
  //OR U209bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U209bar (
    .O(ybar[142]),
    .I0(abar[8]),
    .I1(bbar[14])
  );
  //AND U210
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U210 (
    .O(y[141]),
    .I0(a[8]),
    .I1(b[13])
  );
  //OR U210bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U210bar (
    .O(ybar[141]),
    .I0(abar[8]),
    .I1(bbar[13])
  );
  //AND U211
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U211 (
    .O(y[140]),
    .I0(a[8]),
    .I1(b[12])
  );
  //OR U211bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U211bar (
    .O(ybar[140]),
    .I0(abar[8]),
    .I1(bbar[12])
  );
  //AND U212
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U212 (
    .O(y[13]),
    .I0(b[13]),
    .I1(a[0])
  );
  //OR U212bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U212bar (
    .O(ybar[13]),
    .I0(bbar[13]),
    .I1(abar[0])
  );
  //AND U213
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U213 (
    .O(y[139]),
    .I0(a[8]),
    .I1(b[11])
  );
  //OR U213bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U213bar (
    .O(ybar[139]),
    .I0(abar[8]),
    .I1(bbar[11])
  );
  //AND U214
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U214 (
    .O(y[138]),
    .I0(a[8]),
    .I1(b[10])
  );
  //OR U214bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U214bar (
    .O(ybar[138]),
    .I0(abar[8]),
    .I1(bbar[10])
  );
  //AND U215
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U215 (
    .O(y[137]),
    .I0(a[8]),
    .I1(b[9])
  );
  //OR U215bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U215bar (
    .O(ybar[137]),
    .I0(abar[8]),
    .I1(bbar[9])
  );
  //AND U216
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U216 (
    .O(y[136]),
    .I0(a[8]),
    .I1(b[8])
  );
  //OR U216bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U216bar (
    .O(ybar[136]),
    .I0(abar[8]),
    .I1(bbar[8])
  );
  //AND U217
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U217 (
    .O(y[135]),
    .I0(a[8]),
    .I1(b[7])
  );
  //OR U217bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U217bar (
    .O(ybar[135]),
    .I0(abar[8]),
    .I1(bbar[7])
  );
  //AND U218
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U218 (
    .O(y[134]),
    .I0(a[8]),
    .I1(b[6])
  );
  //OR U218bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U218bar (
    .O(ybar[134]),
    .I0(abar[8]),
    .I1(bbar[6])
  );
  //AND U219
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U219 (
    .O(y[133]),
    .I0(a[8]),
    .I1(b[5])
  );
  //OR U219bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U219bar (
    .O(ybar[133]),
    .I0(abar[8]),
    .I1(bbar[5])
  );
  //AND U220
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U220 (
    .O(y[132]),
    .I0(a[8]),
    .I1(b[4])
  );
  //OR U220bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U220bar (
    .O(ybar[132]),
    .I0(abar[8]),
    .I1(bbar[4])
  );
  //AND U221
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U221 (
    .O(y[131]),
    .I0(a[8]),
    .I1(b[3])
  );
  //OR U221bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U221bar (
    .O(ybar[131]),
    .I0(abar[8]),
    .I1(bbar[3])
  );
  //AND U222
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U222 (
    .O(y[130]),
    .I0(a[8]),
    .I1(b[2])
  );
  //OR U222bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U222bar (
    .O(ybar[130]),
    .I0(abar[8]),
    .I1(bbar[2])
  );
  //AND U223
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U223 (
    .O(y[12]),
    .I0(b[12]),
    .I1(a[0])
  );
  //OR U223bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U223bar (
    .O(ybar[12]),
    .I0(bbar[12]),
    .I1(abar[0])
  );
  //AND U224
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U224 (
    .O(y[129]),
    .I0(a[8]),
    .I1(b[1])
  );
  //OR U224bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U224bar (
    .O(ybar[129]),
    .I0(abar[8]),
    .I1(bbar[1])
  );
  //AND U225
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U225 (
    .O(y[128]),
    .I0(a[8]),
    .I1(b[0])
  );
  //OR U225bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U225bar (
    .O(ybar[128]),
    .I0(abar[8]),
    .I1(bbar[0])
  );
  //AND U226
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U226 (
    .O(y[127]),
    .I0(a[7]),
    .I1(b[15])
  );
  //OR U226bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U226bar (
    .O(ybar[127]),
    .I0(abar[7]),
    .I1(bbar[15])
  );
  //AND U227
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U227 (
    .O(y[126]),
    .I0(a[7]),
    .I1(b[14])
  );
  //OR U227bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U227bar (
    .O(ybar[126]),
    .I0(abar[7]),
    .I1(bbar[14])
  );
  //AND U228
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U228 (
    .O(y[125]),
    .I0(a[7]),
    .I1(b[13])
  );
  //OR U228bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U228bar (
    .O(ybar[125]),
    .I0(abar[7]),
    .I1(bbar[13])
  );
  //AND U229
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U229 (
    .O(y[124]),
    .I0(a[7]),
    .I1(b[12])
  );
  //OR U229bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U229bar (
    .O(ybar[124]),
    .I0(abar[7]),
    .I1(bbar[12])
  );
  //AND U230
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U230 (
    .O(y[123]),
    .I0(a[7]),
    .I1(b[11])
  );
  //OR U230bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U230bar (
    .O(ybar[123]),
    .I0(abar[7]),
    .I1(bbar[11])
  );
  //AND U231
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U231 (
    .O(y[122]),
    .I0(a[7]),
    .I1(b[10])
  );
  //OR U231bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U231bar (
    .O(ybar[122]),
    .I0(abar[7]),
    .I1(bbar[10])
  );
  //AND U232
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U232 (
    .O(y[121]),
    .I0(a[7]),
    .I1(b[9])
  );
  //OR U232bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U232bar (
    .O(ybar[121]),
    .I0(abar[7]),
    .I1(bbar[9])
  );
  //AND U233
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U233 (
    .O(y[120]),
    .I0(a[7]),
    .I1(b[8])
  );
  //OR U233bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U233bar (
    .O(ybar[120]),
    .I0(abar[7]),
    .I1(bbar[8])
  );
  //AND U234
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U234 (
    .O(y[11]),
    .I0(b[11]),
    .I1(a[0])
  );
  //OR U234bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U234bar (
    .O(ybar[11]),
    .I0(bbar[11]),
    .I1(abar[0])
  );
  //AND U235
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U235 (
    .O(y[119]),
    .I0(a[7]),
    .I1(b[7])
  );
  //OR U235bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U235bar (
    .O(ybar[119]),
    .I0(abar[7]),
    .I1(bbar[7])
  );
  //AND U236
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U236 (
    .O(y[118]),
    .I0(a[7]),
    .I1(b[6])
  );
  //OR U236bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U236bar (
    .O(ybar[118]),
    .I0(abar[7]),
    .I1(bbar[6])
  );
  //AND U237
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U237 (
    .O(y[117]),
    .I0(a[7]),
    .I1(b[5])
  );
  //OR U237bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U237bar (
    .O(ybar[117]),
    .I0(abar[7]),
    .I1(bbar[5])
  );
  //AND U238
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U238 (
    .O(y[116]),
    .I0(a[7]),
    .I1(b[4])
  );
  //OR U238bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U238bar (
    .O(ybar[116]),
    .I0(abar[7]),
    .I1(bbar[4])
  );
  //AND U239
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U239 (
    .O(y[115]),
    .I0(a[7]),
    .I1(b[3])
  );
  //OR U239bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U239bar (
    .O(ybar[115]),
    .I0(abar[7]),
    .I1(bbar[3])
  );
  //AND U240
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U240 (
    .O(y[114]),
    .I0(a[7]),
    .I1(b[2])
  );
  //OR U240bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U240bar (
    .O(ybar[114]),
    .I0(abar[7]),
    .I1(bbar[2])
  );
  //AND U241
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U241 (
    .O(y[113]),
    .I0(a[7]),
    .I1(b[1])
  );
  //OR U241bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U241bar (
    .O(ybar[113]),
    .I0(abar[7]),
    .I1(bbar[1])
  );
  //AND U242
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U242 (
    .O(y[112]),
    .I0(a[7]),
    .I1(b[0])
  );
  //OR U242bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U242bar (
    .O(ybar[112]),
    .I0(abar[7]),
    .I1(bbar[0])
  );
  //AND U243
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U243 (
    .O(y[111]),
    .I0(b[15]),
    .I1(a[6])
  );
  //OR U243bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U243bar (
    .O(ybar[111]),
    .I0(bbar[15]),
    .I1(abar[6])
  );
  //AND U244
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U244 (
    .O(y[110]),
    .I0(b[14]),
    .I1(a[6])
  );
  //OR U244bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U244bar (
    .O(ybar[110]),
    .I0(bbar[14]),
    .I1(abar[6])
  );
  //AND U245
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U245 (
    .O(y[10]),
    .I0(b[10]),
    .I1(a[0])
  );
  //OR U245bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U245bar (
    .O(ybar[10]),
    .I0(bbar[10]),
    .I1(abar[0])
  );
  //AND U246
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U246 (
    .O(y[109]),
    .I0(b[13]),
    .I1(a[6])
  );
  //OR U246bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U246bar (
    .O(ybar[109]),
    .I0(bbar[13]),
    .I1(abar[6])
  );
  //AND U247
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U247 (
    .O(y[108]),
    .I0(b[12]),
    .I1(a[6])
  );
  //OR U247bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U247bar (
    .O(ybar[108]),
    .I0(bbar[12]),
    .I1(abar[6])
  );
  //AND U248
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U248 (
    .O(y[107]),
    .I0(b[11]),
    .I1(a[6])
  );
  //OR U248bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U248bar (
    .O(ybar[107]),
    .I0(bbar[11]),
    .I1(abar[6])
  );
  //AND U249
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U249 (
    .O(y[106]),
    .I0(b[10]),
    .I1(a[6])
  );
  //OR U249bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U249bar (
    .O(ybar[106]),
    .I0(bbar[10]),
    .I1(abar[6])
  );
  //AND U250
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U250 (
    .O(y[105]),
    .I0(a[6]),
    .I1(b[9])
  );
  //OR U250bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U250bar (
    .O(ybar[105]),
    .I0(abar[6]),
    .I1(bbar[9])
  );
  //AND U251
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U251 (
    .O(y[104]),
    .I0(b[8]),
    .I1(a[6])
  );
  //OR U251bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U251bar (
    .O(ybar[104]),
    .I0(bbar[8]),
    .I1(abar[6])
  );
  //AND U252
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U252 (
    .O(y[103]),
    .I0(b[7]),
    .I1(a[6])
  );
  //OR U252bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U252bar (
    .O(ybar[103]),
    .I0(bbar[7]),
    .I1(abar[6])
  );
  //AND U253
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U253 (
    .O(y[102]),
    .I0(b[6]),
    .I1(a[6])
  );
  //OR U253bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U253bar (
    .O(ybar[102]),
    .I0(bbar[6]),
    .I1(abar[6])
  );
  //AND U254
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U254 (
    .O(y[101]),
    .I0(b[5]),
    .I1(a[6])
  );
  //OR U254bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U254bar (
    .O(ybar[101]),
    .I0(bbar[5]),
    .I1(abar[6])
  );
  //AND U255
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U255 (
    .O(y[100]),
    .I0(b[4]),
    .I1(a[6])
  );
  //OR U255bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U255bar (
    .O(ybar[100]),
    .I0(bbar[4]),
    .I1(abar[6])
  );
  //AND U256
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U256 (
    .O(y[0]),
    .I0(b[0]),
    .I1(a[0])
  );
  //OR U256bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U256bar (
    .O(ybar[0]),
    .I0(bbar[0]),
    .I1(abar[0])
  );
endmodule

module decode_5 ( in, out );

  input wire [7:0] in;
//input_done

  output wire [255:0] out;
//output_done

  wire [15:0] level1;
  wire [31:0] level2;
//wire_done

  CD2_20 cd_l1_1 ( .a(in[1]), .b(in[0]), .y(level1[3:0]) );
  CD2_19 cd_l1_2 ( .a(in[3]), .b(in[2]), .y(level1[7:4]) );
  CD2_18 cd_l1_3 ( .a(in[5]), .b(in[4]), .y(level1[11:8]) );
  CD2_17 cd_l1_4 ( .a(in[7]), .b(in[6]), .y(level1[15:12]) );
  CD4_10 cd_l2_1 ( .a(level1[7:4]), .b(level1[3:0]), .y(level2[15:0]) );
  CD4_9 cd_l2_2 ( .a(level1[15:12]), .b(level1[11:8]), .y(level2[31:16]) );
  CD16_5 cd_l3 ( .a(level2[31:16]), .b(level2[15:0]), .y(out) );
endmodule

module encode_5 ( in, out );

  input wire [255:0] in;
  wire [255:0] inbar;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
  assign inbar[8] = ~in[8];
  assign inbar[9] = ~in[9];
  assign inbar[10] = ~in[10];
  assign inbar[11] = ~in[11];
  assign inbar[12] = ~in[12];
  assign inbar[13] = ~in[13];
  assign inbar[14] = ~in[14];
  assign inbar[15] = ~in[15];
  assign inbar[16] = ~in[16];
  assign inbar[17] = ~in[17];
  assign inbar[18] = ~in[18];
  assign inbar[19] = ~in[19];
  assign inbar[20] = ~in[20];
  assign inbar[21] = ~in[21];
  assign inbar[22] = ~in[22];
  assign inbar[23] = ~in[23];
  assign inbar[24] = ~in[24];
  assign inbar[25] = ~in[25];
  assign inbar[26] = ~in[26];
  assign inbar[27] = ~in[27];
  assign inbar[28] = ~in[28];
  assign inbar[29] = ~in[29];
  assign inbar[30] = ~in[30];
  assign inbar[31] = ~in[31];
  assign inbar[32] = ~in[32];
  assign inbar[33] = ~in[33];
  assign inbar[34] = ~in[34];
  assign inbar[35] = ~in[35];
  assign inbar[36] = ~in[36];
  assign inbar[37] = ~in[37];
  assign inbar[38] = ~in[38];
  assign inbar[39] = ~in[39];
  assign inbar[40] = ~in[40];
  assign inbar[41] = ~in[41];
  assign inbar[42] = ~in[42];
  assign inbar[43] = ~in[43];
  assign inbar[44] = ~in[44];
  assign inbar[45] = ~in[45];
  assign inbar[46] = ~in[46];
  assign inbar[47] = ~in[47];
  assign inbar[48] = ~in[48];
  assign inbar[49] = ~in[49];
  assign inbar[50] = ~in[50];
  assign inbar[51] = ~in[51];
  assign inbar[52] = ~in[52];
  assign inbar[53] = ~in[53];
  assign inbar[54] = ~in[54];
  assign inbar[55] = ~in[55];
  assign inbar[56] = ~in[56];
  assign inbar[57] = ~in[57];
  assign inbar[58] = ~in[58];
  assign inbar[59] = ~in[59];
  assign inbar[60] = ~in[60];
  assign inbar[61] = ~in[61];
  assign inbar[62] = ~in[62];
  assign inbar[63] = ~in[63];
  assign inbar[64] = ~in[64];
  assign inbar[65] = ~in[65];
  assign inbar[66] = ~in[66];
  assign inbar[67] = ~in[67];
  assign inbar[68] = ~in[68];
  assign inbar[69] = ~in[69];
  assign inbar[70] = ~in[70];
  assign inbar[71] = ~in[71];
  assign inbar[72] = ~in[72];
  assign inbar[73] = ~in[73];
  assign inbar[74] = ~in[74];
  assign inbar[75] = ~in[75];
  assign inbar[76] = ~in[76];
  assign inbar[77] = ~in[77];
  assign inbar[78] = ~in[78];
  assign inbar[79] = ~in[79];
  assign inbar[80] = ~in[80];
  assign inbar[81] = ~in[81];
  assign inbar[82] = ~in[82];
  assign inbar[83] = ~in[83];
  assign inbar[84] = ~in[84];
  assign inbar[85] = ~in[85];
  assign inbar[86] = ~in[86];
  assign inbar[87] = ~in[87];
  assign inbar[88] = ~in[88];
  assign inbar[89] = ~in[89];
  assign inbar[90] = ~in[90];
  assign inbar[91] = ~in[91];
  assign inbar[92] = ~in[92];
  assign inbar[93] = ~in[93];
  assign inbar[94] = ~in[94];
  assign inbar[95] = ~in[95];
  assign inbar[96] = ~in[96];
  assign inbar[97] = ~in[97];
  assign inbar[98] = ~in[98];
  assign inbar[99] = ~in[99];
  assign inbar[100] = ~in[100];
  assign inbar[101] = ~in[101];
  assign inbar[102] = ~in[102];
  assign inbar[103] = ~in[103];
  assign inbar[104] = ~in[104];
  assign inbar[105] = ~in[105];
  assign inbar[106] = ~in[106];
  assign inbar[107] = ~in[107];
  assign inbar[108] = ~in[108];
  assign inbar[109] = ~in[109];
  assign inbar[110] = ~in[110];
  assign inbar[111] = ~in[111];
  assign inbar[112] = ~in[112];
  assign inbar[113] = ~in[113];
  assign inbar[114] = ~in[114];
  assign inbar[115] = ~in[115];
  assign inbar[116] = ~in[116];
  assign inbar[117] = ~in[117];
  assign inbar[118] = ~in[118];
  assign inbar[119] = ~in[119];
  assign inbar[120] = ~in[120];
  assign inbar[121] = ~in[121];
  assign inbar[122] = ~in[122];
  assign inbar[123] = ~in[123];
  assign inbar[124] = ~in[124];
  assign inbar[125] = ~in[125];
  assign inbar[126] = ~in[126];
  assign inbar[127] = ~in[127];
  assign inbar[128] = ~in[128];
  assign inbar[129] = ~in[129];
  assign inbar[130] = ~in[130];
  assign inbar[131] = ~in[131];
  assign inbar[132] = ~in[132];
  assign inbar[133] = ~in[133];
  assign inbar[134] = ~in[134];
  assign inbar[135] = ~in[135];
  assign inbar[136] = ~in[136];
  assign inbar[137] = ~in[137];
  assign inbar[138] = ~in[138];
  assign inbar[139] = ~in[139];
  assign inbar[140] = ~in[140];
  assign inbar[141] = ~in[141];
  assign inbar[142] = ~in[142];
  assign inbar[143] = ~in[143];
  assign inbar[144] = ~in[144];
  assign inbar[145] = ~in[145];
  assign inbar[146] = ~in[146];
  assign inbar[147] = ~in[147];
  assign inbar[148] = ~in[148];
  assign inbar[149] = ~in[149];
  assign inbar[150] = ~in[150];
  assign inbar[151] = ~in[151];
  assign inbar[152] = ~in[152];
  assign inbar[153] = ~in[153];
  assign inbar[154] = ~in[154];
  assign inbar[155] = ~in[155];
  assign inbar[156] = ~in[156];
  assign inbar[157] = ~in[157];
  assign inbar[158] = ~in[158];
  assign inbar[159] = ~in[159];
  assign inbar[160] = ~in[160];
  assign inbar[161] = ~in[161];
  assign inbar[162] = ~in[162];
  assign inbar[163] = ~in[163];
  assign inbar[164] = ~in[164];
  assign inbar[165] = ~in[165];
  assign inbar[166] = ~in[166];
  assign inbar[167] = ~in[167];
  assign inbar[168] = ~in[168];
  assign inbar[169] = ~in[169];
  assign inbar[170] = ~in[170];
  assign inbar[171] = ~in[171];
  assign inbar[172] = ~in[172];
  assign inbar[173] = ~in[173];
  assign inbar[174] = ~in[174];
  assign inbar[175] = ~in[175];
  assign inbar[176] = ~in[176];
  assign inbar[177] = ~in[177];
  assign inbar[178] = ~in[178];
  assign inbar[179] = ~in[179];
  assign inbar[180] = ~in[180];
  assign inbar[181] = ~in[181];
  assign inbar[182] = ~in[182];
  assign inbar[183] = ~in[183];
  assign inbar[184] = ~in[184];
  assign inbar[185] = ~in[185];
  assign inbar[186] = ~in[186];
  assign inbar[187] = ~in[187];
  assign inbar[188] = ~in[188];
  assign inbar[189] = ~in[189];
  assign inbar[190] = ~in[190];
  assign inbar[191] = ~in[191];
  assign inbar[192] = ~in[192];
  assign inbar[193] = ~in[193];
  assign inbar[194] = ~in[194];
  assign inbar[195] = ~in[195];
  assign inbar[196] = ~in[196];
  assign inbar[197] = ~in[197];
  assign inbar[198] = ~in[198];
  assign inbar[199] = ~in[199];
  assign inbar[200] = ~in[200];
  assign inbar[201] = ~in[201];
  assign inbar[202] = ~in[202];
  assign inbar[203] = ~in[203];
  assign inbar[204] = ~in[204];
  assign inbar[205] = ~in[205];
  assign inbar[206] = ~in[206];
  assign inbar[207] = ~in[207];
  assign inbar[208] = ~in[208];
  assign inbar[209] = ~in[209];
  assign inbar[210] = ~in[210];
  assign inbar[211] = ~in[211];
  assign inbar[212] = ~in[212];
  assign inbar[213] = ~in[213];
  assign inbar[214] = ~in[214];
  assign inbar[215] = ~in[215];
  assign inbar[216] = ~in[216];
  assign inbar[217] = ~in[217];
  assign inbar[218] = ~in[218];
  assign inbar[219] = ~in[219];
  assign inbar[220] = ~in[220];
  assign inbar[221] = ~in[221];
  assign inbar[222] = ~in[222];
  assign inbar[223] = ~in[223];
  assign inbar[224] = ~in[224];
  assign inbar[225] = ~in[225];
  assign inbar[226] = ~in[226];
  assign inbar[227] = ~in[227];
  assign inbar[228] = ~in[228];
  assign inbar[229] = ~in[229];
  assign inbar[230] = ~in[230];
  assign inbar[231] = ~in[231];
  assign inbar[232] = ~in[232];
  assign inbar[233] = ~in[233];
  assign inbar[234] = ~in[234];
  assign inbar[235] = ~in[235];
  assign inbar[236] = ~in[236];
  assign inbar[237] = ~in[237];
  assign inbar[238] = ~in[238];
  assign inbar[239] = ~in[239];
  assign inbar[240] = ~in[240];
  assign inbar[241] = ~in[241];
  assign inbar[242] = ~in[242];
  assign inbar[243] = ~in[243];
  assign inbar[244] = ~in[244];
  assign inbar[245] = ~in[245];
  assign inbar[246] = ~in[246];
  assign inbar[247] = ~in[247];
  assign inbar[248] = ~in[248];
  assign inbar[249] = ~in[249];
  assign inbar[250] = ~in[250];
  assign inbar[251] = ~in[251];
  assign inbar[252] = ~in[252];
  assign inbar[253] = ~in[253];
  assign inbar[254] = ~in[254];
  assign inbar[255] = ~in[255];
//input_done

  output wire [7:0] out;
  wire [7:0] outbar;
//output_done

  wire in_81;
  wire in_80;
  wire in_79;
  wire in_78;
  wire in_77;
  wire in_76;
  wire in_75;
  wire in_74;
  wire in_73;
  wire in_72;
  wire in_71;
  wire in_70;
  wire in_69;
  wire in_68;
  wire in_67;
  wire in_66;
  wire in_65;
  wire in_64;
  wire in_63;
  wire in_62;
  wire in_61;
  wire in_60;
  wire in_59;
  wire in_58;
  wire in_57;
  wire in_56;
  wire in_55;
  wire in_54;
  wire in_53;
  wire in_52;
  wire in_51;
  wire in_50;
  wire in_49;
  wire in_48;
  wire in_47;
  wire in_46;
  wire in_45;
  wire in_44;
  wire in_43;
  wire in_42;
  wire in_41;
  wire in_40;
  wire in_39;
  wire in_38;
  wire in_37;
  wire in_36;
  wire in_35;
  wire in_34;
  wire in_33;
  wire in_32;
  wire in_31;
  wire in_30;
  wire in_29;
  wire in_28;
  wire in_27;
  wire in_26;
  wire in_25;
  wire in_24;
  wire in_23;
  wire in_22;
  wire in_21;
  wire in_20;
  wire in_19;
  wire in_18;
  wire in_17;
  wire in_16;
  wire in_15;
  wire in_14;
  wire in_13;
  wire in_12;
  wire in_11;
  wire in_10;
  wire in_9;
  wire in_8;
  wire in_7;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_3;
  wire in_2;
  wire in_1;
  wire in_0;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire in_81bar;
  wire in_80bar;
  wire in_79bar;
  wire in_78bar;
  wire in_77bar;
  wire in_76bar;
  wire in_75bar;
  wire in_74bar;
  wire in_73bar;
  wire in_72bar;
  wire in_71bar;
  wire in_70bar;
  wire in_69bar;
  wire in_68bar;
  wire in_67bar;
  wire in_66bar;
  wire in_65bar;
  wire in_64bar;
  wire in_63bar;
  wire in_62bar;
  wire in_61bar;
  wire in_60bar;
  wire in_59bar;
  wire in_58bar;
  wire in_57bar;
  wire in_56bar;
  wire in_55bar;
  wire in_54bar;
  wire in_53bar;
  wire in_52bar;
  wire in_51bar;
  wire in_50bar;
  wire in_49bar;
  wire in_48bar;
  wire in_47bar;
  wire in_46bar;
  wire in_45bar;
  wire in_44bar;
  wire in_43bar;
  wire in_42bar;
  wire in_41bar;
  wire in_40bar;
  wire in_39bar;
  wire in_38bar;
  wire in_37bar;
  wire in_36bar;
  wire in_35bar;
  wire in_34bar;
  wire in_33bar;
  wire in_32bar;
  wire in_31bar;
  wire in_30bar;
  wire in_29bar;
  wire in_28bar;
  wire in_27bar;
  wire in_26bar;
  wire in_25bar;
  wire in_24bar;
  wire in_23bar;
  wire in_22bar;
  wire in_21bar;
  wire in_20bar;
  wire in_19bar;
  wire in_18bar;
  wire in_17bar;
  wire in_16bar;
  wire in_15bar;
  wire in_14bar;
  wire in_13bar;
  wire in_12bar;
  wire in_11bar;
  wire in_10bar;
  wire in_9bar;
  wire in_8bar;
  wire in_7bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_3bar;
  wire in_2bar;
  wire in_1bar;
  wire in_0bar;
  wire n487bar;
  wire n488bar;
  wire n489bar;
  wire n490bar;
  wire n491bar;
  wire n492bar;
  wire n493bar;
  wire n494bar;
  wire n495bar;
  wire n496bar;
  wire n497bar;
  wire n498bar;
  wire n499bar;
  wire n500bar;
  wire n501bar;
  wire n502bar;
  wire n503bar;
  wire n504bar;
  wire n505bar;
  wire n506bar;
  wire n507bar;
  wire n508bar;
  wire n509bar;
  wire n510bar;
  wire n511bar;
  wire n512bar;
  wire n513bar;
  wire n514bar;
  wire n515bar;
  wire n516bar;
  wire n517bar;
  wire n518bar;
  wire n519bar;
  wire n520bar;
  wire n521bar;
  wire n522bar;
  wire n523bar;
  wire n524bar;
  wire n525bar;
  wire n526bar;
  wire n527bar;
  wire n528bar;
  wire n529bar;
  wire n530bar;
  wire n531bar;
  wire n532bar;
  wire n533bar;
  wire n534bar;
  wire n535bar;
  wire n536bar;
  wire n537bar;
  wire n538bar;
  wire n539bar;
  wire n540bar;
  wire n541bar;
  wire n542bar;
  wire n543bar;
  wire n544bar;
  wire n545bar;
  wire n546bar;
  wire n547bar;
  wire n548bar;
  wire n549bar;
  wire n550bar;
  wire n551bar;
  wire n552bar;
  wire n553bar;
  wire n554bar;
  wire n555bar;
  wire n556bar;
  wire n557bar;
  wire n558bar;
  wire n559bar;
  wire n560bar;
  wire n561bar;
  wire n562bar;
  wire n563bar;
  wire n564bar;
  wire n565bar;
  wire n566bar;
  wire n567bar;
  wire n568bar;
  wire n569bar;
  wire n570bar;
  wire n571bar;
  wire n572bar;
  wire n573bar;
  wire n574bar;
  wire n575bar;
  wire n576bar;
  wire n577bar;
  wire n578bar;
  wire n579bar;
  wire n580bar;
  wire n581bar;
  wire n582bar;
  wire n583bar;
  wire n584bar;
  wire n585bar;
  wire n586bar;
  wire n587bar;
  wire n588bar;
  wire n589bar;
  wire n590bar;
  wire n591bar;
  wire n592bar;
  wire n593bar;
  wire n594bar;
  wire n595bar;
  wire n596bar;
  wire n597bar;
  wire n598bar;
  wire n599bar;
  wire n600bar;
  wire n601bar;
  wire n602bar;
  wire n603bar;
  wire n604bar;
  wire n605bar;
  wire n606bar;
  wire n607bar;
  wire n608bar;
  wire n609bar;
  wire n610bar;
  wire n611bar;
  wire n612bar;
  wire n613bar;
  wire n614bar;
  wire n615bar;
  wire n616bar;
  wire n617bar;
  wire n618bar;
  wire n619bar;
  wire n620bar;
  wire n621bar;
  wire n622bar;
  wire n623bar;
  wire n624bar;
  wire n625bar;
  wire n626bar;
  wire n627bar;
  wire n628bar;
  wire n629bar;
  wire n630bar;
  wire n631bar;
  wire n632bar;
  wire n633bar;
  wire n634bar;
  wire n635bar;
  wire n636bar;
  wire n637bar;
  wire n638bar;
  wire n639bar;
  wire n640bar;
  wire n641bar;
  wire n642bar;
  wire n643bar;
  wire n644bar;
  wire n645bar;
  wire n646bar;
  wire n647bar;
  wire n648bar;
  wire n649bar;
  wire n650bar;
  wire n651bar;
  wire n652bar;
  wire n653bar;
  wire n654bar;
  wire n655bar;
  wire n656bar;
  wire n657bar;
  wire n658bar;
  wire n659bar;
  wire n660bar;
  wire n661bar;
  wire n662bar;
  wire n663bar;
  wire n664bar;
  wire n665bar;
  wire n666bar;
  wire n667bar;
  wire n668bar;
  wire n669bar;
  wire n670bar;
  wire n671bar;
  wire n672bar;
  wire n673bar;
  wire n674bar;
  wire n675bar;
  wire n676bar;
  wire n677bar;
  wire n678bar;
  wire n679bar;
  wire n680bar;
  wire n681bar;
  wire n682bar;
  wire n683bar;
  wire n684bar;
  wire n685bar;
  wire n686bar;
  wire n687bar;
  wire n688bar;
  wire n689bar;
  wire n690bar;
  wire n691bar;
  wire n692bar;
  wire n693bar;
  wire n694bar;
  wire n695bar;
  wire n696bar;
  wire n697bar;
  wire n698bar;
  wire n699bar;
  wire n700bar;
  wire n701bar;
  wire n702bar;
  wire n703bar;
  wire n704bar;
  wire n705bar;
  wire n706bar;
  wire n707bar;
  wire n708bar;
  wire n709bar;
  wire n710bar;
  wire n711bar;
  wire n712bar;
  wire n713bar;
  wire n714bar;
  wire n715bar;
  wire n716bar;
  wire n717bar;
  wire n718bar;
  wire n719bar;
  wire n720bar;
  wire n721bar;
  wire n722bar;
  wire n723bar;
  wire n724bar;
  wire n725bar;
  wire n726bar;
  wire n727bar;
  wire n728bar;
  wire n729bar;
  wire n730bar;
  wire n731bar;
  wire n732bar;
  wire n733bar;
  wire n734bar;
  wire n735bar;
  wire n736bar;
  wire n737bar;
  wire n738bar;
  wire n739bar;
  wire n740bar;
  wire n741bar;
  wire n742bar;
  wire n743bar;
  wire n744bar;
  wire n745bar;
  wire n746bar;
  wire n747bar;
  wire n748bar;
  wire n749bar;
  wire n750bar;
  wire n751bar;
  wire n752bar;
  wire n753bar;
  wire n754bar;
  wire n755bar;
  wire n756bar;
  wire n757bar;
  wire n758bar;
  wire n759bar;
  wire n760bar;
  wire n761bar;
  wire n762bar;
  wire n763bar;
  wire n764bar;
  wire n765bar;
  wire n766bar;
  wire n767bar;
  wire n768bar;
  wire n769bar;
  wire n770bar;
  wire n771bar;
  wire n772bar;
  wire n773bar;
  wire n774bar;
  wire n775bar;
  wire n776bar;
  wire n777bar;
  wire n778bar;
  wire n779bar;
  wire n780bar;
  wire n781bar;
  wire n782bar;
  wire n783bar;
  wire n784bar;
  wire n785bar;
  wire n786bar;
  wire n787bar;
  wire n788bar;
  wire n789bar;
  wire n790bar;
  wire n791bar;
  wire n792bar;
  wire n793bar;
  wire n794bar;
  wire n795bar;
  wire n796bar;
  wire n797bar;
  wire n798bar;
  wire n799bar;
  wire n800bar;
  wire n801bar;
  wire n802bar;
  wire n803bar;
  wire n804bar;
  wire n805bar;
  wire n806bar;
  wire n807bar;
  wire n808bar;
  wire n809bar;
  wire n810bar;
  wire n811bar;
  wire n812bar;
  wire n813bar;
  wire n814bar;
  wire n815bar;
  wire n816bar;
  wire n817bar;
  wire n818bar;
  wire n819bar;
  wire n820bar;
  wire n821bar;
  wire n822bar;
  wire n823bar;
  wire n824bar;
  wire n825bar;
  wire n826bar;
  wire n827bar;
  wire n828bar;
  wire n829bar;
  wire n830bar;
  wire n831bar;
  wire n832bar;
  wire n833bar;
  wire n834bar;
  wire n835bar;
  wire n836bar;
  wire n837bar;
  wire n838bar;
  wire n839bar;
  wire n840bar;
  wire n841bar;
  wire n842bar;
  wire n843bar;
  wire n844bar;
  wire n845bar;
  wire n846bar;
  wire n847bar;
  wire n848bar;
  wire n849bar;
  wire n850bar;
  wire n851bar;
  wire n852bar;
  wire n853bar;
  wire n854bar;
  wire n855bar;
  wire n856bar;
  wire n857bar;
  wire n858bar;
  wire n859bar;
  wire n860bar;
  wire n861bar;
  wire n862bar;
  wire n863bar;
  wire n864bar;
  wire n865bar;
  wire n866bar;
  wire n867bar;
  wire n868bar;
  wire n869bar;
  wire n870bar;
  wire n871bar;
  wire n872bar;
  wire n873bar;
  wire n874bar;
  wire n875bar;
  wire n876bar;
  wire n877bar;
  wire n878bar;
  wire n879bar;
  wire n880bar;
  wire n881bar;
  wire n882bar;
  wire n883bar;
  wire n884bar;
  wire n885bar;
  wire n886bar;
  wire n887bar;
  wire n888bar;
  wire n889bar;
  wire n890bar;
  wire n891bar;
  wire n892bar;
  wire n893bar;
  wire n894bar;
  wire n895bar;
  wire n896bar;
  wire n897bar;
  wire n898bar;
  wire n899bar;
  wire n900bar;
  wire n901bar;
  wire n902bar;
  wire n903bar;
  wire n904bar;
  wire n905bar;
  wire n906bar;
  wire n907bar;
  wire n908bar;
  wire n909bar;
  wire n910bar;
  wire n911bar;
  wire n912bar;
  wire n913bar;
  wire n914bar;
  wire n915bar;
  wire n916bar;
  wire n917bar;
  wire n918bar;
  wire n919bar;
  wire n920bar;
  wire n921bar;
  wire n922bar;
  wire n923bar;
  wire n924bar;
  wire n925bar;
  wire n926bar;
  wire n927bar;
  wire n928bar;
  wire n929bar;
  wire n930bar;
  wire n931bar;
  wire n932bar;
  wire n933bar;
  wire n934bar;
  wire n935bar;
  wire n936bar;
  wire n937bar;
  wire n938bar;
  wire n939bar;
  wire n940bar;
  wire n941bar;
  wire n942bar;
  wire n943bar;
  wire n944bar;
  wire n945bar;
  wire n946bar;
  wire n947bar;
  wire n948bar;
  wire n949bar;
  wire n950bar;
  wire n951bar;
  wire n952bar;
  wire n953bar;
  wire n954bar;
  wire n955bar;
  wire n956bar;
  wire n957bar;
  wire n958bar;
  wire n959bar;
  wire n960bar;
  wire n961bar;
  wire n962bar;
  wire n963bar;
  wire n964bar;
  wire n965bar;
  wire n966bar;
  wire n967bar;
  wire n968bar;
  wire n969bar;
  wire n970bar;
  wire n971bar;
  wire n972bar;
//wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];
  //OR U1
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1 (
    .O(out[7]),
    .I0(n972),
    .I1(n971)
  );
  //AND U1bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1bar (
    .O(outbar[7]),
    .I0(n972bar),
    .I1(n971bar)
  );
  //OR U2
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2 (
    .O(n971),
    .I0(n970),
    .I1(n969)
  );
  //AND U2bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2bar (
    .O(n971bar),
    .I0(n970bar),
    .I1(n969bar)
  );
  //OR U3
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3 (
    .O(n969),
    .I0(n968),
    .I1(n967)
  );
  //AND U3bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3bar (
    .O(n969bar),
    .I0(n968bar),
    .I1(n967bar)
  );
  //OR U4
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4 (
    .O(n967),
    .I0(n966),
    .I1(n965)
  );
  //AND U4bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4bar (
    .O(n967bar),
    .I0(n966bar),
    .I1(n965bar)
  );
  //OR U5
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5 (
    .O(n968),
    .I0(n964),
    .I1(n963)
  );
  //AND U5bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5bar (
    .O(n968bar),
    .I0(n964bar),
    .I1(n963bar)
  );
  //OR U6
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6 (
    .O(n963),
    .I0(in[116]),
    .I1(n962)
  );
  //AND U6bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6bar (
    .O(n963bar),
    .I0(inbar[116]),
    .I1(n962bar)
  );
  //OR U7
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7 (
    .O(n970),
    .I0(n961),
    .I1(n960)
  );
  //AND U7bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7bar (
    .O(n970bar),
    .I0(n961bar),
    .I1(n960bar)
  );
  //OR U8
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8 (
    .O(n960),
    .I0(in[150]),
    .I1(in[127])
  );
  //AND U8bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8bar (
    .O(n960bar),
    .I0(inbar[150]),
    .I1(inbar[127])
  );
  //OR U9
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9 (
    .O(n961),
    .I0(in[160]),
    .I1(n959)
  );
  //AND U9bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9bar (
    .O(n961bar),
    .I0(inbar[160]),
    .I1(n959bar)
  );
  //OR U10
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10 (
    .O(n959),
    .I0(in[252]),
    .I1(in[168])
  );
  //AND U10bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10bar (
    .O(n959bar),
    .I0(inbar[252]),
    .I1(inbar[168])
  );
  //OR U11
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11 (
    .O(n972),
    .I0(n958),
    .I1(n957)
  );
  //AND U11bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11bar (
    .O(n972bar),
    .I0(n958bar),
    .I1(n957bar)
  );
  //OR U12
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12 (
    .O(n957),
    .I0(n956),
    .I1(n955)
  );
  //AND U12bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12bar (
    .O(n957bar),
    .I0(n956bar),
    .I1(n955bar)
  );
  //OR U13
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13 (
    .O(n955),
    .I0(in_17),
    .I1(in[96])
  );
  //AND U13bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13bar (
    .O(n955bar),
    .I0(in_17bar),
    .I1(inbar[96])
  );
  //OR U14
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14 (
    .O(n956),
    .I0(in_23),
    .I1(n954)
  );
  //AND U14bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14bar (
    .O(n956bar),
    .I0(in_23bar),
    .I1(n954bar)
  );
  //OR U15
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15 (
    .O(n954),
    .I0(in_31),
    .I1(in_26)
  );
  //AND U15bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15bar (
    .O(n954bar),
    .I0(in_31bar),
    .I1(in_26bar)
  );
  //OR U16
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16 (
    .O(n958),
    .I0(n953),
    .I1(n952)
  );
  //AND U16bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16bar (
    .O(n958bar),
    .I0(n953bar),
    .I1(n952bar)
  );
  //OR U17
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U17 (
    .O(n952),
    .I0(in_58),
    .I1(in_4)
  );
  //AND U17bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U17bar (
    .O(n952bar),
    .I0(in_58bar),
    .I1(in_4bar)
  );
  //OR U18
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U18 (
    .O(n953),
    .I0(in_59),
    .I1(n951)
  );
  //AND U18bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U18bar (
    .O(n953bar),
    .I0(in_59bar),
    .I1(n951bar)
  );
  //OR U19
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U19 (
    .O(n951),
    .I0(in_71),
    .I1(in_62)
  );
  //AND U19bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U19bar (
    .O(n951bar),
    .I0(in_71bar),
    .I1(in_62bar)
  );
  //OR U20
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U20 (
    .O(out[6]),
    .I0(n950),
    .I1(n949)
  );
  //AND U20bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U20bar (
    .O(outbar[6]),
    .I0(n950bar),
    .I1(n949bar)
  );
  //OR U21
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U21 (
    .O(n949),
    .I0(n948),
    .I1(n947)
  );
  //AND U21bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U21bar (
    .O(n949bar),
    .I0(n948bar),
    .I1(n947bar)
  );
  //OR U22
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U22 (
    .O(n947),
    .I0(n946),
    .I1(n945)
  );
  //AND U22bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U22bar (
    .O(n947bar),
    .I0(n946bar),
    .I1(n945bar)
  );
  //OR U23
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U23 (
    .O(n945),
    .I0(n944),
    .I1(n943)
  );
  //AND U23bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U23bar (
    .O(n945bar),
    .I0(n944bar),
    .I1(n943bar)
  );
  //OR U24
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U24 (
    .O(n946),
    .I0(n942),
    .I1(n941)
  );
  //AND U24bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U24bar (
    .O(n946bar),
    .I0(n942bar),
    .I1(n941bar)
  );
  //OR U25
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U25 (
    .O(n941),
    .I0(in[101]),
    .I1(n940)
  );
  //AND U25bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U25bar (
    .O(n941bar),
    .I0(inbar[101]),
    .I1(n940bar)
  );
  //OR U26
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U26 (
    .O(n948),
    .I0(n939),
    .I1(n938)
  );
  //AND U26bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U26bar (
    .O(n948bar),
    .I0(n939bar),
    .I1(n938bar)
  );
  //OR U27
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U27 (
    .O(n938),
    .I0(in[114]),
    .I1(in[104])
  );
  //AND U27bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U27bar (
    .O(n938bar),
    .I0(inbar[114]),
    .I1(inbar[104])
  );
  //OR U28
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U28 (
    .O(n939),
    .I0(in[128]),
    .I1(n937)
  );
  //AND U28bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U28bar (
    .O(n939bar),
    .I0(inbar[128]),
    .I1(n937bar)
  );
  //OR U29
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U29 (
    .O(n937),
    .I0(in[136]),
    .I1(in[134])
  );
  //AND U29bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U29bar (
    .O(n937bar),
    .I0(inbar[136]),
    .I1(inbar[134])
  );
  //OR U30
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U30 (
    .O(n950),
    .I0(n936),
    .I1(n935)
  );
  //AND U30bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U30bar (
    .O(n950bar),
    .I0(n936bar),
    .I1(n935bar)
  );
  //OR U31
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U31 (
    .O(n935),
    .I0(n934),
    .I1(n933)
  );
  //AND U31bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U31bar (
    .O(n935bar),
    .I0(n934bar),
    .I1(n933bar)
  );
  //OR U32
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U32 (
    .O(n933),
    .I0(in[177]),
    .I1(in[164])
  );
  //AND U32bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U32bar (
    .O(n933bar),
    .I0(inbar[177]),
    .I1(inbar[164])
  );
  //OR U33
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U33 (
    .O(n934),
    .I0(in[212]),
    .I1(n932)
  );
  //AND U33bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U33bar (
    .O(n934bar),
    .I0(inbar[212]),
    .I1(n932bar)
  );
  //OR U34
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U34 (
    .O(n932),
    .I0(in[248]),
    .I1(in[221])
  );
  //AND U34bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U34bar (
    .O(n932bar),
    .I0(inbar[248]),
    .I1(inbar[221])
  );
  //OR U35
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U35 (
    .O(n936),
    .I0(n931),
    .I1(n930)
  );
  //AND U35bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U35bar (
    .O(n936bar),
    .I0(n931bar),
    .I1(n930bar)
  );
  //OR U36
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U36 (
    .O(n930),
    .I0(in_18),
    .I1(in[93])
  );
  //AND U36bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U36bar (
    .O(n930bar),
    .I0(in_18bar),
    .I1(inbar[93])
  );
  //OR U37
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U37 (
    .O(n931),
    .I0(in_31),
    .I1(n929)
  );
  //AND U37bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U37bar (
    .O(n931bar),
    .I0(in_31bar),
    .I1(n929bar)
  );
  //OR U38
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U38 (
    .O(n929),
    .I0(in_7),
    .I1(in_39)
  );
  //AND U38bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U38bar (
    .O(n929bar),
    .I0(in_7bar),
    .I1(in_39bar)
  );
  //OR U39
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U39 (
    .O(out[5]),
    .I0(n928),
    .I1(n927)
  );
  //AND U39bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U39bar (
    .O(outbar[5]),
    .I0(n928bar),
    .I1(n927bar)
  );
  //OR U40
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U40 (
    .O(n927),
    .I0(n926),
    .I1(n925)
  );
  //AND U40bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U40bar (
    .O(n927bar),
    .I0(n926bar),
    .I1(n925bar)
  );
  //OR U41
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U41 (
    .O(n925),
    .I0(n924),
    .I1(n923)
  );
  //AND U41bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U41bar (
    .O(n925bar),
    .I0(n924bar),
    .I1(n923bar)
  );
  //OR U42
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U42 (
    .O(n923),
    .I0(n922),
    .I1(n921)
  );
  //AND U42bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U42bar (
    .O(n923bar),
    .I0(n922bar),
    .I1(n921bar)
  );
  //OR U43
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U43 (
    .O(n924),
    .I0(n940),
    .I1(n920)
  );
  //AND U43bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U43bar (
    .O(n924bar),
    .I0(n940bar),
    .I1(n920bar)
  );
  //OR U44
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U44 (
    .O(n920),
    .I0(in[111]),
    .I1(n919)
  );
  //AND U44bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U44bar (
    .O(n920bar),
    .I0(inbar[111]),
    .I1(n919bar)
  );
  //OR U45
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U45 (
    .O(n940),
    .I0(n918),
    .I1(n917)
  );
  //AND U45bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U45bar (
    .O(n940bar),
    .I0(n918bar),
    .I1(n917bar)
  );
  //OR U46
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U46 (
    .O(n917),
    .I0(n916),
    .I1(n915)
  );
  //AND U46bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U46bar (
    .O(n917bar),
    .I0(n916bar),
    .I1(n915bar)
  );
  //OR U47
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U47 (
    .O(n915),
    .I0(n914),
    .I1(n913)
  );
  //AND U47bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U47bar (
    .O(n915bar),
    .I0(n914bar),
    .I1(n913bar)
  );
  //OR U48
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U48 (
    .O(n913),
    .I0(in[140]),
    .I1(in[131])
  );
  //AND U48bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U48bar (
    .O(n913bar),
    .I0(inbar[140]),
    .I1(inbar[131])
  );
  //OR U49
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U49 (
    .O(n914),
    .I0(in[160]),
    .I1(in[144])
  );
  //AND U49bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U49bar (
    .O(n914bar),
    .I0(inbar[160]),
    .I1(inbar[144])
  );
  //OR U50
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U50 (
    .O(n916),
    .I0(n912),
    .I1(n911)
  );
  //AND U50bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U50bar (
    .O(n916bar),
    .I0(n912bar),
    .I1(n911bar)
  );
  //OR U51
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U51 (
    .O(n911),
    .I0(in[179]),
    .I1(in[174])
  );
  //AND U51bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U51bar (
    .O(n911bar),
    .I0(inbar[179]),
    .I1(inbar[174])
  );
  //OR U52
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U52 (
    .O(n912),
    .I0(in[188]),
    .I1(in[184])
  );
  //AND U52bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U52bar (
    .O(n912bar),
    .I0(inbar[188]),
    .I1(inbar[184])
  );
  //OR U53
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U53 (
    .O(n918),
    .I0(n910),
    .I1(n909)
  );
  //AND U53bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U53bar (
    .O(n918bar),
    .I0(n910bar),
    .I1(n909bar)
  );
  //OR U54
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U54 (
    .O(n909),
    .I0(n908),
    .I1(n907)
  );
  //AND U54bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U54bar (
    .O(n909bar),
    .I0(n908bar),
    .I1(n907bar)
  );
  //OR U55
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U55 (
    .O(n907),
    .I0(in[216]),
    .I1(in[200])
  );
  //AND U55bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U55bar (
    .O(n907bar),
    .I0(inbar[216]),
    .I1(inbar[200])
  );
  //OR U56
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U56 (
    .O(n908),
    .I0(in[228]),
    .I1(in[224])
  );
  //AND U56bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U56bar (
    .O(n908bar),
    .I0(inbar[228]),
    .I1(inbar[224])
  );
  //OR U57
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U57 (
    .O(n910),
    .I0(n906),
    .I1(n905)
  );
  //AND U57bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U57bar (
    .O(n910bar),
    .I0(n906bar),
    .I1(n905bar)
  );
  //OR U58
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U58 (
    .O(n905),
    .I0(in[247]),
    .I1(in[235])
  );
  //AND U58bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U58bar (
    .O(n905bar),
    .I0(inbar[247]),
    .I1(inbar[235])
  );
  //OR U59
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U59 (
    .O(n906),
    .I0(in_42),
    .I1(in[83])
  );
  //AND U59bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U59bar (
    .O(n906bar),
    .I0(in_42bar),
    .I1(inbar[83])
  );
  //OR U60
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U60 (
    .O(n926),
    .I0(n904),
    .I1(n903)
  );
  //AND U60bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U60bar (
    .O(n926bar),
    .I0(n904bar),
    .I1(n903bar)
  );
  //OR U61
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U61 (
    .O(n903),
    .I0(in[166]),
    .I1(in[123])
  );
  //AND U61bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U61bar (
    .O(n903bar),
    .I0(inbar[166]),
    .I1(inbar[123])
  );
  //OR U62
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U62 (
    .O(n904),
    .I0(in[170]),
    .I1(n902)
  );
  //AND U62bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U62bar (
    .O(n904bar),
    .I0(inbar[170]),
    .I1(n902bar)
  );
  //OR U63
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U63 (
    .O(n902),
    .I0(in[194]),
    .I1(in[183])
  );
  //AND U63bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U63bar (
    .O(n902bar),
    .I0(inbar[194]),
    .I1(inbar[183])
  );
  //OR U64
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U64 (
    .O(n928),
    .I0(n901),
    .I1(n900)
  );
  //AND U64bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U64bar (
    .O(n928bar),
    .I0(n901bar),
    .I1(n900bar)
  );
  //OR U65
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U65 (
    .O(n900),
    .I0(n899),
    .I1(n898)
  );
  //AND U65bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U65bar (
    .O(n900bar),
    .I0(n899bar),
    .I1(n898bar)
  );
  //OR U66
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U66 (
    .O(n898),
    .I0(in[241]),
    .I1(in[238])
  );
  //AND U66bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U66bar (
    .O(n898bar),
    .I0(inbar[241]),
    .I1(inbar[238])
  );
  //OR U67
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U67 (
    .O(n899),
    .I0(in[250]),
    .I1(n897)
  );
  //AND U67bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U67bar (
    .O(n899bar),
    .I0(inbar[250]),
    .I1(n897bar)
  );
  //OR U68
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U68 (
    .O(n897),
    .I0(in_24),
    .I1(in[84])
  );
  //AND U68bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U68bar (
    .O(n897bar),
    .I0(in_24bar),
    .I1(inbar[84])
  );
  //OR U69
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U69 (
    .O(n901),
    .I0(n896),
    .I1(n895)
  );
  //AND U69bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U69bar (
    .O(n901bar),
    .I0(n896bar),
    .I1(n895bar)
  );
  //OR U70
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U70 (
    .O(n895),
    .I0(in_41),
    .I1(in_29)
  );
  //AND U70bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U70bar (
    .O(n895bar),
    .I0(in_41bar),
    .I1(in_29bar)
  );
  //OR U71
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U71 (
    .O(n896),
    .I0(in_66),
    .I1(n894)
  );
  //AND U71bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U71bar (
    .O(n896bar),
    .I0(in_66bar),
    .I1(n894bar)
  );
  //OR U72
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U72 (
    .O(n894),
    .I0(in_76),
    .I1(in_71)
  );
  //AND U72bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U72bar (
    .O(n894bar),
    .I0(in_76bar),
    .I1(in_71bar)
  );
  //OR U73
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U73 (
    .O(out[4]),
    .I0(n893),
    .I1(n892)
  );
  //AND U73bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U73bar (
    .O(outbar[4]),
    .I0(n893bar),
    .I1(n892bar)
  );
  //OR U74
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U74 (
    .O(n892),
    .I0(n891),
    .I1(n890)
  );
  //AND U74bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U74bar (
    .O(n892bar),
    .I0(n891bar),
    .I1(n890bar)
  );
  //OR U75
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U75 (
    .O(n890),
    .I0(n889),
    .I1(n888)
  );
  //AND U75bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U75bar (
    .O(n890bar),
    .I0(n889bar),
    .I1(n888bar)
  );
  //OR U76
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U76 (
    .O(n888),
    .I0(n922),
    .I1(n887)
  );
  //AND U76bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U76bar (
    .O(n888bar),
    .I0(n922bar),
    .I1(n887bar)
  );
  //OR U77
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U77 (
    .O(n922),
    .I0(n886),
    .I1(n885)
  );
  //AND U77bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U77bar (
    .O(n922bar),
    .I0(n886bar),
    .I1(n885bar)
  );
  //OR U78
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U78 (
    .O(n885),
    .I0(n884),
    .I1(n883)
  );
  //AND U78bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U78bar (
    .O(n885bar),
    .I0(n884bar),
    .I1(n883bar)
  );
  //OR U79
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U79 (
    .O(n883),
    .I0(n882),
    .I1(n881)
  );
  //AND U79bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U79bar (
    .O(n883bar),
    .I0(n882bar),
    .I1(n881bar)
  );
  //OR U80
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U80 (
    .O(n881),
    .I0(in[118]),
    .I1(in[109])
  );
  //AND U80bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U80bar (
    .O(n881bar),
    .I0(inbar[118]),
    .I1(inbar[109])
  );
  //OR U81
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U81 (
    .O(n882),
    .I0(in[139]),
    .I1(in[120])
  );
  //AND U81bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U81bar (
    .O(n882bar),
    .I0(inbar[139]),
    .I1(inbar[120])
  );
  //OR U82
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U82 (
    .O(n884),
    .I0(n880),
    .I1(n879)
  );
  //AND U82bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U82bar (
    .O(n884bar),
    .I0(n880bar),
    .I1(n879bar)
  );
  //OR U83
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U83 (
    .O(n879),
    .I0(in[198]),
    .I1(in[154])
  );
  //AND U83bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U83bar (
    .O(n879bar),
    .I0(inbar[198]),
    .I1(inbar[154])
  );
  //OR U84
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U84 (
    .O(n880),
    .I0(in[210]),
    .I1(in[205])
  );
  //AND U84bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U84bar (
    .O(n880bar),
    .I0(inbar[210]),
    .I1(inbar[205])
  );
  //OR U85
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U85 (
    .O(n886),
    .I0(n878),
    .I1(n877)
  );
  //AND U85bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U85bar (
    .O(n886bar),
    .I0(n878bar),
    .I1(n877bar)
  );
  //OR U86
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U86 (
    .O(n877),
    .I0(n876),
    .I1(n875)
  );
  //AND U86bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U86bar (
    .O(n877bar),
    .I0(n876bar),
    .I1(n875bar)
  );
  //OR U87
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U87 (
    .O(n875),
    .I0(in[219]),
    .I1(in[217])
  );
  //AND U87bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U87bar (
    .O(n875bar),
    .I0(inbar[219]),
    .I1(inbar[217])
  );
  //OR U88
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U88 (
    .O(n876),
    .I0(in[86]),
    .I1(in[252])
  );
  //AND U88bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U88bar (
    .O(n876bar),
    .I0(inbar[86]),
    .I1(inbar[252])
  );
  //OR U89
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U89 (
    .O(n878),
    .I0(n874),
    .I1(n873)
  );
  //AND U89bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U89bar (
    .O(n878bar),
    .I0(n874bar),
    .I1(n873bar)
  );
  //OR U90
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U90 (
    .O(n873),
    .I0(in_40),
    .I1(in[91])
  );
  //AND U90bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U90bar (
    .O(n873bar),
    .I0(in_40bar),
    .I1(inbar[91])
  );
  //OR U91
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U91 (
    .O(n874),
    .I0(in_8),
    .I1(in_46)
  );
  //AND U91bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U91bar (
    .O(n874bar),
    .I0(in_8bar),
    .I1(in_46bar)
  );
  //OR U92
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U92 (
    .O(n889),
    .I0(n872),
    .I1(n871)
  );
  //AND U92bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U92bar (
    .O(n889bar),
    .I0(n872bar),
    .I1(n871bar)
  );
  //OR U93
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U93 (
    .O(n871),
    .I0(in[117]),
    .I1(n943)
  );
  //AND U93bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U93bar (
    .O(n871bar),
    .I0(inbar[117]),
    .I1(n943bar)
  );
  //OR U94
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U94 (
    .O(n943),
    .I0(n870),
    .I1(n869)
  );
  //AND U94bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U94bar (
    .O(n943bar),
    .I0(n870bar),
    .I1(n869bar)
  );
  //OR U95
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U95 (
    .O(n869),
    .I0(n868),
    .I1(n867)
  );
  //AND U95bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U95bar (
    .O(n869bar),
    .I0(n868bar),
    .I1(n867bar)
  );
  //OR U96
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U96 (
    .O(n867),
    .I0(n866),
    .I1(n865)
  );
  //AND U96bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U96bar (
    .O(n867bar),
    .I0(n866bar),
    .I1(n865bar)
  );
  //OR U97
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U97 (
    .O(n865),
    .I0(n864),
    .I1(n863)
  );
  //AND U97bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U97bar (
    .O(n865bar),
    .I0(n864bar),
    .I1(n863bar)
  );
  //OR U98
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U98 (
    .O(n866),
    .I0(in[108]),
    .I1(n919)
  );
  //AND U98bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U98bar (
    .O(n866bar),
    .I0(inbar[108]),
    .I1(n919bar)
  );
  //OR U99
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U99 (
    .O(n919),
    .I0(n862),
    .I1(n861)
  );
  //AND U99bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U99bar (
    .O(n919bar),
    .I0(n862bar),
    .I1(n861bar)
  );
  //OR U100
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U100 (
    .O(n861),
    .I0(n860),
    .I1(n859)
  );
  //AND U100bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U100bar (
    .O(n861bar),
    .I0(n860bar),
    .I1(n859bar)
  );
  //OR U101
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U101 (
    .O(n859),
    .I0(n858),
    .I1(n857)
  );
  //AND U101bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U101bar (
    .O(n859bar),
    .I0(n858bar),
    .I1(n857bar)
  );
  //OR U102
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U102 (
    .O(n857),
    .I0(in[119]),
    .I1(in[105])
  );
  //AND U102bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U102bar (
    .O(n857bar),
    .I0(inbar[119]),
    .I1(inbar[105])
  );
  //OR U103
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U103 (
    .O(n858),
    .I0(in[186]),
    .I1(in[175])
  );
  //AND U103bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U103bar (
    .O(n858bar),
    .I0(inbar[186]),
    .I1(inbar[175])
  );
  //OR U104
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U104 (
    .O(n860),
    .I0(n856),
    .I1(n855)
  );
  //AND U104bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U104bar (
    .O(n860bar),
    .I0(n856bar),
    .I1(n855bar)
  );
  //OR U105
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U105 (
    .O(n855),
    .I0(in[202]),
    .I1(in[193])
  );
  //AND U105bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U105bar (
    .O(n855bar),
    .I0(inbar[202]),
    .I1(inbar[193])
  );
  //OR U106
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U106 (
    .O(n856),
    .I0(in[225]),
    .I1(in[208])
  );
  //AND U106bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U106bar (
    .O(n856bar),
    .I0(inbar[225]),
    .I1(inbar[208])
  );
  //OR U107
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U107 (
    .O(n862),
    .I0(n854),
    .I1(n853)
  );
  //AND U107bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U107bar (
    .O(n862bar),
    .I0(n854bar),
    .I1(n853bar)
  );
  //OR U108
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U108 (
    .O(n853),
    .I0(n852),
    .I1(n851)
  );
  //AND U108bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U108bar (
    .O(n853bar),
    .I0(n852bar),
    .I1(n851bar)
  );
  //OR U109
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U109 (
    .O(n851),
    .I0(in_1),
    .I1(in[85])
  );
  //AND U109bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U109bar (
    .O(n851bar),
    .I0(in_1bar),
    .I1(inbar[85])
  );
  //OR U110
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U110 (
    .O(n852),
    .I0(in_23),
    .I1(in_19)
  );
  //AND U110bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U110bar (
    .O(n852bar),
    .I0(in_23bar),
    .I1(in_19bar)
  );
  //OR U111
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U111 (
    .O(n854),
    .I0(n850),
    .I1(n849)
  );
  //AND U111bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U111bar (
    .O(n854bar),
    .I0(n850bar),
    .I1(n849bar)
  );
  //OR U112
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U112 (
    .O(n849),
    .I0(in_43),
    .I1(in_33)
  );
  //AND U112bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U112bar (
    .O(n849bar),
    .I0(in_43bar),
    .I1(in_33bar)
  );
  //OR U113
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U113 (
    .O(n850),
    .I0(in_63),
    .I1(in_44)
  );
  //AND U113bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U113bar (
    .O(n850bar),
    .I0(in_63bar),
    .I1(in_44bar)
  );
  //OR U114
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U114 (
    .O(n868),
    .I0(n848),
    .I1(n847)
  );
  //AND U114bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U114bar (
    .O(n868bar),
    .I0(n848bar),
    .I1(n847bar)
  );
  //OR U115
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U115 (
    .O(n847),
    .I0(in[141]),
    .I1(in[112])
  );
  //AND U115bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U115bar (
    .O(n847bar),
    .I0(inbar[141]),
    .I1(inbar[112])
  );
  //OR U116
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U116 (
    .O(n848),
    .I0(in[147]),
    .I1(n846)
  );
  //AND U116bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U116bar (
    .O(n848bar),
    .I0(inbar[147]),
    .I1(n846bar)
  );
  //OR U117
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U117 (
    .O(n846),
    .I0(in[181]),
    .I1(in[167])
  );
  //AND U117bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U117bar (
    .O(n846bar),
    .I0(inbar[181]),
    .I1(inbar[167])
  );
  //OR U118
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U118 (
    .O(n870),
    .I0(n845),
    .I1(n844)
  );
  //AND U118bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U118bar (
    .O(n870bar),
    .I0(n845bar),
    .I1(n844bar)
  );
  //OR U119
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U119 (
    .O(n844),
    .I0(n843),
    .I1(n842)
  );
  //AND U119bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U119bar (
    .O(n844bar),
    .I0(n843bar),
    .I1(n842bar)
  );
  //OR U120
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U120 (
    .O(n842),
    .I0(in[229]),
    .I1(in[201])
  );
  //AND U120bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U120bar (
    .O(n842bar),
    .I0(inbar[229]),
    .I1(inbar[201])
  );
  //OR U121
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U121 (
    .O(n843),
    .I0(in[237]),
    .I1(n841)
  );
  //AND U121bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U121bar (
    .O(n843bar),
    .I0(inbar[237]),
    .I1(n841bar)
  );
  //OR U122
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U122 (
    .O(n841),
    .I0(in[94]),
    .I1(in[253])
  );
  //AND U122bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U122bar (
    .O(n841bar),
    .I0(inbar[94]),
    .I1(inbar[253])
  );
  //OR U123
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U123 (
    .O(n845),
    .I0(n840),
    .I1(n839)
  );
  //AND U123bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U123bar (
    .O(n845bar),
    .I0(n840bar),
    .I1(n839bar)
  );
  //OR U124
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U124 (
    .O(n839),
    .I0(in_21),
    .I1(in[96])
  );
  //AND U124bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U124bar (
    .O(n839bar),
    .I0(in_21bar),
    .I1(inbar[96])
  );
  //OR U125
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U125 (
    .O(n840),
    .I0(in_25),
    .I1(n838)
  );
  //AND U125bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U125bar (
    .O(n840bar),
    .I0(in_25bar),
    .I1(n838bar)
  );
  //OR U126
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U126 (
    .O(n838),
    .I0(in_81),
    .I1(in_45)
  );
  //AND U126bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U126bar (
    .O(n838bar),
    .I0(in_81bar),
    .I1(in_45bar)
  );
  //OR U127
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U127 (
    .O(n891),
    .I0(n837),
    .I1(n836)
  );
  //AND U127bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U127bar (
    .O(n891bar),
    .I0(n837bar),
    .I1(n836bar)
  );
  //OR U128
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U128 (
    .O(n836),
    .I0(in[142]),
    .I1(in[124])
  );
  //AND U128bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U128bar (
    .O(n836bar),
    .I0(inbar[142]),
    .I1(inbar[124])
  );
  //OR U129
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U129 (
    .O(n837),
    .I0(in[150]),
    .I1(n835)
  );
  //AND U129bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U129bar (
    .O(n837bar),
    .I0(inbar[150]),
    .I1(n835bar)
  );
  //OR U130
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U130 (
    .O(n835),
    .I0(in[172]),
    .I1(in[155])
  );
  //AND U130bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U130bar (
    .O(n835bar),
    .I0(inbar[172]),
    .I1(inbar[155])
  );
  //OR U131
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U131 (
    .O(n893),
    .I0(n834),
    .I1(n833)
  );
  //AND U131bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U131bar (
    .O(n893bar),
    .I0(n834bar),
    .I1(n833bar)
  );
  //OR U132
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U132 (
    .O(n833),
    .I0(n832),
    .I1(n831)
  );
  //AND U132bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U132bar (
    .O(n833bar),
    .I0(n832bar),
    .I1(n831bar)
  );
  //OR U133
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U133 (
    .O(n831),
    .I0(in[196]),
    .I1(in[173])
  );
  //AND U133bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U133bar (
    .O(n831bar),
    .I0(inbar[196]),
    .I1(inbar[173])
  );
  //OR U134
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U134 (
    .O(n832),
    .I0(in[222]),
    .I1(n830)
  );
  //AND U134bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U134bar (
    .O(n832bar),
    .I0(inbar[222]),
    .I1(n830bar)
  );
  //OR U135
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U135 (
    .O(n830),
    .I0(in[227]),
    .I1(in[226])
  );
  //AND U135bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U135bar (
    .O(n830bar),
    .I0(inbar[227]),
    .I1(inbar[226])
  );
  //OR U136
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U136 (
    .O(n834),
    .I0(n829),
    .I1(n828)
  );
  //AND U136bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U136bar (
    .O(n834bar),
    .I0(n829bar),
    .I1(n828bar)
  );
  //OR U137
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U137 (
    .O(n828),
    .I0(in[249]),
    .I1(in[231])
  );
  //AND U137bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U137bar (
    .O(n828bar),
    .I0(inbar[249]),
    .I1(inbar[231])
  );
  //OR U138
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U138 (
    .O(n829),
    .I0(in_28),
    .I1(n827)
  );
  //AND U138bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U138bar (
    .O(n829bar),
    .I0(in_28bar),
    .I1(n827bar)
  );
  //OR U139
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U139 (
    .O(n827),
    .I0(in_52),
    .I1(in_47)
  );
  //AND U139bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U139bar (
    .O(n827bar),
    .I0(in_52bar),
    .I1(in_47bar)
  );
  //OR U140
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U140 (
    .O(out[3]),
    .I0(n826),
    .I1(n825)
  );
  //AND U140bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U140bar (
    .O(outbar[3]),
    .I0(n826bar),
    .I1(n825bar)
  );
  //OR U141
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U141 (
    .O(n825),
    .I0(n824),
    .I1(n823)
  );
  //AND U141bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U141bar (
    .O(n825bar),
    .I0(n824bar),
    .I1(n823bar)
  );
  //OR U142
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U142 (
    .O(n823),
    .I0(n822),
    .I1(n821)
  );
  //AND U142bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U142bar (
    .O(n823bar),
    .I0(n822bar),
    .I1(n821bar)
  );
  //OR U143
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U143 (
    .O(n821),
    .I0(n820),
    .I1(n819)
  );
  //AND U143bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U143bar (
    .O(n821bar),
    .I0(n820bar),
    .I1(n819bar)
  );
  //OR U144
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U144 (
    .O(n822),
    .I0(n964),
    .I1(n818)
  );
  //AND U144bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U144bar (
    .O(n822bar),
    .I0(n964bar),
    .I1(n818bar)
  );
  //OR U145
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U145 (
    .O(n818),
    .I0(in[118]),
    .I1(n817)
  );
  //AND U145bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U145bar (
    .O(n818bar),
    .I0(inbar[118]),
    .I1(n817bar)
  );
  //OR U146
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U146 (
    .O(n964),
    .I0(n816),
    .I1(n815)
  );
  //AND U146bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U146bar (
    .O(n964bar),
    .I0(n816bar),
    .I1(n815bar)
  );
  //OR U147
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U147 (
    .O(n815),
    .I0(n814),
    .I1(n813)
  );
  //AND U147bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U147bar (
    .O(n815bar),
    .I0(n814bar),
    .I1(n813bar)
  );
  //OR U148
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U148 (
    .O(n813),
    .I0(n812),
    .I1(n811)
  );
  //AND U148bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U148bar (
    .O(n813bar),
    .I0(n812bar),
    .I1(n811bar)
  );
  //OR U149
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U149 (
    .O(n811),
    .I0(in[122]),
    .I1(in[111])
  );
  //AND U149bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U149bar (
    .O(n811bar),
    .I0(inbar[122]),
    .I1(inbar[111])
  );
  //OR U150
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U150 (
    .O(n812),
    .I0(in[154]),
    .I1(in[151])
  );
  //AND U150bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U150bar (
    .O(n812bar),
    .I0(inbar[154]),
    .I1(inbar[151])
  );
  //OR U151
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U151 (
    .O(n814),
    .I0(n810),
    .I1(n809)
  );
  //AND U151bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U151bar (
    .O(n814bar),
    .I0(n810bar),
    .I1(n809bar)
  );
  //OR U152
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U152 (
    .O(n809),
    .I0(in[187]),
    .I1(in[177])
  );
  //AND U152bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U152bar (
    .O(n809bar),
    .I0(inbar[187]),
    .I1(inbar[177])
  );
  //OR U153
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U153 (
    .O(n810),
    .I0(in[200]),
    .I1(in[192])
  );
  //AND U153bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U153bar (
    .O(n810bar),
    .I0(inbar[200]),
    .I1(inbar[192])
  );
  //OR U154
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U154 (
    .O(n816),
    .I0(n808),
    .I1(n807)
  );
  //AND U154bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U154bar (
    .O(n816bar),
    .I0(n808bar),
    .I1(n807bar)
  );
  //OR U155
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U155 (
    .O(n807),
    .I0(n806),
    .I1(n805)
  );
  //AND U155bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U155bar (
    .O(n807bar),
    .I0(n806bar),
    .I1(n805bar)
  );
  //OR U156
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U156 (
    .O(n805),
    .I0(in[225]),
    .I1(in[207])
  );
  //AND U156bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U156bar (
    .O(n805bar),
    .I0(inbar[225]),
    .I1(inbar[207])
  );
  //OR U157
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U157 (
    .O(n806),
    .I0(in[98]),
    .I1(in[226])
  );
  //AND U157bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U157bar (
    .O(n806bar),
    .I0(inbar[98]),
    .I1(inbar[226])
  );
  //OR U158
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U158 (
    .O(n808),
    .I0(n804),
    .I1(n803)
  );
  //AND U158bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U158bar (
    .O(n808bar),
    .I0(n804bar),
    .I1(n803bar)
  );
  //OR U159
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U159 (
    .O(n803),
    .I0(in_20),
    .I1(in_16)
  );
  //AND U159bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U159bar (
    .O(n803bar),
    .I0(in_20bar),
    .I1(in_16bar)
  );
  //OR U160
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U160 (
    .O(n804),
    .I0(in_55),
    .I1(in_45)
  );
  //AND U160bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U160bar (
    .O(n804bar),
    .I0(in_55bar),
    .I1(in_45bar)
  );
  //OR U161
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U161 (
    .O(n824),
    .I0(n802),
    .I1(n801)
  );
  //AND U161bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U161bar (
    .O(n824bar),
    .I0(n802bar),
    .I1(n801bar)
  );
  //OR U162
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U162 (
    .O(n801),
    .I0(in[162]),
    .I1(in[149])
  );
  //AND U162bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U162bar (
    .O(n801bar),
    .I0(inbar[162]),
    .I1(inbar[149])
  );
  //OR U163
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U163 (
    .O(n802),
    .I0(in[163]),
    .I1(n800)
  );
  //AND U163bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U163bar (
    .O(n802bar),
    .I0(inbar[163]),
    .I1(n800bar)
  );
  //OR U164
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U164 (
    .O(n800),
    .I0(in[191]),
    .I1(in[189])
  );
  //AND U164bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U164bar (
    .O(n800bar),
    .I0(inbar[191]),
    .I1(inbar[189])
  );
  //OR U165
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U165 (
    .O(n826),
    .I0(n799),
    .I1(n798)
  );
  //AND U165bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U165bar (
    .O(n826bar),
    .I0(n799bar),
    .I1(n798bar)
  );
  //OR U166
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U166 (
    .O(n798),
    .I0(n797),
    .I1(n796)
  );
  //AND U166bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U166bar (
    .O(n798bar),
    .I0(n797bar),
    .I1(n796bar)
  );
  //OR U167
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U167 (
    .O(n796),
    .I0(in[212]),
    .I1(in[193])
  );
  //AND U167bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U167bar (
    .O(n796bar),
    .I0(inbar[212]),
    .I1(inbar[193])
  );
  //OR U168
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U168 (
    .O(n797),
    .I0(in[238]),
    .I1(n795)
  );
  //AND U168bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U168bar (
    .O(n797bar),
    .I0(inbar[238]),
    .I1(n795bar)
  );
  //OR U169
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U169 (
    .O(n795),
    .I0(in[88]),
    .I1(in[247])
  );
  //AND U169bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U169bar (
    .O(n795bar),
    .I0(inbar[88]),
    .I1(inbar[247])
  );
  //OR U170
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U170 (
    .O(n799),
    .I0(n794),
    .I1(n793)
  );
  //AND U170bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U170bar (
    .O(n799bar),
    .I0(n794bar),
    .I1(n793bar)
  );
  //OR U171
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U171 (
    .O(n793),
    .I0(in[94]),
    .I1(in[92])
  );
  //AND U171bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U171bar (
    .O(n793bar),
    .I0(inbar[94]),
    .I1(inbar[92])
  );
  //OR U172
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U172 (
    .O(n794),
    .I0(in_52),
    .I1(n792)
  );
  //AND U172bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U172bar (
    .O(n794bar),
    .I0(in_52bar),
    .I1(n792bar)
  );
  //OR U173
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U173 (
    .O(n792),
    .I0(in_70),
    .I1(in_67)
  );
  //AND U173bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U173bar (
    .O(n792bar),
    .I0(in_70bar),
    .I1(in_67bar)
  );
  //OR U174
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U174 (
    .O(out[2]),
    .I0(n791),
    .I1(n790)
  );
  //AND U174bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U174bar (
    .O(outbar[2]),
    .I0(n791bar),
    .I1(n790bar)
  );
  //OR U175
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U175 (
    .O(n790),
    .I0(n789),
    .I1(n788)
  );
  //AND U175bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U175bar (
    .O(n790bar),
    .I0(n789bar),
    .I1(n788bar)
  );
  //OR U176
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U176 (
    .O(n788),
    .I0(n787),
    .I1(n786)
  );
  //AND U176bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U176bar (
    .O(n788bar),
    .I0(n787bar),
    .I1(n786bar)
  );
  //OR U177
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U177 (
    .O(n786),
    .I0(n819),
    .I1(n785)
  );
  //AND U177bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U177bar (
    .O(n786bar),
    .I0(n819bar),
    .I1(n785bar)
  );
  //OR U178
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U178 (
    .O(n819),
    .I0(n784),
    .I1(n783)
  );
  //AND U178bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U178bar (
    .O(n819bar),
    .I0(n784bar),
    .I1(n783bar)
  );
  //OR U179
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U179 (
    .O(n783),
    .I0(n782),
    .I1(n781)
  );
  //AND U179bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U179bar (
    .O(n783bar),
    .I0(n782bar),
    .I1(n781bar)
  );
  //OR U180
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U180 (
    .O(n781),
    .I0(n780),
    .I1(n779)
  );
  //AND U180bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U180bar (
    .O(n781bar),
    .I0(n780bar),
    .I1(n779bar)
  );
  //OR U181
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U181 (
    .O(n779),
    .I0(n962),
    .I1(n778)
  );
  //AND U181bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U181bar (
    .O(n779bar),
    .I0(n962bar),
    .I1(n778bar)
  );
  //OR U182
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U182 (
    .O(n962),
    .I0(n777),
    .I1(n776)
  );
  //AND U182bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U182bar (
    .O(n962bar),
    .I0(n777bar),
    .I1(n776bar)
  );
  //OR U183
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U183 (
    .O(n776),
    .I0(n775),
    .I1(n774)
  );
  //AND U183bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U183bar (
    .O(n776bar),
    .I0(n775bar),
    .I1(n774bar)
  );
  //OR U184
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U184 (
    .O(n774),
    .I0(n773),
    .I1(n772)
  );
  //AND U184bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U184bar (
    .O(n774bar),
    .I0(n773bar),
    .I1(n772bar)
  );
  //OR U185
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U185 (
    .O(n772),
    .I0(in[131]),
    .I1(in[120])
  );
  //AND U185bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U185bar (
    .O(n772bar),
    .I0(inbar[131]),
    .I1(inbar[120])
  );
  //OR U186
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U186 (
    .O(n773),
    .I0(in[153]),
    .I1(in[147])
  );
  //AND U186bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U186bar (
    .O(n773bar),
    .I0(inbar[153]),
    .I1(inbar[147])
  );
  //OR U187
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U187 (
    .O(n775),
    .I0(n771),
    .I1(n770)
  );
  //AND U187bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U187bar (
    .O(n775bar),
    .I0(n771bar),
    .I1(n770bar)
  );
  //OR U188
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U188 (
    .O(n770),
    .I0(in[170]),
    .I1(in[156])
  );
  //AND U188bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U188bar (
    .O(n770bar),
    .I0(inbar[170]),
    .I1(inbar[156])
  );
  //OR U189
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U189 (
    .O(n771),
    .I0(in[223]),
    .I1(in[190])
  );
  //AND U189bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U189bar (
    .O(n771bar),
    .I0(inbar[223]),
    .I1(inbar[190])
  );
  //OR U190
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U190 (
    .O(n777),
    .I0(n769),
    .I1(n768)
  );
  //AND U190bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U190bar (
    .O(n777bar),
    .I0(n769bar),
    .I1(n768bar)
  );
  //OR U191
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U191 (
    .O(n768),
    .I0(n767),
    .I1(n766)
  );
  //AND U191bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U191bar (
    .O(n768bar),
    .I0(n767bar),
    .I1(n766bar)
  );
  //OR U192
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U192 (
    .O(n766),
    .I0(in[236]),
    .I1(in[230])
  );
  //AND U192bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U192bar (
    .O(n766bar),
    .I0(inbar[236]),
    .I1(inbar[230])
  );
  //OR U193
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U193 (
    .O(n767),
    .I0(in[85]),
    .I1(in[240])
  );
  //AND U193bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U193bar (
    .O(n767bar),
    .I0(inbar[85]),
    .I1(inbar[240])
  );
  //OR U194
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U194 (
    .O(n769),
    .I0(n765),
    .I1(n764)
  );
  //AND U194bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U194bar (
    .O(n769bar),
    .I0(n765bar),
    .I1(n764bar)
  );
  //OR U195
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U195 (
    .O(n764),
    .I0(in_12),
    .I1(in[90])
  );
  //AND U195bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U195bar (
    .O(n764bar),
    .I0(in_12bar),
    .I1(inbar[90])
  );
  //OR U196
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U196 (
    .O(n765),
    .I0(in_39),
    .I1(in_28)
  );
  //AND U196bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U196bar (
    .O(n765bar),
    .I0(in_39bar),
    .I1(in_28bar)
  );
  //OR U197
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U197 (
    .O(n780),
    .I0(in[109]),
    .I1(n763)
  );
  //AND U197bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U197bar (
    .O(n780bar),
    .I0(inbar[109]),
    .I1(n763bar)
  );
  //OR U198
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U198 (
    .O(n782),
    .I0(n762),
    .I1(n761)
  );
  //AND U198bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U198bar (
    .O(n782bar),
    .I0(n762bar),
    .I1(n761bar)
  );
  //OR U199
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U199 (
    .O(n761),
    .I0(in[138]),
    .I1(in[129])
  );
  //AND U199bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U199bar (
    .O(n761bar),
    .I0(inbar[138]),
    .I1(inbar[129])
  );
  //OR U200
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U200 (
    .O(n762),
    .I0(in[157]),
    .I1(n760)
  );
  //AND U200bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U200bar (
    .O(n762bar),
    .I0(inbar[157]),
    .I1(n760bar)
  );
  //OR U201
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U201 (
    .O(n760),
    .I0(in[182]),
    .I1(in[167])
  );
  //AND U201bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U201bar (
    .O(n760bar),
    .I0(inbar[182]),
    .I1(inbar[167])
  );
  //OR U202
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U202 (
    .O(n784),
    .I0(n759),
    .I1(n758)
  );
  //AND U202bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U202bar (
    .O(n784bar),
    .I0(n759bar),
    .I1(n758bar)
  );
  //OR U203
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U203 (
    .O(n758),
    .I0(n757),
    .I1(n756)
  );
  //AND U203bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U203bar (
    .O(n758bar),
    .I0(n757bar),
    .I1(n756bar)
  );
  //OR U204
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U204 (
    .O(n756),
    .I0(in[195]),
    .I1(in[184])
  );
  //AND U204bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U204bar (
    .O(n756bar),
    .I0(inbar[195]),
    .I1(inbar[184])
  );
  //OR U205
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U205 (
    .O(n757),
    .I0(in[196]),
    .I1(n755)
  );
  //AND U205bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U205bar (
    .O(n757bar),
    .I0(inbar[196]),
    .I1(n755bar)
  );
  //OR U206
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U206 (
    .O(n755),
    .I0(in[215]),
    .I1(in[209])
  );
  //AND U206bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U206bar (
    .O(n755bar),
    .I0(inbar[215]),
    .I1(inbar[209])
  );
  //OR U207
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U207 (
    .O(n759),
    .I0(n754),
    .I1(n753)
  );
  //AND U207bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U207bar (
    .O(n759bar),
    .I0(n754bar),
    .I1(n753bar)
  );
  //OR U208
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U208 (
    .O(n753),
    .I0(in[93]),
    .I1(in[233])
  );
  //AND U208bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U208bar (
    .O(n753bar),
    .I0(inbar[93]),
    .I1(inbar[233])
  );
  //OR U209
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U209 (
    .O(n754),
    .I0(in_1),
    .I1(n752)
  );
  //AND U209bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U209bar (
    .O(n754bar),
    .I0(in_1bar),
    .I1(n752bar)
  );
  //OR U210
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U210 (
    .O(n752),
    .I0(in_69),
    .I1(in_66)
  );
  //AND U210bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U210bar (
    .O(n752bar),
    .I0(in_69bar),
    .I1(in_66bar)
  );
  //OR U211
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U211 (
    .O(n787),
    .I0(n966),
    .I1(n751)
  );
  //AND U211bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U211bar (
    .O(n787bar),
    .I0(n966bar),
    .I1(n751bar)
  );
  //OR U212
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U212 (
    .O(n751),
    .I0(in[134]),
    .I1(n750)
  );
  //AND U212bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U212bar (
    .O(n751bar),
    .I0(inbar[134]),
    .I1(n750bar)
  );
  //OR U213
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U213 (
    .O(n966),
    .I0(n749),
    .I1(n748)
  );
  //AND U213bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U213bar (
    .O(n966bar),
    .I0(n749bar),
    .I1(n748bar)
  );
  //OR U214
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U214 (
    .O(n748),
    .I0(n747),
    .I1(n746)
  );
  //AND U214bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U214bar (
    .O(n748bar),
    .I0(n747bar),
    .I1(n746bar)
  );
  //OR U215
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U215 (
    .O(n746),
    .I0(n745),
    .I1(n744)
  );
  //AND U215bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U215bar (
    .O(n746bar),
    .I0(n745bar),
    .I1(n744bar)
  );
  //OR U216
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U216 (
    .O(n744),
    .I0(in[136]),
    .I1(in[121])
  );
  //AND U216bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U216bar (
    .O(n744bar),
    .I0(inbar[136]),
    .I1(inbar[121])
  );
  //OR U217
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U217 (
    .O(n745),
    .I0(in[186]),
    .I1(in[174])
  );
  //AND U217bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U217bar (
    .O(n745bar),
    .I0(inbar[186]),
    .I1(inbar[174])
  );
  //OR U218
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U218 (
    .O(n747),
    .I0(n743),
    .I1(n742)
  );
  //AND U218bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U218bar (
    .O(n747bar),
    .I0(n743bar),
    .I1(n742bar)
  );
  //OR U219
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U219 (
    .O(n742),
    .I0(in[198]),
    .I1(in[197])
  );
  //AND U219bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U219bar (
    .O(n742bar),
    .I0(inbar[198]),
    .I1(inbar[197])
  );
  //OR U220
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U220 (
    .O(n743),
    .I0(in[214]),
    .I1(in[199])
  );
  //AND U220bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U220bar (
    .O(n743bar),
    .I0(inbar[214]),
    .I1(inbar[199])
  );
  //OR U221
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U221 (
    .O(n749),
    .I0(n741),
    .I1(n740)
  );
  //AND U221bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U221bar (
    .O(n749bar),
    .I0(n741bar),
    .I1(n740bar)
  );
  //OR U222
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U222 (
    .O(n740),
    .I0(n739),
    .I1(n738)
  );
  //AND U222bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U222bar (
    .O(n740bar),
    .I0(n739bar),
    .I1(n738bar)
  );
  //OR U223
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U223 (
    .O(n738),
    .I0(in[231]),
    .I1(in[220])
  );
  //AND U223bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U223bar (
    .O(n738bar),
    .I0(inbar[231]),
    .I1(inbar[220])
  );
  //OR U224
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U224 (
    .O(n739),
    .I0(in_25),
    .I1(in[245])
  );
  //AND U224bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U224bar (
    .O(n739bar),
    .I0(in_25bar),
    .I1(inbar[245])
  );
  //OR U225
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U225 (
    .O(n741),
    .I0(n737),
    .I1(n736)
  );
  //AND U225bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U225bar (
    .O(n741bar),
    .I0(n737bar),
    .I1(n736bar)
  );
  //OR U226
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U226 (
    .O(n736),
    .I0(in_53),
    .I1(in_29)
  );
  //AND U226bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U226bar (
    .O(n736bar),
    .I0(in_53bar),
    .I1(in_29bar)
  );
  //OR U227
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U227 (
    .O(n737),
    .I0(in_79),
    .I1(in_74)
  );
  //AND U227bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U227bar (
    .O(n737bar),
    .I0(in_79bar),
    .I1(in_74bar)
  );
  //OR U228
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U228 (
    .O(n789),
    .I0(n735),
    .I1(n734)
  );
  //AND U228bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U228bar (
    .O(n789bar),
    .I0(n735bar),
    .I1(n734bar)
  );
  //OR U229
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U229 (
    .O(n734),
    .I0(in[152]),
    .I1(in[140])
  );
  //AND U229bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U229bar (
    .O(n734bar),
    .I0(inbar[152]),
    .I1(inbar[140])
  );
  //OR U230
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U230 (
    .O(n735),
    .I0(in[155]),
    .I1(n733)
  );
  //AND U230bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U230bar (
    .O(n735bar),
    .I0(inbar[155]),
    .I1(n733bar)
  );
  //OR U231
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U231 (
    .O(n733),
    .I0(in[166]),
    .I1(in[165])
  );
  //AND U231bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U231bar (
    .O(n733bar),
    .I0(inbar[166]),
    .I1(inbar[165])
  );
  //OR U232
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U232 (
    .O(n791),
    .I0(n732),
    .I1(n731)
  );
  //AND U232bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U232bar (
    .O(n791bar),
    .I0(n732bar),
    .I1(n731bar)
  );
  //OR U233
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U233 (
    .O(n731),
    .I0(n730),
    .I1(n729)
  );
  //AND U233bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U233bar (
    .O(n731bar),
    .I0(n730bar),
    .I1(n729bar)
  );
  //OR U234
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U234 (
    .O(n729),
    .I0(in[202]),
    .I1(in[185])
  );
  //AND U234bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U234bar (
    .O(n729bar),
    .I0(inbar[202]),
    .I1(inbar[185])
  );
  //OR U235
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U235 (
    .O(n730),
    .I0(in[211]),
    .I1(n728)
  );
  //AND U235bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U235bar (
    .O(n730bar),
    .I0(inbar[211]),
    .I1(n728bar)
  );
  //OR U236
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U236 (
    .O(n728),
    .I0(in[255]),
    .I1(in[253])
  );
  //AND U236bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U236bar (
    .O(n728bar),
    .I0(inbar[255]),
    .I1(inbar[253])
  );
  //OR U237
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U237 (
    .O(n732),
    .I0(n727),
    .I1(n726)
  );
  //AND U237bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U237bar (
    .O(n732bar),
    .I0(n727bar),
    .I1(n726bar)
  );
  //OR U238
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U238 (
    .O(n726),
    .I0(in_35),
    .I1(in_15)
  );
  //AND U238bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U238bar (
    .O(n726bar),
    .I0(in_35bar),
    .I1(in_15bar)
  );
  //OR U239
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U239 (
    .O(n727),
    .I0(in_36),
    .I1(n725)
  );
  //AND U239bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U239bar (
    .O(n727bar),
    .I0(in_36bar),
    .I1(n725bar)
  );
  //OR U240
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U240 (
    .O(n725),
    .I0(in_48),
    .I1(in_40)
  );
  //AND U240bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U240bar (
    .O(n725bar),
    .I0(in_48bar),
    .I1(in_40bar)
  );
  //OR U241
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U241 (
    .O(out[1]),
    .I0(n724),
    .I1(n723)
  );
  //AND U241bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U241bar (
    .O(outbar[1]),
    .I0(n724bar),
    .I1(n723bar)
  );
  //OR U242
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U242 (
    .O(n723),
    .I0(n722),
    .I1(n721)
  );
  //AND U242bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U242bar (
    .O(n723bar),
    .I0(n722bar),
    .I1(n721bar)
  );
  //OR U243
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U243 (
    .O(n721),
    .I0(n720),
    .I1(n719)
  );
  //AND U243bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U243bar (
    .O(n721bar),
    .I0(n720bar),
    .I1(n719bar)
  );
  //OR U244
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U244 (
    .O(n719),
    .I0(n921),
    .I1(n887)
  );
  //AND U244bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U244bar (
    .O(n719bar),
    .I0(n921bar),
    .I1(n887bar)
  );
  //OR U245
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U245 (
    .O(n887),
    .I0(n718),
    .I1(n717)
  );
  //AND U245bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U245bar (
    .O(n887bar),
    .I0(n718bar),
    .I1(n717bar)
  );
  //OR U246
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U246 (
    .O(n717),
    .I0(n716),
    .I1(n715)
  );
  //AND U246bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U246bar (
    .O(n717bar),
    .I0(n716bar),
    .I1(n715bar)
  );
  //OR U247
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U247 (
    .O(n715),
    .I0(n714),
    .I1(n713)
  );
  //AND U247bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U247bar (
    .O(n715bar),
    .I0(n714bar),
    .I1(n713bar)
  );
  //OR U248
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U248 (
    .O(n713),
    .I0(in[116]),
    .I1(in[110])
  );
  //AND U248bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U248bar (
    .O(n713bar),
    .I0(inbar[116]),
    .I1(inbar[110])
  );
  //OR U249
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U249 (
    .O(n714),
    .I0(in[133]),
    .I1(in[130])
  );
  //AND U249bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U249bar (
    .O(n714bar),
    .I0(inbar[133]),
    .I1(inbar[130])
  );
  //OR U250
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U250 (
    .O(n716),
    .I0(n712),
    .I1(n711)
  );
  //AND U250bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U250bar (
    .O(n716bar),
    .I0(n712bar),
    .I1(n711bar)
  );
  //OR U251
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U251 (
    .O(n711),
    .I0(in[203]),
    .I1(in[135])
  );
  //AND U251bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U251bar (
    .O(n711bar),
    .I0(inbar[203]),
    .I1(inbar[135])
  );
  //OR U252
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U252 (
    .O(n712),
    .I0(in[232]),
    .I1(in[223])
  );
  //AND U252bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U252bar (
    .O(n712bar),
    .I0(inbar[232]),
    .I1(inbar[223])
  );
  //OR U253
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U253 (
    .O(n718),
    .I0(n710),
    .I1(n709)
  );
  //AND U253bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U253bar (
    .O(n718bar),
    .I0(n710bar),
    .I1(n709bar)
  );
  //OR U254
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U254 (
    .O(n709),
    .I0(n708),
    .I1(n707)
  );
  //AND U254bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U254bar (
    .O(n709bar),
    .I0(n708bar),
    .I1(n707bar)
  );
  //OR U255
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U255 (
    .O(n707),
    .I0(in[255]),
    .I1(in[233])
  );
  //AND U255bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U255bar (
    .O(n707bar),
    .I0(inbar[255]),
    .I1(inbar[233])
  );
  //OR U256
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U256 (
    .O(n708),
    .I0(in_53),
    .I1(in_34)
  );
  //AND U256bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U256bar (
    .O(n708bar),
    .I0(in_53bar),
    .I1(in_34bar)
  );
  //OR U257
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U257 (
    .O(n710),
    .I0(n706),
    .I1(n705)
  );
  //AND U257bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U257bar (
    .O(n710bar),
    .I0(n706bar),
    .I1(n705bar)
  );
  //OR U258
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U258 (
    .O(n705),
    .I0(in_57),
    .I1(in_55)
  );
  //AND U258bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U258bar (
    .O(n705bar),
    .I0(in_57bar),
    .I1(in_55bar)
  );
  //OR U259
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U259 (
    .O(n706),
    .I0(in_68),
    .I1(in_67)
  );
  //AND U259bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U259bar (
    .O(n706bar),
    .I0(in_68bar),
    .I1(in_67bar)
  );
  //OR U260
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U260 (
    .O(n921),
    .I0(n704),
    .I1(n703)
  );
  //AND U260bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U260bar (
    .O(n921bar),
    .I0(n704bar),
    .I1(n703bar)
  );
  //OR U261
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U261 (
    .O(n703),
    .I0(n702),
    .I1(n701)
  );
  //AND U261bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U261bar (
    .O(n703bar),
    .I0(n702bar),
    .I1(n701bar)
  );
  //OR U262
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U262 (
    .O(n701),
    .I0(n700),
    .I1(n699)
  );
  //AND U262bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U262bar (
    .O(n701bar),
    .I0(n700bar),
    .I1(n699bar)
  );
  //OR U263
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U263 (
    .O(n699),
    .I0(n944),
    .I1(n872)
  );
  //AND U263bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U263bar (
    .O(n699bar),
    .I0(n944bar),
    .I1(n872bar)
  );
  //OR U264
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U264 (
    .O(n872),
    .I0(n698),
    .I1(n697)
  );
  //AND U264bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U264bar (
    .O(n872bar),
    .I0(n698bar),
    .I1(n697bar)
  );
  //OR U265
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U265 (
    .O(n697),
    .I0(n696),
    .I1(n695)
  );
  //AND U265bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U265bar (
    .O(n697bar),
    .I0(n696bar),
    .I1(n695bar)
  );
  //OR U266
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U266 (
    .O(n695),
    .I0(n694),
    .I1(n693)
  );
  //AND U266bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U266bar (
    .O(n695bar),
    .I0(n694bar),
    .I1(n693bar)
  );
  //OR U267
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U267 (
    .O(n693),
    .I0(in[121]),
    .I1(in[102])
  );
  //AND U267bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U267bar (
    .O(n693bar),
    .I0(inbar[121]),
    .I1(inbar[102])
  );
  //OR U268
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U268 (
    .O(n694),
    .I0(in[162]),
    .I1(in[161])
  );
  //AND U268bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U268bar (
    .O(n694bar),
    .I0(inbar[162]),
    .I1(inbar[161])
  );
  //OR U269
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U269 (
    .O(n696),
    .I0(n692),
    .I1(n691)
  );
  //AND U269bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U269bar (
    .O(n696bar),
    .I0(n692bar),
    .I1(n691bar)
  );
  //OR U270
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U270 (
    .O(n691),
    .I0(in[192]),
    .I1(in[178])
  );
  //AND U270bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U270bar (
    .O(n691bar),
    .I0(inbar[192]),
    .I1(inbar[178])
  );
  //OR U271
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U271 (
    .O(n692),
    .I0(in[244]),
    .I1(in[209])
  );
  //AND U271bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U271bar (
    .O(n692bar),
    .I0(inbar[244]),
    .I1(inbar[209])
  );
  //OR U272
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U272 (
    .O(n698),
    .I0(n690),
    .I1(n689)
  );
  //AND U272bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U272bar (
    .O(n698bar),
    .I0(n690bar),
    .I1(n689bar)
  );
  //OR U273
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U273 (
    .O(n689),
    .I0(n688),
    .I1(n687)
  );
  //AND U273bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U273bar (
    .O(n689bar),
    .I0(n688bar),
    .I1(n687bar)
  );
  //OR U274
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U274 (
    .O(n687),
    .I0(in[90]),
    .I1(in[254])
  );
  //AND U274bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U274bar (
    .O(n687bar),
    .I0(inbar[90]),
    .I1(inbar[254])
  );
  //OR U275
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U275 (
    .O(n688),
    .I0(in_36),
    .I1(in_32)
  );
  //AND U275bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U275bar (
    .O(n688bar),
    .I0(in_36bar),
    .I1(in_32bar)
  );
  //OR U276
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U276 (
    .O(n690),
    .I0(n686),
    .I1(n685)
  );
  //AND U276bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U276bar (
    .O(n690bar),
    .I0(n686bar),
    .I1(n685bar)
  );
  //OR U277
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U277 (
    .O(n685),
    .I0(in_62),
    .I1(in_37)
  );
  //AND U277bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U277bar (
    .O(n685bar),
    .I0(in_62bar),
    .I1(in_37bar)
  );
  //OR U278
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U278 (
    .O(n686),
    .I0(in_75),
    .I1(in_73)
  );
  //AND U278bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U278bar (
    .O(n686bar),
    .I0(in_75bar),
    .I1(in_73bar)
  );
  //OR U279
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U279 (
    .O(n944),
    .I0(n684),
    .I1(n683)
  );
  //AND U279bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U279bar (
    .O(n944bar),
    .I0(n684bar),
    .I1(n683bar)
  );
  //OR U280
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U280 (
    .O(n683),
    .I0(n682),
    .I1(n681)
  );
  //AND U280bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U280bar (
    .O(n683bar),
    .I0(n682bar),
    .I1(n681bar)
  );
  //OR U281
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U281 (
    .O(n681),
    .I0(n680),
    .I1(n679)
  );
  //AND U281bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U281bar (
    .O(n681bar),
    .I0(n680bar),
    .I1(n679bar)
  );
  //OR U282
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U282 (
    .O(n679),
    .I0(in[171]),
    .I1(in[153])
  );
  //AND U282bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U282bar (
    .O(n679bar),
    .I0(inbar[171]),
    .I1(inbar[153])
  );
  //OR U283
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U283 (
    .O(n680),
    .I0(in[187]),
    .I1(in[176])
  );
  //AND U283bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U283bar (
    .O(n680bar),
    .I0(inbar[187]),
    .I1(inbar[176])
  );
  //OR U284
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U284 (
    .O(n682),
    .I0(n678),
    .I1(n677)
  );
  //AND U284bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U284bar (
    .O(n682bar),
    .I0(n678bar),
    .I1(n677bar)
  );
  //OR U285
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U285 (
    .O(n677),
    .I0(in[245]),
    .I1(in[211])
  );
  //AND U285bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U285bar (
    .O(n677bar),
    .I0(inbar[245]),
    .I1(inbar[211])
  );
  //OR U286
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U286 (
    .O(n678),
    .I0(in[97]),
    .I1(in[88])
  );
  //AND U286bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U286bar (
    .O(n678bar),
    .I0(inbar[97]),
    .I1(inbar[88])
  );
  //OR U287
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U287 (
    .O(n684),
    .I0(n676),
    .I1(n675)
  );
  //AND U287bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U287bar (
    .O(n684bar),
    .I0(n676bar),
    .I1(n675bar)
  );
  //OR U288
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U288 (
    .O(n675),
    .I0(n674),
    .I1(n673)
  );
  //AND U288bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U288bar (
    .O(n675bar),
    .I0(n674bar),
    .I1(n673bar)
  );
  //OR U289
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U289 (
    .O(n673),
    .I0(in_10),
    .I1(in_0)
  );
  //AND U289bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U289bar (
    .O(n673bar),
    .I0(in_10bar),
    .I1(in_0bar)
  );
  //OR U290
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U290 (
    .O(n674),
    .I0(in_59),
    .I1(in_5)
  );
  //AND U290bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U290bar (
    .O(n674bar),
    .I0(in_59bar),
    .I1(in_5bar)
  );
  //OR U291
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U291 (
    .O(n676),
    .I0(n672),
    .I1(n671)
  );
  //AND U291bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U291bar (
    .O(n676bar),
    .I0(n672bar),
    .I1(n671bar)
  );
  //OR U292
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U292 (
    .O(n671),
    .I0(in_60),
    .I1(in_6)
  );
  //AND U292bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U292bar (
    .O(n671bar),
    .I0(in_60bar),
    .I1(in_6bar)
  );
  //OR U293
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U293 (
    .O(n672),
    .I0(in_77),
    .I1(in_69)
  );
  //AND U293bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U293bar (
    .O(n672bar),
    .I0(in_77bar),
    .I1(in_69bar)
  );
  //OR U294
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U294 (
    .O(n700),
    .I0(in[113]),
    .I1(n864)
  );
  //AND U294bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U294bar (
    .O(n700bar),
    .I0(inbar[113]),
    .I1(n864bar)
  );
  //OR U295
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U295 (
    .O(n864),
    .I0(n670),
    .I1(n669)
  );
  //AND U295bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U295bar (
    .O(n864bar),
    .I0(n670bar),
    .I1(n669bar)
  );
  //OR U296
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U296 (
    .O(n669),
    .I0(n668),
    .I1(n667)
  );
  //AND U296bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U296bar (
    .O(n669bar),
    .I0(n668bar),
    .I1(n667bar)
  );
  //OR U297
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U297 (
    .O(n667),
    .I0(n666),
    .I1(n665)
  );
  //AND U297bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U297bar (
    .O(n667bar),
    .I0(n666bar),
    .I1(n665bar)
  );
  //OR U298
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U298 (
    .O(n665),
    .I0(in[125]),
    .I1(in[107])
  );
  //AND U298bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U298bar (
    .O(n665bar),
    .I0(inbar[125]),
    .I1(inbar[107])
  );
  //OR U299
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U299 (
    .O(n666),
    .I0(in[138]),
    .I1(in[126])
  );
  //AND U299bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U299bar (
    .O(n666bar),
    .I0(inbar[138]),
    .I1(inbar[126])
  );
  //OR U300
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U300 (
    .O(n668),
    .I0(n664),
    .I1(n663)
  );
  //AND U300bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U300bar (
    .O(n668bar),
    .I0(n664bar),
    .I1(n663bar)
  );
  //OR U301
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U301 (
    .O(n663),
    .I0(in[189]),
    .I1(in[143])
  );
  //AND U301bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U301bar (
    .O(n663bar),
    .I0(inbar[189]),
    .I1(inbar[143])
  );
  //OR U302
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U302 (
    .O(n664),
    .I0(in[99]),
    .I1(in[214])
  );
  //AND U302bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U302bar (
    .O(n664bar),
    .I0(inbar[99]),
    .I1(inbar[214])
  );
  //OR U303
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U303 (
    .O(n670),
    .I0(n662),
    .I1(n661)
  );
  //AND U303bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U303bar (
    .O(n670bar),
    .I0(n662bar),
    .I1(n661bar)
  );
  //OR U304
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U304 (
    .O(n661),
    .I0(n660),
    .I1(n659)
  );
  //AND U304bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U304bar (
    .O(n661bar),
    .I0(n660bar),
    .I1(n659bar)
  );
  //OR U305
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U305 (
    .O(n659),
    .I0(in_15),
    .I1(in_12)
  );
  //AND U305bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U305bar (
    .O(n659bar),
    .I0(in_15bar),
    .I1(in_12bar)
  );
  //OR U306
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U306 (
    .O(n660),
    .I0(in_20),
    .I1(in_2)
  );
  //AND U306bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U306bar (
    .O(n660bar),
    .I0(in_20bar),
    .I1(in_2bar)
  );
  //OR U307
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U307 (
    .O(n662),
    .I0(n658),
    .I1(n657)
  );
  //AND U307bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U307bar (
    .O(n662bar),
    .I0(n658bar),
    .I1(n657bar)
  );
  //OR U308
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U308 (
    .O(n657),
    .I0(in_30),
    .I1(in_3)
  );
  //AND U308bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U308bar (
    .O(n657bar),
    .I0(in_30bar),
    .I1(in_3bar)
  );
  //OR U309
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U309 (
    .O(n658),
    .I0(in_4),
    .I1(in_38)
  );
  //AND U309bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U309bar (
    .O(n658bar),
    .I0(in_4bar),
    .I1(in_38bar)
  );
  //OR U310
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U310 (
    .O(n702),
    .I0(n656),
    .I1(n655)
  );
  //AND U310bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U310bar (
    .O(n702bar),
    .I0(n656bar),
    .I1(n655bar)
  );
  //OR U311
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U311 (
    .O(n655),
    .I0(in[148]),
    .I1(in[137])
  );
  //AND U311bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U311bar (
    .O(n655bar),
    .I0(inbar[148]),
    .I1(inbar[137])
  );
  //OR U312
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U312 (
    .O(n656),
    .I0(in[149]),
    .I1(n654)
  );
  //AND U312bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U312bar (
    .O(n656bar),
    .I0(inbar[149]),
    .I1(n654bar)
  );
  //OR U313
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U313 (
    .O(n654),
    .I0(in[195]),
    .I1(in[190])
  );
  //AND U313bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U313bar (
    .O(n654bar),
    .I0(inbar[195]),
    .I1(inbar[190])
  );
  //OR U314
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U314 (
    .O(n704),
    .I0(n653),
    .I1(n652)
  );
  //AND U314bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U314bar (
    .O(n704bar),
    .I0(n653bar),
    .I1(n652bar)
  );
  //OR U315
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U315 (
    .O(n652),
    .I0(n651),
    .I1(n650)
  );
  //AND U315bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U315bar (
    .O(n652bar),
    .I0(n651bar),
    .I1(n650bar)
  );
  //OR U316
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U316 (
    .O(n650),
    .I0(in[98]),
    .I1(in[197])
  );
  //AND U316bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U316bar (
    .O(n650bar),
    .I0(inbar[98]),
    .I1(inbar[197])
  );
  //OR U317
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U317 (
    .O(n651),
    .I0(in_11),
    .I1(n649)
  );
  //AND U317bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U317bar (
    .O(n651bar),
    .I0(in_11bar),
    .I1(n649bar)
  );
  //OR U318
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U318 (
    .O(n649),
    .I0(in_26),
    .I1(in_14)
  );
  //AND U318bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U318bar (
    .O(n649bar),
    .I0(in_26bar),
    .I1(in_14bar)
  );
  //OR U319
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U319 (
    .O(n653),
    .I0(n648),
    .I1(n647)
  );
  //AND U319bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U319bar (
    .O(n653bar),
    .I0(n648bar),
    .I1(n647bar)
  );
  //OR U320
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U320 (
    .O(n647),
    .I0(in_35),
    .I1(in_27)
  );
  //AND U320bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U320bar (
    .O(n647bar),
    .I0(in_35bar),
    .I1(in_27bar)
  );
  //OR U321
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U321 (
    .O(n648),
    .I0(in_50),
    .I1(n646)
  );
  //AND U321bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U321bar (
    .O(n648bar),
    .I0(in_50bar),
    .I1(n646bar)
  );
  //OR U322
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U322 (
    .O(n646),
    .I0(in_78),
    .I1(in_61)
  );
  //AND U322bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U322bar (
    .O(n646bar),
    .I0(in_78bar),
    .I1(in_61bar)
  );
  //OR U323
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U323 (
    .O(n720),
    .I0(n942),
    .I1(n645)
  );
  //AND U323bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U323bar (
    .O(n720bar),
    .I0(n942bar),
    .I1(n645bar)
  );
  //OR U324
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U324 (
    .O(n645),
    .I0(in[106]),
    .I1(n863)
  );
  //AND U324bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U324bar (
    .O(n645bar),
    .I0(inbar[106]),
    .I1(n863bar)
  );
  //OR U325
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U325 (
    .O(n863),
    .I0(n644),
    .I1(n643)
  );
  //AND U325bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U325bar (
    .O(n863bar),
    .I0(n644bar),
    .I1(n643bar)
  );
  //OR U326
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U326 (
    .O(n643),
    .I0(n642),
    .I1(n641)
  );
  //AND U326bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U326bar (
    .O(n643bar),
    .I0(n642bar),
    .I1(n641bar)
  );
  //OR U327
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U327 (
    .O(n641),
    .I0(n640),
    .I1(n639)
  );
  //AND U327bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U327bar (
    .O(n641bar),
    .I0(n640bar),
    .I1(n639bar)
  );
  //OR U328
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U328 (
    .O(n639),
    .I0(in[127]),
    .I1(in[122])
  );
  //AND U328bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U328bar (
    .O(n639bar),
    .I0(inbar[127]),
    .I1(inbar[122])
  );
  //OR U329
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U329 (
    .O(n640),
    .I0(in[156]),
    .I1(in[132])
  );
  //AND U329bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U329bar (
    .O(n640bar),
    .I0(inbar[156]),
    .I1(inbar[132])
  );
  //OR U330
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U330 (
    .O(n642),
    .I0(n638),
    .I1(n637)
  );
  //AND U330bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U330bar (
    .O(n642bar),
    .I0(n638bar),
    .I1(n637bar)
  );
  //OR U331
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U331 (
    .O(n637),
    .I0(in[159]),
    .I1(in[157])
  );
  //AND U331bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U331bar (
    .O(n637bar),
    .I0(inbar[159]),
    .I1(inbar[157])
  );
  //OR U332
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U332 (
    .O(n638),
    .I0(in[185]),
    .I1(in[169])
  );
  //AND U332bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U332bar (
    .O(n638bar),
    .I0(inbar[185]),
    .I1(inbar[169])
  );
  //OR U333
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U333 (
    .O(n644),
    .I0(n636),
    .I1(n635)
  );
  //AND U333bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U333bar (
    .O(n644bar),
    .I0(n636bar),
    .I1(n635bar)
  );
  //OR U334
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U334 (
    .O(n635),
    .I0(n634),
    .I1(n633)
  );
  //AND U334bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U334bar (
    .O(n635bar),
    .I0(n634bar),
    .I1(n633bar)
  );
  //OR U335
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U335 (
    .O(n633),
    .I0(in[239]),
    .I1(in[218])
  );
  //AND U335bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U335bar (
    .O(n633bar),
    .I0(inbar[239]),
    .I1(inbar[218])
  );
  //OR U336
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U336 (
    .O(n634),
    .I0(in_13),
    .I1(in[87])
  );
  //AND U336bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U336bar (
    .O(n634bar),
    .I0(in_13bar),
    .I1(inbar[87])
  );
  //OR U337
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U337 (
    .O(n636),
    .I0(n632),
    .I1(n631)
  );
  //AND U337bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U337bar (
    .O(n636bar),
    .I0(n632bar),
    .I1(n631bar)
  );
  //OR U338
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U338 (
    .O(n631),
    .I0(in_72),
    .I1(in_70)
  );
  //AND U338bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U338bar (
    .O(n631bar),
    .I0(in_72bar),
    .I1(in_70bar)
  );
  //OR U339
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U339 (
    .O(n632),
    .I0(in_80),
    .I1(in_74)
  );
  //AND U339bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U339bar (
    .O(n632bar),
    .I0(in_80bar),
    .I1(in_74bar)
  );
  //OR U340
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U340 (
    .O(n942),
    .I0(n630),
    .I1(n629)
  );
  //AND U340bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U340bar (
    .O(n942bar),
    .I0(n630bar),
    .I1(n629bar)
  );
  //OR U341
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U341 (
    .O(n629),
    .I0(n628),
    .I1(n627)
  );
  //AND U341bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U341bar (
    .O(n629bar),
    .I0(n628bar),
    .I1(n627bar)
  );
  //OR U342
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U342 (
    .O(n627),
    .I0(n626),
    .I1(n625)
  );
  //AND U342bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U342bar (
    .O(n627bar),
    .I0(n626bar),
    .I1(n625bar)
  );
  //OR U343
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U343 (
    .O(n625),
    .I0(in[146]),
    .I1(in[100])
  );
  //AND U343bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U343bar (
    .O(n625bar),
    .I0(inbar[146]),
    .I1(inbar[100])
  );
  //OR U344
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U344 (
    .O(n626),
    .I0(in[168]),
    .I1(in[152])
  );
  //AND U344bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U344bar (
    .O(n626bar),
    .I0(inbar[168]),
    .I1(inbar[152])
  );
  //OR U345
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U345 (
    .O(n628),
    .I0(n624),
    .I1(n623)
  );
  //AND U345bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U345bar (
    .O(n628bar),
    .I0(n624bar),
    .I1(n623bar)
  );
  //OR U346
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U346 (
    .O(n623),
    .I0(in[199]),
    .I1(in[182])
  );
  //AND U346bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U346bar (
    .O(n623bar),
    .I0(inbar[199]),
    .I1(inbar[182])
  );
  //OR U347
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U347 (
    .O(n624),
    .I0(in[236]),
    .I1(in[204])
  );
  //AND U347bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U347bar (
    .O(n624bar),
    .I0(inbar[236]),
    .I1(inbar[204])
  );
  //OR U348
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U348 (
    .O(n630),
    .I0(n622),
    .I1(n621)
  );
  //AND U348bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U348bar (
    .O(n630bar),
    .I0(n622bar),
    .I1(n621bar)
  );
  //OR U349
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U349 (
    .O(n621),
    .I0(n620),
    .I1(n619)
  );
  //AND U349bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U349bar (
    .O(n621bar),
    .I0(n620bar),
    .I1(n619bar)
  );
  //OR U350
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U350 (
    .O(n619),
    .I0(in[89]),
    .I1(in[246])
  );
  //AND U350bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U350bar (
    .O(n619bar),
    .I0(inbar[89]),
    .I1(inbar[246])
  );
  //OR U351
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U351 (
    .O(n620),
    .I0(in[95]),
    .I1(in[92])
  );
  //AND U351bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U351bar (
    .O(n620bar),
    .I0(inbar[95]),
    .I1(inbar[92])
  );
  //OR U352
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U352 (
    .O(n622),
    .I0(n618),
    .I1(n617)
  );
  //AND U352bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U352bar (
    .O(n622bar),
    .I0(n618bar),
    .I1(n617bar)
  );
  //OR U353
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U353 (
    .O(n617),
    .I0(in_22),
    .I1(in_16)
  );
  //AND U353bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U353bar (
    .O(n617bar),
    .I0(in_22bar),
    .I1(in_16bar)
  );
  //OR U354
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U354 (
    .O(n618),
    .I0(in_51),
    .I1(in_49)
  );
  //AND U354bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U354bar (
    .O(n618bar),
    .I0(in_51bar),
    .I1(in_49bar)
  );
  //OR U355
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U355 (
    .O(n722),
    .I0(n616),
    .I1(n615)
  );
  //AND U355bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U355bar (
    .O(n722bar),
    .I0(n616bar),
    .I1(n615bar)
  );
  //OR U356
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U356 (
    .O(n615),
    .I0(in[158]),
    .I1(in[115])
  );
  //AND U356bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U356bar (
    .O(n615bar),
    .I0(inbar[158]),
    .I1(inbar[115])
  );
  //OR U357
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U357 (
    .O(n616),
    .I0(in[163]),
    .I1(n614)
  );
  //AND U357bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U357bar (
    .O(n616bar),
    .I0(inbar[163]),
    .I1(n614bar)
  );
  //OR U358
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U358 (
    .O(n614),
    .I0(in[206]),
    .I1(in[165])
  );
  //AND U358bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U358bar (
    .O(n614bar),
    .I0(inbar[206]),
    .I1(inbar[165])
  );
  //OR U359
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U359 (
    .O(n724),
    .I0(n613),
    .I1(n612)
  );
  //AND U359bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U359bar (
    .O(n724bar),
    .I0(n613bar),
    .I1(n612bar)
  );
  //OR U360
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U360 (
    .O(n612),
    .I0(n611),
    .I1(n610)
  );
  //AND U360bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U360bar (
    .O(n612bar),
    .I0(n611bar),
    .I1(n610bar)
  );
  //OR U361
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U361 (
    .O(n610),
    .I0(in[213]),
    .I1(in[207])
  );
  //AND U361bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U361bar (
    .O(n610bar),
    .I0(inbar[213]),
    .I1(inbar[207])
  );
  //OR U362
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U362 (
    .O(n611),
    .I0(in[215]),
    .I1(n609)
  );
  //AND U362bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U362bar (
    .O(n611bar),
    .I0(inbar[215]),
    .I1(n609bar)
  );
  //OR U363
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U363 (
    .O(n609),
    .I0(in[230]),
    .I1(in[220])
  );
  //AND U363bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U363bar (
    .O(n609bar),
    .I0(inbar[230]),
    .I1(inbar[220])
  );
  //OR U364
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U364 (
    .O(n613),
    .I0(n608),
    .I1(n607)
  );
  //AND U364bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U364bar (
    .O(n613bar),
    .I0(n608bar),
    .I1(n607bar)
  );
  //OR U365
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U365 (
    .O(n607),
    .I0(in[251]),
    .I1(in[234])
  );
  //AND U365bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U365bar (
    .O(n607bar),
    .I0(inbar[251]),
    .I1(inbar[234])
  );
  //OR U366
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U366 (
    .O(n608),
    .I0(in_17),
    .I1(n606)
  );
  //AND U366bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U366bar (
    .O(n608bar),
    .I0(in_17bar),
    .I1(n606bar)
  );
  //OR U367
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U367 (
    .O(n606),
    .I0(in_65),
    .I1(in_56)
  );
  //AND U367bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U367bar (
    .O(n606bar),
    .I0(in_65bar),
    .I1(in_56bar)
  );
  //OR U368
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U368 (
    .O(out[0]),
    .I0(n605),
    .I1(n604)
  );
  //AND U368bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U368bar (
    .O(outbar[0]),
    .I0(n605bar),
    .I1(n604bar)
  );
  //OR U369
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U369 (
    .O(n604),
    .I0(n603),
    .I1(n602)
  );
  //AND U369bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U369bar (
    .O(n604bar),
    .I0(n603bar),
    .I1(n602bar)
  );
  //OR U370
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U370 (
    .O(n602),
    .I0(n601),
    .I1(n600)
  );
  //AND U370bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U370bar (
    .O(n602bar),
    .I0(n601bar),
    .I1(n600bar)
  );
  //OR U371
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U371 (
    .O(n600),
    .I0(n820),
    .I1(n785)
  );
  //AND U371bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U371bar (
    .O(n600bar),
    .I0(n820bar),
    .I1(n785bar)
  );
  //OR U372
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U372 (
    .O(n785),
    .I0(n599),
    .I1(n598)
  );
  //AND U372bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U372bar (
    .O(n785bar),
    .I0(n599bar),
    .I1(n598bar)
  );
  //OR U373
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U373 (
    .O(n598),
    .I0(n597),
    .I1(n596)
  );
  //AND U373bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U373bar (
    .O(n598bar),
    .I0(n597bar),
    .I1(n596bar)
  );
  //OR U374
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U374 (
    .O(n596),
    .I0(n595),
    .I1(n594)
  );
  //AND U374bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U374bar (
    .O(n596bar),
    .I0(n595bar),
    .I1(n594bar)
  );
  //OR U375
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U375 (
    .O(n594),
    .I0(in[135]),
    .I1(in[104])
  );
  //AND U375bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U375bar (
    .O(n594bar),
    .I0(inbar[135]),
    .I1(inbar[104])
  );
  //OR U376
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U376 (
    .O(n595),
    .I0(in[188]),
    .I1(in[178])
  );
  //AND U376bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U376bar (
    .O(n595bar),
    .I0(inbar[188]),
    .I1(inbar[178])
  );
  //OR U377
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U377 (
    .O(n597),
    .I0(n593),
    .I1(n592)
  );
  //AND U377bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U377bar (
    .O(n597bar),
    .I0(n593bar),
    .I1(n592bar)
  );
  //OR U378
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U378 (
    .O(n592),
    .I0(in[217]),
    .I1(in[194])
  );
  //AND U378bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U378bar (
    .O(n592bar),
    .I0(inbar[217]),
    .I1(inbar[194])
  );
  //OR U379
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U379 (
    .O(n593),
    .I0(in[237]),
    .I1(in[218])
  );
  //AND U379bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U379bar (
    .O(n593bar),
    .I0(inbar[237]),
    .I1(inbar[218])
  );
  //OR U380
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U380 (
    .O(n599),
    .I0(n591),
    .I1(n590)
  );
  //AND U380bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U380bar (
    .O(n599bar),
    .I0(n591bar),
    .I1(n590bar)
  );
  //OR U381
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U381 (
    .O(n590),
    .I0(n589),
    .I1(n588)
  );
  //AND U381bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U381bar (
    .O(n590bar),
    .I0(n589bar),
    .I1(n588bar)
  );
  //OR U382
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U382 (
    .O(n588),
    .I0(in_2),
    .I1(in_10)
  );
  //AND U382bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U382bar (
    .O(n588bar),
    .I0(in_2bar),
    .I1(in_10bar)
  );
  //OR U383
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U383 (
    .O(n589),
    .I0(in_47),
    .I1(in_22)
  );
  //AND U383bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U383bar (
    .O(n589bar),
    .I0(in_47bar),
    .I1(in_22bar)
  );
  //OR U384
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U384 (
    .O(n591),
    .I0(n587),
    .I1(n586)
  );
  //AND U384bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U384bar (
    .O(n591bar),
    .I0(n587bar),
    .I1(n586bar)
  );
  //OR U385
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U385 (
    .O(n586),
    .I0(in_56),
    .I1(in_54)
  );
  //AND U385bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U385bar (
    .O(n586bar),
    .I0(in_56bar),
    .I1(in_54bar)
  );
  //OR U386
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U386 (
    .O(n587),
    .I0(in_63),
    .I1(in_61)
  );
  //AND U386bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U386bar (
    .O(n587bar),
    .I0(in_63bar),
    .I1(in_61bar)
  );
  //OR U387
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U387 (
    .O(n820),
    .I0(n585),
    .I1(n584)
  );
  //AND U387bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U387bar (
    .O(n820bar),
    .I0(n585bar),
    .I1(n584bar)
  );
  //OR U388
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U388 (
    .O(n584),
    .I0(n583),
    .I1(n582)
  );
  //AND U388bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U388bar (
    .O(n584bar),
    .I0(n583bar),
    .I1(n582bar)
  );
  //OR U389
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U389 (
    .O(n582),
    .I0(n581),
    .I1(n580)
  );
  //AND U389bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U389bar (
    .O(n582bar),
    .I0(n581bar),
    .I1(n580bar)
  );
  //OR U390
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U390 (
    .O(n580),
    .I0(in[158]),
    .I1(in[142])
  );
  //AND U390bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U390bar (
    .O(n580bar),
    .I0(inbar[158]),
    .I1(inbar[142])
  );
  //OR U391
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U391 (
    .O(n581),
    .I0(in[175]),
    .I1(in[164])
  );
  //AND U391bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U391bar (
    .O(n581bar),
    .I0(inbar[175]),
    .I1(inbar[164])
  );
  //OR U392
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U392 (
    .O(n583),
    .I0(n579),
    .I1(n578)
  );
  //AND U392bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U392bar (
    .O(n583bar),
    .I0(n579bar),
    .I1(n578bar)
  );
  //OR U393
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U393 (
    .O(n578),
    .I0(in[228]),
    .I1(in[204])
  );
  //AND U393bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U393bar (
    .O(n578bar),
    .I0(inbar[228]),
    .I1(inbar[204])
  );
  //OR U394
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U394 (
    .O(n579),
    .I0(in[91]),
    .I1(in[87])
  );
  //AND U394bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U394bar (
    .O(n579bar),
    .I0(inbar[91]),
    .I1(inbar[87])
  );
  //OR U395
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U395 (
    .O(n585),
    .I0(n577),
    .I1(n576)
  );
  //AND U395bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U395bar (
    .O(n585bar),
    .I0(n577bar),
    .I1(n576bar)
  );
  //OR U396
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U396 (
    .O(n576),
    .I0(n575),
    .I1(n574)
  );
  //AND U396bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U396bar (
    .O(n576bar),
    .I0(n575bar),
    .I1(n574bar)
  );
  //OR U397
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U397 (
    .O(n574),
    .I0(in_21),
    .I1(in_11)
  );
  //AND U397bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U397bar (
    .O(n574bar),
    .I0(in_21bar),
    .I1(in_11bar)
  );
  //OR U398
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U398 (
    .O(n575),
    .I0(in_5),
    .I1(in_3)
  );
  //AND U398bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U398bar (
    .O(n575bar),
    .I0(in_5bar),
    .I1(in_3bar)
  );
  //OR U399
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U399 (
    .O(n577),
    .I0(n573),
    .I1(n572)
  );
  //AND U399bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U399bar (
    .O(n577bar),
    .I0(n573bar),
    .I1(n572bar)
  );
  //OR U400
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U400 (
    .O(n572),
    .I0(in_68),
    .I1(in_64)
  );
  //AND U400bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U400bar (
    .O(n572bar),
    .I0(in_68bar),
    .I1(in_64bar)
  );
  //OR U401
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U401 (
    .O(n573),
    .I0(in_76),
    .I1(in_73)
  );
  //AND U401bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U401bar (
    .O(n573bar),
    .I0(in_76bar),
    .I1(in_73bar)
  );
  //OR U402
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U402 (
    .O(n601),
    .I0(n778),
    .I1(n571)
  );
  //AND U402bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U402bar (
    .O(n601bar),
    .I0(n778bar),
    .I1(n571bar)
  );
  //OR U403
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U403 (
    .O(n571),
    .I0(in[100]),
    .I1(n965)
  );
  //AND U403bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U403bar (
    .O(n571bar),
    .I0(inbar[100]),
    .I1(n965bar)
  );
  //OR U404
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U404 (
    .O(n965),
    .I0(n570),
    .I1(n569)
  );
  //AND U404bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U404bar (
    .O(n965bar),
    .I0(n570bar),
    .I1(n569bar)
  );
  //OR U405
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U405 (
    .O(n569),
    .I0(n568),
    .I1(n567)
  );
  //AND U405bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U405bar (
    .O(n569bar),
    .I0(n568bar),
    .I1(n567bar)
  );
  //OR U406
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U406 (
    .O(n567),
    .I0(n566),
    .I1(n565)
  );
  //AND U406bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U406bar (
    .O(n567bar),
    .I0(n566bar),
    .I1(n565bar)
  );
  //OR U407
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U407 (
    .O(n565),
    .I0(n817),
    .I1(n750)
  );
  //AND U407bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U407bar (
    .O(n565bar),
    .I0(n817bar),
    .I1(n750bar)
  );
  //OR U408
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U408 (
    .O(n750),
    .I0(n564),
    .I1(n563)
  );
  //AND U408bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U408bar (
    .O(n750bar),
    .I0(n564bar),
    .I1(n563bar)
  );
  //OR U409
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U409 (
    .O(n563),
    .I0(n562),
    .I1(n561)
  );
  //AND U409bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U409bar (
    .O(n563bar),
    .I0(n562bar),
    .I1(n561bar)
  );
  //OR U410
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U410 (
    .O(n561),
    .I0(n560),
    .I1(n559)
  );
  //AND U410bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U410bar (
    .O(n561bar),
    .I0(n560bar),
    .I1(n559bar)
  );
  //OR U411
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U411 (
    .O(n559),
    .I0(in[119]),
    .I1(in[103])
  );
  //AND U411bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U411bar (
    .O(n559bar),
    .I0(inbar[119]),
    .I1(inbar[103])
  );
  //OR U412
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U412 (
    .O(n560),
    .I0(in[137]),
    .I1(in[133])
  );
  //AND U412bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U412bar (
    .O(n560bar),
    .I0(inbar[137]),
    .I1(inbar[133])
  );
  //OR U413
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U413 (
    .O(n562),
    .I0(n558),
    .I1(n557)
  );
  //AND U413bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U413bar (
    .O(n562bar),
    .I0(n558bar),
    .I1(n557bar)
  );
  //OR U414
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U414 (
    .O(n557),
    .I0(in[176]),
    .I1(in[173])
  );
  //AND U414bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U414bar (
    .O(n557bar),
    .I0(inbar[176]),
    .I1(inbar[173])
  );
  //OR U415
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U415 (
    .O(n558),
    .I0(in[210]),
    .I1(in[181])
  );
  //AND U415bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U415bar (
    .O(n558bar),
    .I0(inbar[210]),
    .I1(inbar[181])
  );
  //OR U416
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U416 (
    .O(n564),
    .I0(n556),
    .I1(n555)
  );
  //AND U416bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U416bar (
    .O(n564bar),
    .I0(n556bar),
    .I1(n555bar)
  );
  //OR U417
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U417 (
    .O(n555),
    .I0(n554),
    .I1(n553)
  );
  //AND U417bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U417bar (
    .O(n555bar),
    .I0(n554bar),
    .I1(n553bar)
  );
  //OR U418
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U418 (
    .O(n553),
    .I0(in_13),
    .I1(in[234])
  );
  //AND U418bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U418bar (
    .O(n553bar),
    .I0(in_13bar),
    .I1(inbar[234])
  );
  //OR U419
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U419 (
    .O(n554),
    .I0(in_38),
    .I1(in_32)
  );
  //AND U419bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U419bar (
    .O(n554bar),
    .I0(in_38bar),
    .I1(in_32bar)
  );
  //OR U420
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U420 (
    .O(n556),
    .I0(n552),
    .I1(n551)
  );
  //AND U420bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U420bar (
    .O(n556bar),
    .I0(n552bar),
    .I1(n551bar)
  );
  //OR U421
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U421 (
    .O(n551),
    .I0(in_42),
    .I1(in_41)
  );
  //AND U421bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U421bar (
    .O(n551bar),
    .I0(in_42bar),
    .I1(in_41bar)
  );
  //OR U422
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U422 (
    .O(n552),
    .I0(in_7),
    .I1(in_49)
  );
  //AND U422bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U422bar (
    .O(n552bar),
    .I0(in_7bar),
    .I1(in_49bar)
  );
  //OR U423
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U423 (
    .O(n817),
    .I0(n550),
    .I1(n549)
  );
  //AND U423bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U423bar (
    .O(n817bar),
    .I0(n550bar),
    .I1(n549bar)
  );
  //OR U424
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U424 (
    .O(n549),
    .I0(n548),
    .I1(n547)
  );
  //AND U424bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U424bar (
    .O(n549bar),
    .I0(n548bar),
    .I1(n547bar)
  );
  //OR U425
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U425 (
    .O(n547),
    .I0(n546),
    .I1(n545)
  );
  //AND U425bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U425bar (
    .O(n547bar),
    .I0(n546bar),
    .I1(n545bar)
  );
  //OR U426
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U426 (
    .O(n545),
    .I0(in[159]),
    .I1(in[105])
  );
  //AND U426bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U426bar (
    .O(n545bar),
    .I0(inbar[159]),
    .I1(inbar[105])
  );
  //OR U427
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U427 (
    .O(n546),
    .I0(in[206]),
    .I1(in[183])
  );
  //AND U427bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U427bar (
    .O(n546bar),
    .I0(inbar[206]),
    .I1(inbar[183])
  );
  //OR U428
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U428 (
    .O(n548),
    .I0(n544),
    .I1(n543)
  );
  //AND U428bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U428bar (
    .O(n548bar),
    .I0(n544bar),
    .I1(n543bar)
  );
  //OR U429
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U429 (
    .O(n543),
    .I0(in[229]),
    .I1(in[219])
  );
  //AND U429bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U429bar (
    .O(n543bar),
    .I0(inbar[229]),
    .I1(inbar[219])
  );
  //OR U430
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U430 (
    .O(n544),
    .I0(in[235]),
    .I1(in[232])
  );
  //AND U430bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U430bar (
    .O(n544bar),
    .I0(inbar[235]),
    .I1(inbar[232])
  );
  //OR U431
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U431 (
    .O(n550),
    .I0(n542),
    .I1(n541)
  );
  //AND U431bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U431bar (
    .O(n550bar),
    .I0(n542bar),
    .I1(n541bar)
  );
  //OR U432
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U432 (
    .O(n541),
    .I0(n540),
    .I1(n539)
  );
  //AND U432bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U432bar (
    .O(n541bar),
    .I0(n540bar),
    .I1(n539bar)
  );
  //OR U433
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U433 (
    .O(n539),
    .I0(in[249]),
    .I1(in[242])
  );
  //AND U433bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U433bar (
    .O(n539bar),
    .I0(inbar[249]),
    .I1(inbar[242])
  );
  //OR U434
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U434 (
    .O(n540),
    .I0(in[89]),
    .I1(in[254])
  );
  //AND U434bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U434bar (
    .O(n540bar),
    .I0(inbar[89]),
    .I1(inbar[254])
  );
  //OR U435
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U435 (
    .O(n542),
    .I0(n538),
    .I1(n537)
  );
  //AND U435bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U435bar (
    .O(n542bar),
    .I0(n538bar),
    .I1(n537bar)
  );
  //OR U436
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U436 (
    .O(n537),
    .I0(in_14),
    .I1(in[99])
  );
  //AND U436bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U436bar (
    .O(n537bar),
    .I0(in_14bar),
    .I1(inbar[99])
  );
  //OR U437
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U437 (
    .O(n538),
    .I0(in_60),
    .I1(in_18)
  );
  //AND U437bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U437bar (
    .O(n538bar),
    .I0(in_60bar),
    .I1(in_18bar)
  );
  //OR U438
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U438 (
    .O(n566),
    .I0(in[113]),
    .I1(n763)
  );
  //AND U438bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U438bar (
    .O(n566bar),
    .I0(inbar[113]),
    .I1(n763bar)
  );
  //OR U439
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U439 (
    .O(n763),
    .I0(n536),
    .I1(n535)
  );
  //AND U439bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U439bar (
    .O(n763bar),
    .I0(n536bar),
    .I1(n535bar)
  );
  //OR U440
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U440 (
    .O(n535),
    .I0(n534),
    .I1(n533)
  );
  //AND U440bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U440bar (
    .O(n535bar),
    .I0(n534bar),
    .I1(n533bar)
  );
  //OR U441
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U441 (
    .O(n533),
    .I0(n532),
    .I1(n531)
  );
  //AND U441bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U441bar (
    .O(n533bar),
    .I0(n532bar),
    .I1(n531bar)
  );
  //OR U442
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U442 (
    .O(n531),
    .I0(in[115]),
    .I1(in[110])
  );
  //AND U442bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U442bar (
    .O(n531bar),
    .I0(inbar[115]),
    .I1(inbar[110])
  );
  //OR U443
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U443 (
    .O(n532),
    .I0(in[125]),
    .I1(in[117])
  );
  //AND U443bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U443bar (
    .O(n532bar),
    .I0(inbar[125]),
    .I1(inbar[117])
  );
  //OR U444
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U444 (
    .O(n534),
    .I0(n530),
    .I1(n529)
  );
  //AND U444bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U444bar (
    .O(n534bar),
    .I0(n530bar),
    .I1(n529bar)
  );
  //OR U445
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U445 (
    .O(n529),
    .I0(in[180]),
    .I1(in[128])
  );
  //AND U445bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U445bar (
    .O(n529bar),
    .I0(inbar[180]),
    .I1(inbar[128])
  );
  //OR U446
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U446 (
    .O(n530),
    .I0(in[205]),
    .I1(in[201])
  );
  //AND U446bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U446bar (
    .O(n530bar),
    .I0(inbar[205]),
    .I1(inbar[201])
  );
  //OR U447
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U447 (
    .O(n536),
    .I0(n528),
    .I1(n527)
  );
  //AND U447bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U447bar (
    .O(n536bar),
    .I0(n528bar),
    .I1(n527bar)
  );
  //OR U448
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U448 (
    .O(n527),
    .I0(n526),
    .I1(n525)
  );
  //AND U448bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U448bar (
    .O(n527bar),
    .I0(n526bar),
    .I1(n525bar)
  );
  //OR U449
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U449 (
    .O(n525),
    .I0(in[244]),
    .I1(in[239])
  );
  //AND U449bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U449bar (
    .O(n525bar),
    .I0(inbar[244]),
    .I1(inbar[239])
  );
  //OR U450
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U450 (
    .O(n526),
    .I0(in[95]),
    .I1(in[83])
  );
  //AND U450bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U450bar (
    .O(n526bar),
    .I0(inbar[95]),
    .I1(inbar[83])
  );
  //OR U451
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U451 (
    .O(n528),
    .I0(n524),
    .I1(n523)
  );
  //AND U451bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U451bar (
    .O(n528bar),
    .I0(n524bar),
    .I1(n523bar)
  );
  //OR U452
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U452 (
    .O(n523),
    .I0(in_24),
    .I1(in[97])
  );
  //AND U452bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U452bar (
    .O(n523bar),
    .I0(in_24bar),
    .I1(inbar[97])
  );
  //OR U453
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U453 (
    .O(n524),
    .I0(in_33),
    .I1(in_27)
  );
  //AND U453bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U453bar (
    .O(n524bar),
    .I0(in_33bar),
    .I1(in_27bar)
  );
  //OR U454
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U454 (
    .O(n568),
    .I0(n522),
    .I1(n521)
  );
  //AND U454bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U454bar (
    .O(n568bar),
    .I0(n522bar),
    .I1(n521bar)
  );
  //OR U455
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U455 (
    .O(n521),
    .I0(in[145]),
    .I1(in[126])
  );
  //AND U455bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U455bar (
    .O(n521bar),
    .I0(inbar[145]),
    .I1(inbar[126])
  );
  //OR U456
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U456 (
    .O(n522),
    .I0(in[169]),
    .I1(n520)
  );
  //AND U456bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U456bar (
    .O(n522bar),
    .I0(inbar[169]),
    .I1(n520bar)
  );
  //OR U457
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U457 (
    .O(n520),
    .I0(in[221]),
    .I1(in[172])
  );
  //AND U457bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U457bar (
    .O(n520bar),
    .I0(inbar[221]),
    .I1(inbar[172])
  );
  //OR U458
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U458 (
    .O(n570),
    .I0(n519),
    .I1(n518)
  );
  //AND U458bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U458bar (
    .O(n570bar),
    .I0(n519bar),
    .I1(n518bar)
  );
  //OR U459
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U459 (
    .O(n518),
    .I0(n517),
    .I1(n516)
  );
  //AND U459bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U459bar (
    .O(n518bar),
    .I0(n517bar),
    .I1(n516bar)
  );
  //OR U460
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U460 (
    .O(n516),
    .I0(in[241]),
    .I1(in[224])
  );
  //AND U460bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U460bar (
    .O(n516bar),
    .I0(inbar[241]),
    .I1(inbar[224])
  );
  //OR U461
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U461 (
    .O(n517),
    .I0(in[86]),
    .I1(n515)
  );
  //AND U461bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U461bar (
    .O(n517bar),
    .I0(inbar[86]),
    .I1(n515bar)
  );
  //OR U462
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U462 (
    .O(n515),
    .I0(in_43),
    .I1(in_34)
  );
  //AND U462bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U462bar (
    .O(n515bar),
    .I0(in_43bar),
    .I1(in_34bar)
  );
  //OR U463
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U463 (
    .O(n519),
    .I0(n514),
    .I1(n513)
  );
  //AND U463bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U463bar (
    .O(n519bar),
    .I0(n514bar),
    .I1(n513bar)
  );
  //OR U464
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U464 (
    .O(n513),
    .I0(in_65),
    .I1(in_51)
  );
  //AND U464bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U464bar (
    .O(n513bar),
    .I0(in_65bar),
    .I1(in_51bar)
  );
  //OR U465
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U465 (
    .O(n514),
    .I0(in_75),
    .I1(n512)
  );
  //AND U465bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U465bar (
    .O(n514bar),
    .I0(in_75bar),
    .I1(n512bar)
  );
  //OR U466
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U466 (
    .O(n512),
    .I0(in_81),
    .I1(in_77)
  );
  //AND U466bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U466bar (
    .O(n512bar),
    .I0(in_81bar),
    .I1(in_77bar)
  );
  //OR U467
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U467 (
    .O(n778),
    .I0(n511),
    .I1(n510)
  );
  //AND U467bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U467bar (
    .O(n778bar),
    .I0(n511bar),
    .I1(n510bar)
  );
  //OR U468
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U468 (
    .O(n510),
    .I0(n509),
    .I1(n508)
  );
  //AND U468bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U468bar (
    .O(n510bar),
    .I0(n509bar),
    .I1(n508bar)
  );
  //OR U469
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U469 (
    .O(n508),
    .I0(n507),
    .I1(n506)
  );
  //AND U469bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U469bar (
    .O(n508bar),
    .I0(n507bar),
    .I1(n506bar)
  );
  //OR U470
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U470 (
    .O(n506),
    .I0(in[107]),
    .I1(in[101])
  );
  //AND U470bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U470bar (
    .O(n506bar),
    .I0(inbar[107]),
    .I1(inbar[101])
  );
  //OR U471
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U471 (
    .O(n507),
    .I0(in[139]),
    .I1(in[132])
  );
  //AND U471bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U471bar (
    .O(n507bar),
    .I0(inbar[139]),
    .I1(inbar[132])
  );
  //OR U472
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U472 (
    .O(n509),
    .I0(n505),
    .I1(n504)
  );
  //AND U472bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U472bar (
    .O(n509bar),
    .I0(n505bar),
    .I1(n504bar)
  );
  //OR U473
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U473 (
    .O(n504),
    .I0(in[146]),
    .I1(in[141])
  );
  //AND U473bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U473bar (
    .O(n504bar),
    .I0(inbar[146]),
    .I1(inbar[141])
  );
  //OR U474
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U474 (
    .O(n505),
    .I0(in[203]),
    .I1(in[179])
  );
  //AND U474bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U474bar (
    .O(n505bar),
    .I0(inbar[203]),
    .I1(inbar[179])
  );
  //OR U475
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U475 (
    .O(n511),
    .I0(n503),
    .I1(n502)
  );
  //AND U475bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U475bar (
    .O(n511bar),
    .I0(n503bar),
    .I1(n502bar)
  );
  //OR U476
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U476 (
    .O(n502),
    .I0(n501),
    .I1(n500)
  );
  //AND U476bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U476bar (
    .O(n502bar),
    .I0(n501bar),
    .I1(n500bar)
  );
  //OR U477
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U477 (
    .O(n500),
    .I0(in[243]),
    .I1(in[222])
  );
  //AND U477bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U477bar (
    .O(n500bar),
    .I0(inbar[243]),
    .I1(inbar[222])
  );
  //OR U478
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U478 (
    .O(n501),
    .I0(in[251]),
    .I1(in[250])
  );
  //AND U478bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U478bar (
    .O(n501bar),
    .I0(inbar[251]),
    .I1(inbar[250])
  );
  //OR U479
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U479 (
    .O(n503),
    .I0(n499),
    .I1(n498)
  );
  //AND U479bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U479bar (
    .O(n503bar),
    .I0(n499bar),
    .I1(n498bar)
  );
  //OR U480
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U480 (
    .O(n498),
    .I0(in_37),
    .I1(in_19)
  );
  //AND U480bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U480bar (
    .O(n498bar),
    .I0(in_37bar),
    .I1(in_19bar)
  );
  //OR U481
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U481 (
    .O(n499),
    .I0(in_78),
    .I1(in_6)
  );
  //AND U481bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U481bar (
    .O(n499bar),
    .I0(in_78bar),
    .I1(in_6bar)
  );
  //OR U482
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U482 (
    .O(n603),
    .I0(n497),
    .I1(n496)
  );
  //AND U482bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U482bar (
    .O(n603bar),
    .I0(n497bar),
    .I1(n496bar)
  );
  //OR U483
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U483 (
    .O(n496),
    .I0(in[112]),
    .I1(in[102])
  );
  //AND U483bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U483bar (
    .O(n496bar),
    .I0(inbar[112]),
    .I1(inbar[102])
  );
  //OR U484
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U484 (
    .O(n497),
    .I0(in[123]),
    .I1(n495)
  );
  //AND U484bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U484bar (
    .O(n497bar),
    .I0(inbar[123]),
    .I1(n495bar)
  );
  //OR U485
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U485 (
    .O(n495),
    .I0(in[143]),
    .I1(in[130])
  );
  //AND U485bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U485bar (
    .O(n495bar),
    .I0(inbar[143]),
    .I1(inbar[130])
  );
  //OR U486
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U486 (
    .O(n605),
    .I0(n494),
    .I1(n493)
  );
  //AND U486bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U486bar (
    .O(n605bar),
    .I0(n494bar),
    .I1(n493bar)
  );
  //OR U487
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U487 (
    .O(n493),
    .I0(n492),
    .I1(n491)
  );
  //AND U487bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U487bar (
    .O(n493bar),
    .I0(n492bar),
    .I1(n491bar)
  );
  //OR U488
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U488 (
    .O(n491),
    .I0(in[216]),
    .I1(in[213])
  );
  //AND U488bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U488bar (
    .O(n491bar),
    .I0(inbar[216]),
    .I1(inbar[213])
  );
  //OR U489
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U489 (
    .O(n492),
    .I0(in[227]),
    .I1(n490)
  );
  //AND U489bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U489bar (
    .O(n492bar),
    .I0(inbar[227]),
    .I1(n490bar)
  );
  //OR U490
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U490 (
    .O(n490),
    .I0(in_0),
    .I1(in[248])
  );
  //AND U490bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U490bar (
    .O(n490bar),
    .I0(in_0bar),
    .I1(inbar[248])
  );
  //OR U491
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U491 (
    .O(n494),
    .I0(n489),
    .I1(n488)
  );
  //AND U491bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U491bar (
    .O(n494bar),
    .I0(n489bar),
    .I1(n488bar)
  );
  //OR U492
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U492 (
    .O(n488),
    .I0(in_46),
    .I1(in_44)
  );
  //AND U492bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U492bar (
    .O(n488bar),
    .I0(in_46bar),
    .I1(in_44bar)
  );
  //OR U493
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U493 (
    .O(n489),
    .I0(in_50),
    .I1(n487)
  );
  //AND U493bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U493bar (
    .O(n489bar),
    .I0(in_50bar),
    .I1(n487bar)
  );
  //OR U494
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U494 (
    .O(n487),
    .I0(in_9),
    .I1(in_80)
  );
  //AND U494bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U494bar (
    .O(n487bar),
    .I0(in_9bar),
    .I1(in_80bar)
  );
endmodule

module sBox_5 ( in, out );

  input wire [7:0] in;
//input_done

  output wire [7:0] out;
//output_done

  wire [255:0] decodeOut;
//wire_done

  decode_5 dec ( .in(in), .out(decodeOut) );
  encode_5 enc ( .in(decodeOut), .out(out) );
endmodule

module CD2_21 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD2_22 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD2_23 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD2_24 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD4_11 ( a, b, y );

  input wire [3:0] a;
  input wire [3:0] b;
  wire [3:0] abar;
  wire [3:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
//input_done

  output wire [15:0] y;
  wire [15:0] ybar;
//output_done

//wire_done

  //AND U1
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1 (
    .O(y[9]),
    .I0(b[1]),
    .I1(a[2])
  );
  //OR U1bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1bar (
    .O(ybar[9]),
    .I0(bbar[1]),
    .I1(abar[2])
  );
  //AND U2
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2 (
    .O(y[8]),
    .I0(b[0]),
    .I1(a[2])
  );
  //OR U2bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2bar (
    .O(ybar[8]),
    .I0(bbar[0]),
    .I1(abar[2])
  );
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[7]),
    .I0(b[3]),
    .I1(a[1])
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[7]),
    .I0(bbar[3]),
    .I1(abar[1])
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[6]),
    .I0(b[2]),
    .I1(a[1])
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[6]),
    .I0(bbar[2]),
    .I1(abar[1])
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[5]),
    .I0(a[1]),
    .I1(b[1])
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[5]),
    .I0(abar[1]),
    .I1(bbar[1])
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[4]),
    .I0(a[1]),
    .I1(b[0])
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[4]),
    .I0(abar[1]),
    .I1(bbar[0])
  );
  //AND U7
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7 (
    .O(y[3]),
    .I0(a[0]),
    .I1(b[3])
  );
  //OR U7bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7bar (
    .O(ybar[3]),
    .I0(abar[0]),
    .I1(bbar[3])
  );
  //AND U8
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8 (
    .O(y[2]),
    .I0(a[0]),
    .I1(b[2])
  );
  //OR U8bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8bar (
    .O(ybar[2]),
    .I0(abar[0]),
    .I1(bbar[2])
  );
  //AND U9
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9 (
    .O(y[1]),
    .I0(a[0]),
    .I1(b[1])
  );
  //OR U9bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9bar (
    .O(ybar[1]),
    .I0(abar[0]),
    .I1(bbar[1])
  );
  //AND U10
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10 (
    .O(y[15]),
    .I0(a[3]),
    .I1(b[3])
  );
  //OR U10bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10bar (
    .O(ybar[15]),
    .I0(abar[3]),
    .I1(bbar[3])
  );
  //AND U11
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11 (
    .O(y[14]),
    .I0(a[3]),
    .I1(b[2])
  );
  //OR U11bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11bar (
    .O(ybar[14]),
    .I0(abar[3]),
    .I1(bbar[2])
  );
  //AND U12
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12 (
    .O(y[13]),
    .I0(a[3]),
    .I1(b[1])
  );
  //OR U12bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12bar (
    .O(ybar[13]),
    .I0(abar[3]),
    .I1(bbar[1])
  );
  //AND U13
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13 (
    .O(y[12]),
    .I0(a[3]),
    .I1(b[0])
  );
  //OR U13bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13bar (
    .O(ybar[12]),
    .I0(abar[3]),
    .I1(bbar[0])
  );
  //AND U14
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14 (
    .O(y[11]),
    .I0(b[3]),
    .I1(a[2])
  );
  //OR U14bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14bar (
    .O(ybar[11]),
    .I0(bbar[3]),
    .I1(abar[2])
  );
  //AND U15
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15 (
    .O(y[10]),
    .I0(b[2]),
    .I1(a[2])
  );
  //OR U15bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15bar (
    .O(ybar[10]),
    .I0(bbar[2]),
    .I1(abar[2])
  );
  //AND U16
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16 (
    .O(y[0]),
    .I0(a[0]),
    .I1(b[0])
  );
  //OR U16bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16bar (
    .O(ybar[0]),
    .I0(abar[0]),
    .I1(bbar[0])
  );
endmodule

module CD4_12 ( a, b, y );

  input wire [3:0] a;
  input wire [3:0] b;
  wire [3:0] abar;
  wire [3:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
//input_done

  output wire [15:0] y;
  wire [15:0] ybar;
//output_done

//wire_done

  //AND U1
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1 (
    .O(y[9]),
    .I0(b[1]),
    .I1(a[2])
  );
  //OR U1bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1bar (
    .O(ybar[9]),
    .I0(bbar[1]),
    .I1(abar[2])
  );
  //AND U2
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2 (
    .O(y[8]),
    .I0(b[0]),
    .I1(a[2])
  );
  //OR U2bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2bar (
    .O(ybar[8]),
    .I0(bbar[0]),
    .I1(abar[2])
  );
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[7]),
    .I0(b[3]),
    .I1(a[1])
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[7]),
    .I0(bbar[3]),
    .I1(abar[1])
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[6]),
    .I0(b[2]),
    .I1(a[1])
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[6]),
    .I0(bbar[2]),
    .I1(abar[1])
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[5]),
    .I0(a[1]),
    .I1(b[1])
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[5]),
    .I0(abar[1]),
    .I1(bbar[1])
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[4]),
    .I0(a[1]),
    .I1(b[0])
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[4]),
    .I0(abar[1]),
    .I1(bbar[0])
  );
  //AND U7
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7 (
    .O(y[3]),
    .I0(a[0]),
    .I1(b[3])
  );
  //OR U7bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7bar (
    .O(ybar[3]),
    .I0(abar[0]),
    .I1(bbar[3])
  );
  //AND U8
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8 (
    .O(y[2]),
    .I0(a[0]),
    .I1(b[2])
  );
  //OR U8bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8bar (
    .O(ybar[2]),
    .I0(abar[0]),
    .I1(bbar[2])
  );
  //AND U9
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9 (
    .O(y[1]),
    .I0(a[0]),
    .I1(b[1])
  );
  //OR U9bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9bar (
    .O(ybar[1]),
    .I0(abar[0]),
    .I1(bbar[1])
  );
  //AND U10
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10 (
    .O(y[15]),
    .I0(a[3]),
    .I1(b[3])
  );
  //OR U10bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10bar (
    .O(ybar[15]),
    .I0(abar[3]),
    .I1(bbar[3])
  );
  //AND U11
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11 (
    .O(y[14]),
    .I0(a[3]),
    .I1(b[2])
  );
  //OR U11bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11bar (
    .O(ybar[14]),
    .I0(abar[3]),
    .I1(bbar[2])
  );
  //AND U12
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12 (
    .O(y[13]),
    .I0(a[3]),
    .I1(b[1])
  );
  //OR U12bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12bar (
    .O(ybar[13]),
    .I0(abar[3]),
    .I1(bbar[1])
  );
  //AND U13
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13 (
    .O(y[12]),
    .I0(a[3]),
    .I1(b[0])
  );
  //OR U13bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13bar (
    .O(ybar[12]),
    .I0(abar[3]),
    .I1(bbar[0])
  );
  //AND U14
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14 (
    .O(y[11]),
    .I0(b[3]),
    .I1(a[2])
  );
  //OR U14bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14bar (
    .O(ybar[11]),
    .I0(bbar[3]),
    .I1(abar[2])
  );
  //AND U15
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15 (
    .O(y[10]),
    .I0(b[2]),
    .I1(a[2])
  );
  //OR U15bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15bar (
    .O(ybar[10]),
    .I0(bbar[2]),
    .I1(abar[2])
  );
  //AND U16
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16 (
    .O(y[0]),
    .I0(a[0]),
    .I1(b[0])
  );
  //OR U16bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16bar (
    .O(ybar[0]),
    .I0(abar[0]),
    .I1(bbar[0])
  );
endmodule

module CD16_6 ( a, b, y );

  input wire [15:0] a;
  input wire [15:0] b;
  wire [15:0] abar;
  wire [15:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign abar[8] = ~a[8];
  assign abar[9] = ~a[9];
  assign abar[10] = ~a[10];
  assign abar[11] = ~a[11];
  assign abar[12] = ~a[12];
  assign abar[13] = ~a[13];
  assign abar[14] = ~a[14];
  assign abar[15] = ~a[15];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign bbar[8] = ~b[8];
  assign bbar[9] = ~b[9];
  assign bbar[10] = ~b[10];
  assign bbar[11] = ~b[11];
  assign bbar[12] = ~b[12];
  assign bbar[13] = ~b[13];
  assign bbar[14] = ~b[14];
  assign bbar[15] = ~b[15];
//input_done

  output wire [255:0] y;
  wire [255:0] ybar;
//output_done

//wire_done

  //AND U1
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1 (
    .O(y[9]),
    .I0(b[9]),
    .I1(a[0])
  );
  //OR U1bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1bar (
    .O(ybar[9]),
    .I0(bbar[9]),
    .I1(abar[0])
  );
  //AND U2
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2 (
    .O(y[99]),
    .I0(b[3]),
    .I1(a[6])
  );
  //OR U2bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2bar (
    .O(ybar[99]),
    .I0(bbar[3]),
    .I1(abar[6])
  );
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[98]),
    .I0(b[2]),
    .I1(a[6])
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[98]),
    .I0(bbar[2]),
    .I1(abar[6])
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[97]),
    .I0(b[1]),
    .I1(a[6])
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[97]),
    .I0(bbar[1]),
    .I1(abar[6])
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[96]),
    .I0(b[0]),
    .I1(a[6])
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[96]),
    .I0(bbar[0]),
    .I1(abar[6])
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[95]),
    .I0(b[15]),
    .I1(a[5])
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[95]),
    .I0(bbar[15]),
    .I1(abar[5])
  );
  //AND U7
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7 (
    .O(y[94]),
    .I0(b[14]),
    .I1(a[5])
  );
  //OR U7bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7bar (
    .O(ybar[94]),
    .I0(bbar[14]),
    .I1(abar[5])
  );
  //AND U8
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8 (
    .O(y[93]),
    .I0(b[13]),
    .I1(a[5])
  );
  //OR U8bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8bar (
    .O(ybar[93]),
    .I0(bbar[13]),
    .I1(abar[5])
  );
  //AND U9
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9 (
    .O(y[92]),
    .I0(b[12]),
    .I1(a[5])
  );
  //OR U9bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9bar (
    .O(ybar[92]),
    .I0(bbar[12]),
    .I1(abar[5])
  );
  //AND U10
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10 (
    .O(y[91]),
    .I0(b[11]),
    .I1(a[5])
  );
  //OR U10bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10bar (
    .O(ybar[91]),
    .I0(bbar[11]),
    .I1(abar[5])
  );
  //AND U11
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11 (
    .O(y[90]),
    .I0(b[10]),
    .I1(a[5])
  );
  //OR U11bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11bar (
    .O(ybar[90]),
    .I0(bbar[10]),
    .I1(abar[5])
  );
  //AND U12
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12 (
    .O(y[8]),
    .I0(b[8]),
    .I1(a[0])
  );
  //OR U12bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12bar (
    .O(ybar[8]),
    .I0(bbar[8]),
    .I1(abar[0])
  );
  //AND U13
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13 (
    .O(y[89]),
    .I0(a[5]),
    .I1(b[9])
  );
  //OR U13bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13bar (
    .O(ybar[89]),
    .I0(abar[5]),
    .I1(bbar[9])
  );
  //AND U14
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14 (
    .O(y[88]),
    .I0(b[8]),
    .I1(a[5])
  );
  //OR U14bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14bar (
    .O(ybar[88]),
    .I0(bbar[8]),
    .I1(abar[5])
  );
  //AND U15
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15 (
    .O(y[87]),
    .I0(b[7]),
    .I1(a[5])
  );
  //OR U15bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15bar (
    .O(ybar[87]),
    .I0(bbar[7]),
    .I1(abar[5])
  );
  //AND U16
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16 (
    .O(y[86]),
    .I0(b[6]),
    .I1(a[5])
  );
  //OR U16bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16bar (
    .O(ybar[86]),
    .I0(bbar[6]),
    .I1(abar[5])
  );
  //AND U17
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U17 (
    .O(y[85]),
    .I0(b[5]),
    .I1(a[5])
  );
  //OR U17bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U17bar (
    .O(ybar[85]),
    .I0(bbar[5]),
    .I1(abar[5])
  );
  //AND U18
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U18 (
    .O(y[84]),
    .I0(b[4]),
    .I1(a[5])
  );
  //OR U18bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U18bar (
    .O(ybar[84]),
    .I0(bbar[4]),
    .I1(abar[5])
  );
  //AND U19
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U19 (
    .O(y[83]),
    .I0(a[5]),
    .I1(b[3])
  );
  //OR U19bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U19bar (
    .O(ybar[83]),
    .I0(abar[5]),
    .I1(bbar[3])
  );
  //AND U20
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U20 (
    .O(y[82]),
    .I0(a[5]),
    .I1(b[2])
  );
  //OR U20bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U20bar (
    .O(ybar[82]),
    .I0(abar[5]),
    .I1(bbar[2])
  );
  //AND U21
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U21 (
    .O(y[81]),
    .I0(a[5]),
    .I1(b[1])
  );
  //OR U21bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U21bar (
    .O(ybar[81]),
    .I0(abar[5]),
    .I1(bbar[1])
  );
  //AND U22
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U22 (
    .O(y[80]),
    .I0(a[5]),
    .I1(b[0])
  );
  //OR U22bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U22bar (
    .O(ybar[80]),
    .I0(abar[5]),
    .I1(bbar[0])
  );
  //AND U23
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U23 (
    .O(y[7]),
    .I0(b[7]),
    .I1(a[0])
  );
  //OR U23bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U23bar (
    .O(ybar[7]),
    .I0(bbar[7]),
    .I1(abar[0])
  );
  //AND U24
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U24 (
    .O(y[79]),
    .I0(a[4]),
    .I1(b[15])
  );
  //OR U24bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U24bar (
    .O(ybar[79]),
    .I0(abar[4]),
    .I1(bbar[15])
  );
  //AND U25
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U25 (
    .O(y[78]),
    .I0(a[4]),
    .I1(b[14])
  );
  //OR U25bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U25bar (
    .O(ybar[78]),
    .I0(abar[4]),
    .I1(bbar[14])
  );
  //AND U26
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U26 (
    .O(y[77]),
    .I0(a[4]),
    .I1(b[13])
  );
  //OR U26bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U26bar (
    .O(ybar[77]),
    .I0(abar[4]),
    .I1(bbar[13])
  );
  //AND U27
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U27 (
    .O(y[76]),
    .I0(a[4]),
    .I1(b[12])
  );
  //OR U27bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U27bar (
    .O(ybar[76]),
    .I0(abar[4]),
    .I1(bbar[12])
  );
  //AND U28
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U28 (
    .O(y[75]),
    .I0(a[4]),
    .I1(b[11])
  );
  //OR U28bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U28bar (
    .O(ybar[75]),
    .I0(abar[4]),
    .I1(bbar[11])
  );
  //AND U29
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U29 (
    .O(y[74]),
    .I0(a[4]),
    .I1(b[10])
  );
  //OR U29bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U29bar (
    .O(ybar[74]),
    .I0(abar[4]),
    .I1(bbar[10])
  );
  //AND U30
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U30 (
    .O(y[73]),
    .I0(a[4]),
    .I1(b[9])
  );
  //OR U30bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U30bar (
    .O(ybar[73]),
    .I0(abar[4]),
    .I1(bbar[9])
  );
  //AND U31
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U31 (
    .O(y[72]),
    .I0(a[4]),
    .I1(b[8])
  );
  //OR U31bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U31bar (
    .O(ybar[72]),
    .I0(abar[4]),
    .I1(bbar[8])
  );
  //AND U32
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U32 (
    .O(y[71]),
    .I0(a[4]),
    .I1(b[7])
  );
  //OR U32bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U32bar (
    .O(ybar[71]),
    .I0(abar[4]),
    .I1(bbar[7])
  );
  //AND U33
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U33 (
    .O(y[70]),
    .I0(a[4]),
    .I1(b[6])
  );
  //OR U33bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U33bar (
    .O(ybar[70]),
    .I0(abar[4]),
    .I1(bbar[6])
  );
  //AND U34
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U34 (
    .O(y[6]),
    .I0(b[6]),
    .I1(a[0])
  );
  //OR U34bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U34bar (
    .O(ybar[6]),
    .I0(bbar[6]),
    .I1(abar[0])
  );
  //AND U35
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U35 (
    .O(y[69]),
    .I0(a[4]),
    .I1(b[5])
  );
  //OR U35bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U35bar (
    .O(ybar[69]),
    .I0(abar[4]),
    .I1(bbar[5])
  );
  //AND U36
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U36 (
    .O(y[68]),
    .I0(a[4]),
    .I1(b[4])
  );
  //OR U36bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U36bar (
    .O(ybar[68]),
    .I0(abar[4]),
    .I1(bbar[4])
  );
  //AND U37
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U37 (
    .O(y[67]),
    .I0(a[4]),
    .I1(b[3])
  );
  //OR U37bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U37bar (
    .O(ybar[67]),
    .I0(abar[4]),
    .I1(bbar[3])
  );
  //AND U38
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U38 (
    .O(y[66]),
    .I0(a[4]),
    .I1(b[2])
  );
  //OR U38bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U38bar (
    .O(ybar[66]),
    .I0(abar[4]),
    .I1(bbar[2])
  );
  //AND U39
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U39 (
    .O(y[65]),
    .I0(a[4]),
    .I1(b[1])
  );
  //OR U39bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U39bar (
    .O(ybar[65]),
    .I0(abar[4]),
    .I1(bbar[1])
  );
  //AND U40
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U40 (
    .O(y[64]),
    .I0(a[4]),
    .I1(b[0])
  );
  //OR U40bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U40bar (
    .O(ybar[64]),
    .I0(abar[4]),
    .I1(bbar[0])
  );
  //AND U41
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U41 (
    .O(y[63]),
    .I0(a[3]),
    .I1(b[15])
  );
  //OR U41bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U41bar (
    .O(ybar[63]),
    .I0(abar[3]),
    .I1(bbar[15])
  );
  //AND U42
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U42 (
    .O(y[62]),
    .I0(a[3]),
    .I1(b[14])
  );
  //OR U42bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U42bar (
    .O(ybar[62]),
    .I0(abar[3]),
    .I1(bbar[14])
  );
  //AND U43
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U43 (
    .O(y[61]),
    .I0(a[3]),
    .I1(b[13])
  );
  //OR U43bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U43bar (
    .O(ybar[61]),
    .I0(abar[3]),
    .I1(bbar[13])
  );
  //AND U44
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U44 (
    .O(y[60]),
    .I0(a[3]),
    .I1(b[12])
  );
  //OR U44bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U44bar (
    .O(ybar[60]),
    .I0(abar[3]),
    .I1(bbar[12])
  );
  //AND U45
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U45 (
    .O(y[5]),
    .I0(b[5]),
    .I1(a[0])
  );
  //OR U45bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U45bar (
    .O(ybar[5]),
    .I0(bbar[5]),
    .I1(abar[0])
  );
  //AND U46
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U46 (
    .O(y[59]),
    .I0(a[3]),
    .I1(b[11])
  );
  //OR U46bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U46bar (
    .O(ybar[59]),
    .I0(abar[3]),
    .I1(bbar[11])
  );
  //AND U47
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U47 (
    .O(y[58]),
    .I0(a[3]),
    .I1(b[10])
  );
  //OR U47bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U47bar (
    .O(ybar[58]),
    .I0(abar[3]),
    .I1(bbar[10])
  );
  //AND U48
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U48 (
    .O(y[57]),
    .I0(a[3]),
    .I1(b[9])
  );
  //OR U48bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U48bar (
    .O(ybar[57]),
    .I0(abar[3]),
    .I1(bbar[9])
  );
  //AND U49
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U49 (
    .O(y[56]),
    .I0(a[3]),
    .I1(b[8])
  );
  //OR U49bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U49bar (
    .O(ybar[56]),
    .I0(abar[3]),
    .I1(bbar[8])
  );
  //AND U50
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U50 (
    .O(y[55]),
    .I0(a[3]),
    .I1(b[7])
  );
  //OR U50bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U50bar (
    .O(ybar[55]),
    .I0(abar[3]),
    .I1(bbar[7])
  );
  //AND U51
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U51 (
    .O(y[54]),
    .I0(a[3]),
    .I1(b[6])
  );
  //OR U51bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U51bar (
    .O(ybar[54]),
    .I0(abar[3]),
    .I1(bbar[6])
  );
  //AND U52
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U52 (
    .O(y[53]),
    .I0(a[3]),
    .I1(b[5])
  );
  //OR U52bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U52bar (
    .O(ybar[53]),
    .I0(abar[3]),
    .I1(bbar[5])
  );
  //AND U53
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U53 (
    .O(y[52]),
    .I0(a[3]),
    .I1(b[4])
  );
  //OR U53bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U53bar (
    .O(ybar[52]),
    .I0(abar[3]),
    .I1(bbar[4])
  );
  //AND U54
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U54 (
    .O(y[51]),
    .I0(a[3]),
    .I1(b[3])
  );
  //OR U54bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U54bar (
    .O(ybar[51]),
    .I0(abar[3]),
    .I1(bbar[3])
  );
  //AND U55
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U55 (
    .O(y[50]),
    .I0(a[3]),
    .I1(b[2])
  );
  //OR U55bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U55bar (
    .O(ybar[50]),
    .I0(abar[3]),
    .I1(bbar[2])
  );
  //AND U56
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U56 (
    .O(y[4]),
    .I0(b[4]),
    .I1(a[0])
  );
  //OR U56bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U56bar (
    .O(ybar[4]),
    .I0(bbar[4]),
    .I1(abar[0])
  );
  //AND U57
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U57 (
    .O(y[49]),
    .I0(a[3]),
    .I1(b[1])
  );
  //OR U57bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U57bar (
    .O(ybar[49]),
    .I0(abar[3]),
    .I1(bbar[1])
  );
  //AND U58
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U58 (
    .O(y[48]),
    .I0(a[3]),
    .I1(b[0])
  );
  //OR U58bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U58bar (
    .O(ybar[48]),
    .I0(abar[3]),
    .I1(bbar[0])
  );
  //AND U59
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U59 (
    .O(y[47]),
    .I0(a[2]),
    .I1(b[15])
  );
  //OR U59bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U59bar (
    .O(ybar[47]),
    .I0(abar[2]),
    .I1(bbar[15])
  );
  //AND U60
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U60 (
    .O(y[46]),
    .I0(a[2]),
    .I1(b[14])
  );
  //OR U60bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U60bar (
    .O(ybar[46]),
    .I0(abar[2]),
    .I1(bbar[14])
  );
  //AND U61
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U61 (
    .O(y[45]),
    .I0(a[2]),
    .I1(b[13])
  );
  //OR U61bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U61bar (
    .O(ybar[45]),
    .I0(abar[2]),
    .I1(bbar[13])
  );
  //AND U62
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U62 (
    .O(y[44]),
    .I0(a[2]),
    .I1(b[12])
  );
  //OR U62bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U62bar (
    .O(ybar[44]),
    .I0(abar[2]),
    .I1(bbar[12])
  );
  //AND U63
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U63 (
    .O(y[43]),
    .I0(a[2]),
    .I1(b[11])
  );
  //OR U63bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U63bar (
    .O(ybar[43]),
    .I0(abar[2]),
    .I1(bbar[11])
  );
  //AND U64
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U64 (
    .O(y[42]),
    .I0(a[2]),
    .I1(b[10])
  );
  //OR U64bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U64bar (
    .O(ybar[42]),
    .I0(abar[2]),
    .I1(bbar[10])
  );
  //AND U65
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U65 (
    .O(y[41]),
    .I0(a[2]),
    .I1(b[9])
  );
  //OR U65bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U65bar (
    .O(ybar[41]),
    .I0(abar[2]),
    .I1(bbar[9])
  );
  //AND U66
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U66 (
    .O(y[40]),
    .I0(a[2]),
    .I1(b[8])
  );
  //OR U66bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U66bar (
    .O(ybar[40]),
    .I0(abar[2]),
    .I1(bbar[8])
  );
  //AND U67
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U67 (
    .O(y[3]),
    .I0(b[3]),
    .I1(a[0])
  );
  //OR U67bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U67bar (
    .O(ybar[3]),
    .I0(bbar[3]),
    .I1(abar[0])
  );
  //AND U68
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U68 (
    .O(y[39]),
    .I0(a[2]),
    .I1(b[7])
  );
  //OR U68bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U68bar (
    .O(ybar[39]),
    .I0(abar[2]),
    .I1(bbar[7])
  );
  //AND U69
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U69 (
    .O(y[38]),
    .I0(a[2]),
    .I1(b[6])
  );
  //OR U69bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U69bar (
    .O(ybar[38]),
    .I0(abar[2]),
    .I1(bbar[6])
  );
  //AND U70
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U70 (
    .O(y[37]),
    .I0(a[2]),
    .I1(b[5])
  );
  //OR U70bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U70bar (
    .O(ybar[37]),
    .I0(abar[2]),
    .I1(bbar[5])
  );
  //AND U71
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U71 (
    .O(y[36]),
    .I0(a[2]),
    .I1(b[4])
  );
  //OR U71bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U71bar (
    .O(ybar[36]),
    .I0(abar[2]),
    .I1(bbar[4])
  );
  //AND U72
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U72 (
    .O(y[35]),
    .I0(a[2]),
    .I1(b[3])
  );
  //OR U72bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U72bar (
    .O(ybar[35]),
    .I0(abar[2]),
    .I1(bbar[3])
  );
  //AND U73
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U73 (
    .O(y[34]),
    .I0(a[2]),
    .I1(b[2])
  );
  //OR U73bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U73bar (
    .O(ybar[34]),
    .I0(abar[2]),
    .I1(bbar[2])
  );
  //AND U74
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U74 (
    .O(y[33]),
    .I0(a[2]),
    .I1(b[1])
  );
  //OR U74bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U74bar (
    .O(ybar[33]),
    .I0(abar[2]),
    .I1(bbar[1])
  );
  //AND U75
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U75 (
    .O(y[32]),
    .I0(a[2]),
    .I1(b[0])
  );
  //OR U75bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U75bar (
    .O(ybar[32]),
    .I0(abar[2]),
    .I1(bbar[0])
  );
  //AND U76
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U76 (
    .O(y[31]),
    .I0(a[1]),
    .I1(b[15])
  );
  //OR U76bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U76bar (
    .O(ybar[31]),
    .I0(abar[1]),
    .I1(bbar[15])
  );
  //AND U77
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U77 (
    .O(y[30]),
    .I0(a[1]),
    .I1(b[14])
  );
  //OR U77bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U77bar (
    .O(ybar[30]),
    .I0(abar[1]),
    .I1(bbar[14])
  );
  //AND U78
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U78 (
    .O(y[2]),
    .I0(b[2]),
    .I1(a[0])
  );
  //OR U78bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U78bar (
    .O(ybar[2]),
    .I0(bbar[2]),
    .I1(abar[0])
  );
  //AND U79
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U79 (
    .O(y[29]),
    .I0(a[1]),
    .I1(b[13])
  );
  //OR U79bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U79bar (
    .O(ybar[29]),
    .I0(abar[1]),
    .I1(bbar[13])
  );
  //AND U80
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U80 (
    .O(y[28]),
    .I0(a[1]),
    .I1(b[12])
  );
  //OR U80bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U80bar (
    .O(ybar[28]),
    .I0(abar[1]),
    .I1(bbar[12])
  );
  //AND U81
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U81 (
    .O(y[27]),
    .I0(a[1]),
    .I1(b[11])
  );
  //OR U81bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U81bar (
    .O(ybar[27]),
    .I0(abar[1]),
    .I1(bbar[11])
  );
  //AND U82
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U82 (
    .O(y[26]),
    .I0(a[1]),
    .I1(b[10])
  );
  //OR U82bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U82bar (
    .O(ybar[26]),
    .I0(abar[1]),
    .I1(bbar[10])
  );
  //AND U83
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U83 (
    .O(y[25]),
    .I0(a[1]),
    .I1(b[9])
  );
  //OR U83bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U83bar (
    .O(ybar[25]),
    .I0(abar[1]),
    .I1(bbar[9])
  );
  //AND U84
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U84 (
    .O(y[255]),
    .I0(a[15]),
    .I1(b[15])
  );
  //OR U84bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U84bar (
    .O(ybar[255]),
    .I0(abar[15]),
    .I1(bbar[15])
  );
  //AND U85
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U85 (
    .O(y[254]),
    .I0(a[15]),
    .I1(b[14])
  );
  //OR U85bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U85bar (
    .O(ybar[254]),
    .I0(abar[15]),
    .I1(bbar[14])
  );
  //AND U86
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U86 (
    .O(y[253]),
    .I0(a[15]),
    .I1(b[13])
  );
  //OR U86bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U86bar (
    .O(ybar[253]),
    .I0(abar[15]),
    .I1(bbar[13])
  );
  //AND U87
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U87 (
    .O(y[252]),
    .I0(a[15]),
    .I1(b[12])
  );
  //OR U87bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U87bar (
    .O(ybar[252]),
    .I0(abar[15]),
    .I1(bbar[12])
  );
  //AND U88
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U88 (
    .O(y[251]),
    .I0(a[15]),
    .I1(b[11])
  );
  //OR U88bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U88bar (
    .O(ybar[251]),
    .I0(abar[15]),
    .I1(bbar[11])
  );
  //AND U89
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U89 (
    .O(y[250]),
    .I0(a[15]),
    .I1(b[10])
  );
  //OR U89bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U89bar (
    .O(ybar[250]),
    .I0(abar[15]),
    .I1(bbar[10])
  );
  //AND U90
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U90 (
    .O(y[24]),
    .I0(a[1]),
    .I1(b[8])
  );
  //OR U90bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U90bar (
    .O(ybar[24]),
    .I0(abar[1]),
    .I1(bbar[8])
  );
  //AND U91
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U91 (
    .O(y[249]),
    .I0(a[15]),
    .I1(b[9])
  );
  //OR U91bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U91bar (
    .O(ybar[249]),
    .I0(abar[15]),
    .I1(bbar[9])
  );
  //AND U92
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U92 (
    .O(y[248]),
    .I0(a[15]),
    .I1(b[8])
  );
  //OR U92bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U92bar (
    .O(ybar[248]),
    .I0(abar[15]),
    .I1(bbar[8])
  );
  //AND U93
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U93 (
    .O(y[247]),
    .I0(a[15]),
    .I1(b[7])
  );
  //OR U93bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U93bar (
    .O(ybar[247]),
    .I0(abar[15]),
    .I1(bbar[7])
  );
  //AND U94
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U94 (
    .O(y[246]),
    .I0(a[15]),
    .I1(b[6])
  );
  //OR U94bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U94bar (
    .O(ybar[246]),
    .I0(abar[15]),
    .I1(bbar[6])
  );
  //AND U95
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U95 (
    .O(y[245]),
    .I0(a[15]),
    .I1(b[5])
  );
  //OR U95bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U95bar (
    .O(ybar[245]),
    .I0(abar[15]),
    .I1(bbar[5])
  );
  //AND U96
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U96 (
    .O(y[244]),
    .I0(a[15]),
    .I1(b[4])
  );
  //OR U96bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U96bar (
    .O(ybar[244]),
    .I0(abar[15]),
    .I1(bbar[4])
  );
  //AND U97
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U97 (
    .O(y[243]),
    .I0(a[15]),
    .I1(b[3])
  );
  //OR U97bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U97bar (
    .O(ybar[243]),
    .I0(abar[15]),
    .I1(bbar[3])
  );
  //AND U98
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U98 (
    .O(y[242]),
    .I0(a[15]),
    .I1(b[2])
  );
  //OR U98bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U98bar (
    .O(ybar[242]),
    .I0(abar[15]),
    .I1(bbar[2])
  );
  //AND U99
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U99 (
    .O(y[241]),
    .I0(a[15]),
    .I1(b[1])
  );
  //OR U99bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U99bar (
    .O(ybar[241]),
    .I0(abar[15]),
    .I1(bbar[1])
  );
  //AND U100
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U100 (
    .O(y[240]),
    .I0(a[15]),
    .I1(b[0])
  );
  //OR U100bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U100bar (
    .O(ybar[240]),
    .I0(abar[15]),
    .I1(bbar[0])
  );
  //AND U101
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U101 (
    .O(y[23]),
    .I0(a[1]),
    .I1(b[7])
  );
  //OR U101bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U101bar (
    .O(ybar[23]),
    .I0(abar[1]),
    .I1(bbar[7])
  );
  //AND U102
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U102 (
    .O(y[239]),
    .I0(a[14]),
    .I1(b[15])
  );
  //OR U102bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U102bar (
    .O(ybar[239]),
    .I0(abar[14]),
    .I1(bbar[15])
  );
  //AND U103
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U103 (
    .O(y[238]),
    .I0(a[14]),
    .I1(b[14])
  );
  //OR U103bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U103bar (
    .O(ybar[238]),
    .I0(abar[14]),
    .I1(bbar[14])
  );
  //AND U104
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U104 (
    .O(y[237]),
    .I0(a[14]),
    .I1(b[13])
  );
  //OR U104bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U104bar (
    .O(ybar[237]),
    .I0(abar[14]),
    .I1(bbar[13])
  );
  //AND U105
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U105 (
    .O(y[236]),
    .I0(a[14]),
    .I1(b[12])
  );
  //OR U105bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U105bar (
    .O(ybar[236]),
    .I0(abar[14]),
    .I1(bbar[12])
  );
  //AND U106
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U106 (
    .O(y[235]),
    .I0(a[14]),
    .I1(b[11])
  );
  //OR U106bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U106bar (
    .O(ybar[235]),
    .I0(abar[14]),
    .I1(bbar[11])
  );
  //AND U107
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U107 (
    .O(y[234]),
    .I0(a[14]),
    .I1(b[10])
  );
  //OR U107bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U107bar (
    .O(ybar[234]),
    .I0(abar[14]),
    .I1(bbar[10])
  );
  //AND U108
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U108 (
    .O(y[233]),
    .I0(a[14]),
    .I1(b[9])
  );
  //OR U108bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U108bar (
    .O(ybar[233]),
    .I0(abar[14]),
    .I1(bbar[9])
  );
  //AND U109
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U109 (
    .O(y[232]),
    .I0(a[14]),
    .I1(b[8])
  );
  //OR U109bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U109bar (
    .O(ybar[232]),
    .I0(abar[14]),
    .I1(bbar[8])
  );
  //AND U110
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U110 (
    .O(y[231]),
    .I0(a[14]),
    .I1(b[7])
  );
  //OR U110bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U110bar (
    .O(ybar[231]),
    .I0(abar[14]),
    .I1(bbar[7])
  );
  //AND U111
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U111 (
    .O(y[230]),
    .I0(a[14]),
    .I1(b[6])
  );
  //OR U111bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U111bar (
    .O(ybar[230]),
    .I0(abar[14]),
    .I1(bbar[6])
  );
  //AND U112
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U112 (
    .O(y[22]),
    .I0(a[1]),
    .I1(b[6])
  );
  //OR U112bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U112bar (
    .O(ybar[22]),
    .I0(abar[1]),
    .I1(bbar[6])
  );
  //AND U113
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U113 (
    .O(y[229]),
    .I0(a[14]),
    .I1(b[5])
  );
  //OR U113bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U113bar (
    .O(ybar[229]),
    .I0(abar[14]),
    .I1(bbar[5])
  );
  //AND U114
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U114 (
    .O(y[228]),
    .I0(a[14]),
    .I1(b[4])
  );
  //OR U114bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U114bar (
    .O(ybar[228]),
    .I0(abar[14]),
    .I1(bbar[4])
  );
  //AND U115
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U115 (
    .O(y[227]),
    .I0(a[14]),
    .I1(b[3])
  );
  //OR U115bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U115bar (
    .O(ybar[227]),
    .I0(abar[14]),
    .I1(bbar[3])
  );
  //AND U116
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U116 (
    .O(y[226]),
    .I0(a[14]),
    .I1(b[2])
  );
  //OR U116bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U116bar (
    .O(ybar[226]),
    .I0(abar[14]),
    .I1(bbar[2])
  );
  //AND U117
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U117 (
    .O(y[225]),
    .I0(a[14]),
    .I1(b[1])
  );
  //OR U117bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U117bar (
    .O(ybar[225]),
    .I0(abar[14]),
    .I1(bbar[1])
  );
  //AND U118
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U118 (
    .O(y[224]),
    .I0(a[14]),
    .I1(b[0])
  );
  //OR U118bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U118bar (
    .O(ybar[224]),
    .I0(abar[14]),
    .I1(bbar[0])
  );
  //AND U119
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U119 (
    .O(y[223]),
    .I0(a[13]),
    .I1(b[15])
  );
  //OR U119bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U119bar (
    .O(ybar[223]),
    .I0(abar[13]),
    .I1(bbar[15])
  );
  //AND U120
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U120 (
    .O(y[222]),
    .I0(a[13]),
    .I1(b[14])
  );
  //OR U120bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U120bar (
    .O(ybar[222]),
    .I0(abar[13]),
    .I1(bbar[14])
  );
  //AND U121
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U121 (
    .O(y[221]),
    .I0(a[13]),
    .I1(b[13])
  );
  //OR U121bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U121bar (
    .O(ybar[221]),
    .I0(abar[13]),
    .I1(bbar[13])
  );
  //AND U122
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U122 (
    .O(y[220]),
    .I0(a[13]),
    .I1(b[12])
  );
  //OR U122bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U122bar (
    .O(ybar[220]),
    .I0(abar[13]),
    .I1(bbar[12])
  );
  //AND U123
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U123 (
    .O(y[21]),
    .I0(a[1]),
    .I1(b[5])
  );
  //OR U123bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U123bar (
    .O(ybar[21]),
    .I0(abar[1]),
    .I1(bbar[5])
  );
  //AND U124
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U124 (
    .O(y[219]),
    .I0(a[13]),
    .I1(b[11])
  );
  //OR U124bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U124bar (
    .O(ybar[219]),
    .I0(abar[13]),
    .I1(bbar[11])
  );
  //AND U125
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U125 (
    .O(y[218]),
    .I0(a[13]),
    .I1(b[10])
  );
  //OR U125bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U125bar (
    .O(ybar[218]),
    .I0(abar[13]),
    .I1(bbar[10])
  );
  //AND U126
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U126 (
    .O(y[217]),
    .I0(a[13]),
    .I1(b[9])
  );
  //OR U126bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U126bar (
    .O(ybar[217]),
    .I0(abar[13]),
    .I1(bbar[9])
  );
  //AND U127
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U127 (
    .O(y[216]),
    .I0(a[13]),
    .I1(b[8])
  );
  //OR U127bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U127bar (
    .O(ybar[216]),
    .I0(abar[13]),
    .I1(bbar[8])
  );
  //AND U128
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U128 (
    .O(y[215]),
    .I0(a[13]),
    .I1(b[7])
  );
  //OR U128bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U128bar (
    .O(ybar[215]),
    .I0(abar[13]),
    .I1(bbar[7])
  );
  //AND U129
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U129 (
    .O(y[214]),
    .I0(a[13]),
    .I1(b[6])
  );
  //OR U129bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U129bar (
    .O(ybar[214]),
    .I0(abar[13]),
    .I1(bbar[6])
  );
  //AND U130
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U130 (
    .O(y[213]),
    .I0(a[13]),
    .I1(b[5])
  );
  //OR U130bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U130bar (
    .O(ybar[213]),
    .I0(abar[13]),
    .I1(bbar[5])
  );
  //AND U131
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U131 (
    .O(y[212]),
    .I0(a[13]),
    .I1(b[4])
  );
  //OR U131bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U131bar (
    .O(ybar[212]),
    .I0(abar[13]),
    .I1(bbar[4])
  );
  //AND U132
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U132 (
    .O(y[211]),
    .I0(a[13]),
    .I1(b[3])
  );
  //OR U132bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U132bar (
    .O(ybar[211]),
    .I0(abar[13]),
    .I1(bbar[3])
  );
  //AND U133
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U133 (
    .O(y[210]),
    .I0(a[13]),
    .I1(b[2])
  );
  //OR U133bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U133bar (
    .O(ybar[210]),
    .I0(abar[13]),
    .I1(bbar[2])
  );
  //AND U134
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U134 (
    .O(y[20]),
    .I0(a[1]),
    .I1(b[4])
  );
  //OR U134bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U134bar (
    .O(ybar[20]),
    .I0(abar[1]),
    .I1(bbar[4])
  );
  //AND U135
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U135 (
    .O(y[209]),
    .I0(a[13]),
    .I1(b[1])
  );
  //OR U135bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U135bar (
    .O(ybar[209]),
    .I0(abar[13]),
    .I1(bbar[1])
  );
  //AND U136
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U136 (
    .O(y[208]),
    .I0(a[13]),
    .I1(b[0])
  );
  //OR U136bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U136bar (
    .O(ybar[208]),
    .I0(abar[13]),
    .I1(bbar[0])
  );
  //AND U137
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U137 (
    .O(y[207]),
    .I0(a[12]),
    .I1(b[15])
  );
  //OR U137bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U137bar (
    .O(ybar[207]),
    .I0(abar[12]),
    .I1(bbar[15])
  );
  //AND U138
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U138 (
    .O(y[206]),
    .I0(a[12]),
    .I1(b[14])
  );
  //OR U138bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U138bar (
    .O(ybar[206]),
    .I0(abar[12]),
    .I1(bbar[14])
  );
  //AND U139
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U139 (
    .O(y[205]),
    .I0(a[12]),
    .I1(b[13])
  );
  //OR U139bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U139bar (
    .O(ybar[205]),
    .I0(abar[12]),
    .I1(bbar[13])
  );
  //AND U140
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U140 (
    .O(y[204]),
    .I0(a[12]),
    .I1(b[12])
  );
  //OR U140bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U140bar (
    .O(ybar[204]),
    .I0(abar[12]),
    .I1(bbar[12])
  );
  //AND U141
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U141 (
    .O(y[203]),
    .I0(a[12]),
    .I1(b[11])
  );
  //OR U141bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U141bar (
    .O(ybar[203]),
    .I0(abar[12]),
    .I1(bbar[11])
  );
  //AND U142
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U142 (
    .O(y[202]),
    .I0(a[12]),
    .I1(b[10])
  );
  //OR U142bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U142bar (
    .O(ybar[202]),
    .I0(abar[12]),
    .I1(bbar[10])
  );
  //AND U143
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U143 (
    .O(y[201]),
    .I0(a[12]),
    .I1(b[9])
  );
  //OR U143bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U143bar (
    .O(ybar[201]),
    .I0(abar[12]),
    .I1(bbar[9])
  );
  //AND U144
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U144 (
    .O(y[200]),
    .I0(a[12]),
    .I1(b[8])
  );
  //OR U144bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U144bar (
    .O(ybar[200]),
    .I0(abar[12]),
    .I1(bbar[8])
  );
  //AND U145
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U145 (
    .O(y[1]),
    .I0(b[1]),
    .I1(a[0])
  );
  //OR U145bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U145bar (
    .O(ybar[1]),
    .I0(bbar[1]),
    .I1(abar[0])
  );
  //AND U146
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U146 (
    .O(y[19]),
    .I0(a[1]),
    .I1(b[3])
  );
  //OR U146bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U146bar (
    .O(ybar[19]),
    .I0(abar[1]),
    .I1(bbar[3])
  );
  //AND U147
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U147 (
    .O(y[199]),
    .I0(a[12]),
    .I1(b[7])
  );
  //OR U147bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U147bar (
    .O(ybar[199]),
    .I0(abar[12]),
    .I1(bbar[7])
  );
  //AND U148
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U148 (
    .O(y[198]),
    .I0(a[12]),
    .I1(b[6])
  );
  //OR U148bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U148bar (
    .O(ybar[198]),
    .I0(abar[12]),
    .I1(bbar[6])
  );
  //AND U149
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U149 (
    .O(y[197]),
    .I0(a[12]),
    .I1(b[5])
  );
  //OR U149bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U149bar (
    .O(ybar[197]),
    .I0(abar[12]),
    .I1(bbar[5])
  );
  //AND U150
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U150 (
    .O(y[196]),
    .I0(a[12]),
    .I1(b[4])
  );
  //OR U150bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U150bar (
    .O(ybar[196]),
    .I0(abar[12]),
    .I1(bbar[4])
  );
  //AND U151
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U151 (
    .O(y[195]),
    .I0(a[12]),
    .I1(b[3])
  );
  //OR U151bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U151bar (
    .O(ybar[195]),
    .I0(abar[12]),
    .I1(bbar[3])
  );
  //AND U152
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U152 (
    .O(y[194]),
    .I0(a[12]),
    .I1(b[2])
  );
  //OR U152bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U152bar (
    .O(ybar[194]),
    .I0(abar[12]),
    .I1(bbar[2])
  );
  //AND U153
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U153 (
    .O(y[193]),
    .I0(a[12]),
    .I1(b[1])
  );
  //OR U153bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U153bar (
    .O(ybar[193]),
    .I0(abar[12]),
    .I1(bbar[1])
  );
  //AND U154
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U154 (
    .O(y[192]),
    .I0(a[12]),
    .I1(b[0])
  );
  //OR U154bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U154bar (
    .O(ybar[192]),
    .I0(abar[12]),
    .I1(bbar[0])
  );
  //AND U155
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U155 (
    .O(y[191]),
    .I0(a[11]),
    .I1(b[15])
  );
  //OR U155bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U155bar (
    .O(ybar[191]),
    .I0(abar[11]),
    .I1(bbar[15])
  );
  //AND U156
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U156 (
    .O(y[190]),
    .I0(a[11]),
    .I1(b[14])
  );
  //OR U156bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U156bar (
    .O(ybar[190]),
    .I0(abar[11]),
    .I1(bbar[14])
  );
  //AND U157
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U157 (
    .O(y[18]),
    .I0(a[1]),
    .I1(b[2])
  );
  //OR U157bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U157bar (
    .O(ybar[18]),
    .I0(abar[1]),
    .I1(bbar[2])
  );
  //AND U158
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U158 (
    .O(y[189]),
    .I0(a[11]),
    .I1(b[13])
  );
  //OR U158bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U158bar (
    .O(ybar[189]),
    .I0(abar[11]),
    .I1(bbar[13])
  );
  //AND U159
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U159 (
    .O(y[188]),
    .I0(a[11]),
    .I1(b[12])
  );
  //OR U159bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U159bar (
    .O(ybar[188]),
    .I0(abar[11]),
    .I1(bbar[12])
  );
  //AND U160
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U160 (
    .O(y[187]),
    .I0(a[11]),
    .I1(b[11])
  );
  //OR U160bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U160bar (
    .O(ybar[187]),
    .I0(abar[11]),
    .I1(bbar[11])
  );
  //AND U161
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U161 (
    .O(y[186]),
    .I0(a[11]),
    .I1(b[10])
  );
  //OR U161bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U161bar (
    .O(ybar[186]),
    .I0(abar[11]),
    .I1(bbar[10])
  );
  //AND U162
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U162 (
    .O(y[185]),
    .I0(a[11]),
    .I1(b[9])
  );
  //OR U162bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U162bar (
    .O(ybar[185]),
    .I0(abar[11]),
    .I1(bbar[9])
  );
  //AND U163
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U163 (
    .O(y[184]),
    .I0(a[11]),
    .I1(b[8])
  );
  //OR U163bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U163bar (
    .O(ybar[184]),
    .I0(abar[11]),
    .I1(bbar[8])
  );
  //AND U164
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U164 (
    .O(y[183]),
    .I0(a[11]),
    .I1(b[7])
  );
  //OR U164bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U164bar (
    .O(ybar[183]),
    .I0(abar[11]),
    .I1(bbar[7])
  );
  //AND U165
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U165 (
    .O(y[182]),
    .I0(a[11]),
    .I1(b[6])
  );
  //OR U165bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U165bar (
    .O(ybar[182]),
    .I0(abar[11]),
    .I1(bbar[6])
  );
  //AND U166
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U166 (
    .O(y[181]),
    .I0(a[11]),
    .I1(b[5])
  );
  //OR U166bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U166bar (
    .O(ybar[181]),
    .I0(abar[11]),
    .I1(bbar[5])
  );
  //AND U167
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U167 (
    .O(y[180]),
    .I0(a[11]),
    .I1(b[4])
  );
  //OR U167bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U167bar (
    .O(ybar[180]),
    .I0(abar[11]),
    .I1(bbar[4])
  );
  //AND U168
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U168 (
    .O(y[17]),
    .I0(a[1]),
    .I1(b[1])
  );
  //OR U168bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U168bar (
    .O(ybar[17]),
    .I0(abar[1]),
    .I1(bbar[1])
  );
  //AND U169
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U169 (
    .O(y[179]),
    .I0(a[11]),
    .I1(b[3])
  );
  //OR U169bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U169bar (
    .O(ybar[179]),
    .I0(abar[11]),
    .I1(bbar[3])
  );
  //AND U170
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U170 (
    .O(y[178]),
    .I0(a[11]),
    .I1(b[2])
  );
  //OR U170bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U170bar (
    .O(ybar[178]),
    .I0(abar[11]),
    .I1(bbar[2])
  );
  //AND U171
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U171 (
    .O(y[177]),
    .I0(a[11]),
    .I1(b[1])
  );
  //OR U171bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U171bar (
    .O(ybar[177]),
    .I0(abar[11]),
    .I1(bbar[1])
  );
  //AND U172
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U172 (
    .O(y[176]),
    .I0(a[11]),
    .I1(b[0])
  );
  //OR U172bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U172bar (
    .O(ybar[176]),
    .I0(abar[11]),
    .I1(bbar[0])
  );
  //AND U173
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U173 (
    .O(y[175]),
    .I0(a[10]),
    .I1(b[15])
  );
  //OR U173bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U173bar (
    .O(ybar[175]),
    .I0(abar[10]),
    .I1(bbar[15])
  );
  //AND U174
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U174 (
    .O(y[174]),
    .I0(a[10]),
    .I1(b[14])
  );
  //OR U174bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U174bar (
    .O(ybar[174]),
    .I0(abar[10]),
    .I1(bbar[14])
  );
  //AND U175
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U175 (
    .O(y[173]),
    .I0(a[10]),
    .I1(b[13])
  );
  //OR U175bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U175bar (
    .O(ybar[173]),
    .I0(abar[10]),
    .I1(bbar[13])
  );
  //AND U176
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U176 (
    .O(y[172]),
    .I0(a[10]),
    .I1(b[12])
  );
  //OR U176bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U176bar (
    .O(ybar[172]),
    .I0(abar[10]),
    .I1(bbar[12])
  );
  //AND U177
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U177 (
    .O(y[171]),
    .I0(a[10]),
    .I1(b[11])
  );
  //OR U177bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U177bar (
    .O(ybar[171]),
    .I0(abar[10]),
    .I1(bbar[11])
  );
  //AND U178
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U178 (
    .O(y[170]),
    .I0(a[10]),
    .I1(b[10])
  );
  //OR U178bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U178bar (
    .O(ybar[170]),
    .I0(abar[10]),
    .I1(bbar[10])
  );
  //AND U179
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U179 (
    .O(y[16]),
    .I0(a[1]),
    .I1(b[0])
  );
  //OR U179bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U179bar (
    .O(ybar[16]),
    .I0(abar[1]),
    .I1(bbar[0])
  );
  //AND U180
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U180 (
    .O(y[169]),
    .I0(a[10]),
    .I1(b[9])
  );
  //OR U180bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U180bar (
    .O(ybar[169]),
    .I0(abar[10]),
    .I1(bbar[9])
  );
  //AND U181
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U181 (
    .O(y[168]),
    .I0(a[10]),
    .I1(b[8])
  );
  //OR U181bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U181bar (
    .O(ybar[168]),
    .I0(abar[10]),
    .I1(bbar[8])
  );
  //AND U182
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U182 (
    .O(y[167]),
    .I0(a[10]),
    .I1(b[7])
  );
  //OR U182bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U182bar (
    .O(ybar[167]),
    .I0(abar[10]),
    .I1(bbar[7])
  );
  //AND U183
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U183 (
    .O(y[166]),
    .I0(a[10]),
    .I1(b[6])
  );
  //OR U183bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U183bar (
    .O(ybar[166]),
    .I0(abar[10]),
    .I1(bbar[6])
  );
  //AND U184
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U184 (
    .O(y[165]),
    .I0(a[10]),
    .I1(b[5])
  );
  //OR U184bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U184bar (
    .O(ybar[165]),
    .I0(abar[10]),
    .I1(bbar[5])
  );
  //AND U185
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U185 (
    .O(y[164]),
    .I0(a[10]),
    .I1(b[4])
  );
  //OR U185bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U185bar (
    .O(ybar[164]),
    .I0(abar[10]),
    .I1(bbar[4])
  );
  //AND U186
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U186 (
    .O(y[163]),
    .I0(a[10]),
    .I1(b[3])
  );
  //OR U186bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U186bar (
    .O(ybar[163]),
    .I0(abar[10]),
    .I1(bbar[3])
  );
  //AND U187
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U187 (
    .O(y[162]),
    .I0(a[10]),
    .I1(b[2])
  );
  //OR U187bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U187bar (
    .O(ybar[162]),
    .I0(abar[10]),
    .I1(bbar[2])
  );
  //AND U188
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U188 (
    .O(y[161]),
    .I0(a[10]),
    .I1(b[1])
  );
  //OR U188bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U188bar (
    .O(ybar[161]),
    .I0(abar[10]),
    .I1(bbar[1])
  );
  //AND U189
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U189 (
    .O(y[160]),
    .I0(a[10]),
    .I1(b[0])
  );
  //OR U189bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U189bar (
    .O(ybar[160]),
    .I0(abar[10]),
    .I1(bbar[0])
  );
  //AND U190
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U190 (
    .O(y[15]),
    .I0(b[15]),
    .I1(a[0])
  );
  //OR U190bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U190bar (
    .O(ybar[15]),
    .I0(bbar[15]),
    .I1(abar[0])
  );
  //AND U191
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U191 (
    .O(y[159]),
    .I0(a[9]),
    .I1(b[15])
  );
  //OR U191bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U191bar (
    .O(ybar[159]),
    .I0(abar[9]),
    .I1(bbar[15])
  );
  //AND U192
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U192 (
    .O(y[158]),
    .I0(a[9]),
    .I1(b[14])
  );
  //OR U192bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U192bar (
    .O(ybar[158]),
    .I0(abar[9]),
    .I1(bbar[14])
  );
  //AND U193
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U193 (
    .O(y[157]),
    .I0(a[9]),
    .I1(b[13])
  );
  //OR U193bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U193bar (
    .O(ybar[157]),
    .I0(abar[9]),
    .I1(bbar[13])
  );
  //AND U194
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U194 (
    .O(y[156]),
    .I0(a[9]),
    .I1(b[12])
  );
  //OR U194bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U194bar (
    .O(ybar[156]),
    .I0(abar[9]),
    .I1(bbar[12])
  );
  //AND U195
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U195 (
    .O(y[155]),
    .I0(a[9]),
    .I1(b[11])
  );
  //OR U195bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U195bar (
    .O(ybar[155]),
    .I0(abar[9]),
    .I1(bbar[11])
  );
  //AND U196
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U196 (
    .O(y[154]),
    .I0(a[9]),
    .I1(b[10])
  );
  //OR U196bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U196bar (
    .O(ybar[154]),
    .I0(abar[9]),
    .I1(bbar[10])
  );
  //AND U197
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U197 (
    .O(y[153]),
    .I0(a[9]),
    .I1(b[9])
  );
  //OR U197bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U197bar (
    .O(ybar[153]),
    .I0(abar[9]),
    .I1(bbar[9])
  );
  //AND U198
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U198 (
    .O(y[152]),
    .I0(a[9]),
    .I1(b[8])
  );
  //OR U198bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U198bar (
    .O(ybar[152]),
    .I0(abar[9]),
    .I1(bbar[8])
  );
  //AND U199
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U199 (
    .O(y[151]),
    .I0(a[9]),
    .I1(b[7])
  );
  //OR U199bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U199bar (
    .O(ybar[151]),
    .I0(abar[9]),
    .I1(bbar[7])
  );
  //AND U200
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U200 (
    .O(y[150]),
    .I0(a[9]),
    .I1(b[6])
  );
  //OR U200bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U200bar (
    .O(ybar[150]),
    .I0(abar[9]),
    .I1(bbar[6])
  );
  //AND U201
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U201 (
    .O(y[14]),
    .I0(b[14]),
    .I1(a[0])
  );
  //OR U201bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U201bar (
    .O(ybar[14]),
    .I0(bbar[14]),
    .I1(abar[0])
  );
  //AND U202
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U202 (
    .O(y[149]),
    .I0(a[9]),
    .I1(b[5])
  );
  //OR U202bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U202bar (
    .O(ybar[149]),
    .I0(abar[9]),
    .I1(bbar[5])
  );
  //AND U203
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U203 (
    .O(y[148]),
    .I0(a[9]),
    .I1(b[4])
  );
  //OR U203bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U203bar (
    .O(ybar[148]),
    .I0(abar[9]),
    .I1(bbar[4])
  );
  //AND U204
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U204 (
    .O(y[147]),
    .I0(a[9]),
    .I1(b[3])
  );
  //OR U204bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U204bar (
    .O(ybar[147]),
    .I0(abar[9]),
    .I1(bbar[3])
  );
  //AND U205
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U205 (
    .O(y[146]),
    .I0(a[9]),
    .I1(b[2])
  );
  //OR U205bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U205bar (
    .O(ybar[146]),
    .I0(abar[9]),
    .I1(bbar[2])
  );
  //AND U206
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U206 (
    .O(y[145]),
    .I0(a[9]),
    .I1(b[1])
  );
  //OR U206bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U206bar (
    .O(ybar[145]),
    .I0(abar[9]),
    .I1(bbar[1])
  );
  //AND U207
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U207 (
    .O(y[144]),
    .I0(a[9]),
    .I1(b[0])
  );
  //OR U207bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U207bar (
    .O(ybar[144]),
    .I0(abar[9]),
    .I1(bbar[0])
  );
  //AND U208
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U208 (
    .O(y[143]),
    .I0(a[8]),
    .I1(b[15])
  );
  //OR U208bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U208bar (
    .O(ybar[143]),
    .I0(abar[8]),
    .I1(bbar[15])
  );
  //AND U209
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U209 (
    .O(y[142]),
    .I0(a[8]),
    .I1(b[14])
  );
  //OR U209bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U209bar (
    .O(ybar[142]),
    .I0(abar[8]),
    .I1(bbar[14])
  );
  //AND U210
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U210 (
    .O(y[141]),
    .I0(a[8]),
    .I1(b[13])
  );
  //OR U210bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U210bar (
    .O(ybar[141]),
    .I0(abar[8]),
    .I1(bbar[13])
  );
  //AND U211
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U211 (
    .O(y[140]),
    .I0(a[8]),
    .I1(b[12])
  );
  //OR U211bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U211bar (
    .O(ybar[140]),
    .I0(abar[8]),
    .I1(bbar[12])
  );
  //AND U212
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U212 (
    .O(y[13]),
    .I0(b[13]),
    .I1(a[0])
  );
  //OR U212bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U212bar (
    .O(ybar[13]),
    .I0(bbar[13]),
    .I1(abar[0])
  );
  //AND U213
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U213 (
    .O(y[139]),
    .I0(a[8]),
    .I1(b[11])
  );
  //OR U213bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U213bar (
    .O(ybar[139]),
    .I0(abar[8]),
    .I1(bbar[11])
  );
  //AND U214
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U214 (
    .O(y[138]),
    .I0(a[8]),
    .I1(b[10])
  );
  //OR U214bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U214bar (
    .O(ybar[138]),
    .I0(abar[8]),
    .I1(bbar[10])
  );
  //AND U215
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U215 (
    .O(y[137]),
    .I0(a[8]),
    .I1(b[9])
  );
  //OR U215bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U215bar (
    .O(ybar[137]),
    .I0(abar[8]),
    .I1(bbar[9])
  );
  //AND U216
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U216 (
    .O(y[136]),
    .I0(a[8]),
    .I1(b[8])
  );
  //OR U216bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U216bar (
    .O(ybar[136]),
    .I0(abar[8]),
    .I1(bbar[8])
  );
  //AND U217
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U217 (
    .O(y[135]),
    .I0(a[8]),
    .I1(b[7])
  );
  //OR U217bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U217bar (
    .O(ybar[135]),
    .I0(abar[8]),
    .I1(bbar[7])
  );
  //AND U218
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U218 (
    .O(y[134]),
    .I0(a[8]),
    .I1(b[6])
  );
  //OR U218bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U218bar (
    .O(ybar[134]),
    .I0(abar[8]),
    .I1(bbar[6])
  );
  //AND U219
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U219 (
    .O(y[133]),
    .I0(a[8]),
    .I1(b[5])
  );
  //OR U219bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U219bar (
    .O(ybar[133]),
    .I0(abar[8]),
    .I1(bbar[5])
  );
  //AND U220
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U220 (
    .O(y[132]),
    .I0(a[8]),
    .I1(b[4])
  );
  //OR U220bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U220bar (
    .O(ybar[132]),
    .I0(abar[8]),
    .I1(bbar[4])
  );
  //AND U221
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U221 (
    .O(y[131]),
    .I0(a[8]),
    .I1(b[3])
  );
  //OR U221bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U221bar (
    .O(ybar[131]),
    .I0(abar[8]),
    .I1(bbar[3])
  );
  //AND U222
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U222 (
    .O(y[130]),
    .I0(a[8]),
    .I1(b[2])
  );
  //OR U222bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U222bar (
    .O(ybar[130]),
    .I0(abar[8]),
    .I1(bbar[2])
  );
  //AND U223
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U223 (
    .O(y[12]),
    .I0(b[12]),
    .I1(a[0])
  );
  //OR U223bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U223bar (
    .O(ybar[12]),
    .I0(bbar[12]),
    .I1(abar[0])
  );
  //AND U224
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U224 (
    .O(y[129]),
    .I0(a[8]),
    .I1(b[1])
  );
  //OR U224bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U224bar (
    .O(ybar[129]),
    .I0(abar[8]),
    .I1(bbar[1])
  );
  //AND U225
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U225 (
    .O(y[128]),
    .I0(a[8]),
    .I1(b[0])
  );
  //OR U225bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U225bar (
    .O(ybar[128]),
    .I0(abar[8]),
    .I1(bbar[0])
  );
  //AND U226
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U226 (
    .O(y[127]),
    .I0(a[7]),
    .I1(b[15])
  );
  //OR U226bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U226bar (
    .O(ybar[127]),
    .I0(abar[7]),
    .I1(bbar[15])
  );
  //AND U227
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U227 (
    .O(y[126]),
    .I0(a[7]),
    .I1(b[14])
  );
  //OR U227bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U227bar (
    .O(ybar[126]),
    .I0(abar[7]),
    .I1(bbar[14])
  );
  //AND U228
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U228 (
    .O(y[125]),
    .I0(a[7]),
    .I1(b[13])
  );
  //OR U228bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U228bar (
    .O(ybar[125]),
    .I0(abar[7]),
    .I1(bbar[13])
  );
  //AND U229
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U229 (
    .O(y[124]),
    .I0(a[7]),
    .I1(b[12])
  );
  //OR U229bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U229bar (
    .O(ybar[124]),
    .I0(abar[7]),
    .I1(bbar[12])
  );
  //AND U230
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U230 (
    .O(y[123]),
    .I0(a[7]),
    .I1(b[11])
  );
  //OR U230bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U230bar (
    .O(ybar[123]),
    .I0(abar[7]),
    .I1(bbar[11])
  );
  //AND U231
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U231 (
    .O(y[122]),
    .I0(a[7]),
    .I1(b[10])
  );
  //OR U231bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U231bar (
    .O(ybar[122]),
    .I0(abar[7]),
    .I1(bbar[10])
  );
  //AND U232
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U232 (
    .O(y[121]),
    .I0(a[7]),
    .I1(b[9])
  );
  //OR U232bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U232bar (
    .O(ybar[121]),
    .I0(abar[7]),
    .I1(bbar[9])
  );
  //AND U233
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U233 (
    .O(y[120]),
    .I0(a[7]),
    .I1(b[8])
  );
  //OR U233bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U233bar (
    .O(ybar[120]),
    .I0(abar[7]),
    .I1(bbar[8])
  );
  //AND U234
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U234 (
    .O(y[11]),
    .I0(b[11]),
    .I1(a[0])
  );
  //OR U234bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U234bar (
    .O(ybar[11]),
    .I0(bbar[11]),
    .I1(abar[0])
  );
  //AND U235
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U235 (
    .O(y[119]),
    .I0(a[7]),
    .I1(b[7])
  );
  //OR U235bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U235bar (
    .O(ybar[119]),
    .I0(abar[7]),
    .I1(bbar[7])
  );
  //AND U236
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U236 (
    .O(y[118]),
    .I0(a[7]),
    .I1(b[6])
  );
  //OR U236bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U236bar (
    .O(ybar[118]),
    .I0(abar[7]),
    .I1(bbar[6])
  );
  //AND U237
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U237 (
    .O(y[117]),
    .I0(a[7]),
    .I1(b[5])
  );
  //OR U237bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U237bar (
    .O(ybar[117]),
    .I0(abar[7]),
    .I1(bbar[5])
  );
  //AND U238
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U238 (
    .O(y[116]),
    .I0(a[7]),
    .I1(b[4])
  );
  //OR U238bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U238bar (
    .O(ybar[116]),
    .I0(abar[7]),
    .I1(bbar[4])
  );
  //AND U239
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U239 (
    .O(y[115]),
    .I0(a[7]),
    .I1(b[3])
  );
  //OR U239bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U239bar (
    .O(ybar[115]),
    .I0(abar[7]),
    .I1(bbar[3])
  );
  //AND U240
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U240 (
    .O(y[114]),
    .I0(a[7]),
    .I1(b[2])
  );
  //OR U240bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U240bar (
    .O(ybar[114]),
    .I0(abar[7]),
    .I1(bbar[2])
  );
  //AND U241
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U241 (
    .O(y[113]),
    .I0(a[7]),
    .I1(b[1])
  );
  //OR U241bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U241bar (
    .O(ybar[113]),
    .I0(abar[7]),
    .I1(bbar[1])
  );
  //AND U242
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U242 (
    .O(y[112]),
    .I0(a[7]),
    .I1(b[0])
  );
  //OR U242bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U242bar (
    .O(ybar[112]),
    .I0(abar[7]),
    .I1(bbar[0])
  );
  //AND U243
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U243 (
    .O(y[111]),
    .I0(b[15]),
    .I1(a[6])
  );
  //OR U243bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U243bar (
    .O(ybar[111]),
    .I0(bbar[15]),
    .I1(abar[6])
  );
  //AND U244
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U244 (
    .O(y[110]),
    .I0(b[14]),
    .I1(a[6])
  );
  //OR U244bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U244bar (
    .O(ybar[110]),
    .I0(bbar[14]),
    .I1(abar[6])
  );
  //AND U245
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U245 (
    .O(y[10]),
    .I0(b[10]),
    .I1(a[0])
  );
  //OR U245bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U245bar (
    .O(ybar[10]),
    .I0(bbar[10]),
    .I1(abar[0])
  );
  //AND U246
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U246 (
    .O(y[109]),
    .I0(b[13]),
    .I1(a[6])
  );
  //OR U246bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U246bar (
    .O(ybar[109]),
    .I0(bbar[13]),
    .I1(abar[6])
  );
  //AND U247
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U247 (
    .O(y[108]),
    .I0(b[12]),
    .I1(a[6])
  );
  //OR U247bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U247bar (
    .O(ybar[108]),
    .I0(bbar[12]),
    .I1(abar[6])
  );
  //AND U248
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U248 (
    .O(y[107]),
    .I0(b[11]),
    .I1(a[6])
  );
  //OR U248bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U248bar (
    .O(ybar[107]),
    .I0(bbar[11]),
    .I1(abar[6])
  );
  //AND U249
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U249 (
    .O(y[106]),
    .I0(b[10]),
    .I1(a[6])
  );
  //OR U249bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U249bar (
    .O(ybar[106]),
    .I0(bbar[10]),
    .I1(abar[6])
  );
  //AND U250
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U250 (
    .O(y[105]),
    .I0(a[6]),
    .I1(b[9])
  );
  //OR U250bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U250bar (
    .O(ybar[105]),
    .I0(abar[6]),
    .I1(bbar[9])
  );
  //AND U251
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U251 (
    .O(y[104]),
    .I0(b[8]),
    .I1(a[6])
  );
  //OR U251bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U251bar (
    .O(ybar[104]),
    .I0(bbar[8]),
    .I1(abar[6])
  );
  //AND U252
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U252 (
    .O(y[103]),
    .I0(b[7]),
    .I1(a[6])
  );
  //OR U252bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U252bar (
    .O(ybar[103]),
    .I0(bbar[7]),
    .I1(abar[6])
  );
  //AND U253
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U253 (
    .O(y[102]),
    .I0(b[6]),
    .I1(a[6])
  );
  //OR U253bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U253bar (
    .O(ybar[102]),
    .I0(bbar[6]),
    .I1(abar[6])
  );
  //AND U254
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U254 (
    .O(y[101]),
    .I0(b[5]),
    .I1(a[6])
  );
  //OR U254bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U254bar (
    .O(ybar[101]),
    .I0(bbar[5]),
    .I1(abar[6])
  );
  //AND U255
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U255 (
    .O(y[100]),
    .I0(b[4]),
    .I1(a[6])
  );
  //OR U255bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U255bar (
    .O(ybar[100]),
    .I0(bbar[4]),
    .I1(abar[6])
  );
  //AND U256
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U256 (
    .O(y[0]),
    .I0(b[0]),
    .I1(a[0])
  );
  //OR U256bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U256bar (
    .O(ybar[0]),
    .I0(bbar[0]),
    .I1(abar[0])
  );
endmodule

module decode_6 ( in, out );

  input wire [7:0] in;
//input_done

  output wire [255:0] out;
//output_done

  wire [15:0] level1;
  wire [31:0] level2;
//wire_done

  CD2_24 cd_l1_1 ( .a(in[1]), .b(in[0]), .y(level1[3:0]) );
  CD2_23 cd_l1_2 ( .a(in[3]), .b(in[2]), .y(level1[7:4]) );
  CD2_22 cd_l1_3 ( .a(in[5]), .b(in[4]), .y(level1[11:8]) );
  CD2_21 cd_l1_4 ( .a(in[7]), .b(in[6]), .y(level1[15:12]) );
  CD4_12 cd_l2_1 ( .a(level1[7:4]), .b(level1[3:0]), .y(level2[15:0]) );
  CD4_11 cd_l2_2 ( .a(level1[15:12]), .b(level1[11:8]), .y(level2[31:16]) );
  CD16_6 cd_l3 ( .a(level2[31:16]), .b(level2[15:0]), .y(out) );
endmodule

module encode_6 ( in, out );

  input wire [255:0] in;
  wire [255:0] inbar;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
  assign inbar[8] = ~in[8];
  assign inbar[9] = ~in[9];
  assign inbar[10] = ~in[10];
  assign inbar[11] = ~in[11];
  assign inbar[12] = ~in[12];
  assign inbar[13] = ~in[13];
  assign inbar[14] = ~in[14];
  assign inbar[15] = ~in[15];
  assign inbar[16] = ~in[16];
  assign inbar[17] = ~in[17];
  assign inbar[18] = ~in[18];
  assign inbar[19] = ~in[19];
  assign inbar[20] = ~in[20];
  assign inbar[21] = ~in[21];
  assign inbar[22] = ~in[22];
  assign inbar[23] = ~in[23];
  assign inbar[24] = ~in[24];
  assign inbar[25] = ~in[25];
  assign inbar[26] = ~in[26];
  assign inbar[27] = ~in[27];
  assign inbar[28] = ~in[28];
  assign inbar[29] = ~in[29];
  assign inbar[30] = ~in[30];
  assign inbar[31] = ~in[31];
  assign inbar[32] = ~in[32];
  assign inbar[33] = ~in[33];
  assign inbar[34] = ~in[34];
  assign inbar[35] = ~in[35];
  assign inbar[36] = ~in[36];
  assign inbar[37] = ~in[37];
  assign inbar[38] = ~in[38];
  assign inbar[39] = ~in[39];
  assign inbar[40] = ~in[40];
  assign inbar[41] = ~in[41];
  assign inbar[42] = ~in[42];
  assign inbar[43] = ~in[43];
  assign inbar[44] = ~in[44];
  assign inbar[45] = ~in[45];
  assign inbar[46] = ~in[46];
  assign inbar[47] = ~in[47];
  assign inbar[48] = ~in[48];
  assign inbar[49] = ~in[49];
  assign inbar[50] = ~in[50];
  assign inbar[51] = ~in[51];
  assign inbar[52] = ~in[52];
  assign inbar[53] = ~in[53];
  assign inbar[54] = ~in[54];
  assign inbar[55] = ~in[55];
  assign inbar[56] = ~in[56];
  assign inbar[57] = ~in[57];
  assign inbar[58] = ~in[58];
  assign inbar[59] = ~in[59];
  assign inbar[60] = ~in[60];
  assign inbar[61] = ~in[61];
  assign inbar[62] = ~in[62];
  assign inbar[63] = ~in[63];
  assign inbar[64] = ~in[64];
  assign inbar[65] = ~in[65];
  assign inbar[66] = ~in[66];
  assign inbar[67] = ~in[67];
  assign inbar[68] = ~in[68];
  assign inbar[69] = ~in[69];
  assign inbar[70] = ~in[70];
  assign inbar[71] = ~in[71];
  assign inbar[72] = ~in[72];
  assign inbar[73] = ~in[73];
  assign inbar[74] = ~in[74];
  assign inbar[75] = ~in[75];
  assign inbar[76] = ~in[76];
  assign inbar[77] = ~in[77];
  assign inbar[78] = ~in[78];
  assign inbar[79] = ~in[79];
  assign inbar[80] = ~in[80];
  assign inbar[81] = ~in[81];
  assign inbar[82] = ~in[82];
  assign inbar[83] = ~in[83];
  assign inbar[84] = ~in[84];
  assign inbar[85] = ~in[85];
  assign inbar[86] = ~in[86];
  assign inbar[87] = ~in[87];
  assign inbar[88] = ~in[88];
  assign inbar[89] = ~in[89];
  assign inbar[90] = ~in[90];
  assign inbar[91] = ~in[91];
  assign inbar[92] = ~in[92];
  assign inbar[93] = ~in[93];
  assign inbar[94] = ~in[94];
  assign inbar[95] = ~in[95];
  assign inbar[96] = ~in[96];
  assign inbar[97] = ~in[97];
  assign inbar[98] = ~in[98];
  assign inbar[99] = ~in[99];
  assign inbar[100] = ~in[100];
  assign inbar[101] = ~in[101];
  assign inbar[102] = ~in[102];
  assign inbar[103] = ~in[103];
  assign inbar[104] = ~in[104];
  assign inbar[105] = ~in[105];
  assign inbar[106] = ~in[106];
  assign inbar[107] = ~in[107];
  assign inbar[108] = ~in[108];
  assign inbar[109] = ~in[109];
  assign inbar[110] = ~in[110];
  assign inbar[111] = ~in[111];
  assign inbar[112] = ~in[112];
  assign inbar[113] = ~in[113];
  assign inbar[114] = ~in[114];
  assign inbar[115] = ~in[115];
  assign inbar[116] = ~in[116];
  assign inbar[117] = ~in[117];
  assign inbar[118] = ~in[118];
  assign inbar[119] = ~in[119];
  assign inbar[120] = ~in[120];
  assign inbar[121] = ~in[121];
  assign inbar[122] = ~in[122];
  assign inbar[123] = ~in[123];
  assign inbar[124] = ~in[124];
  assign inbar[125] = ~in[125];
  assign inbar[126] = ~in[126];
  assign inbar[127] = ~in[127];
  assign inbar[128] = ~in[128];
  assign inbar[129] = ~in[129];
  assign inbar[130] = ~in[130];
  assign inbar[131] = ~in[131];
  assign inbar[132] = ~in[132];
  assign inbar[133] = ~in[133];
  assign inbar[134] = ~in[134];
  assign inbar[135] = ~in[135];
  assign inbar[136] = ~in[136];
  assign inbar[137] = ~in[137];
  assign inbar[138] = ~in[138];
  assign inbar[139] = ~in[139];
  assign inbar[140] = ~in[140];
  assign inbar[141] = ~in[141];
  assign inbar[142] = ~in[142];
  assign inbar[143] = ~in[143];
  assign inbar[144] = ~in[144];
  assign inbar[145] = ~in[145];
  assign inbar[146] = ~in[146];
  assign inbar[147] = ~in[147];
  assign inbar[148] = ~in[148];
  assign inbar[149] = ~in[149];
  assign inbar[150] = ~in[150];
  assign inbar[151] = ~in[151];
  assign inbar[152] = ~in[152];
  assign inbar[153] = ~in[153];
  assign inbar[154] = ~in[154];
  assign inbar[155] = ~in[155];
  assign inbar[156] = ~in[156];
  assign inbar[157] = ~in[157];
  assign inbar[158] = ~in[158];
  assign inbar[159] = ~in[159];
  assign inbar[160] = ~in[160];
  assign inbar[161] = ~in[161];
  assign inbar[162] = ~in[162];
  assign inbar[163] = ~in[163];
  assign inbar[164] = ~in[164];
  assign inbar[165] = ~in[165];
  assign inbar[166] = ~in[166];
  assign inbar[167] = ~in[167];
  assign inbar[168] = ~in[168];
  assign inbar[169] = ~in[169];
  assign inbar[170] = ~in[170];
  assign inbar[171] = ~in[171];
  assign inbar[172] = ~in[172];
  assign inbar[173] = ~in[173];
  assign inbar[174] = ~in[174];
  assign inbar[175] = ~in[175];
  assign inbar[176] = ~in[176];
  assign inbar[177] = ~in[177];
  assign inbar[178] = ~in[178];
  assign inbar[179] = ~in[179];
  assign inbar[180] = ~in[180];
  assign inbar[181] = ~in[181];
  assign inbar[182] = ~in[182];
  assign inbar[183] = ~in[183];
  assign inbar[184] = ~in[184];
  assign inbar[185] = ~in[185];
  assign inbar[186] = ~in[186];
  assign inbar[187] = ~in[187];
  assign inbar[188] = ~in[188];
  assign inbar[189] = ~in[189];
  assign inbar[190] = ~in[190];
  assign inbar[191] = ~in[191];
  assign inbar[192] = ~in[192];
  assign inbar[193] = ~in[193];
  assign inbar[194] = ~in[194];
  assign inbar[195] = ~in[195];
  assign inbar[196] = ~in[196];
  assign inbar[197] = ~in[197];
  assign inbar[198] = ~in[198];
  assign inbar[199] = ~in[199];
  assign inbar[200] = ~in[200];
  assign inbar[201] = ~in[201];
  assign inbar[202] = ~in[202];
  assign inbar[203] = ~in[203];
  assign inbar[204] = ~in[204];
  assign inbar[205] = ~in[205];
  assign inbar[206] = ~in[206];
  assign inbar[207] = ~in[207];
  assign inbar[208] = ~in[208];
  assign inbar[209] = ~in[209];
  assign inbar[210] = ~in[210];
  assign inbar[211] = ~in[211];
  assign inbar[212] = ~in[212];
  assign inbar[213] = ~in[213];
  assign inbar[214] = ~in[214];
  assign inbar[215] = ~in[215];
  assign inbar[216] = ~in[216];
  assign inbar[217] = ~in[217];
  assign inbar[218] = ~in[218];
  assign inbar[219] = ~in[219];
  assign inbar[220] = ~in[220];
  assign inbar[221] = ~in[221];
  assign inbar[222] = ~in[222];
  assign inbar[223] = ~in[223];
  assign inbar[224] = ~in[224];
  assign inbar[225] = ~in[225];
  assign inbar[226] = ~in[226];
  assign inbar[227] = ~in[227];
  assign inbar[228] = ~in[228];
  assign inbar[229] = ~in[229];
  assign inbar[230] = ~in[230];
  assign inbar[231] = ~in[231];
  assign inbar[232] = ~in[232];
  assign inbar[233] = ~in[233];
  assign inbar[234] = ~in[234];
  assign inbar[235] = ~in[235];
  assign inbar[236] = ~in[236];
  assign inbar[237] = ~in[237];
  assign inbar[238] = ~in[238];
  assign inbar[239] = ~in[239];
  assign inbar[240] = ~in[240];
  assign inbar[241] = ~in[241];
  assign inbar[242] = ~in[242];
  assign inbar[243] = ~in[243];
  assign inbar[244] = ~in[244];
  assign inbar[245] = ~in[245];
  assign inbar[246] = ~in[246];
  assign inbar[247] = ~in[247];
  assign inbar[248] = ~in[248];
  assign inbar[249] = ~in[249];
  assign inbar[250] = ~in[250];
  assign inbar[251] = ~in[251];
  assign inbar[252] = ~in[252];
  assign inbar[253] = ~in[253];
  assign inbar[254] = ~in[254];
  assign inbar[255] = ~in[255];
//input_done

  output wire [7:0] out;
  wire [7:0] outbar;
//output_done

  wire in_81;
  wire in_80;
  wire in_79;
  wire in_78;
  wire in_77;
  wire in_76;
  wire in_75;
  wire in_74;
  wire in_73;
  wire in_72;
  wire in_71;
  wire in_70;
  wire in_69;
  wire in_68;
  wire in_67;
  wire in_66;
  wire in_65;
  wire in_64;
  wire in_63;
  wire in_62;
  wire in_61;
  wire in_60;
  wire in_59;
  wire in_58;
  wire in_57;
  wire in_56;
  wire in_55;
  wire in_54;
  wire in_53;
  wire in_52;
  wire in_51;
  wire in_50;
  wire in_49;
  wire in_48;
  wire in_47;
  wire in_46;
  wire in_45;
  wire in_44;
  wire in_43;
  wire in_42;
  wire in_41;
  wire in_40;
  wire in_39;
  wire in_38;
  wire in_37;
  wire in_36;
  wire in_35;
  wire in_34;
  wire in_33;
  wire in_32;
  wire in_31;
  wire in_30;
  wire in_29;
  wire in_28;
  wire in_27;
  wire in_26;
  wire in_25;
  wire in_24;
  wire in_23;
  wire in_22;
  wire in_21;
  wire in_20;
  wire in_19;
  wire in_18;
  wire in_17;
  wire in_16;
  wire in_15;
  wire in_14;
  wire in_13;
  wire in_12;
  wire in_11;
  wire in_10;
  wire in_9;
  wire in_8;
  wire in_7;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_3;
  wire in_2;
  wire in_1;
  wire in_0;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire in_81bar;
  wire in_80bar;
  wire in_79bar;
  wire in_78bar;
  wire in_77bar;
  wire in_76bar;
  wire in_75bar;
  wire in_74bar;
  wire in_73bar;
  wire in_72bar;
  wire in_71bar;
  wire in_70bar;
  wire in_69bar;
  wire in_68bar;
  wire in_67bar;
  wire in_66bar;
  wire in_65bar;
  wire in_64bar;
  wire in_63bar;
  wire in_62bar;
  wire in_61bar;
  wire in_60bar;
  wire in_59bar;
  wire in_58bar;
  wire in_57bar;
  wire in_56bar;
  wire in_55bar;
  wire in_54bar;
  wire in_53bar;
  wire in_52bar;
  wire in_51bar;
  wire in_50bar;
  wire in_49bar;
  wire in_48bar;
  wire in_47bar;
  wire in_46bar;
  wire in_45bar;
  wire in_44bar;
  wire in_43bar;
  wire in_42bar;
  wire in_41bar;
  wire in_40bar;
  wire in_39bar;
  wire in_38bar;
  wire in_37bar;
  wire in_36bar;
  wire in_35bar;
  wire in_34bar;
  wire in_33bar;
  wire in_32bar;
  wire in_31bar;
  wire in_30bar;
  wire in_29bar;
  wire in_28bar;
  wire in_27bar;
  wire in_26bar;
  wire in_25bar;
  wire in_24bar;
  wire in_23bar;
  wire in_22bar;
  wire in_21bar;
  wire in_20bar;
  wire in_19bar;
  wire in_18bar;
  wire in_17bar;
  wire in_16bar;
  wire in_15bar;
  wire in_14bar;
  wire in_13bar;
  wire in_12bar;
  wire in_11bar;
  wire in_10bar;
  wire in_9bar;
  wire in_8bar;
  wire in_7bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_3bar;
  wire in_2bar;
  wire in_1bar;
  wire in_0bar;
  wire n487bar;
  wire n488bar;
  wire n489bar;
  wire n490bar;
  wire n491bar;
  wire n492bar;
  wire n493bar;
  wire n494bar;
  wire n495bar;
  wire n496bar;
  wire n497bar;
  wire n498bar;
  wire n499bar;
  wire n500bar;
  wire n501bar;
  wire n502bar;
  wire n503bar;
  wire n504bar;
  wire n505bar;
  wire n506bar;
  wire n507bar;
  wire n508bar;
  wire n509bar;
  wire n510bar;
  wire n511bar;
  wire n512bar;
  wire n513bar;
  wire n514bar;
  wire n515bar;
  wire n516bar;
  wire n517bar;
  wire n518bar;
  wire n519bar;
  wire n520bar;
  wire n521bar;
  wire n522bar;
  wire n523bar;
  wire n524bar;
  wire n525bar;
  wire n526bar;
  wire n527bar;
  wire n528bar;
  wire n529bar;
  wire n530bar;
  wire n531bar;
  wire n532bar;
  wire n533bar;
  wire n534bar;
  wire n535bar;
  wire n536bar;
  wire n537bar;
  wire n538bar;
  wire n539bar;
  wire n540bar;
  wire n541bar;
  wire n542bar;
  wire n543bar;
  wire n544bar;
  wire n545bar;
  wire n546bar;
  wire n547bar;
  wire n548bar;
  wire n549bar;
  wire n550bar;
  wire n551bar;
  wire n552bar;
  wire n553bar;
  wire n554bar;
  wire n555bar;
  wire n556bar;
  wire n557bar;
  wire n558bar;
  wire n559bar;
  wire n560bar;
  wire n561bar;
  wire n562bar;
  wire n563bar;
  wire n564bar;
  wire n565bar;
  wire n566bar;
  wire n567bar;
  wire n568bar;
  wire n569bar;
  wire n570bar;
  wire n571bar;
  wire n572bar;
  wire n573bar;
  wire n574bar;
  wire n575bar;
  wire n576bar;
  wire n577bar;
  wire n578bar;
  wire n579bar;
  wire n580bar;
  wire n581bar;
  wire n582bar;
  wire n583bar;
  wire n584bar;
  wire n585bar;
  wire n586bar;
  wire n587bar;
  wire n588bar;
  wire n589bar;
  wire n590bar;
  wire n591bar;
  wire n592bar;
  wire n593bar;
  wire n594bar;
  wire n595bar;
  wire n596bar;
  wire n597bar;
  wire n598bar;
  wire n599bar;
  wire n600bar;
  wire n601bar;
  wire n602bar;
  wire n603bar;
  wire n604bar;
  wire n605bar;
  wire n606bar;
  wire n607bar;
  wire n608bar;
  wire n609bar;
  wire n610bar;
  wire n611bar;
  wire n612bar;
  wire n613bar;
  wire n614bar;
  wire n615bar;
  wire n616bar;
  wire n617bar;
  wire n618bar;
  wire n619bar;
  wire n620bar;
  wire n621bar;
  wire n622bar;
  wire n623bar;
  wire n624bar;
  wire n625bar;
  wire n626bar;
  wire n627bar;
  wire n628bar;
  wire n629bar;
  wire n630bar;
  wire n631bar;
  wire n632bar;
  wire n633bar;
  wire n634bar;
  wire n635bar;
  wire n636bar;
  wire n637bar;
  wire n638bar;
  wire n639bar;
  wire n640bar;
  wire n641bar;
  wire n642bar;
  wire n643bar;
  wire n644bar;
  wire n645bar;
  wire n646bar;
  wire n647bar;
  wire n648bar;
  wire n649bar;
  wire n650bar;
  wire n651bar;
  wire n652bar;
  wire n653bar;
  wire n654bar;
  wire n655bar;
  wire n656bar;
  wire n657bar;
  wire n658bar;
  wire n659bar;
  wire n660bar;
  wire n661bar;
  wire n662bar;
  wire n663bar;
  wire n664bar;
  wire n665bar;
  wire n666bar;
  wire n667bar;
  wire n668bar;
  wire n669bar;
  wire n670bar;
  wire n671bar;
  wire n672bar;
  wire n673bar;
  wire n674bar;
  wire n675bar;
  wire n676bar;
  wire n677bar;
  wire n678bar;
  wire n679bar;
  wire n680bar;
  wire n681bar;
  wire n682bar;
  wire n683bar;
  wire n684bar;
  wire n685bar;
  wire n686bar;
  wire n687bar;
  wire n688bar;
  wire n689bar;
  wire n690bar;
  wire n691bar;
  wire n692bar;
  wire n693bar;
  wire n694bar;
  wire n695bar;
  wire n696bar;
  wire n697bar;
  wire n698bar;
  wire n699bar;
  wire n700bar;
  wire n701bar;
  wire n702bar;
  wire n703bar;
  wire n704bar;
  wire n705bar;
  wire n706bar;
  wire n707bar;
  wire n708bar;
  wire n709bar;
  wire n710bar;
  wire n711bar;
  wire n712bar;
  wire n713bar;
  wire n714bar;
  wire n715bar;
  wire n716bar;
  wire n717bar;
  wire n718bar;
  wire n719bar;
  wire n720bar;
  wire n721bar;
  wire n722bar;
  wire n723bar;
  wire n724bar;
  wire n725bar;
  wire n726bar;
  wire n727bar;
  wire n728bar;
  wire n729bar;
  wire n730bar;
  wire n731bar;
  wire n732bar;
  wire n733bar;
  wire n734bar;
  wire n735bar;
  wire n736bar;
  wire n737bar;
  wire n738bar;
  wire n739bar;
  wire n740bar;
  wire n741bar;
  wire n742bar;
  wire n743bar;
  wire n744bar;
  wire n745bar;
  wire n746bar;
  wire n747bar;
  wire n748bar;
  wire n749bar;
  wire n750bar;
  wire n751bar;
  wire n752bar;
  wire n753bar;
  wire n754bar;
  wire n755bar;
  wire n756bar;
  wire n757bar;
  wire n758bar;
  wire n759bar;
  wire n760bar;
  wire n761bar;
  wire n762bar;
  wire n763bar;
  wire n764bar;
  wire n765bar;
  wire n766bar;
  wire n767bar;
  wire n768bar;
  wire n769bar;
  wire n770bar;
  wire n771bar;
  wire n772bar;
  wire n773bar;
  wire n774bar;
  wire n775bar;
  wire n776bar;
  wire n777bar;
  wire n778bar;
  wire n779bar;
  wire n780bar;
  wire n781bar;
  wire n782bar;
  wire n783bar;
  wire n784bar;
  wire n785bar;
  wire n786bar;
  wire n787bar;
  wire n788bar;
  wire n789bar;
  wire n790bar;
  wire n791bar;
  wire n792bar;
  wire n793bar;
  wire n794bar;
  wire n795bar;
  wire n796bar;
  wire n797bar;
  wire n798bar;
  wire n799bar;
  wire n800bar;
  wire n801bar;
  wire n802bar;
  wire n803bar;
  wire n804bar;
  wire n805bar;
  wire n806bar;
  wire n807bar;
  wire n808bar;
  wire n809bar;
  wire n810bar;
  wire n811bar;
  wire n812bar;
  wire n813bar;
  wire n814bar;
  wire n815bar;
  wire n816bar;
  wire n817bar;
  wire n818bar;
  wire n819bar;
  wire n820bar;
  wire n821bar;
  wire n822bar;
  wire n823bar;
  wire n824bar;
  wire n825bar;
  wire n826bar;
  wire n827bar;
  wire n828bar;
  wire n829bar;
  wire n830bar;
  wire n831bar;
  wire n832bar;
  wire n833bar;
  wire n834bar;
  wire n835bar;
  wire n836bar;
  wire n837bar;
  wire n838bar;
  wire n839bar;
  wire n840bar;
  wire n841bar;
  wire n842bar;
  wire n843bar;
  wire n844bar;
  wire n845bar;
  wire n846bar;
  wire n847bar;
  wire n848bar;
  wire n849bar;
  wire n850bar;
  wire n851bar;
  wire n852bar;
  wire n853bar;
  wire n854bar;
  wire n855bar;
  wire n856bar;
  wire n857bar;
  wire n858bar;
  wire n859bar;
  wire n860bar;
  wire n861bar;
  wire n862bar;
  wire n863bar;
  wire n864bar;
  wire n865bar;
  wire n866bar;
  wire n867bar;
  wire n868bar;
  wire n869bar;
  wire n870bar;
  wire n871bar;
  wire n872bar;
  wire n873bar;
  wire n874bar;
  wire n875bar;
  wire n876bar;
  wire n877bar;
  wire n878bar;
  wire n879bar;
  wire n880bar;
  wire n881bar;
  wire n882bar;
  wire n883bar;
  wire n884bar;
  wire n885bar;
  wire n886bar;
  wire n887bar;
  wire n888bar;
  wire n889bar;
  wire n890bar;
  wire n891bar;
  wire n892bar;
  wire n893bar;
  wire n894bar;
  wire n895bar;
  wire n896bar;
  wire n897bar;
  wire n898bar;
  wire n899bar;
  wire n900bar;
  wire n901bar;
  wire n902bar;
  wire n903bar;
  wire n904bar;
  wire n905bar;
  wire n906bar;
  wire n907bar;
  wire n908bar;
  wire n909bar;
  wire n910bar;
  wire n911bar;
  wire n912bar;
  wire n913bar;
  wire n914bar;
  wire n915bar;
  wire n916bar;
  wire n917bar;
  wire n918bar;
  wire n919bar;
  wire n920bar;
  wire n921bar;
  wire n922bar;
  wire n923bar;
  wire n924bar;
  wire n925bar;
  wire n926bar;
  wire n927bar;
  wire n928bar;
  wire n929bar;
  wire n930bar;
  wire n931bar;
  wire n932bar;
  wire n933bar;
  wire n934bar;
  wire n935bar;
  wire n936bar;
  wire n937bar;
  wire n938bar;
  wire n939bar;
  wire n940bar;
  wire n941bar;
  wire n942bar;
  wire n943bar;
  wire n944bar;
  wire n945bar;
  wire n946bar;
  wire n947bar;
  wire n948bar;
  wire n949bar;
  wire n950bar;
  wire n951bar;
  wire n952bar;
  wire n953bar;
  wire n954bar;
  wire n955bar;
  wire n956bar;
  wire n957bar;
  wire n958bar;
  wire n959bar;
  wire n960bar;
  wire n961bar;
  wire n962bar;
  wire n963bar;
  wire n964bar;
  wire n965bar;
  wire n966bar;
  wire n967bar;
  wire n968bar;
  wire n969bar;
  wire n970bar;
  wire n971bar;
  wire n972bar;
//wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];
  //OR U1
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1 (
    .O(out[7]),
    .I0(n972),
    .I1(n971)
  );
  //AND U1bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1bar (
    .O(outbar[7]),
    .I0(n972bar),
    .I1(n971bar)
  );
  //OR U2
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2 (
    .O(n971),
    .I0(n970),
    .I1(n969)
  );
  //AND U2bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2bar (
    .O(n971bar),
    .I0(n970bar),
    .I1(n969bar)
  );
  //OR U3
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3 (
    .O(n969),
    .I0(n968),
    .I1(n967)
  );
  //AND U3bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3bar (
    .O(n969bar),
    .I0(n968bar),
    .I1(n967bar)
  );
  //OR U4
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4 (
    .O(n967),
    .I0(n966),
    .I1(n965)
  );
  //AND U4bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4bar (
    .O(n967bar),
    .I0(n966bar),
    .I1(n965bar)
  );
  //OR U5
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5 (
    .O(n968),
    .I0(n964),
    .I1(n963)
  );
  //AND U5bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5bar (
    .O(n968bar),
    .I0(n964bar),
    .I1(n963bar)
  );
  //OR U6
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6 (
    .O(n963),
    .I0(in[116]),
    .I1(n962)
  );
  //AND U6bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6bar (
    .O(n963bar),
    .I0(inbar[116]),
    .I1(n962bar)
  );
  //OR U7
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7 (
    .O(n970),
    .I0(n961),
    .I1(n960)
  );
  //AND U7bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7bar (
    .O(n970bar),
    .I0(n961bar),
    .I1(n960bar)
  );
  //OR U8
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8 (
    .O(n960),
    .I0(in[150]),
    .I1(in[127])
  );
  //AND U8bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8bar (
    .O(n960bar),
    .I0(inbar[150]),
    .I1(inbar[127])
  );
  //OR U9
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9 (
    .O(n961),
    .I0(in[160]),
    .I1(n959)
  );
  //AND U9bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9bar (
    .O(n961bar),
    .I0(inbar[160]),
    .I1(n959bar)
  );
  //OR U10
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10 (
    .O(n959),
    .I0(in[252]),
    .I1(in[168])
  );
  //AND U10bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10bar (
    .O(n959bar),
    .I0(inbar[252]),
    .I1(inbar[168])
  );
  //OR U11
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11 (
    .O(n972),
    .I0(n958),
    .I1(n957)
  );
  //AND U11bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11bar (
    .O(n972bar),
    .I0(n958bar),
    .I1(n957bar)
  );
  //OR U12
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12 (
    .O(n957),
    .I0(n956),
    .I1(n955)
  );
  //AND U12bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12bar (
    .O(n957bar),
    .I0(n956bar),
    .I1(n955bar)
  );
  //OR U13
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13 (
    .O(n955),
    .I0(in_17),
    .I1(in[96])
  );
  //AND U13bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13bar (
    .O(n955bar),
    .I0(in_17bar),
    .I1(inbar[96])
  );
  //OR U14
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14 (
    .O(n956),
    .I0(in_23),
    .I1(n954)
  );
  //AND U14bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14bar (
    .O(n956bar),
    .I0(in_23bar),
    .I1(n954bar)
  );
  //OR U15
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15 (
    .O(n954),
    .I0(in_31),
    .I1(in_26)
  );
  //AND U15bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15bar (
    .O(n954bar),
    .I0(in_31bar),
    .I1(in_26bar)
  );
  //OR U16
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16 (
    .O(n958),
    .I0(n953),
    .I1(n952)
  );
  //AND U16bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16bar (
    .O(n958bar),
    .I0(n953bar),
    .I1(n952bar)
  );
  //OR U17
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U17 (
    .O(n952),
    .I0(in_58),
    .I1(in_4)
  );
  //AND U17bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U17bar (
    .O(n952bar),
    .I0(in_58bar),
    .I1(in_4bar)
  );
  //OR U18
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U18 (
    .O(n953),
    .I0(in_59),
    .I1(n951)
  );
  //AND U18bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U18bar (
    .O(n953bar),
    .I0(in_59bar),
    .I1(n951bar)
  );
  //OR U19
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U19 (
    .O(n951),
    .I0(in_71),
    .I1(in_62)
  );
  //AND U19bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U19bar (
    .O(n951bar),
    .I0(in_71bar),
    .I1(in_62bar)
  );
  //OR U20
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U20 (
    .O(out[6]),
    .I0(n950),
    .I1(n949)
  );
  //AND U20bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U20bar (
    .O(outbar[6]),
    .I0(n950bar),
    .I1(n949bar)
  );
  //OR U21
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U21 (
    .O(n949),
    .I0(n948),
    .I1(n947)
  );
  //AND U21bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U21bar (
    .O(n949bar),
    .I0(n948bar),
    .I1(n947bar)
  );
  //OR U22
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U22 (
    .O(n947),
    .I0(n946),
    .I1(n945)
  );
  //AND U22bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U22bar (
    .O(n947bar),
    .I0(n946bar),
    .I1(n945bar)
  );
  //OR U23
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U23 (
    .O(n945),
    .I0(n944),
    .I1(n943)
  );
  //AND U23bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U23bar (
    .O(n945bar),
    .I0(n944bar),
    .I1(n943bar)
  );
  //OR U24
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U24 (
    .O(n946),
    .I0(n942),
    .I1(n941)
  );
  //AND U24bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U24bar (
    .O(n946bar),
    .I0(n942bar),
    .I1(n941bar)
  );
  //OR U25
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U25 (
    .O(n941),
    .I0(in[101]),
    .I1(n940)
  );
  //AND U25bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U25bar (
    .O(n941bar),
    .I0(inbar[101]),
    .I1(n940bar)
  );
  //OR U26
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U26 (
    .O(n948),
    .I0(n939),
    .I1(n938)
  );
  //AND U26bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U26bar (
    .O(n948bar),
    .I0(n939bar),
    .I1(n938bar)
  );
  //OR U27
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U27 (
    .O(n938),
    .I0(in[114]),
    .I1(in[104])
  );
  //AND U27bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U27bar (
    .O(n938bar),
    .I0(inbar[114]),
    .I1(inbar[104])
  );
  //OR U28
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U28 (
    .O(n939),
    .I0(in[128]),
    .I1(n937)
  );
  //AND U28bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U28bar (
    .O(n939bar),
    .I0(inbar[128]),
    .I1(n937bar)
  );
  //OR U29
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U29 (
    .O(n937),
    .I0(in[136]),
    .I1(in[134])
  );
  //AND U29bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U29bar (
    .O(n937bar),
    .I0(inbar[136]),
    .I1(inbar[134])
  );
  //OR U30
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U30 (
    .O(n950),
    .I0(n936),
    .I1(n935)
  );
  //AND U30bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U30bar (
    .O(n950bar),
    .I0(n936bar),
    .I1(n935bar)
  );
  //OR U31
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U31 (
    .O(n935),
    .I0(n934),
    .I1(n933)
  );
  //AND U31bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U31bar (
    .O(n935bar),
    .I0(n934bar),
    .I1(n933bar)
  );
  //OR U32
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U32 (
    .O(n933),
    .I0(in[177]),
    .I1(in[164])
  );
  //AND U32bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U32bar (
    .O(n933bar),
    .I0(inbar[177]),
    .I1(inbar[164])
  );
  //OR U33
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U33 (
    .O(n934),
    .I0(in[212]),
    .I1(n932)
  );
  //AND U33bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U33bar (
    .O(n934bar),
    .I0(inbar[212]),
    .I1(n932bar)
  );
  //OR U34
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U34 (
    .O(n932),
    .I0(in[248]),
    .I1(in[221])
  );
  //AND U34bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U34bar (
    .O(n932bar),
    .I0(inbar[248]),
    .I1(inbar[221])
  );
  //OR U35
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U35 (
    .O(n936),
    .I0(n931),
    .I1(n930)
  );
  //AND U35bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U35bar (
    .O(n936bar),
    .I0(n931bar),
    .I1(n930bar)
  );
  //OR U36
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U36 (
    .O(n930),
    .I0(in_18),
    .I1(in[93])
  );
  //AND U36bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U36bar (
    .O(n930bar),
    .I0(in_18bar),
    .I1(inbar[93])
  );
  //OR U37
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U37 (
    .O(n931),
    .I0(in_31),
    .I1(n929)
  );
  //AND U37bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U37bar (
    .O(n931bar),
    .I0(in_31bar),
    .I1(n929bar)
  );
  //OR U38
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U38 (
    .O(n929),
    .I0(in_7),
    .I1(in_39)
  );
  //AND U38bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U38bar (
    .O(n929bar),
    .I0(in_7bar),
    .I1(in_39bar)
  );
  //OR U39
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U39 (
    .O(out[5]),
    .I0(n928),
    .I1(n927)
  );
  //AND U39bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U39bar (
    .O(outbar[5]),
    .I0(n928bar),
    .I1(n927bar)
  );
  //OR U40
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U40 (
    .O(n927),
    .I0(n926),
    .I1(n925)
  );
  //AND U40bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U40bar (
    .O(n927bar),
    .I0(n926bar),
    .I1(n925bar)
  );
  //OR U41
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U41 (
    .O(n925),
    .I0(n924),
    .I1(n923)
  );
  //AND U41bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U41bar (
    .O(n925bar),
    .I0(n924bar),
    .I1(n923bar)
  );
  //OR U42
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U42 (
    .O(n923),
    .I0(n922),
    .I1(n921)
  );
  //AND U42bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U42bar (
    .O(n923bar),
    .I0(n922bar),
    .I1(n921bar)
  );
  //OR U43
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U43 (
    .O(n924),
    .I0(n940),
    .I1(n920)
  );
  //AND U43bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U43bar (
    .O(n924bar),
    .I0(n940bar),
    .I1(n920bar)
  );
  //OR U44
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U44 (
    .O(n920),
    .I0(in[111]),
    .I1(n919)
  );
  //AND U44bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U44bar (
    .O(n920bar),
    .I0(inbar[111]),
    .I1(n919bar)
  );
  //OR U45
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U45 (
    .O(n940),
    .I0(n918),
    .I1(n917)
  );
  //AND U45bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U45bar (
    .O(n940bar),
    .I0(n918bar),
    .I1(n917bar)
  );
  //OR U46
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U46 (
    .O(n917),
    .I0(n916),
    .I1(n915)
  );
  //AND U46bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U46bar (
    .O(n917bar),
    .I0(n916bar),
    .I1(n915bar)
  );
  //OR U47
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U47 (
    .O(n915),
    .I0(n914),
    .I1(n913)
  );
  //AND U47bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U47bar (
    .O(n915bar),
    .I0(n914bar),
    .I1(n913bar)
  );
  //OR U48
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U48 (
    .O(n913),
    .I0(in[140]),
    .I1(in[131])
  );
  //AND U48bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U48bar (
    .O(n913bar),
    .I0(inbar[140]),
    .I1(inbar[131])
  );
  //OR U49
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U49 (
    .O(n914),
    .I0(in[160]),
    .I1(in[144])
  );
  //AND U49bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U49bar (
    .O(n914bar),
    .I0(inbar[160]),
    .I1(inbar[144])
  );
  //OR U50
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U50 (
    .O(n916),
    .I0(n912),
    .I1(n911)
  );
  //AND U50bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U50bar (
    .O(n916bar),
    .I0(n912bar),
    .I1(n911bar)
  );
  //OR U51
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U51 (
    .O(n911),
    .I0(in[179]),
    .I1(in[174])
  );
  //AND U51bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U51bar (
    .O(n911bar),
    .I0(inbar[179]),
    .I1(inbar[174])
  );
  //OR U52
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U52 (
    .O(n912),
    .I0(in[188]),
    .I1(in[184])
  );
  //AND U52bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U52bar (
    .O(n912bar),
    .I0(inbar[188]),
    .I1(inbar[184])
  );
  //OR U53
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U53 (
    .O(n918),
    .I0(n910),
    .I1(n909)
  );
  //AND U53bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U53bar (
    .O(n918bar),
    .I0(n910bar),
    .I1(n909bar)
  );
  //OR U54
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U54 (
    .O(n909),
    .I0(n908),
    .I1(n907)
  );
  //AND U54bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U54bar (
    .O(n909bar),
    .I0(n908bar),
    .I1(n907bar)
  );
  //OR U55
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U55 (
    .O(n907),
    .I0(in[216]),
    .I1(in[200])
  );
  //AND U55bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U55bar (
    .O(n907bar),
    .I0(inbar[216]),
    .I1(inbar[200])
  );
  //OR U56
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U56 (
    .O(n908),
    .I0(in[228]),
    .I1(in[224])
  );
  //AND U56bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U56bar (
    .O(n908bar),
    .I0(inbar[228]),
    .I1(inbar[224])
  );
  //OR U57
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U57 (
    .O(n910),
    .I0(n906),
    .I1(n905)
  );
  //AND U57bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U57bar (
    .O(n910bar),
    .I0(n906bar),
    .I1(n905bar)
  );
  //OR U58
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U58 (
    .O(n905),
    .I0(in[247]),
    .I1(in[235])
  );
  //AND U58bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U58bar (
    .O(n905bar),
    .I0(inbar[247]),
    .I1(inbar[235])
  );
  //OR U59
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U59 (
    .O(n906),
    .I0(in_42),
    .I1(in[83])
  );
  //AND U59bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U59bar (
    .O(n906bar),
    .I0(in_42bar),
    .I1(inbar[83])
  );
  //OR U60
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U60 (
    .O(n926),
    .I0(n904),
    .I1(n903)
  );
  //AND U60bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U60bar (
    .O(n926bar),
    .I0(n904bar),
    .I1(n903bar)
  );
  //OR U61
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U61 (
    .O(n903),
    .I0(in[166]),
    .I1(in[123])
  );
  //AND U61bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U61bar (
    .O(n903bar),
    .I0(inbar[166]),
    .I1(inbar[123])
  );
  //OR U62
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U62 (
    .O(n904),
    .I0(in[170]),
    .I1(n902)
  );
  //AND U62bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U62bar (
    .O(n904bar),
    .I0(inbar[170]),
    .I1(n902bar)
  );
  //OR U63
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U63 (
    .O(n902),
    .I0(in[194]),
    .I1(in[183])
  );
  //AND U63bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U63bar (
    .O(n902bar),
    .I0(inbar[194]),
    .I1(inbar[183])
  );
  //OR U64
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U64 (
    .O(n928),
    .I0(n901),
    .I1(n900)
  );
  //AND U64bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U64bar (
    .O(n928bar),
    .I0(n901bar),
    .I1(n900bar)
  );
  //OR U65
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U65 (
    .O(n900),
    .I0(n899),
    .I1(n898)
  );
  //AND U65bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U65bar (
    .O(n900bar),
    .I0(n899bar),
    .I1(n898bar)
  );
  //OR U66
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U66 (
    .O(n898),
    .I0(in[241]),
    .I1(in[238])
  );
  //AND U66bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U66bar (
    .O(n898bar),
    .I0(inbar[241]),
    .I1(inbar[238])
  );
  //OR U67
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U67 (
    .O(n899),
    .I0(in[250]),
    .I1(n897)
  );
  //AND U67bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U67bar (
    .O(n899bar),
    .I0(inbar[250]),
    .I1(n897bar)
  );
  //OR U68
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U68 (
    .O(n897),
    .I0(in_24),
    .I1(in[84])
  );
  //AND U68bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U68bar (
    .O(n897bar),
    .I0(in_24bar),
    .I1(inbar[84])
  );
  //OR U69
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U69 (
    .O(n901),
    .I0(n896),
    .I1(n895)
  );
  //AND U69bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U69bar (
    .O(n901bar),
    .I0(n896bar),
    .I1(n895bar)
  );
  //OR U70
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U70 (
    .O(n895),
    .I0(in_41),
    .I1(in_29)
  );
  //AND U70bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U70bar (
    .O(n895bar),
    .I0(in_41bar),
    .I1(in_29bar)
  );
  //OR U71
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U71 (
    .O(n896),
    .I0(in_66),
    .I1(n894)
  );
  //AND U71bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U71bar (
    .O(n896bar),
    .I0(in_66bar),
    .I1(n894bar)
  );
  //OR U72
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U72 (
    .O(n894),
    .I0(in_76),
    .I1(in_71)
  );
  //AND U72bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U72bar (
    .O(n894bar),
    .I0(in_76bar),
    .I1(in_71bar)
  );
  //OR U73
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U73 (
    .O(out[4]),
    .I0(n893),
    .I1(n892)
  );
  //AND U73bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U73bar (
    .O(outbar[4]),
    .I0(n893bar),
    .I1(n892bar)
  );
  //OR U74
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U74 (
    .O(n892),
    .I0(n891),
    .I1(n890)
  );
  //AND U74bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U74bar (
    .O(n892bar),
    .I0(n891bar),
    .I1(n890bar)
  );
  //OR U75
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U75 (
    .O(n890),
    .I0(n889),
    .I1(n888)
  );
  //AND U75bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U75bar (
    .O(n890bar),
    .I0(n889bar),
    .I1(n888bar)
  );
  //OR U76
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U76 (
    .O(n888),
    .I0(n922),
    .I1(n887)
  );
  //AND U76bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U76bar (
    .O(n888bar),
    .I0(n922bar),
    .I1(n887bar)
  );
  //OR U77
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U77 (
    .O(n922),
    .I0(n886),
    .I1(n885)
  );
  //AND U77bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U77bar (
    .O(n922bar),
    .I0(n886bar),
    .I1(n885bar)
  );
  //OR U78
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U78 (
    .O(n885),
    .I0(n884),
    .I1(n883)
  );
  //AND U78bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U78bar (
    .O(n885bar),
    .I0(n884bar),
    .I1(n883bar)
  );
  //OR U79
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U79 (
    .O(n883),
    .I0(n882),
    .I1(n881)
  );
  //AND U79bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U79bar (
    .O(n883bar),
    .I0(n882bar),
    .I1(n881bar)
  );
  //OR U80
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U80 (
    .O(n881),
    .I0(in[118]),
    .I1(in[109])
  );
  //AND U80bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U80bar (
    .O(n881bar),
    .I0(inbar[118]),
    .I1(inbar[109])
  );
  //OR U81
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U81 (
    .O(n882),
    .I0(in[139]),
    .I1(in[120])
  );
  //AND U81bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U81bar (
    .O(n882bar),
    .I0(inbar[139]),
    .I1(inbar[120])
  );
  //OR U82
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U82 (
    .O(n884),
    .I0(n880),
    .I1(n879)
  );
  //AND U82bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U82bar (
    .O(n884bar),
    .I0(n880bar),
    .I1(n879bar)
  );
  //OR U83
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U83 (
    .O(n879),
    .I0(in[198]),
    .I1(in[154])
  );
  //AND U83bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U83bar (
    .O(n879bar),
    .I0(inbar[198]),
    .I1(inbar[154])
  );
  //OR U84
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U84 (
    .O(n880),
    .I0(in[210]),
    .I1(in[205])
  );
  //AND U84bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U84bar (
    .O(n880bar),
    .I0(inbar[210]),
    .I1(inbar[205])
  );
  //OR U85
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U85 (
    .O(n886),
    .I0(n878),
    .I1(n877)
  );
  //AND U85bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U85bar (
    .O(n886bar),
    .I0(n878bar),
    .I1(n877bar)
  );
  //OR U86
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U86 (
    .O(n877),
    .I0(n876),
    .I1(n875)
  );
  //AND U86bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U86bar (
    .O(n877bar),
    .I0(n876bar),
    .I1(n875bar)
  );
  //OR U87
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U87 (
    .O(n875),
    .I0(in[219]),
    .I1(in[217])
  );
  //AND U87bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U87bar (
    .O(n875bar),
    .I0(inbar[219]),
    .I1(inbar[217])
  );
  //OR U88
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U88 (
    .O(n876),
    .I0(in[86]),
    .I1(in[252])
  );
  //AND U88bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U88bar (
    .O(n876bar),
    .I0(inbar[86]),
    .I1(inbar[252])
  );
  //OR U89
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U89 (
    .O(n878),
    .I0(n874),
    .I1(n873)
  );
  //AND U89bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U89bar (
    .O(n878bar),
    .I0(n874bar),
    .I1(n873bar)
  );
  //OR U90
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U90 (
    .O(n873),
    .I0(in_40),
    .I1(in[91])
  );
  //AND U90bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U90bar (
    .O(n873bar),
    .I0(in_40bar),
    .I1(inbar[91])
  );
  //OR U91
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U91 (
    .O(n874),
    .I0(in_8),
    .I1(in_46)
  );
  //AND U91bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U91bar (
    .O(n874bar),
    .I0(in_8bar),
    .I1(in_46bar)
  );
  //OR U92
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U92 (
    .O(n889),
    .I0(n872),
    .I1(n871)
  );
  //AND U92bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U92bar (
    .O(n889bar),
    .I0(n872bar),
    .I1(n871bar)
  );
  //OR U93
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U93 (
    .O(n871),
    .I0(in[117]),
    .I1(n943)
  );
  //AND U93bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U93bar (
    .O(n871bar),
    .I0(inbar[117]),
    .I1(n943bar)
  );
  //OR U94
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U94 (
    .O(n943),
    .I0(n870),
    .I1(n869)
  );
  //AND U94bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U94bar (
    .O(n943bar),
    .I0(n870bar),
    .I1(n869bar)
  );
  //OR U95
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U95 (
    .O(n869),
    .I0(n868),
    .I1(n867)
  );
  //AND U95bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U95bar (
    .O(n869bar),
    .I0(n868bar),
    .I1(n867bar)
  );
  //OR U96
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U96 (
    .O(n867),
    .I0(n866),
    .I1(n865)
  );
  //AND U96bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U96bar (
    .O(n867bar),
    .I0(n866bar),
    .I1(n865bar)
  );
  //OR U97
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U97 (
    .O(n865),
    .I0(n864),
    .I1(n863)
  );
  //AND U97bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U97bar (
    .O(n865bar),
    .I0(n864bar),
    .I1(n863bar)
  );
  //OR U98
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U98 (
    .O(n866),
    .I0(in[108]),
    .I1(n919)
  );
  //AND U98bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U98bar (
    .O(n866bar),
    .I0(inbar[108]),
    .I1(n919bar)
  );
  //OR U99
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U99 (
    .O(n919),
    .I0(n862),
    .I1(n861)
  );
  //AND U99bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U99bar (
    .O(n919bar),
    .I0(n862bar),
    .I1(n861bar)
  );
  //OR U100
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U100 (
    .O(n861),
    .I0(n860),
    .I1(n859)
  );
  //AND U100bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U100bar (
    .O(n861bar),
    .I0(n860bar),
    .I1(n859bar)
  );
  //OR U101
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U101 (
    .O(n859),
    .I0(n858),
    .I1(n857)
  );
  //AND U101bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U101bar (
    .O(n859bar),
    .I0(n858bar),
    .I1(n857bar)
  );
  //OR U102
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U102 (
    .O(n857),
    .I0(in[119]),
    .I1(in[105])
  );
  //AND U102bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U102bar (
    .O(n857bar),
    .I0(inbar[119]),
    .I1(inbar[105])
  );
  //OR U103
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U103 (
    .O(n858),
    .I0(in[186]),
    .I1(in[175])
  );
  //AND U103bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U103bar (
    .O(n858bar),
    .I0(inbar[186]),
    .I1(inbar[175])
  );
  //OR U104
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U104 (
    .O(n860),
    .I0(n856),
    .I1(n855)
  );
  //AND U104bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U104bar (
    .O(n860bar),
    .I0(n856bar),
    .I1(n855bar)
  );
  //OR U105
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U105 (
    .O(n855),
    .I0(in[202]),
    .I1(in[193])
  );
  //AND U105bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U105bar (
    .O(n855bar),
    .I0(inbar[202]),
    .I1(inbar[193])
  );
  //OR U106
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U106 (
    .O(n856),
    .I0(in[225]),
    .I1(in[208])
  );
  //AND U106bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U106bar (
    .O(n856bar),
    .I0(inbar[225]),
    .I1(inbar[208])
  );
  //OR U107
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U107 (
    .O(n862),
    .I0(n854),
    .I1(n853)
  );
  //AND U107bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U107bar (
    .O(n862bar),
    .I0(n854bar),
    .I1(n853bar)
  );
  //OR U108
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U108 (
    .O(n853),
    .I0(n852),
    .I1(n851)
  );
  //AND U108bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U108bar (
    .O(n853bar),
    .I0(n852bar),
    .I1(n851bar)
  );
  //OR U109
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U109 (
    .O(n851),
    .I0(in_1),
    .I1(in[85])
  );
  //AND U109bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U109bar (
    .O(n851bar),
    .I0(in_1bar),
    .I1(inbar[85])
  );
  //OR U110
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U110 (
    .O(n852),
    .I0(in_23),
    .I1(in_19)
  );
  //AND U110bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U110bar (
    .O(n852bar),
    .I0(in_23bar),
    .I1(in_19bar)
  );
  //OR U111
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U111 (
    .O(n854),
    .I0(n850),
    .I1(n849)
  );
  //AND U111bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U111bar (
    .O(n854bar),
    .I0(n850bar),
    .I1(n849bar)
  );
  //OR U112
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U112 (
    .O(n849),
    .I0(in_43),
    .I1(in_33)
  );
  //AND U112bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U112bar (
    .O(n849bar),
    .I0(in_43bar),
    .I1(in_33bar)
  );
  //OR U113
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U113 (
    .O(n850),
    .I0(in_63),
    .I1(in_44)
  );
  //AND U113bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U113bar (
    .O(n850bar),
    .I0(in_63bar),
    .I1(in_44bar)
  );
  //OR U114
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U114 (
    .O(n868),
    .I0(n848),
    .I1(n847)
  );
  //AND U114bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U114bar (
    .O(n868bar),
    .I0(n848bar),
    .I1(n847bar)
  );
  //OR U115
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U115 (
    .O(n847),
    .I0(in[141]),
    .I1(in[112])
  );
  //AND U115bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U115bar (
    .O(n847bar),
    .I0(inbar[141]),
    .I1(inbar[112])
  );
  //OR U116
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U116 (
    .O(n848),
    .I0(in[147]),
    .I1(n846)
  );
  //AND U116bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U116bar (
    .O(n848bar),
    .I0(inbar[147]),
    .I1(n846bar)
  );
  //OR U117
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U117 (
    .O(n846),
    .I0(in[181]),
    .I1(in[167])
  );
  //AND U117bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U117bar (
    .O(n846bar),
    .I0(inbar[181]),
    .I1(inbar[167])
  );
  //OR U118
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U118 (
    .O(n870),
    .I0(n845),
    .I1(n844)
  );
  //AND U118bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U118bar (
    .O(n870bar),
    .I0(n845bar),
    .I1(n844bar)
  );
  //OR U119
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U119 (
    .O(n844),
    .I0(n843),
    .I1(n842)
  );
  //AND U119bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U119bar (
    .O(n844bar),
    .I0(n843bar),
    .I1(n842bar)
  );
  //OR U120
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U120 (
    .O(n842),
    .I0(in[229]),
    .I1(in[201])
  );
  //AND U120bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U120bar (
    .O(n842bar),
    .I0(inbar[229]),
    .I1(inbar[201])
  );
  //OR U121
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U121 (
    .O(n843),
    .I0(in[237]),
    .I1(n841)
  );
  //AND U121bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U121bar (
    .O(n843bar),
    .I0(inbar[237]),
    .I1(n841bar)
  );
  //OR U122
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U122 (
    .O(n841),
    .I0(in[94]),
    .I1(in[253])
  );
  //AND U122bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U122bar (
    .O(n841bar),
    .I0(inbar[94]),
    .I1(inbar[253])
  );
  //OR U123
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U123 (
    .O(n845),
    .I0(n840),
    .I1(n839)
  );
  //AND U123bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U123bar (
    .O(n845bar),
    .I0(n840bar),
    .I1(n839bar)
  );
  //OR U124
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U124 (
    .O(n839),
    .I0(in_21),
    .I1(in[96])
  );
  //AND U124bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U124bar (
    .O(n839bar),
    .I0(in_21bar),
    .I1(inbar[96])
  );
  //OR U125
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U125 (
    .O(n840),
    .I0(in_25),
    .I1(n838)
  );
  //AND U125bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U125bar (
    .O(n840bar),
    .I0(in_25bar),
    .I1(n838bar)
  );
  //OR U126
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U126 (
    .O(n838),
    .I0(in_81),
    .I1(in_45)
  );
  //AND U126bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U126bar (
    .O(n838bar),
    .I0(in_81bar),
    .I1(in_45bar)
  );
  //OR U127
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U127 (
    .O(n891),
    .I0(n837),
    .I1(n836)
  );
  //AND U127bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U127bar (
    .O(n891bar),
    .I0(n837bar),
    .I1(n836bar)
  );
  //OR U128
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U128 (
    .O(n836),
    .I0(in[142]),
    .I1(in[124])
  );
  //AND U128bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U128bar (
    .O(n836bar),
    .I0(inbar[142]),
    .I1(inbar[124])
  );
  //OR U129
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U129 (
    .O(n837),
    .I0(in[150]),
    .I1(n835)
  );
  //AND U129bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U129bar (
    .O(n837bar),
    .I0(inbar[150]),
    .I1(n835bar)
  );
  //OR U130
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U130 (
    .O(n835),
    .I0(in[172]),
    .I1(in[155])
  );
  //AND U130bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U130bar (
    .O(n835bar),
    .I0(inbar[172]),
    .I1(inbar[155])
  );
  //OR U131
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U131 (
    .O(n893),
    .I0(n834),
    .I1(n833)
  );
  //AND U131bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U131bar (
    .O(n893bar),
    .I0(n834bar),
    .I1(n833bar)
  );
  //OR U132
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U132 (
    .O(n833),
    .I0(n832),
    .I1(n831)
  );
  //AND U132bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U132bar (
    .O(n833bar),
    .I0(n832bar),
    .I1(n831bar)
  );
  //OR U133
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U133 (
    .O(n831),
    .I0(in[196]),
    .I1(in[173])
  );
  //AND U133bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U133bar (
    .O(n831bar),
    .I0(inbar[196]),
    .I1(inbar[173])
  );
  //OR U134
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U134 (
    .O(n832),
    .I0(in[222]),
    .I1(n830)
  );
  //AND U134bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U134bar (
    .O(n832bar),
    .I0(inbar[222]),
    .I1(n830bar)
  );
  //OR U135
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U135 (
    .O(n830),
    .I0(in[227]),
    .I1(in[226])
  );
  //AND U135bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U135bar (
    .O(n830bar),
    .I0(inbar[227]),
    .I1(inbar[226])
  );
  //OR U136
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U136 (
    .O(n834),
    .I0(n829),
    .I1(n828)
  );
  //AND U136bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U136bar (
    .O(n834bar),
    .I0(n829bar),
    .I1(n828bar)
  );
  //OR U137
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U137 (
    .O(n828),
    .I0(in[249]),
    .I1(in[231])
  );
  //AND U137bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U137bar (
    .O(n828bar),
    .I0(inbar[249]),
    .I1(inbar[231])
  );
  //OR U138
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U138 (
    .O(n829),
    .I0(in_28),
    .I1(n827)
  );
  //AND U138bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U138bar (
    .O(n829bar),
    .I0(in_28bar),
    .I1(n827bar)
  );
  //OR U139
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U139 (
    .O(n827),
    .I0(in_52),
    .I1(in_47)
  );
  //AND U139bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U139bar (
    .O(n827bar),
    .I0(in_52bar),
    .I1(in_47bar)
  );
  //OR U140
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U140 (
    .O(out[3]),
    .I0(n826),
    .I1(n825)
  );
  //AND U140bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U140bar (
    .O(outbar[3]),
    .I0(n826bar),
    .I1(n825bar)
  );
  //OR U141
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U141 (
    .O(n825),
    .I0(n824),
    .I1(n823)
  );
  //AND U141bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U141bar (
    .O(n825bar),
    .I0(n824bar),
    .I1(n823bar)
  );
  //OR U142
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U142 (
    .O(n823),
    .I0(n822),
    .I1(n821)
  );
  //AND U142bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U142bar (
    .O(n823bar),
    .I0(n822bar),
    .I1(n821bar)
  );
  //OR U143
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U143 (
    .O(n821),
    .I0(n820),
    .I1(n819)
  );
  //AND U143bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U143bar (
    .O(n821bar),
    .I0(n820bar),
    .I1(n819bar)
  );
  //OR U144
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U144 (
    .O(n822),
    .I0(n964),
    .I1(n818)
  );
  //AND U144bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U144bar (
    .O(n822bar),
    .I0(n964bar),
    .I1(n818bar)
  );
  //OR U145
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U145 (
    .O(n818),
    .I0(in[118]),
    .I1(n817)
  );
  //AND U145bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U145bar (
    .O(n818bar),
    .I0(inbar[118]),
    .I1(n817bar)
  );
  //OR U146
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U146 (
    .O(n964),
    .I0(n816),
    .I1(n815)
  );
  //AND U146bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U146bar (
    .O(n964bar),
    .I0(n816bar),
    .I1(n815bar)
  );
  //OR U147
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U147 (
    .O(n815),
    .I0(n814),
    .I1(n813)
  );
  //AND U147bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U147bar (
    .O(n815bar),
    .I0(n814bar),
    .I1(n813bar)
  );
  //OR U148
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U148 (
    .O(n813),
    .I0(n812),
    .I1(n811)
  );
  //AND U148bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U148bar (
    .O(n813bar),
    .I0(n812bar),
    .I1(n811bar)
  );
  //OR U149
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U149 (
    .O(n811),
    .I0(in[122]),
    .I1(in[111])
  );
  //AND U149bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U149bar (
    .O(n811bar),
    .I0(inbar[122]),
    .I1(inbar[111])
  );
  //OR U150
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U150 (
    .O(n812),
    .I0(in[154]),
    .I1(in[151])
  );
  //AND U150bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U150bar (
    .O(n812bar),
    .I0(inbar[154]),
    .I1(inbar[151])
  );
  //OR U151
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U151 (
    .O(n814),
    .I0(n810),
    .I1(n809)
  );
  //AND U151bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U151bar (
    .O(n814bar),
    .I0(n810bar),
    .I1(n809bar)
  );
  //OR U152
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U152 (
    .O(n809),
    .I0(in[187]),
    .I1(in[177])
  );
  //AND U152bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U152bar (
    .O(n809bar),
    .I0(inbar[187]),
    .I1(inbar[177])
  );
  //OR U153
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U153 (
    .O(n810),
    .I0(in[200]),
    .I1(in[192])
  );
  //AND U153bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U153bar (
    .O(n810bar),
    .I0(inbar[200]),
    .I1(inbar[192])
  );
  //OR U154
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U154 (
    .O(n816),
    .I0(n808),
    .I1(n807)
  );
  //AND U154bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U154bar (
    .O(n816bar),
    .I0(n808bar),
    .I1(n807bar)
  );
  //OR U155
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U155 (
    .O(n807),
    .I0(n806),
    .I1(n805)
  );
  //AND U155bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U155bar (
    .O(n807bar),
    .I0(n806bar),
    .I1(n805bar)
  );
  //OR U156
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U156 (
    .O(n805),
    .I0(in[225]),
    .I1(in[207])
  );
  //AND U156bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U156bar (
    .O(n805bar),
    .I0(inbar[225]),
    .I1(inbar[207])
  );
  //OR U157
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U157 (
    .O(n806),
    .I0(in[98]),
    .I1(in[226])
  );
  //AND U157bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U157bar (
    .O(n806bar),
    .I0(inbar[98]),
    .I1(inbar[226])
  );
  //OR U158
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U158 (
    .O(n808),
    .I0(n804),
    .I1(n803)
  );
  //AND U158bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U158bar (
    .O(n808bar),
    .I0(n804bar),
    .I1(n803bar)
  );
  //OR U159
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U159 (
    .O(n803),
    .I0(in_20),
    .I1(in_16)
  );
  //AND U159bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U159bar (
    .O(n803bar),
    .I0(in_20bar),
    .I1(in_16bar)
  );
  //OR U160
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U160 (
    .O(n804),
    .I0(in_55),
    .I1(in_45)
  );
  //AND U160bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U160bar (
    .O(n804bar),
    .I0(in_55bar),
    .I1(in_45bar)
  );
  //OR U161
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U161 (
    .O(n824),
    .I0(n802),
    .I1(n801)
  );
  //AND U161bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U161bar (
    .O(n824bar),
    .I0(n802bar),
    .I1(n801bar)
  );
  //OR U162
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U162 (
    .O(n801),
    .I0(in[162]),
    .I1(in[149])
  );
  //AND U162bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U162bar (
    .O(n801bar),
    .I0(inbar[162]),
    .I1(inbar[149])
  );
  //OR U163
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U163 (
    .O(n802),
    .I0(in[163]),
    .I1(n800)
  );
  //AND U163bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U163bar (
    .O(n802bar),
    .I0(inbar[163]),
    .I1(n800bar)
  );
  //OR U164
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U164 (
    .O(n800),
    .I0(in[191]),
    .I1(in[189])
  );
  //AND U164bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U164bar (
    .O(n800bar),
    .I0(inbar[191]),
    .I1(inbar[189])
  );
  //OR U165
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U165 (
    .O(n826),
    .I0(n799),
    .I1(n798)
  );
  //AND U165bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U165bar (
    .O(n826bar),
    .I0(n799bar),
    .I1(n798bar)
  );
  //OR U166
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U166 (
    .O(n798),
    .I0(n797),
    .I1(n796)
  );
  //AND U166bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U166bar (
    .O(n798bar),
    .I0(n797bar),
    .I1(n796bar)
  );
  //OR U167
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U167 (
    .O(n796),
    .I0(in[212]),
    .I1(in[193])
  );
  //AND U167bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U167bar (
    .O(n796bar),
    .I0(inbar[212]),
    .I1(inbar[193])
  );
  //OR U168
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U168 (
    .O(n797),
    .I0(in[238]),
    .I1(n795)
  );
  //AND U168bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U168bar (
    .O(n797bar),
    .I0(inbar[238]),
    .I1(n795bar)
  );
  //OR U169
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U169 (
    .O(n795),
    .I0(in[88]),
    .I1(in[247])
  );
  //AND U169bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U169bar (
    .O(n795bar),
    .I0(inbar[88]),
    .I1(inbar[247])
  );
  //OR U170
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U170 (
    .O(n799),
    .I0(n794),
    .I1(n793)
  );
  //AND U170bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U170bar (
    .O(n799bar),
    .I0(n794bar),
    .I1(n793bar)
  );
  //OR U171
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U171 (
    .O(n793),
    .I0(in[94]),
    .I1(in[92])
  );
  //AND U171bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U171bar (
    .O(n793bar),
    .I0(inbar[94]),
    .I1(inbar[92])
  );
  //OR U172
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U172 (
    .O(n794),
    .I0(in_52),
    .I1(n792)
  );
  //AND U172bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U172bar (
    .O(n794bar),
    .I0(in_52bar),
    .I1(n792bar)
  );
  //OR U173
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U173 (
    .O(n792),
    .I0(in_70),
    .I1(in_67)
  );
  //AND U173bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U173bar (
    .O(n792bar),
    .I0(in_70bar),
    .I1(in_67bar)
  );
  //OR U174
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U174 (
    .O(out[2]),
    .I0(n791),
    .I1(n790)
  );
  //AND U174bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U174bar (
    .O(outbar[2]),
    .I0(n791bar),
    .I1(n790bar)
  );
  //OR U175
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U175 (
    .O(n790),
    .I0(n789),
    .I1(n788)
  );
  //AND U175bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U175bar (
    .O(n790bar),
    .I0(n789bar),
    .I1(n788bar)
  );
  //OR U176
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U176 (
    .O(n788),
    .I0(n787),
    .I1(n786)
  );
  //AND U176bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U176bar (
    .O(n788bar),
    .I0(n787bar),
    .I1(n786bar)
  );
  //OR U177
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U177 (
    .O(n786),
    .I0(n819),
    .I1(n785)
  );
  //AND U177bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U177bar (
    .O(n786bar),
    .I0(n819bar),
    .I1(n785bar)
  );
  //OR U178
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U178 (
    .O(n819),
    .I0(n784),
    .I1(n783)
  );
  //AND U178bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U178bar (
    .O(n819bar),
    .I0(n784bar),
    .I1(n783bar)
  );
  //OR U179
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U179 (
    .O(n783),
    .I0(n782),
    .I1(n781)
  );
  //AND U179bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U179bar (
    .O(n783bar),
    .I0(n782bar),
    .I1(n781bar)
  );
  //OR U180
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U180 (
    .O(n781),
    .I0(n780),
    .I1(n779)
  );
  //AND U180bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U180bar (
    .O(n781bar),
    .I0(n780bar),
    .I1(n779bar)
  );
  //OR U181
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U181 (
    .O(n779),
    .I0(n962),
    .I1(n778)
  );
  //AND U181bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U181bar (
    .O(n779bar),
    .I0(n962bar),
    .I1(n778bar)
  );
  //OR U182
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U182 (
    .O(n962),
    .I0(n777),
    .I1(n776)
  );
  //AND U182bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U182bar (
    .O(n962bar),
    .I0(n777bar),
    .I1(n776bar)
  );
  //OR U183
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U183 (
    .O(n776),
    .I0(n775),
    .I1(n774)
  );
  //AND U183bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U183bar (
    .O(n776bar),
    .I0(n775bar),
    .I1(n774bar)
  );
  //OR U184
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U184 (
    .O(n774),
    .I0(n773),
    .I1(n772)
  );
  //AND U184bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U184bar (
    .O(n774bar),
    .I0(n773bar),
    .I1(n772bar)
  );
  //OR U185
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U185 (
    .O(n772),
    .I0(in[131]),
    .I1(in[120])
  );
  //AND U185bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U185bar (
    .O(n772bar),
    .I0(inbar[131]),
    .I1(inbar[120])
  );
  //OR U186
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U186 (
    .O(n773),
    .I0(in[153]),
    .I1(in[147])
  );
  //AND U186bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U186bar (
    .O(n773bar),
    .I0(inbar[153]),
    .I1(inbar[147])
  );
  //OR U187
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U187 (
    .O(n775),
    .I0(n771),
    .I1(n770)
  );
  //AND U187bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U187bar (
    .O(n775bar),
    .I0(n771bar),
    .I1(n770bar)
  );
  //OR U188
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U188 (
    .O(n770),
    .I0(in[170]),
    .I1(in[156])
  );
  //AND U188bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U188bar (
    .O(n770bar),
    .I0(inbar[170]),
    .I1(inbar[156])
  );
  //OR U189
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U189 (
    .O(n771),
    .I0(in[223]),
    .I1(in[190])
  );
  //AND U189bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U189bar (
    .O(n771bar),
    .I0(inbar[223]),
    .I1(inbar[190])
  );
  //OR U190
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U190 (
    .O(n777),
    .I0(n769),
    .I1(n768)
  );
  //AND U190bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U190bar (
    .O(n777bar),
    .I0(n769bar),
    .I1(n768bar)
  );
  //OR U191
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U191 (
    .O(n768),
    .I0(n767),
    .I1(n766)
  );
  //AND U191bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U191bar (
    .O(n768bar),
    .I0(n767bar),
    .I1(n766bar)
  );
  //OR U192
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U192 (
    .O(n766),
    .I0(in[236]),
    .I1(in[230])
  );
  //AND U192bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U192bar (
    .O(n766bar),
    .I0(inbar[236]),
    .I1(inbar[230])
  );
  //OR U193
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U193 (
    .O(n767),
    .I0(in[85]),
    .I1(in[240])
  );
  //AND U193bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U193bar (
    .O(n767bar),
    .I0(inbar[85]),
    .I1(inbar[240])
  );
  //OR U194
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U194 (
    .O(n769),
    .I0(n765),
    .I1(n764)
  );
  //AND U194bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U194bar (
    .O(n769bar),
    .I0(n765bar),
    .I1(n764bar)
  );
  //OR U195
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U195 (
    .O(n764),
    .I0(in_12),
    .I1(in[90])
  );
  //AND U195bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U195bar (
    .O(n764bar),
    .I0(in_12bar),
    .I1(inbar[90])
  );
  //OR U196
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U196 (
    .O(n765),
    .I0(in_39),
    .I1(in_28)
  );
  //AND U196bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U196bar (
    .O(n765bar),
    .I0(in_39bar),
    .I1(in_28bar)
  );
  //OR U197
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U197 (
    .O(n780),
    .I0(in[109]),
    .I1(n763)
  );
  //AND U197bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U197bar (
    .O(n780bar),
    .I0(inbar[109]),
    .I1(n763bar)
  );
  //OR U198
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U198 (
    .O(n782),
    .I0(n762),
    .I1(n761)
  );
  //AND U198bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U198bar (
    .O(n782bar),
    .I0(n762bar),
    .I1(n761bar)
  );
  //OR U199
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U199 (
    .O(n761),
    .I0(in[138]),
    .I1(in[129])
  );
  //AND U199bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U199bar (
    .O(n761bar),
    .I0(inbar[138]),
    .I1(inbar[129])
  );
  //OR U200
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U200 (
    .O(n762),
    .I0(in[157]),
    .I1(n760)
  );
  //AND U200bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U200bar (
    .O(n762bar),
    .I0(inbar[157]),
    .I1(n760bar)
  );
  //OR U201
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U201 (
    .O(n760),
    .I0(in[182]),
    .I1(in[167])
  );
  //AND U201bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U201bar (
    .O(n760bar),
    .I0(inbar[182]),
    .I1(inbar[167])
  );
  //OR U202
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U202 (
    .O(n784),
    .I0(n759),
    .I1(n758)
  );
  //AND U202bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U202bar (
    .O(n784bar),
    .I0(n759bar),
    .I1(n758bar)
  );
  //OR U203
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U203 (
    .O(n758),
    .I0(n757),
    .I1(n756)
  );
  //AND U203bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U203bar (
    .O(n758bar),
    .I0(n757bar),
    .I1(n756bar)
  );
  //OR U204
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U204 (
    .O(n756),
    .I0(in[195]),
    .I1(in[184])
  );
  //AND U204bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U204bar (
    .O(n756bar),
    .I0(inbar[195]),
    .I1(inbar[184])
  );
  //OR U205
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U205 (
    .O(n757),
    .I0(in[196]),
    .I1(n755)
  );
  //AND U205bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U205bar (
    .O(n757bar),
    .I0(inbar[196]),
    .I1(n755bar)
  );
  //OR U206
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U206 (
    .O(n755),
    .I0(in[215]),
    .I1(in[209])
  );
  //AND U206bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U206bar (
    .O(n755bar),
    .I0(inbar[215]),
    .I1(inbar[209])
  );
  //OR U207
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U207 (
    .O(n759),
    .I0(n754),
    .I1(n753)
  );
  //AND U207bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U207bar (
    .O(n759bar),
    .I0(n754bar),
    .I1(n753bar)
  );
  //OR U208
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U208 (
    .O(n753),
    .I0(in[93]),
    .I1(in[233])
  );
  //AND U208bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U208bar (
    .O(n753bar),
    .I0(inbar[93]),
    .I1(inbar[233])
  );
  //OR U209
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U209 (
    .O(n754),
    .I0(in_1),
    .I1(n752)
  );
  //AND U209bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U209bar (
    .O(n754bar),
    .I0(in_1bar),
    .I1(n752bar)
  );
  //OR U210
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U210 (
    .O(n752),
    .I0(in_69),
    .I1(in_66)
  );
  //AND U210bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U210bar (
    .O(n752bar),
    .I0(in_69bar),
    .I1(in_66bar)
  );
  //OR U211
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U211 (
    .O(n787),
    .I0(n966),
    .I1(n751)
  );
  //AND U211bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U211bar (
    .O(n787bar),
    .I0(n966bar),
    .I1(n751bar)
  );
  //OR U212
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U212 (
    .O(n751),
    .I0(in[134]),
    .I1(n750)
  );
  //AND U212bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U212bar (
    .O(n751bar),
    .I0(inbar[134]),
    .I1(n750bar)
  );
  //OR U213
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U213 (
    .O(n966),
    .I0(n749),
    .I1(n748)
  );
  //AND U213bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U213bar (
    .O(n966bar),
    .I0(n749bar),
    .I1(n748bar)
  );
  //OR U214
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U214 (
    .O(n748),
    .I0(n747),
    .I1(n746)
  );
  //AND U214bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U214bar (
    .O(n748bar),
    .I0(n747bar),
    .I1(n746bar)
  );
  //OR U215
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U215 (
    .O(n746),
    .I0(n745),
    .I1(n744)
  );
  //AND U215bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U215bar (
    .O(n746bar),
    .I0(n745bar),
    .I1(n744bar)
  );
  //OR U216
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U216 (
    .O(n744),
    .I0(in[136]),
    .I1(in[121])
  );
  //AND U216bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U216bar (
    .O(n744bar),
    .I0(inbar[136]),
    .I1(inbar[121])
  );
  //OR U217
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U217 (
    .O(n745),
    .I0(in[186]),
    .I1(in[174])
  );
  //AND U217bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U217bar (
    .O(n745bar),
    .I0(inbar[186]),
    .I1(inbar[174])
  );
  //OR U218
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U218 (
    .O(n747),
    .I0(n743),
    .I1(n742)
  );
  //AND U218bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U218bar (
    .O(n747bar),
    .I0(n743bar),
    .I1(n742bar)
  );
  //OR U219
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U219 (
    .O(n742),
    .I0(in[198]),
    .I1(in[197])
  );
  //AND U219bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U219bar (
    .O(n742bar),
    .I0(inbar[198]),
    .I1(inbar[197])
  );
  //OR U220
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U220 (
    .O(n743),
    .I0(in[214]),
    .I1(in[199])
  );
  //AND U220bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U220bar (
    .O(n743bar),
    .I0(inbar[214]),
    .I1(inbar[199])
  );
  //OR U221
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U221 (
    .O(n749),
    .I0(n741),
    .I1(n740)
  );
  //AND U221bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U221bar (
    .O(n749bar),
    .I0(n741bar),
    .I1(n740bar)
  );
  //OR U222
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U222 (
    .O(n740),
    .I0(n739),
    .I1(n738)
  );
  //AND U222bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U222bar (
    .O(n740bar),
    .I0(n739bar),
    .I1(n738bar)
  );
  //OR U223
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U223 (
    .O(n738),
    .I0(in[231]),
    .I1(in[220])
  );
  //AND U223bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U223bar (
    .O(n738bar),
    .I0(inbar[231]),
    .I1(inbar[220])
  );
  //OR U224
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U224 (
    .O(n739),
    .I0(in_25),
    .I1(in[245])
  );
  //AND U224bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U224bar (
    .O(n739bar),
    .I0(in_25bar),
    .I1(inbar[245])
  );
  //OR U225
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U225 (
    .O(n741),
    .I0(n737),
    .I1(n736)
  );
  //AND U225bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U225bar (
    .O(n741bar),
    .I0(n737bar),
    .I1(n736bar)
  );
  //OR U226
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U226 (
    .O(n736),
    .I0(in_53),
    .I1(in_29)
  );
  //AND U226bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U226bar (
    .O(n736bar),
    .I0(in_53bar),
    .I1(in_29bar)
  );
  //OR U227
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U227 (
    .O(n737),
    .I0(in_79),
    .I1(in_74)
  );
  //AND U227bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U227bar (
    .O(n737bar),
    .I0(in_79bar),
    .I1(in_74bar)
  );
  //OR U228
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U228 (
    .O(n789),
    .I0(n735),
    .I1(n734)
  );
  //AND U228bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U228bar (
    .O(n789bar),
    .I0(n735bar),
    .I1(n734bar)
  );
  //OR U229
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U229 (
    .O(n734),
    .I0(in[152]),
    .I1(in[140])
  );
  //AND U229bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U229bar (
    .O(n734bar),
    .I0(inbar[152]),
    .I1(inbar[140])
  );
  //OR U230
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U230 (
    .O(n735),
    .I0(in[155]),
    .I1(n733)
  );
  //AND U230bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U230bar (
    .O(n735bar),
    .I0(inbar[155]),
    .I1(n733bar)
  );
  //OR U231
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U231 (
    .O(n733),
    .I0(in[166]),
    .I1(in[165])
  );
  //AND U231bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U231bar (
    .O(n733bar),
    .I0(inbar[166]),
    .I1(inbar[165])
  );
  //OR U232
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U232 (
    .O(n791),
    .I0(n732),
    .I1(n731)
  );
  //AND U232bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U232bar (
    .O(n791bar),
    .I0(n732bar),
    .I1(n731bar)
  );
  //OR U233
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U233 (
    .O(n731),
    .I0(n730),
    .I1(n729)
  );
  //AND U233bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U233bar (
    .O(n731bar),
    .I0(n730bar),
    .I1(n729bar)
  );
  //OR U234
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U234 (
    .O(n729),
    .I0(in[202]),
    .I1(in[185])
  );
  //AND U234bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U234bar (
    .O(n729bar),
    .I0(inbar[202]),
    .I1(inbar[185])
  );
  //OR U235
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U235 (
    .O(n730),
    .I0(in[211]),
    .I1(n728)
  );
  //AND U235bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U235bar (
    .O(n730bar),
    .I0(inbar[211]),
    .I1(n728bar)
  );
  //OR U236
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U236 (
    .O(n728),
    .I0(in[255]),
    .I1(in[253])
  );
  //AND U236bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U236bar (
    .O(n728bar),
    .I0(inbar[255]),
    .I1(inbar[253])
  );
  //OR U237
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U237 (
    .O(n732),
    .I0(n727),
    .I1(n726)
  );
  //AND U237bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U237bar (
    .O(n732bar),
    .I0(n727bar),
    .I1(n726bar)
  );
  //OR U238
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U238 (
    .O(n726),
    .I0(in_35),
    .I1(in_15)
  );
  //AND U238bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U238bar (
    .O(n726bar),
    .I0(in_35bar),
    .I1(in_15bar)
  );
  //OR U239
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U239 (
    .O(n727),
    .I0(in_36),
    .I1(n725)
  );
  //AND U239bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U239bar (
    .O(n727bar),
    .I0(in_36bar),
    .I1(n725bar)
  );
  //OR U240
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U240 (
    .O(n725),
    .I0(in_48),
    .I1(in_40)
  );
  //AND U240bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U240bar (
    .O(n725bar),
    .I0(in_48bar),
    .I1(in_40bar)
  );
  //OR U241
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U241 (
    .O(out[1]),
    .I0(n724),
    .I1(n723)
  );
  //AND U241bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U241bar (
    .O(outbar[1]),
    .I0(n724bar),
    .I1(n723bar)
  );
  //OR U242
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U242 (
    .O(n723),
    .I0(n722),
    .I1(n721)
  );
  //AND U242bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U242bar (
    .O(n723bar),
    .I0(n722bar),
    .I1(n721bar)
  );
  //OR U243
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U243 (
    .O(n721),
    .I0(n720),
    .I1(n719)
  );
  //AND U243bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U243bar (
    .O(n721bar),
    .I0(n720bar),
    .I1(n719bar)
  );
  //OR U244
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U244 (
    .O(n719),
    .I0(n921),
    .I1(n887)
  );
  //AND U244bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U244bar (
    .O(n719bar),
    .I0(n921bar),
    .I1(n887bar)
  );
  //OR U245
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U245 (
    .O(n887),
    .I0(n718),
    .I1(n717)
  );
  //AND U245bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U245bar (
    .O(n887bar),
    .I0(n718bar),
    .I1(n717bar)
  );
  //OR U246
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U246 (
    .O(n717),
    .I0(n716),
    .I1(n715)
  );
  //AND U246bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U246bar (
    .O(n717bar),
    .I0(n716bar),
    .I1(n715bar)
  );
  //OR U247
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U247 (
    .O(n715),
    .I0(n714),
    .I1(n713)
  );
  //AND U247bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U247bar (
    .O(n715bar),
    .I0(n714bar),
    .I1(n713bar)
  );
  //OR U248
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U248 (
    .O(n713),
    .I0(in[116]),
    .I1(in[110])
  );
  //AND U248bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U248bar (
    .O(n713bar),
    .I0(inbar[116]),
    .I1(inbar[110])
  );
  //OR U249
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U249 (
    .O(n714),
    .I0(in[133]),
    .I1(in[130])
  );
  //AND U249bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U249bar (
    .O(n714bar),
    .I0(inbar[133]),
    .I1(inbar[130])
  );
  //OR U250
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U250 (
    .O(n716),
    .I0(n712),
    .I1(n711)
  );
  //AND U250bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U250bar (
    .O(n716bar),
    .I0(n712bar),
    .I1(n711bar)
  );
  //OR U251
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U251 (
    .O(n711),
    .I0(in[203]),
    .I1(in[135])
  );
  //AND U251bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U251bar (
    .O(n711bar),
    .I0(inbar[203]),
    .I1(inbar[135])
  );
  //OR U252
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U252 (
    .O(n712),
    .I0(in[232]),
    .I1(in[223])
  );
  //AND U252bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U252bar (
    .O(n712bar),
    .I0(inbar[232]),
    .I1(inbar[223])
  );
  //OR U253
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U253 (
    .O(n718),
    .I0(n710),
    .I1(n709)
  );
  //AND U253bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U253bar (
    .O(n718bar),
    .I0(n710bar),
    .I1(n709bar)
  );
  //OR U254
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U254 (
    .O(n709),
    .I0(n708),
    .I1(n707)
  );
  //AND U254bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U254bar (
    .O(n709bar),
    .I0(n708bar),
    .I1(n707bar)
  );
  //OR U255
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U255 (
    .O(n707),
    .I0(in[255]),
    .I1(in[233])
  );
  //AND U255bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U255bar (
    .O(n707bar),
    .I0(inbar[255]),
    .I1(inbar[233])
  );
  //OR U256
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U256 (
    .O(n708),
    .I0(in_53),
    .I1(in_34)
  );
  //AND U256bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U256bar (
    .O(n708bar),
    .I0(in_53bar),
    .I1(in_34bar)
  );
  //OR U257
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U257 (
    .O(n710),
    .I0(n706),
    .I1(n705)
  );
  //AND U257bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U257bar (
    .O(n710bar),
    .I0(n706bar),
    .I1(n705bar)
  );
  //OR U258
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U258 (
    .O(n705),
    .I0(in_57),
    .I1(in_55)
  );
  //AND U258bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U258bar (
    .O(n705bar),
    .I0(in_57bar),
    .I1(in_55bar)
  );
  //OR U259
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U259 (
    .O(n706),
    .I0(in_68),
    .I1(in_67)
  );
  //AND U259bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U259bar (
    .O(n706bar),
    .I0(in_68bar),
    .I1(in_67bar)
  );
  //OR U260
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U260 (
    .O(n921),
    .I0(n704),
    .I1(n703)
  );
  //AND U260bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U260bar (
    .O(n921bar),
    .I0(n704bar),
    .I1(n703bar)
  );
  //OR U261
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U261 (
    .O(n703),
    .I0(n702),
    .I1(n701)
  );
  //AND U261bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U261bar (
    .O(n703bar),
    .I0(n702bar),
    .I1(n701bar)
  );
  //OR U262
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U262 (
    .O(n701),
    .I0(n700),
    .I1(n699)
  );
  //AND U262bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U262bar (
    .O(n701bar),
    .I0(n700bar),
    .I1(n699bar)
  );
  //OR U263
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U263 (
    .O(n699),
    .I0(n944),
    .I1(n872)
  );
  //AND U263bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U263bar (
    .O(n699bar),
    .I0(n944bar),
    .I1(n872bar)
  );
  //OR U264
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U264 (
    .O(n872),
    .I0(n698),
    .I1(n697)
  );
  //AND U264bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U264bar (
    .O(n872bar),
    .I0(n698bar),
    .I1(n697bar)
  );
  //OR U265
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U265 (
    .O(n697),
    .I0(n696),
    .I1(n695)
  );
  //AND U265bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U265bar (
    .O(n697bar),
    .I0(n696bar),
    .I1(n695bar)
  );
  //OR U266
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U266 (
    .O(n695),
    .I0(n694),
    .I1(n693)
  );
  //AND U266bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U266bar (
    .O(n695bar),
    .I0(n694bar),
    .I1(n693bar)
  );
  //OR U267
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U267 (
    .O(n693),
    .I0(in[121]),
    .I1(in[102])
  );
  //AND U267bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U267bar (
    .O(n693bar),
    .I0(inbar[121]),
    .I1(inbar[102])
  );
  //OR U268
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U268 (
    .O(n694),
    .I0(in[162]),
    .I1(in[161])
  );
  //AND U268bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U268bar (
    .O(n694bar),
    .I0(inbar[162]),
    .I1(inbar[161])
  );
  //OR U269
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U269 (
    .O(n696),
    .I0(n692),
    .I1(n691)
  );
  //AND U269bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U269bar (
    .O(n696bar),
    .I0(n692bar),
    .I1(n691bar)
  );
  //OR U270
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U270 (
    .O(n691),
    .I0(in[192]),
    .I1(in[178])
  );
  //AND U270bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U270bar (
    .O(n691bar),
    .I0(inbar[192]),
    .I1(inbar[178])
  );
  //OR U271
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U271 (
    .O(n692),
    .I0(in[244]),
    .I1(in[209])
  );
  //AND U271bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U271bar (
    .O(n692bar),
    .I0(inbar[244]),
    .I1(inbar[209])
  );
  //OR U272
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U272 (
    .O(n698),
    .I0(n690),
    .I1(n689)
  );
  //AND U272bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U272bar (
    .O(n698bar),
    .I0(n690bar),
    .I1(n689bar)
  );
  //OR U273
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U273 (
    .O(n689),
    .I0(n688),
    .I1(n687)
  );
  //AND U273bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U273bar (
    .O(n689bar),
    .I0(n688bar),
    .I1(n687bar)
  );
  //OR U274
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U274 (
    .O(n687),
    .I0(in[90]),
    .I1(in[254])
  );
  //AND U274bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U274bar (
    .O(n687bar),
    .I0(inbar[90]),
    .I1(inbar[254])
  );
  //OR U275
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U275 (
    .O(n688),
    .I0(in_36),
    .I1(in_32)
  );
  //AND U275bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U275bar (
    .O(n688bar),
    .I0(in_36bar),
    .I1(in_32bar)
  );
  //OR U276
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U276 (
    .O(n690),
    .I0(n686),
    .I1(n685)
  );
  //AND U276bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U276bar (
    .O(n690bar),
    .I0(n686bar),
    .I1(n685bar)
  );
  //OR U277
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U277 (
    .O(n685),
    .I0(in_62),
    .I1(in_37)
  );
  //AND U277bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U277bar (
    .O(n685bar),
    .I0(in_62bar),
    .I1(in_37bar)
  );
  //OR U278
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U278 (
    .O(n686),
    .I0(in_75),
    .I1(in_73)
  );
  //AND U278bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U278bar (
    .O(n686bar),
    .I0(in_75bar),
    .I1(in_73bar)
  );
  //OR U279
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U279 (
    .O(n944),
    .I0(n684),
    .I1(n683)
  );
  //AND U279bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U279bar (
    .O(n944bar),
    .I0(n684bar),
    .I1(n683bar)
  );
  //OR U280
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U280 (
    .O(n683),
    .I0(n682),
    .I1(n681)
  );
  //AND U280bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U280bar (
    .O(n683bar),
    .I0(n682bar),
    .I1(n681bar)
  );
  //OR U281
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U281 (
    .O(n681),
    .I0(n680),
    .I1(n679)
  );
  //AND U281bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U281bar (
    .O(n681bar),
    .I0(n680bar),
    .I1(n679bar)
  );
  //OR U282
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U282 (
    .O(n679),
    .I0(in[171]),
    .I1(in[153])
  );
  //AND U282bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U282bar (
    .O(n679bar),
    .I0(inbar[171]),
    .I1(inbar[153])
  );
  //OR U283
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U283 (
    .O(n680),
    .I0(in[187]),
    .I1(in[176])
  );
  //AND U283bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U283bar (
    .O(n680bar),
    .I0(inbar[187]),
    .I1(inbar[176])
  );
  //OR U284
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U284 (
    .O(n682),
    .I0(n678),
    .I1(n677)
  );
  //AND U284bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U284bar (
    .O(n682bar),
    .I0(n678bar),
    .I1(n677bar)
  );
  //OR U285
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U285 (
    .O(n677),
    .I0(in[245]),
    .I1(in[211])
  );
  //AND U285bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U285bar (
    .O(n677bar),
    .I0(inbar[245]),
    .I1(inbar[211])
  );
  //OR U286
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U286 (
    .O(n678),
    .I0(in[97]),
    .I1(in[88])
  );
  //AND U286bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U286bar (
    .O(n678bar),
    .I0(inbar[97]),
    .I1(inbar[88])
  );
  //OR U287
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U287 (
    .O(n684),
    .I0(n676),
    .I1(n675)
  );
  //AND U287bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U287bar (
    .O(n684bar),
    .I0(n676bar),
    .I1(n675bar)
  );
  //OR U288
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U288 (
    .O(n675),
    .I0(n674),
    .I1(n673)
  );
  //AND U288bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U288bar (
    .O(n675bar),
    .I0(n674bar),
    .I1(n673bar)
  );
  //OR U289
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U289 (
    .O(n673),
    .I0(in_10),
    .I1(in_0)
  );
  //AND U289bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U289bar (
    .O(n673bar),
    .I0(in_10bar),
    .I1(in_0bar)
  );
  //OR U290
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U290 (
    .O(n674),
    .I0(in_59),
    .I1(in_5)
  );
  //AND U290bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U290bar (
    .O(n674bar),
    .I0(in_59bar),
    .I1(in_5bar)
  );
  //OR U291
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U291 (
    .O(n676),
    .I0(n672),
    .I1(n671)
  );
  //AND U291bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U291bar (
    .O(n676bar),
    .I0(n672bar),
    .I1(n671bar)
  );
  //OR U292
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U292 (
    .O(n671),
    .I0(in_60),
    .I1(in_6)
  );
  //AND U292bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U292bar (
    .O(n671bar),
    .I0(in_60bar),
    .I1(in_6bar)
  );
  //OR U293
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U293 (
    .O(n672),
    .I0(in_77),
    .I1(in_69)
  );
  //AND U293bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U293bar (
    .O(n672bar),
    .I0(in_77bar),
    .I1(in_69bar)
  );
  //OR U294
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U294 (
    .O(n700),
    .I0(in[113]),
    .I1(n864)
  );
  //AND U294bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U294bar (
    .O(n700bar),
    .I0(inbar[113]),
    .I1(n864bar)
  );
  //OR U295
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U295 (
    .O(n864),
    .I0(n670),
    .I1(n669)
  );
  //AND U295bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U295bar (
    .O(n864bar),
    .I0(n670bar),
    .I1(n669bar)
  );
  //OR U296
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U296 (
    .O(n669),
    .I0(n668),
    .I1(n667)
  );
  //AND U296bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U296bar (
    .O(n669bar),
    .I0(n668bar),
    .I1(n667bar)
  );
  //OR U297
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U297 (
    .O(n667),
    .I0(n666),
    .I1(n665)
  );
  //AND U297bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U297bar (
    .O(n667bar),
    .I0(n666bar),
    .I1(n665bar)
  );
  //OR U298
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U298 (
    .O(n665),
    .I0(in[125]),
    .I1(in[107])
  );
  //AND U298bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U298bar (
    .O(n665bar),
    .I0(inbar[125]),
    .I1(inbar[107])
  );
  //OR U299
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U299 (
    .O(n666),
    .I0(in[138]),
    .I1(in[126])
  );
  //AND U299bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U299bar (
    .O(n666bar),
    .I0(inbar[138]),
    .I1(inbar[126])
  );
  //OR U300
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U300 (
    .O(n668),
    .I0(n664),
    .I1(n663)
  );
  //AND U300bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U300bar (
    .O(n668bar),
    .I0(n664bar),
    .I1(n663bar)
  );
  //OR U301
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U301 (
    .O(n663),
    .I0(in[189]),
    .I1(in[143])
  );
  //AND U301bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U301bar (
    .O(n663bar),
    .I0(inbar[189]),
    .I1(inbar[143])
  );
  //OR U302
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U302 (
    .O(n664),
    .I0(in[99]),
    .I1(in[214])
  );
  //AND U302bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U302bar (
    .O(n664bar),
    .I0(inbar[99]),
    .I1(inbar[214])
  );
  //OR U303
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U303 (
    .O(n670),
    .I0(n662),
    .I1(n661)
  );
  //AND U303bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U303bar (
    .O(n670bar),
    .I0(n662bar),
    .I1(n661bar)
  );
  //OR U304
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U304 (
    .O(n661),
    .I0(n660),
    .I1(n659)
  );
  //AND U304bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U304bar (
    .O(n661bar),
    .I0(n660bar),
    .I1(n659bar)
  );
  //OR U305
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U305 (
    .O(n659),
    .I0(in_15),
    .I1(in_12)
  );
  //AND U305bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U305bar (
    .O(n659bar),
    .I0(in_15bar),
    .I1(in_12bar)
  );
  //OR U306
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U306 (
    .O(n660),
    .I0(in_20),
    .I1(in_2)
  );
  //AND U306bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U306bar (
    .O(n660bar),
    .I0(in_20bar),
    .I1(in_2bar)
  );
  //OR U307
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U307 (
    .O(n662),
    .I0(n658),
    .I1(n657)
  );
  //AND U307bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U307bar (
    .O(n662bar),
    .I0(n658bar),
    .I1(n657bar)
  );
  //OR U308
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U308 (
    .O(n657),
    .I0(in_30),
    .I1(in_3)
  );
  //AND U308bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U308bar (
    .O(n657bar),
    .I0(in_30bar),
    .I1(in_3bar)
  );
  //OR U309
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U309 (
    .O(n658),
    .I0(in_4),
    .I1(in_38)
  );
  //AND U309bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U309bar (
    .O(n658bar),
    .I0(in_4bar),
    .I1(in_38bar)
  );
  //OR U310
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U310 (
    .O(n702),
    .I0(n656),
    .I1(n655)
  );
  //AND U310bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U310bar (
    .O(n702bar),
    .I0(n656bar),
    .I1(n655bar)
  );
  //OR U311
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U311 (
    .O(n655),
    .I0(in[148]),
    .I1(in[137])
  );
  //AND U311bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U311bar (
    .O(n655bar),
    .I0(inbar[148]),
    .I1(inbar[137])
  );
  //OR U312
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U312 (
    .O(n656),
    .I0(in[149]),
    .I1(n654)
  );
  //AND U312bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U312bar (
    .O(n656bar),
    .I0(inbar[149]),
    .I1(n654bar)
  );
  //OR U313
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U313 (
    .O(n654),
    .I0(in[195]),
    .I1(in[190])
  );
  //AND U313bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U313bar (
    .O(n654bar),
    .I0(inbar[195]),
    .I1(inbar[190])
  );
  //OR U314
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U314 (
    .O(n704),
    .I0(n653),
    .I1(n652)
  );
  //AND U314bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U314bar (
    .O(n704bar),
    .I0(n653bar),
    .I1(n652bar)
  );
  //OR U315
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U315 (
    .O(n652),
    .I0(n651),
    .I1(n650)
  );
  //AND U315bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U315bar (
    .O(n652bar),
    .I0(n651bar),
    .I1(n650bar)
  );
  //OR U316
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U316 (
    .O(n650),
    .I0(in[98]),
    .I1(in[197])
  );
  //AND U316bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U316bar (
    .O(n650bar),
    .I0(inbar[98]),
    .I1(inbar[197])
  );
  //OR U317
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U317 (
    .O(n651),
    .I0(in_11),
    .I1(n649)
  );
  //AND U317bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U317bar (
    .O(n651bar),
    .I0(in_11bar),
    .I1(n649bar)
  );
  //OR U318
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U318 (
    .O(n649),
    .I0(in_26),
    .I1(in_14)
  );
  //AND U318bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U318bar (
    .O(n649bar),
    .I0(in_26bar),
    .I1(in_14bar)
  );
  //OR U319
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U319 (
    .O(n653),
    .I0(n648),
    .I1(n647)
  );
  //AND U319bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U319bar (
    .O(n653bar),
    .I0(n648bar),
    .I1(n647bar)
  );
  //OR U320
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U320 (
    .O(n647),
    .I0(in_35),
    .I1(in_27)
  );
  //AND U320bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U320bar (
    .O(n647bar),
    .I0(in_35bar),
    .I1(in_27bar)
  );
  //OR U321
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U321 (
    .O(n648),
    .I0(in_50),
    .I1(n646)
  );
  //AND U321bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U321bar (
    .O(n648bar),
    .I0(in_50bar),
    .I1(n646bar)
  );
  //OR U322
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U322 (
    .O(n646),
    .I0(in_78),
    .I1(in_61)
  );
  //AND U322bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U322bar (
    .O(n646bar),
    .I0(in_78bar),
    .I1(in_61bar)
  );
  //OR U323
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U323 (
    .O(n720),
    .I0(n942),
    .I1(n645)
  );
  //AND U323bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U323bar (
    .O(n720bar),
    .I0(n942bar),
    .I1(n645bar)
  );
  //OR U324
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U324 (
    .O(n645),
    .I0(in[106]),
    .I1(n863)
  );
  //AND U324bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U324bar (
    .O(n645bar),
    .I0(inbar[106]),
    .I1(n863bar)
  );
  //OR U325
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U325 (
    .O(n863),
    .I0(n644),
    .I1(n643)
  );
  //AND U325bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U325bar (
    .O(n863bar),
    .I0(n644bar),
    .I1(n643bar)
  );
  //OR U326
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U326 (
    .O(n643),
    .I0(n642),
    .I1(n641)
  );
  //AND U326bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U326bar (
    .O(n643bar),
    .I0(n642bar),
    .I1(n641bar)
  );
  //OR U327
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U327 (
    .O(n641),
    .I0(n640),
    .I1(n639)
  );
  //AND U327bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U327bar (
    .O(n641bar),
    .I0(n640bar),
    .I1(n639bar)
  );
  //OR U328
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U328 (
    .O(n639),
    .I0(in[127]),
    .I1(in[122])
  );
  //AND U328bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U328bar (
    .O(n639bar),
    .I0(inbar[127]),
    .I1(inbar[122])
  );
  //OR U329
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U329 (
    .O(n640),
    .I0(in[156]),
    .I1(in[132])
  );
  //AND U329bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U329bar (
    .O(n640bar),
    .I0(inbar[156]),
    .I1(inbar[132])
  );
  //OR U330
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U330 (
    .O(n642),
    .I0(n638),
    .I1(n637)
  );
  //AND U330bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U330bar (
    .O(n642bar),
    .I0(n638bar),
    .I1(n637bar)
  );
  //OR U331
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U331 (
    .O(n637),
    .I0(in[159]),
    .I1(in[157])
  );
  //AND U331bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U331bar (
    .O(n637bar),
    .I0(inbar[159]),
    .I1(inbar[157])
  );
  //OR U332
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U332 (
    .O(n638),
    .I0(in[185]),
    .I1(in[169])
  );
  //AND U332bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U332bar (
    .O(n638bar),
    .I0(inbar[185]),
    .I1(inbar[169])
  );
  //OR U333
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U333 (
    .O(n644),
    .I0(n636),
    .I1(n635)
  );
  //AND U333bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U333bar (
    .O(n644bar),
    .I0(n636bar),
    .I1(n635bar)
  );
  //OR U334
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U334 (
    .O(n635),
    .I0(n634),
    .I1(n633)
  );
  //AND U334bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U334bar (
    .O(n635bar),
    .I0(n634bar),
    .I1(n633bar)
  );
  //OR U335
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U335 (
    .O(n633),
    .I0(in[239]),
    .I1(in[218])
  );
  //AND U335bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U335bar (
    .O(n633bar),
    .I0(inbar[239]),
    .I1(inbar[218])
  );
  //OR U336
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U336 (
    .O(n634),
    .I0(in_13),
    .I1(in[87])
  );
  //AND U336bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U336bar (
    .O(n634bar),
    .I0(in_13bar),
    .I1(inbar[87])
  );
  //OR U337
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U337 (
    .O(n636),
    .I0(n632),
    .I1(n631)
  );
  //AND U337bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U337bar (
    .O(n636bar),
    .I0(n632bar),
    .I1(n631bar)
  );
  //OR U338
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U338 (
    .O(n631),
    .I0(in_72),
    .I1(in_70)
  );
  //AND U338bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U338bar (
    .O(n631bar),
    .I0(in_72bar),
    .I1(in_70bar)
  );
  //OR U339
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U339 (
    .O(n632),
    .I0(in_80),
    .I1(in_74)
  );
  //AND U339bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U339bar (
    .O(n632bar),
    .I0(in_80bar),
    .I1(in_74bar)
  );
  //OR U340
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U340 (
    .O(n942),
    .I0(n630),
    .I1(n629)
  );
  //AND U340bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U340bar (
    .O(n942bar),
    .I0(n630bar),
    .I1(n629bar)
  );
  //OR U341
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U341 (
    .O(n629),
    .I0(n628),
    .I1(n627)
  );
  //AND U341bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U341bar (
    .O(n629bar),
    .I0(n628bar),
    .I1(n627bar)
  );
  //OR U342
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U342 (
    .O(n627),
    .I0(n626),
    .I1(n625)
  );
  //AND U342bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U342bar (
    .O(n627bar),
    .I0(n626bar),
    .I1(n625bar)
  );
  //OR U343
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U343 (
    .O(n625),
    .I0(in[146]),
    .I1(in[100])
  );
  //AND U343bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U343bar (
    .O(n625bar),
    .I0(inbar[146]),
    .I1(inbar[100])
  );
  //OR U344
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U344 (
    .O(n626),
    .I0(in[168]),
    .I1(in[152])
  );
  //AND U344bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U344bar (
    .O(n626bar),
    .I0(inbar[168]),
    .I1(inbar[152])
  );
  //OR U345
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U345 (
    .O(n628),
    .I0(n624),
    .I1(n623)
  );
  //AND U345bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U345bar (
    .O(n628bar),
    .I0(n624bar),
    .I1(n623bar)
  );
  //OR U346
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U346 (
    .O(n623),
    .I0(in[199]),
    .I1(in[182])
  );
  //AND U346bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U346bar (
    .O(n623bar),
    .I0(inbar[199]),
    .I1(inbar[182])
  );
  //OR U347
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U347 (
    .O(n624),
    .I0(in[236]),
    .I1(in[204])
  );
  //AND U347bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U347bar (
    .O(n624bar),
    .I0(inbar[236]),
    .I1(inbar[204])
  );
  //OR U348
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U348 (
    .O(n630),
    .I0(n622),
    .I1(n621)
  );
  //AND U348bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U348bar (
    .O(n630bar),
    .I0(n622bar),
    .I1(n621bar)
  );
  //OR U349
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U349 (
    .O(n621),
    .I0(n620),
    .I1(n619)
  );
  //AND U349bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U349bar (
    .O(n621bar),
    .I0(n620bar),
    .I1(n619bar)
  );
  //OR U350
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U350 (
    .O(n619),
    .I0(in[89]),
    .I1(in[246])
  );
  //AND U350bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U350bar (
    .O(n619bar),
    .I0(inbar[89]),
    .I1(inbar[246])
  );
  //OR U351
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U351 (
    .O(n620),
    .I0(in[95]),
    .I1(in[92])
  );
  //AND U351bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U351bar (
    .O(n620bar),
    .I0(inbar[95]),
    .I1(inbar[92])
  );
  //OR U352
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U352 (
    .O(n622),
    .I0(n618),
    .I1(n617)
  );
  //AND U352bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U352bar (
    .O(n622bar),
    .I0(n618bar),
    .I1(n617bar)
  );
  //OR U353
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U353 (
    .O(n617),
    .I0(in_22),
    .I1(in_16)
  );
  //AND U353bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U353bar (
    .O(n617bar),
    .I0(in_22bar),
    .I1(in_16bar)
  );
  //OR U354
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U354 (
    .O(n618),
    .I0(in_51),
    .I1(in_49)
  );
  //AND U354bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U354bar (
    .O(n618bar),
    .I0(in_51bar),
    .I1(in_49bar)
  );
  //OR U355
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U355 (
    .O(n722),
    .I0(n616),
    .I1(n615)
  );
  //AND U355bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U355bar (
    .O(n722bar),
    .I0(n616bar),
    .I1(n615bar)
  );
  //OR U356
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U356 (
    .O(n615),
    .I0(in[158]),
    .I1(in[115])
  );
  //AND U356bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U356bar (
    .O(n615bar),
    .I0(inbar[158]),
    .I1(inbar[115])
  );
  //OR U357
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U357 (
    .O(n616),
    .I0(in[163]),
    .I1(n614)
  );
  //AND U357bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U357bar (
    .O(n616bar),
    .I0(inbar[163]),
    .I1(n614bar)
  );
  //OR U358
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U358 (
    .O(n614),
    .I0(in[206]),
    .I1(in[165])
  );
  //AND U358bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U358bar (
    .O(n614bar),
    .I0(inbar[206]),
    .I1(inbar[165])
  );
  //OR U359
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U359 (
    .O(n724),
    .I0(n613),
    .I1(n612)
  );
  //AND U359bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U359bar (
    .O(n724bar),
    .I0(n613bar),
    .I1(n612bar)
  );
  //OR U360
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U360 (
    .O(n612),
    .I0(n611),
    .I1(n610)
  );
  //AND U360bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U360bar (
    .O(n612bar),
    .I0(n611bar),
    .I1(n610bar)
  );
  //OR U361
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U361 (
    .O(n610),
    .I0(in[213]),
    .I1(in[207])
  );
  //AND U361bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U361bar (
    .O(n610bar),
    .I0(inbar[213]),
    .I1(inbar[207])
  );
  //OR U362
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U362 (
    .O(n611),
    .I0(in[215]),
    .I1(n609)
  );
  //AND U362bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U362bar (
    .O(n611bar),
    .I0(inbar[215]),
    .I1(n609bar)
  );
  //OR U363
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U363 (
    .O(n609),
    .I0(in[230]),
    .I1(in[220])
  );
  //AND U363bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U363bar (
    .O(n609bar),
    .I0(inbar[230]),
    .I1(inbar[220])
  );
  //OR U364
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U364 (
    .O(n613),
    .I0(n608),
    .I1(n607)
  );
  //AND U364bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U364bar (
    .O(n613bar),
    .I0(n608bar),
    .I1(n607bar)
  );
  //OR U365
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U365 (
    .O(n607),
    .I0(in[251]),
    .I1(in[234])
  );
  //AND U365bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U365bar (
    .O(n607bar),
    .I0(inbar[251]),
    .I1(inbar[234])
  );
  //OR U366
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U366 (
    .O(n608),
    .I0(in_17),
    .I1(n606)
  );
  //AND U366bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U366bar (
    .O(n608bar),
    .I0(in_17bar),
    .I1(n606bar)
  );
  //OR U367
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U367 (
    .O(n606),
    .I0(in_65),
    .I1(in_56)
  );
  //AND U367bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U367bar (
    .O(n606bar),
    .I0(in_65bar),
    .I1(in_56bar)
  );
  //OR U368
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U368 (
    .O(out[0]),
    .I0(n605),
    .I1(n604)
  );
  //AND U368bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U368bar (
    .O(outbar[0]),
    .I0(n605bar),
    .I1(n604bar)
  );
  //OR U369
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U369 (
    .O(n604),
    .I0(n603),
    .I1(n602)
  );
  //AND U369bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U369bar (
    .O(n604bar),
    .I0(n603bar),
    .I1(n602bar)
  );
  //OR U370
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U370 (
    .O(n602),
    .I0(n601),
    .I1(n600)
  );
  //AND U370bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U370bar (
    .O(n602bar),
    .I0(n601bar),
    .I1(n600bar)
  );
  //OR U371
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U371 (
    .O(n600),
    .I0(n820),
    .I1(n785)
  );
  //AND U371bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U371bar (
    .O(n600bar),
    .I0(n820bar),
    .I1(n785bar)
  );
  //OR U372
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U372 (
    .O(n785),
    .I0(n599),
    .I1(n598)
  );
  //AND U372bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U372bar (
    .O(n785bar),
    .I0(n599bar),
    .I1(n598bar)
  );
  //OR U373
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U373 (
    .O(n598),
    .I0(n597),
    .I1(n596)
  );
  //AND U373bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U373bar (
    .O(n598bar),
    .I0(n597bar),
    .I1(n596bar)
  );
  //OR U374
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U374 (
    .O(n596),
    .I0(n595),
    .I1(n594)
  );
  //AND U374bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U374bar (
    .O(n596bar),
    .I0(n595bar),
    .I1(n594bar)
  );
  //OR U375
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U375 (
    .O(n594),
    .I0(in[135]),
    .I1(in[104])
  );
  //AND U375bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U375bar (
    .O(n594bar),
    .I0(inbar[135]),
    .I1(inbar[104])
  );
  //OR U376
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U376 (
    .O(n595),
    .I0(in[188]),
    .I1(in[178])
  );
  //AND U376bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U376bar (
    .O(n595bar),
    .I0(inbar[188]),
    .I1(inbar[178])
  );
  //OR U377
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U377 (
    .O(n597),
    .I0(n593),
    .I1(n592)
  );
  //AND U377bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U377bar (
    .O(n597bar),
    .I0(n593bar),
    .I1(n592bar)
  );
  //OR U378
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U378 (
    .O(n592),
    .I0(in[217]),
    .I1(in[194])
  );
  //AND U378bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U378bar (
    .O(n592bar),
    .I0(inbar[217]),
    .I1(inbar[194])
  );
  //OR U379
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U379 (
    .O(n593),
    .I0(in[237]),
    .I1(in[218])
  );
  //AND U379bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U379bar (
    .O(n593bar),
    .I0(inbar[237]),
    .I1(inbar[218])
  );
  //OR U380
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U380 (
    .O(n599),
    .I0(n591),
    .I1(n590)
  );
  //AND U380bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U380bar (
    .O(n599bar),
    .I0(n591bar),
    .I1(n590bar)
  );
  //OR U381
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U381 (
    .O(n590),
    .I0(n589),
    .I1(n588)
  );
  //AND U381bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U381bar (
    .O(n590bar),
    .I0(n589bar),
    .I1(n588bar)
  );
  //OR U382
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U382 (
    .O(n588),
    .I0(in_2),
    .I1(in_10)
  );
  //AND U382bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U382bar (
    .O(n588bar),
    .I0(in_2bar),
    .I1(in_10bar)
  );
  //OR U383
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U383 (
    .O(n589),
    .I0(in_47),
    .I1(in_22)
  );
  //AND U383bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U383bar (
    .O(n589bar),
    .I0(in_47bar),
    .I1(in_22bar)
  );
  //OR U384
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U384 (
    .O(n591),
    .I0(n587),
    .I1(n586)
  );
  //AND U384bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U384bar (
    .O(n591bar),
    .I0(n587bar),
    .I1(n586bar)
  );
  //OR U385
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U385 (
    .O(n586),
    .I0(in_56),
    .I1(in_54)
  );
  //AND U385bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U385bar (
    .O(n586bar),
    .I0(in_56bar),
    .I1(in_54bar)
  );
  //OR U386
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U386 (
    .O(n587),
    .I0(in_63),
    .I1(in_61)
  );
  //AND U386bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U386bar (
    .O(n587bar),
    .I0(in_63bar),
    .I1(in_61bar)
  );
  //OR U387
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U387 (
    .O(n820),
    .I0(n585),
    .I1(n584)
  );
  //AND U387bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U387bar (
    .O(n820bar),
    .I0(n585bar),
    .I1(n584bar)
  );
  //OR U388
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U388 (
    .O(n584),
    .I0(n583),
    .I1(n582)
  );
  //AND U388bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U388bar (
    .O(n584bar),
    .I0(n583bar),
    .I1(n582bar)
  );
  //OR U389
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U389 (
    .O(n582),
    .I0(n581),
    .I1(n580)
  );
  //AND U389bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U389bar (
    .O(n582bar),
    .I0(n581bar),
    .I1(n580bar)
  );
  //OR U390
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U390 (
    .O(n580),
    .I0(in[158]),
    .I1(in[142])
  );
  //AND U390bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U390bar (
    .O(n580bar),
    .I0(inbar[158]),
    .I1(inbar[142])
  );
  //OR U391
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U391 (
    .O(n581),
    .I0(in[175]),
    .I1(in[164])
  );
  //AND U391bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U391bar (
    .O(n581bar),
    .I0(inbar[175]),
    .I1(inbar[164])
  );
  //OR U392
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U392 (
    .O(n583),
    .I0(n579),
    .I1(n578)
  );
  //AND U392bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U392bar (
    .O(n583bar),
    .I0(n579bar),
    .I1(n578bar)
  );
  //OR U393
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U393 (
    .O(n578),
    .I0(in[228]),
    .I1(in[204])
  );
  //AND U393bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U393bar (
    .O(n578bar),
    .I0(inbar[228]),
    .I1(inbar[204])
  );
  //OR U394
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U394 (
    .O(n579),
    .I0(in[91]),
    .I1(in[87])
  );
  //AND U394bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U394bar (
    .O(n579bar),
    .I0(inbar[91]),
    .I1(inbar[87])
  );
  //OR U395
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U395 (
    .O(n585),
    .I0(n577),
    .I1(n576)
  );
  //AND U395bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U395bar (
    .O(n585bar),
    .I0(n577bar),
    .I1(n576bar)
  );
  //OR U396
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U396 (
    .O(n576),
    .I0(n575),
    .I1(n574)
  );
  //AND U396bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U396bar (
    .O(n576bar),
    .I0(n575bar),
    .I1(n574bar)
  );
  //OR U397
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U397 (
    .O(n574),
    .I0(in_21),
    .I1(in_11)
  );
  //AND U397bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U397bar (
    .O(n574bar),
    .I0(in_21bar),
    .I1(in_11bar)
  );
  //OR U398
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U398 (
    .O(n575),
    .I0(in_5),
    .I1(in_3)
  );
  //AND U398bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U398bar (
    .O(n575bar),
    .I0(in_5bar),
    .I1(in_3bar)
  );
  //OR U399
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U399 (
    .O(n577),
    .I0(n573),
    .I1(n572)
  );
  //AND U399bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U399bar (
    .O(n577bar),
    .I0(n573bar),
    .I1(n572bar)
  );
  //OR U400
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U400 (
    .O(n572),
    .I0(in_68),
    .I1(in_64)
  );
  //AND U400bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U400bar (
    .O(n572bar),
    .I0(in_68bar),
    .I1(in_64bar)
  );
  //OR U401
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U401 (
    .O(n573),
    .I0(in_76),
    .I1(in_73)
  );
  //AND U401bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U401bar (
    .O(n573bar),
    .I0(in_76bar),
    .I1(in_73bar)
  );
  //OR U402
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U402 (
    .O(n601),
    .I0(n778),
    .I1(n571)
  );
  //AND U402bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U402bar (
    .O(n601bar),
    .I0(n778bar),
    .I1(n571bar)
  );
  //OR U403
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U403 (
    .O(n571),
    .I0(in[100]),
    .I1(n965)
  );
  //AND U403bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U403bar (
    .O(n571bar),
    .I0(inbar[100]),
    .I1(n965bar)
  );
  //OR U404
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U404 (
    .O(n965),
    .I0(n570),
    .I1(n569)
  );
  //AND U404bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U404bar (
    .O(n965bar),
    .I0(n570bar),
    .I1(n569bar)
  );
  //OR U405
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U405 (
    .O(n569),
    .I0(n568),
    .I1(n567)
  );
  //AND U405bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U405bar (
    .O(n569bar),
    .I0(n568bar),
    .I1(n567bar)
  );
  //OR U406
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U406 (
    .O(n567),
    .I0(n566),
    .I1(n565)
  );
  //AND U406bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U406bar (
    .O(n567bar),
    .I0(n566bar),
    .I1(n565bar)
  );
  //OR U407
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U407 (
    .O(n565),
    .I0(n817),
    .I1(n750)
  );
  //AND U407bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U407bar (
    .O(n565bar),
    .I0(n817bar),
    .I1(n750bar)
  );
  //OR U408
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U408 (
    .O(n750),
    .I0(n564),
    .I1(n563)
  );
  //AND U408bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U408bar (
    .O(n750bar),
    .I0(n564bar),
    .I1(n563bar)
  );
  //OR U409
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U409 (
    .O(n563),
    .I0(n562),
    .I1(n561)
  );
  //AND U409bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U409bar (
    .O(n563bar),
    .I0(n562bar),
    .I1(n561bar)
  );
  //OR U410
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U410 (
    .O(n561),
    .I0(n560),
    .I1(n559)
  );
  //AND U410bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U410bar (
    .O(n561bar),
    .I0(n560bar),
    .I1(n559bar)
  );
  //OR U411
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U411 (
    .O(n559),
    .I0(in[119]),
    .I1(in[103])
  );
  //AND U411bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U411bar (
    .O(n559bar),
    .I0(inbar[119]),
    .I1(inbar[103])
  );
  //OR U412
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U412 (
    .O(n560),
    .I0(in[137]),
    .I1(in[133])
  );
  //AND U412bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U412bar (
    .O(n560bar),
    .I0(inbar[137]),
    .I1(inbar[133])
  );
  //OR U413
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U413 (
    .O(n562),
    .I0(n558),
    .I1(n557)
  );
  //AND U413bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U413bar (
    .O(n562bar),
    .I0(n558bar),
    .I1(n557bar)
  );
  //OR U414
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U414 (
    .O(n557),
    .I0(in[176]),
    .I1(in[173])
  );
  //AND U414bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U414bar (
    .O(n557bar),
    .I0(inbar[176]),
    .I1(inbar[173])
  );
  //OR U415
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U415 (
    .O(n558),
    .I0(in[210]),
    .I1(in[181])
  );
  //AND U415bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U415bar (
    .O(n558bar),
    .I0(inbar[210]),
    .I1(inbar[181])
  );
  //OR U416
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U416 (
    .O(n564),
    .I0(n556),
    .I1(n555)
  );
  //AND U416bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U416bar (
    .O(n564bar),
    .I0(n556bar),
    .I1(n555bar)
  );
  //OR U417
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U417 (
    .O(n555),
    .I0(n554),
    .I1(n553)
  );
  //AND U417bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U417bar (
    .O(n555bar),
    .I0(n554bar),
    .I1(n553bar)
  );
  //OR U418
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U418 (
    .O(n553),
    .I0(in_13),
    .I1(in[234])
  );
  //AND U418bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U418bar (
    .O(n553bar),
    .I0(in_13bar),
    .I1(inbar[234])
  );
  //OR U419
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U419 (
    .O(n554),
    .I0(in_38),
    .I1(in_32)
  );
  //AND U419bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U419bar (
    .O(n554bar),
    .I0(in_38bar),
    .I1(in_32bar)
  );
  //OR U420
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U420 (
    .O(n556),
    .I0(n552),
    .I1(n551)
  );
  //AND U420bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U420bar (
    .O(n556bar),
    .I0(n552bar),
    .I1(n551bar)
  );
  //OR U421
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U421 (
    .O(n551),
    .I0(in_42),
    .I1(in_41)
  );
  //AND U421bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U421bar (
    .O(n551bar),
    .I0(in_42bar),
    .I1(in_41bar)
  );
  //OR U422
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U422 (
    .O(n552),
    .I0(in_7),
    .I1(in_49)
  );
  //AND U422bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U422bar (
    .O(n552bar),
    .I0(in_7bar),
    .I1(in_49bar)
  );
  //OR U423
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U423 (
    .O(n817),
    .I0(n550),
    .I1(n549)
  );
  //AND U423bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U423bar (
    .O(n817bar),
    .I0(n550bar),
    .I1(n549bar)
  );
  //OR U424
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U424 (
    .O(n549),
    .I0(n548),
    .I1(n547)
  );
  //AND U424bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U424bar (
    .O(n549bar),
    .I0(n548bar),
    .I1(n547bar)
  );
  //OR U425
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U425 (
    .O(n547),
    .I0(n546),
    .I1(n545)
  );
  //AND U425bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U425bar (
    .O(n547bar),
    .I0(n546bar),
    .I1(n545bar)
  );
  //OR U426
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U426 (
    .O(n545),
    .I0(in[159]),
    .I1(in[105])
  );
  //AND U426bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U426bar (
    .O(n545bar),
    .I0(inbar[159]),
    .I1(inbar[105])
  );
  //OR U427
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U427 (
    .O(n546),
    .I0(in[206]),
    .I1(in[183])
  );
  //AND U427bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U427bar (
    .O(n546bar),
    .I0(inbar[206]),
    .I1(inbar[183])
  );
  //OR U428
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U428 (
    .O(n548),
    .I0(n544),
    .I1(n543)
  );
  //AND U428bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U428bar (
    .O(n548bar),
    .I0(n544bar),
    .I1(n543bar)
  );
  //OR U429
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U429 (
    .O(n543),
    .I0(in[229]),
    .I1(in[219])
  );
  //AND U429bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U429bar (
    .O(n543bar),
    .I0(inbar[229]),
    .I1(inbar[219])
  );
  //OR U430
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U430 (
    .O(n544),
    .I0(in[235]),
    .I1(in[232])
  );
  //AND U430bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U430bar (
    .O(n544bar),
    .I0(inbar[235]),
    .I1(inbar[232])
  );
  //OR U431
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U431 (
    .O(n550),
    .I0(n542),
    .I1(n541)
  );
  //AND U431bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U431bar (
    .O(n550bar),
    .I0(n542bar),
    .I1(n541bar)
  );
  //OR U432
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U432 (
    .O(n541),
    .I0(n540),
    .I1(n539)
  );
  //AND U432bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U432bar (
    .O(n541bar),
    .I0(n540bar),
    .I1(n539bar)
  );
  //OR U433
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U433 (
    .O(n539),
    .I0(in[249]),
    .I1(in[242])
  );
  //AND U433bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U433bar (
    .O(n539bar),
    .I0(inbar[249]),
    .I1(inbar[242])
  );
  //OR U434
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U434 (
    .O(n540),
    .I0(in[89]),
    .I1(in[254])
  );
  //AND U434bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U434bar (
    .O(n540bar),
    .I0(inbar[89]),
    .I1(inbar[254])
  );
  //OR U435
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U435 (
    .O(n542),
    .I0(n538),
    .I1(n537)
  );
  //AND U435bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U435bar (
    .O(n542bar),
    .I0(n538bar),
    .I1(n537bar)
  );
  //OR U436
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U436 (
    .O(n537),
    .I0(in_14),
    .I1(in[99])
  );
  //AND U436bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U436bar (
    .O(n537bar),
    .I0(in_14bar),
    .I1(inbar[99])
  );
  //OR U437
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U437 (
    .O(n538),
    .I0(in_60),
    .I1(in_18)
  );
  //AND U437bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U437bar (
    .O(n538bar),
    .I0(in_60bar),
    .I1(in_18bar)
  );
  //OR U438
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U438 (
    .O(n566),
    .I0(in[113]),
    .I1(n763)
  );
  //AND U438bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U438bar (
    .O(n566bar),
    .I0(inbar[113]),
    .I1(n763bar)
  );
  //OR U439
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U439 (
    .O(n763),
    .I0(n536),
    .I1(n535)
  );
  //AND U439bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U439bar (
    .O(n763bar),
    .I0(n536bar),
    .I1(n535bar)
  );
  //OR U440
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U440 (
    .O(n535),
    .I0(n534),
    .I1(n533)
  );
  //AND U440bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U440bar (
    .O(n535bar),
    .I0(n534bar),
    .I1(n533bar)
  );
  //OR U441
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U441 (
    .O(n533),
    .I0(n532),
    .I1(n531)
  );
  //AND U441bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U441bar (
    .O(n533bar),
    .I0(n532bar),
    .I1(n531bar)
  );
  //OR U442
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U442 (
    .O(n531),
    .I0(in[115]),
    .I1(in[110])
  );
  //AND U442bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U442bar (
    .O(n531bar),
    .I0(inbar[115]),
    .I1(inbar[110])
  );
  //OR U443
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U443 (
    .O(n532),
    .I0(in[125]),
    .I1(in[117])
  );
  //AND U443bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U443bar (
    .O(n532bar),
    .I0(inbar[125]),
    .I1(inbar[117])
  );
  //OR U444
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U444 (
    .O(n534),
    .I0(n530),
    .I1(n529)
  );
  //AND U444bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U444bar (
    .O(n534bar),
    .I0(n530bar),
    .I1(n529bar)
  );
  //OR U445
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U445 (
    .O(n529),
    .I0(in[180]),
    .I1(in[128])
  );
  //AND U445bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U445bar (
    .O(n529bar),
    .I0(inbar[180]),
    .I1(inbar[128])
  );
  //OR U446
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U446 (
    .O(n530),
    .I0(in[205]),
    .I1(in[201])
  );
  //AND U446bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U446bar (
    .O(n530bar),
    .I0(inbar[205]),
    .I1(inbar[201])
  );
  //OR U447
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U447 (
    .O(n536),
    .I0(n528),
    .I1(n527)
  );
  //AND U447bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U447bar (
    .O(n536bar),
    .I0(n528bar),
    .I1(n527bar)
  );
  //OR U448
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U448 (
    .O(n527),
    .I0(n526),
    .I1(n525)
  );
  //AND U448bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U448bar (
    .O(n527bar),
    .I0(n526bar),
    .I1(n525bar)
  );
  //OR U449
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U449 (
    .O(n525),
    .I0(in[244]),
    .I1(in[239])
  );
  //AND U449bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U449bar (
    .O(n525bar),
    .I0(inbar[244]),
    .I1(inbar[239])
  );
  //OR U450
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U450 (
    .O(n526),
    .I0(in[95]),
    .I1(in[83])
  );
  //AND U450bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U450bar (
    .O(n526bar),
    .I0(inbar[95]),
    .I1(inbar[83])
  );
  //OR U451
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U451 (
    .O(n528),
    .I0(n524),
    .I1(n523)
  );
  //AND U451bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U451bar (
    .O(n528bar),
    .I0(n524bar),
    .I1(n523bar)
  );
  //OR U452
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U452 (
    .O(n523),
    .I0(in_24),
    .I1(in[97])
  );
  //AND U452bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U452bar (
    .O(n523bar),
    .I0(in_24bar),
    .I1(inbar[97])
  );
  //OR U453
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U453 (
    .O(n524),
    .I0(in_33),
    .I1(in_27)
  );
  //AND U453bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U453bar (
    .O(n524bar),
    .I0(in_33bar),
    .I1(in_27bar)
  );
  //OR U454
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U454 (
    .O(n568),
    .I0(n522),
    .I1(n521)
  );
  //AND U454bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U454bar (
    .O(n568bar),
    .I0(n522bar),
    .I1(n521bar)
  );
  //OR U455
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U455 (
    .O(n521),
    .I0(in[145]),
    .I1(in[126])
  );
  //AND U455bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U455bar (
    .O(n521bar),
    .I0(inbar[145]),
    .I1(inbar[126])
  );
  //OR U456
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U456 (
    .O(n522),
    .I0(in[169]),
    .I1(n520)
  );
  //AND U456bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U456bar (
    .O(n522bar),
    .I0(inbar[169]),
    .I1(n520bar)
  );
  //OR U457
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U457 (
    .O(n520),
    .I0(in[221]),
    .I1(in[172])
  );
  //AND U457bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U457bar (
    .O(n520bar),
    .I0(inbar[221]),
    .I1(inbar[172])
  );
  //OR U458
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U458 (
    .O(n570),
    .I0(n519),
    .I1(n518)
  );
  //AND U458bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U458bar (
    .O(n570bar),
    .I0(n519bar),
    .I1(n518bar)
  );
  //OR U459
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U459 (
    .O(n518),
    .I0(n517),
    .I1(n516)
  );
  //AND U459bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U459bar (
    .O(n518bar),
    .I0(n517bar),
    .I1(n516bar)
  );
  //OR U460
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U460 (
    .O(n516),
    .I0(in[241]),
    .I1(in[224])
  );
  //AND U460bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U460bar (
    .O(n516bar),
    .I0(inbar[241]),
    .I1(inbar[224])
  );
  //OR U461
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U461 (
    .O(n517),
    .I0(in[86]),
    .I1(n515)
  );
  //AND U461bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U461bar (
    .O(n517bar),
    .I0(inbar[86]),
    .I1(n515bar)
  );
  //OR U462
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U462 (
    .O(n515),
    .I0(in_43),
    .I1(in_34)
  );
  //AND U462bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U462bar (
    .O(n515bar),
    .I0(in_43bar),
    .I1(in_34bar)
  );
  //OR U463
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U463 (
    .O(n519),
    .I0(n514),
    .I1(n513)
  );
  //AND U463bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U463bar (
    .O(n519bar),
    .I0(n514bar),
    .I1(n513bar)
  );
  //OR U464
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U464 (
    .O(n513),
    .I0(in_65),
    .I1(in_51)
  );
  //AND U464bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U464bar (
    .O(n513bar),
    .I0(in_65bar),
    .I1(in_51bar)
  );
  //OR U465
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U465 (
    .O(n514),
    .I0(in_75),
    .I1(n512)
  );
  //AND U465bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U465bar (
    .O(n514bar),
    .I0(in_75bar),
    .I1(n512bar)
  );
  //OR U466
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U466 (
    .O(n512),
    .I0(in_81),
    .I1(in_77)
  );
  //AND U466bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U466bar (
    .O(n512bar),
    .I0(in_81bar),
    .I1(in_77bar)
  );
  //OR U467
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U467 (
    .O(n778),
    .I0(n511),
    .I1(n510)
  );
  //AND U467bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U467bar (
    .O(n778bar),
    .I0(n511bar),
    .I1(n510bar)
  );
  //OR U468
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U468 (
    .O(n510),
    .I0(n509),
    .I1(n508)
  );
  //AND U468bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U468bar (
    .O(n510bar),
    .I0(n509bar),
    .I1(n508bar)
  );
  //OR U469
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U469 (
    .O(n508),
    .I0(n507),
    .I1(n506)
  );
  //AND U469bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U469bar (
    .O(n508bar),
    .I0(n507bar),
    .I1(n506bar)
  );
  //OR U470
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U470 (
    .O(n506),
    .I0(in[107]),
    .I1(in[101])
  );
  //AND U470bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U470bar (
    .O(n506bar),
    .I0(inbar[107]),
    .I1(inbar[101])
  );
  //OR U471
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U471 (
    .O(n507),
    .I0(in[139]),
    .I1(in[132])
  );
  //AND U471bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U471bar (
    .O(n507bar),
    .I0(inbar[139]),
    .I1(inbar[132])
  );
  //OR U472
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U472 (
    .O(n509),
    .I0(n505),
    .I1(n504)
  );
  //AND U472bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U472bar (
    .O(n509bar),
    .I0(n505bar),
    .I1(n504bar)
  );
  //OR U473
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U473 (
    .O(n504),
    .I0(in[146]),
    .I1(in[141])
  );
  //AND U473bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U473bar (
    .O(n504bar),
    .I0(inbar[146]),
    .I1(inbar[141])
  );
  //OR U474
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U474 (
    .O(n505),
    .I0(in[203]),
    .I1(in[179])
  );
  //AND U474bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U474bar (
    .O(n505bar),
    .I0(inbar[203]),
    .I1(inbar[179])
  );
  //OR U475
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U475 (
    .O(n511),
    .I0(n503),
    .I1(n502)
  );
  //AND U475bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U475bar (
    .O(n511bar),
    .I0(n503bar),
    .I1(n502bar)
  );
  //OR U476
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U476 (
    .O(n502),
    .I0(n501),
    .I1(n500)
  );
  //AND U476bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U476bar (
    .O(n502bar),
    .I0(n501bar),
    .I1(n500bar)
  );
  //OR U477
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U477 (
    .O(n500),
    .I0(in[243]),
    .I1(in[222])
  );
  //AND U477bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U477bar (
    .O(n500bar),
    .I0(inbar[243]),
    .I1(inbar[222])
  );
  //OR U478
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U478 (
    .O(n501),
    .I0(in[251]),
    .I1(in[250])
  );
  //AND U478bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U478bar (
    .O(n501bar),
    .I0(inbar[251]),
    .I1(inbar[250])
  );
  //OR U479
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U479 (
    .O(n503),
    .I0(n499),
    .I1(n498)
  );
  //AND U479bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U479bar (
    .O(n503bar),
    .I0(n499bar),
    .I1(n498bar)
  );
  //OR U480
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U480 (
    .O(n498),
    .I0(in_37),
    .I1(in_19)
  );
  //AND U480bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U480bar (
    .O(n498bar),
    .I0(in_37bar),
    .I1(in_19bar)
  );
  //OR U481
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U481 (
    .O(n499),
    .I0(in_78),
    .I1(in_6)
  );
  //AND U481bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U481bar (
    .O(n499bar),
    .I0(in_78bar),
    .I1(in_6bar)
  );
  //OR U482
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U482 (
    .O(n603),
    .I0(n497),
    .I1(n496)
  );
  //AND U482bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U482bar (
    .O(n603bar),
    .I0(n497bar),
    .I1(n496bar)
  );
  //OR U483
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U483 (
    .O(n496),
    .I0(in[112]),
    .I1(in[102])
  );
  //AND U483bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U483bar (
    .O(n496bar),
    .I0(inbar[112]),
    .I1(inbar[102])
  );
  //OR U484
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U484 (
    .O(n497),
    .I0(in[123]),
    .I1(n495)
  );
  //AND U484bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U484bar (
    .O(n497bar),
    .I0(inbar[123]),
    .I1(n495bar)
  );
  //OR U485
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U485 (
    .O(n495),
    .I0(in[143]),
    .I1(in[130])
  );
  //AND U485bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U485bar (
    .O(n495bar),
    .I0(inbar[143]),
    .I1(inbar[130])
  );
  //OR U486
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U486 (
    .O(n605),
    .I0(n494),
    .I1(n493)
  );
  //AND U486bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U486bar (
    .O(n605bar),
    .I0(n494bar),
    .I1(n493bar)
  );
  //OR U487
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U487 (
    .O(n493),
    .I0(n492),
    .I1(n491)
  );
  //AND U487bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U487bar (
    .O(n493bar),
    .I0(n492bar),
    .I1(n491bar)
  );
  //OR U488
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U488 (
    .O(n491),
    .I0(in[216]),
    .I1(in[213])
  );
  //AND U488bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U488bar (
    .O(n491bar),
    .I0(inbar[216]),
    .I1(inbar[213])
  );
  //OR U489
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U489 (
    .O(n492),
    .I0(in[227]),
    .I1(n490)
  );
  //AND U489bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U489bar (
    .O(n492bar),
    .I0(inbar[227]),
    .I1(n490bar)
  );
  //OR U490
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U490 (
    .O(n490),
    .I0(in_0),
    .I1(in[248])
  );
  //AND U490bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U490bar (
    .O(n490bar),
    .I0(in_0bar),
    .I1(inbar[248])
  );
  //OR U491
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U491 (
    .O(n494),
    .I0(n489),
    .I1(n488)
  );
  //AND U491bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U491bar (
    .O(n494bar),
    .I0(n489bar),
    .I1(n488bar)
  );
  //OR U492
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U492 (
    .O(n488),
    .I0(in_46),
    .I1(in_44)
  );
  //AND U492bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U492bar (
    .O(n488bar),
    .I0(in_46bar),
    .I1(in_44bar)
  );
  //OR U493
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U493 (
    .O(n489),
    .I0(in_50),
    .I1(n487)
  );
  //AND U493bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U493bar (
    .O(n489bar),
    .I0(in_50bar),
    .I1(n487bar)
  );
  //OR U494
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U494 (
    .O(n487),
    .I0(in_9),
    .I1(in_80)
  );
  //AND U494bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U494bar (
    .O(n487bar),
    .I0(in_9bar),
    .I1(in_80bar)
  );
endmodule

module sBox_6 ( in, out );

  input wire [7:0] in;
//input_done

  output wire [7:0] out;
//output_done

  wire [255:0] decodeOut;
//wire_done

  decode_6 dec ( .in(in), .out(decodeOut) );
  encode_6 enc ( .in(decodeOut), .out(out) );
endmodule

module CD2_25 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD2_26 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD2_27 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD2_28 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD4_13 ( a, b, y );

  input wire [3:0] a;
  input wire [3:0] b;
  wire [3:0] abar;
  wire [3:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
//input_done

  output wire [15:0] y;
  wire [15:0] ybar;
//output_done

//wire_done

  //AND U1
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1 (
    .O(y[9]),
    .I0(b[1]),
    .I1(a[2])
  );
  //OR U1bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1bar (
    .O(ybar[9]),
    .I0(bbar[1]),
    .I1(abar[2])
  );
  //AND U2
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2 (
    .O(y[8]),
    .I0(b[0]),
    .I1(a[2])
  );
  //OR U2bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2bar (
    .O(ybar[8]),
    .I0(bbar[0]),
    .I1(abar[2])
  );
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[7]),
    .I0(b[3]),
    .I1(a[1])
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[7]),
    .I0(bbar[3]),
    .I1(abar[1])
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[6]),
    .I0(b[2]),
    .I1(a[1])
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[6]),
    .I0(bbar[2]),
    .I1(abar[1])
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[5]),
    .I0(a[1]),
    .I1(b[1])
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[5]),
    .I0(abar[1]),
    .I1(bbar[1])
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[4]),
    .I0(a[1]),
    .I1(b[0])
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[4]),
    .I0(abar[1]),
    .I1(bbar[0])
  );
  //AND U7
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7 (
    .O(y[3]),
    .I0(a[0]),
    .I1(b[3])
  );
  //OR U7bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7bar (
    .O(ybar[3]),
    .I0(abar[0]),
    .I1(bbar[3])
  );
  //AND U8
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8 (
    .O(y[2]),
    .I0(a[0]),
    .I1(b[2])
  );
  //OR U8bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8bar (
    .O(ybar[2]),
    .I0(abar[0]),
    .I1(bbar[2])
  );
  //AND U9
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9 (
    .O(y[1]),
    .I0(a[0]),
    .I1(b[1])
  );
  //OR U9bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9bar (
    .O(ybar[1]),
    .I0(abar[0]),
    .I1(bbar[1])
  );
  //AND U10
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10 (
    .O(y[15]),
    .I0(a[3]),
    .I1(b[3])
  );
  //OR U10bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10bar (
    .O(ybar[15]),
    .I0(abar[3]),
    .I1(bbar[3])
  );
  //AND U11
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11 (
    .O(y[14]),
    .I0(a[3]),
    .I1(b[2])
  );
  //OR U11bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11bar (
    .O(ybar[14]),
    .I0(abar[3]),
    .I1(bbar[2])
  );
  //AND U12
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12 (
    .O(y[13]),
    .I0(a[3]),
    .I1(b[1])
  );
  //OR U12bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12bar (
    .O(ybar[13]),
    .I0(abar[3]),
    .I1(bbar[1])
  );
  //AND U13
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13 (
    .O(y[12]),
    .I0(a[3]),
    .I1(b[0])
  );
  //OR U13bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13bar (
    .O(ybar[12]),
    .I0(abar[3]),
    .I1(bbar[0])
  );
  //AND U14
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14 (
    .O(y[11]),
    .I0(b[3]),
    .I1(a[2])
  );
  //OR U14bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14bar (
    .O(ybar[11]),
    .I0(bbar[3]),
    .I1(abar[2])
  );
  //AND U15
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15 (
    .O(y[10]),
    .I0(b[2]),
    .I1(a[2])
  );
  //OR U15bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15bar (
    .O(ybar[10]),
    .I0(bbar[2]),
    .I1(abar[2])
  );
  //AND U16
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16 (
    .O(y[0]),
    .I0(a[0]),
    .I1(b[0])
  );
  //OR U16bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16bar (
    .O(ybar[0]),
    .I0(abar[0]),
    .I1(bbar[0])
  );
endmodule

module CD4_14 ( a, b, y );

  input wire [3:0] a;
  input wire [3:0] b;
  wire [3:0] abar;
  wire [3:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
//input_done

  output wire [15:0] y;
  wire [15:0] ybar;
//output_done

//wire_done

  //AND U1
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1 (
    .O(y[9]),
    .I0(b[1]),
    .I1(a[2])
  );
  //OR U1bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1bar (
    .O(ybar[9]),
    .I0(bbar[1]),
    .I1(abar[2])
  );
  //AND U2
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2 (
    .O(y[8]),
    .I0(b[0]),
    .I1(a[2])
  );
  //OR U2bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2bar (
    .O(ybar[8]),
    .I0(bbar[0]),
    .I1(abar[2])
  );
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[7]),
    .I0(b[3]),
    .I1(a[1])
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[7]),
    .I0(bbar[3]),
    .I1(abar[1])
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[6]),
    .I0(b[2]),
    .I1(a[1])
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[6]),
    .I0(bbar[2]),
    .I1(abar[1])
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[5]),
    .I0(a[1]),
    .I1(b[1])
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[5]),
    .I0(abar[1]),
    .I1(bbar[1])
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[4]),
    .I0(a[1]),
    .I1(b[0])
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[4]),
    .I0(abar[1]),
    .I1(bbar[0])
  );
  //AND U7
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7 (
    .O(y[3]),
    .I0(a[0]),
    .I1(b[3])
  );
  //OR U7bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7bar (
    .O(ybar[3]),
    .I0(abar[0]),
    .I1(bbar[3])
  );
  //AND U8
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8 (
    .O(y[2]),
    .I0(a[0]),
    .I1(b[2])
  );
  //OR U8bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8bar (
    .O(ybar[2]),
    .I0(abar[0]),
    .I1(bbar[2])
  );
  //AND U9
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9 (
    .O(y[1]),
    .I0(a[0]),
    .I1(b[1])
  );
  //OR U9bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9bar (
    .O(ybar[1]),
    .I0(abar[0]),
    .I1(bbar[1])
  );
  //AND U10
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10 (
    .O(y[15]),
    .I0(a[3]),
    .I1(b[3])
  );
  //OR U10bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10bar (
    .O(ybar[15]),
    .I0(abar[3]),
    .I1(bbar[3])
  );
  //AND U11
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11 (
    .O(y[14]),
    .I0(a[3]),
    .I1(b[2])
  );
  //OR U11bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11bar (
    .O(ybar[14]),
    .I0(abar[3]),
    .I1(bbar[2])
  );
  //AND U12
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12 (
    .O(y[13]),
    .I0(a[3]),
    .I1(b[1])
  );
  //OR U12bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12bar (
    .O(ybar[13]),
    .I0(abar[3]),
    .I1(bbar[1])
  );
  //AND U13
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13 (
    .O(y[12]),
    .I0(a[3]),
    .I1(b[0])
  );
  //OR U13bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13bar (
    .O(ybar[12]),
    .I0(abar[3]),
    .I1(bbar[0])
  );
  //AND U14
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14 (
    .O(y[11]),
    .I0(b[3]),
    .I1(a[2])
  );
  //OR U14bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14bar (
    .O(ybar[11]),
    .I0(bbar[3]),
    .I1(abar[2])
  );
  //AND U15
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15 (
    .O(y[10]),
    .I0(b[2]),
    .I1(a[2])
  );
  //OR U15bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15bar (
    .O(ybar[10]),
    .I0(bbar[2]),
    .I1(abar[2])
  );
  //AND U16
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16 (
    .O(y[0]),
    .I0(a[0]),
    .I1(b[0])
  );
  //OR U16bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16bar (
    .O(ybar[0]),
    .I0(abar[0]),
    .I1(bbar[0])
  );
endmodule

module CD16_7 ( a, b, y );

  input wire [15:0] a;
  input wire [15:0] b;
  wire [15:0] abar;
  wire [15:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign abar[8] = ~a[8];
  assign abar[9] = ~a[9];
  assign abar[10] = ~a[10];
  assign abar[11] = ~a[11];
  assign abar[12] = ~a[12];
  assign abar[13] = ~a[13];
  assign abar[14] = ~a[14];
  assign abar[15] = ~a[15];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign bbar[8] = ~b[8];
  assign bbar[9] = ~b[9];
  assign bbar[10] = ~b[10];
  assign bbar[11] = ~b[11];
  assign bbar[12] = ~b[12];
  assign bbar[13] = ~b[13];
  assign bbar[14] = ~b[14];
  assign bbar[15] = ~b[15];
//input_done

  output wire [255:0] y;
  wire [255:0] ybar;
//output_done

//wire_done

  //AND U1
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1 (
    .O(y[9]),
    .I0(b[9]),
    .I1(a[0])
  );
  //OR U1bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1bar (
    .O(ybar[9]),
    .I0(bbar[9]),
    .I1(abar[0])
  );
  //AND U2
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2 (
    .O(y[99]),
    .I0(b[3]),
    .I1(a[6])
  );
  //OR U2bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2bar (
    .O(ybar[99]),
    .I0(bbar[3]),
    .I1(abar[6])
  );
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[98]),
    .I0(b[2]),
    .I1(a[6])
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[98]),
    .I0(bbar[2]),
    .I1(abar[6])
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[97]),
    .I0(b[1]),
    .I1(a[6])
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[97]),
    .I0(bbar[1]),
    .I1(abar[6])
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[96]),
    .I0(b[0]),
    .I1(a[6])
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[96]),
    .I0(bbar[0]),
    .I1(abar[6])
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[95]),
    .I0(b[15]),
    .I1(a[5])
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[95]),
    .I0(bbar[15]),
    .I1(abar[5])
  );
  //AND U7
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7 (
    .O(y[94]),
    .I0(b[14]),
    .I1(a[5])
  );
  //OR U7bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7bar (
    .O(ybar[94]),
    .I0(bbar[14]),
    .I1(abar[5])
  );
  //AND U8
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8 (
    .O(y[93]),
    .I0(b[13]),
    .I1(a[5])
  );
  //OR U8bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8bar (
    .O(ybar[93]),
    .I0(bbar[13]),
    .I1(abar[5])
  );
  //AND U9
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9 (
    .O(y[92]),
    .I0(b[12]),
    .I1(a[5])
  );
  //OR U9bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9bar (
    .O(ybar[92]),
    .I0(bbar[12]),
    .I1(abar[5])
  );
  //AND U10
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10 (
    .O(y[91]),
    .I0(b[11]),
    .I1(a[5])
  );
  //OR U10bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10bar (
    .O(ybar[91]),
    .I0(bbar[11]),
    .I1(abar[5])
  );
  //AND U11
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11 (
    .O(y[90]),
    .I0(b[10]),
    .I1(a[5])
  );
  //OR U11bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11bar (
    .O(ybar[90]),
    .I0(bbar[10]),
    .I1(abar[5])
  );
  //AND U12
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12 (
    .O(y[8]),
    .I0(b[8]),
    .I1(a[0])
  );
  //OR U12bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12bar (
    .O(ybar[8]),
    .I0(bbar[8]),
    .I1(abar[0])
  );
  //AND U13
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13 (
    .O(y[89]),
    .I0(a[5]),
    .I1(b[9])
  );
  //OR U13bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13bar (
    .O(ybar[89]),
    .I0(abar[5]),
    .I1(bbar[9])
  );
  //AND U14
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14 (
    .O(y[88]),
    .I0(b[8]),
    .I1(a[5])
  );
  //OR U14bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14bar (
    .O(ybar[88]),
    .I0(bbar[8]),
    .I1(abar[5])
  );
  //AND U15
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15 (
    .O(y[87]),
    .I0(b[7]),
    .I1(a[5])
  );
  //OR U15bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15bar (
    .O(ybar[87]),
    .I0(bbar[7]),
    .I1(abar[5])
  );
  //AND U16
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16 (
    .O(y[86]),
    .I0(b[6]),
    .I1(a[5])
  );
  //OR U16bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16bar (
    .O(ybar[86]),
    .I0(bbar[6]),
    .I1(abar[5])
  );
  //AND U17
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U17 (
    .O(y[85]),
    .I0(b[5]),
    .I1(a[5])
  );
  //OR U17bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U17bar (
    .O(ybar[85]),
    .I0(bbar[5]),
    .I1(abar[5])
  );
  //AND U18
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U18 (
    .O(y[84]),
    .I0(b[4]),
    .I1(a[5])
  );
  //OR U18bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U18bar (
    .O(ybar[84]),
    .I0(bbar[4]),
    .I1(abar[5])
  );
  //AND U19
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U19 (
    .O(y[83]),
    .I0(a[5]),
    .I1(b[3])
  );
  //OR U19bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U19bar (
    .O(ybar[83]),
    .I0(abar[5]),
    .I1(bbar[3])
  );
  //AND U20
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U20 (
    .O(y[82]),
    .I0(a[5]),
    .I1(b[2])
  );
  //OR U20bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U20bar (
    .O(ybar[82]),
    .I0(abar[5]),
    .I1(bbar[2])
  );
  //AND U21
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U21 (
    .O(y[81]),
    .I0(a[5]),
    .I1(b[1])
  );
  //OR U21bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U21bar (
    .O(ybar[81]),
    .I0(abar[5]),
    .I1(bbar[1])
  );
  //AND U22
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U22 (
    .O(y[80]),
    .I0(a[5]),
    .I1(b[0])
  );
  //OR U22bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U22bar (
    .O(ybar[80]),
    .I0(abar[5]),
    .I1(bbar[0])
  );
  //AND U23
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U23 (
    .O(y[7]),
    .I0(b[7]),
    .I1(a[0])
  );
  //OR U23bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U23bar (
    .O(ybar[7]),
    .I0(bbar[7]),
    .I1(abar[0])
  );
  //AND U24
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U24 (
    .O(y[79]),
    .I0(a[4]),
    .I1(b[15])
  );
  //OR U24bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U24bar (
    .O(ybar[79]),
    .I0(abar[4]),
    .I1(bbar[15])
  );
  //AND U25
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U25 (
    .O(y[78]),
    .I0(a[4]),
    .I1(b[14])
  );
  //OR U25bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U25bar (
    .O(ybar[78]),
    .I0(abar[4]),
    .I1(bbar[14])
  );
  //AND U26
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U26 (
    .O(y[77]),
    .I0(a[4]),
    .I1(b[13])
  );
  //OR U26bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U26bar (
    .O(ybar[77]),
    .I0(abar[4]),
    .I1(bbar[13])
  );
  //AND U27
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U27 (
    .O(y[76]),
    .I0(a[4]),
    .I1(b[12])
  );
  //OR U27bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U27bar (
    .O(ybar[76]),
    .I0(abar[4]),
    .I1(bbar[12])
  );
  //AND U28
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U28 (
    .O(y[75]),
    .I0(a[4]),
    .I1(b[11])
  );
  //OR U28bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U28bar (
    .O(ybar[75]),
    .I0(abar[4]),
    .I1(bbar[11])
  );
  //AND U29
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U29 (
    .O(y[74]),
    .I0(a[4]),
    .I1(b[10])
  );
  //OR U29bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U29bar (
    .O(ybar[74]),
    .I0(abar[4]),
    .I1(bbar[10])
  );
  //AND U30
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U30 (
    .O(y[73]),
    .I0(a[4]),
    .I1(b[9])
  );
  //OR U30bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U30bar (
    .O(ybar[73]),
    .I0(abar[4]),
    .I1(bbar[9])
  );
  //AND U31
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U31 (
    .O(y[72]),
    .I0(a[4]),
    .I1(b[8])
  );
  //OR U31bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U31bar (
    .O(ybar[72]),
    .I0(abar[4]),
    .I1(bbar[8])
  );
  //AND U32
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U32 (
    .O(y[71]),
    .I0(a[4]),
    .I1(b[7])
  );
  //OR U32bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U32bar (
    .O(ybar[71]),
    .I0(abar[4]),
    .I1(bbar[7])
  );
  //AND U33
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U33 (
    .O(y[70]),
    .I0(a[4]),
    .I1(b[6])
  );
  //OR U33bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U33bar (
    .O(ybar[70]),
    .I0(abar[4]),
    .I1(bbar[6])
  );
  //AND U34
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U34 (
    .O(y[6]),
    .I0(b[6]),
    .I1(a[0])
  );
  //OR U34bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U34bar (
    .O(ybar[6]),
    .I0(bbar[6]),
    .I1(abar[0])
  );
  //AND U35
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U35 (
    .O(y[69]),
    .I0(a[4]),
    .I1(b[5])
  );
  //OR U35bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U35bar (
    .O(ybar[69]),
    .I0(abar[4]),
    .I1(bbar[5])
  );
  //AND U36
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U36 (
    .O(y[68]),
    .I0(a[4]),
    .I1(b[4])
  );
  //OR U36bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U36bar (
    .O(ybar[68]),
    .I0(abar[4]),
    .I1(bbar[4])
  );
  //AND U37
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U37 (
    .O(y[67]),
    .I0(a[4]),
    .I1(b[3])
  );
  //OR U37bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U37bar (
    .O(ybar[67]),
    .I0(abar[4]),
    .I1(bbar[3])
  );
  //AND U38
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U38 (
    .O(y[66]),
    .I0(a[4]),
    .I1(b[2])
  );
  //OR U38bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U38bar (
    .O(ybar[66]),
    .I0(abar[4]),
    .I1(bbar[2])
  );
  //AND U39
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U39 (
    .O(y[65]),
    .I0(a[4]),
    .I1(b[1])
  );
  //OR U39bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U39bar (
    .O(ybar[65]),
    .I0(abar[4]),
    .I1(bbar[1])
  );
  //AND U40
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U40 (
    .O(y[64]),
    .I0(a[4]),
    .I1(b[0])
  );
  //OR U40bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U40bar (
    .O(ybar[64]),
    .I0(abar[4]),
    .I1(bbar[0])
  );
  //AND U41
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U41 (
    .O(y[63]),
    .I0(a[3]),
    .I1(b[15])
  );
  //OR U41bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U41bar (
    .O(ybar[63]),
    .I0(abar[3]),
    .I1(bbar[15])
  );
  //AND U42
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U42 (
    .O(y[62]),
    .I0(a[3]),
    .I1(b[14])
  );
  //OR U42bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U42bar (
    .O(ybar[62]),
    .I0(abar[3]),
    .I1(bbar[14])
  );
  //AND U43
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U43 (
    .O(y[61]),
    .I0(a[3]),
    .I1(b[13])
  );
  //OR U43bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U43bar (
    .O(ybar[61]),
    .I0(abar[3]),
    .I1(bbar[13])
  );
  //AND U44
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U44 (
    .O(y[60]),
    .I0(a[3]),
    .I1(b[12])
  );
  //OR U44bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U44bar (
    .O(ybar[60]),
    .I0(abar[3]),
    .I1(bbar[12])
  );
  //AND U45
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U45 (
    .O(y[5]),
    .I0(b[5]),
    .I1(a[0])
  );
  //OR U45bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U45bar (
    .O(ybar[5]),
    .I0(bbar[5]),
    .I1(abar[0])
  );
  //AND U46
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U46 (
    .O(y[59]),
    .I0(a[3]),
    .I1(b[11])
  );
  //OR U46bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U46bar (
    .O(ybar[59]),
    .I0(abar[3]),
    .I1(bbar[11])
  );
  //AND U47
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U47 (
    .O(y[58]),
    .I0(a[3]),
    .I1(b[10])
  );
  //OR U47bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U47bar (
    .O(ybar[58]),
    .I0(abar[3]),
    .I1(bbar[10])
  );
  //AND U48
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U48 (
    .O(y[57]),
    .I0(a[3]),
    .I1(b[9])
  );
  //OR U48bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U48bar (
    .O(ybar[57]),
    .I0(abar[3]),
    .I1(bbar[9])
  );
  //AND U49
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U49 (
    .O(y[56]),
    .I0(a[3]),
    .I1(b[8])
  );
  //OR U49bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U49bar (
    .O(ybar[56]),
    .I0(abar[3]),
    .I1(bbar[8])
  );
  //AND U50
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U50 (
    .O(y[55]),
    .I0(a[3]),
    .I1(b[7])
  );
  //OR U50bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U50bar (
    .O(ybar[55]),
    .I0(abar[3]),
    .I1(bbar[7])
  );
  //AND U51
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U51 (
    .O(y[54]),
    .I0(a[3]),
    .I1(b[6])
  );
  //OR U51bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U51bar (
    .O(ybar[54]),
    .I0(abar[3]),
    .I1(bbar[6])
  );
  //AND U52
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U52 (
    .O(y[53]),
    .I0(a[3]),
    .I1(b[5])
  );
  //OR U52bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U52bar (
    .O(ybar[53]),
    .I0(abar[3]),
    .I1(bbar[5])
  );
  //AND U53
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U53 (
    .O(y[52]),
    .I0(a[3]),
    .I1(b[4])
  );
  //OR U53bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U53bar (
    .O(ybar[52]),
    .I0(abar[3]),
    .I1(bbar[4])
  );
  //AND U54
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U54 (
    .O(y[51]),
    .I0(a[3]),
    .I1(b[3])
  );
  //OR U54bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U54bar (
    .O(ybar[51]),
    .I0(abar[3]),
    .I1(bbar[3])
  );
  //AND U55
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U55 (
    .O(y[50]),
    .I0(a[3]),
    .I1(b[2])
  );
  //OR U55bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U55bar (
    .O(ybar[50]),
    .I0(abar[3]),
    .I1(bbar[2])
  );
  //AND U56
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U56 (
    .O(y[4]),
    .I0(b[4]),
    .I1(a[0])
  );
  //OR U56bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U56bar (
    .O(ybar[4]),
    .I0(bbar[4]),
    .I1(abar[0])
  );
  //AND U57
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U57 (
    .O(y[49]),
    .I0(a[3]),
    .I1(b[1])
  );
  //OR U57bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U57bar (
    .O(ybar[49]),
    .I0(abar[3]),
    .I1(bbar[1])
  );
  //AND U58
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U58 (
    .O(y[48]),
    .I0(a[3]),
    .I1(b[0])
  );
  //OR U58bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U58bar (
    .O(ybar[48]),
    .I0(abar[3]),
    .I1(bbar[0])
  );
  //AND U59
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U59 (
    .O(y[47]),
    .I0(a[2]),
    .I1(b[15])
  );
  //OR U59bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U59bar (
    .O(ybar[47]),
    .I0(abar[2]),
    .I1(bbar[15])
  );
  //AND U60
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U60 (
    .O(y[46]),
    .I0(a[2]),
    .I1(b[14])
  );
  //OR U60bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U60bar (
    .O(ybar[46]),
    .I0(abar[2]),
    .I1(bbar[14])
  );
  //AND U61
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U61 (
    .O(y[45]),
    .I0(a[2]),
    .I1(b[13])
  );
  //OR U61bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U61bar (
    .O(ybar[45]),
    .I0(abar[2]),
    .I1(bbar[13])
  );
  //AND U62
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U62 (
    .O(y[44]),
    .I0(a[2]),
    .I1(b[12])
  );
  //OR U62bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U62bar (
    .O(ybar[44]),
    .I0(abar[2]),
    .I1(bbar[12])
  );
  //AND U63
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U63 (
    .O(y[43]),
    .I0(a[2]),
    .I1(b[11])
  );
  //OR U63bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U63bar (
    .O(ybar[43]),
    .I0(abar[2]),
    .I1(bbar[11])
  );
  //AND U64
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U64 (
    .O(y[42]),
    .I0(a[2]),
    .I1(b[10])
  );
  //OR U64bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U64bar (
    .O(ybar[42]),
    .I0(abar[2]),
    .I1(bbar[10])
  );
  //AND U65
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U65 (
    .O(y[41]),
    .I0(a[2]),
    .I1(b[9])
  );
  //OR U65bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U65bar (
    .O(ybar[41]),
    .I0(abar[2]),
    .I1(bbar[9])
  );
  //AND U66
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U66 (
    .O(y[40]),
    .I0(a[2]),
    .I1(b[8])
  );
  //OR U66bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U66bar (
    .O(ybar[40]),
    .I0(abar[2]),
    .I1(bbar[8])
  );
  //AND U67
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U67 (
    .O(y[3]),
    .I0(b[3]),
    .I1(a[0])
  );
  //OR U67bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U67bar (
    .O(ybar[3]),
    .I0(bbar[3]),
    .I1(abar[0])
  );
  //AND U68
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U68 (
    .O(y[39]),
    .I0(a[2]),
    .I1(b[7])
  );
  //OR U68bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U68bar (
    .O(ybar[39]),
    .I0(abar[2]),
    .I1(bbar[7])
  );
  //AND U69
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U69 (
    .O(y[38]),
    .I0(a[2]),
    .I1(b[6])
  );
  //OR U69bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U69bar (
    .O(ybar[38]),
    .I0(abar[2]),
    .I1(bbar[6])
  );
  //AND U70
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U70 (
    .O(y[37]),
    .I0(a[2]),
    .I1(b[5])
  );
  //OR U70bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U70bar (
    .O(ybar[37]),
    .I0(abar[2]),
    .I1(bbar[5])
  );
  //AND U71
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U71 (
    .O(y[36]),
    .I0(a[2]),
    .I1(b[4])
  );
  //OR U71bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U71bar (
    .O(ybar[36]),
    .I0(abar[2]),
    .I1(bbar[4])
  );
  //AND U72
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U72 (
    .O(y[35]),
    .I0(a[2]),
    .I1(b[3])
  );
  //OR U72bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U72bar (
    .O(ybar[35]),
    .I0(abar[2]),
    .I1(bbar[3])
  );
  //AND U73
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U73 (
    .O(y[34]),
    .I0(a[2]),
    .I1(b[2])
  );
  //OR U73bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U73bar (
    .O(ybar[34]),
    .I0(abar[2]),
    .I1(bbar[2])
  );
  //AND U74
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U74 (
    .O(y[33]),
    .I0(a[2]),
    .I1(b[1])
  );
  //OR U74bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U74bar (
    .O(ybar[33]),
    .I0(abar[2]),
    .I1(bbar[1])
  );
  //AND U75
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U75 (
    .O(y[32]),
    .I0(a[2]),
    .I1(b[0])
  );
  //OR U75bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U75bar (
    .O(ybar[32]),
    .I0(abar[2]),
    .I1(bbar[0])
  );
  //AND U76
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U76 (
    .O(y[31]),
    .I0(a[1]),
    .I1(b[15])
  );
  //OR U76bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U76bar (
    .O(ybar[31]),
    .I0(abar[1]),
    .I1(bbar[15])
  );
  //AND U77
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U77 (
    .O(y[30]),
    .I0(a[1]),
    .I1(b[14])
  );
  //OR U77bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U77bar (
    .O(ybar[30]),
    .I0(abar[1]),
    .I1(bbar[14])
  );
  //AND U78
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U78 (
    .O(y[2]),
    .I0(b[2]),
    .I1(a[0])
  );
  //OR U78bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U78bar (
    .O(ybar[2]),
    .I0(bbar[2]),
    .I1(abar[0])
  );
  //AND U79
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U79 (
    .O(y[29]),
    .I0(a[1]),
    .I1(b[13])
  );
  //OR U79bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U79bar (
    .O(ybar[29]),
    .I0(abar[1]),
    .I1(bbar[13])
  );
  //AND U80
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U80 (
    .O(y[28]),
    .I0(a[1]),
    .I1(b[12])
  );
  //OR U80bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U80bar (
    .O(ybar[28]),
    .I0(abar[1]),
    .I1(bbar[12])
  );
  //AND U81
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U81 (
    .O(y[27]),
    .I0(a[1]),
    .I1(b[11])
  );
  //OR U81bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U81bar (
    .O(ybar[27]),
    .I0(abar[1]),
    .I1(bbar[11])
  );
  //AND U82
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U82 (
    .O(y[26]),
    .I0(a[1]),
    .I1(b[10])
  );
  //OR U82bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U82bar (
    .O(ybar[26]),
    .I0(abar[1]),
    .I1(bbar[10])
  );
  //AND U83
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U83 (
    .O(y[25]),
    .I0(a[1]),
    .I1(b[9])
  );
  //OR U83bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U83bar (
    .O(ybar[25]),
    .I0(abar[1]),
    .I1(bbar[9])
  );
  //AND U84
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U84 (
    .O(y[255]),
    .I0(a[15]),
    .I1(b[15])
  );
  //OR U84bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U84bar (
    .O(ybar[255]),
    .I0(abar[15]),
    .I1(bbar[15])
  );
  //AND U85
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U85 (
    .O(y[254]),
    .I0(a[15]),
    .I1(b[14])
  );
  //OR U85bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U85bar (
    .O(ybar[254]),
    .I0(abar[15]),
    .I1(bbar[14])
  );
  //AND U86
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U86 (
    .O(y[253]),
    .I0(a[15]),
    .I1(b[13])
  );
  //OR U86bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U86bar (
    .O(ybar[253]),
    .I0(abar[15]),
    .I1(bbar[13])
  );
  //AND U87
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U87 (
    .O(y[252]),
    .I0(a[15]),
    .I1(b[12])
  );
  //OR U87bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U87bar (
    .O(ybar[252]),
    .I0(abar[15]),
    .I1(bbar[12])
  );
  //AND U88
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U88 (
    .O(y[251]),
    .I0(a[15]),
    .I1(b[11])
  );
  //OR U88bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U88bar (
    .O(ybar[251]),
    .I0(abar[15]),
    .I1(bbar[11])
  );
  //AND U89
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U89 (
    .O(y[250]),
    .I0(a[15]),
    .I1(b[10])
  );
  //OR U89bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U89bar (
    .O(ybar[250]),
    .I0(abar[15]),
    .I1(bbar[10])
  );
  //AND U90
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U90 (
    .O(y[24]),
    .I0(a[1]),
    .I1(b[8])
  );
  //OR U90bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U90bar (
    .O(ybar[24]),
    .I0(abar[1]),
    .I1(bbar[8])
  );
  //AND U91
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U91 (
    .O(y[249]),
    .I0(a[15]),
    .I1(b[9])
  );
  //OR U91bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U91bar (
    .O(ybar[249]),
    .I0(abar[15]),
    .I1(bbar[9])
  );
  //AND U92
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U92 (
    .O(y[248]),
    .I0(a[15]),
    .I1(b[8])
  );
  //OR U92bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U92bar (
    .O(ybar[248]),
    .I0(abar[15]),
    .I1(bbar[8])
  );
  //AND U93
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U93 (
    .O(y[247]),
    .I0(a[15]),
    .I1(b[7])
  );
  //OR U93bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U93bar (
    .O(ybar[247]),
    .I0(abar[15]),
    .I1(bbar[7])
  );
  //AND U94
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U94 (
    .O(y[246]),
    .I0(a[15]),
    .I1(b[6])
  );
  //OR U94bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U94bar (
    .O(ybar[246]),
    .I0(abar[15]),
    .I1(bbar[6])
  );
  //AND U95
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U95 (
    .O(y[245]),
    .I0(a[15]),
    .I1(b[5])
  );
  //OR U95bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U95bar (
    .O(ybar[245]),
    .I0(abar[15]),
    .I1(bbar[5])
  );
  //AND U96
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U96 (
    .O(y[244]),
    .I0(a[15]),
    .I1(b[4])
  );
  //OR U96bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U96bar (
    .O(ybar[244]),
    .I0(abar[15]),
    .I1(bbar[4])
  );
  //AND U97
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U97 (
    .O(y[243]),
    .I0(a[15]),
    .I1(b[3])
  );
  //OR U97bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U97bar (
    .O(ybar[243]),
    .I0(abar[15]),
    .I1(bbar[3])
  );
  //AND U98
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U98 (
    .O(y[242]),
    .I0(a[15]),
    .I1(b[2])
  );
  //OR U98bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U98bar (
    .O(ybar[242]),
    .I0(abar[15]),
    .I1(bbar[2])
  );
  //AND U99
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U99 (
    .O(y[241]),
    .I0(a[15]),
    .I1(b[1])
  );
  //OR U99bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U99bar (
    .O(ybar[241]),
    .I0(abar[15]),
    .I1(bbar[1])
  );
  //AND U100
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U100 (
    .O(y[240]),
    .I0(a[15]),
    .I1(b[0])
  );
  //OR U100bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U100bar (
    .O(ybar[240]),
    .I0(abar[15]),
    .I1(bbar[0])
  );
  //AND U101
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U101 (
    .O(y[23]),
    .I0(a[1]),
    .I1(b[7])
  );
  //OR U101bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U101bar (
    .O(ybar[23]),
    .I0(abar[1]),
    .I1(bbar[7])
  );
  //AND U102
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U102 (
    .O(y[239]),
    .I0(a[14]),
    .I1(b[15])
  );
  //OR U102bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U102bar (
    .O(ybar[239]),
    .I0(abar[14]),
    .I1(bbar[15])
  );
  //AND U103
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U103 (
    .O(y[238]),
    .I0(a[14]),
    .I1(b[14])
  );
  //OR U103bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U103bar (
    .O(ybar[238]),
    .I0(abar[14]),
    .I1(bbar[14])
  );
  //AND U104
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U104 (
    .O(y[237]),
    .I0(a[14]),
    .I1(b[13])
  );
  //OR U104bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U104bar (
    .O(ybar[237]),
    .I0(abar[14]),
    .I1(bbar[13])
  );
  //AND U105
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U105 (
    .O(y[236]),
    .I0(a[14]),
    .I1(b[12])
  );
  //OR U105bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U105bar (
    .O(ybar[236]),
    .I0(abar[14]),
    .I1(bbar[12])
  );
  //AND U106
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U106 (
    .O(y[235]),
    .I0(a[14]),
    .I1(b[11])
  );
  //OR U106bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U106bar (
    .O(ybar[235]),
    .I0(abar[14]),
    .I1(bbar[11])
  );
  //AND U107
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U107 (
    .O(y[234]),
    .I0(a[14]),
    .I1(b[10])
  );
  //OR U107bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U107bar (
    .O(ybar[234]),
    .I0(abar[14]),
    .I1(bbar[10])
  );
  //AND U108
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U108 (
    .O(y[233]),
    .I0(a[14]),
    .I1(b[9])
  );
  //OR U108bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U108bar (
    .O(ybar[233]),
    .I0(abar[14]),
    .I1(bbar[9])
  );
  //AND U109
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U109 (
    .O(y[232]),
    .I0(a[14]),
    .I1(b[8])
  );
  //OR U109bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U109bar (
    .O(ybar[232]),
    .I0(abar[14]),
    .I1(bbar[8])
  );
  //AND U110
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U110 (
    .O(y[231]),
    .I0(a[14]),
    .I1(b[7])
  );
  //OR U110bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U110bar (
    .O(ybar[231]),
    .I0(abar[14]),
    .I1(bbar[7])
  );
  //AND U111
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U111 (
    .O(y[230]),
    .I0(a[14]),
    .I1(b[6])
  );
  //OR U111bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U111bar (
    .O(ybar[230]),
    .I0(abar[14]),
    .I1(bbar[6])
  );
  //AND U112
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U112 (
    .O(y[22]),
    .I0(a[1]),
    .I1(b[6])
  );
  //OR U112bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U112bar (
    .O(ybar[22]),
    .I0(abar[1]),
    .I1(bbar[6])
  );
  //AND U113
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U113 (
    .O(y[229]),
    .I0(a[14]),
    .I1(b[5])
  );
  //OR U113bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U113bar (
    .O(ybar[229]),
    .I0(abar[14]),
    .I1(bbar[5])
  );
  //AND U114
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U114 (
    .O(y[228]),
    .I0(a[14]),
    .I1(b[4])
  );
  //OR U114bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U114bar (
    .O(ybar[228]),
    .I0(abar[14]),
    .I1(bbar[4])
  );
  //AND U115
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U115 (
    .O(y[227]),
    .I0(a[14]),
    .I1(b[3])
  );
  //OR U115bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U115bar (
    .O(ybar[227]),
    .I0(abar[14]),
    .I1(bbar[3])
  );
  //AND U116
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U116 (
    .O(y[226]),
    .I0(a[14]),
    .I1(b[2])
  );
  //OR U116bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U116bar (
    .O(ybar[226]),
    .I0(abar[14]),
    .I1(bbar[2])
  );
  //AND U117
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U117 (
    .O(y[225]),
    .I0(a[14]),
    .I1(b[1])
  );
  //OR U117bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U117bar (
    .O(ybar[225]),
    .I0(abar[14]),
    .I1(bbar[1])
  );
  //AND U118
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U118 (
    .O(y[224]),
    .I0(a[14]),
    .I1(b[0])
  );
  //OR U118bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U118bar (
    .O(ybar[224]),
    .I0(abar[14]),
    .I1(bbar[0])
  );
  //AND U119
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U119 (
    .O(y[223]),
    .I0(a[13]),
    .I1(b[15])
  );
  //OR U119bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U119bar (
    .O(ybar[223]),
    .I0(abar[13]),
    .I1(bbar[15])
  );
  //AND U120
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U120 (
    .O(y[222]),
    .I0(a[13]),
    .I1(b[14])
  );
  //OR U120bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U120bar (
    .O(ybar[222]),
    .I0(abar[13]),
    .I1(bbar[14])
  );
  //AND U121
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U121 (
    .O(y[221]),
    .I0(a[13]),
    .I1(b[13])
  );
  //OR U121bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U121bar (
    .O(ybar[221]),
    .I0(abar[13]),
    .I1(bbar[13])
  );
  //AND U122
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U122 (
    .O(y[220]),
    .I0(a[13]),
    .I1(b[12])
  );
  //OR U122bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U122bar (
    .O(ybar[220]),
    .I0(abar[13]),
    .I1(bbar[12])
  );
  //AND U123
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U123 (
    .O(y[21]),
    .I0(a[1]),
    .I1(b[5])
  );
  //OR U123bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U123bar (
    .O(ybar[21]),
    .I0(abar[1]),
    .I1(bbar[5])
  );
  //AND U124
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U124 (
    .O(y[219]),
    .I0(a[13]),
    .I1(b[11])
  );
  //OR U124bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U124bar (
    .O(ybar[219]),
    .I0(abar[13]),
    .I1(bbar[11])
  );
  //AND U125
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U125 (
    .O(y[218]),
    .I0(a[13]),
    .I1(b[10])
  );
  //OR U125bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U125bar (
    .O(ybar[218]),
    .I0(abar[13]),
    .I1(bbar[10])
  );
  //AND U126
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U126 (
    .O(y[217]),
    .I0(a[13]),
    .I1(b[9])
  );
  //OR U126bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U126bar (
    .O(ybar[217]),
    .I0(abar[13]),
    .I1(bbar[9])
  );
  //AND U127
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U127 (
    .O(y[216]),
    .I0(a[13]),
    .I1(b[8])
  );
  //OR U127bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U127bar (
    .O(ybar[216]),
    .I0(abar[13]),
    .I1(bbar[8])
  );
  //AND U128
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U128 (
    .O(y[215]),
    .I0(a[13]),
    .I1(b[7])
  );
  //OR U128bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U128bar (
    .O(ybar[215]),
    .I0(abar[13]),
    .I1(bbar[7])
  );
  //AND U129
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U129 (
    .O(y[214]),
    .I0(a[13]),
    .I1(b[6])
  );
  //OR U129bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U129bar (
    .O(ybar[214]),
    .I0(abar[13]),
    .I1(bbar[6])
  );
  //AND U130
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U130 (
    .O(y[213]),
    .I0(a[13]),
    .I1(b[5])
  );
  //OR U130bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U130bar (
    .O(ybar[213]),
    .I0(abar[13]),
    .I1(bbar[5])
  );
  //AND U131
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U131 (
    .O(y[212]),
    .I0(a[13]),
    .I1(b[4])
  );
  //OR U131bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U131bar (
    .O(ybar[212]),
    .I0(abar[13]),
    .I1(bbar[4])
  );
  //AND U132
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U132 (
    .O(y[211]),
    .I0(a[13]),
    .I1(b[3])
  );
  //OR U132bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U132bar (
    .O(ybar[211]),
    .I0(abar[13]),
    .I1(bbar[3])
  );
  //AND U133
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U133 (
    .O(y[210]),
    .I0(a[13]),
    .I1(b[2])
  );
  //OR U133bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U133bar (
    .O(ybar[210]),
    .I0(abar[13]),
    .I1(bbar[2])
  );
  //AND U134
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U134 (
    .O(y[20]),
    .I0(a[1]),
    .I1(b[4])
  );
  //OR U134bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U134bar (
    .O(ybar[20]),
    .I0(abar[1]),
    .I1(bbar[4])
  );
  //AND U135
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U135 (
    .O(y[209]),
    .I0(a[13]),
    .I1(b[1])
  );
  //OR U135bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U135bar (
    .O(ybar[209]),
    .I0(abar[13]),
    .I1(bbar[1])
  );
  //AND U136
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U136 (
    .O(y[208]),
    .I0(a[13]),
    .I1(b[0])
  );
  //OR U136bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U136bar (
    .O(ybar[208]),
    .I0(abar[13]),
    .I1(bbar[0])
  );
  //AND U137
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U137 (
    .O(y[207]),
    .I0(a[12]),
    .I1(b[15])
  );
  //OR U137bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U137bar (
    .O(ybar[207]),
    .I0(abar[12]),
    .I1(bbar[15])
  );
  //AND U138
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U138 (
    .O(y[206]),
    .I0(a[12]),
    .I1(b[14])
  );
  //OR U138bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U138bar (
    .O(ybar[206]),
    .I0(abar[12]),
    .I1(bbar[14])
  );
  //AND U139
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U139 (
    .O(y[205]),
    .I0(a[12]),
    .I1(b[13])
  );
  //OR U139bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U139bar (
    .O(ybar[205]),
    .I0(abar[12]),
    .I1(bbar[13])
  );
  //AND U140
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U140 (
    .O(y[204]),
    .I0(a[12]),
    .I1(b[12])
  );
  //OR U140bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U140bar (
    .O(ybar[204]),
    .I0(abar[12]),
    .I1(bbar[12])
  );
  //AND U141
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U141 (
    .O(y[203]),
    .I0(a[12]),
    .I1(b[11])
  );
  //OR U141bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U141bar (
    .O(ybar[203]),
    .I0(abar[12]),
    .I1(bbar[11])
  );
  //AND U142
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U142 (
    .O(y[202]),
    .I0(a[12]),
    .I1(b[10])
  );
  //OR U142bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U142bar (
    .O(ybar[202]),
    .I0(abar[12]),
    .I1(bbar[10])
  );
  //AND U143
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U143 (
    .O(y[201]),
    .I0(a[12]),
    .I1(b[9])
  );
  //OR U143bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U143bar (
    .O(ybar[201]),
    .I0(abar[12]),
    .I1(bbar[9])
  );
  //AND U144
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U144 (
    .O(y[200]),
    .I0(a[12]),
    .I1(b[8])
  );
  //OR U144bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U144bar (
    .O(ybar[200]),
    .I0(abar[12]),
    .I1(bbar[8])
  );
  //AND U145
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U145 (
    .O(y[1]),
    .I0(b[1]),
    .I1(a[0])
  );
  //OR U145bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U145bar (
    .O(ybar[1]),
    .I0(bbar[1]),
    .I1(abar[0])
  );
  //AND U146
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U146 (
    .O(y[19]),
    .I0(a[1]),
    .I1(b[3])
  );
  //OR U146bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U146bar (
    .O(ybar[19]),
    .I0(abar[1]),
    .I1(bbar[3])
  );
  //AND U147
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U147 (
    .O(y[199]),
    .I0(a[12]),
    .I1(b[7])
  );
  //OR U147bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U147bar (
    .O(ybar[199]),
    .I0(abar[12]),
    .I1(bbar[7])
  );
  //AND U148
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U148 (
    .O(y[198]),
    .I0(a[12]),
    .I1(b[6])
  );
  //OR U148bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U148bar (
    .O(ybar[198]),
    .I0(abar[12]),
    .I1(bbar[6])
  );
  //AND U149
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U149 (
    .O(y[197]),
    .I0(a[12]),
    .I1(b[5])
  );
  //OR U149bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U149bar (
    .O(ybar[197]),
    .I0(abar[12]),
    .I1(bbar[5])
  );
  //AND U150
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U150 (
    .O(y[196]),
    .I0(a[12]),
    .I1(b[4])
  );
  //OR U150bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U150bar (
    .O(ybar[196]),
    .I0(abar[12]),
    .I1(bbar[4])
  );
  //AND U151
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U151 (
    .O(y[195]),
    .I0(a[12]),
    .I1(b[3])
  );
  //OR U151bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U151bar (
    .O(ybar[195]),
    .I0(abar[12]),
    .I1(bbar[3])
  );
  //AND U152
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U152 (
    .O(y[194]),
    .I0(a[12]),
    .I1(b[2])
  );
  //OR U152bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U152bar (
    .O(ybar[194]),
    .I0(abar[12]),
    .I1(bbar[2])
  );
  //AND U153
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U153 (
    .O(y[193]),
    .I0(a[12]),
    .I1(b[1])
  );
  //OR U153bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U153bar (
    .O(ybar[193]),
    .I0(abar[12]),
    .I1(bbar[1])
  );
  //AND U154
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U154 (
    .O(y[192]),
    .I0(a[12]),
    .I1(b[0])
  );
  //OR U154bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U154bar (
    .O(ybar[192]),
    .I0(abar[12]),
    .I1(bbar[0])
  );
  //AND U155
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U155 (
    .O(y[191]),
    .I0(a[11]),
    .I1(b[15])
  );
  //OR U155bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U155bar (
    .O(ybar[191]),
    .I0(abar[11]),
    .I1(bbar[15])
  );
  //AND U156
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U156 (
    .O(y[190]),
    .I0(a[11]),
    .I1(b[14])
  );
  //OR U156bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U156bar (
    .O(ybar[190]),
    .I0(abar[11]),
    .I1(bbar[14])
  );
  //AND U157
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U157 (
    .O(y[18]),
    .I0(a[1]),
    .I1(b[2])
  );
  //OR U157bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U157bar (
    .O(ybar[18]),
    .I0(abar[1]),
    .I1(bbar[2])
  );
  //AND U158
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U158 (
    .O(y[189]),
    .I0(a[11]),
    .I1(b[13])
  );
  //OR U158bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U158bar (
    .O(ybar[189]),
    .I0(abar[11]),
    .I1(bbar[13])
  );
  //AND U159
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U159 (
    .O(y[188]),
    .I0(a[11]),
    .I1(b[12])
  );
  //OR U159bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U159bar (
    .O(ybar[188]),
    .I0(abar[11]),
    .I1(bbar[12])
  );
  //AND U160
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U160 (
    .O(y[187]),
    .I0(a[11]),
    .I1(b[11])
  );
  //OR U160bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U160bar (
    .O(ybar[187]),
    .I0(abar[11]),
    .I1(bbar[11])
  );
  //AND U161
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U161 (
    .O(y[186]),
    .I0(a[11]),
    .I1(b[10])
  );
  //OR U161bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U161bar (
    .O(ybar[186]),
    .I0(abar[11]),
    .I1(bbar[10])
  );
  //AND U162
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U162 (
    .O(y[185]),
    .I0(a[11]),
    .I1(b[9])
  );
  //OR U162bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U162bar (
    .O(ybar[185]),
    .I0(abar[11]),
    .I1(bbar[9])
  );
  //AND U163
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U163 (
    .O(y[184]),
    .I0(a[11]),
    .I1(b[8])
  );
  //OR U163bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U163bar (
    .O(ybar[184]),
    .I0(abar[11]),
    .I1(bbar[8])
  );
  //AND U164
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U164 (
    .O(y[183]),
    .I0(a[11]),
    .I1(b[7])
  );
  //OR U164bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U164bar (
    .O(ybar[183]),
    .I0(abar[11]),
    .I1(bbar[7])
  );
  //AND U165
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U165 (
    .O(y[182]),
    .I0(a[11]),
    .I1(b[6])
  );
  //OR U165bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U165bar (
    .O(ybar[182]),
    .I0(abar[11]),
    .I1(bbar[6])
  );
  //AND U166
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U166 (
    .O(y[181]),
    .I0(a[11]),
    .I1(b[5])
  );
  //OR U166bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U166bar (
    .O(ybar[181]),
    .I0(abar[11]),
    .I1(bbar[5])
  );
  //AND U167
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U167 (
    .O(y[180]),
    .I0(a[11]),
    .I1(b[4])
  );
  //OR U167bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U167bar (
    .O(ybar[180]),
    .I0(abar[11]),
    .I1(bbar[4])
  );
  //AND U168
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U168 (
    .O(y[17]),
    .I0(a[1]),
    .I1(b[1])
  );
  //OR U168bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U168bar (
    .O(ybar[17]),
    .I0(abar[1]),
    .I1(bbar[1])
  );
  //AND U169
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U169 (
    .O(y[179]),
    .I0(a[11]),
    .I1(b[3])
  );
  //OR U169bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U169bar (
    .O(ybar[179]),
    .I0(abar[11]),
    .I1(bbar[3])
  );
  //AND U170
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U170 (
    .O(y[178]),
    .I0(a[11]),
    .I1(b[2])
  );
  //OR U170bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U170bar (
    .O(ybar[178]),
    .I0(abar[11]),
    .I1(bbar[2])
  );
  //AND U171
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U171 (
    .O(y[177]),
    .I0(a[11]),
    .I1(b[1])
  );
  //OR U171bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U171bar (
    .O(ybar[177]),
    .I0(abar[11]),
    .I1(bbar[1])
  );
  //AND U172
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U172 (
    .O(y[176]),
    .I0(a[11]),
    .I1(b[0])
  );
  //OR U172bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U172bar (
    .O(ybar[176]),
    .I0(abar[11]),
    .I1(bbar[0])
  );
  //AND U173
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U173 (
    .O(y[175]),
    .I0(a[10]),
    .I1(b[15])
  );
  //OR U173bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U173bar (
    .O(ybar[175]),
    .I0(abar[10]),
    .I1(bbar[15])
  );
  //AND U174
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U174 (
    .O(y[174]),
    .I0(a[10]),
    .I1(b[14])
  );
  //OR U174bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U174bar (
    .O(ybar[174]),
    .I0(abar[10]),
    .I1(bbar[14])
  );
  //AND U175
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U175 (
    .O(y[173]),
    .I0(a[10]),
    .I1(b[13])
  );
  //OR U175bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U175bar (
    .O(ybar[173]),
    .I0(abar[10]),
    .I1(bbar[13])
  );
  //AND U176
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U176 (
    .O(y[172]),
    .I0(a[10]),
    .I1(b[12])
  );
  //OR U176bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U176bar (
    .O(ybar[172]),
    .I0(abar[10]),
    .I1(bbar[12])
  );
  //AND U177
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U177 (
    .O(y[171]),
    .I0(a[10]),
    .I1(b[11])
  );
  //OR U177bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U177bar (
    .O(ybar[171]),
    .I0(abar[10]),
    .I1(bbar[11])
  );
  //AND U178
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U178 (
    .O(y[170]),
    .I0(a[10]),
    .I1(b[10])
  );
  //OR U178bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U178bar (
    .O(ybar[170]),
    .I0(abar[10]),
    .I1(bbar[10])
  );
  //AND U179
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U179 (
    .O(y[16]),
    .I0(a[1]),
    .I1(b[0])
  );
  //OR U179bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U179bar (
    .O(ybar[16]),
    .I0(abar[1]),
    .I1(bbar[0])
  );
  //AND U180
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U180 (
    .O(y[169]),
    .I0(a[10]),
    .I1(b[9])
  );
  //OR U180bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U180bar (
    .O(ybar[169]),
    .I0(abar[10]),
    .I1(bbar[9])
  );
  //AND U181
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U181 (
    .O(y[168]),
    .I0(a[10]),
    .I1(b[8])
  );
  //OR U181bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U181bar (
    .O(ybar[168]),
    .I0(abar[10]),
    .I1(bbar[8])
  );
  //AND U182
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U182 (
    .O(y[167]),
    .I0(a[10]),
    .I1(b[7])
  );
  //OR U182bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U182bar (
    .O(ybar[167]),
    .I0(abar[10]),
    .I1(bbar[7])
  );
  //AND U183
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U183 (
    .O(y[166]),
    .I0(a[10]),
    .I1(b[6])
  );
  //OR U183bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U183bar (
    .O(ybar[166]),
    .I0(abar[10]),
    .I1(bbar[6])
  );
  //AND U184
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U184 (
    .O(y[165]),
    .I0(a[10]),
    .I1(b[5])
  );
  //OR U184bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U184bar (
    .O(ybar[165]),
    .I0(abar[10]),
    .I1(bbar[5])
  );
  //AND U185
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U185 (
    .O(y[164]),
    .I0(a[10]),
    .I1(b[4])
  );
  //OR U185bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U185bar (
    .O(ybar[164]),
    .I0(abar[10]),
    .I1(bbar[4])
  );
  //AND U186
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U186 (
    .O(y[163]),
    .I0(a[10]),
    .I1(b[3])
  );
  //OR U186bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U186bar (
    .O(ybar[163]),
    .I0(abar[10]),
    .I1(bbar[3])
  );
  //AND U187
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U187 (
    .O(y[162]),
    .I0(a[10]),
    .I1(b[2])
  );
  //OR U187bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U187bar (
    .O(ybar[162]),
    .I0(abar[10]),
    .I1(bbar[2])
  );
  //AND U188
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U188 (
    .O(y[161]),
    .I0(a[10]),
    .I1(b[1])
  );
  //OR U188bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U188bar (
    .O(ybar[161]),
    .I0(abar[10]),
    .I1(bbar[1])
  );
  //AND U189
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U189 (
    .O(y[160]),
    .I0(a[10]),
    .I1(b[0])
  );
  //OR U189bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U189bar (
    .O(ybar[160]),
    .I0(abar[10]),
    .I1(bbar[0])
  );
  //AND U190
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U190 (
    .O(y[15]),
    .I0(b[15]),
    .I1(a[0])
  );
  //OR U190bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U190bar (
    .O(ybar[15]),
    .I0(bbar[15]),
    .I1(abar[0])
  );
  //AND U191
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U191 (
    .O(y[159]),
    .I0(a[9]),
    .I1(b[15])
  );
  //OR U191bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U191bar (
    .O(ybar[159]),
    .I0(abar[9]),
    .I1(bbar[15])
  );
  //AND U192
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U192 (
    .O(y[158]),
    .I0(a[9]),
    .I1(b[14])
  );
  //OR U192bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U192bar (
    .O(ybar[158]),
    .I0(abar[9]),
    .I1(bbar[14])
  );
  //AND U193
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U193 (
    .O(y[157]),
    .I0(a[9]),
    .I1(b[13])
  );
  //OR U193bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U193bar (
    .O(ybar[157]),
    .I0(abar[9]),
    .I1(bbar[13])
  );
  //AND U194
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U194 (
    .O(y[156]),
    .I0(a[9]),
    .I1(b[12])
  );
  //OR U194bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U194bar (
    .O(ybar[156]),
    .I0(abar[9]),
    .I1(bbar[12])
  );
  //AND U195
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U195 (
    .O(y[155]),
    .I0(a[9]),
    .I1(b[11])
  );
  //OR U195bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U195bar (
    .O(ybar[155]),
    .I0(abar[9]),
    .I1(bbar[11])
  );
  //AND U196
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U196 (
    .O(y[154]),
    .I0(a[9]),
    .I1(b[10])
  );
  //OR U196bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U196bar (
    .O(ybar[154]),
    .I0(abar[9]),
    .I1(bbar[10])
  );
  //AND U197
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U197 (
    .O(y[153]),
    .I0(a[9]),
    .I1(b[9])
  );
  //OR U197bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U197bar (
    .O(ybar[153]),
    .I0(abar[9]),
    .I1(bbar[9])
  );
  //AND U198
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U198 (
    .O(y[152]),
    .I0(a[9]),
    .I1(b[8])
  );
  //OR U198bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U198bar (
    .O(ybar[152]),
    .I0(abar[9]),
    .I1(bbar[8])
  );
  //AND U199
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U199 (
    .O(y[151]),
    .I0(a[9]),
    .I1(b[7])
  );
  //OR U199bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U199bar (
    .O(ybar[151]),
    .I0(abar[9]),
    .I1(bbar[7])
  );
  //AND U200
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U200 (
    .O(y[150]),
    .I0(a[9]),
    .I1(b[6])
  );
  //OR U200bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U200bar (
    .O(ybar[150]),
    .I0(abar[9]),
    .I1(bbar[6])
  );
  //AND U201
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U201 (
    .O(y[14]),
    .I0(b[14]),
    .I1(a[0])
  );
  //OR U201bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U201bar (
    .O(ybar[14]),
    .I0(bbar[14]),
    .I1(abar[0])
  );
  //AND U202
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U202 (
    .O(y[149]),
    .I0(a[9]),
    .I1(b[5])
  );
  //OR U202bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U202bar (
    .O(ybar[149]),
    .I0(abar[9]),
    .I1(bbar[5])
  );
  //AND U203
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U203 (
    .O(y[148]),
    .I0(a[9]),
    .I1(b[4])
  );
  //OR U203bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U203bar (
    .O(ybar[148]),
    .I0(abar[9]),
    .I1(bbar[4])
  );
  //AND U204
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U204 (
    .O(y[147]),
    .I0(a[9]),
    .I1(b[3])
  );
  //OR U204bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U204bar (
    .O(ybar[147]),
    .I0(abar[9]),
    .I1(bbar[3])
  );
  //AND U205
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U205 (
    .O(y[146]),
    .I0(a[9]),
    .I1(b[2])
  );
  //OR U205bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U205bar (
    .O(ybar[146]),
    .I0(abar[9]),
    .I1(bbar[2])
  );
  //AND U206
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U206 (
    .O(y[145]),
    .I0(a[9]),
    .I1(b[1])
  );
  //OR U206bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U206bar (
    .O(ybar[145]),
    .I0(abar[9]),
    .I1(bbar[1])
  );
  //AND U207
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U207 (
    .O(y[144]),
    .I0(a[9]),
    .I1(b[0])
  );
  //OR U207bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U207bar (
    .O(ybar[144]),
    .I0(abar[9]),
    .I1(bbar[0])
  );
  //AND U208
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U208 (
    .O(y[143]),
    .I0(a[8]),
    .I1(b[15])
  );
  //OR U208bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U208bar (
    .O(ybar[143]),
    .I0(abar[8]),
    .I1(bbar[15])
  );
  //AND U209
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U209 (
    .O(y[142]),
    .I0(a[8]),
    .I1(b[14])
  );
  //OR U209bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U209bar (
    .O(ybar[142]),
    .I0(abar[8]),
    .I1(bbar[14])
  );
  //AND U210
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U210 (
    .O(y[141]),
    .I0(a[8]),
    .I1(b[13])
  );
  //OR U210bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U210bar (
    .O(ybar[141]),
    .I0(abar[8]),
    .I1(bbar[13])
  );
  //AND U211
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U211 (
    .O(y[140]),
    .I0(a[8]),
    .I1(b[12])
  );
  //OR U211bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U211bar (
    .O(ybar[140]),
    .I0(abar[8]),
    .I1(bbar[12])
  );
  //AND U212
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U212 (
    .O(y[13]),
    .I0(b[13]),
    .I1(a[0])
  );
  //OR U212bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U212bar (
    .O(ybar[13]),
    .I0(bbar[13]),
    .I1(abar[0])
  );
  //AND U213
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U213 (
    .O(y[139]),
    .I0(a[8]),
    .I1(b[11])
  );
  //OR U213bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U213bar (
    .O(ybar[139]),
    .I0(abar[8]),
    .I1(bbar[11])
  );
  //AND U214
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U214 (
    .O(y[138]),
    .I0(a[8]),
    .I1(b[10])
  );
  //OR U214bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U214bar (
    .O(ybar[138]),
    .I0(abar[8]),
    .I1(bbar[10])
  );
  //AND U215
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U215 (
    .O(y[137]),
    .I0(a[8]),
    .I1(b[9])
  );
  //OR U215bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U215bar (
    .O(ybar[137]),
    .I0(abar[8]),
    .I1(bbar[9])
  );
  //AND U216
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U216 (
    .O(y[136]),
    .I0(a[8]),
    .I1(b[8])
  );
  //OR U216bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U216bar (
    .O(ybar[136]),
    .I0(abar[8]),
    .I1(bbar[8])
  );
  //AND U217
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U217 (
    .O(y[135]),
    .I0(a[8]),
    .I1(b[7])
  );
  //OR U217bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U217bar (
    .O(ybar[135]),
    .I0(abar[8]),
    .I1(bbar[7])
  );
  //AND U218
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U218 (
    .O(y[134]),
    .I0(a[8]),
    .I1(b[6])
  );
  //OR U218bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U218bar (
    .O(ybar[134]),
    .I0(abar[8]),
    .I1(bbar[6])
  );
  //AND U219
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U219 (
    .O(y[133]),
    .I0(a[8]),
    .I1(b[5])
  );
  //OR U219bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U219bar (
    .O(ybar[133]),
    .I0(abar[8]),
    .I1(bbar[5])
  );
  //AND U220
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U220 (
    .O(y[132]),
    .I0(a[8]),
    .I1(b[4])
  );
  //OR U220bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U220bar (
    .O(ybar[132]),
    .I0(abar[8]),
    .I1(bbar[4])
  );
  //AND U221
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U221 (
    .O(y[131]),
    .I0(a[8]),
    .I1(b[3])
  );
  //OR U221bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U221bar (
    .O(ybar[131]),
    .I0(abar[8]),
    .I1(bbar[3])
  );
  //AND U222
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U222 (
    .O(y[130]),
    .I0(a[8]),
    .I1(b[2])
  );
  //OR U222bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U222bar (
    .O(ybar[130]),
    .I0(abar[8]),
    .I1(bbar[2])
  );
  //AND U223
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U223 (
    .O(y[12]),
    .I0(b[12]),
    .I1(a[0])
  );
  //OR U223bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U223bar (
    .O(ybar[12]),
    .I0(bbar[12]),
    .I1(abar[0])
  );
  //AND U224
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U224 (
    .O(y[129]),
    .I0(a[8]),
    .I1(b[1])
  );
  //OR U224bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U224bar (
    .O(ybar[129]),
    .I0(abar[8]),
    .I1(bbar[1])
  );
  //AND U225
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U225 (
    .O(y[128]),
    .I0(a[8]),
    .I1(b[0])
  );
  //OR U225bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U225bar (
    .O(ybar[128]),
    .I0(abar[8]),
    .I1(bbar[0])
  );
  //AND U226
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U226 (
    .O(y[127]),
    .I0(a[7]),
    .I1(b[15])
  );
  //OR U226bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U226bar (
    .O(ybar[127]),
    .I0(abar[7]),
    .I1(bbar[15])
  );
  //AND U227
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U227 (
    .O(y[126]),
    .I0(a[7]),
    .I1(b[14])
  );
  //OR U227bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U227bar (
    .O(ybar[126]),
    .I0(abar[7]),
    .I1(bbar[14])
  );
  //AND U228
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U228 (
    .O(y[125]),
    .I0(a[7]),
    .I1(b[13])
  );
  //OR U228bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U228bar (
    .O(ybar[125]),
    .I0(abar[7]),
    .I1(bbar[13])
  );
  //AND U229
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U229 (
    .O(y[124]),
    .I0(a[7]),
    .I1(b[12])
  );
  //OR U229bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U229bar (
    .O(ybar[124]),
    .I0(abar[7]),
    .I1(bbar[12])
  );
  //AND U230
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U230 (
    .O(y[123]),
    .I0(a[7]),
    .I1(b[11])
  );
  //OR U230bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U230bar (
    .O(ybar[123]),
    .I0(abar[7]),
    .I1(bbar[11])
  );
  //AND U231
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U231 (
    .O(y[122]),
    .I0(a[7]),
    .I1(b[10])
  );
  //OR U231bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U231bar (
    .O(ybar[122]),
    .I0(abar[7]),
    .I1(bbar[10])
  );
  //AND U232
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U232 (
    .O(y[121]),
    .I0(a[7]),
    .I1(b[9])
  );
  //OR U232bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U232bar (
    .O(ybar[121]),
    .I0(abar[7]),
    .I1(bbar[9])
  );
  //AND U233
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U233 (
    .O(y[120]),
    .I0(a[7]),
    .I1(b[8])
  );
  //OR U233bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U233bar (
    .O(ybar[120]),
    .I0(abar[7]),
    .I1(bbar[8])
  );
  //AND U234
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U234 (
    .O(y[11]),
    .I0(b[11]),
    .I1(a[0])
  );
  //OR U234bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U234bar (
    .O(ybar[11]),
    .I0(bbar[11]),
    .I1(abar[0])
  );
  //AND U235
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U235 (
    .O(y[119]),
    .I0(a[7]),
    .I1(b[7])
  );
  //OR U235bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U235bar (
    .O(ybar[119]),
    .I0(abar[7]),
    .I1(bbar[7])
  );
  //AND U236
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U236 (
    .O(y[118]),
    .I0(a[7]),
    .I1(b[6])
  );
  //OR U236bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U236bar (
    .O(ybar[118]),
    .I0(abar[7]),
    .I1(bbar[6])
  );
  //AND U237
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U237 (
    .O(y[117]),
    .I0(a[7]),
    .I1(b[5])
  );
  //OR U237bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U237bar (
    .O(ybar[117]),
    .I0(abar[7]),
    .I1(bbar[5])
  );
  //AND U238
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U238 (
    .O(y[116]),
    .I0(a[7]),
    .I1(b[4])
  );
  //OR U238bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U238bar (
    .O(ybar[116]),
    .I0(abar[7]),
    .I1(bbar[4])
  );
  //AND U239
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U239 (
    .O(y[115]),
    .I0(a[7]),
    .I1(b[3])
  );
  //OR U239bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U239bar (
    .O(ybar[115]),
    .I0(abar[7]),
    .I1(bbar[3])
  );
  //AND U240
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U240 (
    .O(y[114]),
    .I0(a[7]),
    .I1(b[2])
  );
  //OR U240bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U240bar (
    .O(ybar[114]),
    .I0(abar[7]),
    .I1(bbar[2])
  );
  //AND U241
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U241 (
    .O(y[113]),
    .I0(a[7]),
    .I1(b[1])
  );
  //OR U241bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U241bar (
    .O(ybar[113]),
    .I0(abar[7]),
    .I1(bbar[1])
  );
  //AND U242
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U242 (
    .O(y[112]),
    .I0(a[7]),
    .I1(b[0])
  );
  //OR U242bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U242bar (
    .O(ybar[112]),
    .I0(abar[7]),
    .I1(bbar[0])
  );
  //AND U243
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U243 (
    .O(y[111]),
    .I0(b[15]),
    .I1(a[6])
  );
  //OR U243bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U243bar (
    .O(ybar[111]),
    .I0(bbar[15]),
    .I1(abar[6])
  );
  //AND U244
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U244 (
    .O(y[110]),
    .I0(b[14]),
    .I1(a[6])
  );
  //OR U244bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U244bar (
    .O(ybar[110]),
    .I0(bbar[14]),
    .I1(abar[6])
  );
  //AND U245
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U245 (
    .O(y[10]),
    .I0(b[10]),
    .I1(a[0])
  );
  //OR U245bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U245bar (
    .O(ybar[10]),
    .I0(bbar[10]),
    .I1(abar[0])
  );
  //AND U246
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U246 (
    .O(y[109]),
    .I0(b[13]),
    .I1(a[6])
  );
  //OR U246bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U246bar (
    .O(ybar[109]),
    .I0(bbar[13]),
    .I1(abar[6])
  );
  //AND U247
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U247 (
    .O(y[108]),
    .I0(b[12]),
    .I1(a[6])
  );
  //OR U247bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U247bar (
    .O(ybar[108]),
    .I0(bbar[12]),
    .I1(abar[6])
  );
  //AND U248
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U248 (
    .O(y[107]),
    .I0(b[11]),
    .I1(a[6])
  );
  //OR U248bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U248bar (
    .O(ybar[107]),
    .I0(bbar[11]),
    .I1(abar[6])
  );
  //AND U249
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U249 (
    .O(y[106]),
    .I0(b[10]),
    .I1(a[6])
  );
  //OR U249bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U249bar (
    .O(ybar[106]),
    .I0(bbar[10]),
    .I1(abar[6])
  );
  //AND U250
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U250 (
    .O(y[105]),
    .I0(a[6]),
    .I1(b[9])
  );
  //OR U250bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U250bar (
    .O(ybar[105]),
    .I0(abar[6]),
    .I1(bbar[9])
  );
  //AND U251
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U251 (
    .O(y[104]),
    .I0(b[8]),
    .I1(a[6])
  );
  //OR U251bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U251bar (
    .O(ybar[104]),
    .I0(bbar[8]),
    .I1(abar[6])
  );
  //AND U252
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U252 (
    .O(y[103]),
    .I0(b[7]),
    .I1(a[6])
  );
  //OR U252bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U252bar (
    .O(ybar[103]),
    .I0(bbar[7]),
    .I1(abar[6])
  );
  //AND U253
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U253 (
    .O(y[102]),
    .I0(b[6]),
    .I1(a[6])
  );
  //OR U253bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U253bar (
    .O(ybar[102]),
    .I0(bbar[6]),
    .I1(abar[6])
  );
  //AND U254
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U254 (
    .O(y[101]),
    .I0(b[5]),
    .I1(a[6])
  );
  //OR U254bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U254bar (
    .O(ybar[101]),
    .I0(bbar[5]),
    .I1(abar[6])
  );
  //AND U255
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U255 (
    .O(y[100]),
    .I0(b[4]),
    .I1(a[6])
  );
  //OR U255bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U255bar (
    .O(ybar[100]),
    .I0(bbar[4]),
    .I1(abar[6])
  );
  //AND U256
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U256 (
    .O(y[0]),
    .I0(b[0]),
    .I1(a[0])
  );
  //OR U256bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U256bar (
    .O(ybar[0]),
    .I0(bbar[0]),
    .I1(abar[0])
  );
endmodule

module decode_7 ( in, out );

  input wire [7:0] in;
//input_done

  output wire [255:0] out;
//output_done

  wire [15:0] level1;
  wire [31:0] level2;
//wire_done

  CD2_28 cd_l1_1 ( .a(in[1]), .b(in[0]), .y(level1[3:0]) );
  CD2_27 cd_l1_2 ( .a(in[3]), .b(in[2]), .y(level1[7:4]) );
  CD2_26 cd_l1_3 ( .a(in[5]), .b(in[4]), .y(level1[11:8]) );
  CD2_25 cd_l1_4 ( .a(in[7]), .b(in[6]), .y(level1[15:12]) );
  CD4_14 cd_l2_1 ( .a(level1[7:4]), .b(level1[3:0]), .y(level2[15:0]) );
  CD4_13 cd_l2_2 ( .a(level1[15:12]), .b(level1[11:8]), .y(level2[31:16]) );
  CD16_7 cd_l3 ( .a(level2[31:16]), .b(level2[15:0]), .y(out) );
endmodule

module encode_7 ( in, out );

  input wire [255:0] in;
  wire [255:0] inbar;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
  assign inbar[8] = ~in[8];
  assign inbar[9] = ~in[9];
  assign inbar[10] = ~in[10];
  assign inbar[11] = ~in[11];
  assign inbar[12] = ~in[12];
  assign inbar[13] = ~in[13];
  assign inbar[14] = ~in[14];
  assign inbar[15] = ~in[15];
  assign inbar[16] = ~in[16];
  assign inbar[17] = ~in[17];
  assign inbar[18] = ~in[18];
  assign inbar[19] = ~in[19];
  assign inbar[20] = ~in[20];
  assign inbar[21] = ~in[21];
  assign inbar[22] = ~in[22];
  assign inbar[23] = ~in[23];
  assign inbar[24] = ~in[24];
  assign inbar[25] = ~in[25];
  assign inbar[26] = ~in[26];
  assign inbar[27] = ~in[27];
  assign inbar[28] = ~in[28];
  assign inbar[29] = ~in[29];
  assign inbar[30] = ~in[30];
  assign inbar[31] = ~in[31];
  assign inbar[32] = ~in[32];
  assign inbar[33] = ~in[33];
  assign inbar[34] = ~in[34];
  assign inbar[35] = ~in[35];
  assign inbar[36] = ~in[36];
  assign inbar[37] = ~in[37];
  assign inbar[38] = ~in[38];
  assign inbar[39] = ~in[39];
  assign inbar[40] = ~in[40];
  assign inbar[41] = ~in[41];
  assign inbar[42] = ~in[42];
  assign inbar[43] = ~in[43];
  assign inbar[44] = ~in[44];
  assign inbar[45] = ~in[45];
  assign inbar[46] = ~in[46];
  assign inbar[47] = ~in[47];
  assign inbar[48] = ~in[48];
  assign inbar[49] = ~in[49];
  assign inbar[50] = ~in[50];
  assign inbar[51] = ~in[51];
  assign inbar[52] = ~in[52];
  assign inbar[53] = ~in[53];
  assign inbar[54] = ~in[54];
  assign inbar[55] = ~in[55];
  assign inbar[56] = ~in[56];
  assign inbar[57] = ~in[57];
  assign inbar[58] = ~in[58];
  assign inbar[59] = ~in[59];
  assign inbar[60] = ~in[60];
  assign inbar[61] = ~in[61];
  assign inbar[62] = ~in[62];
  assign inbar[63] = ~in[63];
  assign inbar[64] = ~in[64];
  assign inbar[65] = ~in[65];
  assign inbar[66] = ~in[66];
  assign inbar[67] = ~in[67];
  assign inbar[68] = ~in[68];
  assign inbar[69] = ~in[69];
  assign inbar[70] = ~in[70];
  assign inbar[71] = ~in[71];
  assign inbar[72] = ~in[72];
  assign inbar[73] = ~in[73];
  assign inbar[74] = ~in[74];
  assign inbar[75] = ~in[75];
  assign inbar[76] = ~in[76];
  assign inbar[77] = ~in[77];
  assign inbar[78] = ~in[78];
  assign inbar[79] = ~in[79];
  assign inbar[80] = ~in[80];
  assign inbar[81] = ~in[81];
  assign inbar[82] = ~in[82];
  assign inbar[83] = ~in[83];
  assign inbar[84] = ~in[84];
  assign inbar[85] = ~in[85];
  assign inbar[86] = ~in[86];
  assign inbar[87] = ~in[87];
  assign inbar[88] = ~in[88];
  assign inbar[89] = ~in[89];
  assign inbar[90] = ~in[90];
  assign inbar[91] = ~in[91];
  assign inbar[92] = ~in[92];
  assign inbar[93] = ~in[93];
  assign inbar[94] = ~in[94];
  assign inbar[95] = ~in[95];
  assign inbar[96] = ~in[96];
  assign inbar[97] = ~in[97];
  assign inbar[98] = ~in[98];
  assign inbar[99] = ~in[99];
  assign inbar[100] = ~in[100];
  assign inbar[101] = ~in[101];
  assign inbar[102] = ~in[102];
  assign inbar[103] = ~in[103];
  assign inbar[104] = ~in[104];
  assign inbar[105] = ~in[105];
  assign inbar[106] = ~in[106];
  assign inbar[107] = ~in[107];
  assign inbar[108] = ~in[108];
  assign inbar[109] = ~in[109];
  assign inbar[110] = ~in[110];
  assign inbar[111] = ~in[111];
  assign inbar[112] = ~in[112];
  assign inbar[113] = ~in[113];
  assign inbar[114] = ~in[114];
  assign inbar[115] = ~in[115];
  assign inbar[116] = ~in[116];
  assign inbar[117] = ~in[117];
  assign inbar[118] = ~in[118];
  assign inbar[119] = ~in[119];
  assign inbar[120] = ~in[120];
  assign inbar[121] = ~in[121];
  assign inbar[122] = ~in[122];
  assign inbar[123] = ~in[123];
  assign inbar[124] = ~in[124];
  assign inbar[125] = ~in[125];
  assign inbar[126] = ~in[126];
  assign inbar[127] = ~in[127];
  assign inbar[128] = ~in[128];
  assign inbar[129] = ~in[129];
  assign inbar[130] = ~in[130];
  assign inbar[131] = ~in[131];
  assign inbar[132] = ~in[132];
  assign inbar[133] = ~in[133];
  assign inbar[134] = ~in[134];
  assign inbar[135] = ~in[135];
  assign inbar[136] = ~in[136];
  assign inbar[137] = ~in[137];
  assign inbar[138] = ~in[138];
  assign inbar[139] = ~in[139];
  assign inbar[140] = ~in[140];
  assign inbar[141] = ~in[141];
  assign inbar[142] = ~in[142];
  assign inbar[143] = ~in[143];
  assign inbar[144] = ~in[144];
  assign inbar[145] = ~in[145];
  assign inbar[146] = ~in[146];
  assign inbar[147] = ~in[147];
  assign inbar[148] = ~in[148];
  assign inbar[149] = ~in[149];
  assign inbar[150] = ~in[150];
  assign inbar[151] = ~in[151];
  assign inbar[152] = ~in[152];
  assign inbar[153] = ~in[153];
  assign inbar[154] = ~in[154];
  assign inbar[155] = ~in[155];
  assign inbar[156] = ~in[156];
  assign inbar[157] = ~in[157];
  assign inbar[158] = ~in[158];
  assign inbar[159] = ~in[159];
  assign inbar[160] = ~in[160];
  assign inbar[161] = ~in[161];
  assign inbar[162] = ~in[162];
  assign inbar[163] = ~in[163];
  assign inbar[164] = ~in[164];
  assign inbar[165] = ~in[165];
  assign inbar[166] = ~in[166];
  assign inbar[167] = ~in[167];
  assign inbar[168] = ~in[168];
  assign inbar[169] = ~in[169];
  assign inbar[170] = ~in[170];
  assign inbar[171] = ~in[171];
  assign inbar[172] = ~in[172];
  assign inbar[173] = ~in[173];
  assign inbar[174] = ~in[174];
  assign inbar[175] = ~in[175];
  assign inbar[176] = ~in[176];
  assign inbar[177] = ~in[177];
  assign inbar[178] = ~in[178];
  assign inbar[179] = ~in[179];
  assign inbar[180] = ~in[180];
  assign inbar[181] = ~in[181];
  assign inbar[182] = ~in[182];
  assign inbar[183] = ~in[183];
  assign inbar[184] = ~in[184];
  assign inbar[185] = ~in[185];
  assign inbar[186] = ~in[186];
  assign inbar[187] = ~in[187];
  assign inbar[188] = ~in[188];
  assign inbar[189] = ~in[189];
  assign inbar[190] = ~in[190];
  assign inbar[191] = ~in[191];
  assign inbar[192] = ~in[192];
  assign inbar[193] = ~in[193];
  assign inbar[194] = ~in[194];
  assign inbar[195] = ~in[195];
  assign inbar[196] = ~in[196];
  assign inbar[197] = ~in[197];
  assign inbar[198] = ~in[198];
  assign inbar[199] = ~in[199];
  assign inbar[200] = ~in[200];
  assign inbar[201] = ~in[201];
  assign inbar[202] = ~in[202];
  assign inbar[203] = ~in[203];
  assign inbar[204] = ~in[204];
  assign inbar[205] = ~in[205];
  assign inbar[206] = ~in[206];
  assign inbar[207] = ~in[207];
  assign inbar[208] = ~in[208];
  assign inbar[209] = ~in[209];
  assign inbar[210] = ~in[210];
  assign inbar[211] = ~in[211];
  assign inbar[212] = ~in[212];
  assign inbar[213] = ~in[213];
  assign inbar[214] = ~in[214];
  assign inbar[215] = ~in[215];
  assign inbar[216] = ~in[216];
  assign inbar[217] = ~in[217];
  assign inbar[218] = ~in[218];
  assign inbar[219] = ~in[219];
  assign inbar[220] = ~in[220];
  assign inbar[221] = ~in[221];
  assign inbar[222] = ~in[222];
  assign inbar[223] = ~in[223];
  assign inbar[224] = ~in[224];
  assign inbar[225] = ~in[225];
  assign inbar[226] = ~in[226];
  assign inbar[227] = ~in[227];
  assign inbar[228] = ~in[228];
  assign inbar[229] = ~in[229];
  assign inbar[230] = ~in[230];
  assign inbar[231] = ~in[231];
  assign inbar[232] = ~in[232];
  assign inbar[233] = ~in[233];
  assign inbar[234] = ~in[234];
  assign inbar[235] = ~in[235];
  assign inbar[236] = ~in[236];
  assign inbar[237] = ~in[237];
  assign inbar[238] = ~in[238];
  assign inbar[239] = ~in[239];
  assign inbar[240] = ~in[240];
  assign inbar[241] = ~in[241];
  assign inbar[242] = ~in[242];
  assign inbar[243] = ~in[243];
  assign inbar[244] = ~in[244];
  assign inbar[245] = ~in[245];
  assign inbar[246] = ~in[246];
  assign inbar[247] = ~in[247];
  assign inbar[248] = ~in[248];
  assign inbar[249] = ~in[249];
  assign inbar[250] = ~in[250];
  assign inbar[251] = ~in[251];
  assign inbar[252] = ~in[252];
  assign inbar[253] = ~in[253];
  assign inbar[254] = ~in[254];
  assign inbar[255] = ~in[255];
//input_done

  output wire [7:0] out;
  wire [7:0] outbar;
//output_done

  wire in_81;
  wire in_80;
  wire in_79;
  wire in_78;
  wire in_77;
  wire in_76;
  wire in_75;
  wire in_74;
  wire in_73;
  wire in_72;
  wire in_71;
  wire in_70;
  wire in_69;
  wire in_68;
  wire in_67;
  wire in_66;
  wire in_65;
  wire in_64;
  wire in_63;
  wire in_62;
  wire in_61;
  wire in_60;
  wire in_59;
  wire in_58;
  wire in_57;
  wire in_56;
  wire in_55;
  wire in_54;
  wire in_53;
  wire in_52;
  wire in_51;
  wire in_50;
  wire in_49;
  wire in_48;
  wire in_47;
  wire in_46;
  wire in_45;
  wire in_44;
  wire in_43;
  wire in_42;
  wire in_41;
  wire in_40;
  wire in_39;
  wire in_38;
  wire in_37;
  wire in_36;
  wire in_35;
  wire in_34;
  wire in_33;
  wire in_32;
  wire in_31;
  wire in_30;
  wire in_29;
  wire in_28;
  wire in_27;
  wire in_26;
  wire in_25;
  wire in_24;
  wire in_23;
  wire in_22;
  wire in_21;
  wire in_20;
  wire in_19;
  wire in_18;
  wire in_17;
  wire in_16;
  wire in_15;
  wire in_14;
  wire in_13;
  wire in_12;
  wire in_11;
  wire in_10;
  wire in_9;
  wire in_8;
  wire in_7;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_3;
  wire in_2;
  wire in_1;
  wire in_0;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire in_81bar;
  wire in_80bar;
  wire in_79bar;
  wire in_78bar;
  wire in_77bar;
  wire in_76bar;
  wire in_75bar;
  wire in_74bar;
  wire in_73bar;
  wire in_72bar;
  wire in_71bar;
  wire in_70bar;
  wire in_69bar;
  wire in_68bar;
  wire in_67bar;
  wire in_66bar;
  wire in_65bar;
  wire in_64bar;
  wire in_63bar;
  wire in_62bar;
  wire in_61bar;
  wire in_60bar;
  wire in_59bar;
  wire in_58bar;
  wire in_57bar;
  wire in_56bar;
  wire in_55bar;
  wire in_54bar;
  wire in_53bar;
  wire in_52bar;
  wire in_51bar;
  wire in_50bar;
  wire in_49bar;
  wire in_48bar;
  wire in_47bar;
  wire in_46bar;
  wire in_45bar;
  wire in_44bar;
  wire in_43bar;
  wire in_42bar;
  wire in_41bar;
  wire in_40bar;
  wire in_39bar;
  wire in_38bar;
  wire in_37bar;
  wire in_36bar;
  wire in_35bar;
  wire in_34bar;
  wire in_33bar;
  wire in_32bar;
  wire in_31bar;
  wire in_30bar;
  wire in_29bar;
  wire in_28bar;
  wire in_27bar;
  wire in_26bar;
  wire in_25bar;
  wire in_24bar;
  wire in_23bar;
  wire in_22bar;
  wire in_21bar;
  wire in_20bar;
  wire in_19bar;
  wire in_18bar;
  wire in_17bar;
  wire in_16bar;
  wire in_15bar;
  wire in_14bar;
  wire in_13bar;
  wire in_12bar;
  wire in_11bar;
  wire in_10bar;
  wire in_9bar;
  wire in_8bar;
  wire in_7bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_3bar;
  wire in_2bar;
  wire in_1bar;
  wire in_0bar;
  wire n487bar;
  wire n488bar;
  wire n489bar;
  wire n490bar;
  wire n491bar;
  wire n492bar;
  wire n493bar;
  wire n494bar;
  wire n495bar;
  wire n496bar;
  wire n497bar;
  wire n498bar;
  wire n499bar;
  wire n500bar;
  wire n501bar;
  wire n502bar;
  wire n503bar;
  wire n504bar;
  wire n505bar;
  wire n506bar;
  wire n507bar;
  wire n508bar;
  wire n509bar;
  wire n510bar;
  wire n511bar;
  wire n512bar;
  wire n513bar;
  wire n514bar;
  wire n515bar;
  wire n516bar;
  wire n517bar;
  wire n518bar;
  wire n519bar;
  wire n520bar;
  wire n521bar;
  wire n522bar;
  wire n523bar;
  wire n524bar;
  wire n525bar;
  wire n526bar;
  wire n527bar;
  wire n528bar;
  wire n529bar;
  wire n530bar;
  wire n531bar;
  wire n532bar;
  wire n533bar;
  wire n534bar;
  wire n535bar;
  wire n536bar;
  wire n537bar;
  wire n538bar;
  wire n539bar;
  wire n540bar;
  wire n541bar;
  wire n542bar;
  wire n543bar;
  wire n544bar;
  wire n545bar;
  wire n546bar;
  wire n547bar;
  wire n548bar;
  wire n549bar;
  wire n550bar;
  wire n551bar;
  wire n552bar;
  wire n553bar;
  wire n554bar;
  wire n555bar;
  wire n556bar;
  wire n557bar;
  wire n558bar;
  wire n559bar;
  wire n560bar;
  wire n561bar;
  wire n562bar;
  wire n563bar;
  wire n564bar;
  wire n565bar;
  wire n566bar;
  wire n567bar;
  wire n568bar;
  wire n569bar;
  wire n570bar;
  wire n571bar;
  wire n572bar;
  wire n573bar;
  wire n574bar;
  wire n575bar;
  wire n576bar;
  wire n577bar;
  wire n578bar;
  wire n579bar;
  wire n580bar;
  wire n581bar;
  wire n582bar;
  wire n583bar;
  wire n584bar;
  wire n585bar;
  wire n586bar;
  wire n587bar;
  wire n588bar;
  wire n589bar;
  wire n590bar;
  wire n591bar;
  wire n592bar;
  wire n593bar;
  wire n594bar;
  wire n595bar;
  wire n596bar;
  wire n597bar;
  wire n598bar;
  wire n599bar;
  wire n600bar;
  wire n601bar;
  wire n602bar;
  wire n603bar;
  wire n604bar;
  wire n605bar;
  wire n606bar;
  wire n607bar;
  wire n608bar;
  wire n609bar;
  wire n610bar;
  wire n611bar;
  wire n612bar;
  wire n613bar;
  wire n614bar;
  wire n615bar;
  wire n616bar;
  wire n617bar;
  wire n618bar;
  wire n619bar;
  wire n620bar;
  wire n621bar;
  wire n622bar;
  wire n623bar;
  wire n624bar;
  wire n625bar;
  wire n626bar;
  wire n627bar;
  wire n628bar;
  wire n629bar;
  wire n630bar;
  wire n631bar;
  wire n632bar;
  wire n633bar;
  wire n634bar;
  wire n635bar;
  wire n636bar;
  wire n637bar;
  wire n638bar;
  wire n639bar;
  wire n640bar;
  wire n641bar;
  wire n642bar;
  wire n643bar;
  wire n644bar;
  wire n645bar;
  wire n646bar;
  wire n647bar;
  wire n648bar;
  wire n649bar;
  wire n650bar;
  wire n651bar;
  wire n652bar;
  wire n653bar;
  wire n654bar;
  wire n655bar;
  wire n656bar;
  wire n657bar;
  wire n658bar;
  wire n659bar;
  wire n660bar;
  wire n661bar;
  wire n662bar;
  wire n663bar;
  wire n664bar;
  wire n665bar;
  wire n666bar;
  wire n667bar;
  wire n668bar;
  wire n669bar;
  wire n670bar;
  wire n671bar;
  wire n672bar;
  wire n673bar;
  wire n674bar;
  wire n675bar;
  wire n676bar;
  wire n677bar;
  wire n678bar;
  wire n679bar;
  wire n680bar;
  wire n681bar;
  wire n682bar;
  wire n683bar;
  wire n684bar;
  wire n685bar;
  wire n686bar;
  wire n687bar;
  wire n688bar;
  wire n689bar;
  wire n690bar;
  wire n691bar;
  wire n692bar;
  wire n693bar;
  wire n694bar;
  wire n695bar;
  wire n696bar;
  wire n697bar;
  wire n698bar;
  wire n699bar;
  wire n700bar;
  wire n701bar;
  wire n702bar;
  wire n703bar;
  wire n704bar;
  wire n705bar;
  wire n706bar;
  wire n707bar;
  wire n708bar;
  wire n709bar;
  wire n710bar;
  wire n711bar;
  wire n712bar;
  wire n713bar;
  wire n714bar;
  wire n715bar;
  wire n716bar;
  wire n717bar;
  wire n718bar;
  wire n719bar;
  wire n720bar;
  wire n721bar;
  wire n722bar;
  wire n723bar;
  wire n724bar;
  wire n725bar;
  wire n726bar;
  wire n727bar;
  wire n728bar;
  wire n729bar;
  wire n730bar;
  wire n731bar;
  wire n732bar;
  wire n733bar;
  wire n734bar;
  wire n735bar;
  wire n736bar;
  wire n737bar;
  wire n738bar;
  wire n739bar;
  wire n740bar;
  wire n741bar;
  wire n742bar;
  wire n743bar;
  wire n744bar;
  wire n745bar;
  wire n746bar;
  wire n747bar;
  wire n748bar;
  wire n749bar;
  wire n750bar;
  wire n751bar;
  wire n752bar;
  wire n753bar;
  wire n754bar;
  wire n755bar;
  wire n756bar;
  wire n757bar;
  wire n758bar;
  wire n759bar;
  wire n760bar;
  wire n761bar;
  wire n762bar;
  wire n763bar;
  wire n764bar;
  wire n765bar;
  wire n766bar;
  wire n767bar;
  wire n768bar;
  wire n769bar;
  wire n770bar;
  wire n771bar;
  wire n772bar;
  wire n773bar;
  wire n774bar;
  wire n775bar;
  wire n776bar;
  wire n777bar;
  wire n778bar;
  wire n779bar;
  wire n780bar;
  wire n781bar;
  wire n782bar;
  wire n783bar;
  wire n784bar;
  wire n785bar;
  wire n786bar;
  wire n787bar;
  wire n788bar;
  wire n789bar;
  wire n790bar;
  wire n791bar;
  wire n792bar;
  wire n793bar;
  wire n794bar;
  wire n795bar;
  wire n796bar;
  wire n797bar;
  wire n798bar;
  wire n799bar;
  wire n800bar;
  wire n801bar;
  wire n802bar;
  wire n803bar;
  wire n804bar;
  wire n805bar;
  wire n806bar;
  wire n807bar;
  wire n808bar;
  wire n809bar;
  wire n810bar;
  wire n811bar;
  wire n812bar;
  wire n813bar;
  wire n814bar;
  wire n815bar;
  wire n816bar;
  wire n817bar;
  wire n818bar;
  wire n819bar;
  wire n820bar;
  wire n821bar;
  wire n822bar;
  wire n823bar;
  wire n824bar;
  wire n825bar;
  wire n826bar;
  wire n827bar;
  wire n828bar;
  wire n829bar;
  wire n830bar;
  wire n831bar;
  wire n832bar;
  wire n833bar;
  wire n834bar;
  wire n835bar;
  wire n836bar;
  wire n837bar;
  wire n838bar;
  wire n839bar;
  wire n840bar;
  wire n841bar;
  wire n842bar;
  wire n843bar;
  wire n844bar;
  wire n845bar;
  wire n846bar;
  wire n847bar;
  wire n848bar;
  wire n849bar;
  wire n850bar;
  wire n851bar;
  wire n852bar;
  wire n853bar;
  wire n854bar;
  wire n855bar;
  wire n856bar;
  wire n857bar;
  wire n858bar;
  wire n859bar;
  wire n860bar;
  wire n861bar;
  wire n862bar;
  wire n863bar;
  wire n864bar;
  wire n865bar;
  wire n866bar;
  wire n867bar;
  wire n868bar;
  wire n869bar;
  wire n870bar;
  wire n871bar;
  wire n872bar;
  wire n873bar;
  wire n874bar;
  wire n875bar;
  wire n876bar;
  wire n877bar;
  wire n878bar;
  wire n879bar;
  wire n880bar;
  wire n881bar;
  wire n882bar;
  wire n883bar;
  wire n884bar;
  wire n885bar;
  wire n886bar;
  wire n887bar;
  wire n888bar;
  wire n889bar;
  wire n890bar;
  wire n891bar;
  wire n892bar;
  wire n893bar;
  wire n894bar;
  wire n895bar;
  wire n896bar;
  wire n897bar;
  wire n898bar;
  wire n899bar;
  wire n900bar;
  wire n901bar;
  wire n902bar;
  wire n903bar;
  wire n904bar;
  wire n905bar;
  wire n906bar;
  wire n907bar;
  wire n908bar;
  wire n909bar;
  wire n910bar;
  wire n911bar;
  wire n912bar;
  wire n913bar;
  wire n914bar;
  wire n915bar;
  wire n916bar;
  wire n917bar;
  wire n918bar;
  wire n919bar;
  wire n920bar;
  wire n921bar;
  wire n922bar;
  wire n923bar;
  wire n924bar;
  wire n925bar;
  wire n926bar;
  wire n927bar;
  wire n928bar;
  wire n929bar;
  wire n930bar;
  wire n931bar;
  wire n932bar;
  wire n933bar;
  wire n934bar;
  wire n935bar;
  wire n936bar;
  wire n937bar;
  wire n938bar;
  wire n939bar;
  wire n940bar;
  wire n941bar;
  wire n942bar;
  wire n943bar;
  wire n944bar;
  wire n945bar;
  wire n946bar;
  wire n947bar;
  wire n948bar;
  wire n949bar;
  wire n950bar;
  wire n951bar;
  wire n952bar;
  wire n953bar;
  wire n954bar;
  wire n955bar;
  wire n956bar;
  wire n957bar;
  wire n958bar;
  wire n959bar;
  wire n960bar;
  wire n961bar;
  wire n962bar;
  wire n963bar;
  wire n964bar;
  wire n965bar;
  wire n966bar;
  wire n967bar;
  wire n968bar;
  wire n969bar;
  wire n970bar;
  wire n971bar;
  wire n972bar;
//wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];
  //OR U1
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1 (
    .O(out[7]),
    .I0(n972),
    .I1(n971)
  );
  //AND U1bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1bar (
    .O(outbar[7]),
    .I0(n972bar),
    .I1(n971bar)
  );
  //OR U2
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2 (
    .O(n971),
    .I0(n970),
    .I1(n969)
  );
  //AND U2bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2bar (
    .O(n971bar),
    .I0(n970bar),
    .I1(n969bar)
  );
  //OR U3
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3 (
    .O(n969),
    .I0(n968),
    .I1(n967)
  );
  //AND U3bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3bar (
    .O(n969bar),
    .I0(n968bar),
    .I1(n967bar)
  );
  //OR U4
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4 (
    .O(n967),
    .I0(n966),
    .I1(n965)
  );
  //AND U4bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4bar (
    .O(n967bar),
    .I0(n966bar),
    .I1(n965bar)
  );
  //OR U5
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5 (
    .O(n968),
    .I0(n964),
    .I1(n963)
  );
  //AND U5bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5bar (
    .O(n968bar),
    .I0(n964bar),
    .I1(n963bar)
  );
  //OR U6
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6 (
    .O(n963),
    .I0(in[116]),
    .I1(n962)
  );
  //AND U6bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6bar (
    .O(n963bar),
    .I0(inbar[116]),
    .I1(n962bar)
  );
  //OR U7
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7 (
    .O(n970),
    .I0(n961),
    .I1(n960)
  );
  //AND U7bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7bar (
    .O(n970bar),
    .I0(n961bar),
    .I1(n960bar)
  );
  //OR U8
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8 (
    .O(n960),
    .I0(in[150]),
    .I1(in[127])
  );
  //AND U8bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8bar (
    .O(n960bar),
    .I0(inbar[150]),
    .I1(inbar[127])
  );
  //OR U9
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9 (
    .O(n961),
    .I0(in[160]),
    .I1(n959)
  );
  //AND U9bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9bar (
    .O(n961bar),
    .I0(inbar[160]),
    .I1(n959bar)
  );
  //OR U10
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10 (
    .O(n959),
    .I0(in[252]),
    .I1(in[168])
  );
  //AND U10bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10bar (
    .O(n959bar),
    .I0(inbar[252]),
    .I1(inbar[168])
  );
  //OR U11
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11 (
    .O(n972),
    .I0(n958),
    .I1(n957)
  );
  //AND U11bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11bar (
    .O(n972bar),
    .I0(n958bar),
    .I1(n957bar)
  );
  //OR U12
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12 (
    .O(n957),
    .I0(n956),
    .I1(n955)
  );
  //AND U12bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12bar (
    .O(n957bar),
    .I0(n956bar),
    .I1(n955bar)
  );
  //OR U13
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13 (
    .O(n955),
    .I0(in_17),
    .I1(in[96])
  );
  //AND U13bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13bar (
    .O(n955bar),
    .I0(in_17bar),
    .I1(inbar[96])
  );
  //OR U14
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14 (
    .O(n956),
    .I0(in_23),
    .I1(n954)
  );
  //AND U14bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14bar (
    .O(n956bar),
    .I0(in_23bar),
    .I1(n954bar)
  );
  //OR U15
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15 (
    .O(n954),
    .I0(in_31),
    .I1(in_26)
  );
  //AND U15bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15bar (
    .O(n954bar),
    .I0(in_31bar),
    .I1(in_26bar)
  );
  //OR U16
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16 (
    .O(n958),
    .I0(n953),
    .I1(n952)
  );
  //AND U16bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16bar (
    .O(n958bar),
    .I0(n953bar),
    .I1(n952bar)
  );
  //OR U17
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U17 (
    .O(n952),
    .I0(in_58),
    .I1(in_4)
  );
  //AND U17bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U17bar (
    .O(n952bar),
    .I0(in_58bar),
    .I1(in_4bar)
  );
  //OR U18
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U18 (
    .O(n953),
    .I0(in_59),
    .I1(n951)
  );
  //AND U18bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U18bar (
    .O(n953bar),
    .I0(in_59bar),
    .I1(n951bar)
  );
  //OR U19
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U19 (
    .O(n951),
    .I0(in_71),
    .I1(in_62)
  );
  //AND U19bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U19bar (
    .O(n951bar),
    .I0(in_71bar),
    .I1(in_62bar)
  );
  //OR U20
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U20 (
    .O(out[6]),
    .I0(n950),
    .I1(n949)
  );
  //AND U20bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U20bar (
    .O(outbar[6]),
    .I0(n950bar),
    .I1(n949bar)
  );
  //OR U21
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U21 (
    .O(n949),
    .I0(n948),
    .I1(n947)
  );
  //AND U21bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U21bar (
    .O(n949bar),
    .I0(n948bar),
    .I1(n947bar)
  );
  //OR U22
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U22 (
    .O(n947),
    .I0(n946),
    .I1(n945)
  );
  //AND U22bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U22bar (
    .O(n947bar),
    .I0(n946bar),
    .I1(n945bar)
  );
  //OR U23
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U23 (
    .O(n945),
    .I0(n944),
    .I1(n943)
  );
  //AND U23bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U23bar (
    .O(n945bar),
    .I0(n944bar),
    .I1(n943bar)
  );
  //OR U24
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U24 (
    .O(n946),
    .I0(n942),
    .I1(n941)
  );
  //AND U24bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U24bar (
    .O(n946bar),
    .I0(n942bar),
    .I1(n941bar)
  );
  //OR U25
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U25 (
    .O(n941),
    .I0(in[101]),
    .I1(n940)
  );
  //AND U25bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U25bar (
    .O(n941bar),
    .I0(inbar[101]),
    .I1(n940bar)
  );
  //OR U26
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U26 (
    .O(n948),
    .I0(n939),
    .I1(n938)
  );
  //AND U26bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U26bar (
    .O(n948bar),
    .I0(n939bar),
    .I1(n938bar)
  );
  //OR U27
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U27 (
    .O(n938),
    .I0(in[114]),
    .I1(in[104])
  );
  //AND U27bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U27bar (
    .O(n938bar),
    .I0(inbar[114]),
    .I1(inbar[104])
  );
  //OR U28
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U28 (
    .O(n939),
    .I0(in[128]),
    .I1(n937)
  );
  //AND U28bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U28bar (
    .O(n939bar),
    .I0(inbar[128]),
    .I1(n937bar)
  );
  //OR U29
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U29 (
    .O(n937),
    .I0(in[136]),
    .I1(in[134])
  );
  //AND U29bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U29bar (
    .O(n937bar),
    .I0(inbar[136]),
    .I1(inbar[134])
  );
  //OR U30
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U30 (
    .O(n950),
    .I0(n936),
    .I1(n935)
  );
  //AND U30bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U30bar (
    .O(n950bar),
    .I0(n936bar),
    .I1(n935bar)
  );
  //OR U31
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U31 (
    .O(n935),
    .I0(n934),
    .I1(n933)
  );
  //AND U31bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U31bar (
    .O(n935bar),
    .I0(n934bar),
    .I1(n933bar)
  );
  //OR U32
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U32 (
    .O(n933),
    .I0(in[177]),
    .I1(in[164])
  );
  //AND U32bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U32bar (
    .O(n933bar),
    .I0(inbar[177]),
    .I1(inbar[164])
  );
  //OR U33
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U33 (
    .O(n934),
    .I0(in[212]),
    .I1(n932)
  );
  //AND U33bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U33bar (
    .O(n934bar),
    .I0(inbar[212]),
    .I1(n932bar)
  );
  //OR U34
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U34 (
    .O(n932),
    .I0(in[248]),
    .I1(in[221])
  );
  //AND U34bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U34bar (
    .O(n932bar),
    .I0(inbar[248]),
    .I1(inbar[221])
  );
  //OR U35
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U35 (
    .O(n936),
    .I0(n931),
    .I1(n930)
  );
  //AND U35bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U35bar (
    .O(n936bar),
    .I0(n931bar),
    .I1(n930bar)
  );
  //OR U36
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U36 (
    .O(n930),
    .I0(in_18),
    .I1(in[93])
  );
  //AND U36bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U36bar (
    .O(n930bar),
    .I0(in_18bar),
    .I1(inbar[93])
  );
  //OR U37
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U37 (
    .O(n931),
    .I0(in_31),
    .I1(n929)
  );
  //AND U37bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U37bar (
    .O(n931bar),
    .I0(in_31bar),
    .I1(n929bar)
  );
  //OR U38
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U38 (
    .O(n929),
    .I0(in_7),
    .I1(in_39)
  );
  //AND U38bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U38bar (
    .O(n929bar),
    .I0(in_7bar),
    .I1(in_39bar)
  );
  //OR U39
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U39 (
    .O(out[5]),
    .I0(n928),
    .I1(n927)
  );
  //AND U39bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U39bar (
    .O(outbar[5]),
    .I0(n928bar),
    .I1(n927bar)
  );
  //OR U40
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U40 (
    .O(n927),
    .I0(n926),
    .I1(n925)
  );
  //AND U40bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U40bar (
    .O(n927bar),
    .I0(n926bar),
    .I1(n925bar)
  );
  //OR U41
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U41 (
    .O(n925),
    .I0(n924),
    .I1(n923)
  );
  //AND U41bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U41bar (
    .O(n925bar),
    .I0(n924bar),
    .I1(n923bar)
  );
  //OR U42
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U42 (
    .O(n923),
    .I0(n922),
    .I1(n921)
  );
  //AND U42bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U42bar (
    .O(n923bar),
    .I0(n922bar),
    .I1(n921bar)
  );
  //OR U43
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U43 (
    .O(n924),
    .I0(n940),
    .I1(n920)
  );
  //AND U43bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U43bar (
    .O(n924bar),
    .I0(n940bar),
    .I1(n920bar)
  );
  //OR U44
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U44 (
    .O(n920),
    .I0(in[111]),
    .I1(n919)
  );
  //AND U44bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U44bar (
    .O(n920bar),
    .I0(inbar[111]),
    .I1(n919bar)
  );
  //OR U45
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U45 (
    .O(n940),
    .I0(n918),
    .I1(n917)
  );
  //AND U45bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U45bar (
    .O(n940bar),
    .I0(n918bar),
    .I1(n917bar)
  );
  //OR U46
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U46 (
    .O(n917),
    .I0(n916),
    .I1(n915)
  );
  //AND U46bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U46bar (
    .O(n917bar),
    .I0(n916bar),
    .I1(n915bar)
  );
  //OR U47
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U47 (
    .O(n915),
    .I0(n914),
    .I1(n913)
  );
  //AND U47bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U47bar (
    .O(n915bar),
    .I0(n914bar),
    .I1(n913bar)
  );
  //OR U48
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U48 (
    .O(n913),
    .I0(in[140]),
    .I1(in[131])
  );
  //AND U48bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U48bar (
    .O(n913bar),
    .I0(inbar[140]),
    .I1(inbar[131])
  );
  //OR U49
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U49 (
    .O(n914),
    .I0(in[160]),
    .I1(in[144])
  );
  //AND U49bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U49bar (
    .O(n914bar),
    .I0(inbar[160]),
    .I1(inbar[144])
  );
  //OR U50
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U50 (
    .O(n916),
    .I0(n912),
    .I1(n911)
  );
  //AND U50bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U50bar (
    .O(n916bar),
    .I0(n912bar),
    .I1(n911bar)
  );
  //OR U51
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U51 (
    .O(n911),
    .I0(in[179]),
    .I1(in[174])
  );
  //AND U51bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U51bar (
    .O(n911bar),
    .I0(inbar[179]),
    .I1(inbar[174])
  );
  //OR U52
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U52 (
    .O(n912),
    .I0(in[188]),
    .I1(in[184])
  );
  //AND U52bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U52bar (
    .O(n912bar),
    .I0(inbar[188]),
    .I1(inbar[184])
  );
  //OR U53
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U53 (
    .O(n918),
    .I0(n910),
    .I1(n909)
  );
  //AND U53bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U53bar (
    .O(n918bar),
    .I0(n910bar),
    .I1(n909bar)
  );
  //OR U54
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U54 (
    .O(n909),
    .I0(n908),
    .I1(n907)
  );
  //AND U54bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U54bar (
    .O(n909bar),
    .I0(n908bar),
    .I1(n907bar)
  );
  //OR U55
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U55 (
    .O(n907),
    .I0(in[216]),
    .I1(in[200])
  );
  //AND U55bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U55bar (
    .O(n907bar),
    .I0(inbar[216]),
    .I1(inbar[200])
  );
  //OR U56
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U56 (
    .O(n908),
    .I0(in[228]),
    .I1(in[224])
  );
  //AND U56bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U56bar (
    .O(n908bar),
    .I0(inbar[228]),
    .I1(inbar[224])
  );
  //OR U57
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U57 (
    .O(n910),
    .I0(n906),
    .I1(n905)
  );
  //AND U57bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U57bar (
    .O(n910bar),
    .I0(n906bar),
    .I1(n905bar)
  );
  //OR U58
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U58 (
    .O(n905),
    .I0(in[247]),
    .I1(in[235])
  );
  //AND U58bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U58bar (
    .O(n905bar),
    .I0(inbar[247]),
    .I1(inbar[235])
  );
  //OR U59
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U59 (
    .O(n906),
    .I0(in_42),
    .I1(in[83])
  );
  //AND U59bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U59bar (
    .O(n906bar),
    .I0(in_42bar),
    .I1(inbar[83])
  );
  //OR U60
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U60 (
    .O(n926),
    .I0(n904),
    .I1(n903)
  );
  //AND U60bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U60bar (
    .O(n926bar),
    .I0(n904bar),
    .I1(n903bar)
  );
  //OR U61
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U61 (
    .O(n903),
    .I0(in[166]),
    .I1(in[123])
  );
  //AND U61bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U61bar (
    .O(n903bar),
    .I0(inbar[166]),
    .I1(inbar[123])
  );
  //OR U62
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U62 (
    .O(n904),
    .I0(in[170]),
    .I1(n902)
  );
  //AND U62bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U62bar (
    .O(n904bar),
    .I0(inbar[170]),
    .I1(n902bar)
  );
  //OR U63
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U63 (
    .O(n902),
    .I0(in[194]),
    .I1(in[183])
  );
  //AND U63bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U63bar (
    .O(n902bar),
    .I0(inbar[194]),
    .I1(inbar[183])
  );
  //OR U64
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U64 (
    .O(n928),
    .I0(n901),
    .I1(n900)
  );
  //AND U64bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U64bar (
    .O(n928bar),
    .I0(n901bar),
    .I1(n900bar)
  );
  //OR U65
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U65 (
    .O(n900),
    .I0(n899),
    .I1(n898)
  );
  //AND U65bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U65bar (
    .O(n900bar),
    .I0(n899bar),
    .I1(n898bar)
  );
  //OR U66
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U66 (
    .O(n898),
    .I0(in[241]),
    .I1(in[238])
  );
  //AND U66bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U66bar (
    .O(n898bar),
    .I0(inbar[241]),
    .I1(inbar[238])
  );
  //OR U67
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U67 (
    .O(n899),
    .I0(in[250]),
    .I1(n897)
  );
  //AND U67bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U67bar (
    .O(n899bar),
    .I0(inbar[250]),
    .I1(n897bar)
  );
  //OR U68
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U68 (
    .O(n897),
    .I0(in_24),
    .I1(in[84])
  );
  //AND U68bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U68bar (
    .O(n897bar),
    .I0(in_24bar),
    .I1(inbar[84])
  );
  //OR U69
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U69 (
    .O(n901),
    .I0(n896),
    .I1(n895)
  );
  //AND U69bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U69bar (
    .O(n901bar),
    .I0(n896bar),
    .I1(n895bar)
  );
  //OR U70
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U70 (
    .O(n895),
    .I0(in_41),
    .I1(in_29)
  );
  //AND U70bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U70bar (
    .O(n895bar),
    .I0(in_41bar),
    .I1(in_29bar)
  );
  //OR U71
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U71 (
    .O(n896),
    .I0(in_66),
    .I1(n894)
  );
  //AND U71bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U71bar (
    .O(n896bar),
    .I0(in_66bar),
    .I1(n894bar)
  );
  //OR U72
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U72 (
    .O(n894),
    .I0(in_76),
    .I1(in_71)
  );
  //AND U72bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U72bar (
    .O(n894bar),
    .I0(in_76bar),
    .I1(in_71bar)
  );
  //OR U73
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U73 (
    .O(out[4]),
    .I0(n893),
    .I1(n892)
  );
  //AND U73bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U73bar (
    .O(outbar[4]),
    .I0(n893bar),
    .I1(n892bar)
  );
  //OR U74
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U74 (
    .O(n892),
    .I0(n891),
    .I1(n890)
  );
  //AND U74bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U74bar (
    .O(n892bar),
    .I0(n891bar),
    .I1(n890bar)
  );
  //OR U75
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U75 (
    .O(n890),
    .I0(n889),
    .I1(n888)
  );
  //AND U75bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U75bar (
    .O(n890bar),
    .I0(n889bar),
    .I1(n888bar)
  );
  //OR U76
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U76 (
    .O(n888),
    .I0(n922),
    .I1(n887)
  );
  //AND U76bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U76bar (
    .O(n888bar),
    .I0(n922bar),
    .I1(n887bar)
  );
  //OR U77
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U77 (
    .O(n922),
    .I0(n886),
    .I1(n885)
  );
  //AND U77bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U77bar (
    .O(n922bar),
    .I0(n886bar),
    .I1(n885bar)
  );
  //OR U78
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U78 (
    .O(n885),
    .I0(n884),
    .I1(n883)
  );
  //AND U78bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U78bar (
    .O(n885bar),
    .I0(n884bar),
    .I1(n883bar)
  );
  //OR U79
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U79 (
    .O(n883),
    .I0(n882),
    .I1(n881)
  );
  //AND U79bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U79bar (
    .O(n883bar),
    .I0(n882bar),
    .I1(n881bar)
  );
  //OR U80
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U80 (
    .O(n881),
    .I0(in[118]),
    .I1(in[109])
  );
  //AND U80bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U80bar (
    .O(n881bar),
    .I0(inbar[118]),
    .I1(inbar[109])
  );
  //OR U81
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U81 (
    .O(n882),
    .I0(in[139]),
    .I1(in[120])
  );
  //AND U81bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U81bar (
    .O(n882bar),
    .I0(inbar[139]),
    .I1(inbar[120])
  );
  //OR U82
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U82 (
    .O(n884),
    .I0(n880),
    .I1(n879)
  );
  //AND U82bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U82bar (
    .O(n884bar),
    .I0(n880bar),
    .I1(n879bar)
  );
  //OR U83
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U83 (
    .O(n879),
    .I0(in[198]),
    .I1(in[154])
  );
  //AND U83bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U83bar (
    .O(n879bar),
    .I0(inbar[198]),
    .I1(inbar[154])
  );
  //OR U84
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U84 (
    .O(n880),
    .I0(in[210]),
    .I1(in[205])
  );
  //AND U84bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U84bar (
    .O(n880bar),
    .I0(inbar[210]),
    .I1(inbar[205])
  );
  //OR U85
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U85 (
    .O(n886),
    .I0(n878),
    .I1(n877)
  );
  //AND U85bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U85bar (
    .O(n886bar),
    .I0(n878bar),
    .I1(n877bar)
  );
  //OR U86
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U86 (
    .O(n877),
    .I0(n876),
    .I1(n875)
  );
  //AND U86bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U86bar (
    .O(n877bar),
    .I0(n876bar),
    .I1(n875bar)
  );
  //OR U87
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U87 (
    .O(n875),
    .I0(in[219]),
    .I1(in[217])
  );
  //AND U87bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U87bar (
    .O(n875bar),
    .I0(inbar[219]),
    .I1(inbar[217])
  );
  //OR U88
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U88 (
    .O(n876),
    .I0(in[86]),
    .I1(in[252])
  );
  //AND U88bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U88bar (
    .O(n876bar),
    .I0(inbar[86]),
    .I1(inbar[252])
  );
  //OR U89
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U89 (
    .O(n878),
    .I0(n874),
    .I1(n873)
  );
  //AND U89bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U89bar (
    .O(n878bar),
    .I0(n874bar),
    .I1(n873bar)
  );
  //OR U90
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U90 (
    .O(n873),
    .I0(in_40),
    .I1(in[91])
  );
  //AND U90bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U90bar (
    .O(n873bar),
    .I0(in_40bar),
    .I1(inbar[91])
  );
  //OR U91
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U91 (
    .O(n874),
    .I0(in_8),
    .I1(in_46)
  );
  //AND U91bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U91bar (
    .O(n874bar),
    .I0(in_8bar),
    .I1(in_46bar)
  );
  //OR U92
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U92 (
    .O(n889),
    .I0(n872),
    .I1(n871)
  );
  //AND U92bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U92bar (
    .O(n889bar),
    .I0(n872bar),
    .I1(n871bar)
  );
  //OR U93
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U93 (
    .O(n871),
    .I0(in[117]),
    .I1(n943)
  );
  //AND U93bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U93bar (
    .O(n871bar),
    .I0(inbar[117]),
    .I1(n943bar)
  );
  //OR U94
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U94 (
    .O(n943),
    .I0(n870),
    .I1(n869)
  );
  //AND U94bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U94bar (
    .O(n943bar),
    .I0(n870bar),
    .I1(n869bar)
  );
  //OR U95
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U95 (
    .O(n869),
    .I0(n868),
    .I1(n867)
  );
  //AND U95bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U95bar (
    .O(n869bar),
    .I0(n868bar),
    .I1(n867bar)
  );
  //OR U96
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U96 (
    .O(n867),
    .I0(n866),
    .I1(n865)
  );
  //AND U96bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U96bar (
    .O(n867bar),
    .I0(n866bar),
    .I1(n865bar)
  );
  //OR U97
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U97 (
    .O(n865),
    .I0(n864),
    .I1(n863)
  );
  //AND U97bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U97bar (
    .O(n865bar),
    .I0(n864bar),
    .I1(n863bar)
  );
  //OR U98
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U98 (
    .O(n866),
    .I0(in[108]),
    .I1(n919)
  );
  //AND U98bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U98bar (
    .O(n866bar),
    .I0(inbar[108]),
    .I1(n919bar)
  );
  //OR U99
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U99 (
    .O(n919),
    .I0(n862),
    .I1(n861)
  );
  //AND U99bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U99bar (
    .O(n919bar),
    .I0(n862bar),
    .I1(n861bar)
  );
  //OR U100
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U100 (
    .O(n861),
    .I0(n860),
    .I1(n859)
  );
  //AND U100bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U100bar (
    .O(n861bar),
    .I0(n860bar),
    .I1(n859bar)
  );
  //OR U101
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U101 (
    .O(n859),
    .I0(n858),
    .I1(n857)
  );
  //AND U101bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U101bar (
    .O(n859bar),
    .I0(n858bar),
    .I1(n857bar)
  );
  //OR U102
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U102 (
    .O(n857),
    .I0(in[119]),
    .I1(in[105])
  );
  //AND U102bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U102bar (
    .O(n857bar),
    .I0(inbar[119]),
    .I1(inbar[105])
  );
  //OR U103
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U103 (
    .O(n858),
    .I0(in[186]),
    .I1(in[175])
  );
  //AND U103bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U103bar (
    .O(n858bar),
    .I0(inbar[186]),
    .I1(inbar[175])
  );
  //OR U104
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U104 (
    .O(n860),
    .I0(n856),
    .I1(n855)
  );
  //AND U104bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U104bar (
    .O(n860bar),
    .I0(n856bar),
    .I1(n855bar)
  );
  //OR U105
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U105 (
    .O(n855),
    .I0(in[202]),
    .I1(in[193])
  );
  //AND U105bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U105bar (
    .O(n855bar),
    .I0(inbar[202]),
    .I1(inbar[193])
  );
  //OR U106
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U106 (
    .O(n856),
    .I0(in[225]),
    .I1(in[208])
  );
  //AND U106bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U106bar (
    .O(n856bar),
    .I0(inbar[225]),
    .I1(inbar[208])
  );
  //OR U107
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U107 (
    .O(n862),
    .I0(n854),
    .I1(n853)
  );
  //AND U107bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U107bar (
    .O(n862bar),
    .I0(n854bar),
    .I1(n853bar)
  );
  //OR U108
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U108 (
    .O(n853),
    .I0(n852),
    .I1(n851)
  );
  //AND U108bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U108bar (
    .O(n853bar),
    .I0(n852bar),
    .I1(n851bar)
  );
  //OR U109
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U109 (
    .O(n851),
    .I0(in_1),
    .I1(in[85])
  );
  //AND U109bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U109bar (
    .O(n851bar),
    .I0(in_1bar),
    .I1(inbar[85])
  );
  //OR U110
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U110 (
    .O(n852),
    .I0(in_23),
    .I1(in_19)
  );
  //AND U110bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U110bar (
    .O(n852bar),
    .I0(in_23bar),
    .I1(in_19bar)
  );
  //OR U111
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U111 (
    .O(n854),
    .I0(n850),
    .I1(n849)
  );
  //AND U111bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U111bar (
    .O(n854bar),
    .I0(n850bar),
    .I1(n849bar)
  );
  //OR U112
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U112 (
    .O(n849),
    .I0(in_43),
    .I1(in_33)
  );
  //AND U112bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U112bar (
    .O(n849bar),
    .I0(in_43bar),
    .I1(in_33bar)
  );
  //OR U113
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U113 (
    .O(n850),
    .I0(in_63),
    .I1(in_44)
  );
  //AND U113bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U113bar (
    .O(n850bar),
    .I0(in_63bar),
    .I1(in_44bar)
  );
  //OR U114
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U114 (
    .O(n868),
    .I0(n848),
    .I1(n847)
  );
  //AND U114bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U114bar (
    .O(n868bar),
    .I0(n848bar),
    .I1(n847bar)
  );
  //OR U115
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U115 (
    .O(n847),
    .I0(in[141]),
    .I1(in[112])
  );
  //AND U115bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U115bar (
    .O(n847bar),
    .I0(inbar[141]),
    .I1(inbar[112])
  );
  //OR U116
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U116 (
    .O(n848),
    .I0(in[147]),
    .I1(n846)
  );
  //AND U116bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U116bar (
    .O(n848bar),
    .I0(inbar[147]),
    .I1(n846bar)
  );
  //OR U117
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U117 (
    .O(n846),
    .I0(in[181]),
    .I1(in[167])
  );
  //AND U117bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U117bar (
    .O(n846bar),
    .I0(inbar[181]),
    .I1(inbar[167])
  );
  //OR U118
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U118 (
    .O(n870),
    .I0(n845),
    .I1(n844)
  );
  //AND U118bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U118bar (
    .O(n870bar),
    .I0(n845bar),
    .I1(n844bar)
  );
  //OR U119
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U119 (
    .O(n844),
    .I0(n843),
    .I1(n842)
  );
  //AND U119bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U119bar (
    .O(n844bar),
    .I0(n843bar),
    .I1(n842bar)
  );
  //OR U120
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U120 (
    .O(n842),
    .I0(in[229]),
    .I1(in[201])
  );
  //AND U120bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U120bar (
    .O(n842bar),
    .I0(inbar[229]),
    .I1(inbar[201])
  );
  //OR U121
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U121 (
    .O(n843),
    .I0(in[237]),
    .I1(n841)
  );
  //AND U121bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U121bar (
    .O(n843bar),
    .I0(inbar[237]),
    .I1(n841bar)
  );
  //OR U122
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U122 (
    .O(n841),
    .I0(in[94]),
    .I1(in[253])
  );
  //AND U122bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U122bar (
    .O(n841bar),
    .I0(inbar[94]),
    .I1(inbar[253])
  );
  //OR U123
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U123 (
    .O(n845),
    .I0(n840),
    .I1(n839)
  );
  //AND U123bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U123bar (
    .O(n845bar),
    .I0(n840bar),
    .I1(n839bar)
  );
  //OR U124
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U124 (
    .O(n839),
    .I0(in_21),
    .I1(in[96])
  );
  //AND U124bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U124bar (
    .O(n839bar),
    .I0(in_21bar),
    .I1(inbar[96])
  );
  //OR U125
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U125 (
    .O(n840),
    .I0(in_25),
    .I1(n838)
  );
  //AND U125bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U125bar (
    .O(n840bar),
    .I0(in_25bar),
    .I1(n838bar)
  );
  //OR U126
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U126 (
    .O(n838),
    .I0(in_81),
    .I1(in_45)
  );
  //AND U126bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U126bar (
    .O(n838bar),
    .I0(in_81bar),
    .I1(in_45bar)
  );
  //OR U127
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U127 (
    .O(n891),
    .I0(n837),
    .I1(n836)
  );
  //AND U127bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U127bar (
    .O(n891bar),
    .I0(n837bar),
    .I1(n836bar)
  );
  //OR U128
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U128 (
    .O(n836),
    .I0(in[142]),
    .I1(in[124])
  );
  //AND U128bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U128bar (
    .O(n836bar),
    .I0(inbar[142]),
    .I1(inbar[124])
  );
  //OR U129
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U129 (
    .O(n837),
    .I0(in[150]),
    .I1(n835)
  );
  //AND U129bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U129bar (
    .O(n837bar),
    .I0(inbar[150]),
    .I1(n835bar)
  );
  //OR U130
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U130 (
    .O(n835),
    .I0(in[172]),
    .I1(in[155])
  );
  //AND U130bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U130bar (
    .O(n835bar),
    .I0(inbar[172]),
    .I1(inbar[155])
  );
  //OR U131
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U131 (
    .O(n893),
    .I0(n834),
    .I1(n833)
  );
  //AND U131bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U131bar (
    .O(n893bar),
    .I0(n834bar),
    .I1(n833bar)
  );
  //OR U132
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U132 (
    .O(n833),
    .I0(n832),
    .I1(n831)
  );
  //AND U132bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U132bar (
    .O(n833bar),
    .I0(n832bar),
    .I1(n831bar)
  );
  //OR U133
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U133 (
    .O(n831),
    .I0(in[196]),
    .I1(in[173])
  );
  //AND U133bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U133bar (
    .O(n831bar),
    .I0(inbar[196]),
    .I1(inbar[173])
  );
  //OR U134
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U134 (
    .O(n832),
    .I0(in[222]),
    .I1(n830)
  );
  //AND U134bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U134bar (
    .O(n832bar),
    .I0(inbar[222]),
    .I1(n830bar)
  );
  //OR U135
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U135 (
    .O(n830),
    .I0(in[227]),
    .I1(in[226])
  );
  //AND U135bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U135bar (
    .O(n830bar),
    .I0(inbar[227]),
    .I1(inbar[226])
  );
  //OR U136
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U136 (
    .O(n834),
    .I0(n829),
    .I1(n828)
  );
  //AND U136bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U136bar (
    .O(n834bar),
    .I0(n829bar),
    .I1(n828bar)
  );
  //OR U137
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U137 (
    .O(n828),
    .I0(in[249]),
    .I1(in[231])
  );
  //AND U137bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U137bar (
    .O(n828bar),
    .I0(inbar[249]),
    .I1(inbar[231])
  );
  //OR U138
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U138 (
    .O(n829),
    .I0(in_28),
    .I1(n827)
  );
  //AND U138bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U138bar (
    .O(n829bar),
    .I0(in_28bar),
    .I1(n827bar)
  );
  //OR U139
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U139 (
    .O(n827),
    .I0(in_52),
    .I1(in_47)
  );
  //AND U139bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U139bar (
    .O(n827bar),
    .I0(in_52bar),
    .I1(in_47bar)
  );
  //OR U140
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U140 (
    .O(out[3]),
    .I0(n826),
    .I1(n825)
  );
  //AND U140bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U140bar (
    .O(outbar[3]),
    .I0(n826bar),
    .I1(n825bar)
  );
  //OR U141
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U141 (
    .O(n825),
    .I0(n824),
    .I1(n823)
  );
  //AND U141bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U141bar (
    .O(n825bar),
    .I0(n824bar),
    .I1(n823bar)
  );
  //OR U142
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U142 (
    .O(n823),
    .I0(n822),
    .I1(n821)
  );
  //AND U142bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U142bar (
    .O(n823bar),
    .I0(n822bar),
    .I1(n821bar)
  );
  //OR U143
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U143 (
    .O(n821),
    .I0(n820),
    .I1(n819)
  );
  //AND U143bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U143bar (
    .O(n821bar),
    .I0(n820bar),
    .I1(n819bar)
  );
  //OR U144
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U144 (
    .O(n822),
    .I0(n964),
    .I1(n818)
  );
  //AND U144bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U144bar (
    .O(n822bar),
    .I0(n964bar),
    .I1(n818bar)
  );
  //OR U145
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U145 (
    .O(n818),
    .I0(in[118]),
    .I1(n817)
  );
  //AND U145bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U145bar (
    .O(n818bar),
    .I0(inbar[118]),
    .I1(n817bar)
  );
  //OR U146
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U146 (
    .O(n964),
    .I0(n816),
    .I1(n815)
  );
  //AND U146bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U146bar (
    .O(n964bar),
    .I0(n816bar),
    .I1(n815bar)
  );
  //OR U147
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U147 (
    .O(n815),
    .I0(n814),
    .I1(n813)
  );
  //AND U147bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U147bar (
    .O(n815bar),
    .I0(n814bar),
    .I1(n813bar)
  );
  //OR U148
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U148 (
    .O(n813),
    .I0(n812),
    .I1(n811)
  );
  //AND U148bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U148bar (
    .O(n813bar),
    .I0(n812bar),
    .I1(n811bar)
  );
  //OR U149
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U149 (
    .O(n811),
    .I0(in[122]),
    .I1(in[111])
  );
  //AND U149bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U149bar (
    .O(n811bar),
    .I0(inbar[122]),
    .I1(inbar[111])
  );
  //OR U150
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U150 (
    .O(n812),
    .I0(in[154]),
    .I1(in[151])
  );
  //AND U150bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U150bar (
    .O(n812bar),
    .I0(inbar[154]),
    .I1(inbar[151])
  );
  //OR U151
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U151 (
    .O(n814),
    .I0(n810),
    .I1(n809)
  );
  //AND U151bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U151bar (
    .O(n814bar),
    .I0(n810bar),
    .I1(n809bar)
  );
  //OR U152
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U152 (
    .O(n809),
    .I0(in[187]),
    .I1(in[177])
  );
  //AND U152bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U152bar (
    .O(n809bar),
    .I0(inbar[187]),
    .I1(inbar[177])
  );
  //OR U153
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U153 (
    .O(n810),
    .I0(in[200]),
    .I1(in[192])
  );
  //AND U153bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U153bar (
    .O(n810bar),
    .I0(inbar[200]),
    .I1(inbar[192])
  );
  //OR U154
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U154 (
    .O(n816),
    .I0(n808),
    .I1(n807)
  );
  //AND U154bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U154bar (
    .O(n816bar),
    .I0(n808bar),
    .I1(n807bar)
  );
  //OR U155
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U155 (
    .O(n807),
    .I0(n806),
    .I1(n805)
  );
  //AND U155bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U155bar (
    .O(n807bar),
    .I0(n806bar),
    .I1(n805bar)
  );
  //OR U156
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U156 (
    .O(n805),
    .I0(in[225]),
    .I1(in[207])
  );
  //AND U156bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U156bar (
    .O(n805bar),
    .I0(inbar[225]),
    .I1(inbar[207])
  );
  //OR U157
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U157 (
    .O(n806),
    .I0(in[98]),
    .I1(in[226])
  );
  //AND U157bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U157bar (
    .O(n806bar),
    .I0(inbar[98]),
    .I1(inbar[226])
  );
  //OR U158
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U158 (
    .O(n808),
    .I0(n804),
    .I1(n803)
  );
  //AND U158bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U158bar (
    .O(n808bar),
    .I0(n804bar),
    .I1(n803bar)
  );
  //OR U159
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U159 (
    .O(n803),
    .I0(in_20),
    .I1(in_16)
  );
  //AND U159bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U159bar (
    .O(n803bar),
    .I0(in_20bar),
    .I1(in_16bar)
  );
  //OR U160
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U160 (
    .O(n804),
    .I0(in_55),
    .I1(in_45)
  );
  //AND U160bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U160bar (
    .O(n804bar),
    .I0(in_55bar),
    .I1(in_45bar)
  );
  //OR U161
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U161 (
    .O(n824),
    .I0(n802),
    .I1(n801)
  );
  //AND U161bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U161bar (
    .O(n824bar),
    .I0(n802bar),
    .I1(n801bar)
  );
  //OR U162
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U162 (
    .O(n801),
    .I0(in[162]),
    .I1(in[149])
  );
  //AND U162bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U162bar (
    .O(n801bar),
    .I0(inbar[162]),
    .I1(inbar[149])
  );
  //OR U163
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U163 (
    .O(n802),
    .I0(in[163]),
    .I1(n800)
  );
  //AND U163bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U163bar (
    .O(n802bar),
    .I0(inbar[163]),
    .I1(n800bar)
  );
  //OR U164
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U164 (
    .O(n800),
    .I0(in[191]),
    .I1(in[189])
  );
  //AND U164bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U164bar (
    .O(n800bar),
    .I0(inbar[191]),
    .I1(inbar[189])
  );
  //OR U165
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U165 (
    .O(n826),
    .I0(n799),
    .I1(n798)
  );
  //AND U165bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U165bar (
    .O(n826bar),
    .I0(n799bar),
    .I1(n798bar)
  );
  //OR U166
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U166 (
    .O(n798),
    .I0(n797),
    .I1(n796)
  );
  //AND U166bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U166bar (
    .O(n798bar),
    .I0(n797bar),
    .I1(n796bar)
  );
  //OR U167
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U167 (
    .O(n796),
    .I0(in[212]),
    .I1(in[193])
  );
  //AND U167bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U167bar (
    .O(n796bar),
    .I0(inbar[212]),
    .I1(inbar[193])
  );
  //OR U168
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U168 (
    .O(n797),
    .I0(in[238]),
    .I1(n795)
  );
  //AND U168bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U168bar (
    .O(n797bar),
    .I0(inbar[238]),
    .I1(n795bar)
  );
  //OR U169
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U169 (
    .O(n795),
    .I0(in[88]),
    .I1(in[247])
  );
  //AND U169bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U169bar (
    .O(n795bar),
    .I0(inbar[88]),
    .I1(inbar[247])
  );
  //OR U170
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U170 (
    .O(n799),
    .I0(n794),
    .I1(n793)
  );
  //AND U170bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U170bar (
    .O(n799bar),
    .I0(n794bar),
    .I1(n793bar)
  );
  //OR U171
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U171 (
    .O(n793),
    .I0(in[94]),
    .I1(in[92])
  );
  //AND U171bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U171bar (
    .O(n793bar),
    .I0(inbar[94]),
    .I1(inbar[92])
  );
  //OR U172
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U172 (
    .O(n794),
    .I0(in_52),
    .I1(n792)
  );
  //AND U172bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U172bar (
    .O(n794bar),
    .I0(in_52bar),
    .I1(n792bar)
  );
  //OR U173
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U173 (
    .O(n792),
    .I0(in_70),
    .I1(in_67)
  );
  //AND U173bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U173bar (
    .O(n792bar),
    .I0(in_70bar),
    .I1(in_67bar)
  );
  //OR U174
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U174 (
    .O(out[2]),
    .I0(n791),
    .I1(n790)
  );
  //AND U174bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U174bar (
    .O(outbar[2]),
    .I0(n791bar),
    .I1(n790bar)
  );
  //OR U175
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U175 (
    .O(n790),
    .I0(n789),
    .I1(n788)
  );
  //AND U175bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U175bar (
    .O(n790bar),
    .I0(n789bar),
    .I1(n788bar)
  );
  //OR U176
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U176 (
    .O(n788),
    .I0(n787),
    .I1(n786)
  );
  //AND U176bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U176bar (
    .O(n788bar),
    .I0(n787bar),
    .I1(n786bar)
  );
  //OR U177
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U177 (
    .O(n786),
    .I0(n819),
    .I1(n785)
  );
  //AND U177bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U177bar (
    .O(n786bar),
    .I0(n819bar),
    .I1(n785bar)
  );
  //OR U178
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U178 (
    .O(n819),
    .I0(n784),
    .I1(n783)
  );
  //AND U178bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U178bar (
    .O(n819bar),
    .I0(n784bar),
    .I1(n783bar)
  );
  //OR U179
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U179 (
    .O(n783),
    .I0(n782),
    .I1(n781)
  );
  //AND U179bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U179bar (
    .O(n783bar),
    .I0(n782bar),
    .I1(n781bar)
  );
  //OR U180
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U180 (
    .O(n781),
    .I0(n780),
    .I1(n779)
  );
  //AND U180bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U180bar (
    .O(n781bar),
    .I0(n780bar),
    .I1(n779bar)
  );
  //OR U181
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U181 (
    .O(n779),
    .I0(n962),
    .I1(n778)
  );
  //AND U181bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U181bar (
    .O(n779bar),
    .I0(n962bar),
    .I1(n778bar)
  );
  //OR U182
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U182 (
    .O(n962),
    .I0(n777),
    .I1(n776)
  );
  //AND U182bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U182bar (
    .O(n962bar),
    .I0(n777bar),
    .I1(n776bar)
  );
  //OR U183
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U183 (
    .O(n776),
    .I0(n775),
    .I1(n774)
  );
  //AND U183bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U183bar (
    .O(n776bar),
    .I0(n775bar),
    .I1(n774bar)
  );
  //OR U184
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U184 (
    .O(n774),
    .I0(n773),
    .I1(n772)
  );
  //AND U184bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U184bar (
    .O(n774bar),
    .I0(n773bar),
    .I1(n772bar)
  );
  //OR U185
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U185 (
    .O(n772),
    .I0(in[131]),
    .I1(in[120])
  );
  //AND U185bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U185bar (
    .O(n772bar),
    .I0(inbar[131]),
    .I1(inbar[120])
  );
  //OR U186
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U186 (
    .O(n773),
    .I0(in[153]),
    .I1(in[147])
  );
  //AND U186bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U186bar (
    .O(n773bar),
    .I0(inbar[153]),
    .I1(inbar[147])
  );
  //OR U187
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U187 (
    .O(n775),
    .I0(n771),
    .I1(n770)
  );
  //AND U187bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U187bar (
    .O(n775bar),
    .I0(n771bar),
    .I1(n770bar)
  );
  //OR U188
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U188 (
    .O(n770),
    .I0(in[170]),
    .I1(in[156])
  );
  //AND U188bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U188bar (
    .O(n770bar),
    .I0(inbar[170]),
    .I1(inbar[156])
  );
  //OR U189
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U189 (
    .O(n771),
    .I0(in[223]),
    .I1(in[190])
  );
  //AND U189bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U189bar (
    .O(n771bar),
    .I0(inbar[223]),
    .I1(inbar[190])
  );
  //OR U190
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U190 (
    .O(n777),
    .I0(n769),
    .I1(n768)
  );
  //AND U190bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U190bar (
    .O(n777bar),
    .I0(n769bar),
    .I1(n768bar)
  );
  //OR U191
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U191 (
    .O(n768),
    .I0(n767),
    .I1(n766)
  );
  //AND U191bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U191bar (
    .O(n768bar),
    .I0(n767bar),
    .I1(n766bar)
  );
  //OR U192
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U192 (
    .O(n766),
    .I0(in[236]),
    .I1(in[230])
  );
  //AND U192bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U192bar (
    .O(n766bar),
    .I0(inbar[236]),
    .I1(inbar[230])
  );
  //OR U193
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U193 (
    .O(n767),
    .I0(in[85]),
    .I1(in[240])
  );
  //AND U193bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U193bar (
    .O(n767bar),
    .I0(inbar[85]),
    .I1(inbar[240])
  );
  //OR U194
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U194 (
    .O(n769),
    .I0(n765),
    .I1(n764)
  );
  //AND U194bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U194bar (
    .O(n769bar),
    .I0(n765bar),
    .I1(n764bar)
  );
  //OR U195
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U195 (
    .O(n764),
    .I0(in_12),
    .I1(in[90])
  );
  //AND U195bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U195bar (
    .O(n764bar),
    .I0(in_12bar),
    .I1(inbar[90])
  );
  //OR U196
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U196 (
    .O(n765),
    .I0(in_39),
    .I1(in_28)
  );
  //AND U196bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U196bar (
    .O(n765bar),
    .I0(in_39bar),
    .I1(in_28bar)
  );
  //OR U197
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U197 (
    .O(n780),
    .I0(in[109]),
    .I1(n763)
  );
  //AND U197bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U197bar (
    .O(n780bar),
    .I0(inbar[109]),
    .I1(n763bar)
  );
  //OR U198
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U198 (
    .O(n782),
    .I0(n762),
    .I1(n761)
  );
  //AND U198bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U198bar (
    .O(n782bar),
    .I0(n762bar),
    .I1(n761bar)
  );
  //OR U199
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U199 (
    .O(n761),
    .I0(in[138]),
    .I1(in[129])
  );
  //AND U199bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U199bar (
    .O(n761bar),
    .I0(inbar[138]),
    .I1(inbar[129])
  );
  //OR U200
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U200 (
    .O(n762),
    .I0(in[157]),
    .I1(n760)
  );
  //AND U200bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U200bar (
    .O(n762bar),
    .I0(inbar[157]),
    .I1(n760bar)
  );
  //OR U201
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U201 (
    .O(n760),
    .I0(in[182]),
    .I1(in[167])
  );
  //AND U201bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U201bar (
    .O(n760bar),
    .I0(inbar[182]),
    .I1(inbar[167])
  );
  //OR U202
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U202 (
    .O(n784),
    .I0(n759),
    .I1(n758)
  );
  //AND U202bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U202bar (
    .O(n784bar),
    .I0(n759bar),
    .I1(n758bar)
  );
  //OR U203
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U203 (
    .O(n758),
    .I0(n757),
    .I1(n756)
  );
  //AND U203bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U203bar (
    .O(n758bar),
    .I0(n757bar),
    .I1(n756bar)
  );
  //OR U204
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U204 (
    .O(n756),
    .I0(in[195]),
    .I1(in[184])
  );
  //AND U204bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U204bar (
    .O(n756bar),
    .I0(inbar[195]),
    .I1(inbar[184])
  );
  //OR U205
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U205 (
    .O(n757),
    .I0(in[196]),
    .I1(n755)
  );
  //AND U205bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U205bar (
    .O(n757bar),
    .I0(inbar[196]),
    .I1(n755bar)
  );
  //OR U206
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U206 (
    .O(n755),
    .I0(in[215]),
    .I1(in[209])
  );
  //AND U206bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U206bar (
    .O(n755bar),
    .I0(inbar[215]),
    .I1(inbar[209])
  );
  //OR U207
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U207 (
    .O(n759),
    .I0(n754),
    .I1(n753)
  );
  //AND U207bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U207bar (
    .O(n759bar),
    .I0(n754bar),
    .I1(n753bar)
  );
  //OR U208
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U208 (
    .O(n753),
    .I0(in[93]),
    .I1(in[233])
  );
  //AND U208bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U208bar (
    .O(n753bar),
    .I0(inbar[93]),
    .I1(inbar[233])
  );
  //OR U209
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U209 (
    .O(n754),
    .I0(in_1),
    .I1(n752)
  );
  //AND U209bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U209bar (
    .O(n754bar),
    .I0(in_1bar),
    .I1(n752bar)
  );
  //OR U210
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U210 (
    .O(n752),
    .I0(in_69),
    .I1(in_66)
  );
  //AND U210bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U210bar (
    .O(n752bar),
    .I0(in_69bar),
    .I1(in_66bar)
  );
  //OR U211
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U211 (
    .O(n787),
    .I0(n966),
    .I1(n751)
  );
  //AND U211bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U211bar (
    .O(n787bar),
    .I0(n966bar),
    .I1(n751bar)
  );
  //OR U212
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U212 (
    .O(n751),
    .I0(in[134]),
    .I1(n750)
  );
  //AND U212bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U212bar (
    .O(n751bar),
    .I0(inbar[134]),
    .I1(n750bar)
  );
  //OR U213
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U213 (
    .O(n966),
    .I0(n749),
    .I1(n748)
  );
  //AND U213bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U213bar (
    .O(n966bar),
    .I0(n749bar),
    .I1(n748bar)
  );
  //OR U214
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U214 (
    .O(n748),
    .I0(n747),
    .I1(n746)
  );
  //AND U214bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U214bar (
    .O(n748bar),
    .I0(n747bar),
    .I1(n746bar)
  );
  //OR U215
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U215 (
    .O(n746),
    .I0(n745),
    .I1(n744)
  );
  //AND U215bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U215bar (
    .O(n746bar),
    .I0(n745bar),
    .I1(n744bar)
  );
  //OR U216
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U216 (
    .O(n744),
    .I0(in[136]),
    .I1(in[121])
  );
  //AND U216bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U216bar (
    .O(n744bar),
    .I0(inbar[136]),
    .I1(inbar[121])
  );
  //OR U217
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U217 (
    .O(n745),
    .I0(in[186]),
    .I1(in[174])
  );
  //AND U217bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U217bar (
    .O(n745bar),
    .I0(inbar[186]),
    .I1(inbar[174])
  );
  //OR U218
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U218 (
    .O(n747),
    .I0(n743),
    .I1(n742)
  );
  //AND U218bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U218bar (
    .O(n747bar),
    .I0(n743bar),
    .I1(n742bar)
  );
  //OR U219
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U219 (
    .O(n742),
    .I0(in[198]),
    .I1(in[197])
  );
  //AND U219bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U219bar (
    .O(n742bar),
    .I0(inbar[198]),
    .I1(inbar[197])
  );
  //OR U220
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U220 (
    .O(n743),
    .I0(in[214]),
    .I1(in[199])
  );
  //AND U220bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U220bar (
    .O(n743bar),
    .I0(inbar[214]),
    .I1(inbar[199])
  );
  //OR U221
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U221 (
    .O(n749),
    .I0(n741),
    .I1(n740)
  );
  //AND U221bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U221bar (
    .O(n749bar),
    .I0(n741bar),
    .I1(n740bar)
  );
  //OR U222
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U222 (
    .O(n740),
    .I0(n739),
    .I1(n738)
  );
  //AND U222bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U222bar (
    .O(n740bar),
    .I0(n739bar),
    .I1(n738bar)
  );
  //OR U223
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U223 (
    .O(n738),
    .I0(in[231]),
    .I1(in[220])
  );
  //AND U223bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U223bar (
    .O(n738bar),
    .I0(inbar[231]),
    .I1(inbar[220])
  );
  //OR U224
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U224 (
    .O(n739),
    .I0(in_25),
    .I1(in[245])
  );
  //AND U224bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U224bar (
    .O(n739bar),
    .I0(in_25bar),
    .I1(inbar[245])
  );
  //OR U225
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U225 (
    .O(n741),
    .I0(n737),
    .I1(n736)
  );
  //AND U225bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U225bar (
    .O(n741bar),
    .I0(n737bar),
    .I1(n736bar)
  );
  //OR U226
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U226 (
    .O(n736),
    .I0(in_53),
    .I1(in_29)
  );
  //AND U226bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U226bar (
    .O(n736bar),
    .I0(in_53bar),
    .I1(in_29bar)
  );
  //OR U227
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U227 (
    .O(n737),
    .I0(in_79),
    .I1(in_74)
  );
  //AND U227bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U227bar (
    .O(n737bar),
    .I0(in_79bar),
    .I1(in_74bar)
  );
  //OR U228
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U228 (
    .O(n789),
    .I0(n735),
    .I1(n734)
  );
  //AND U228bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U228bar (
    .O(n789bar),
    .I0(n735bar),
    .I1(n734bar)
  );
  //OR U229
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U229 (
    .O(n734),
    .I0(in[152]),
    .I1(in[140])
  );
  //AND U229bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U229bar (
    .O(n734bar),
    .I0(inbar[152]),
    .I1(inbar[140])
  );
  //OR U230
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U230 (
    .O(n735),
    .I0(in[155]),
    .I1(n733)
  );
  //AND U230bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U230bar (
    .O(n735bar),
    .I0(inbar[155]),
    .I1(n733bar)
  );
  //OR U231
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U231 (
    .O(n733),
    .I0(in[166]),
    .I1(in[165])
  );
  //AND U231bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U231bar (
    .O(n733bar),
    .I0(inbar[166]),
    .I1(inbar[165])
  );
  //OR U232
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U232 (
    .O(n791),
    .I0(n732),
    .I1(n731)
  );
  //AND U232bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U232bar (
    .O(n791bar),
    .I0(n732bar),
    .I1(n731bar)
  );
  //OR U233
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U233 (
    .O(n731),
    .I0(n730),
    .I1(n729)
  );
  //AND U233bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U233bar (
    .O(n731bar),
    .I0(n730bar),
    .I1(n729bar)
  );
  //OR U234
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U234 (
    .O(n729),
    .I0(in[202]),
    .I1(in[185])
  );
  //AND U234bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U234bar (
    .O(n729bar),
    .I0(inbar[202]),
    .I1(inbar[185])
  );
  //OR U235
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U235 (
    .O(n730),
    .I0(in[211]),
    .I1(n728)
  );
  //AND U235bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U235bar (
    .O(n730bar),
    .I0(inbar[211]),
    .I1(n728bar)
  );
  //OR U236
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U236 (
    .O(n728),
    .I0(in[255]),
    .I1(in[253])
  );
  //AND U236bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U236bar (
    .O(n728bar),
    .I0(inbar[255]),
    .I1(inbar[253])
  );
  //OR U237
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U237 (
    .O(n732),
    .I0(n727),
    .I1(n726)
  );
  //AND U237bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U237bar (
    .O(n732bar),
    .I0(n727bar),
    .I1(n726bar)
  );
  //OR U238
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U238 (
    .O(n726),
    .I0(in_35),
    .I1(in_15)
  );
  //AND U238bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U238bar (
    .O(n726bar),
    .I0(in_35bar),
    .I1(in_15bar)
  );
  //OR U239
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U239 (
    .O(n727),
    .I0(in_36),
    .I1(n725)
  );
  //AND U239bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U239bar (
    .O(n727bar),
    .I0(in_36bar),
    .I1(n725bar)
  );
  //OR U240
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U240 (
    .O(n725),
    .I0(in_48),
    .I1(in_40)
  );
  //AND U240bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U240bar (
    .O(n725bar),
    .I0(in_48bar),
    .I1(in_40bar)
  );
  //OR U241
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U241 (
    .O(out[1]),
    .I0(n724),
    .I1(n723)
  );
  //AND U241bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U241bar (
    .O(outbar[1]),
    .I0(n724bar),
    .I1(n723bar)
  );
  //OR U242
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U242 (
    .O(n723),
    .I0(n722),
    .I1(n721)
  );
  //AND U242bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U242bar (
    .O(n723bar),
    .I0(n722bar),
    .I1(n721bar)
  );
  //OR U243
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U243 (
    .O(n721),
    .I0(n720),
    .I1(n719)
  );
  //AND U243bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U243bar (
    .O(n721bar),
    .I0(n720bar),
    .I1(n719bar)
  );
  //OR U244
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U244 (
    .O(n719),
    .I0(n921),
    .I1(n887)
  );
  //AND U244bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U244bar (
    .O(n719bar),
    .I0(n921bar),
    .I1(n887bar)
  );
  //OR U245
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U245 (
    .O(n887),
    .I0(n718),
    .I1(n717)
  );
  //AND U245bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U245bar (
    .O(n887bar),
    .I0(n718bar),
    .I1(n717bar)
  );
  //OR U246
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U246 (
    .O(n717),
    .I0(n716),
    .I1(n715)
  );
  //AND U246bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U246bar (
    .O(n717bar),
    .I0(n716bar),
    .I1(n715bar)
  );
  //OR U247
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U247 (
    .O(n715),
    .I0(n714),
    .I1(n713)
  );
  //AND U247bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U247bar (
    .O(n715bar),
    .I0(n714bar),
    .I1(n713bar)
  );
  //OR U248
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U248 (
    .O(n713),
    .I0(in[116]),
    .I1(in[110])
  );
  //AND U248bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U248bar (
    .O(n713bar),
    .I0(inbar[116]),
    .I1(inbar[110])
  );
  //OR U249
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U249 (
    .O(n714),
    .I0(in[133]),
    .I1(in[130])
  );
  //AND U249bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U249bar (
    .O(n714bar),
    .I0(inbar[133]),
    .I1(inbar[130])
  );
  //OR U250
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U250 (
    .O(n716),
    .I0(n712),
    .I1(n711)
  );
  //AND U250bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U250bar (
    .O(n716bar),
    .I0(n712bar),
    .I1(n711bar)
  );
  //OR U251
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U251 (
    .O(n711),
    .I0(in[203]),
    .I1(in[135])
  );
  //AND U251bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U251bar (
    .O(n711bar),
    .I0(inbar[203]),
    .I1(inbar[135])
  );
  //OR U252
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U252 (
    .O(n712),
    .I0(in[232]),
    .I1(in[223])
  );
  //AND U252bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U252bar (
    .O(n712bar),
    .I0(inbar[232]),
    .I1(inbar[223])
  );
  //OR U253
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U253 (
    .O(n718),
    .I0(n710),
    .I1(n709)
  );
  //AND U253bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U253bar (
    .O(n718bar),
    .I0(n710bar),
    .I1(n709bar)
  );
  //OR U254
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U254 (
    .O(n709),
    .I0(n708),
    .I1(n707)
  );
  //AND U254bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U254bar (
    .O(n709bar),
    .I0(n708bar),
    .I1(n707bar)
  );
  //OR U255
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U255 (
    .O(n707),
    .I0(in[255]),
    .I1(in[233])
  );
  //AND U255bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U255bar (
    .O(n707bar),
    .I0(inbar[255]),
    .I1(inbar[233])
  );
  //OR U256
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U256 (
    .O(n708),
    .I0(in_53),
    .I1(in_34)
  );
  //AND U256bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U256bar (
    .O(n708bar),
    .I0(in_53bar),
    .I1(in_34bar)
  );
  //OR U257
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U257 (
    .O(n710),
    .I0(n706),
    .I1(n705)
  );
  //AND U257bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U257bar (
    .O(n710bar),
    .I0(n706bar),
    .I1(n705bar)
  );
  //OR U258
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U258 (
    .O(n705),
    .I0(in_57),
    .I1(in_55)
  );
  //AND U258bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U258bar (
    .O(n705bar),
    .I0(in_57bar),
    .I1(in_55bar)
  );
  //OR U259
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U259 (
    .O(n706),
    .I0(in_68),
    .I1(in_67)
  );
  //AND U259bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U259bar (
    .O(n706bar),
    .I0(in_68bar),
    .I1(in_67bar)
  );
  //OR U260
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U260 (
    .O(n921),
    .I0(n704),
    .I1(n703)
  );
  //AND U260bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U260bar (
    .O(n921bar),
    .I0(n704bar),
    .I1(n703bar)
  );
  //OR U261
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U261 (
    .O(n703),
    .I0(n702),
    .I1(n701)
  );
  //AND U261bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U261bar (
    .O(n703bar),
    .I0(n702bar),
    .I1(n701bar)
  );
  //OR U262
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U262 (
    .O(n701),
    .I0(n700),
    .I1(n699)
  );
  //AND U262bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U262bar (
    .O(n701bar),
    .I0(n700bar),
    .I1(n699bar)
  );
  //OR U263
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U263 (
    .O(n699),
    .I0(n944),
    .I1(n872)
  );
  //AND U263bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U263bar (
    .O(n699bar),
    .I0(n944bar),
    .I1(n872bar)
  );
  //OR U264
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U264 (
    .O(n872),
    .I0(n698),
    .I1(n697)
  );
  //AND U264bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U264bar (
    .O(n872bar),
    .I0(n698bar),
    .I1(n697bar)
  );
  //OR U265
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U265 (
    .O(n697),
    .I0(n696),
    .I1(n695)
  );
  //AND U265bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U265bar (
    .O(n697bar),
    .I0(n696bar),
    .I1(n695bar)
  );
  //OR U266
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U266 (
    .O(n695),
    .I0(n694),
    .I1(n693)
  );
  //AND U266bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U266bar (
    .O(n695bar),
    .I0(n694bar),
    .I1(n693bar)
  );
  //OR U267
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U267 (
    .O(n693),
    .I0(in[121]),
    .I1(in[102])
  );
  //AND U267bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U267bar (
    .O(n693bar),
    .I0(inbar[121]),
    .I1(inbar[102])
  );
  //OR U268
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U268 (
    .O(n694),
    .I0(in[162]),
    .I1(in[161])
  );
  //AND U268bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U268bar (
    .O(n694bar),
    .I0(inbar[162]),
    .I1(inbar[161])
  );
  //OR U269
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U269 (
    .O(n696),
    .I0(n692),
    .I1(n691)
  );
  //AND U269bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U269bar (
    .O(n696bar),
    .I0(n692bar),
    .I1(n691bar)
  );
  //OR U270
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U270 (
    .O(n691),
    .I0(in[192]),
    .I1(in[178])
  );
  //AND U270bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U270bar (
    .O(n691bar),
    .I0(inbar[192]),
    .I1(inbar[178])
  );
  //OR U271
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U271 (
    .O(n692),
    .I0(in[244]),
    .I1(in[209])
  );
  //AND U271bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U271bar (
    .O(n692bar),
    .I0(inbar[244]),
    .I1(inbar[209])
  );
  //OR U272
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U272 (
    .O(n698),
    .I0(n690),
    .I1(n689)
  );
  //AND U272bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U272bar (
    .O(n698bar),
    .I0(n690bar),
    .I1(n689bar)
  );
  //OR U273
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U273 (
    .O(n689),
    .I0(n688),
    .I1(n687)
  );
  //AND U273bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U273bar (
    .O(n689bar),
    .I0(n688bar),
    .I1(n687bar)
  );
  //OR U274
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U274 (
    .O(n687),
    .I0(in[90]),
    .I1(in[254])
  );
  //AND U274bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U274bar (
    .O(n687bar),
    .I0(inbar[90]),
    .I1(inbar[254])
  );
  //OR U275
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U275 (
    .O(n688),
    .I0(in_36),
    .I1(in_32)
  );
  //AND U275bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U275bar (
    .O(n688bar),
    .I0(in_36bar),
    .I1(in_32bar)
  );
  //OR U276
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U276 (
    .O(n690),
    .I0(n686),
    .I1(n685)
  );
  //AND U276bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U276bar (
    .O(n690bar),
    .I0(n686bar),
    .I1(n685bar)
  );
  //OR U277
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U277 (
    .O(n685),
    .I0(in_62),
    .I1(in_37)
  );
  //AND U277bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U277bar (
    .O(n685bar),
    .I0(in_62bar),
    .I1(in_37bar)
  );
  //OR U278
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U278 (
    .O(n686),
    .I0(in_75),
    .I1(in_73)
  );
  //AND U278bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U278bar (
    .O(n686bar),
    .I0(in_75bar),
    .I1(in_73bar)
  );
  //OR U279
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U279 (
    .O(n944),
    .I0(n684),
    .I1(n683)
  );
  //AND U279bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U279bar (
    .O(n944bar),
    .I0(n684bar),
    .I1(n683bar)
  );
  //OR U280
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U280 (
    .O(n683),
    .I0(n682),
    .I1(n681)
  );
  //AND U280bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U280bar (
    .O(n683bar),
    .I0(n682bar),
    .I1(n681bar)
  );
  //OR U281
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U281 (
    .O(n681),
    .I0(n680),
    .I1(n679)
  );
  //AND U281bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U281bar (
    .O(n681bar),
    .I0(n680bar),
    .I1(n679bar)
  );
  //OR U282
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U282 (
    .O(n679),
    .I0(in[171]),
    .I1(in[153])
  );
  //AND U282bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U282bar (
    .O(n679bar),
    .I0(inbar[171]),
    .I1(inbar[153])
  );
  //OR U283
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U283 (
    .O(n680),
    .I0(in[187]),
    .I1(in[176])
  );
  //AND U283bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U283bar (
    .O(n680bar),
    .I0(inbar[187]),
    .I1(inbar[176])
  );
  //OR U284
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U284 (
    .O(n682),
    .I0(n678),
    .I1(n677)
  );
  //AND U284bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U284bar (
    .O(n682bar),
    .I0(n678bar),
    .I1(n677bar)
  );
  //OR U285
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U285 (
    .O(n677),
    .I0(in[245]),
    .I1(in[211])
  );
  //AND U285bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U285bar (
    .O(n677bar),
    .I0(inbar[245]),
    .I1(inbar[211])
  );
  //OR U286
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U286 (
    .O(n678),
    .I0(in[97]),
    .I1(in[88])
  );
  //AND U286bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U286bar (
    .O(n678bar),
    .I0(inbar[97]),
    .I1(inbar[88])
  );
  //OR U287
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U287 (
    .O(n684),
    .I0(n676),
    .I1(n675)
  );
  //AND U287bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U287bar (
    .O(n684bar),
    .I0(n676bar),
    .I1(n675bar)
  );
  //OR U288
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U288 (
    .O(n675),
    .I0(n674),
    .I1(n673)
  );
  //AND U288bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U288bar (
    .O(n675bar),
    .I0(n674bar),
    .I1(n673bar)
  );
  //OR U289
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U289 (
    .O(n673),
    .I0(in_10),
    .I1(in_0)
  );
  //AND U289bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U289bar (
    .O(n673bar),
    .I0(in_10bar),
    .I1(in_0bar)
  );
  //OR U290
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U290 (
    .O(n674),
    .I0(in_59),
    .I1(in_5)
  );
  //AND U290bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U290bar (
    .O(n674bar),
    .I0(in_59bar),
    .I1(in_5bar)
  );
  //OR U291
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U291 (
    .O(n676),
    .I0(n672),
    .I1(n671)
  );
  //AND U291bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U291bar (
    .O(n676bar),
    .I0(n672bar),
    .I1(n671bar)
  );
  //OR U292
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U292 (
    .O(n671),
    .I0(in_60),
    .I1(in_6)
  );
  //AND U292bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U292bar (
    .O(n671bar),
    .I0(in_60bar),
    .I1(in_6bar)
  );
  //OR U293
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U293 (
    .O(n672),
    .I0(in_77),
    .I1(in_69)
  );
  //AND U293bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U293bar (
    .O(n672bar),
    .I0(in_77bar),
    .I1(in_69bar)
  );
  //OR U294
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U294 (
    .O(n700),
    .I0(in[113]),
    .I1(n864)
  );
  //AND U294bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U294bar (
    .O(n700bar),
    .I0(inbar[113]),
    .I1(n864bar)
  );
  //OR U295
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U295 (
    .O(n864),
    .I0(n670),
    .I1(n669)
  );
  //AND U295bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U295bar (
    .O(n864bar),
    .I0(n670bar),
    .I1(n669bar)
  );
  //OR U296
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U296 (
    .O(n669),
    .I0(n668),
    .I1(n667)
  );
  //AND U296bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U296bar (
    .O(n669bar),
    .I0(n668bar),
    .I1(n667bar)
  );
  //OR U297
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U297 (
    .O(n667),
    .I0(n666),
    .I1(n665)
  );
  //AND U297bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U297bar (
    .O(n667bar),
    .I0(n666bar),
    .I1(n665bar)
  );
  //OR U298
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U298 (
    .O(n665),
    .I0(in[125]),
    .I1(in[107])
  );
  //AND U298bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U298bar (
    .O(n665bar),
    .I0(inbar[125]),
    .I1(inbar[107])
  );
  //OR U299
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U299 (
    .O(n666),
    .I0(in[138]),
    .I1(in[126])
  );
  //AND U299bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U299bar (
    .O(n666bar),
    .I0(inbar[138]),
    .I1(inbar[126])
  );
  //OR U300
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U300 (
    .O(n668),
    .I0(n664),
    .I1(n663)
  );
  //AND U300bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U300bar (
    .O(n668bar),
    .I0(n664bar),
    .I1(n663bar)
  );
  //OR U301
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U301 (
    .O(n663),
    .I0(in[189]),
    .I1(in[143])
  );
  //AND U301bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U301bar (
    .O(n663bar),
    .I0(inbar[189]),
    .I1(inbar[143])
  );
  //OR U302
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U302 (
    .O(n664),
    .I0(in[99]),
    .I1(in[214])
  );
  //AND U302bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U302bar (
    .O(n664bar),
    .I0(inbar[99]),
    .I1(inbar[214])
  );
  //OR U303
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U303 (
    .O(n670),
    .I0(n662),
    .I1(n661)
  );
  //AND U303bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U303bar (
    .O(n670bar),
    .I0(n662bar),
    .I1(n661bar)
  );
  //OR U304
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U304 (
    .O(n661),
    .I0(n660),
    .I1(n659)
  );
  //AND U304bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U304bar (
    .O(n661bar),
    .I0(n660bar),
    .I1(n659bar)
  );
  //OR U305
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U305 (
    .O(n659),
    .I0(in_15),
    .I1(in_12)
  );
  //AND U305bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U305bar (
    .O(n659bar),
    .I0(in_15bar),
    .I1(in_12bar)
  );
  //OR U306
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U306 (
    .O(n660),
    .I0(in_20),
    .I1(in_2)
  );
  //AND U306bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U306bar (
    .O(n660bar),
    .I0(in_20bar),
    .I1(in_2bar)
  );
  //OR U307
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U307 (
    .O(n662),
    .I0(n658),
    .I1(n657)
  );
  //AND U307bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U307bar (
    .O(n662bar),
    .I0(n658bar),
    .I1(n657bar)
  );
  //OR U308
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U308 (
    .O(n657),
    .I0(in_30),
    .I1(in_3)
  );
  //AND U308bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U308bar (
    .O(n657bar),
    .I0(in_30bar),
    .I1(in_3bar)
  );
  //OR U309
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U309 (
    .O(n658),
    .I0(in_4),
    .I1(in_38)
  );
  //AND U309bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U309bar (
    .O(n658bar),
    .I0(in_4bar),
    .I1(in_38bar)
  );
  //OR U310
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U310 (
    .O(n702),
    .I0(n656),
    .I1(n655)
  );
  //AND U310bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U310bar (
    .O(n702bar),
    .I0(n656bar),
    .I1(n655bar)
  );
  //OR U311
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U311 (
    .O(n655),
    .I0(in[148]),
    .I1(in[137])
  );
  //AND U311bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U311bar (
    .O(n655bar),
    .I0(inbar[148]),
    .I1(inbar[137])
  );
  //OR U312
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U312 (
    .O(n656),
    .I0(in[149]),
    .I1(n654)
  );
  //AND U312bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U312bar (
    .O(n656bar),
    .I0(inbar[149]),
    .I1(n654bar)
  );
  //OR U313
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U313 (
    .O(n654),
    .I0(in[195]),
    .I1(in[190])
  );
  //AND U313bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U313bar (
    .O(n654bar),
    .I0(inbar[195]),
    .I1(inbar[190])
  );
  //OR U314
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U314 (
    .O(n704),
    .I0(n653),
    .I1(n652)
  );
  //AND U314bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U314bar (
    .O(n704bar),
    .I0(n653bar),
    .I1(n652bar)
  );
  //OR U315
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U315 (
    .O(n652),
    .I0(n651),
    .I1(n650)
  );
  //AND U315bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U315bar (
    .O(n652bar),
    .I0(n651bar),
    .I1(n650bar)
  );
  //OR U316
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U316 (
    .O(n650),
    .I0(in[98]),
    .I1(in[197])
  );
  //AND U316bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U316bar (
    .O(n650bar),
    .I0(inbar[98]),
    .I1(inbar[197])
  );
  //OR U317
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U317 (
    .O(n651),
    .I0(in_11),
    .I1(n649)
  );
  //AND U317bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U317bar (
    .O(n651bar),
    .I0(in_11bar),
    .I1(n649bar)
  );
  //OR U318
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U318 (
    .O(n649),
    .I0(in_26),
    .I1(in_14)
  );
  //AND U318bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U318bar (
    .O(n649bar),
    .I0(in_26bar),
    .I1(in_14bar)
  );
  //OR U319
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U319 (
    .O(n653),
    .I0(n648),
    .I1(n647)
  );
  //AND U319bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U319bar (
    .O(n653bar),
    .I0(n648bar),
    .I1(n647bar)
  );
  //OR U320
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U320 (
    .O(n647),
    .I0(in_35),
    .I1(in_27)
  );
  //AND U320bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U320bar (
    .O(n647bar),
    .I0(in_35bar),
    .I1(in_27bar)
  );
  //OR U321
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U321 (
    .O(n648),
    .I0(in_50),
    .I1(n646)
  );
  //AND U321bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U321bar (
    .O(n648bar),
    .I0(in_50bar),
    .I1(n646bar)
  );
  //OR U322
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U322 (
    .O(n646),
    .I0(in_78),
    .I1(in_61)
  );
  //AND U322bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U322bar (
    .O(n646bar),
    .I0(in_78bar),
    .I1(in_61bar)
  );
  //OR U323
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U323 (
    .O(n720),
    .I0(n942),
    .I1(n645)
  );
  //AND U323bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U323bar (
    .O(n720bar),
    .I0(n942bar),
    .I1(n645bar)
  );
  //OR U324
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U324 (
    .O(n645),
    .I0(in[106]),
    .I1(n863)
  );
  //AND U324bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U324bar (
    .O(n645bar),
    .I0(inbar[106]),
    .I1(n863bar)
  );
  //OR U325
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U325 (
    .O(n863),
    .I0(n644),
    .I1(n643)
  );
  //AND U325bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U325bar (
    .O(n863bar),
    .I0(n644bar),
    .I1(n643bar)
  );
  //OR U326
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U326 (
    .O(n643),
    .I0(n642),
    .I1(n641)
  );
  //AND U326bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U326bar (
    .O(n643bar),
    .I0(n642bar),
    .I1(n641bar)
  );
  //OR U327
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U327 (
    .O(n641),
    .I0(n640),
    .I1(n639)
  );
  //AND U327bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U327bar (
    .O(n641bar),
    .I0(n640bar),
    .I1(n639bar)
  );
  //OR U328
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U328 (
    .O(n639),
    .I0(in[127]),
    .I1(in[122])
  );
  //AND U328bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U328bar (
    .O(n639bar),
    .I0(inbar[127]),
    .I1(inbar[122])
  );
  //OR U329
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U329 (
    .O(n640),
    .I0(in[156]),
    .I1(in[132])
  );
  //AND U329bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U329bar (
    .O(n640bar),
    .I0(inbar[156]),
    .I1(inbar[132])
  );
  //OR U330
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U330 (
    .O(n642),
    .I0(n638),
    .I1(n637)
  );
  //AND U330bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U330bar (
    .O(n642bar),
    .I0(n638bar),
    .I1(n637bar)
  );
  //OR U331
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U331 (
    .O(n637),
    .I0(in[159]),
    .I1(in[157])
  );
  //AND U331bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U331bar (
    .O(n637bar),
    .I0(inbar[159]),
    .I1(inbar[157])
  );
  //OR U332
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U332 (
    .O(n638),
    .I0(in[185]),
    .I1(in[169])
  );
  //AND U332bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U332bar (
    .O(n638bar),
    .I0(inbar[185]),
    .I1(inbar[169])
  );
  //OR U333
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U333 (
    .O(n644),
    .I0(n636),
    .I1(n635)
  );
  //AND U333bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U333bar (
    .O(n644bar),
    .I0(n636bar),
    .I1(n635bar)
  );
  //OR U334
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U334 (
    .O(n635),
    .I0(n634),
    .I1(n633)
  );
  //AND U334bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U334bar (
    .O(n635bar),
    .I0(n634bar),
    .I1(n633bar)
  );
  //OR U335
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U335 (
    .O(n633),
    .I0(in[239]),
    .I1(in[218])
  );
  //AND U335bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U335bar (
    .O(n633bar),
    .I0(inbar[239]),
    .I1(inbar[218])
  );
  //OR U336
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U336 (
    .O(n634),
    .I0(in_13),
    .I1(in[87])
  );
  //AND U336bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U336bar (
    .O(n634bar),
    .I0(in_13bar),
    .I1(inbar[87])
  );
  //OR U337
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U337 (
    .O(n636),
    .I0(n632),
    .I1(n631)
  );
  //AND U337bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U337bar (
    .O(n636bar),
    .I0(n632bar),
    .I1(n631bar)
  );
  //OR U338
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U338 (
    .O(n631),
    .I0(in_72),
    .I1(in_70)
  );
  //AND U338bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U338bar (
    .O(n631bar),
    .I0(in_72bar),
    .I1(in_70bar)
  );
  //OR U339
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U339 (
    .O(n632),
    .I0(in_80),
    .I1(in_74)
  );
  //AND U339bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U339bar (
    .O(n632bar),
    .I0(in_80bar),
    .I1(in_74bar)
  );
  //OR U340
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U340 (
    .O(n942),
    .I0(n630),
    .I1(n629)
  );
  //AND U340bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U340bar (
    .O(n942bar),
    .I0(n630bar),
    .I1(n629bar)
  );
  //OR U341
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U341 (
    .O(n629),
    .I0(n628),
    .I1(n627)
  );
  //AND U341bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U341bar (
    .O(n629bar),
    .I0(n628bar),
    .I1(n627bar)
  );
  //OR U342
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U342 (
    .O(n627),
    .I0(n626),
    .I1(n625)
  );
  //AND U342bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U342bar (
    .O(n627bar),
    .I0(n626bar),
    .I1(n625bar)
  );
  //OR U343
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U343 (
    .O(n625),
    .I0(in[146]),
    .I1(in[100])
  );
  //AND U343bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U343bar (
    .O(n625bar),
    .I0(inbar[146]),
    .I1(inbar[100])
  );
  //OR U344
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U344 (
    .O(n626),
    .I0(in[168]),
    .I1(in[152])
  );
  //AND U344bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U344bar (
    .O(n626bar),
    .I0(inbar[168]),
    .I1(inbar[152])
  );
  //OR U345
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U345 (
    .O(n628),
    .I0(n624),
    .I1(n623)
  );
  //AND U345bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U345bar (
    .O(n628bar),
    .I0(n624bar),
    .I1(n623bar)
  );
  //OR U346
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U346 (
    .O(n623),
    .I0(in[199]),
    .I1(in[182])
  );
  //AND U346bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U346bar (
    .O(n623bar),
    .I0(inbar[199]),
    .I1(inbar[182])
  );
  //OR U347
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U347 (
    .O(n624),
    .I0(in[236]),
    .I1(in[204])
  );
  //AND U347bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U347bar (
    .O(n624bar),
    .I0(inbar[236]),
    .I1(inbar[204])
  );
  //OR U348
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U348 (
    .O(n630),
    .I0(n622),
    .I1(n621)
  );
  //AND U348bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U348bar (
    .O(n630bar),
    .I0(n622bar),
    .I1(n621bar)
  );
  //OR U349
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U349 (
    .O(n621),
    .I0(n620),
    .I1(n619)
  );
  //AND U349bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U349bar (
    .O(n621bar),
    .I0(n620bar),
    .I1(n619bar)
  );
  //OR U350
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U350 (
    .O(n619),
    .I0(in[89]),
    .I1(in[246])
  );
  //AND U350bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U350bar (
    .O(n619bar),
    .I0(inbar[89]),
    .I1(inbar[246])
  );
  //OR U351
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U351 (
    .O(n620),
    .I0(in[95]),
    .I1(in[92])
  );
  //AND U351bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U351bar (
    .O(n620bar),
    .I0(inbar[95]),
    .I1(inbar[92])
  );
  //OR U352
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U352 (
    .O(n622),
    .I0(n618),
    .I1(n617)
  );
  //AND U352bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U352bar (
    .O(n622bar),
    .I0(n618bar),
    .I1(n617bar)
  );
  //OR U353
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U353 (
    .O(n617),
    .I0(in_22),
    .I1(in_16)
  );
  //AND U353bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U353bar (
    .O(n617bar),
    .I0(in_22bar),
    .I1(in_16bar)
  );
  //OR U354
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U354 (
    .O(n618),
    .I0(in_51),
    .I1(in_49)
  );
  //AND U354bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U354bar (
    .O(n618bar),
    .I0(in_51bar),
    .I1(in_49bar)
  );
  //OR U355
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U355 (
    .O(n722),
    .I0(n616),
    .I1(n615)
  );
  //AND U355bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U355bar (
    .O(n722bar),
    .I0(n616bar),
    .I1(n615bar)
  );
  //OR U356
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U356 (
    .O(n615),
    .I0(in[158]),
    .I1(in[115])
  );
  //AND U356bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U356bar (
    .O(n615bar),
    .I0(inbar[158]),
    .I1(inbar[115])
  );
  //OR U357
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U357 (
    .O(n616),
    .I0(in[163]),
    .I1(n614)
  );
  //AND U357bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U357bar (
    .O(n616bar),
    .I0(inbar[163]),
    .I1(n614bar)
  );
  //OR U358
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U358 (
    .O(n614),
    .I0(in[206]),
    .I1(in[165])
  );
  //AND U358bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U358bar (
    .O(n614bar),
    .I0(inbar[206]),
    .I1(inbar[165])
  );
  //OR U359
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U359 (
    .O(n724),
    .I0(n613),
    .I1(n612)
  );
  //AND U359bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U359bar (
    .O(n724bar),
    .I0(n613bar),
    .I1(n612bar)
  );
  //OR U360
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U360 (
    .O(n612),
    .I0(n611),
    .I1(n610)
  );
  //AND U360bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U360bar (
    .O(n612bar),
    .I0(n611bar),
    .I1(n610bar)
  );
  //OR U361
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U361 (
    .O(n610),
    .I0(in[213]),
    .I1(in[207])
  );
  //AND U361bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U361bar (
    .O(n610bar),
    .I0(inbar[213]),
    .I1(inbar[207])
  );
  //OR U362
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U362 (
    .O(n611),
    .I0(in[215]),
    .I1(n609)
  );
  //AND U362bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U362bar (
    .O(n611bar),
    .I0(inbar[215]),
    .I1(n609bar)
  );
  //OR U363
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U363 (
    .O(n609),
    .I0(in[230]),
    .I1(in[220])
  );
  //AND U363bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U363bar (
    .O(n609bar),
    .I0(inbar[230]),
    .I1(inbar[220])
  );
  //OR U364
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U364 (
    .O(n613),
    .I0(n608),
    .I1(n607)
  );
  //AND U364bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U364bar (
    .O(n613bar),
    .I0(n608bar),
    .I1(n607bar)
  );
  //OR U365
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U365 (
    .O(n607),
    .I0(in[251]),
    .I1(in[234])
  );
  //AND U365bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U365bar (
    .O(n607bar),
    .I0(inbar[251]),
    .I1(inbar[234])
  );
  //OR U366
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U366 (
    .O(n608),
    .I0(in_17),
    .I1(n606)
  );
  //AND U366bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U366bar (
    .O(n608bar),
    .I0(in_17bar),
    .I1(n606bar)
  );
  //OR U367
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U367 (
    .O(n606),
    .I0(in_65),
    .I1(in_56)
  );
  //AND U367bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U367bar (
    .O(n606bar),
    .I0(in_65bar),
    .I1(in_56bar)
  );
  //OR U368
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U368 (
    .O(out[0]),
    .I0(n605),
    .I1(n604)
  );
  //AND U368bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U368bar (
    .O(outbar[0]),
    .I0(n605bar),
    .I1(n604bar)
  );
  //OR U369
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U369 (
    .O(n604),
    .I0(n603),
    .I1(n602)
  );
  //AND U369bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U369bar (
    .O(n604bar),
    .I0(n603bar),
    .I1(n602bar)
  );
  //OR U370
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U370 (
    .O(n602),
    .I0(n601),
    .I1(n600)
  );
  //AND U370bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U370bar (
    .O(n602bar),
    .I0(n601bar),
    .I1(n600bar)
  );
  //OR U371
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U371 (
    .O(n600),
    .I0(n820),
    .I1(n785)
  );
  //AND U371bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U371bar (
    .O(n600bar),
    .I0(n820bar),
    .I1(n785bar)
  );
  //OR U372
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U372 (
    .O(n785),
    .I0(n599),
    .I1(n598)
  );
  //AND U372bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U372bar (
    .O(n785bar),
    .I0(n599bar),
    .I1(n598bar)
  );
  //OR U373
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U373 (
    .O(n598),
    .I0(n597),
    .I1(n596)
  );
  //AND U373bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U373bar (
    .O(n598bar),
    .I0(n597bar),
    .I1(n596bar)
  );
  //OR U374
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U374 (
    .O(n596),
    .I0(n595),
    .I1(n594)
  );
  //AND U374bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U374bar (
    .O(n596bar),
    .I0(n595bar),
    .I1(n594bar)
  );
  //OR U375
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U375 (
    .O(n594),
    .I0(in[135]),
    .I1(in[104])
  );
  //AND U375bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U375bar (
    .O(n594bar),
    .I0(inbar[135]),
    .I1(inbar[104])
  );
  //OR U376
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U376 (
    .O(n595),
    .I0(in[188]),
    .I1(in[178])
  );
  //AND U376bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U376bar (
    .O(n595bar),
    .I0(inbar[188]),
    .I1(inbar[178])
  );
  //OR U377
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U377 (
    .O(n597),
    .I0(n593),
    .I1(n592)
  );
  //AND U377bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U377bar (
    .O(n597bar),
    .I0(n593bar),
    .I1(n592bar)
  );
  //OR U378
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U378 (
    .O(n592),
    .I0(in[217]),
    .I1(in[194])
  );
  //AND U378bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U378bar (
    .O(n592bar),
    .I0(inbar[217]),
    .I1(inbar[194])
  );
  //OR U379
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U379 (
    .O(n593),
    .I0(in[237]),
    .I1(in[218])
  );
  //AND U379bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U379bar (
    .O(n593bar),
    .I0(inbar[237]),
    .I1(inbar[218])
  );
  //OR U380
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U380 (
    .O(n599),
    .I0(n591),
    .I1(n590)
  );
  //AND U380bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U380bar (
    .O(n599bar),
    .I0(n591bar),
    .I1(n590bar)
  );
  //OR U381
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U381 (
    .O(n590),
    .I0(n589),
    .I1(n588)
  );
  //AND U381bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U381bar (
    .O(n590bar),
    .I0(n589bar),
    .I1(n588bar)
  );
  //OR U382
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U382 (
    .O(n588),
    .I0(in_2),
    .I1(in_10)
  );
  //AND U382bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U382bar (
    .O(n588bar),
    .I0(in_2bar),
    .I1(in_10bar)
  );
  //OR U383
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U383 (
    .O(n589),
    .I0(in_47),
    .I1(in_22)
  );
  //AND U383bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U383bar (
    .O(n589bar),
    .I0(in_47bar),
    .I1(in_22bar)
  );
  //OR U384
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U384 (
    .O(n591),
    .I0(n587),
    .I1(n586)
  );
  //AND U384bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U384bar (
    .O(n591bar),
    .I0(n587bar),
    .I1(n586bar)
  );
  //OR U385
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U385 (
    .O(n586),
    .I0(in_56),
    .I1(in_54)
  );
  //AND U385bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U385bar (
    .O(n586bar),
    .I0(in_56bar),
    .I1(in_54bar)
  );
  //OR U386
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U386 (
    .O(n587),
    .I0(in_63),
    .I1(in_61)
  );
  //AND U386bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U386bar (
    .O(n587bar),
    .I0(in_63bar),
    .I1(in_61bar)
  );
  //OR U387
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U387 (
    .O(n820),
    .I0(n585),
    .I1(n584)
  );
  //AND U387bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U387bar (
    .O(n820bar),
    .I0(n585bar),
    .I1(n584bar)
  );
  //OR U388
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U388 (
    .O(n584),
    .I0(n583),
    .I1(n582)
  );
  //AND U388bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U388bar (
    .O(n584bar),
    .I0(n583bar),
    .I1(n582bar)
  );
  //OR U389
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U389 (
    .O(n582),
    .I0(n581),
    .I1(n580)
  );
  //AND U389bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U389bar (
    .O(n582bar),
    .I0(n581bar),
    .I1(n580bar)
  );
  //OR U390
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U390 (
    .O(n580),
    .I0(in[158]),
    .I1(in[142])
  );
  //AND U390bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U390bar (
    .O(n580bar),
    .I0(inbar[158]),
    .I1(inbar[142])
  );
  //OR U391
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U391 (
    .O(n581),
    .I0(in[175]),
    .I1(in[164])
  );
  //AND U391bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U391bar (
    .O(n581bar),
    .I0(inbar[175]),
    .I1(inbar[164])
  );
  //OR U392
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U392 (
    .O(n583),
    .I0(n579),
    .I1(n578)
  );
  //AND U392bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U392bar (
    .O(n583bar),
    .I0(n579bar),
    .I1(n578bar)
  );
  //OR U393
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U393 (
    .O(n578),
    .I0(in[228]),
    .I1(in[204])
  );
  //AND U393bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U393bar (
    .O(n578bar),
    .I0(inbar[228]),
    .I1(inbar[204])
  );
  //OR U394
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U394 (
    .O(n579),
    .I0(in[91]),
    .I1(in[87])
  );
  //AND U394bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U394bar (
    .O(n579bar),
    .I0(inbar[91]),
    .I1(inbar[87])
  );
  //OR U395
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U395 (
    .O(n585),
    .I0(n577),
    .I1(n576)
  );
  //AND U395bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U395bar (
    .O(n585bar),
    .I0(n577bar),
    .I1(n576bar)
  );
  //OR U396
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U396 (
    .O(n576),
    .I0(n575),
    .I1(n574)
  );
  //AND U396bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U396bar (
    .O(n576bar),
    .I0(n575bar),
    .I1(n574bar)
  );
  //OR U397
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U397 (
    .O(n574),
    .I0(in_21),
    .I1(in_11)
  );
  //AND U397bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U397bar (
    .O(n574bar),
    .I0(in_21bar),
    .I1(in_11bar)
  );
  //OR U398
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U398 (
    .O(n575),
    .I0(in_5),
    .I1(in_3)
  );
  //AND U398bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U398bar (
    .O(n575bar),
    .I0(in_5bar),
    .I1(in_3bar)
  );
  //OR U399
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U399 (
    .O(n577),
    .I0(n573),
    .I1(n572)
  );
  //AND U399bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U399bar (
    .O(n577bar),
    .I0(n573bar),
    .I1(n572bar)
  );
  //OR U400
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U400 (
    .O(n572),
    .I0(in_68),
    .I1(in_64)
  );
  //AND U400bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U400bar (
    .O(n572bar),
    .I0(in_68bar),
    .I1(in_64bar)
  );
  //OR U401
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U401 (
    .O(n573),
    .I0(in_76),
    .I1(in_73)
  );
  //AND U401bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U401bar (
    .O(n573bar),
    .I0(in_76bar),
    .I1(in_73bar)
  );
  //OR U402
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U402 (
    .O(n601),
    .I0(n778),
    .I1(n571)
  );
  //AND U402bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U402bar (
    .O(n601bar),
    .I0(n778bar),
    .I1(n571bar)
  );
  //OR U403
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U403 (
    .O(n571),
    .I0(in[100]),
    .I1(n965)
  );
  //AND U403bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U403bar (
    .O(n571bar),
    .I0(inbar[100]),
    .I1(n965bar)
  );
  //OR U404
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U404 (
    .O(n965),
    .I0(n570),
    .I1(n569)
  );
  //AND U404bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U404bar (
    .O(n965bar),
    .I0(n570bar),
    .I1(n569bar)
  );
  //OR U405
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U405 (
    .O(n569),
    .I0(n568),
    .I1(n567)
  );
  //AND U405bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U405bar (
    .O(n569bar),
    .I0(n568bar),
    .I1(n567bar)
  );
  //OR U406
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U406 (
    .O(n567),
    .I0(n566),
    .I1(n565)
  );
  //AND U406bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U406bar (
    .O(n567bar),
    .I0(n566bar),
    .I1(n565bar)
  );
  //OR U407
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U407 (
    .O(n565),
    .I0(n817),
    .I1(n750)
  );
  //AND U407bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U407bar (
    .O(n565bar),
    .I0(n817bar),
    .I1(n750bar)
  );
  //OR U408
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U408 (
    .O(n750),
    .I0(n564),
    .I1(n563)
  );
  //AND U408bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U408bar (
    .O(n750bar),
    .I0(n564bar),
    .I1(n563bar)
  );
  //OR U409
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U409 (
    .O(n563),
    .I0(n562),
    .I1(n561)
  );
  //AND U409bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U409bar (
    .O(n563bar),
    .I0(n562bar),
    .I1(n561bar)
  );
  //OR U410
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U410 (
    .O(n561),
    .I0(n560),
    .I1(n559)
  );
  //AND U410bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U410bar (
    .O(n561bar),
    .I0(n560bar),
    .I1(n559bar)
  );
  //OR U411
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U411 (
    .O(n559),
    .I0(in[119]),
    .I1(in[103])
  );
  //AND U411bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U411bar (
    .O(n559bar),
    .I0(inbar[119]),
    .I1(inbar[103])
  );
  //OR U412
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U412 (
    .O(n560),
    .I0(in[137]),
    .I1(in[133])
  );
  //AND U412bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U412bar (
    .O(n560bar),
    .I0(inbar[137]),
    .I1(inbar[133])
  );
  //OR U413
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U413 (
    .O(n562),
    .I0(n558),
    .I1(n557)
  );
  //AND U413bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U413bar (
    .O(n562bar),
    .I0(n558bar),
    .I1(n557bar)
  );
  //OR U414
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U414 (
    .O(n557),
    .I0(in[176]),
    .I1(in[173])
  );
  //AND U414bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U414bar (
    .O(n557bar),
    .I0(inbar[176]),
    .I1(inbar[173])
  );
  //OR U415
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U415 (
    .O(n558),
    .I0(in[210]),
    .I1(in[181])
  );
  //AND U415bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U415bar (
    .O(n558bar),
    .I0(inbar[210]),
    .I1(inbar[181])
  );
  //OR U416
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U416 (
    .O(n564),
    .I0(n556),
    .I1(n555)
  );
  //AND U416bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U416bar (
    .O(n564bar),
    .I0(n556bar),
    .I1(n555bar)
  );
  //OR U417
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U417 (
    .O(n555),
    .I0(n554),
    .I1(n553)
  );
  //AND U417bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U417bar (
    .O(n555bar),
    .I0(n554bar),
    .I1(n553bar)
  );
  //OR U418
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U418 (
    .O(n553),
    .I0(in_13),
    .I1(in[234])
  );
  //AND U418bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U418bar (
    .O(n553bar),
    .I0(in_13bar),
    .I1(inbar[234])
  );
  //OR U419
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U419 (
    .O(n554),
    .I0(in_38),
    .I1(in_32)
  );
  //AND U419bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U419bar (
    .O(n554bar),
    .I0(in_38bar),
    .I1(in_32bar)
  );
  //OR U420
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U420 (
    .O(n556),
    .I0(n552),
    .I1(n551)
  );
  //AND U420bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U420bar (
    .O(n556bar),
    .I0(n552bar),
    .I1(n551bar)
  );
  //OR U421
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U421 (
    .O(n551),
    .I0(in_42),
    .I1(in_41)
  );
  //AND U421bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U421bar (
    .O(n551bar),
    .I0(in_42bar),
    .I1(in_41bar)
  );
  //OR U422
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U422 (
    .O(n552),
    .I0(in_7),
    .I1(in_49)
  );
  //AND U422bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U422bar (
    .O(n552bar),
    .I0(in_7bar),
    .I1(in_49bar)
  );
  //OR U423
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U423 (
    .O(n817),
    .I0(n550),
    .I1(n549)
  );
  //AND U423bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U423bar (
    .O(n817bar),
    .I0(n550bar),
    .I1(n549bar)
  );
  //OR U424
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U424 (
    .O(n549),
    .I0(n548),
    .I1(n547)
  );
  //AND U424bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U424bar (
    .O(n549bar),
    .I0(n548bar),
    .I1(n547bar)
  );
  //OR U425
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U425 (
    .O(n547),
    .I0(n546),
    .I1(n545)
  );
  //AND U425bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U425bar (
    .O(n547bar),
    .I0(n546bar),
    .I1(n545bar)
  );
  //OR U426
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U426 (
    .O(n545),
    .I0(in[159]),
    .I1(in[105])
  );
  //AND U426bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U426bar (
    .O(n545bar),
    .I0(inbar[159]),
    .I1(inbar[105])
  );
  //OR U427
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U427 (
    .O(n546),
    .I0(in[206]),
    .I1(in[183])
  );
  //AND U427bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U427bar (
    .O(n546bar),
    .I0(inbar[206]),
    .I1(inbar[183])
  );
  //OR U428
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U428 (
    .O(n548),
    .I0(n544),
    .I1(n543)
  );
  //AND U428bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U428bar (
    .O(n548bar),
    .I0(n544bar),
    .I1(n543bar)
  );
  //OR U429
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U429 (
    .O(n543),
    .I0(in[229]),
    .I1(in[219])
  );
  //AND U429bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U429bar (
    .O(n543bar),
    .I0(inbar[229]),
    .I1(inbar[219])
  );
  //OR U430
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U430 (
    .O(n544),
    .I0(in[235]),
    .I1(in[232])
  );
  //AND U430bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U430bar (
    .O(n544bar),
    .I0(inbar[235]),
    .I1(inbar[232])
  );
  //OR U431
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U431 (
    .O(n550),
    .I0(n542),
    .I1(n541)
  );
  //AND U431bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U431bar (
    .O(n550bar),
    .I0(n542bar),
    .I1(n541bar)
  );
  //OR U432
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U432 (
    .O(n541),
    .I0(n540),
    .I1(n539)
  );
  //AND U432bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U432bar (
    .O(n541bar),
    .I0(n540bar),
    .I1(n539bar)
  );
  //OR U433
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U433 (
    .O(n539),
    .I0(in[249]),
    .I1(in[242])
  );
  //AND U433bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U433bar (
    .O(n539bar),
    .I0(inbar[249]),
    .I1(inbar[242])
  );
  //OR U434
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U434 (
    .O(n540),
    .I0(in[89]),
    .I1(in[254])
  );
  //AND U434bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U434bar (
    .O(n540bar),
    .I0(inbar[89]),
    .I1(inbar[254])
  );
  //OR U435
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U435 (
    .O(n542),
    .I0(n538),
    .I1(n537)
  );
  //AND U435bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U435bar (
    .O(n542bar),
    .I0(n538bar),
    .I1(n537bar)
  );
  //OR U436
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U436 (
    .O(n537),
    .I0(in_14),
    .I1(in[99])
  );
  //AND U436bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U436bar (
    .O(n537bar),
    .I0(in_14bar),
    .I1(inbar[99])
  );
  //OR U437
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U437 (
    .O(n538),
    .I0(in_60),
    .I1(in_18)
  );
  //AND U437bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U437bar (
    .O(n538bar),
    .I0(in_60bar),
    .I1(in_18bar)
  );
  //OR U438
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U438 (
    .O(n566),
    .I0(in[113]),
    .I1(n763)
  );
  //AND U438bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U438bar (
    .O(n566bar),
    .I0(inbar[113]),
    .I1(n763bar)
  );
  //OR U439
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U439 (
    .O(n763),
    .I0(n536),
    .I1(n535)
  );
  //AND U439bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U439bar (
    .O(n763bar),
    .I0(n536bar),
    .I1(n535bar)
  );
  //OR U440
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U440 (
    .O(n535),
    .I0(n534),
    .I1(n533)
  );
  //AND U440bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U440bar (
    .O(n535bar),
    .I0(n534bar),
    .I1(n533bar)
  );
  //OR U441
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U441 (
    .O(n533),
    .I0(n532),
    .I1(n531)
  );
  //AND U441bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U441bar (
    .O(n533bar),
    .I0(n532bar),
    .I1(n531bar)
  );
  //OR U442
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U442 (
    .O(n531),
    .I0(in[115]),
    .I1(in[110])
  );
  //AND U442bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U442bar (
    .O(n531bar),
    .I0(inbar[115]),
    .I1(inbar[110])
  );
  //OR U443
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U443 (
    .O(n532),
    .I0(in[125]),
    .I1(in[117])
  );
  //AND U443bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U443bar (
    .O(n532bar),
    .I0(inbar[125]),
    .I1(inbar[117])
  );
  //OR U444
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U444 (
    .O(n534),
    .I0(n530),
    .I1(n529)
  );
  //AND U444bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U444bar (
    .O(n534bar),
    .I0(n530bar),
    .I1(n529bar)
  );
  //OR U445
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U445 (
    .O(n529),
    .I0(in[180]),
    .I1(in[128])
  );
  //AND U445bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U445bar (
    .O(n529bar),
    .I0(inbar[180]),
    .I1(inbar[128])
  );
  //OR U446
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U446 (
    .O(n530),
    .I0(in[205]),
    .I1(in[201])
  );
  //AND U446bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U446bar (
    .O(n530bar),
    .I0(inbar[205]),
    .I1(inbar[201])
  );
  //OR U447
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U447 (
    .O(n536),
    .I0(n528),
    .I1(n527)
  );
  //AND U447bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U447bar (
    .O(n536bar),
    .I0(n528bar),
    .I1(n527bar)
  );
  //OR U448
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U448 (
    .O(n527),
    .I0(n526),
    .I1(n525)
  );
  //AND U448bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U448bar (
    .O(n527bar),
    .I0(n526bar),
    .I1(n525bar)
  );
  //OR U449
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U449 (
    .O(n525),
    .I0(in[244]),
    .I1(in[239])
  );
  //AND U449bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U449bar (
    .O(n525bar),
    .I0(inbar[244]),
    .I1(inbar[239])
  );
  //OR U450
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U450 (
    .O(n526),
    .I0(in[95]),
    .I1(in[83])
  );
  //AND U450bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U450bar (
    .O(n526bar),
    .I0(inbar[95]),
    .I1(inbar[83])
  );
  //OR U451
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U451 (
    .O(n528),
    .I0(n524),
    .I1(n523)
  );
  //AND U451bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U451bar (
    .O(n528bar),
    .I0(n524bar),
    .I1(n523bar)
  );
  //OR U452
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U452 (
    .O(n523),
    .I0(in_24),
    .I1(in[97])
  );
  //AND U452bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U452bar (
    .O(n523bar),
    .I0(in_24bar),
    .I1(inbar[97])
  );
  //OR U453
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U453 (
    .O(n524),
    .I0(in_33),
    .I1(in_27)
  );
  //AND U453bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U453bar (
    .O(n524bar),
    .I0(in_33bar),
    .I1(in_27bar)
  );
  //OR U454
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U454 (
    .O(n568),
    .I0(n522),
    .I1(n521)
  );
  //AND U454bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U454bar (
    .O(n568bar),
    .I0(n522bar),
    .I1(n521bar)
  );
  //OR U455
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U455 (
    .O(n521),
    .I0(in[145]),
    .I1(in[126])
  );
  //AND U455bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U455bar (
    .O(n521bar),
    .I0(inbar[145]),
    .I1(inbar[126])
  );
  //OR U456
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U456 (
    .O(n522),
    .I0(in[169]),
    .I1(n520)
  );
  //AND U456bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U456bar (
    .O(n522bar),
    .I0(inbar[169]),
    .I1(n520bar)
  );
  //OR U457
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U457 (
    .O(n520),
    .I0(in[221]),
    .I1(in[172])
  );
  //AND U457bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U457bar (
    .O(n520bar),
    .I0(inbar[221]),
    .I1(inbar[172])
  );
  //OR U458
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U458 (
    .O(n570),
    .I0(n519),
    .I1(n518)
  );
  //AND U458bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U458bar (
    .O(n570bar),
    .I0(n519bar),
    .I1(n518bar)
  );
  //OR U459
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U459 (
    .O(n518),
    .I0(n517),
    .I1(n516)
  );
  //AND U459bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U459bar (
    .O(n518bar),
    .I0(n517bar),
    .I1(n516bar)
  );
  //OR U460
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U460 (
    .O(n516),
    .I0(in[241]),
    .I1(in[224])
  );
  //AND U460bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U460bar (
    .O(n516bar),
    .I0(inbar[241]),
    .I1(inbar[224])
  );
  //OR U461
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U461 (
    .O(n517),
    .I0(in[86]),
    .I1(n515)
  );
  //AND U461bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U461bar (
    .O(n517bar),
    .I0(inbar[86]),
    .I1(n515bar)
  );
  //OR U462
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U462 (
    .O(n515),
    .I0(in_43),
    .I1(in_34)
  );
  //AND U462bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U462bar (
    .O(n515bar),
    .I0(in_43bar),
    .I1(in_34bar)
  );
  //OR U463
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U463 (
    .O(n519),
    .I0(n514),
    .I1(n513)
  );
  //AND U463bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U463bar (
    .O(n519bar),
    .I0(n514bar),
    .I1(n513bar)
  );
  //OR U464
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U464 (
    .O(n513),
    .I0(in_65),
    .I1(in_51)
  );
  //AND U464bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U464bar (
    .O(n513bar),
    .I0(in_65bar),
    .I1(in_51bar)
  );
  //OR U465
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U465 (
    .O(n514),
    .I0(in_75),
    .I1(n512)
  );
  //AND U465bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U465bar (
    .O(n514bar),
    .I0(in_75bar),
    .I1(n512bar)
  );
  //OR U466
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U466 (
    .O(n512),
    .I0(in_81),
    .I1(in_77)
  );
  //AND U466bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U466bar (
    .O(n512bar),
    .I0(in_81bar),
    .I1(in_77bar)
  );
  //OR U467
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U467 (
    .O(n778),
    .I0(n511),
    .I1(n510)
  );
  //AND U467bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U467bar (
    .O(n778bar),
    .I0(n511bar),
    .I1(n510bar)
  );
  //OR U468
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U468 (
    .O(n510),
    .I0(n509),
    .I1(n508)
  );
  //AND U468bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U468bar (
    .O(n510bar),
    .I0(n509bar),
    .I1(n508bar)
  );
  //OR U469
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U469 (
    .O(n508),
    .I0(n507),
    .I1(n506)
  );
  //AND U469bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U469bar (
    .O(n508bar),
    .I0(n507bar),
    .I1(n506bar)
  );
  //OR U470
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U470 (
    .O(n506),
    .I0(in[107]),
    .I1(in[101])
  );
  //AND U470bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U470bar (
    .O(n506bar),
    .I0(inbar[107]),
    .I1(inbar[101])
  );
  //OR U471
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U471 (
    .O(n507),
    .I0(in[139]),
    .I1(in[132])
  );
  //AND U471bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U471bar (
    .O(n507bar),
    .I0(inbar[139]),
    .I1(inbar[132])
  );
  //OR U472
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U472 (
    .O(n509),
    .I0(n505),
    .I1(n504)
  );
  //AND U472bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U472bar (
    .O(n509bar),
    .I0(n505bar),
    .I1(n504bar)
  );
  //OR U473
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U473 (
    .O(n504),
    .I0(in[146]),
    .I1(in[141])
  );
  //AND U473bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U473bar (
    .O(n504bar),
    .I0(inbar[146]),
    .I1(inbar[141])
  );
  //OR U474
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U474 (
    .O(n505),
    .I0(in[203]),
    .I1(in[179])
  );
  //AND U474bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U474bar (
    .O(n505bar),
    .I0(inbar[203]),
    .I1(inbar[179])
  );
  //OR U475
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U475 (
    .O(n511),
    .I0(n503),
    .I1(n502)
  );
  //AND U475bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U475bar (
    .O(n511bar),
    .I0(n503bar),
    .I1(n502bar)
  );
  //OR U476
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U476 (
    .O(n502),
    .I0(n501),
    .I1(n500)
  );
  //AND U476bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U476bar (
    .O(n502bar),
    .I0(n501bar),
    .I1(n500bar)
  );
  //OR U477
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U477 (
    .O(n500),
    .I0(in[243]),
    .I1(in[222])
  );
  //AND U477bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U477bar (
    .O(n500bar),
    .I0(inbar[243]),
    .I1(inbar[222])
  );
  //OR U478
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U478 (
    .O(n501),
    .I0(in[251]),
    .I1(in[250])
  );
  //AND U478bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U478bar (
    .O(n501bar),
    .I0(inbar[251]),
    .I1(inbar[250])
  );
  //OR U479
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U479 (
    .O(n503),
    .I0(n499),
    .I1(n498)
  );
  //AND U479bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U479bar (
    .O(n503bar),
    .I0(n499bar),
    .I1(n498bar)
  );
  //OR U480
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U480 (
    .O(n498),
    .I0(in_37),
    .I1(in_19)
  );
  //AND U480bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U480bar (
    .O(n498bar),
    .I0(in_37bar),
    .I1(in_19bar)
  );
  //OR U481
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U481 (
    .O(n499),
    .I0(in_78),
    .I1(in_6)
  );
  //AND U481bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U481bar (
    .O(n499bar),
    .I0(in_78bar),
    .I1(in_6bar)
  );
  //OR U482
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U482 (
    .O(n603),
    .I0(n497),
    .I1(n496)
  );
  //AND U482bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U482bar (
    .O(n603bar),
    .I0(n497bar),
    .I1(n496bar)
  );
  //OR U483
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U483 (
    .O(n496),
    .I0(in[112]),
    .I1(in[102])
  );
  //AND U483bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U483bar (
    .O(n496bar),
    .I0(inbar[112]),
    .I1(inbar[102])
  );
  //OR U484
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U484 (
    .O(n497),
    .I0(in[123]),
    .I1(n495)
  );
  //AND U484bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U484bar (
    .O(n497bar),
    .I0(inbar[123]),
    .I1(n495bar)
  );
  //OR U485
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U485 (
    .O(n495),
    .I0(in[143]),
    .I1(in[130])
  );
  //AND U485bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U485bar (
    .O(n495bar),
    .I0(inbar[143]),
    .I1(inbar[130])
  );
  //OR U486
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U486 (
    .O(n605),
    .I0(n494),
    .I1(n493)
  );
  //AND U486bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U486bar (
    .O(n605bar),
    .I0(n494bar),
    .I1(n493bar)
  );
  //OR U487
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U487 (
    .O(n493),
    .I0(n492),
    .I1(n491)
  );
  //AND U487bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U487bar (
    .O(n493bar),
    .I0(n492bar),
    .I1(n491bar)
  );
  //OR U488
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U488 (
    .O(n491),
    .I0(in[216]),
    .I1(in[213])
  );
  //AND U488bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U488bar (
    .O(n491bar),
    .I0(inbar[216]),
    .I1(inbar[213])
  );
  //OR U489
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U489 (
    .O(n492),
    .I0(in[227]),
    .I1(n490)
  );
  //AND U489bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U489bar (
    .O(n492bar),
    .I0(inbar[227]),
    .I1(n490bar)
  );
  //OR U490
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U490 (
    .O(n490),
    .I0(in_0),
    .I1(in[248])
  );
  //AND U490bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U490bar (
    .O(n490bar),
    .I0(in_0bar),
    .I1(inbar[248])
  );
  //OR U491
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U491 (
    .O(n494),
    .I0(n489),
    .I1(n488)
  );
  //AND U491bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U491bar (
    .O(n494bar),
    .I0(n489bar),
    .I1(n488bar)
  );
  //OR U492
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U492 (
    .O(n488),
    .I0(in_46),
    .I1(in_44)
  );
  //AND U492bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U492bar (
    .O(n488bar),
    .I0(in_46bar),
    .I1(in_44bar)
  );
  //OR U493
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U493 (
    .O(n489),
    .I0(in_50),
    .I1(n487)
  );
  //AND U493bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U493bar (
    .O(n489bar),
    .I0(in_50bar),
    .I1(n487bar)
  );
  //OR U494
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U494 (
    .O(n487),
    .I0(in_9),
    .I1(in_80)
  );
  //AND U494bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U494bar (
    .O(n487bar),
    .I0(in_9bar),
    .I1(in_80bar)
  );
endmodule

module sBox_7 ( in, out );

  input wire [7:0] in;
//input_done

  output wire [7:0] out;
//output_done

  wire [255:0] decodeOut;
//wire_done

  decode_7 dec ( .in(in), .out(decodeOut) );
  encode_7 enc ( .in(decodeOut), .out(out) );
endmodule

module CD2_29 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD2_30 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD2_31 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD2_32 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD4_15 ( a, b, y );

  input wire [3:0] a;
  input wire [3:0] b;
  wire [3:0] abar;
  wire [3:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
//input_done

  output wire [15:0] y;
  wire [15:0] ybar;
//output_done

//wire_done

  //AND U1
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1 (
    .O(y[9]),
    .I0(b[1]),
    .I1(a[2])
  );
  //OR U1bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1bar (
    .O(ybar[9]),
    .I0(bbar[1]),
    .I1(abar[2])
  );
  //AND U2
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2 (
    .O(y[8]),
    .I0(b[0]),
    .I1(a[2])
  );
  //OR U2bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2bar (
    .O(ybar[8]),
    .I0(bbar[0]),
    .I1(abar[2])
  );
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[7]),
    .I0(b[3]),
    .I1(a[1])
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[7]),
    .I0(bbar[3]),
    .I1(abar[1])
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[6]),
    .I0(b[2]),
    .I1(a[1])
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[6]),
    .I0(bbar[2]),
    .I1(abar[1])
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[5]),
    .I0(a[1]),
    .I1(b[1])
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[5]),
    .I0(abar[1]),
    .I1(bbar[1])
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[4]),
    .I0(a[1]),
    .I1(b[0])
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[4]),
    .I0(abar[1]),
    .I1(bbar[0])
  );
  //AND U7
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7 (
    .O(y[3]),
    .I0(a[0]),
    .I1(b[3])
  );
  //OR U7bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7bar (
    .O(ybar[3]),
    .I0(abar[0]),
    .I1(bbar[3])
  );
  //AND U8
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8 (
    .O(y[2]),
    .I0(a[0]),
    .I1(b[2])
  );
  //OR U8bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8bar (
    .O(ybar[2]),
    .I0(abar[0]),
    .I1(bbar[2])
  );
  //AND U9
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9 (
    .O(y[1]),
    .I0(a[0]),
    .I1(b[1])
  );
  //OR U9bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9bar (
    .O(ybar[1]),
    .I0(abar[0]),
    .I1(bbar[1])
  );
  //AND U10
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10 (
    .O(y[15]),
    .I0(a[3]),
    .I1(b[3])
  );
  //OR U10bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10bar (
    .O(ybar[15]),
    .I0(abar[3]),
    .I1(bbar[3])
  );
  //AND U11
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11 (
    .O(y[14]),
    .I0(a[3]),
    .I1(b[2])
  );
  //OR U11bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11bar (
    .O(ybar[14]),
    .I0(abar[3]),
    .I1(bbar[2])
  );
  //AND U12
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12 (
    .O(y[13]),
    .I0(a[3]),
    .I1(b[1])
  );
  //OR U12bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12bar (
    .O(ybar[13]),
    .I0(abar[3]),
    .I1(bbar[1])
  );
  //AND U13
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13 (
    .O(y[12]),
    .I0(a[3]),
    .I1(b[0])
  );
  //OR U13bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13bar (
    .O(ybar[12]),
    .I0(abar[3]),
    .I1(bbar[0])
  );
  //AND U14
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14 (
    .O(y[11]),
    .I0(b[3]),
    .I1(a[2])
  );
  //OR U14bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14bar (
    .O(ybar[11]),
    .I0(bbar[3]),
    .I1(abar[2])
  );
  //AND U15
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15 (
    .O(y[10]),
    .I0(b[2]),
    .I1(a[2])
  );
  //OR U15bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15bar (
    .O(ybar[10]),
    .I0(bbar[2]),
    .I1(abar[2])
  );
  //AND U16
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16 (
    .O(y[0]),
    .I0(a[0]),
    .I1(b[0])
  );
  //OR U16bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16bar (
    .O(ybar[0]),
    .I0(abar[0]),
    .I1(bbar[0])
  );
endmodule

module CD4_16 ( a, b, y );

  input wire [3:0] a;
  input wire [3:0] b;
  wire [3:0] abar;
  wire [3:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
//input_done

  output wire [15:0] y;
  wire [15:0] ybar;
//output_done

//wire_done

  //AND U1
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1 (
    .O(y[9]),
    .I0(b[1]),
    .I1(a[2])
  );
  //OR U1bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1bar (
    .O(ybar[9]),
    .I0(bbar[1]),
    .I1(abar[2])
  );
  //AND U2
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2 (
    .O(y[8]),
    .I0(b[0]),
    .I1(a[2])
  );
  //OR U2bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2bar (
    .O(ybar[8]),
    .I0(bbar[0]),
    .I1(abar[2])
  );
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[7]),
    .I0(b[3]),
    .I1(a[1])
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[7]),
    .I0(bbar[3]),
    .I1(abar[1])
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[6]),
    .I0(b[2]),
    .I1(a[1])
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[6]),
    .I0(bbar[2]),
    .I1(abar[1])
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[5]),
    .I0(a[1]),
    .I1(b[1])
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[5]),
    .I0(abar[1]),
    .I1(bbar[1])
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[4]),
    .I0(a[1]),
    .I1(b[0])
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[4]),
    .I0(abar[1]),
    .I1(bbar[0])
  );
  //AND U7
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7 (
    .O(y[3]),
    .I0(a[0]),
    .I1(b[3])
  );
  //OR U7bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7bar (
    .O(ybar[3]),
    .I0(abar[0]),
    .I1(bbar[3])
  );
  //AND U8
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8 (
    .O(y[2]),
    .I0(a[0]),
    .I1(b[2])
  );
  //OR U8bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8bar (
    .O(ybar[2]),
    .I0(abar[0]),
    .I1(bbar[2])
  );
  //AND U9
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9 (
    .O(y[1]),
    .I0(a[0]),
    .I1(b[1])
  );
  //OR U9bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9bar (
    .O(ybar[1]),
    .I0(abar[0]),
    .I1(bbar[1])
  );
  //AND U10
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10 (
    .O(y[15]),
    .I0(a[3]),
    .I1(b[3])
  );
  //OR U10bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10bar (
    .O(ybar[15]),
    .I0(abar[3]),
    .I1(bbar[3])
  );
  //AND U11
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11 (
    .O(y[14]),
    .I0(a[3]),
    .I1(b[2])
  );
  //OR U11bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11bar (
    .O(ybar[14]),
    .I0(abar[3]),
    .I1(bbar[2])
  );
  //AND U12
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12 (
    .O(y[13]),
    .I0(a[3]),
    .I1(b[1])
  );
  //OR U12bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12bar (
    .O(ybar[13]),
    .I0(abar[3]),
    .I1(bbar[1])
  );
  //AND U13
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13 (
    .O(y[12]),
    .I0(a[3]),
    .I1(b[0])
  );
  //OR U13bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13bar (
    .O(ybar[12]),
    .I0(abar[3]),
    .I1(bbar[0])
  );
  //AND U14
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14 (
    .O(y[11]),
    .I0(b[3]),
    .I1(a[2])
  );
  //OR U14bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14bar (
    .O(ybar[11]),
    .I0(bbar[3]),
    .I1(abar[2])
  );
  //AND U15
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15 (
    .O(y[10]),
    .I0(b[2]),
    .I1(a[2])
  );
  //OR U15bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15bar (
    .O(ybar[10]),
    .I0(bbar[2]),
    .I1(abar[2])
  );
  //AND U16
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16 (
    .O(y[0]),
    .I0(a[0]),
    .I1(b[0])
  );
  //OR U16bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16bar (
    .O(ybar[0]),
    .I0(abar[0]),
    .I1(bbar[0])
  );
endmodule

module CD16_8 ( a, b, y );

  input wire [15:0] a;
  input wire [15:0] b;
  wire [15:0] abar;
  wire [15:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign abar[8] = ~a[8];
  assign abar[9] = ~a[9];
  assign abar[10] = ~a[10];
  assign abar[11] = ~a[11];
  assign abar[12] = ~a[12];
  assign abar[13] = ~a[13];
  assign abar[14] = ~a[14];
  assign abar[15] = ~a[15];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign bbar[8] = ~b[8];
  assign bbar[9] = ~b[9];
  assign bbar[10] = ~b[10];
  assign bbar[11] = ~b[11];
  assign bbar[12] = ~b[12];
  assign bbar[13] = ~b[13];
  assign bbar[14] = ~b[14];
  assign bbar[15] = ~b[15];
//input_done

  output wire [255:0] y;
  wire [255:0] ybar;
//output_done

//wire_done

  //AND U1
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1 (
    .O(y[9]),
    .I0(b[9]),
    .I1(a[0])
  );
  //OR U1bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1bar (
    .O(ybar[9]),
    .I0(bbar[9]),
    .I1(abar[0])
  );
  //AND U2
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2 (
    .O(y[99]),
    .I0(b[3]),
    .I1(a[6])
  );
  //OR U2bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2bar (
    .O(ybar[99]),
    .I0(bbar[3]),
    .I1(abar[6])
  );
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[98]),
    .I0(b[2]),
    .I1(a[6])
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[98]),
    .I0(bbar[2]),
    .I1(abar[6])
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[97]),
    .I0(b[1]),
    .I1(a[6])
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[97]),
    .I0(bbar[1]),
    .I1(abar[6])
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[96]),
    .I0(b[0]),
    .I1(a[6])
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[96]),
    .I0(bbar[0]),
    .I1(abar[6])
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[95]),
    .I0(b[15]),
    .I1(a[5])
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[95]),
    .I0(bbar[15]),
    .I1(abar[5])
  );
  //AND U7
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7 (
    .O(y[94]),
    .I0(b[14]),
    .I1(a[5])
  );
  //OR U7bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7bar (
    .O(ybar[94]),
    .I0(bbar[14]),
    .I1(abar[5])
  );
  //AND U8
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8 (
    .O(y[93]),
    .I0(b[13]),
    .I1(a[5])
  );
  //OR U8bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8bar (
    .O(ybar[93]),
    .I0(bbar[13]),
    .I1(abar[5])
  );
  //AND U9
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9 (
    .O(y[92]),
    .I0(b[12]),
    .I1(a[5])
  );
  //OR U9bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9bar (
    .O(ybar[92]),
    .I0(bbar[12]),
    .I1(abar[5])
  );
  //AND U10
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10 (
    .O(y[91]),
    .I0(b[11]),
    .I1(a[5])
  );
  //OR U10bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10bar (
    .O(ybar[91]),
    .I0(bbar[11]),
    .I1(abar[5])
  );
  //AND U11
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11 (
    .O(y[90]),
    .I0(b[10]),
    .I1(a[5])
  );
  //OR U11bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11bar (
    .O(ybar[90]),
    .I0(bbar[10]),
    .I1(abar[5])
  );
  //AND U12
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12 (
    .O(y[8]),
    .I0(b[8]),
    .I1(a[0])
  );
  //OR U12bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12bar (
    .O(ybar[8]),
    .I0(bbar[8]),
    .I1(abar[0])
  );
  //AND U13
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13 (
    .O(y[89]),
    .I0(a[5]),
    .I1(b[9])
  );
  //OR U13bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13bar (
    .O(ybar[89]),
    .I0(abar[5]),
    .I1(bbar[9])
  );
  //AND U14
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14 (
    .O(y[88]),
    .I0(b[8]),
    .I1(a[5])
  );
  //OR U14bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14bar (
    .O(ybar[88]),
    .I0(bbar[8]),
    .I1(abar[5])
  );
  //AND U15
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15 (
    .O(y[87]),
    .I0(b[7]),
    .I1(a[5])
  );
  //OR U15bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15bar (
    .O(ybar[87]),
    .I0(bbar[7]),
    .I1(abar[5])
  );
  //AND U16
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16 (
    .O(y[86]),
    .I0(b[6]),
    .I1(a[5])
  );
  //OR U16bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16bar (
    .O(ybar[86]),
    .I0(bbar[6]),
    .I1(abar[5])
  );
  //AND U17
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U17 (
    .O(y[85]),
    .I0(b[5]),
    .I1(a[5])
  );
  //OR U17bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U17bar (
    .O(ybar[85]),
    .I0(bbar[5]),
    .I1(abar[5])
  );
  //AND U18
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U18 (
    .O(y[84]),
    .I0(b[4]),
    .I1(a[5])
  );
  //OR U18bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U18bar (
    .O(ybar[84]),
    .I0(bbar[4]),
    .I1(abar[5])
  );
  //AND U19
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U19 (
    .O(y[83]),
    .I0(a[5]),
    .I1(b[3])
  );
  //OR U19bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U19bar (
    .O(ybar[83]),
    .I0(abar[5]),
    .I1(bbar[3])
  );
  //AND U20
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U20 (
    .O(y[82]),
    .I0(a[5]),
    .I1(b[2])
  );
  //OR U20bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U20bar (
    .O(ybar[82]),
    .I0(abar[5]),
    .I1(bbar[2])
  );
  //AND U21
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U21 (
    .O(y[81]),
    .I0(a[5]),
    .I1(b[1])
  );
  //OR U21bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U21bar (
    .O(ybar[81]),
    .I0(abar[5]),
    .I1(bbar[1])
  );
  //AND U22
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U22 (
    .O(y[80]),
    .I0(a[5]),
    .I1(b[0])
  );
  //OR U22bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U22bar (
    .O(ybar[80]),
    .I0(abar[5]),
    .I1(bbar[0])
  );
  //AND U23
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U23 (
    .O(y[7]),
    .I0(b[7]),
    .I1(a[0])
  );
  //OR U23bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U23bar (
    .O(ybar[7]),
    .I0(bbar[7]),
    .I1(abar[0])
  );
  //AND U24
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U24 (
    .O(y[79]),
    .I0(a[4]),
    .I1(b[15])
  );
  //OR U24bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U24bar (
    .O(ybar[79]),
    .I0(abar[4]),
    .I1(bbar[15])
  );
  //AND U25
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U25 (
    .O(y[78]),
    .I0(a[4]),
    .I1(b[14])
  );
  //OR U25bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U25bar (
    .O(ybar[78]),
    .I0(abar[4]),
    .I1(bbar[14])
  );
  //AND U26
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U26 (
    .O(y[77]),
    .I0(a[4]),
    .I1(b[13])
  );
  //OR U26bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U26bar (
    .O(ybar[77]),
    .I0(abar[4]),
    .I1(bbar[13])
  );
  //AND U27
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U27 (
    .O(y[76]),
    .I0(a[4]),
    .I1(b[12])
  );
  //OR U27bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U27bar (
    .O(ybar[76]),
    .I0(abar[4]),
    .I1(bbar[12])
  );
  //AND U28
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U28 (
    .O(y[75]),
    .I0(a[4]),
    .I1(b[11])
  );
  //OR U28bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U28bar (
    .O(ybar[75]),
    .I0(abar[4]),
    .I1(bbar[11])
  );
  //AND U29
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U29 (
    .O(y[74]),
    .I0(a[4]),
    .I1(b[10])
  );
  //OR U29bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U29bar (
    .O(ybar[74]),
    .I0(abar[4]),
    .I1(bbar[10])
  );
  //AND U30
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U30 (
    .O(y[73]),
    .I0(a[4]),
    .I1(b[9])
  );
  //OR U30bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U30bar (
    .O(ybar[73]),
    .I0(abar[4]),
    .I1(bbar[9])
  );
  //AND U31
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U31 (
    .O(y[72]),
    .I0(a[4]),
    .I1(b[8])
  );
  //OR U31bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U31bar (
    .O(ybar[72]),
    .I0(abar[4]),
    .I1(bbar[8])
  );
  //AND U32
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U32 (
    .O(y[71]),
    .I0(a[4]),
    .I1(b[7])
  );
  //OR U32bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U32bar (
    .O(ybar[71]),
    .I0(abar[4]),
    .I1(bbar[7])
  );
  //AND U33
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U33 (
    .O(y[70]),
    .I0(a[4]),
    .I1(b[6])
  );
  //OR U33bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U33bar (
    .O(ybar[70]),
    .I0(abar[4]),
    .I1(bbar[6])
  );
  //AND U34
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U34 (
    .O(y[6]),
    .I0(b[6]),
    .I1(a[0])
  );
  //OR U34bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U34bar (
    .O(ybar[6]),
    .I0(bbar[6]),
    .I1(abar[0])
  );
  //AND U35
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U35 (
    .O(y[69]),
    .I0(a[4]),
    .I1(b[5])
  );
  //OR U35bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U35bar (
    .O(ybar[69]),
    .I0(abar[4]),
    .I1(bbar[5])
  );
  //AND U36
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U36 (
    .O(y[68]),
    .I0(a[4]),
    .I1(b[4])
  );
  //OR U36bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U36bar (
    .O(ybar[68]),
    .I0(abar[4]),
    .I1(bbar[4])
  );
  //AND U37
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U37 (
    .O(y[67]),
    .I0(a[4]),
    .I1(b[3])
  );
  //OR U37bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U37bar (
    .O(ybar[67]),
    .I0(abar[4]),
    .I1(bbar[3])
  );
  //AND U38
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U38 (
    .O(y[66]),
    .I0(a[4]),
    .I1(b[2])
  );
  //OR U38bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U38bar (
    .O(ybar[66]),
    .I0(abar[4]),
    .I1(bbar[2])
  );
  //AND U39
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U39 (
    .O(y[65]),
    .I0(a[4]),
    .I1(b[1])
  );
  //OR U39bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U39bar (
    .O(ybar[65]),
    .I0(abar[4]),
    .I1(bbar[1])
  );
  //AND U40
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U40 (
    .O(y[64]),
    .I0(a[4]),
    .I1(b[0])
  );
  //OR U40bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U40bar (
    .O(ybar[64]),
    .I0(abar[4]),
    .I1(bbar[0])
  );
  //AND U41
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U41 (
    .O(y[63]),
    .I0(a[3]),
    .I1(b[15])
  );
  //OR U41bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U41bar (
    .O(ybar[63]),
    .I0(abar[3]),
    .I1(bbar[15])
  );
  //AND U42
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U42 (
    .O(y[62]),
    .I0(a[3]),
    .I1(b[14])
  );
  //OR U42bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U42bar (
    .O(ybar[62]),
    .I0(abar[3]),
    .I1(bbar[14])
  );
  //AND U43
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U43 (
    .O(y[61]),
    .I0(a[3]),
    .I1(b[13])
  );
  //OR U43bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U43bar (
    .O(ybar[61]),
    .I0(abar[3]),
    .I1(bbar[13])
  );
  //AND U44
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U44 (
    .O(y[60]),
    .I0(a[3]),
    .I1(b[12])
  );
  //OR U44bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U44bar (
    .O(ybar[60]),
    .I0(abar[3]),
    .I1(bbar[12])
  );
  //AND U45
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U45 (
    .O(y[5]),
    .I0(b[5]),
    .I1(a[0])
  );
  //OR U45bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U45bar (
    .O(ybar[5]),
    .I0(bbar[5]),
    .I1(abar[0])
  );
  //AND U46
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U46 (
    .O(y[59]),
    .I0(a[3]),
    .I1(b[11])
  );
  //OR U46bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U46bar (
    .O(ybar[59]),
    .I0(abar[3]),
    .I1(bbar[11])
  );
  //AND U47
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U47 (
    .O(y[58]),
    .I0(a[3]),
    .I1(b[10])
  );
  //OR U47bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U47bar (
    .O(ybar[58]),
    .I0(abar[3]),
    .I1(bbar[10])
  );
  //AND U48
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U48 (
    .O(y[57]),
    .I0(a[3]),
    .I1(b[9])
  );
  //OR U48bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U48bar (
    .O(ybar[57]),
    .I0(abar[3]),
    .I1(bbar[9])
  );
  //AND U49
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U49 (
    .O(y[56]),
    .I0(a[3]),
    .I1(b[8])
  );
  //OR U49bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U49bar (
    .O(ybar[56]),
    .I0(abar[3]),
    .I1(bbar[8])
  );
  //AND U50
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U50 (
    .O(y[55]),
    .I0(a[3]),
    .I1(b[7])
  );
  //OR U50bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U50bar (
    .O(ybar[55]),
    .I0(abar[3]),
    .I1(bbar[7])
  );
  //AND U51
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U51 (
    .O(y[54]),
    .I0(a[3]),
    .I1(b[6])
  );
  //OR U51bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U51bar (
    .O(ybar[54]),
    .I0(abar[3]),
    .I1(bbar[6])
  );
  //AND U52
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U52 (
    .O(y[53]),
    .I0(a[3]),
    .I1(b[5])
  );
  //OR U52bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U52bar (
    .O(ybar[53]),
    .I0(abar[3]),
    .I1(bbar[5])
  );
  //AND U53
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U53 (
    .O(y[52]),
    .I0(a[3]),
    .I1(b[4])
  );
  //OR U53bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U53bar (
    .O(ybar[52]),
    .I0(abar[3]),
    .I1(bbar[4])
  );
  //AND U54
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U54 (
    .O(y[51]),
    .I0(a[3]),
    .I1(b[3])
  );
  //OR U54bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U54bar (
    .O(ybar[51]),
    .I0(abar[3]),
    .I1(bbar[3])
  );
  //AND U55
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U55 (
    .O(y[50]),
    .I0(a[3]),
    .I1(b[2])
  );
  //OR U55bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U55bar (
    .O(ybar[50]),
    .I0(abar[3]),
    .I1(bbar[2])
  );
  //AND U56
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U56 (
    .O(y[4]),
    .I0(b[4]),
    .I1(a[0])
  );
  //OR U56bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U56bar (
    .O(ybar[4]),
    .I0(bbar[4]),
    .I1(abar[0])
  );
  //AND U57
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U57 (
    .O(y[49]),
    .I0(a[3]),
    .I1(b[1])
  );
  //OR U57bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U57bar (
    .O(ybar[49]),
    .I0(abar[3]),
    .I1(bbar[1])
  );
  //AND U58
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U58 (
    .O(y[48]),
    .I0(a[3]),
    .I1(b[0])
  );
  //OR U58bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U58bar (
    .O(ybar[48]),
    .I0(abar[3]),
    .I1(bbar[0])
  );
  //AND U59
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U59 (
    .O(y[47]),
    .I0(a[2]),
    .I1(b[15])
  );
  //OR U59bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U59bar (
    .O(ybar[47]),
    .I0(abar[2]),
    .I1(bbar[15])
  );
  //AND U60
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U60 (
    .O(y[46]),
    .I0(a[2]),
    .I1(b[14])
  );
  //OR U60bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U60bar (
    .O(ybar[46]),
    .I0(abar[2]),
    .I1(bbar[14])
  );
  //AND U61
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U61 (
    .O(y[45]),
    .I0(a[2]),
    .I1(b[13])
  );
  //OR U61bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U61bar (
    .O(ybar[45]),
    .I0(abar[2]),
    .I1(bbar[13])
  );
  //AND U62
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U62 (
    .O(y[44]),
    .I0(a[2]),
    .I1(b[12])
  );
  //OR U62bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U62bar (
    .O(ybar[44]),
    .I0(abar[2]),
    .I1(bbar[12])
  );
  //AND U63
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U63 (
    .O(y[43]),
    .I0(a[2]),
    .I1(b[11])
  );
  //OR U63bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U63bar (
    .O(ybar[43]),
    .I0(abar[2]),
    .I1(bbar[11])
  );
  //AND U64
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U64 (
    .O(y[42]),
    .I0(a[2]),
    .I1(b[10])
  );
  //OR U64bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U64bar (
    .O(ybar[42]),
    .I0(abar[2]),
    .I1(bbar[10])
  );
  //AND U65
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U65 (
    .O(y[41]),
    .I0(a[2]),
    .I1(b[9])
  );
  //OR U65bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U65bar (
    .O(ybar[41]),
    .I0(abar[2]),
    .I1(bbar[9])
  );
  //AND U66
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U66 (
    .O(y[40]),
    .I0(a[2]),
    .I1(b[8])
  );
  //OR U66bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U66bar (
    .O(ybar[40]),
    .I0(abar[2]),
    .I1(bbar[8])
  );
  //AND U67
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U67 (
    .O(y[3]),
    .I0(b[3]),
    .I1(a[0])
  );
  //OR U67bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U67bar (
    .O(ybar[3]),
    .I0(bbar[3]),
    .I1(abar[0])
  );
  //AND U68
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U68 (
    .O(y[39]),
    .I0(a[2]),
    .I1(b[7])
  );
  //OR U68bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U68bar (
    .O(ybar[39]),
    .I0(abar[2]),
    .I1(bbar[7])
  );
  //AND U69
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U69 (
    .O(y[38]),
    .I0(a[2]),
    .I1(b[6])
  );
  //OR U69bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U69bar (
    .O(ybar[38]),
    .I0(abar[2]),
    .I1(bbar[6])
  );
  //AND U70
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U70 (
    .O(y[37]),
    .I0(a[2]),
    .I1(b[5])
  );
  //OR U70bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U70bar (
    .O(ybar[37]),
    .I0(abar[2]),
    .I1(bbar[5])
  );
  //AND U71
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U71 (
    .O(y[36]),
    .I0(a[2]),
    .I1(b[4])
  );
  //OR U71bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U71bar (
    .O(ybar[36]),
    .I0(abar[2]),
    .I1(bbar[4])
  );
  //AND U72
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U72 (
    .O(y[35]),
    .I0(a[2]),
    .I1(b[3])
  );
  //OR U72bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U72bar (
    .O(ybar[35]),
    .I0(abar[2]),
    .I1(bbar[3])
  );
  //AND U73
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U73 (
    .O(y[34]),
    .I0(a[2]),
    .I1(b[2])
  );
  //OR U73bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U73bar (
    .O(ybar[34]),
    .I0(abar[2]),
    .I1(bbar[2])
  );
  //AND U74
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U74 (
    .O(y[33]),
    .I0(a[2]),
    .I1(b[1])
  );
  //OR U74bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U74bar (
    .O(ybar[33]),
    .I0(abar[2]),
    .I1(bbar[1])
  );
  //AND U75
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U75 (
    .O(y[32]),
    .I0(a[2]),
    .I1(b[0])
  );
  //OR U75bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U75bar (
    .O(ybar[32]),
    .I0(abar[2]),
    .I1(bbar[0])
  );
  //AND U76
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U76 (
    .O(y[31]),
    .I0(a[1]),
    .I1(b[15])
  );
  //OR U76bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U76bar (
    .O(ybar[31]),
    .I0(abar[1]),
    .I1(bbar[15])
  );
  //AND U77
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U77 (
    .O(y[30]),
    .I0(a[1]),
    .I1(b[14])
  );
  //OR U77bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U77bar (
    .O(ybar[30]),
    .I0(abar[1]),
    .I1(bbar[14])
  );
  //AND U78
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U78 (
    .O(y[2]),
    .I0(b[2]),
    .I1(a[0])
  );
  //OR U78bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U78bar (
    .O(ybar[2]),
    .I0(bbar[2]),
    .I1(abar[0])
  );
  //AND U79
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U79 (
    .O(y[29]),
    .I0(a[1]),
    .I1(b[13])
  );
  //OR U79bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U79bar (
    .O(ybar[29]),
    .I0(abar[1]),
    .I1(bbar[13])
  );
  //AND U80
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U80 (
    .O(y[28]),
    .I0(a[1]),
    .I1(b[12])
  );
  //OR U80bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U80bar (
    .O(ybar[28]),
    .I0(abar[1]),
    .I1(bbar[12])
  );
  //AND U81
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U81 (
    .O(y[27]),
    .I0(a[1]),
    .I1(b[11])
  );
  //OR U81bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U81bar (
    .O(ybar[27]),
    .I0(abar[1]),
    .I1(bbar[11])
  );
  //AND U82
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U82 (
    .O(y[26]),
    .I0(a[1]),
    .I1(b[10])
  );
  //OR U82bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U82bar (
    .O(ybar[26]),
    .I0(abar[1]),
    .I1(bbar[10])
  );
  //AND U83
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U83 (
    .O(y[25]),
    .I0(a[1]),
    .I1(b[9])
  );
  //OR U83bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U83bar (
    .O(ybar[25]),
    .I0(abar[1]),
    .I1(bbar[9])
  );
  //AND U84
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U84 (
    .O(y[255]),
    .I0(a[15]),
    .I1(b[15])
  );
  //OR U84bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U84bar (
    .O(ybar[255]),
    .I0(abar[15]),
    .I1(bbar[15])
  );
  //AND U85
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U85 (
    .O(y[254]),
    .I0(a[15]),
    .I1(b[14])
  );
  //OR U85bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U85bar (
    .O(ybar[254]),
    .I0(abar[15]),
    .I1(bbar[14])
  );
  //AND U86
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U86 (
    .O(y[253]),
    .I0(a[15]),
    .I1(b[13])
  );
  //OR U86bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U86bar (
    .O(ybar[253]),
    .I0(abar[15]),
    .I1(bbar[13])
  );
  //AND U87
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U87 (
    .O(y[252]),
    .I0(a[15]),
    .I1(b[12])
  );
  //OR U87bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U87bar (
    .O(ybar[252]),
    .I0(abar[15]),
    .I1(bbar[12])
  );
  //AND U88
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U88 (
    .O(y[251]),
    .I0(a[15]),
    .I1(b[11])
  );
  //OR U88bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U88bar (
    .O(ybar[251]),
    .I0(abar[15]),
    .I1(bbar[11])
  );
  //AND U89
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U89 (
    .O(y[250]),
    .I0(a[15]),
    .I1(b[10])
  );
  //OR U89bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U89bar (
    .O(ybar[250]),
    .I0(abar[15]),
    .I1(bbar[10])
  );
  //AND U90
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U90 (
    .O(y[24]),
    .I0(a[1]),
    .I1(b[8])
  );
  //OR U90bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U90bar (
    .O(ybar[24]),
    .I0(abar[1]),
    .I1(bbar[8])
  );
  //AND U91
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U91 (
    .O(y[249]),
    .I0(a[15]),
    .I1(b[9])
  );
  //OR U91bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U91bar (
    .O(ybar[249]),
    .I0(abar[15]),
    .I1(bbar[9])
  );
  //AND U92
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U92 (
    .O(y[248]),
    .I0(a[15]),
    .I1(b[8])
  );
  //OR U92bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U92bar (
    .O(ybar[248]),
    .I0(abar[15]),
    .I1(bbar[8])
  );
  //AND U93
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U93 (
    .O(y[247]),
    .I0(a[15]),
    .I1(b[7])
  );
  //OR U93bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U93bar (
    .O(ybar[247]),
    .I0(abar[15]),
    .I1(bbar[7])
  );
  //AND U94
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U94 (
    .O(y[246]),
    .I0(a[15]),
    .I1(b[6])
  );
  //OR U94bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U94bar (
    .O(ybar[246]),
    .I0(abar[15]),
    .I1(bbar[6])
  );
  //AND U95
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U95 (
    .O(y[245]),
    .I0(a[15]),
    .I1(b[5])
  );
  //OR U95bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U95bar (
    .O(ybar[245]),
    .I0(abar[15]),
    .I1(bbar[5])
  );
  //AND U96
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U96 (
    .O(y[244]),
    .I0(a[15]),
    .I1(b[4])
  );
  //OR U96bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U96bar (
    .O(ybar[244]),
    .I0(abar[15]),
    .I1(bbar[4])
  );
  //AND U97
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U97 (
    .O(y[243]),
    .I0(a[15]),
    .I1(b[3])
  );
  //OR U97bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U97bar (
    .O(ybar[243]),
    .I0(abar[15]),
    .I1(bbar[3])
  );
  //AND U98
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U98 (
    .O(y[242]),
    .I0(a[15]),
    .I1(b[2])
  );
  //OR U98bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U98bar (
    .O(ybar[242]),
    .I0(abar[15]),
    .I1(bbar[2])
  );
  //AND U99
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U99 (
    .O(y[241]),
    .I0(a[15]),
    .I1(b[1])
  );
  //OR U99bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U99bar (
    .O(ybar[241]),
    .I0(abar[15]),
    .I1(bbar[1])
  );
  //AND U100
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U100 (
    .O(y[240]),
    .I0(a[15]),
    .I1(b[0])
  );
  //OR U100bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U100bar (
    .O(ybar[240]),
    .I0(abar[15]),
    .I1(bbar[0])
  );
  //AND U101
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U101 (
    .O(y[23]),
    .I0(a[1]),
    .I1(b[7])
  );
  //OR U101bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U101bar (
    .O(ybar[23]),
    .I0(abar[1]),
    .I1(bbar[7])
  );
  //AND U102
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U102 (
    .O(y[239]),
    .I0(a[14]),
    .I1(b[15])
  );
  //OR U102bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U102bar (
    .O(ybar[239]),
    .I0(abar[14]),
    .I1(bbar[15])
  );
  //AND U103
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U103 (
    .O(y[238]),
    .I0(a[14]),
    .I1(b[14])
  );
  //OR U103bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U103bar (
    .O(ybar[238]),
    .I0(abar[14]),
    .I1(bbar[14])
  );
  //AND U104
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U104 (
    .O(y[237]),
    .I0(a[14]),
    .I1(b[13])
  );
  //OR U104bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U104bar (
    .O(ybar[237]),
    .I0(abar[14]),
    .I1(bbar[13])
  );
  //AND U105
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U105 (
    .O(y[236]),
    .I0(a[14]),
    .I1(b[12])
  );
  //OR U105bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U105bar (
    .O(ybar[236]),
    .I0(abar[14]),
    .I1(bbar[12])
  );
  //AND U106
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U106 (
    .O(y[235]),
    .I0(a[14]),
    .I1(b[11])
  );
  //OR U106bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U106bar (
    .O(ybar[235]),
    .I0(abar[14]),
    .I1(bbar[11])
  );
  //AND U107
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U107 (
    .O(y[234]),
    .I0(a[14]),
    .I1(b[10])
  );
  //OR U107bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U107bar (
    .O(ybar[234]),
    .I0(abar[14]),
    .I1(bbar[10])
  );
  //AND U108
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U108 (
    .O(y[233]),
    .I0(a[14]),
    .I1(b[9])
  );
  //OR U108bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U108bar (
    .O(ybar[233]),
    .I0(abar[14]),
    .I1(bbar[9])
  );
  //AND U109
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U109 (
    .O(y[232]),
    .I0(a[14]),
    .I1(b[8])
  );
  //OR U109bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U109bar (
    .O(ybar[232]),
    .I0(abar[14]),
    .I1(bbar[8])
  );
  //AND U110
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U110 (
    .O(y[231]),
    .I0(a[14]),
    .I1(b[7])
  );
  //OR U110bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U110bar (
    .O(ybar[231]),
    .I0(abar[14]),
    .I1(bbar[7])
  );
  //AND U111
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U111 (
    .O(y[230]),
    .I0(a[14]),
    .I1(b[6])
  );
  //OR U111bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U111bar (
    .O(ybar[230]),
    .I0(abar[14]),
    .I1(bbar[6])
  );
  //AND U112
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U112 (
    .O(y[22]),
    .I0(a[1]),
    .I1(b[6])
  );
  //OR U112bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U112bar (
    .O(ybar[22]),
    .I0(abar[1]),
    .I1(bbar[6])
  );
  //AND U113
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U113 (
    .O(y[229]),
    .I0(a[14]),
    .I1(b[5])
  );
  //OR U113bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U113bar (
    .O(ybar[229]),
    .I0(abar[14]),
    .I1(bbar[5])
  );
  //AND U114
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U114 (
    .O(y[228]),
    .I0(a[14]),
    .I1(b[4])
  );
  //OR U114bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U114bar (
    .O(ybar[228]),
    .I0(abar[14]),
    .I1(bbar[4])
  );
  //AND U115
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U115 (
    .O(y[227]),
    .I0(a[14]),
    .I1(b[3])
  );
  //OR U115bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U115bar (
    .O(ybar[227]),
    .I0(abar[14]),
    .I1(bbar[3])
  );
  //AND U116
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U116 (
    .O(y[226]),
    .I0(a[14]),
    .I1(b[2])
  );
  //OR U116bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U116bar (
    .O(ybar[226]),
    .I0(abar[14]),
    .I1(bbar[2])
  );
  //AND U117
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U117 (
    .O(y[225]),
    .I0(a[14]),
    .I1(b[1])
  );
  //OR U117bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U117bar (
    .O(ybar[225]),
    .I0(abar[14]),
    .I1(bbar[1])
  );
  //AND U118
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U118 (
    .O(y[224]),
    .I0(a[14]),
    .I1(b[0])
  );
  //OR U118bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U118bar (
    .O(ybar[224]),
    .I0(abar[14]),
    .I1(bbar[0])
  );
  //AND U119
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U119 (
    .O(y[223]),
    .I0(a[13]),
    .I1(b[15])
  );
  //OR U119bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U119bar (
    .O(ybar[223]),
    .I0(abar[13]),
    .I1(bbar[15])
  );
  //AND U120
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U120 (
    .O(y[222]),
    .I0(a[13]),
    .I1(b[14])
  );
  //OR U120bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U120bar (
    .O(ybar[222]),
    .I0(abar[13]),
    .I1(bbar[14])
  );
  //AND U121
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U121 (
    .O(y[221]),
    .I0(a[13]),
    .I1(b[13])
  );
  //OR U121bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U121bar (
    .O(ybar[221]),
    .I0(abar[13]),
    .I1(bbar[13])
  );
  //AND U122
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U122 (
    .O(y[220]),
    .I0(a[13]),
    .I1(b[12])
  );
  //OR U122bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U122bar (
    .O(ybar[220]),
    .I0(abar[13]),
    .I1(bbar[12])
  );
  //AND U123
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U123 (
    .O(y[21]),
    .I0(a[1]),
    .I1(b[5])
  );
  //OR U123bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U123bar (
    .O(ybar[21]),
    .I0(abar[1]),
    .I1(bbar[5])
  );
  //AND U124
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U124 (
    .O(y[219]),
    .I0(a[13]),
    .I1(b[11])
  );
  //OR U124bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U124bar (
    .O(ybar[219]),
    .I0(abar[13]),
    .I1(bbar[11])
  );
  //AND U125
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U125 (
    .O(y[218]),
    .I0(a[13]),
    .I1(b[10])
  );
  //OR U125bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U125bar (
    .O(ybar[218]),
    .I0(abar[13]),
    .I1(bbar[10])
  );
  //AND U126
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U126 (
    .O(y[217]),
    .I0(a[13]),
    .I1(b[9])
  );
  //OR U126bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U126bar (
    .O(ybar[217]),
    .I0(abar[13]),
    .I1(bbar[9])
  );
  //AND U127
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U127 (
    .O(y[216]),
    .I0(a[13]),
    .I1(b[8])
  );
  //OR U127bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U127bar (
    .O(ybar[216]),
    .I0(abar[13]),
    .I1(bbar[8])
  );
  //AND U128
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U128 (
    .O(y[215]),
    .I0(a[13]),
    .I1(b[7])
  );
  //OR U128bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U128bar (
    .O(ybar[215]),
    .I0(abar[13]),
    .I1(bbar[7])
  );
  //AND U129
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U129 (
    .O(y[214]),
    .I0(a[13]),
    .I1(b[6])
  );
  //OR U129bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U129bar (
    .O(ybar[214]),
    .I0(abar[13]),
    .I1(bbar[6])
  );
  //AND U130
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U130 (
    .O(y[213]),
    .I0(a[13]),
    .I1(b[5])
  );
  //OR U130bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U130bar (
    .O(ybar[213]),
    .I0(abar[13]),
    .I1(bbar[5])
  );
  //AND U131
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U131 (
    .O(y[212]),
    .I0(a[13]),
    .I1(b[4])
  );
  //OR U131bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U131bar (
    .O(ybar[212]),
    .I0(abar[13]),
    .I1(bbar[4])
  );
  //AND U132
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U132 (
    .O(y[211]),
    .I0(a[13]),
    .I1(b[3])
  );
  //OR U132bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U132bar (
    .O(ybar[211]),
    .I0(abar[13]),
    .I1(bbar[3])
  );
  //AND U133
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U133 (
    .O(y[210]),
    .I0(a[13]),
    .I1(b[2])
  );
  //OR U133bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U133bar (
    .O(ybar[210]),
    .I0(abar[13]),
    .I1(bbar[2])
  );
  //AND U134
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U134 (
    .O(y[20]),
    .I0(a[1]),
    .I1(b[4])
  );
  //OR U134bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U134bar (
    .O(ybar[20]),
    .I0(abar[1]),
    .I1(bbar[4])
  );
  //AND U135
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U135 (
    .O(y[209]),
    .I0(a[13]),
    .I1(b[1])
  );
  //OR U135bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U135bar (
    .O(ybar[209]),
    .I0(abar[13]),
    .I1(bbar[1])
  );
  //AND U136
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U136 (
    .O(y[208]),
    .I0(a[13]),
    .I1(b[0])
  );
  //OR U136bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U136bar (
    .O(ybar[208]),
    .I0(abar[13]),
    .I1(bbar[0])
  );
  //AND U137
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U137 (
    .O(y[207]),
    .I0(a[12]),
    .I1(b[15])
  );
  //OR U137bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U137bar (
    .O(ybar[207]),
    .I0(abar[12]),
    .I1(bbar[15])
  );
  //AND U138
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U138 (
    .O(y[206]),
    .I0(a[12]),
    .I1(b[14])
  );
  //OR U138bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U138bar (
    .O(ybar[206]),
    .I0(abar[12]),
    .I1(bbar[14])
  );
  //AND U139
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U139 (
    .O(y[205]),
    .I0(a[12]),
    .I1(b[13])
  );
  //OR U139bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U139bar (
    .O(ybar[205]),
    .I0(abar[12]),
    .I1(bbar[13])
  );
  //AND U140
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U140 (
    .O(y[204]),
    .I0(a[12]),
    .I1(b[12])
  );
  //OR U140bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U140bar (
    .O(ybar[204]),
    .I0(abar[12]),
    .I1(bbar[12])
  );
  //AND U141
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U141 (
    .O(y[203]),
    .I0(a[12]),
    .I1(b[11])
  );
  //OR U141bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U141bar (
    .O(ybar[203]),
    .I0(abar[12]),
    .I1(bbar[11])
  );
  //AND U142
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U142 (
    .O(y[202]),
    .I0(a[12]),
    .I1(b[10])
  );
  //OR U142bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U142bar (
    .O(ybar[202]),
    .I0(abar[12]),
    .I1(bbar[10])
  );
  //AND U143
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U143 (
    .O(y[201]),
    .I0(a[12]),
    .I1(b[9])
  );
  //OR U143bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U143bar (
    .O(ybar[201]),
    .I0(abar[12]),
    .I1(bbar[9])
  );
  //AND U144
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U144 (
    .O(y[200]),
    .I0(a[12]),
    .I1(b[8])
  );
  //OR U144bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U144bar (
    .O(ybar[200]),
    .I0(abar[12]),
    .I1(bbar[8])
  );
  //AND U145
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U145 (
    .O(y[1]),
    .I0(b[1]),
    .I1(a[0])
  );
  //OR U145bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U145bar (
    .O(ybar[1]),
    .I0(bbar[1]),
    .I1(abar[0])
  );
  //AND U146
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U146 (
    .O(y[19]),
    .I0(a[1]),
    .I1(b[3])
  );
  //OR U146bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U146bar (
    .O(ybar[19]),
    .I0(abar[1]),
    .I1(bbar[3])
  );
  //AND U147
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U147 (
    .O(y[199]),
    .I0(a[12]),
    .I1(b[7])
  );
  //OR U147bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U147bar (
    .O(ybar[199]),
    .I0(abar[12]),
    .I1(bbar[7])
  );
  //AND U148
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U148 (
    .O(y[198]),
    .I0(a[12]),
    .I1(b[6])
  );
  //OR U148bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U148bar (
    .O(ybar[198]),
    .I0(abar[12]),
    .I1(bbar[6])
  );
  //AND U149
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U149 (
    .O(y[197]),
    .I0(a[12]),
    .I1(b[5])
  );
  //OR U149bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U149bar (
    .O(ybar[197]),
    .I0(abar[12]),
    .I1(bbar[5])
  );
  //AND U150
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U150 (
    .O(y[196]),
    .I0(a[12]),
    .I1(b[4])
  );
  //OR U150bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U150bar (
    .O(ybar[196]),
    .I0(abar[12]),
    .I1(bbar[4])
  );
  //AND U151
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U151 (
    .O(y[195]),
    .I0(a[12]),
    .I1(b[3])
  );
  //OR U151bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U151bar (
    .O(ybar[195]),
    .I0(abar[12]),
    .I1(bbar[3])
  );
  //AND U152
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U152 (
    .O(y[194]),
    .I0(a[12]),
    .I1(b[2])
  );
  //OR U152bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U152bar (
    .O(ybar[194]),
    .I0(abar[12]),
    .I1(bbar[2])
  );
  //AND U153
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U153 (
    .O(y[193]),
    .I0(a[12]),
    .I1(b[1])
  );
  //OR U153bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U153bar (
    .O(ybar[193]),
    .I0(abar[12]),
    .I1(bbar[1])
  );
  //AND U154
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U154 (
    .O(y[192]),
    .I0(a[12]),
    .I1(b[0])
  );
  //OR U154bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U154bar (
    .O(ybar[192]),
    .I0(abar[12]),
    .I1(bbar[0])
  );
  //AND U155
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U155 (
    .O(y[191]),
    .I0(a[11]),
    .I1(b[15])
  );
  //OR U155bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U155bar (
    .O(ybar[191]),
    .I0(abar[11]),
    .I1(bbar[15])
  );
  //AND U156
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U156 (
    .O(y[190]),
    .I0(a[11]),
    .I1(b[14])
  );
  //OR U156bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U156bar (
    .O(ybar[190]),
    .I0(abar[11]),
    .I1(bbar[14])
  );
  //AND U157
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U157 (
    .O(y[18]),
    .I0(a[1]),
    .I1(b[2])
  );
  //OR U157bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U157bar (
    .O(ybar[18]),
    .I0(abar[1]),
    .I1(bbar[2])
  );
  //AND U158
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U158 (
    .O(y[189]),
    .I0(a[11]),
    .I1(b[13])
  );
  //OR U158bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U158bar (
    .O(ybar[189]),
    .I0(abar[11]),
    .I1(bbar[13])
  );
  //AND U159
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U159 (
    .O(y[188]),
    .I0(a[11]),
    .I1(b[12])
  );
  //OR U159bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U159bar (
    .O(ybar[188]),
    .I0(abar[11]),
    .I1(bbar[12])
  );
  //AND U160
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U160 (
    .O(y[187]),
    .I0(a[11]),
    .I1(b[11])
  );
  //OR U160bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U160bar (
    .O(ybar[187]),
    .I0(abar[11]),
    .I1(bbar[11])
  );
  //AND U161
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U161 (
    .O(y[186]),
    .I0(a[11]),
    .I1(b[10])
  );
  //OR U161bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U161bar (
    .O(ybar[186]),
    .I0(abar[11]),
    .I1(bbar[10])
  );
  //AND U162
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U162 (
    .O(y[185]),
    .I0(a[11]),
    .I1(b[9])
  );
  //OR U162bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U162bar (
    .O(ybar[185]),
    .I0(abar[11]),
    .I1(bbar[9])
  );
  //AND U163
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U163 (
    .O(y[184]),
    .I0(a[11]),
    .I1(b[8])
  );
  //OR U163bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U163bar (
    .O(ybar[184]),
    .I0(abar[11]),
    .I1(bbar[8])
  );
  //AND U164
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U164 (
    .O(y[183]),
    .I0(a[11]),
    .I1(b[7])
  );
  //OR U164bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U164bar (
    .O(ybar[183]),
    .I0(abar[11]),
    .I1(bbar[7])
  );
  //AND U165
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U165 (
    .O(y[182]),
    .I0(a[11]),
    .I1(b[6])
  );
  //OR U165bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U165bar (
    .O(ybar[182]),
    .I0(abar[11]),
    .I1(bbar[6])
  );
  //AND U166
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U166 (
    .O(y[181]),
    .I0(a[11]),
    .I1(b[5])
  );
  //OR U166bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U166bar (
    .O(ybar[181]),
    .I0(abar[11]),
    .I1(bbar[5])
  );
  //AND U167
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U167 (
    .O(y[180]),
    .I0(a[11]),
    .I1(b[4])
  );
  //OR U167bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U167bar (
    .O(ybar[180]),
    .I0(abar[11]),
    .I1(bbar[4])
  );
  //AND U168
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U168 (
    .O(y[17]),
    .I0(a[1]),
    .I1(b[1])
  );
  //OR U168bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U168bar (
    .O(ybar[17]),
    .I0(abar[1]),
    .I1(bbar[1])
  );
  //AND U169
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U169 (
    .O(y[179]),
    .I0(a[11]),
    .I1(b[3])
  );
  //OR U169bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U169bar (
    .O(ybar[179]),
    .I0(abar[11]),
    .I1(bbar[3])
  );
  //AND U170
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U170 (
    .O(y[178]),
    .I0(a[11]),
    .I1(b[2])
  );
  //OR U170bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U170bar (
    .O(ybar[178]),
    .I0(abar[11]),
    .I1(bbar[2])
  );
  //AND U171
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U171 (
    .O(y[177]),
    .I0(a[11]),
    .I1(b[1])
  );
  //OR U171bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U171bar (
    .O(ybar[177]),
    .I0(abar[11]),
    .I1(bbar[1])
  );
  //AND U172
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U172 (
    .O(y[176]),
    .I0(a[11]),
    .I1(b[0])
  );
  //OR U172bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U172bar (
    .O(ybar[176]),
    .I0(abar[11]),
    .I1(bbar[0])
  );
  //AND U173
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U173 (
    .O(y[175]),
    .I0(a[10]),
    .I1(b[15])
  );
  //OR U173bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U173bar (
    .O(ybar[175]),
    .I0(abar[10]),
    .I1(bbar[15])
  );
  //AND U174
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U174 (
    .O(y[174]),
    .I0(a[10]),
    .I1(b[14])
  );
  //OR U174bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U174bar (
    .O(ybar[174]),
    .I0(abar[10]),
    .I1(bbar[14])
  );
  //AND U175
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U175 (
    .O(y[173]),
    .I0(a[10]),
    .I1(b[13])
  );
  //OR U175bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U175bar (
    .O(ybar[173]),
    .I0(abar[10]),
    .I1(bbar[13])
  );
  //AND U176
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U176 (
    .O(y[172]),
    .I0(a[10]),
    .I1(b[12])
  );
  //OR U176bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U176bar (
    .O(ybar[172]),
    .I0(abar[10]),
    .I1(bbar[12])
  );
  //AND U177
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U177 (
    .O(y[171]),
    .I0(a[10]),
    .I1(b[11])
  );
  //OR U177bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U177bar (
    .O(ybar[171]),
    .I0(abar[10]),
    .I1(bbar[11])
  );
  //AND U178
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U178 (
    .O(y[170]),
    .I0(a[10]),
    .I1(b[10])
  );
  //OR U178bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U178bar (
    .O(ybar[170]),
    .I0(abar[10]),
    .I1(bbar[10])
  );
  //AND U179
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U179 (
    .O(y[16]),
    .I0(a[1]),
    .I1(b[0])
  );
  //OR U179bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U179bar (
    .O(ybar[16]),
    .I0(abar[1]),
    .I1(bbar[0])
  );
  //AND U180
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U180 (
    .O(y[169]),
    .I0(a[10]),
    .I1(b[9])
  );
  //OR U180bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U180bar (
    .O(ybar[169]),
    .I0(abar[10]),
    .I1(bbar[9])
  );
  //AND U181
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U181 (
    .O(y[168]),
    .I0(a[10]),
    .I1(b[8])
  );
  //OR U181bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U181bar (
    .O(ybar[168]),
    .I0(abar[10]),
    .I1(bbar[8])
  );
  //AND U182
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U182 (
    .O(y[167]),
    .I0(a[10]),
    .I1(b[7])
  );
  //OR U182bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U182bar (
    .O(ybar[167]),
    .I0(abar[10]),
    .I1(bbar[7])
  );
  //AND U183
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U183 (
    .O(y[166]),
    .I0(a[10]),
    .I1(b[6])
  );
  //OR U183bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U183bar (
    .O(ybar[166]),
    .I0(abar[10]),
    .I1(bbar[6])
  );
  //AND U184
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U184 (
    .O(y[165]),
    .I0(a[10]),
    .I1(b[5])
  );
  //OR U184bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U184bar (
    .O(ybar[165]),
    .I0(abar[10]),
    .I1(bbar[5])
  );
  //AND U185
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U185 (
    .O(y[164]),
    .I0(a[10]),
    .I1(b[4])
  );
  //OR U185bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U185bar (
    .O(ybar[164]),
    .I0(abar[10]),
    .I1(bbar[4])
  );
  //AND U186
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U186 (
    .O(y[163]),
    .I0(a[10]),
    .I1(b[3])
  );
  //OR U186bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U186bar (
    .O(ybar[163]),
    .I0(abar[10]),
    .I1(bbar[3])
  );
  //AND U187
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U187 (
    .O(y[162]),
    .I0(a[10]),
    .I1(b[2])
  );
  //OR U187bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U187bar (
    .O(ybar[162]),
    .I0(abar[10]),
    .I1(bbar[2])
  );
  //AND U188
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U188 (
    .O(y[161]),
    .I0(a[10]),
    .I1(b[1])
  );
  //OR U188bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U188bar (
    .O(ybar[161]),
    .I0(abar[10]),
    .I1(bbar[1])
  );
  //AND U189
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U189 (
    .O(y[160]),
    .I0(a[10]),
    .I1(b[0])
  );
  //OR U189bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U189bar (
    .O(ybar[160]),
    .I0(abar[10]),
    .I1(bbar[0])
  );
  //AND U190
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U190 (
    .O(y[15]),
    .I0(b[15]),
    .I1(a[0])
  );
  //OR U190bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U190bar (
    .O(ybar[15]),
    .I0(bbar[15]),
    .I1(abar[0])
  );
  //AND U191
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U191 (
    .O(y[159]),
    .I0(a[9]),
    .I1(b[15])
  );
  //OR U191bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U191bar (
    .O(ybar[159]),
    .I0(abar[9]),
    .I1(bbar[15])
  );
  //AND U192
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U192 (
    .O(y[158]),
    .I0(a[9]),
    .I1(b[14])
  );
  //OR U192bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U192bar (
    .O(ybar[158]),
    .I0(abar[9]),
    .I1(bbar[14])
  );
  //AND U193
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U193 (
    .O(y[157]),
    .I0(a[9]),
    .I1(b[13])
  );
  //OR U193bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U193bar (
    .O(ybar[157]),
    .I0(abar[9]),
    .I1(bbar[13])
  );
  //AND U194
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U194 (
    .O(y[156]),
    .I0(a[9]),
    .I1(b[12])
  );
  //OR U194bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U194bar (
    .O(ybar[156]),
    .I0(abar[9]),
    .I1(bbar[12])
  );
  //AND U195
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U195 (
    .O(y[155]),
    .I0(a[9]),
    .I1(b[11])
  );
  //OR U195bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U195bar (
    .O(ybar[155]),
    .I0(abar[9]),
    .I1(bbar[11])
  );
  //AND U196
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U196 (
    .O(y[154]),
    .I0(a[9]),
    .I1(b[10])
  );
  //OR U196bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U196bar (
    .O(ybar[154]),
    .I0(abar[9]),
    .I1(bbar[10])
  );
  //AND U197
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U197 (
    .O(y[153]),
    .I0(a[9]),
    .I1(b[9])
  );
  //OR U197bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U197bar (
    .O(ybar[153]),
    .I0(abar[9]),
    .I1(bbar[9])
  );
  //AND U198
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U198 (
    .O(y[152]),
    .I0(a[9]),
    .I1(b[8])
  );
  //OR U198bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U198bar (
    .O(ybar[152]),
    .I0(abar[9]),
    .I1(bbar[8])
  );
  //AND U199
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U199 (
    .O(y[151]),
    .I0(a[9]),
    .I1(b[7])
  );
  //OR U199bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U199bar (
    .O(ybar[151]),
    .I0(abar[9]),
    .I1(bbar[7])
  );
  //AND U200
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U200 (
    .O(y[150]),
    .I0(a[9]),
    .I1(b[6])
  );
  //OR U200bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U200bar (
    .O(ybar[150]),
    .I0(abar[9]),
    .I1(bbar[6])
  );
  //AND U201
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U201 (
    .O(y[14]),
    .I0(b[14]),
    .I1(a[0])
  );
  //OR U201bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U201bar (
    .O(ybar[14]),
    .I0(bbar[14]),
    .I1(abar[0])
  );
  //AND U202
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U202 (
    .O(y[149]),
    .I0(a[9]),
    .I1(b[5])
  );
  //OR U202bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U202bar (
    .O(ybar[149]),
    .I0(abar[9]),
    .I1(bbar[5])
  );
  //AND U203
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U203 (
    .O(y[148]),
    .I0(a[9]),
    .I1(b[4])
  );
  //OR U203bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U203bar (
    .O(ybar[148]),
    .I0(abar[9]),
    .I1(bbar[4])
  );
  //AND U204
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U204 (
    .O(y[147]),
    .I0(a[9]),
    .I1(b[3])
  );
  //OR U204bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U204bar (
    .O(ybar[147]),
    .I0(abar[9]),
    .I1(bbar[3])
  );
  //AND U205
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U205 (
    .O(y[146]),
    .I0(a[9]),
    .I1(b[2])
  );
  //OR U205bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U205bar (
    .O(ybar[146]),
    .I0(abar[9]),
    .I1(bbar[2])
  );
  //AND U206
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U206 (
    .O(y[145]),
    .I0(a[9]),
    .I1(b[1])
  );
  //OR U206bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U206bar (
    .O(ybar[145]),
    .I0(abar[9]),
    .I1(bbar[1])
  );
  //AND U207
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U207 (
    .O(y[144]),
    .I0(a[9]),
    .I1(b[0])
  );
  //OR U207bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U207bar (
    .O(ybar[144]),
    .I0(abar[9]),
    .I1(bbar[0])
  );
  //AND U208
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U208 (
    .O(y[143]),
    .I0(a[8]),
    .I1(b[15])
  );
  //OR U208bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U208bar (
    .O(ybar[143]),
    .I0(abar[8]),
    .I1(bbar[15])
  );
  //AND U209
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U209 (
    .O(y[142]),
    .I0(a[8]),
    .I1(b[14])
  );
  //OR U209bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U209bar (
    .O(ybar[142]),
    .I0(abar[8]),
    .I1(bbar[14])
  );
  //AND U210
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U210 (
    .O(y[141]),
    .I0(a[8]),
    .I1(b[13])
  );
  //OR U210bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U210bar (
    .O(ybar[141]),
    .I0(abar[8]),
    .I1(bbar[13])
  );
  //AND U211
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U211 (
    .O(y[140]),
    .I0(a[8]),
    .I1(b[12])
  );
  //OR U211bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U211bar (
    .O(ybar[140]),
    .I0(abar[8]),
    .I1(bbar[12])
  );
  //AND U212
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U212 (
    .O(y[13]),
    .I0(b[13]),
    .I1(a[0])
  );
  //OR U212bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U212bar (
    .O(ybar[13]),
    .I0(bbar[13]),
    .I1(abar[0])
  );
  //AND U213
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U213 (
    .O(y[139]),
    .I0(a[8]),
    .I1(b[11])
  );
  //OR U213bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U213bar (
    .O(ybar[139]),
    .I0(abar[8]),
    .I1(bbar[11])
  );
  //AND U214
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U214 (
    .O(y[138]),
    .I0(a[8]),
    .I1(b[10])
  );
  //OR U214bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U214bar (
    .O(ybar[138]),
    .I0(abar[8]),
    .I1(bbar[10])
  );
  //AND U215
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U215 (
    .O(y[137]),
    .I0(a[8]),
    .I1(b[9])
  );
  //OR U215bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U215bar (
    .O(ybar[137]),
    .I0(abar[8]),
    .I1(bbar[9])
  );
  //AND U216
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U216 (
    .O(y[136]),
    .I0(a[8]),
    .I1(b[8])
  );
  //OR U216bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U216bar (
    .O(ybar[136]),
    .I0(abar[8]),
    .I1(bbar[8])
  );
  //AND U217
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U217 (
    .O(y[135]),
    .I0(a[8]),
    .I1(b[7])
  );
  //OR U217bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U217bar (
    .O(ybar[135]),
    .I0(abar[8]),
    .I1(bbar[7])
  );
  //AND U218
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U218 (
    .O(y[134]),
    .I0(a[8]),
    .I1(b[6])
  );
  //OR U218bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U218bar (
    .O(ybar[134]),
    .I0(abar[8]),
    .I1(bbar[6])
  );
  //AND U219
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U219 (
    .O(y[133]),
    .I0(a[8]),
    .I1(b[5])
  );
  //OR U219bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U219bar (
    .O(ybar[133]),
    .I0(abar[8]),
    .I1(bbar[5])
  );
  //AND U220
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U220 (
    .O(y[132]),
    .I0(a[8]),
    .I1(b[4])
  );
  //OR U220bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U220bar (
    .O(ybar[132]),
    .I0(abar[8]),
    .I1(bbar[4])
  );
  //AND U221
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U221 (
    .O(y[131]),
    .I0(a[8]),
    .I1(b[3])
  );
  //OR U221bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U221bar (
    .O(ybar[131]),
    .I0(abar[8]),
    .I1(bbar[3])
  );
  //AND U222
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U222 (
    .O(y[130]),
    .I0(a[8]),
    .I1(b[2])
  );
  //OR U222bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U222bar (
    .O(ybar[130]),
    .I0(abar[8]),
    .I1(bbar[2])
  );
  //AND U223
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U223 (
    .O(y[12]),
    .I0(b[12]),
    .I1(a[0])
  );
  //OR U223bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U223bar (
    .O(ybar[12]),
    .I0(bbar[12]),
    .I1(abar[0])
  );
  //AND U224
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U224 (
    .O(y[129]),
    .I0(a[8]),
    .I1(b[1])
  );
  //OR U224bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U224bar (
    .O(ybar[129]),
    .I0(abar[8]),
    .I1(bbar[1])
  );
  //AND U225
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U225 (
    .O(y[128]),
    .I0(a[8]),
    .I1(b[0])
  );
  //OR U225bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U225bar (
    .O(ybar[128]),
    .I0(abar[8]),
    .I1(bbar[0])
  );
  //AND U226
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U226 (
    .O(y[127]),
    .I0(a[7]),
    .I1(b[15])
  );
  //OR U226bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U226bar (
    .O(ybar[127]),
    .I0(abar[7]),
    .I1(bbar[15])
  );
  //AND U227
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U227 (
    .O(y[126]),
    .I0(a[7]),
    .I1(b[14])
  );
  //OR U227bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U227bar (
    .O(ybar[126]),
    .I0(abar[7]),
    .I1(bbar[14])
  );
  //AND U228
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U228 (
    .O(y[125]),
    .I0(a[7]),
    .I1(b[13])
  );
  //OR U228bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U228bar (
    .O(ybar[125]),
    .I0(abar[7]),
    .I1(bbar[13])
  );
  //AND U229
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U229 (
    .O(y[124]),
    .I0(a[7]),
    .I1(b[12])
  );
  //OR U229bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U229bar (
    .O(ybar[124]),
    .I0(abar[7]),
    .I1(bbar[12])
  );
  //AND U230
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U230 (
    .O(y[123]),
    .I0(a[7]),
    .I1(b[11])
  );
  //OR U230bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U230bar (
    .O(ybar[123]),
    .I0(abar[7]),
    .I1(bbar[11])
  );
  //AND U231
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U231 (
    .O(y[122]),
    .I0(a[7]),
    .I1(b[10])
  );
  //OR U231bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U231bar (
    .O(ybar[122]),
    .I0(abar[7]),
    .I1(bbar[10])
  );
  //AND U232
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U232 (
    .O(y[121]),
    .I0(a[7]),
    .I1(b[9])
  );
  //OR U232bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U232bar (
    .O(ybar[121]),
    .I0(abar[7]),
    .I1(bbar[9])
  );
  //AND U233
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U233 (
    .O(y[120]),
    .I0(a[7]),
    .I1(b[8])
  );
  //OR U233bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U233bar (
    .O(ybar[120]),
    .I0(abar[7]),
    .I1(bbar[8])
  );
  //AND U234
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U234 (
    .O(y[11]),
    .I0(b[11]),
    .I1(a[0])
  );
  //OR U234bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U234bar (
    .O(ybar[11]),
    .I0(bbar[11]),
    .I1(abar[0])
  );
  //AND U235
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U235 (
    .O(y[119]),
    .I0(a[7]),
    .I1(b[7])
  );
  //OR U235bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U235bar (
    .O(ybar[119]),
    .I0(abar[7]),
    .I1(bbar[7])
  );
  //AND U236
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U236 (
    .O(y[118]),
    .I0(a[7]),
    .I1(b[6])
  );
  //OR U236bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U236bar (
    .O(ybar[118]),
    .I0(abar[7]),
    .I1(bbar[6])
  );
  //AND U237
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U237 (
    .O(y[117]),
    .I0(a[7]),
    .I1(b[5])
  );
  //OR U237bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U237bar (
    .O(ybar[117]),
    .I0(abar[7]),
    .I1(bbar[5])
  );
  //AND U238
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U238 (
    .O(y[116]),
    .I0(a[7]),
    .I1(b[4])
  );
  //OR U238bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U238bar (
    .O(ybar[116]),
    .I0(abar[7]),
    .I1(bbar[4])
  );
  //AND U239
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U239 (
    .O(y[115]),
    .I0(a[7]),
    .I1(b[3])
  );
  //OR U239bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U239bar (
    .O(ybar[115]),
    .I0(abar[7]),
    .I1(bbar[3])
  );
  //AND U240
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U240 (
    .O(y[114]),
    .I0(a[7]),
    .I1(b[2])
  );
  //OR U240bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U240bar (
    .O(ybar[114]),
    .I0(abar[7]),
    .I1(bbar[2])
  );
  //AND U241
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U241 (
    .O(y[113]),
    .I0(a[7]),
    .I1(b[1])
  );
  //OR U241bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U241bar (
    .O(ybar[113]),
    .I0(abar[7]),
    .I1(bbar[1])
  );
  //AND U242
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U242 (
    .O(y[112]),
    .I0(a[7]),
    .I1(b[0])
  );
  //OR U242bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U242bar (
    .O(ybar[112]),
    .I0(abar[7]),
    .I1(bbar[0])
  );
  //AND U243
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U243 (
    .O(y[111]),
    .I0(b[15]),
    .I1(a[6])
  );
  //OR U243bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U243bar (
    .O(ybar[111]),
    .I0(bbar[15]),
    .I1(abar[6])
  );
  //AND U244
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U244 (
    .O(y[110]),
    .I0(b[14]),
    .I1(a[6])
  );
  //OR U244bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U244bar (
    .O(ybar[110]),
    .I0(bbar[14]),
    .I1(abar[6])
  );
  //AND U245
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U245 (
    .O(y[10]),
    .I0(b[10]),
    .I1(a[0])
  );
  //OR U245bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U245bar (
    .O(ybar[10]),
    .I0(bbar[10]),
    .I1(abar[0])
  );
  //AND U246
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U246 (
    .O(y[109]),
    .I0(b[13]),
    .I1(a[6])
  );
  //OR U246bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U246bar (
    .O(ybar[109]),
    .I0(bbar[13]),
    .I1(abar[6])
  );
  //AND U247
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U247 (
    .O(y[108]),
    .I0(b[12]),
    .I1(a[6])
  );
  //OR U247bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U247bar (
    .O(ybar[108]),
    .I0(bbar[12]),
    .I1(abar[6])
  );
  //AND U248
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U248 (
    .O(y[107]),
    .I0(b[11]),
    .I1(a[6])
  );
  //OR U248bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U248bar (
    .O(ybar[107]),
    .I0(bbar[11]),
    .I1(abar[6])
  );
  //AND U249
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U249 (
    .O(y[106]),
    .I0(b[10]),
    .I1(a[6])
  );
  //OR U249bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U249bar (
    .O(ybar[106]),
    .I0(bbar[10]),
    .I1(abar[6])
  );
  //AND U250
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U250 (
    .O(y[105]),
    .I0(a[6]),
    .I1(b[9])
  );
  //OR U250bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U250bar (
    .O(ybar[105]),
    .I0(abar[6]),
    .I1(bbar[9])
  );
  //AND U251
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U251 (
    .O(y[104]),
    .I0(b[8]),
    .I1(a[6])
  );
  //OR U251bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U251bar (
    .O(ybar[104]),
    .I0(bbar[8]),
    .I1(abar[6])
  );
  //AND U252
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U252 (
    .O(y[103]),
    .I0(b[7]),
    .I1(a[6])
  );
  //OR U252bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U252bar (
    .O(ybar[103]),
    .I0(bbar[7]),
    .I1(abar[6])
  );
  //AND U253
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U253 (
    .O(y[102]),
    .I0(b[6]),
    .I1(a[6])
  );
  //OR U253bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U253bar (
    .O(ybar[102]),
    .I0(bbar[6]),
    .I1(abar[6])
  );
  //AND U254
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U254 (
    .O(y[101]),
    .I0(b[5]),
    .I1(a[6])
  );
  //OR U254bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U254bar (
    .O(ybar[101]),
    .I0(bbar[5]),
    .I1(abar[6])
  );
  //AND U255
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U255 (
    .O(y[100]),
    .I0(b[4]),
    .I1(a[6])
  );
  //OR U255bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U255bar (
    .O(ybar[100]),
    .I0(bbar[4]),
    .I1(abar[6])
  );
  //AND U256
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U256 (
    .O(y[0]),
    .I0(b[0]),
    .I1(a[0])
  );
  //OR U256bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U256bar (
    .O(ybar[0]),
    .I0(bbar[0]),
    .I1(abar[0])
  );
endmodule

module decode_8 ( in, out );

  input wire [7:0] in;
//input_done

  output wire [255:0] out;
//output_done

  wire [15:0] level1;
  wire [31:0] level2;
//wire_done

  CD2_32 cd_l1_1 ( .a(in[1]), .b(in[0]), .y(level1[3:0]) );
  CD2_31 cd_l1_2 ( .a(in[3]), .b(in[2]), .y(level1[7:4]) );
  CD2_30 cd_l1_3 ( .a(in[5]), .b(in[4]), .y(level1[11:8]) );
  CD2_29 cd_l1_4 ( .a(in[7]), .b(in[6]), .y(level1[15:12]) );
  CD4_16 cd_l2_1 ( .a(level1[7:4]), .b(level1[3:0]), .y(level2[15:0]) );
  CD4_15 cd_l2_2 ( .a(level1[15:12]), .b(level1[11:8]), .y(level2[31:16]) );
  CD16_8 cd_l3 ( .a(level2[31:16]), .b(level2[15:0]), .y(out) );
endmodule

module encode_8 ( in, out );

  input wire [255:0] in;
  wire [255:0] inbar;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
  assign inbar[8] = ~in[8];
  assign inbar[9] = ~in[9];
  assign inbar[10] = ~in[10];
  assign inbar[11] = ~in[11];
  assign inbar[12] = ~in[12];
  assign inbar[13] = ~in[13];
  assign inbar[14] = ~in[14];
  assign inbar[15] = ~in[15];
  assign inbar[16] = ~in[16];
  assign inbar[17] = ~in[17];
  assign inbar[18] = ~in[18];
  assign inbar[19] = ~in[19];
  assign inbar[20] = ~in[20];
  assign inbar[21] = ~in[21];
  assign inbar[22] = ~in[22];
  assign inbar[23] = ~in[23];
  assign inbar[24] = ~in[24];
  assign inbar[25] = ~in[25];
  assign inbar[26] = ~in[26];
  assign inbar[27] = ~in[27];
  assign inbar[28] = ~in[28];
  assign inbar[29] = ~in[29];
  assign inbar[30] = ~in[30];
  assign inbar[31] = ~in[31];
  assign inbar[32] = ~in[32];
  assign inbar[33] = ~in[33];
  assign inbar[34] = ~in[34];
  assign inbar[35] = ~in[35];
  assign inbar[36] = ~in[36];
  assign inbar[37] = ~in[37];
  assign inbar[38] = ~in[38];
  assign inbar[39] = ~in[39];
  assign inbar[40] = ~in[40];
  assign inbar[41] = ~in[41];
  assign inbar[42] = ~in[42];
  assign inbar[43] = ~in[43];
  assign inbar[44] = ~in[44];
  assign inbar[45] = ~in[45];
  assign inbar[46] = ~in[46];
  assign inbar[47] = ~in[47];
  assign inbar[48] = ~in[48];
  assign inbar[49] = ~in[49];
  assign inbar[50] = ~in[50];
  assign inbar[51] = ~in[51];
  assign inbar[52] = ~in[52];
  assign inbar[53] = ~in[53];
  assign inbar[54] = ~in[54];
  assign inbar[55] = ~in[55];
  assign inbar[56] = ~in[56];
  assign inbar[57] = ~in[57];
  assign inbar[58] = ~in[58];
  assign inbar[59] = ~in[59];
  assign inbar[60] = ~in[60];
  assign inbar[61] = ~in[61];
  assign inbar[62] = ~in[62];
  assign inbar[63] = ~in[63];
  assign inbar[64] = ~in[64];
  assign inbar[65] = ~in[65];
  assign inbar[66] = ~in[66];
  assign inbar[67] = ~in[67];
  assign inbar[68] = ~in[68];
  assign inbar[69] = ~in[69];
  assign inbar[70] = ~in[70];
  assign inbar[71] = ~in[71];
  assign inbar[72] = ~in[72];
  assign inbar[73] = ~in[73];
  assign inbar[74] = ~in[74];
  assign inbar[75] = ~in[75];
  assign inbar[76] = ~in[76];
  assign inbar[77] = ~in[77];
  assign inbar[78] = ~in[78];
  assign inbar[79] = ~in[79];
  assign inbar[80] = ~in[80];
  assign inbar[81] = ~in[81];
  assign inbar[82] = ~in[82];
  assign inbar[83] = ~in[83];
  assign inbar[84] = ~in[84];
  assign inbar[85] = ~in[85];
  assign inbar[86] = ~in[86];
  assign inbar[87] = ~in[87];
  assign inbar[88] = ~in[88];
  assign inbar[89] = ~in[89];
  assign inbar[90] = ~in[90];
  assign inbar[91] = ~in[91];
  assign inbar[92] = ~in[92];
  assign inbar[93] = ~in[93];
  assign inbar[94] = ~in[94];
  assign inbar[95] = ~in[95];
  assign inbar[96] = ~in[96];
  assign inbar[97] = ~in[97];
  assign inbar[98] = ~in[98];
  assign inbar[99] = ~in[99];
  assign inbar[100] = ~in[100];
  assign inbar[101] = ~in[101];
  assign inbar[102] = ~in[102];
  assign inbar[103] = ~in[103];
  assign inbar[104] = ~in[104];
  assign inbar[105] = ~in[105];
  assign inbar[106] = ~in[106];
  assign inbar[107] = ~in[107];
  assign inbar[108] = ~in[108];
  assign inbar[109] = ~in[109];
  assign inbar[110] = ~in[110];
  assign inbar[111] = ~in[111];
  assign inbar[112] = ~in[112];
  assign inbar[113] = ~in[113];
  assign inbar[114] = ~in[114];
  assign inbar[115] = ~in[115];
  assign inbar[116] = ~in[116];
  assign inbar[117] = ~in[117];
  assign inbar[118] = ~in[118];
  assign inbar[119] = ~in[119];
  assign inbar[120] = ~in[120];
  assign inbar[121] = ~in[121];
  assign inbar[122] = ~in[122];
  assign inbar[123] = ~in[123];
  assign inbar[124] = ~in[124];
  assign inbar[125] = ~in[125];
  assign inbar[126] = ~in[126];
  assign inbar[127] = ~in[127];
  assign inbar[128] = ~in[128];
  assign inbar[129] = ~in[129];
  assign inbar[130] = ~in[130];
  assign inbar[131] = ~in[131];
  assign inbar[132] = ~in[132];
  assign inbar[133] = ~in[133];
  assign inbar[134] = ~in[134];
  assign inbar[135] = ~in[135];
  assign inbar[136] = ~in[136];
  assign inbar[137] = ~in[137];
  assign inbar[138] = ~in[138];
  assign inbar[139] = ~in[139];
  assign inbar[140] = ~in[140];
  assign inbar[141] = ~in[141];
  assign inbar[142] = ~in[142];
  assign inbar[143] = ~in[143];
  assign inbar[144] = ~in[144];
  assign inbar[145] = ~in[145];
  assign inbar[146] = ~in[146];
  assign inbar[147] = ~in[147];
  assign inbar[148] = ~in[148];
  assign inbar[149] = ~in[149];
  assign inbar[150] = ~in[150];
  assign inbar[151] = ~in[151];
  assign inbar[152] = ~in[152];
  assign inbar[153] = ~in[153];
  assign inbar[154] = ~in[154];
  assign inbar[155] = ~in[155];
  assign inbar[156] = ~in[156];
  assign inbar[157] = ~in[157];
  assign inbar[158] = ~in[158];
  assign inbar[159] = ~in[159];
  assign inbar[160] = ~in[160];
  assign inbar[161] = ~in[161];
  assign inbar[162] = ~in[162];
  assign inbar[163] = ~in[163];
  assign inbar[164] = ~in[164];
  assign inbar[165] = ~in[165];
  assign inbar[166] = ~in[166];
  assign inbar[167] = ~in[167];
  assign inbar[168] = ~in[168];
  assign inbar[169] = ~in[169];
  assign inbar[170] = ~in[170];
  assign inbar[171] = ~in[171];
  assign inbar[172] = ~in[172];
  assign inbar[173] = ~in[173];
  assign inbar[174] = ~in[174];
  assign inbar[175] = ~in[175];
  assign inbar[176] = ~in[176];
  assign inbar[177] = ~in[177];
  assign inbar[178] = ~in[178];
  assign inbar[179] = ~in[179];
  assign inbar[180] = ~in[180];
  assign inbar[181] = ~in[181];
  assign inbar[182] = ~in[182];
  assign inbar[183] = ~in[183];
  assign inbar[184] = ~in[184];
  assign inbar[185] = ~in[185];
  assign inbar[186] = ~in[186];
  assign inbar[187] = ~in[187];
  assign inbar[188] = ~in[188];
  assign inbar[189] = ~in[189];
  assign inbar[190] = ~in[190];
  assign inbar[191] = ~in[191];
  assign inbar[192] = ~in[192];
  assign inbar[193] = ~in[193];
  assign inbar[194] = ~in[194];
  assign inbar[195] = ~in[195];
  assign inbar[196] = ~in[196];
  assign inbar[197] = ~in[197];
  assign inbar[198] = ~in[198];
  assign inbar[199] = ~in[199];
  assign inbar[200] = ~in[200];
  assign inbar[201] = ~in[201];
  assign inbar[202] = ~in[202];
  assign inbar[203] = ~in[203];
  assign inbar[204] = ~in[204];
  assign inbar[205] = ~in[205];
  assign inbar[206] = ~in[206];
  assign inbar[207] = ~in[207];
  assign inbar[208] = ~in[208];
  assign inbar[209] = ~in[209];
  assign inbar[210] = ~in[210];
  assign inbar[211] = ~in[211];
  assign inbar[212] = ~in[212];
  assign inbar[213] = ~in[213];
  assign inbar[214] = ~in[214];
  assign inbar[215] = ~in[215];
  assign inbar[216] = ~in[216];
  assign inbar[217] = ~in[217];
  assign inbar[218] = ~in[218];
  assign inbar[219] = ~in[219];
  assign inbar[220] = ~in[220];
  assign inbar[221] = ~in[221];
  assign inbar[222] = ~in[222];
  assign inbar[223] = ~in[223];
  assign inbar[224] = ~in[224];
  assign inbar[225] = ~in[225];
  assign inbar[226] = ~in[226];
  assign inbar[227] = ~in[227];
  assign inbar[228] = ~in[228];
  assign inbar[229] = ~in[229];
  assign inbar[230] = ~in[230];
  assign inbar[231] = ~in[231];
  assign inbar[232] = ~in[232];
  assign inbar[233] = ~in[233];
  assign inbar[234] = ~in[234];
  assign inbar[235] = ~in[235];
  assign inbar[236] = ~in[236];
  assign inbar[237] = ~in[237];
  assign inbar[238] = ~in[238];
  assign inbar[239] = ~in[239];
  assign inbar[240] = ~in[240];
  assign inbar[241] = ~in[241];
  assign inbar[242] = ~in[242];
  assign inbar[243] = ~in[243];
  assign inbar[244] = ~in[244];
  assign inbar[245] = ~in[245];
  assign inbar[246] = ~in[246];
  assign inbar[247] = ~in[247];
  assign inbar[248] = ~in[248];
  assign inbar[249] = ~in[249];
  assign inbar[250] = ~in[250];
  assign inbar[251] = ~in[251];
  assign inbar[252] = ~in[252];
  assign inbar[253] = ~in[253];
  assign inbar[254] = ~in[254];
  assign inbar[255] = ~in[255];
//input_done

  output wire [7:0] out;
  wire [7:0] outbar;
//output_done

  wire in_81;
  wire in_80;
  wire in_79;
  wire in_78;
  wire in_77;
  wire in_76;
  wire in_75;
  wire in_74;
  wire in_73;
  wire in_72;
  wire in_71;
  wire in_70;
  wire in_69;
  wire in_68;
  wire in_67;
  wire in_66;
  wire in_65;
  wire in_64;
  wire in_63;
  wire in_62;
  wire in_61;
  wire in_60;
  wire in_59;
  wire in_58;
  wire in_57;
  wire in_56;
  wire in_55;
  wire in_54;
  wire in_53;
  wire in_52;
  wire in_51;
  wire in_50;
  wire in_49;
  wire in_48;
  wire in_47;
  wire in_46;
  wire in_45;
  wire in_44;
  wire in_43;
  wire in_42;
  wire in_41;
  wire in_40;
  wire in_39;
  wire in_38;
  wire in_37;
  wire in_36;
  wire in_35;
  wire in_34;
  wire in_33;
  wire in_32;
  wire in_31;
  wire in_30;
  wire in_29;
  wire in_28;
  wire in_27;
  wire in_26;
  wire in_25;
  wire in_24;
  wire in_23;
  wire in_22;
  wire in_21;
  wire in_20;
  wire in_19;
  wire in_18;
  wire in_17;
  wire in_16;
  wire in_15;
  wire in_14;
  wire in_13;
  wire in_12;
  wire in_11;
  wire in_10;
  wire in_9;
  wire in_8;
  wire in_7;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_3;
  wire in_2;
  wire in_1;
  wire in_0;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire in_81bar;
  wire in_80bar;
  wire in_79bar;
  wire in_78bar;
  wire in_77bar;
  wire in_76bar;
  wire in_75bar;
  wire in_74bar;
  wire in_73bar;
  wire in_72bar;
  wire in_71bar;
  wire in_70bar;
  wire in_69bar;
  wire in_68bar;
  wire in_67bar;
  wire in_66bar;
  wire in_65bar;
  wire in_64bar;
  wire in_63bar;
  wire in_62bar;
  wire in_61bar;
  wire in_60bar;
  wire in_59bar;
  wire in_58bar;
  wire in_57bar;
  wire in_56bar;
  wire in_55bar;
  wire in_54bar;
  wire in_53bar;
  wire in_52bar;
  wire in_51bar;
  wire in_50bar;
  wire in_49bar;
  wire in_48bar;
  wire in_47bar;
  wire in_46bar;
  wire in_45bar;
  wire in_44bar;
  wire in_43bar;
  wire in_42bar;
  wire in_41bar;
  wire in_40bar;
  wire in_39bar;
  wire in_38bar;
  wire in_37bar;
  wire in_36bar;
  wire in_35bar;
  wire in_34bar;
  wire in_33bar;
  wire in_32bar;
  wire in_31bar;
  wire in_30bar;
  wire in_29bar;
  wire in_28bar;
  wire in_27bar;
  wire in_26bar;
  wire in_25bar;
  wire in_24bar;
  wire in_23bar;
  wire in_22bar;
  wire in_21bar;
  wire in_20bar;
  wire in_19bar;
  wire in_18bar;
  wire in_17bar;
  wire in_16bar;
  wire in_15bar;
  wire in_14bar;
  wire in_13bar;
  wire in_12bar;
  wire in_11bar;
  wire in_10bar;
  wire in_9bar;
  wire in_8bar;
  wire in_7bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_3bar;
  wire in_2bar;
  wire in_1bar;
  wire in_0bar;
  wire n487bar;
  wire n488bar;
  wire n489bar;
  wire n490bar;
  wire n491bar;
  wire n492bar;
  wire n493bar;
  wire n494bar;
  wire n495bar;
  wire n496bar;
  wire n497bar;
  wire n498bar;
  wire n499bar;
  wire n500bar;
  wire n501bar;
  wire n502bar;
  wire n503bar;
  wire n504bar;
  wire n505bar;
  wire n506bar;
  wire n507bar;
  wire n508bar;
  wire n509bar;
  wire n510bar;
  wire n511bar;
  wire n512bar;
  wire n513bar;
  wire n514bar;
  wire n515bar;
  wire n516bar;
  wire n517bar;
  wire n518bar;
  wire n519bar;
  wire n520bar;
  wire n521bar;
  wire n522bar;
  wire n523bar;
  wire n524bar;
  wire n525bar;
  wire n526bar;
  wire n527bar;
  wire n528bar;
  wire n529bar;
  wire n530bar;
  wire n531bar;
  wire n532bar;
  wire n533bar;
  wire n534bar;
  wire n535bar;
  wire n536bar;
  wire n537bar;
  wire n538bar;
  wire n539bar;
  wire n540bar;
  wire n541bar;
  wire n542bar;
  wire n543bar;
  wire n544bar;
  wire n545bar;
  wire n546bar;
  wire n547bar;
  wire n548bar;
  wire n549bar;
  wire n550bar;
  wire n551bar;
  wire n552bar;
  wire n553bar;
  wire n554bar;
  wire n555bar;
  wire n556bar;
  wire n557bar;
  wire n558bar;
  wire n559bar;
  wire n560bar;
  wire n561bar;
  wire n562bar;
  wire n563bar;
  wire n564bar;
  wire n565bar;
  wire n566bar;
  wire n567bar;
  wire n568bar;
  wire n569bar;
  wire n570bar;
  wire n571bar;
  wire n572bar;
  wire n573bar;
  wire n574bar;
  wire n575bar;
  wire n576bar;
  wire n577bar;
  wire n578bar;
  wire n579bar;
  wire n580bar;
  wire n581bar;
  wire n582bar;
  wire n583bar;
  wire n584bar;
  wire n585bar;
  wire n586bar;
  wire n587bar;
  wire n588bar;
  wire n589bar;
  wire n590bar;
  wire n591bar;
  wire n592bar;
  wire n593bar;
  wire n594bar;
  wire n595bar;
  wire n596bar;
  wire n597bar;
  wire n598bar;
  wire n599bar;
  wire n600bar;
  wire n601bar;
  wire n602bar;
  wire n603bar;
  wire n604bar;
  wire n605bar;
  wire n606bar;
  wire n607bar;
  wire n608bar;
  wire n609bar;
  wire n610bar;
  wire n611bar;
  wire n612bar;
  wire n613bar;
  wire n614bar;
  wire n615bar;
  wire n616bar;
  wire n617bar;
  wire n618bar;
  wire n619bar;
  wire n620bar;
  wire n621bar;
  wire n622bar;
  wire n623bar;
  wire n624bar;
  wire n625bar;
  wire n626bar;
  wire n627bar;
  wire n628bar;
  wire n629bar;
  wire n630bar;
  wire n631bar;
  wire n632bar;
  wire n633bar;
  wire n634bar;
  wire n635bar;
  wire n636bar;
  wire n637bar;
  wire n638bar;
  wire n639bar;
  wire n640bar;
  wire n641bar;
  wire n642bar;
  wire n643bar;
  wire n644bar;
  wire n645bar;
  wire n646bar;
  wire n647bar;
  wire n648bar;
  wire n649bar;
  wire n650bar;
  wire n651bar;
  wire n652bar;
  wire n653bar;
  wire n654bar;
  wire n655bar;
  wire n656bar;
  wire n657bar;
  wire n658bar;
  wire n659bar;
  wire n660bar;
  wire n661bar;
  wire n662bar;
  wire n663bar;
  wire n664bar;
  wire n665bar;
  wire n666bar;
  wire n667bar;
  wire n668bar;
  wire n669bar;
  wire n670bar;
  wire n671bar;
  wire n672bar;
  wire n673bar;
  wire n674bar;
  wire n675bar;
  wire n676bar;
  wire n677bar;
  wire n678bar;
  wire n679bar;
  wire n680bar;
  wire n681bar;
  wire n682bar;
  wire n683bar;
  wire n684bar;
  wire n685bar;
  wire n686bar;
  wire n687bar;
  wire n688bar;
  wire n689bar;
  wire n690bar;
  wire n691bar;
  wire n692bar;
  wire n693bar;
  wire n694bar;
  wire n695bar;
  wire n696bar;
  wire n697bar;
  wire n698bar;
  wire n699bar;
  wire n700bar;
  wire n701bar;
  wire n702bar;
  wire n703bar;
  wire n704bar;
  wire n705bar;
  wire n706bar;
  wire n707bar;
  wire n708bar;
  wire n709bar;
  wire n710bar;
  wire n711bar;
  wire n712bar;
  wire n713bar;
  wire n714bar;
  wire n715bar;
  wire n716bar;
  wire n717bar;
  wire n718bar;
  wire n719bar;
  wire n720bar;
  wire n721bar;
  wire n722bar;
  wire n723bar;
  wire n724bar;
  wire n725bar;
  wire n726bar;
  wire n727bar;
  wire n728bar;
  wire n729bar;
  wire n730bar;
  wire n731bar;
  wire n732bar;
  wire n733bar;
  wire n734bar;
  wire n735bar;
  wire n736bar;
  wire n737bar;
  wire n738bar;
  wire n739bar;
  wire n740bar;
  wire n741bar;
  wire n742bar;
  wire n743bar;
  wire n744bar;
  wire n745bar;
  wire n746bar;
  wire n747bar;
  wire n748bar;
  wire n749bar;
  wire n750bar;
  wire n751bar;
  wire n752bar;
  wire n753bar;
  wire n754bar;
  wire n755bar;
  wire n756bar;
  wire n757bar;
  wire n758bar;
  wire n759bar;
  wire n760bar;
  wire n761bar;
  wire n762bar;
  wire n763bar;
  wire n764bar;
  wire n765bar;
  wire n766bar;
  wire n767bar;
  wire n768bar;
  wire n769bar;
  wire n770bar;
  wire n771bar;
  wire n772bar;
  wire n773bar;
  wire n774bar;
  wire n775bar;
  wire n776bar;
  wire n777bar;
  wire n778bar;
  wire n779bar;
  wire n780bar;
  wire n781bar;
  wire n782bar;
  wire n783bar;
  wire n784bar;
  wire n785bar;
  wire n786bar;
  wire n787bar;
  wire n788bar;
  wire n789bar;
  wire n790bar;
  wire n791bar;
  wire n792bar;
  wire n793bar;
  wire n794bar;
  wire n795bar;
  wire n796bar;
  wire n797bar;
  wire n798bar;
  wire n799bar;
  wire n800bar;
  wire n801bar;
  wire n802bar;
  wire n803bar;
  wire n804bar;
  wire n805bar;
  wire n806bar;
  wire n807bar;
  wire n808bar;
  wire n809bar;
  wire n810bar;
  wire n811bar;
  wire n812bar;
  wire n813bar;
  wire n814bar;
  wire n815bar;
  wire n816bar;
  wire n817bar;
  wire n818bar;
  wire n819bar;
  wire n820bar;
  wire n821bar;
  wire n822bar;
  wire n823bar;
  wire n824bar;
  wire n825bar;
  wire n826bar;
  wire n827bar;
  wire n828bar;
  wire n829bar;
  wire n830bar;
  wire n831bar;
  wire n832bar;
  wire n833bar;
  wire n834bar;
  wire n835bar;
  wire n836bar;
  wire n837bar;
  wire n838bar;
  wire n839bar;
  wire n840bar;
  wire n841bar;
  wire n842bar;
  wire n843bar;
  wire n844bar;
  wire n845bar;
  wire n846bar;
  wire n847bar;
  wire n848bar;
  wire n849bar;
  wire n850bar;
  wire n851bar;
  wire n852bar;
  wire n853bar;
  wire n854bar;
  wire n855bar;
  wire n856bar;
  wire n857bar;
  wire n858bar;
  wire n859bar;
  wire n860bar;
  wire n861bar;
  wire n862bar;
  wire n863bar;
  wire n864bar;
  wire n865bar;
  wire n866bar;
  wire n867bar;
  wire n868bar;
  wire n869bar;
  wire n870bar;
  wire n871bar;
  wire n872bar;
  wire n873bar;
  wire n874bar;
  wire n875bar;
  wire n876bar;
  wire n877bar;
  wire n878bar;
  wire n879bar;
  wire n880bar;
  wire n881bar;
  wire n882bar;
  wire n883bar;
  wire n884bar;
  wire n885bar;
  wire n886bar;
  wire n887bar;
  wire n888bar;
  wire n889bar;
  wire n890bar;
  wire n891bar;
  wire n892bar;
  wire n893bar;
  wire n894bar;
  wire n895bar;
  wire n896bar;
  wire n897bar;
  wire n898bar;
  wire n899bar;
  wire n900bar;
  wire n901bar;
  wire n902bar;
  wire n903bar;
  wire n904bar;
  wire n905bar;
  wire n906bar;
  wire n907bar;
  wire n908bar;
  wire n909bar;
  wire n910bar;
  wire n911bar;
  wire n912bar;
  wire n913bar;
  wire n914bar;
  wire n915bar;
  wire n916bar;
  wire n917bar;
  wire n918bar;
  wire n919bar;
  wire n920bar;
  wire n921bar;
  wire n922bar;
  wire n923bar;
  wire n924bar;
  wire n925bar;
  wire n926bar;
  wire n927bar;
  wire n928bar;
  wire n929bar;
  wire n930bar;
  wire n931bar;
  wire n932bar;
  wire n933bar;
  wire n934bar;
  wire n935bar;
  wire n936bar;
  wire n937bar;
  wire n938bar;
  wire n939bar;
  wire n940bar;
  wire n941bar;
  wire n942bar;
  wire n943bar;
  wire n944bar;
  wire n945bar;
  wire n946bar;
  wire n947bar;
  wire n948bar;
  wire n949bar;
  wire n950bar;
  wire n951bar;
  wire n952bar;
  wire n953bar;
  wire n954bar;
  wire n955bar;
  wire n956bar;
  wire n957bar;
  wire n958bar;
  wire n959bar;
  wire n960bar;
  wire n961bar;
  wire n962bar;
  wire n963bar;
  wire n964bar;
  wire n965bar;
  wire n966bar;
  wire n967bar;
  wire n968bar;
  wire n969bar;
  wire n970bar;
  wire n971bar;
  wire n972bar;
//wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];
  //OR U1
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1 (
    .O(out[7]),
    .I0(n972),
    .I1(n971)
  );
  //AND U1bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1bar (
    .O(outbar[7]),
    .I0(n972bar),
    .I1(n971bar)
  );
  //OR U2
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2 (
    .O(n971),
    .I0(n970),
    .I1(n969)
  );
  //AND U2bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2bar (
    .O(n971bar),
    .I0(n970bar),
    .I1(n969bar)
  );
  //OR U3
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3 (
    .O(n969),
    .I0(n968),
    .I1(n967)
  );
  //AND U3bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3bar (
    .O(n969bar),
    .I0(n968bar),
    .I1(n967bar)
  );
  //OR U4
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4 (
    .O(n967),
    .I0(n966),
    .I1(n965)
  );
  //AND U4bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4bar (
    .O(n967bar),
    .I0(n966bar),
    .I1(n965bar)
  );
  //OR U5
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5 (
    .O(n968),
    .I0(n964),
    .I1(n963)
  );
  //AND U5bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5bar (
    .O(n968bar),
    .I0(n964bar),
    .I1(n963bar)
  );
  //OR U6
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6 (
    .O(n963),
    .I0(in[116]),
    .I1(n962)
  );
  //AND U6bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6bar (
    .O(n963bar),
    .I0(inbar[116]),
    .I1(n962bar)
  );
  //OR U7
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7 (
    .O(n970),
    .I0(n961),
    .I1(n960)
  );
  //AND U7bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7bar (
    .O(n970bar),
    .I0(n961bar),
    .I1(n960bar)
  );
  //OR U8
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8 (
    .O(n960),
    .I0(in[150]),
    .I1(in[127])
  );
  //AND U8bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8bar (
    .O(n960bar),
    .I0(inbar[150]),
    .I1(inbar[127])
  );
  //OR U9
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9 (
    .O(n961),
    .I0(in[160]),
    .I1(n959)
  );
  //AND U9bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9bar (
    .O(n961bar),
    .I0(inbar[160]),
    .I1(n959bar)
  );
  //OR U10
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10 (
    .O(n959),
    .I0(in[252]),
    .I1(in[168])
  );
  //AND U10bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10bar (
    .O(n959bar),
    .I0(inbar[252]),
    .I1(inbar[168])
  );
  //OR U11
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11 (
    .O(n972),
    .I0(n958),
    .I1(n957)
  );
  //AND U11bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11bar (
    .O(n972bar),
    .I0(n958bar),
    .I1(n957bar)
  );
  //OR U12
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12 (
    .O(n957),
    .I0(n956),
    .I1(n955)
  );
  //AND U12bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12bar (
    .O(n957bar),
    .I0(n956bar),
    .I1(n955bar)
  );
  //OR U13
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13 (
    .O(n955),
    .I0(in_17),
    .I1(in[96])
  );
  //AND U13bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13bar (
    .O(n955bar),
    .I0(in_17bar),
    .I1(inbar[96])
  );
  //OR U14
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14 (
    .O(n956),
    .I0(in_23),
    .I1(n954)
  );
  //AND U14bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14bar (
    .O(n956bar),
    .I0(in_23bar),
    .I1(n954bar)
  );
  //OR U15
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15 (
    .O(n954),
    .I0(in_31),
    .I1(in_26)
  );
  //AND U15bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15bar (
    .O(n954bar),
    .I0(in_31bar),
    .I1(in_26bar)
  );
  //OR U16
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16 (
    .O(n958),
    .I0(n953),
    .I1(n952)
  );
  //AND U16bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16bar (
    .O(n958bar),
    .I0(n953bar),
    .I1(n952bar)
  );
  //OR U17
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U17 (
    .O(n952),
    .I0(in_58),
    .I1(in_4)
  );
  //AND U17bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U17bar (
    .O(n952bar),
    .I0(in_58bar),
    .I1(in_4bar)
  );
  //OR U18
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U18 (
    .O(n953),
    .I0(in_59),
    .I1(n951)
  );
  //AND U18bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U18bar (
    .O(n953bar),
    .I0(in_59bar),
    .I1(n951bar)
  );
  //OR U19
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U19 (
    .O(n951),
    .I0(in_71),
    .I1(in_62)
  );
  //AND U19bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U19bar (
    .O(n951bar),
    .I0(in_71bar),
    .I1(in_62bar)
  );
  //OR U20
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U20 (
    .O(out[6]),
    .I0(n950),
    .I1(n949)
  );
  //AND U20bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U20bar (
    .O(outbar[6]),
    .I0(n950bar),
    .I1(n949bar)
  );
  //OR U21
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U21 (
    .O(n949),
    .I0(n948),
    .I1(n947)
  );
  //AND U21bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U21bar (
    .O(n949bar),
    .I0(n948bar),
    .I1(n947bar)
  );
  //OR U22
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U22 (
    .O(n947),
    .I0(n946),
    .I1(n945)
  );
  //AND U22bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U22bar (
    .O(n947bar),
    .I0(n946bar),
    .I1(n945bar)
  );
  //OR U23
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U23 (
    .O(n945),
    .I0(n944),
    .I1(n943)
  );
  //AND U23bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U23bar (
    .O(n945bar),
    .I0(n944bar),
    .I1(n943bar)
  );
  //OR U24
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U24 (
    .O(n946),
    .I0(n942),
    .I1(n941)
  );
  //AND U24bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U24bar (
    .O(n946bar),
    .I0(n942bar),
    .I1(n941bar)
  );
  //OR U25
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U25 (
    .O(n941),
    .I0(in[101]),
    .I1(n940)
  );
  //AND U25bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U25bar (
    .O(n941bar),
    .I0(inbar[101]),
    .I1(n940bar)
  );
  //OR U26
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U26 (
    .O(n948),
    .I0(n939),
    .I1(n938)
  );
  //AND U26bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U26bar (
    .O(n948bar),
    .I0(n939bar),
    .I1(n938bar)
  );
  //OR U27
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U27 (
    .O(n938),
    .I0(in[114]),
    .I1(in[104])
  );
  //AND U27bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U27bar (
    .O(n938bar),
    .I0(inbar[114]),
    .I1(inbar[104])
  );
  //OR U28
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U28 (
    .O(n939),
    .I0(in[128]),
    .I1(n937)
  );
  //AND U28bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U28bar (
    .O(n939bar),
    .I0(inbar[128]),
    .I1(n937bar)
  );
  //OR U29
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U29 (
    .O(n937),
    .I0(in[136]),
    .I1(in[134])
  );
  //AND U29bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U29bar (
    .O(n937bar),
    .I0(inbar[136]),
    .I1(inbar[134])
  );
  //OR U30
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U30 (
    .O(n950),
    .I0(n936),
    .I1(n935)
  );
  //AND U30bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U30bar (
    .O(n950bar),
    .I0(n936bar),
    .I1(n935bar)
  );
  //OR U31
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U31 (
    .O(n935),
    .I0(n934),
    .I1(n933)
  );
  //AND U31bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U31bar (
    .O(n935bar),
    .I0(n934bar),
    .I1(n933bar)
  );
  //OR U32
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U32 (
    .O(n933),
    .I0(in[177]),
    .I1(in[164])
  );
  //AND U32bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U32bar (
    .O(n933bar),
    .I0(inbar[177]),
    .I1(inbar[164])
  );
  //OR U33
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U33 (
    .O(n934),
    .I0(in[212]),
    .I1(n932)
  );
  //AND U33bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U33bar (
    .O(n934bar),
    .I0(inbar[212]),
    .I1(n932bar)
  );
  //OR U34
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U34 (
    .O(n932),
    .I0(in[248]),
    .I1(in[221])
  );
  //AND U34bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U34bar (
    .O(n932bar),
    .I0(inbar[248]),
    .I1(inbar[221])
  );
  //OR U35
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U35 (
    .O(n936),
    .I0(n931),
    .I1(n930)
  );
  //AND U35bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U35bar (
    .O(n936bar),
    .I0(n931bar),
    .I1(n930bar)
  );
  //OR U36
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U36 (
    .O(n930),
    .I0(in_18),
    .I1(in[93])
  );
  //AND U36bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U36bar (
    .O(n930bar),
    .I0(in_18bar),
    .I1(inbar[93])
  );
  //OR U37
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U37 (
    .O(n931),
    .I0(in_31),
    .I1(n929)
  );
  //AND U37bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U37bar (
    .O(n931bar),
    .I0(in_31bar),
    .I1(n929bar)
  );
  //OR U38
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U38 (
    .O(n929),
    .I0(in_7),
    .I1(in_39)
  );
  //AND U38bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U38bar (
    .O(n929bar),
    .I0(in_7bar),
    .I1(in_39bar)
  );
  //OR U39
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U39 (
    .O(out[5]),
    .I0(n928),
    .I1(n927)
  );
  //AND U39bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U39bar (
    .O(outbar[5]),
    .I0(n928bar),
    .I1(n927bar)
  );
  //OR U40
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U40 (
    .O(n927),
    .I0(n926),
    .I1(n925)
  );
  //AND U40bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U40bar (
    .O(n927bar),
    .I0(n926bar),
    .I1(n925bar)
  );
  //OR U41
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U41 (
    .O(n925),
    .I0(n924),
    .I1(n923)
  );
  //AND U41bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U41bar (
    .O(n925bar),
    .I0(n924bar),
    .I1(n923bar)
  );
  //OR U42
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U42 (
    .O(n923),
    .I0(n922),
    .I1(n921)
  );
  //AND U42bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U42bar (
    .O(n923bar),
    .I0(n922bar),
    .I1(n921bar)
  );
  //OR U43
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U43 (
    .O(n924),
    .I0(n940),
    .I1(n920)
  );
  //AND U43bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U43bar (
    .O(n924bar),
    .I0(n940bar),
    .I1(n920bar)
  );
  //OR U44
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U44 (
    .O(n920),
    .I0(in[111]),
    .I1(n919)
  );
  //AND U44bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U44bar (
    .O(n920bar),
    .I0(inbar[111]),
    .I1(n919bar)
  );
  //OR U45
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U45 (
    .O(n940),
    .I0(n918),
    .I1(n917)
  );
  //AND U45bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U45bar (
    .O(n940bar),
    .I0(n918bar),
    .I1(n917bar)
  );
  //OR U46
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U46 (
    .O(n917),
    .I0(n916),
    .I1(n915)
  );
  //AND U46bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U46bar (
    .O(n917bar),
    .I0(n916bar),
    .I1(n915bar)
  );
  //OR U47
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U47 (
    .O(n915),
    .I0(n914),
    .I1(n913)
  );
  //AND U47bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U47bar (
    .O(n915bar),
    .I0(n914bar),
    .I1(n913bar)
  );
  //OR U48
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U48 (
    .O(n913),
    .I0(in[140]),
    .I1(in[131])
  );
  //AND U48bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U48bar (
    .O(n913bar),
    .I0(inbar[140]),
    .I1(inbar[131])
  );
  //OR U49
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U49 (
    .O(n914),
    .I0(in[160]),
    .I1(in[144])
  );
  //AND U49bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U49bar (
    .O(n914bar),
    .I0(inbar[160]),
    .I1(inbar[144])
  );
  //OR U50
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U50 (
    .O(n916),
    .I0(n912),
    .I1(n911)
  );
  //AND U50bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U50bar (
    .O(n916bar),
    .I0(n912bar),
    .I1(n911bar)
  );
  //OR U51
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U51 (
    .O(n911),
    .I0(in[179]),
    .I1(in[174])
  );
  //AND U51bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U51bar (
    .O(n911bar),
    .I0(inbar[179]),
    .I1(inbar[174])
  );
  //OR U52
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U52 (
    .O(n912),
    .I0(in[188]),
    .I1(in[184])
  );
  //AND U52bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U52bar (
    .O(n912bar),
    .I0(inbar[188]),
    .I1(inbar[184])
  );
  //OR U53
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U53 (
    .O(n918),
    .I0(n910),
    .I1(n909)
  );
  //AND U53bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U53bar (
    .O(n918bar),
    .I0(n910bar),
    .I1(n909bar)
  );
  //OR U54
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U54 (
    .O(n909),
    .I0(n908),
    .I1(n907)
  );
  //AND U54bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U54bar (
    .O(n909bar),
    .I0(n908bar),
    .I1(n907bar)
  );
  //OR U55
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U55 (
    .O(n907),
    .I0(in[216]),
    .I1(in[200])
  );
  //AND U55bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U55bar (
    .O(n907bar),
    .I0(inbar[216]),
    .I1(inbar[200])
  );
  //OR U56
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U56 (
    .O(n908),
    .I0(in[228]),
    .I1(in[224])
  );
  //AND U56bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U56bar (
    .O(n908bar),
    .I0(inbar[228]),
    .I1(inbar[224])
  );
  //OR U57
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U57 (
    .O(n910),
    .I0(n906),
    .I1(n905)
  );
  //AND U57bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U57bar (
    .O(n910bar),
    .I0(n906bar),
    .I1(n905bar)
  );
  //OR U58
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U58 (
    .O(n905),
    .I0(in[247]),
    .I1(in[235])
  );
  //AND U58bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U58bar (
    .O(n905bar),
    .I0(inbar[247]),
    .I1(inbar[235])
  );
  //OR U59
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U59 (
    .O(n906),
    .I0(in_42),
    .I1(in[83])
  );
  //AND U59bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U59bar (
    .O(n906bar),
    .I0(in_42bar),
    .I1(inbar[83])
  );
  //OR U60
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U60 (
    .O(n926),
    .I0(n904),
    .I1(n903)
  );
  //AND U60bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U60bar (
    .O(n926bar),
    .I0(n904bar),
    .I1(n903bar)
  );
  //OR U61
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U61 (
    .O(n903),
    .I0(in[166]),
    .I1(in[123])
  );
  //AND U61bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U61bar (
    .O(n903bar),
    .I0(inbar[166]),
    .I1(inbar[123])
  );
  //OR U62
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U62 (
    .O(n904),
    .I0(in[170]),
    .I1(n902)
  );
  //AND U62bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U62bar (
    .O(n904bar),
    .I0(inbar[170]),
    .I1(n902bar)
  );
  //OR U63
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U63 (
    .O(n902),
    .I0(in[194]),
    .I1(in[183])
  );
  //AND U63bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U63bar (
    .O(n902bar),
    .I0(inbar[194]),
    .I1(inbar[183])
  );
  //OR U64
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U64 (
    .O(n928),
    .I0(n901),
    .I1(n900)
  );
  //AND U64bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U64bar (
    .O(n928bar),
    .I0(n901bar),
    .I1(n900bar)
  );
  //OR U65
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U65 (
    .O(n900),
    .I0(n899),
    .I1(n898)
  );
  //AND U65bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U65bar (
    .O(n900bar),
    .I0(n899bar),
    .I1(n898bar)
  );
  //OR U66
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U66 (
    .O(n898),
    .I0(in[241]),
    .I1(in[238])
  );
  //AND U66bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U66bar (
    .O(n898bar),
    .I0(inbar[241]),
    .I1(inbar[238])
  );
  //OR U67
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U67 (
    .O(n899),
    .I0(in[250]),
    .I1(n897)
  );
  //AND U67bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U67bar (
    .O(n899bar),
    .I0(inbar[250]),
    .I1(n897bar)
  );
  //OR U68
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U68 (
    .O(n897),
    .I0(in_24),
    .I1(in[84])
  );
  //AND U68bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U68bar (
    .O(n897bar),
    .I0(in_24bar),
    .I1(inbar[84])
  );
  //OR U69
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U69 (
    .O(n901),
    .I0(n896),
    .I1(n895)
  );
  //AND U69bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U69bar (
    .O(n901bar),
    .I0(n896bar),
    .I1(n895bar)
  );
  //OR U70
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U70 (
    .O(n895),
    .I0(in_41),
    .I1(in_29)
  );
  //AND U70bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U70bar (
    .O(n895bar),
    .I0(in_41bar),
    .I1(in_29bar)
  );
  //OR U71
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U71 (
    .O(n896),
    .I0(in_66),
    .I1(n894)
  );
  //AND U71bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U71bar (
    .O(n896bar),
    .I0(in_66bar),
    .I1(n894bar)
  );
  //OR U72
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U72 (
    .O(n894),
    .I0(in_76),
    .I1(in_71)
  );
  //AND U72bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U72bar (
    .O(n894bar),
    .I0(in_76bar),
    .I1(in_71bar)
  );
  //OR U73
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U73 (
    .O(out[4]),
    .I0(n893),
    .I1(n892)
  );
  //AND U73bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U73bar (
    .O(outbar[4]),
    .I0(n893bar),
    .I1(n892bar)
  );
  //OR U74
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U74 (
    .O(n892),
    .I0(n891),
    .I1(n890)
  );
  //AND U74bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U74bar (
    .O(n892bar),
    .I0(n891bar),
    .I1(n890bar)
  );
  //OR U75
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U75 (
    .O(n890),
    .I0(n889),
    .I1(n888)
  );
  //AND U75bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U75bar (
    .O(n890bar),
    .I0(n889bar),
    .I1(n888bar)
  );
  //OR U76
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U76 (
    .O(n888),
    .I0(n922),
    .I1(n887)
  );
  //AND U76bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U76bar (
    .O(n888bar),
    .I0(n922bar),
    .I1(n887bar)
  );
  //OR U77
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U77 (
    .O(n922),
    .I0(n886),
    .I1(n885)
  );
  //AND U77bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U77bar (
    .O(n922bar),
    .I0(n886bar),
    .I1(n885bar)
  );
  //OR U78
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U78 (
    .O(n885),
    .I0(n884),
    .I1(n883)
  );
  //AND U78bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U78bar (
    .O(n885bar),
    .I0(n884bar),
    .I1(n883bar)
  );
  //OR U79
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U79 (
    .O(n883),
    .I0(n882),
    .I1(n881)
  );
  //AND U79bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U79bar (
    .O(n883bar),
    .I0(n882bar),
    .I1(n881bar)
  );
  //OR U80
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U80 (
    .O(n881),
    .I0(in[118]),
    .I1(in[109])
  );
  //AND U80bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U80bar (
    .O(n881bar),
    .I0(inbar[118]),
    .I1(inbar[109])
  );
  //OR U81
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U81 (
    .O(n882),
    .I0(in[139]),
    .I1(in[120])
  );
  //AND U81bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U81bar (
    .O(n882bar),
    .I0(inbar[139]),
    .I1(inbar[120])
  );
  //OR U82
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U82 (
    .O(n884),
    .I0(n880),
    .I1(n879)
  );
  //AND U82bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U82bar (
    .O(n884bar),
    .I0(n880bar),
    .I1(n879bar)
  );
  //OR U83
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U83 (
    .O(n879),
    .I0(in[198]),
    .I1(in[154])
  );
  //AND U83bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U83bar (
    .O(n879bar),
    .I0(inbar[198]),
    .I1(inbar[154])
  );
  //OR U84
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U84 (
    .O(n880),
    .I0(in[210]),
    .I1(in[205])
  );
  //AND U84bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U84bar (
    .O(n880bar),
    .I0(inbar[210]),
    .I1(inbar[205])
  );
  //OR U85
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U85 (
    .O(n886),
    .I0(n878),
    .I1(n877)
  );
  //AND U85bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U85bar (
    .O(n886bar),
    .I0(n878bar),
    .I1(n877bar)
  );
  //OR U86
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U86 (
    .O(n877),
    .I0(n876),
    .I1(n875)
  );
  //AND U86bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U86bar (
    .O(n877bar),
    .I0(n876bar),
    .I1(n875bar)
  );
  //OR U87
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U87 (
    .O(n875),
    .I0(in[219]),
    .I1(in[217])
  );
  //AND U87bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U87bar (
    .O(n875bar),
    .I0(inbar[219]),
    .I1(inbar[217])
  );
  //OR U88
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U88 (
    .O(n876),
    .I0(in[86]),
    .I1(in[252])
  );
  //AND U88bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U88bar (
    .O(n876bar),
    .I0(inbar[86]),
    .I1(inbar[252])
  );
  //OR U89
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U89 (
    .O(n878),
    .I0(n874),
    .I1(n873)
  );
  //AND U89bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U89bar (
    .O(n878bar),
    .I0(n874bar),
    .I1(n873bar)
  );
  //OR U90
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U90 (
    .O(n873),
    .I0(in_40),
    .I1(in[91])
  );
  //AND U90bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U90bar (
    .O(n873bar),
    .I0(in_40bar),
    .I1(inbar[91])
  );
  //OR U91
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U91 (
    .O(n874),
    .I0(in_8),
    .I1(in_46)
  );
  //AND U91bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U91bar (
    .O(n874bar),
    .I0(in_8bar),
    .I1(in_46bar)
  );
  //OR U92
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U92 (
    .O(n889),
    .I0(n872),
    .I1(n871)
  );
  //AND U92bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U92bar (
    .O(n889bar),
    .I0(n872bar),
    .I1(n871bar)
  );
  //OR U93
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U93 (
    .O(n871),
    .I0(in[117]),
    .I1(n943)
  );
  //AND U93bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U93bar (
    .O(n871bar),
    .I0(inbar[117]),
    .I1(n943bar)
  );
  //OR U94
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U94 (
    .O(n943),
    .I0(n870),
    .I1(n869)
  );
  //AND U94bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U94bar (
    .O(n943bar),
    .I0(n870bar),
    .I1(n869bar)
  );
  //OR U95
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U95 (
    .O(n869),
    .I0(n868),
    .I1(n867)
  );
  //AND U95bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U95bar (
    .O(n869bar),
    .I0(n868bar),
    .I1(n867bar)
  );
  //OR U96
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U96 (
    .O(n867),
    .I0(n866),
    .I1(n865)
  );
  //AND U96bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U96bar (
    .O(n867bar),
    .I0(n866bar),
    .I1(n865bar)
  );
  //OR U97
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U97 (
    .O(n865),
    .I0(n864),
    .I1(n863)
  );
  //AND U97bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U97bar (
    .O(n865bar),
    .I0(n864bar),
    .I1(n863bar)
  );
  //OR U98
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U98 (
    .O(n866),
    .I0(in[108]),
    .I1(n919)
  );
  //AND U98bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U98bar (
    .O(n866bar),
    .I0(inbar[108]),
    .I1(n919bar)
  );
  //OR U99
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U99 (
    .O(n919),
    .I0(n862),
    .I1(n861)
  );
  //AND U99bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U99bar (
    .O(n919bar),
    .I0(n862bar),
    .I1(n861bar)
  );
  //OR U100
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U100 (
    .O(n861),
    .I0(n860),
    .I1(n859)
  );
  //AND U100bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U100bar (
    .O(n861bar),
    .I0(n860bar),
    .I1(n859bar)
  );
  //OR U101
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U101 (
    .O(n859),
    .I0(n858),
    .I1(n857)
  );
  //AND U101bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U101bar (
    .O(n859bar),
    .I0(n858bar),
    .I1(n857bar)
  );
  //OR U102
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U102 (
    .O(n857),
    .I0(in[119]),
    .I1(in[105])
  );
  //AND U102bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U102bar (
    .O(n857bar),
    .I0(inbar[119]),
    .I1(inbar[105])
  );
  //OR U103
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U103 (
    .O(n858),
    .I0(in[186]),
    .I1(in[175])
  );
  //AND U103bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U103bar (
    .O(n858bar),
    .I0(inbar[186]),
    .I1(inbar[175])
  );
  //OR U104
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U104 (
    .O(n860),
    .I0(n856),
    .I1(n855)
  );
  //AND U104bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U104bar (
    .O(n860bar),
    .I0(n856bar),
    .I1(n855bar)
  );
  //OR U105
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U105 (
    .O(n855),
    .I0(in[202]),
    .I1(in[193])
  );
  //AND U105bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U105bar (
    .O(n855bar),
    .I0(inbar[202]),
    .I1(inbar[193])
  );
  //OR U106
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U106 (
    .O(n856),
    .I0(in[225]),
    .I1(in[208])
  );
  //AND U106bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U106bar (
    .O(n856bar),
    .I0(inbar[225]),
    .I1(inbar[208])
  );
  //OR U107
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U107 (
    .O(n862),
    .I0(n854),
    .I1(n853)
  );
  //AND U107bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U107bar (
    .O(n862bar),
    .I0(n854bar),
    .I1(n853bar)
  );
  //OR U108
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U108 (
    .O(n853),
    .I0(n852),
    .I1(n851)
  );
  //AND U108bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U108bar (
    .O(n853bar),
    .I0(n852bar),
    .I1(n851bar)
  );
  //OR U109
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U109 (
    .O(n851),
    .I0(in_1),
    .I1(in[85])
  );
  //AND U109bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U109bar (
    .O(n851bar),
    .I0(in_1bar),
    .I1(inbar[85])
  );
  //OR U110
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U110 (
    .O(n852),
    .I0(in_23),
    .I1(in_19)
  );
  //AND U110bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U110bar (
    .O(n852bar),
    .I0(in_23bar),
    .I1(in_19bar)
  );
  //OR U111
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U111 (
    .O(n854),
    .I0(n850),
    .I1(n849)
  );
  //AND U111bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U111bar (
    .O(n854bar),
    .I0(n850bar),
    .I1(n849bar)
  );
  //OR U112
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U112 (
    .O(n849),
    .I0(in_43),
    .I1(in_33)
  );
  //AND U112bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U112bar (
    .O(n849bar),
    .I0(in_43bar),
    .I1(in_33bar)
  );
  //OR U113
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U113 (
    .O(n850),
    .I0(in_63),
    .I1(in_44)
  );
  //AND U113bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U113bar (
    .O(n850bar),
    .I0(in_63bar),
    .I1(in_44bar)
  );
  //OR U114
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U114 (
    .O(n868),
    .I0(n848),
    .I1(n847)
  );
  //AND U114bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U114bar (
    .O(n868bar),
    .I0(n848bar),
    .I1(n847bar)
  );
  //OR U115
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U115 (
    .O(n847),
    .I0(in[141]),
    .I1(in[112])
  );
  //AND U115bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U115bar (
    .O(n847bar),
    .I0(inbar[141]),
    .I1(inbar[112])
  );
  //OR U116
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U116 (
    .O(n848),
    .I0(in[147]),
    .I1(n846)
  );
  //AND U116bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U116bar (
    .O(n848bar),
    .I0(inbar[147]),
    .I1(n846bar)
  );
  //OR U117
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U117 (
    .O(n846),
    .I0(in[181]),
    .I1(in[167])
  );
  //AND U117bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U117bar (
    .O(n846bar),
    .I0(inbar[181]),
    .I1(inbar[167])
  );
  //OR U118
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U118 (
    .O(n870),
    .I0(n845),
    .I1(n844)
  );
  //AND U118bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U118bar (
    .O(n870bar),
    .I0(n845bar),
    .I1(n844bar)
  );
  //OR U119
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U119 (
    .O(n844),
    .I0(n843),
    .I1(n842)
  );
  //AND U119bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U119bar (
    .O(n844bar),
    .I0(n843bar),
    .I1(n842bar)
  );
  //OR U120
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U120 (
    .O(n842),
    .I0(in[229]),
    .I1(in[201])
  );
  //AND U120bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U120bar (
    .O(n842bar),
    .I0(inbar[229]),
    .I1(inbar[201])
  );
  //OR U121
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U121 (
    .O(n843),
    .I0(in[237]),
    .I1(n841)
  );
  //AND U121bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U121bar (
    .O(n843bar),
    .I0(inbar[237]),
    .I1(n841bar)
  );
  //OR U122
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U122 (
    .O(n841),
    .I0(in[94]),
    .I1(in[253])
  );
  //AND U122bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U122bar (
    .O(n841bar),
    .I0(inbar[94]),
    .I1(inbar[253])
  );
  //OR U123
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U123 (
    .O(n845),
    .I0(n840),
    .I1(n839)
  );
  //AND U123bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U123bar (
    .O(n845bar),
    .I0(n840bar),
    .I1(n839bar)
  );
  //OR U124
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U124 (
    .O(n839),
    .I0(in_21),
    .I1(in[96])
  );
  //AND U124bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U124bar (
    .O(n839bar),
    .I0(in_21bar),
    .I1(inbar[96])
  );
  //OR U125
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U125 (
    .O(n840),
    .I0(in_25),
    .I1(n838)
  );
  //AND U125bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U125bar (
    .O(n840bar),
    .I0(in_25bar),
    .I1(n838bar)
  );
  //OR U126
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U126 (
    .O(n838),
    .I0(in_81),
    .I1(in_45)
  );
  //AND U126bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U126bar (
    .O(n838bar),
    .I0(in_81bar),
    .I1(in_45bar)
  );
  //OR U127
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U127 (
    .O(n891),
    .I0(n837),
    .I1(n836)
  );
  //AND U127bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U127bar (
    .O(n891bar),
    .I0(n837bar),
    .I1(n836bar)
  );
  //OR U128
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U128 (
    .O(n836),
    .I0(in[142]),
    .I1(in[124])
  );
  //AND U128bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U128bar (
    .O(n836bar),
    .I0(inbar[142]),
    .I1(inbar[124])
  );
  //OR U129
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U129 (
    .O(n837),
    .I0(in[150]),
    .I1(n835)
  );
  //AND U129bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U129bar (
    .O(n837bar),
    .I0(inbar[150]),
    .I1(n835bar)
  );
  //OR U130
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U130 (
    .O(n835),
    .I0(in[172]),
    .I1(in[155])
  );
  //AND U130bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U130bar (
    .O(n835bar),
    .I0(inbar[172]),
    .I1(inbar[155])
  );
  //OR U131
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U131 (
    .O(n893),
    .I0(n834),
    .I1(n833)
  );
  //AND U131bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U131bar (
    .O(n893bar),
    .I0(n834bar),
    .I1(n833bar)
  );
  //OR U132
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U132 (
    .O(n833),
    .I0(n832),
    .I1(n831)
  );
  //AND U132bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U132bar (
    .O(n833bar),
    .I0(n832bar),
    .I1(n831bar)
  );
  //OR U133
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U133 (
    .O(n831),
    .I0(in[196]),
    .I1(in[173])
  );
  //AND U133bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U133bar (
    .O(n831bar),
    .I0(inbar[196]),
    .I1(inbar[173])
  );
  //OR U134
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U134 (
    .O(n832),
    .I0(in[222]),
    .I1(n830)
  );
  //AND U134bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U134bar (
    .O(n832bar),
    .I0(inbar[222]),
    .I1(n830bar)
  );
  //OR U135
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U135 (
    .O(n830),
    .I0(in[227]),
    .I1(in[226])
  );
  //AND U135bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U135bar (
    .O(n830bar),
    .I0(inbar[227]),
    .I1(inbar[226])
  );
  //OR U136
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U136 (
    .O(n834),
    .I0(n829),
    .I1(n828)
  );
  //AND U136bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U136bar (
    .O(n834bar),
    .I0(n829bar),
    .I1(n828bar)
  );
  //OR U137
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U137 (
    .O(n828),
    .I0(in[249]),
    .I1(in[231])
  );
  //AND U137bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U137bar (
    .O(n828bar),
    .I0(inbar[249]),
    .I1(inbar[231])
  );
  //OR U138
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U138 (
    .O(n829),
    .I0(in_28),
    .I1(n827)
  );
  //AND U138bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U138bar (
    .O(n829bar),
    .I0(in_28bar),
    .I1(n827bar)
  );
  //OR U139
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U139 (
    .O(n827),
    .I0(in_52),
    .I1(in_47)
  );
  //AND U139bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U139bar (
    .O(n827bar),
    .I0(in_52bar),
    .I1(in_47bar)
  );
  //OR U140
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U140 (
    .O(out[3]),
    .I0(n826),
    .I1(n825)
  );
  //AND U140bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U140bar (
    .O(outbar[3]),
    .I0(n826bar),
    .I1(n825bar)
  );
  //OR U141
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U141 (
    .O(n825),
    .I0(n824),
    .I1(n823)
  );
  //AND U141bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U141bar (
    .O(n825bar),
    .I0(n824bar),
    .I1(n823bar)
  );
  //OR U142
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U142 (
    .O(n823),
    .I0(n822),
    .I1(n821)
  );
  //AND U142bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U142bar (
    .O(n823bar),
    .I0(n822bar),
    .I1(n821bar)
  );
  //OR U143
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U143 (
    .O(n821),
    .I0(n820),
    .I1(n819)
  );
  //AND U143bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U143bar (
    .O(n821bar),
    .I0(n820bar),
    .I1(n819bar)
  );
  //OR U144
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U144 (
    .O(n822),
    .I0(n964),
    .I1(n818)
  );
  //AND U144bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U144bar (
    .O(n822bar),
    .I0(n964bar),
    .I1(n818bar)
  );
  //OR U145
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U145 (
    .O(n818),
    .I0(in[118]),
    .I1(n817)
  );
  //AND U145bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U145bar (
    .O(n818bar),
    .I0(inbar[118]),
    .I1(n817bar)
  );
  //OR U146
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U146 (
    .O(n964),
    .I0(n816),
    .I1(n815)
  );
  //AND U146bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U146bar (
    .O(n964bar),
    .I0(n816bar),
    .I1(n815bar)
  );
  //OR U147
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U147 (
    .O(n815),
    .I0(n814),
    .I1(n813)
  );
  //AND U147bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U147bar (
    .O(n815bar),
    .I0(n814bar),
    .I1(n813bar)
  );
  //OR U148
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U148 (
    .O(n813),
    .I0(n812),
    .I1(n811)
  );
  //AND U148bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U148bar (
    .O(n813bar),
    .I0(n812bar),
    .I1(n811bar)
  );
  //OR U149
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U149 (
    .O(n811),
    .I0(in[122]),
    .I1(in[111])
  );
  //AND U149bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U149bar (
    .O(n811bar),
    .I0(inbar[122]),
    .I1(inbar[111])
  );
  //OR U150
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U150 (
    .O(n812),
    .I0(in[154]),
    .I1(in[151])
  );
  //AND U150bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U150bar (
    .O(n812bar),
    .I0(inbar[154]),
    .I1(inbar[151])
  );
  //OR U151
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U151 (
    .O(n814),
    .I0(n810),
    .I1(n809)
  );
  //AND U151bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U151bar (
    .O(n814bar),
    .I0(n810bar),
    .I1(n809bar)
  );
  //OR U152
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U152 (
    .O(n809),
    .I0(in[187]),
    .I1(in[177])
  );
  //AND U152bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U152bar (
    .O(n809bar),
    .I0(inbar[187]),
    .I1(inbar[177])
  );
  //OR U153
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U153 (
    .O(n810),
    .I0(in[200]),
    .I1(in[192])
  );
  //AND U153bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U153bar (
    .O(n810bar),
    .I0(inbar[200]),
    .I1(inbar[192])
  );
  //OR U154
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U154 (
    .O(n816),
    .I0(n808),
    .I1(n807)
  );
  //AND U154bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U154bar (
    .O(n816bar),
    .I0(n808bar),
    .I1(n807bar)
  );
  //OR U155
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U155 (
    .O(n807),
    .I0(n806),
    .I1(n805)
  );
  //AND U155bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U155bar (
    .O(n807bar),
    .I0(n806bar),
    .I1(n805bar)
  );
  //OR U156
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U156 (
    .O(n805),
    .I0(in[225]),
    .I1(in[207])
  );
  //AND U156bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U156bar (
    .O(n805bar),
    .I0(inbar[225]),
    .I1(inbar[207])
  );
  //OR U157
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U157 (
    .O(n806),
    .I0(in[98]),
    .I1(in[226])
  );
  //AND U157bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U157bar (
    .O(n806bar),
    .I0(inbar[98]),
    .I1(inbar[226])
  );
  //OR U158
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U158 (
    .O(n808),
    .I0(n804),
    .I1(n803)
  );
  //AND U158bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U158bar (
    .O(n808bar),
    .I0(n804bar),
    .I1(n803bar)
  );
  //OR U159
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U159 (
    .O(n803),
    .I0(in_20),
    .I1(in_16)
  );
  //AND U159bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U159bar (
    .O(n803bar),
    .I0(in_20bar),
    .I1(in_16bar)
  );
  //OR U160
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U160 (
    .O(n804),
    .I0(in_55),
    .I1(in_45)
  );
  //AND U160bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U160bar (
    .O(n804bar),
    .I0(in_55bar),
    .I1(in_45bar)
  );
  //OR U161
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U161 (
    .O(n824),
    .I0(n802),
    .I1(n801)
  );
  //AND U161bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U161bar (
    .O(n824bar),
    .I0(n802bar),
    .I1(n801bar)
  );
  //OR U162
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U162 (
    .O(n801),
    .I0(in[162]),
    .I1(in[149])
  );
  //AND U162bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U162bar (
    .O(n801bar),
    .I0(inbar[162]),
    .I1(inbar[149])
  );
  //OR U163
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U163 (
    .O(n802),
    .I0(in[163]),
    .I1(n800)
  );
  //AND U163bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U163bar (
    .O(n802bar),
    .I0(inbar[163]),
    .I1(n800bar)
  );
  //OR U164
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U164 (
    .O(n800),
    .I0(in[191]),
    .I1(in[189])
  );
  //AND U164bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U164bar (
    .O(n800bar),
    .I0(inbar[191]),
    .I1(inbar[189])
  );
  //OR U165
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U165 (
    .O(n826),
    .I0(n799),
    .I1(n798)
  );
  //AND U165bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U165bar (
    .O(n826bar),
    .I0(n799bar),
    .I1(n798bar)
  );
  //OR U166
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U166 (
    .O(n798),
    .I0(n797),
    .I1(n796)
  );
  //AND U166bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U166bar (
    .O(n798bar),
    .I0(n797bar),
    .I1(n796bar)
  );
  //OR U167
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U167 (
    .O(n796),
    .I0(in[212]),
    .I1(in[193])
  );
  //AND U167bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U167bar (
    .O(n796bar),
    .I0(inbar[212]),
    .I1(inbar[193])
  );
  //OR U168
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U168 (
    .O(n797),
    .I0(in[238]),
    .I1(n795)
  );
  //AND U168bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U168bar (
    .O(n797bar),
    .I0(inbar[238]),
    .I1(n795bar)
  );
  //OR U169
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U169 (
    .O(n795),
    .I0(in[88]),
    .I1(in[247])
  );
  //AND U169bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U169bar (
    .O(n795bar),
    .I0(inbar[88]),
    .I1(inbar[247])
  );
  //OR U170
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U170 (
    .O(n799),
    .I0(n794),
    .I1(n793)
  );
  //AND U170bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U170bar (
    .O(n799bar),
    .I0(n794bar),
    .I1(n793bar)
  );
  //OR U171
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U171 (
    .O(n793),
    .I0(in[94]),
    .I1(in[92])
  );
  //AND U171bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U171bar (
    .O(n793bar),
    .I0(inbar[94]),
    .I1(inbar[92])
  );
  //OR U172
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U172 (
    .O(n794),
    .I0(in_52),
    .I1(n792)
  );
  //AND U172bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U172bar (
    .O(n794bar),
    .I0(in_52bar),
    .I1(n792bar)
  );
  //OR U173
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U173 (
    .O(n792),
    .I0(in_70),
    .I1(in_67)
  );
  //AND U173bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U173bar (
    .O(n792bar),
    .I0(in_70bar),
    .I1(in_67bar)
  );
  //OR U174
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U174 (
    .O(out[2]),
    .I0(n791),
    .I1(n790)
  );
  //AND U174bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U174bar (
    .O(outbar[2]),
    .I0(n791bar),
    .I1(n790bar)
  );
  //OR U175
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U175 (
    .O(n790),
    .I0(n789),
    .I1(n788)
  );
  //AND U175bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U175bar (
    .O(n790bar),
    .I0(n789bar),
    .I1(n788bar)
  );
  //OR U176
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U176 (
    .O(n788),
    .I0(n787),
    .I1(n786)
  );
  //AND U176bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U176bar (
    .O(n788bar),
    .I0(n787bar),
    .I1(n786bar)
  );
  //OR U177
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U177 (
    .O(n786),
    .I0(n819),
    .I1(n785)
  );
  //AND U177bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U177bar (
    .O(n786bar),
    .I0(n819bar),
    .I1(n785bar)
  );
  //OR U178
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U178 (
    .O(n819),
    .I0(n784),
    .I1(n783)
  );
  //AND U178bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U178bar (
    .O(n819bar),
    .I0(n784bar),
    .I1(n783bar)
  );
  //OR U179
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U179 (
    .O(n783),
    .I0(n782),
    .I1(n781)
  );
  //AND U179bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U179bar (
    .O(n783bar),
    .I0(n782bar),
    .I1(n781bar)
  );
  //OR U180
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U180 (
    .O(n781),
    .I0(n780),
    .I1(n779)
  );
  //AND U180bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U180bar (
    .O(n781bar),
    .I0(n780bar),
    .I1(n779bar)
  );
  //OR U181
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U181 (
    .O(n779),
    .I0(n962),
    .I1(n778)
  );
  //AND U181bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U181bar (
    .O(n779bar),
    .I0(n962bar),
    .I1(n778bar)
  );
  //OR U182
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U182 (
    .O(n962),
    .I0(n777),
    .I1(n776)
  );
  //AND U182bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U182bar (
    .O(n962bar),
    .I0(n777bar),
    .I1(n776bar)
  );
  //OR U183
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U183 (
    .O(n776),
    .I0(n775),
    .I1(n774)
  );
  //AND U183bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U183bar (
    .O(n776bar),
    .I0(n775bar),
    .I1(n774bar)
  );
  //OR U184
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U184 (
    .O(n774),
    .I0(n773),
    .I1(n772)
  );
  //AND U184bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U184bar (
    .O(n774bar),
    .I0(n773bar),
    .I1(n772bar)
  );
  //OR U185
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U185 (
    .O(n772),
    .I0(in[131]),
    .I1(in[120])
  );
  //AND U185bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U185bar (
    .O(n772bar),
    .I0(inbar[131]),
    .I1(inbar[120])
  );
  //OR U186
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U186 (
    .O(n773),
    .I0(in[153]),
    .I1(in[147])
  );
  //AND U186bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U186bar (
    .O(n773bar),
    .I0(inbar[153]),
    .I1(inbar[147])
  );
  //OR U187
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U187 (
    .O(n775),
    .I0(n771),
    .I1(n770)
  );
  //AND U187bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U187bar (
    .O(n775bar),
    .I0(n771bar),
    .I1(n770bar)
  );
  //OR U188
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U188 (
    .O(n770),
    .I0(in[170]),
    .I1(in[156])
  );
  //AND U188bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U188bar (
    .O(n770bar),
    .I0(inbar[170]),
    .I1(inbar[156])
  );
  //OR U189
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U189 (
    .O(n771),
    .I0(in[223]),
    .I1(in[190])
  );
  //AND U189bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U189bar (
    .O(n771bar),
    .I0(inbar[223]),
    .I1(inbar[190])
  );
  //OR U190
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U190 (
    .O(n777),
    .I0(n769),
    .I1(n768)
  );
  //AND U190bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U190bar (
    .O(n777bar),
    .I0(n769bar),
    .I1(n768bar)
  );
  //OR U191
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U191 (
    .O(n768),
    .I0(n767),
    .I1(n766)
  );
  //AND U191bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U191bar (
    .O(n768bar),
    .I0(n767bar),
    .I1(n766bar)
  );
  //OR U192
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U192 (
    .O(n766),
    .I0(in[236]),
    .I1(in[230])
  );
  //AND U192bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U192bar (
    .O(n766bar),
    .I0(inbar[236]),
    .I1(inbar[230])
  );
  //OR U193
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U193 (
    .O(n767),
    .I0(in[85]),
    .I1(in[240])
  );
  //AND U193bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U193bar (
    .O(n767bar),
    .I0(inbar[85]),
    .I1(inbar[240])
  );
  //OR U194
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U194 (
    .O(n769),
    .I0(n765),
    .I1(n764)
  );
  //AND U194bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U194bar (
    .O(n769bar),
    .I0(n765bar),
    .I1(n764bar)
  );
  //OR U195
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U195 (
    .O(n764),
    .I0(in_12),
    .I1(in[90])
  );
  //AND U195bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U195bar (
    .O(n764bar),
    .I0(in_12bar),
    .I1(inbar[90])
  );
  //OR U196
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U196 (
    .O(n765),
    .I0(in_39),
    .I1(in_28)
  );
  //AND U196bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U196bar (
    .O(n765bar),
    .I0(in_39bar),
    .I1(in_28bar)
  );
  //OR U197
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U197 (
    .O(n780),
    .I0(in[109]),
    .I1(n763)
  );
  //AND U197bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U197bar (
    .O(n780bar),
    .I0(inbar[109]),
    .I1(n763bar)
  );
  //OR U198
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U198 (
    .O(n782),
    .I0(n762),
    .I1(n761)
  );
  //AND U198bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U198bar (
    .O(n782bar),
    .I0(n762bar),
    .I1(n761bar)
  );
  //OR U199
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U199 (
    .O(n761),
    .I0(in[138]),
    .I1(in[129])
  );
  //AND U199bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U199bar (
    .O(n761bar),
    .I0(inbar[138]),
    .I1(inbar[129])
  );
  //OR U200
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U200 (
    .O(n762),
    .I0(in[157]),
    .I1(n760)
  );
  //AND U200bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U200bar (
    .O(n762bar),
    .I0(inbar[157]),
    .I1(n760bar)
  );
  //OR U201
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U201 (
    .O(n760),
    .I0(in[182]),
    .I1(in[167])
  );
  //AND U201bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U201bar (
    .O(n760bar),
    .I0(inbar[182]),
    .I1(inbar[167])
  );
  //OR U202
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U202 (
    .O(n784),
    .I0(n759),
    .I1(n758)
  );
  //AND U202bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U202bar (
    .O(n784bar),
    .I0(n759bar),
    .I1(n758bar)
  );
  //OR U203
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U203 (
    .O(n758),
    .I0(n757),
    .I1(n756)
  );
  //AND U203bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U203bar (
    .O(n758bar),
    .I0(n757bar),
    .I1(n756bar)
  );
  //OR U204
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U204 (
    .O(n756),
    .I0(in[195]),
    .I1(in[184])
  );
  //AND U204bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U204bar (
    .O(n756bar),
    .I0(inbar[195]),
    .I1(inbar[184])
  );
  //OR U205
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U205 (
    .O(n757),
    .I0(in[196]),
    .I1(n755)
  );
  //AND U205bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U205bar (
    .O(n757bar),
    .I0(inbar[196]),
    .I1(n755bar)
  );
  //OR U206
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U206 (
    .O(n755),
    .I0(in[215]),
    .I1(in[209])
  );
  //AND U206bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U206bar (
    .O(n755bar),
    .I0(inbar[215]),
    .I1(inbar[209])
  );
  //OR U207
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U207 (
    .O(n759),
    .I0(n754),
    .I1(n753)
  );
  //AND U207bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U207bar (
    .O(n759bar),
    .I0(n754bar),
    .I1(n753bar)
  );
  //OR U208
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U208 (
    .O(n753),
    .I0(in[93]),
    .I1(in[233])
  );
  //AND U208bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U208bar (
    .O(n753bar),
    .I0(inbar[93]),
    .I1(inbar[233])
  );
  //OR U209
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U209 (
    .O(n754),
    .I0(in_1),
    .I1(n752)
  );
  //AND U209bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U209bar (
    .O(n754bar),
    .I0(in_1bar),
    .I1(n752bar)
  );
  //OR U210
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U210 (
    .O(n752),
    .I0(in_69),
    .I1(in_66)
  );
  //AND U210bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U210bar (
    .O(n752bar),
    .I0(in_69bar),
    .I1(in_66bar)
  );
  //OR U211
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U211 (
    .O(n787),
    .I0(n966),
    .I1(n751)
  );
  //AND U211bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U211bar (
    .O(n787bar),
    .I0(n966bar),
    .I1(n751bar)
  );
  //OR U212
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U212 (
    .O(n751),
    .I0(in[134]),
    .I1(n750)
  );
  //AND U212bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U212bar (
    .O(n751bar),
    .I0(inbar[134]),
    .I1(n750bar)
  );
  //OR U213
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U213 (
    .O(n966),
    .I0(n749),
    .I1(n748)
  );
  //AND U213bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U213bar (
    .O(n966bar),
    .I0(n749bar),
    .I1(n748bar)
  );
  //OR U214
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U214 (
    .O(n748),
    .I0(n747),
    .I1(n746)
  );
  //AND U214bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U214bar (
    .O(n748bar),
    .I0(n747bar),
    .I1(n746bar)
  );
  //OR U215
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U215 (
    .O(n746),
    .I0(n745),
    .I1(n744)
  );
  //AND U215bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U215bar (
    .O(n746bar),
    .I0(n745bar),
    .I1(n744bar)
  );
  //OR U216
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U216 (
    .O(n744),
    .I0(in[136]),
    .I1(in[121])
  );
  //AND U216bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U216bar (
    .O(n744bar),
    .I0(inbar[136]),
    .I1(inbar[121])
  );
  //OR U217
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U217 (
    .O(n745),
    .I0(in[186]),
    .I1(in[174])
  );
  //AND U217bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U217bar (
    .O(n745bar),
    .I0(inbar[186]),
    .I1(inbar[174])
  );
  //OR U218
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U218 (
    .O(n747),
    .I0(n743),
    .I1(n742)
  );
  //AND U218bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U218bar (
    .O(n747bar),
    .I0(n743bar),
    .I1(n742bar)
  );
  //OR U219
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U219 (
    .O(n742),
    .I0(in[198]),
    .I1(in[197])
  );
  //AND U219bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U219bar (
    .O(n742bar),
    .I0(inbar[198]),
    .I1(inbar[197])
  );
  //OR U220
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U220 (
    .O(n743),
    .I0(in[214]),
    .I1(in[199])
  );
  //AND U220bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U220bar (
    .O(n743bar),
    .I0(inbar[214]),
    .I1(inbar[199])
  );
  //OR U221
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U221 (
    .O(n749),
    .I0(n741),
    .I1(n740)
  );
  //AND U221bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U221bar (
    .O(n749bar),
    .I0(n741bar),
    .I1(n740bar)
  );
  //OR U222
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U222 (
    .O(n740),
    .I0(n739),
    .I1(n738)
  );
  //AND U222bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U222bar (
    .O(n740bar),
    .I0(n739bar),
    .I1(n738bar)
  );
  //OR U223
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U223 (
    .O(n738),
    .I0(in[231]),
    .I1(in[220])
  );
  //AND U223bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U223bar (
    .O(n738bar),
    .I0(inbar[231]),
    .I1(inbar[220])
  );
  //OR U224
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U224 (
    .O(n739),
    .I0(in_25),
    .I1(in[245])
  );
  //AND U224bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U224bar (
    .O(n739bar),
    .I0(in_25bar),
    .I1(inbar[245])
  );
  //OR U225
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U225 (
    .O(n741),
    .I0(n737),
    .I1(n736)
  );
  //AND U225bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U225bar (
    .O(n741bar),
    .I0(n737bar),
    .I1(n736bar)
  );
  //OR U226
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U226 (
    .O(n736),
    .I0(in_53),
    .I1(in_29)
  );
  //AND U226bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U226bar (
    .O(n736bar),
    .I0(in_53bar),
    .I1(in_29bar)
  );
  //OR U227
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U227 (
    .O(n737),
    .I0(in_79),
    .I1(in_74)
  );
  //AND U227bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U227bar (
    .O(n737bar),
    .I0(in_79bar),
    .I1(in_74bar)
  );
  //OR U228
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U228 (
    .O(n789),
    .I0(n735),
    .I1(n734)
  );
  //AND U228bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U228bar (
    .O(n789bar),
    .I0(n735bar),
    .I1(n734bar)
  );
  //OR U229
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U229 (
    .O(n734),
    .I0(in[152]),
    .I1(in[140])
  );
  //AND U229bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U229bar (
    .O(n734bar),
    .I0(inbar[152]),
    .I1(inbar[140])
  );
  //OR U230
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U230 (
    .O(n735),
    .I0(in[155]),
    .I1(n733)
  );
  //AND U230bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U230bar (
    .O(n735bar),
    .I0(inbar[155]),
    .I1(n733bar)
  );
  //OR U231
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U231 (
    .O(n733),
    .I0(in[166]),
    .I1(in[165])
  );
  //AND U231bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U231bar (
    .O(n733bar),
    .I0(inbar[166]),
    .I1(inbar[165])
  );
  //OR U232
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U232 (
    .O(n791),
    .I0(n732),
    .I1(n731)
  );
  //AND U232bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U232bar (
    .O(n791bar),
    .I0(n732bar),
    .I1(n731bar)
  );
  //OR U233
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U233 (
    .O(n731),
    .I0(n730),
    .I1(n729)
  );
  //AND U233bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U233bar (
    .O(n731bar),
    .I0(n730bar),
    .I1(n729bar)
  );
  //OR U234
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U234 (
    .O(n729),
    .I0(in[202]),
    .I1(in[185])
  );
  //AND U234bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U234bar (
    .O(n729bar),
    .I0(inbar[202]),
    .I1(inbar[185])
  );
  //OR U235
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U235 (
    .O(n730),
    .I0(in[211]),
    .I1(n728)
  );
  //AND U235bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U235bar (
    .O(n730bar),
    .I0(inbar[211]),
    .I1(n728bar)
  );
  //OR U236
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U236 (
    .O(n728),
    .I0(in[255]),
    .I1(in[253])
  );
  //AND U236bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U236bar (
    .O(n728bar),
    .I0(inbar[255]),
    .I1(inbar[253])
  );
  //OR U237
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U237 (
    .O(n732),
    .I0(n727),
    .I1(n726)
  );
  //AND U237bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U237bar (
    .O(n732bar),
    .I0(n727bar),
    .I1(n726bar)
  );
  //OR U238
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U238 (
    .O(n726),
    .I0(in_35),
    .I1(in_15)
  );
  //AND U238bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U238bar (
    .O(n726bar),
    .I0(in_35bar),
    .I1(in_15bar)
  );
  //OR U239
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U239 (
    .O(n727),
    .I0(in_36),
    .I1(n725)
  );
  //AND U239bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U239bar (
    .O(n727bar),
    .I0(in_36bar),
    .I1(n725bar)
  );
  //OR U240
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U240 (
    .O(n725),
    .I0(in_48),
    .I1(in_40)
  );
  //AND U240bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U240bar (
    .O(n725bar),
    .I0(in_48bar),
    .I1(in_40bar)
  );
  //OR U241
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U241 (
    .O(out[1]),
    .I0(n724),
    .I1(n723)
  );
  //AND U241bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U241bar (
    .O(outbar[1]),
    .I0(n724bar),
    .I1(n723bar)
  );
  //OR U242
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U242 (
    .O(n723),
    .I0(n722),
    .I1(n721)
  );
  //AND U242bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U242bar (
    .O(n723bar),
    .I0(n722bar),
    .I1(n721bar)
  );
  //OR U243
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U243 (
    .O(n721),
    .I0(n720),
    .I1(n719)
  );
  //AND U243bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U243bar (
    .O(n721bar),
    .I0(n720bar),
    .I1(n719bar)
  );
  //OR U244
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U244 (
    .O(n719),
    .I0(n921),
    .I1(n887)
  );
  //AND U244bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U244bar (
    .O(n719bar),
    .I0(n921bar),
    .I1(n887bar)
  );
  //OR U245
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U245 (
    .O(n887),
    .I0(n718),
    .I1(n717)
  );
  //AND U245bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U245bar (
    .O(n887bar),
    .I0(n718bar),
    .I1(n717bar)
  );
  //OR U246
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U246 (
    .O(n717),
    .I0(n716),
    .I1(n715)
  );
  //AND U246bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U246bar (
    .O(n717bar),
    .I0(n716bar),
    .I1(n715bar)
  );
  //OR U247
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U247 (
    .O(n715),
    .I0(n714),
    .I1(n713)
  );
  //AND U247bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U247bar (
    .O(n715bar),
    .I0(n714bar),
    .I1(n713bar)
  );
  //OR U248
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U248 (
    .O(n713),
    .I0(in[116]),
    .I1(in[110])
  );
  //AND U248bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U248bar (
    .O(n713bar),
    .I0(inbar[116]),
    .I1(inbar[110])
  );
  //OR U249
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U249 (
    .O(n714),
    .I0(in[133]),
    .I1(in[130])
  );
  //AND U249bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U249bar (
    .O(n714bar),
    .I0(inbar[133]),
    .I1(inbar[130])
  );
  //OR U250
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U250 (
    .O(n716),
    .I0(n712),
    .I1(n711)
  );
  //AND U250bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U250bar (
    .O(n716bar),
    .I0(n712bar),
    .I1(n711bar)
  );
  //OR U251
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U251 (
    .O(n711),
    .I0(in[203]),
    .I1(in[135])
  );
  //AND U251bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U251bar (
    .O(n711bar),
    .I0(inbar[203]),
    .I1(inbar[135])
  );
  //OR U252
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U252 (
    .O(n712),
    .I0(in[232]),
    .I1(in[223])
  );
  //AND U252bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U252bar (
    .O(n712bar),
    .I0(inbar[232]),
    .I1(inbar[223])
  );
  //OR U253
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U253 (
    .O(n718),
    .I0(n710),
    .I1(n709)
  );
  //AND U253bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U253bar (
    .O(n718bar),
    .I0(n710bar),
    .I1(n709bar)
  );
  //OR U254
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U254 (
    .O(n709),
    .I0(n708),
    .I1(n707)
  );
  //AND U254bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U254bar (
    .O(n709bar),
    .I0(n708bar),
    .I1(n707bar)
  );
  //OR U255
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U255 (
    .O(n707),
    .I0(in[255]),
    .I1(in[233])
  );
  //AND U255bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U255bar (
    .O(n707bar),
    .I0(inbar[255]),
    .I1(inbar[233])
  );
  //OR U256
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U256 (
    .O(n708),
    .I0(in_53),
    .I1(in_34)
  );
  //AND U256bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U256bar (
    .O(n708bar),
    .I0(in_53bar),
    .I1(in_34bar)
  );
  //OR U257
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U257 (
    .O(n710),
    .I0(n706),
    .I1(n705)
  );
  //AND U257bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U257bar (
    .O(n710bar),
    .I0(n706bar),
    .I1(n705bar)
  );
  //OR U258
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U258 (
    .O(n705),
    .I0(in_57),
    .I1(in_55)
  );
  //AND U258bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U258bar (
    .O(n705bar),
    .I0(in_57bar),
    .I1(in_55bar)
  );
  //OR U259
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U259 (
    .O(n706),
    .I0(in_68),
    .I1(in_67)
  );
  //AND U259bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U259bar (
    .O(n706bar),
    .I0(in_68bar),
    .I1(in_67bar)
  );
  //OR U260
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U260 (
    .O(n921),
    .I0(n704),
    .I1(n703)
  );
  //AND U260bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U260bar (
    .O(n921bar),
    .I0(n704bar),
    .I1(n703bar)
  );
  //OR U261
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U261 (
    .O(n703),
    .I0(n702),
    .I1(n701)
  );
  //AND U261bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U261bar (
    .O(n703bar),
    .I0(n702bar),
    .I1(n701bar)
  );
  //OR U262
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U262 (
    .O(n701),
    .I0(n700),
    .I1(n699)
  );
  //AND U262bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U262bar (
    .O(n701bar),
    .I0(n700bar),
    .I1(n699bar)
  );
  //OR U263
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U263 (
    .O(n699),
    .I0(n944),
    .I1(n872)
  );
  //AND U263bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U263bar (
    .O(n699bar),
    .I0(n944bar),
    .I1(n872bar)
  );
  //OR U264
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U264 (
    .O(n872),
    .I0(n698),
    .I1(n697)
  );
  //AND U264bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U264bar (
    .O(n872bar),
    .I0(n698bar),
    .I1(n697bar)
  );
  //OR U265
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U265 (
    .O(n697),
    .I0(n696),
    .I1(n695)
  );
  //AND U265bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U265bar (
    .O(n697bar),
    .I0(n696bar),
    .I1(n695bar)
  );
  //OR U266
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U266 (
    .O(n695),
    .I0(n694),
    .I1(n693)
  );
  //AND U266bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U266bar (
    .O(n695bar),
    .I0(n694bar),
    .I1(n693bar)
  );
  //OR U267
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U267 (
    .O(n693),
    .I0(in[121]),
    .I1(in[102])
  );
  //AND U267bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U267bar (
    .O(n693bar),
    .I0(inbar[121]),
    .I1(inbar[102])
  );
  //OR U268
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U268 (
    .O(n694),
    .I0(in[162]),
    .I1(in[161])
  );
  //AND U268bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U268bar (
    .O(n694bar),
    .I0(inbar[162]),
    .I1(inbar[161])
  );
  //OR U269
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U269 (
    .O(n696),
    .I0(n692),
    .I1(n691)
  );
  //AND U269bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U269bar (
    .O(n696bar),
    .I0(n692bar),
    .I1(n691bar)
  );
  //OR U270
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U270 (
    .O(n691),
    .I0(in[192]),
    .I1(in[178])
  );
  //AND U270bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U270bar (
    .O(n691bar),
    .I0(inbar[192]),
    .I1(inbar[178])
  );
  //OR U271
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U271 (
    .O(n692),
    .I0(in[244]),
    .I1(in[209])
  );
  //AND U271bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U271bar (
    .O(n692bar),
    .I0(inbar[244]),
    .I1(inbar[209])
  );
  //OR U272
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U272 (
    .O(n698),
    .I0(n690),
    .I1(n689)
  );
  //AND U272bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U272bar (
    .O(n698bar),
    .I0(n690bar),
    .I1(n689bar)
  );
  //OR U273
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U273 (
    .O(n689),
    .I0(n688),
    .I1(n687)
  );
  //AND U273bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U273bar (
    .O(n689bar),
    .I0(n688bar),
    .I1(n687bar)
  );
  //OR U274
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U274 (
    .O(n687),
    .I0(in[90]),
    .I1(in[254])
  );
  //AND U274bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U274bar (
    .O(n687bar),
    .I0(inbar[90]),
    .I1(inbar[254])
  );
  //OR U275
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U275 (
    .O(n688),
    .I0(in_36),
    .I1(in_32)
  );
  //AND U275bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U275bar (
    .O(n688bar),
    .I0(in_36bar),
    .I1(in_32bar)
  );
  //OR U276
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U276 (
    .O(n690),
    .I0(n686),
    .I1(n685)
  );
  //AND U276bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U276bar (
    .O(n690bar),
    .I0(n686bar),
    .I1(n685bar)
  );
  //OR U277
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U277 (
    .O(n685),
    .I0(in_62),
    .I1(in_37)
  );
  //AND U277bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U277bar (
    .O(n685bar),
    .I0(in_62bar),
    .I1(in_37bar)
  );
  //OR U278
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U278 (
    .O(n686),
    .I0(in_75),
    .I1(in_73)
  );
  //AND U278bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U278bar (
    .O(n686bar),
    .I0(in_75bar),
    .I1(in_73bar)
  );
  //OR U279
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U279 (
    .O(n944),
    .I0(n684),
    .I1(n683)
  );
  //AND U279bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U279bar (
    .O(n944bar),
    .I0(n684bar),
    .I1(n683bar)
  );
  //OR U280
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U280 (
    .O(n683),
    .I0(n682),
    .I1(n681)
  );
  //AND U280bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U280bar (
    .O(n683bar),
    .I0(n682bar),
    .I1(n681bar)
  );
  //OR U281
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U281 (
    .O(n681),
    .I0(n680),
    .I1(n679)
  );
  //AND U281bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U281bar (
    .O(n681bar),
    .I0(n680bar),
    .I1(n679bar)
  );
  //OR U282
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U282 (
    .O(n679),
    .I0(in[171]),
    .I1(in[153])
  );
  //AND U282bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U282bar (
    .O(n679bar),
    .I0(inbar[171]),
    .I1(inbar[153])
  );
  //OR U283
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U283 (
    .O(n680),
    .I0(in[187]),
    .I1(in[176])
  );
  //AND U283bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U283bar (
    .O(n680bar),
    .I0(inbar[187]),
    .I1(inbar[176])
  );
  //OR U284
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U284 (
    .O(n682),
    .I0(n678),
    .I1(n677)
  );
  //AND U284bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U284bar (
    .O(n682bar),
    .I0(n678bar),
    .I1(n677bar)
  );
  //OR U285
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U285 (
    .O(n677),
    .I0(in[245]),
    .I1(in[211])
  );
  //AND U285bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U285bar (
    .O(n677bar),
    .I0(inbar[245]),
    .I1(inbar[211])
  );
  //OR U286
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U286 (
    .O(n678),
    .I0(in[97]),
    .I1(in[88])
  );
  //AND U286bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U286bar (
    .O(n678bar),
    .I0(inbar[97]),
    .I1(inbar[88])
  );
  //OR U287
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U287 (
    .O(n684),
    .I0(n676),
    .I1(n675)
  );
  //AND U287bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U287bar (
    .O(n684bar),
    .I0(n676bar),
    .I1(n675bar)
  );
  //OR U288
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U288 (
    .O(n675),
    .I0(n674),
    .I1(n673)
  );
  //AND U288bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U288bar (
    .O(n675bar),
    .I0(n674bar),
    .I1(n673bar)
  );
  //OR U289
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U289 (
    .O(n673),
    .I0(in_10),
    .I1(in_0)
  );
  //AND U289bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U289bar (
    .O(n673bar),
    .I0(in_10bar),
    .I1(in_0bar)
  );
  //OR U290
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U290 (
    .O(n674),
    .I0(in_59),
    .I1(in_5)
  );
  //AND U290bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U290bar (
    .O(n674bar),
    .I0(in_59bar),
    .I1(in_5bar)
  );
  //OR U291
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U291 (
    .O(n676),
    .I0(n672),
    .I1(n671)
  );
  //AND U291bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U291bar (
    .O(n676bar),
    .I0(n672bar),
    .I1(n671bar)
  );
  //OR U292
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U292 (
    .O(n671),
    .I0(in_60),
    .I1(in_6)
  );
  //AND U292bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U292bar (
    .O(n671bar),
    .I0(in_60bar),
    .I1(in_6bar)
  );
  //OR U293
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U293 (
    .O(n672),
    .I0(in_77),
    .I1(in_69)
  );
  //AND U293bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U293bar (
    .O(n672bar),
    .I0(in_77bar),
    .I1(in_69bar)
  );
  //OR U294
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U294 (
    .O(n700),
    .I0(in[113]),
    .I1(n864)
  );
  //AND U294bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U294bar (
    .O(n700bar),
    .I0(inbar[113]),
    .I1(n864bar)
  );
  //OR U295
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U295 (
    .O(n864),
    .I0(n670),
    .I1(n669)
  );
  //AND U295bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U295bar (
    .O(n864bar),
    .I0(n670bar),
    .I1(n669bar)
  );
  //OR U296
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U296 (
    .O(n669),
    .I0(n668),
    .I1(n667)
  );
  //AND U296bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U296bar (
    .O(n669bar),
    .I0(n668bar),
    .I1(n667bar)
  );
  //OR U297
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U297 (
    .O(n667),
    .I0(n666),
    .I1(n665)
  );
  //AND U297bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U297bar (
    .O(n667bar),
    .I0(n666bar),
    .I1(n665bar)
  );
  //OR U298
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U298 (
    .O(n665),
    .I0(in[125]),
    .I1(in[107])
  );
  //AND U298bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U298bar (
    .O(n665bar),
    .I0(inbar[125]),
    .I1(inbar[107])
  );
  //OR U299
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U299 (
    .O(n666),
    .I0(in[138]),
    .I1(in[126])
  );
  //AND U299bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U299bar (
    .O(n666bar),
    .I0(inbar[138]),
    .I1(inbar[126])
  );
  //OR U300
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U300 (
    .O(n668),
    .I0(n664),
    .I1(n663)
  );
  //AND U300bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U300bar (
    .O(n668bar),
    .I0(n664bar),
    .I1(n663bar)
  );
  //OR U301
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U301 (
    .O(n663),
    .I0(in[189]),
    .I1(in[143])
  );
  //AND U301bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U301bar (
    .O(n663bar),
    .I0(inbar[189]),
    .I1(inbar[143])
  );
  //OR U302
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U302 (
    .O(n664),
    .I0(in[99]),
    .I1(in[214])
  );
  //AND U302bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U302bar (
    .O(n664bar),
    .I0(inbar[99]),
    .I1(inbar[214])
  );
  //OR U303
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U303 (
    .O(n670),
    .I0(n662),
    .I1(n661)
  );
  //AND U303bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U303bar (
    .O(n670bar),
    .I0(n662bar),
    .I1(n661bar)
  );
  //OR U304
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U304 (
    .O(n661),
    .I0(n660),
    .I1(n659)
  );
  //AND U304bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U304bar (
    .O(n661bar),
    .I0(n660bar),
    .I1(n659bar)
  );
  //OR U305
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U305 (
    .O(n659),
    .I0(in_15),
    .I1(in_12)
  );
  //AND U305bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U305bar (
    .O(n659bar),
    .I0(in_15bar),
    .I1(in_12bar)
  );
  //OR U306
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U306 (
    .O(n660),
    .I0(in_20),
    .I1(in_2)
  );
  //AND U306bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U306bar (
    .O(n660bar),
    .I0(in_20bar),
    .I1(in_2bar)
  );
  //OR U307
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U307 (
    .O(n662),
    .I0(n658),
    .I1(n657)
  );
  //AND U307bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U307bar (
    .O(n662bar),
    .I0(n658bar),
    .I1(n657bar)
  );
  //OR U308
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U308 (
    .O(n657),
    .I0(in_30),
    .I1(in_3)
  );
  //AND U308bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U308bar (
    .O(n657bar),
    .I0(in_30bar),
    .I1(in_3bar)
  );
  //OR U309
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U309 (
    .O(n658),
    .I0(in_4),
    .I1(in_38)
  );
  //AND U309bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U309bar (
    .O(n658bar),
    .I0(in_4bar),
    .I1(in_38bar)
  );
  //OR U310
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U310 (
    .O(n702),
    .I0(n656),
    .I1(n655)
  );
  //AND U310bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U310bar (
    .O(n702bar),
    .I0(n656bar),
    .I1(n655bar)
  );
  //OR U311
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U311 (
    .O(n655),
    .I0(in[148]),
    .I1(in[137])
  );
  //AND U311bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U311bar (
    .O(n655bar),
    .I0(inbar[148]),
    .I1(inbar[137])
  );
  //OR U312
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U312 (
    .O(n656),
    .I0(in[149]),
    .I1(n654)
  );
  //AND U312bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U312bar (
    .O(n656bar),
    .I0(inbar[149]),
    .I1(n654bar)
  );
  //OR U313
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U313 (
    .O(n654),
    .I0(in[195]),
    .I1(in[190])
  );
  //AND U313bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U313bar (
    .O(n654bar),
    .I0(inbar[195]),
    .I1(inbar[190])
  );
  //OR U314
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U314 (
    .O(n704),
    .I0(n653),
    .I1(n652)
  );
  //AND U314bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U314bar (
    .O(n704bar),
    .I0(n653bar),
    .I1(n652bar)
  );
  //OR U315
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U315 (
    .O(n652),
    .I0(n651),
    .I1(n650)
  );
  //AND U315bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U315bar (
    .O(n652bar),
    .I0(n651bar),
    .I1(n650bar)
  );
  //OR U316
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U316 (
    .O(n650),
    .I0(in[98]),
    .I1(in[197])
  );
  //AND U316bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U316bar (
    .O(n650bar),
    .I0(inbar[98]),
    .I1(inbar[197])
  );
  //OR U317
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U317 (
    .O(n651),
    .I0(in_11),
    .I1(n649)
  );
  //AND U317bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U317bar (
    .O(n651bar),
    .I0(in_11bar),
    .I1(n649bar)
  );
  //OR U318
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U318 (
    .O(n649),
    .I0(in_26),
    .I1(in_14)
  );
  //AND U318bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U318bar (
    .O(n649bar),
    .I0(in_26bar),
    .I1(in_14bar)
  );
  //OR U319
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U319 (
    .O(n653),
    .I0(n648),
    .I1(n647)
  );
  //AND U319bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U319bar (
    .O(n653bar),
    .I0(n648bar),
    .I1(n647bar)
  );
  //OR U320
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U320 (
    .O(n647),
    .I0(in_35),
    .I1(in_27)
  );
  //AND U320bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U320bar (
    .O(n647bar),
    .I0(in_35bar),
    .I1(in_27bar)
  );
  //OR U321
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U321 (
    .O(n648),
    .I0(in_50),
    .I1(n646)
  );
  //AND U321bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U321bar (
    .O(n648bar),
    .I0(in_50bar),
    .I1(n646bar)
  );
  //OR U322
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U322 (
    .O(n646),
    .I0(in_78),
    .I1(in_61)
  );
  //AND U322bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U322bar (
    .O(n646bar),
    .I0(in_78bar),
    .I1(in_61bar)
  );
  //OR U323
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U323 (
    .O(n720),
    .I0(n942),
    .I1(n645)
  );
  //AND U323bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U323bar (
    .O(n720bar),
    .I0(n942bar),
    .I1(n645bar)
  );
  //OR U324
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U324 (
    .O(n645),
    .I0(in[106]),
    .I1(n863)
  );
  //AND U324bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U324bar (
    .O(n645bar),
    .I0(inbar[106]),
    .I1(n863bar)
  );
  //OR U325
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U325 (
    .O(n863),
    .I0(n644),
    .I1(n643)
  );
  //AND U325bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U325bar (
    .O(n863bar),
    .I0(n644bar),
    .I1(n643bar)
  );
  //OR U326
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U326 (
    .O(n643),
    .I0(n642),
    .I1(n641)
  );
  //AND U326bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U326bar (
    .O(n643bar),
    .I0(n642bar),
    .I1(n641bar)
  );
  //OR U327
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U327 (
    .O(n641),
    .I0(n640),
    .I1(n639)
  );
  //AND U327bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U327bar (
    .O(n641bar),
    .I0(n640bar),
    .I1(n639bar)
  );
  //OR U328
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U328 (
    .O(n639),
    .I0(in[127]),
    .I1(in[122])
  );
  //AND U328bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U328bar (
    .O(n639bar),
    .I0(inbar[127]),
    .I1(inbar[122])
  );
  //OR U329
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U329 (
    .O(n640),
    .I0(in[156]),
    .I1(in[132])
  );
  //AND U329bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U329bar (
    .O(n640bar),
    .I0(inbar[156]),
    .I1(inbar[132])
  );
  //OR U330
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U330 (
    .O(n642),
    .I0(n638),
    .I1(n637)
  );
  //AND U330bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U330bar (
    .O(n642bar),
    .I0(n638bar),
    .I1(n637bar)
  );
  //OR U331
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U331 (
    .O(n637),
    .I0(in[159]),
    .I1(in[157])
  );
  //AND U331bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U331bar (
    .O(n637bar),
    .I0(inbar[159]),
    .I1(inbar[157])
  );
  //OR U332
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U332 (
    .O(n638),
    .I0(in[185]),
    .I1(in[169])
  );
  //AND U332bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U332bar (
    .O(n638bar),
    .I0(inbar[185]),
    .I1(inbar[169])
  );
  //OR U333
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U333 (
    .O(n644),
    .I0(n636),
    .I1(n635)
  );
  //AND U333bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U333bar (
    .O(n644bar),
    .I0(n636bar),
    .I1(n635bar)
  );
  //OR U334
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U334 (
    .O(n635),
    .I0(n634),
    .I1(n633)
  );
  //AND U334bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U334bar (
    .O(n635bar),
    .I0(n634bar),
    .I1(n633bar)
  );
  //OR U335
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U335 (
    .O(n633),
    .I0(in[239]),
    .I1(in[218])
  );
  //AND U335bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U335bar (
    .O(n633bar),
    .I0(inbar[239]),
    .I1(inbar[218])
  );
  //OR U336
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U336 (
    .O(n634),
    .I0(in_13),
    .I1(in[87])
  );
  //AND U336bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U336bar (
    .O(n634bar),
    .I0(in_13bar),
    .I1(inbar[87])
  );
  //OR U337
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U337 (
    .O(n636),
    .I0(n632),
    .I1(n631)
  );
  //AND U337bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U337bar (
    .O(n636bar),
    .I0(n632bar),
    .I1(n631bar)
  );
  //OR U338
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U338 (
    .O(n631),
    .I0(in_72),
    .I1(in_70)
  );
  //AND U338bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U338bar (
    .O(n631bar),
    .I0(in_72bar),
    .I1(in_70bar)
  );
  //OR U339
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U339 (
    .O(n632),
    .I0(in_80),
    .I1(in_74)
  );
  //AND U339bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U339bar (
    .O(n632bar),
    .I0(in_80bar),
    .I1(in_74bar)
  );
  //OR U340
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U340 (
    .O(n942),
    .I0(n630),
    .I1(n629)
  );
  //AND U340bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U340bar (
    .O(n942bar),
    .I0(n630bar),
    .I1(n629bar)
  );
  //OR U341
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U341 (
    .O(n629),
    .I0(n628),
    .I1(n627)
  );
  //AND U341bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U341bar (
    .O(n629bar),
    .I0(n628bar),
    .I1(n627bar)
  );
  //OR U342
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U342 (
    .O(n627),
    .I0(n626),
    .I1(n625)
  );
  //AND U342bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U342bar (
    .O(n627bar),
    .I0(n626bar),
    .I1(n625bar)
  );
  //OR U343
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U343 (
    .O(n625),
    .I0(in[146]),
    .I1(in[100])
  );
  //AND U343bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U343bar (
    .O(n625bar),
    .I0(inbar[146]),
    .I1(inbar[100])
  );
  //OR U344
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U344 (
    .O(n626),
    .I0(in[168]),
    .I1(in[152])
  );
  //AND U344bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U344bar (
    .O(n626bar),
    .I0(inbar[168]),
    .I1(inbar[152])
  );
  //OR U345
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U345 (
    .O(n628),
    .I0(n624),
    .I1(n623)
  );
  //AND U345bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U345bar (
    .O(n628bar),
    .I0(n624bar),
    .I1(n623bar)
  );
  //OR U346
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U346 (
    .O(n623),
    .I0(in[199]),
    .I1(in[182])
  );
  //AND U346bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U346bar (
    .O(n623bar),
    .I0(inbar[199]),
    .I1(inbar[182])
  );
  //OR U347
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U347 (
    .O(n624),
    .I0(in[236]),
    .I1(in[204])
  );
  //AND U347bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U347bar (
    .O(n624bar),
    .I0(inbar[236]),
    .I1(inbar[204])
  );
  //OR U348
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U348 (
    .O(n630),
    .I0(n622),
    .I1(n621)
  );
  //AND U348bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U348bar (
    .O(n630bar),
    .I0(n622bar),
    .I1(n621bar)
  );
  //OR U349
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U349 (
    .O(n621),
    .I0(n620),
    .I1(n619)
  );
  //AND U349bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U349bar (
    .O(n621bar),
    .I0(n620bar),
    .I1(n619bar)
  );
  //OR U350
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U350 (
    .O(n619),
    .I0(in[89]),
    .I1(in[246])
  );
  //AND U350bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U350bar (
    .O(n619bar),
    .I0(inbar[89]),
    .I1(inbar[246])
  );
  //OR U351
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U351 (
    .O(n620),
    .I0(in[95]),
    .I1(in[92])
  );
  //AND U351bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U351bar (
    .O(n620bar),
    .I0(inbar[95]),
    .I1(inbar[92])
  );
  //OR U352
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U352 (
    .O(n622),
    .I0(n618),
    .I1(n617)
  );
  //AND U352bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U352bar (
    .O(n622bar),
    .I0(n618bar),
    .I1(n617bar)
  );
  //OR U353
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U353 (
    .O(n617),
    .I0(in_22),
    .I1(in_16)
  );
  //AND U353bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U353bar (
    .O(n617bar),
    .I0(in_22bar),
    .I1(in_16bar)
  );
  //OR U354
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U354 (
    .O(n618),
    .I0(in_51),
    .I1(in_49)
  );
  //AND U354bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U354bar (
    .O(n618bar),
    .I0(in_51bar),
    .I1(in_49bar)
  );
  //OR U355
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U355 (
    .O(n722),
    .I0(n616),
    .I1(n615)
  );
  //AND U355bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U355bar (
    .O(n722bar),
    .I0(n616bar),
    .I1(n615bar)
  );
  //OR U356
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U356 (
    .O(n615),
    .I0(in[158]),
    .I1(in[115])
  );
  //AND U356bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U356bar (
    .O(n615bar),
    .I0(inbar[158]),
    .I1(inbar[115])
  );
  //OR U357
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U357 (
    .O(n616),
    .I0(in[163]),
    .I1(n614)
  );
  //AND U357bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U357bar (
    .O(n616bar),
    .I0(inbar[163]),
    .I1(n614bar)
  );
  //OR U358
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U358 (
    .O(n614),
    .I0(in[206]),
    .I1(in[165])
  );
  //AND U358bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U358bar (
    .O(n614bar),
    .I0(inbar[206]),
    .I1(inbar[165])
  );
  //OR U359
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U359 (
    .O(n724),
    .I0(n613),
    .I1(n612)
  );
  //AND U359bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U359bar (
    .O(n724bar),
    .I0(n613bar),
    .I1(n612bar)
  );
  //OR U360
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U360 (
    .O(n612),
    .I0(n611),
    .I1(n610)
  );
  //AND U360bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U360bar (
    .O(n612bar),
    .I0(n611bar),
    .I1(n610bar)
  );
  //OR U361
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U361 (
    .O(n610),
    .I0(in[213]),
    .I1(in[207])
  );
  //AND U361bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U361bar (
    .O(n610bar),
    .I0(inbar[213]),
    .I1(inbar[207])
  );
  //OR U362
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U362 (
    .O(n611),
    .I0(in[215]),
    .I1(n609)
  );
  //AND U362bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U362bar (
    .O(n611bar),
    .I0(inbar[215]),
    .I1(n609bar)
  );
  //OR U363
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U363 (
    .O(n609),
    .I0(in[230]),
    .I1(in[220])
  );
  //AND U363bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U363bar (
    .O(n609bar),
    .I0(inbar[230]),
    .I1(inbar[220])
  );
  //OR U364
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U364 (
    .O(n613),
    .I0(n608),
    .I1(n607)
  );
  //AND U364bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U364bar (
    .O(n613bar),
    .I0(n608bar),
    .I1(n607bar)
  );
  //OR U365
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U365 (
    .O(n607),
    .I0(in[251]),
    .I1(in[234])
  );
  //AND U365bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U365bar (
    .O(n607bar),
    .I0(inbar[251]),
    .I1(inbar[234])
  );
  //OR U366
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U366 (
    .O(n608),
    .I0(in_17),
    .I1(n606)
  );
  //AND U366bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U366bar (
    .O(n608bar),
    .I0(in_17bar),
    .I1(n606bar)
  );
  //OR U367
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U367 (
    .O(n606),
    .I0(in_65),
    .I1(in_56)
  );
  //AND U367bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U367bar (
    .O(n606bar),
    .I0(in_65bar),
    .I1(in_56bar)
  );
  //OR U368
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U368 (
    .O(out[0]),
    .I0(n605),
    .I1(n604)
  );
  //AND U368bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U368bar (
    .O(outbar[0]),
    .I0(n605bar),
    .I1(n604bar)
  );
  //OR U369
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U369 (
    .O(n604),
    .I0(n603),
    .I1(n602)
  );
  //AND U369bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U369bar (
    .O(n604bar),
    .I0(n603bar),
    .I1(n602bar)
  );
  //OR U370
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U370 (
    .O(n602),
    .I0(n601),
    .I1(n600)
  );
  //AND U370bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U370bar (
    .O(n602bar),
    .I0(n601bar),
    .I1(n600bar)
  );
  //OR U371
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U371 (
    .O(n600),
    .I0(n820),
    .I1(n785)
  );
  //AND U371bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U371bar (
    .O(n600bar),
    .I0(n820bar),
    .I1(n785bar)
  );
  //OR U372
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U372 (
    .O(n785),
    .I0(n599),
    .I1(n598)
  );
  //AND U372bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U372bar (
    .O(n785bar),
    .I0(n599bar),
    .I1(n598bar)
  );
  //OR U373
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U373 (
    .O(n598),
    .I0(n597),
    .I1(n596)
  );
  //AND U373bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U373bar (
    .O(n598bar),
    .I0(n597bar),
    .I1(n596bar)
  );
  //OR U374
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U374 (
    .O(n596),
    .I0(n595),
    .I1(n594)
  );
  //AND U374bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U374bar (
    .O(n596bar),
    .I0(n595bar),
    .I1(n594bar)
  );
  //OR U375
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U375 (
    .O(n594),
    .I0(in[135]),
    .I1(in[104])
  );
  //AND U375bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U375bar (
    .O(n594bar),
    .I0(inbar[135]),
    .I1(inbar[104])
  );
  //OR U376
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U376 (
    .O(n595),
    .I0(in[188]),
    .I1(in[178])
  );
  //AND U376bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U376bar (
    .O(n595bar),
    .I0(inbar[188]),
    .I1(inbar[178])
  );
  //OR U377
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U377 (
    .O(n597),
    .I0(n593),
    .I1(n592)
  );
  //AND U377bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U377bar (
    .O(n597bar),
    .I0(n593bar),
    .I1(n592bar)
  );
  //OR U378
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U378 (
    .O(n592),
    .I0(in[217]),
    .I1(in[194])
  );
  //AND U378bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U378bar (
    .O(n592bar),
    .I0(inbar[217]),
    .I1(inbar[194])
  );
  //OR U379
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U379 (
    .O(n593),
    .I0(in[237]),
    .I1(in[218])
  );
  //AND U379bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U379bar (
    .O(n593bar),
    .I0(inbar[237]),
    .I1(inbar[218])
  );
  //OR U380
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U380 (
    .O(n599),
    .I0(n591),
    .I1(n590)
  );
  //AND U380bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U380bar (
    .O(n599bar),
    .I0(n591bar),
    .I1(n590bar)
  );
  //OR U381
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U381 (
    .O(n590),
    .I0(n589),
    .I1(n588)
  );
  //AND U381bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U381bar (
    .O(n590bar),
    .I0(n589bar),
    .I1(n588bar)
  );
  //OR U382
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U382 (
    .O(n588),
    .I0(in_2),
    .I1(in_10)
  );
  //AND U382bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U382bar (
    .O(n588bar),
    .I0(in_2bar),
    .I1(in_10bar)
  );
  //OR U383
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U383 (
    .O(n589),
    .I0(in_47),
    .I1(in_22)
  );
  //AND U383bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U383bar (
    .O(n589bar),
    .I0(in_47bar),
    .I1(in_22bar)
  );
  //OR U384
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U384 (
    .O(n591),
    .I0(n587),
    .I1(n586)
  );
  //AND U384bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U384bar (
    .O(n591bar),
    .I0(n587bar),
    .I1(n586bar)
  );
  //OR U385
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U385 (
    .O(n586),
    .I0(in_56),
    .I1(in_54)
  );
  //AND U385bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U385bar (
    .O(n586bar),
    .I0(in_56bar),
    .I1(in_54bar)
  );
  //OR U386
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U386 (
    .O(n587),
    .I0(in_63),
    .I1(in_61)
  );
  //AND U386bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U386bar (
    .O(n587bar),
    .I0(in_63bar),
    .I1(in_61bar)
  );
  //OR U387
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U387 (
    .O(n820),
    .I0(n585),
    .I1(n584)
  );
  //AND U387bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U387bar (
    .O(n820bar),
    .I0(n585bar),
    .I1(n584bar)
  );
  //OR U388
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U388 (
    .O(n584),
    .I0(n583),
    .I1(n582)
  );
  //AND U388bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U388bar (
    .O(n584bar),
    .I0(n583bar),
    .I1(n582bar)
  );
  //OR U389
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U389 (
    .O(n582),
    .I0(n581),
    .I1(n580)
  );
  //AND U389bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U389bar (
    .O(n582bar),
    .I0(n581bar),
    .I1(n580bar)
  );
  //OR U390
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U390 (
    .O(n580),
    .I0(in[158]),
    .I1(in[142])
  );
  //AND U390bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U390bar (
    .O(n580bar),
    .I0(inbar[158]),
    .I1(inbar[142])
  );
  //OR U391
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U391 (
    .O(n581),
    .I0(in[175]),
    .I1(in[164])
  );
  //AND U391bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U391bar (
    .O(n581bar),
    .I0(inbar[175]),
    .I1(inbar[164])
  );
  //OR U392
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U392 (
    .O(n583),
    .I0(n579),
    .I1(n578)
  );
  //AND U392bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U392bar (
    .O(n583bar),
    .I0(n579bar),
    .I1(n578bar)
  );
  //OR U393
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U393 (
    .O(n578),
    .I0(in[228]),
    .I1(in[204])
  );
  //AND U393bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U393bar (
    .O(n578bar),
    .I0(inbar[228]),
    .I1(inbar[204])
  );
  //OR U394
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U394 (
    .O(n579),
    .I0(in[91]),
    .I1(in[87])
  );
  //AND U394bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U394bar (
    .O(n579bar),
    .I0(inbar[91]),
    .I1(inbar[87])
  );
  //OR U395
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U395 (
    .O(n585),
    .I0(n577),
    .I1(n576)
  );
  //AND U395bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U395bar (
    .O(n585bar),
    .I0(n577bar),
    .I1(n576bar)
  );
  //OR U396
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U396 (
    .O(n576),
    .I0(n575),
    .I1(n574)
  );
  //AND U396bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U396bar (
    .O(n576bar),
    .I0(n575bar),
    .I1(n574bar)
  );
  //OR U397
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U397 (
    .O(n574),
    .I0(in_21),
    .I1(in_11)
  );
  //AND U397bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U397bar (
    .O(n574bar),
    .I0(in_21bar),
    .I1(in_11bar)
  );
  //OR U398
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U398 (
    .O(n575),
    .I0(in_5),
    .I1(in_3)
  );
  //AND U398bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U398bar (
    .O(n575bar),
    .I0(in_5bar),
    .I1(in_3bar)
  );
  //OR U399
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U399 (
    .O(n577),
    .I0(n573),
    .I1(n572)
  );
  //AND U399bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U399bar (
    .O(n577bar),
    .I0(n573bar),
    .I1(n572bar)
  );
  //OR U400
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U400 (
    .O(n572),
    .I0(in_68),
    .I1(in_64)
  );
  //AND U400bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U400bar (
    .O(n572bar),
    .I0(in_68bar),
    .I1(in_64bar)
  );
  //OR U401
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U401 (
    .O(n573),
    .I0(in_76),
    .I1(in_73)
  );
  //AND U401bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U401bar (
    .O(n573bar),
    .I0(in_76bar),
    .I1(in_73bar)
  );
  //OR U402
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U402 (
    .O(n601),
    .I0(n778),
    .I1(n571)
  );
  //AND U402bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U402bar (
    .O(n601bar),
    .I0(n778bar),
    .I1(n571bar)
  );
  //OR U403
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U403 (
    .O(n571),
    .I0(in[100]),
    .I1(n965)
  );
  //AND U403bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U403bar (
    .O(n571bar),
    .I0(inbar[100]),
    .I1(n965bar)
  );
  //OR U404
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U404 (
    .O(n965),
    .I0(n570),
    .I1(n569)
  );
  //AND U404bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U404bar (
    .O(n965bar),
    .I0(n570bar),
    .I1(n569bar)
  );
  //OR U405
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U405 (
    .O(n569),
    .I0(n568),
    .I1(n567)
  );
  //AND U405bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U405bar (
    .O(n569bar),
    .I0(n568bar),
    .I1(n567bar)
  );
  //OR U406
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U406 (
    .O(n567),
    .I0(n566),
    .I1(n565)
  );
  //AND U406bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U406bar (
    .O(n567bar),
    .I0(n566bar),
    .I1(n565bar)
  );
  //OR U407
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U407 (
    .O(n565),
    .I0(n817),
    .I1(n750)
  );
  //AND U407bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U407bar (
    .O(n565bar),
    .I0(n817bar),
    .I1(n750bar)
  );
  //OR U408
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U408 (
    .O(n750),
    .I0(n564),
    .I1(n563)
  );
  //AND U408bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U408bar (
    .O(n750bar),
    .I0(n564bar),
    .I1(n563bar)
  );
  //OR U409
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U409 (
    .O(n563),
    .I0(n562),
    .I1(n561)
  );
  //AND U409bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U409bar (
    .O(n563bar),
    .I0(n562bar),
    .I1(n561bar)
  );
  //OR U410
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U410 (
    .O(n561),
    .I0(n560),
    .I1(n559)
  );
  //AND U410bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U410bar (
    .O(n561bar),
    .I0(n560bar),
    .I1(n559bar)
  );
  //OR U411
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U411 (
    .O(n559),
    .I0(in[119]),
    .I1(in[103])
  );
  //AND U411bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U411bar (
    .O(n559bar),
    .I0(inbar[119]),
    .I1(inbar[103])
  );
  //OR U412
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U412 (
    .O(n560),
    .I0(in[137]),
    .I1(in[133])
  );
  //AND U412bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U412bar (
    .O(n560bar),
    .I0(inbar[137]),
    .I1(inbar[133])
  );
  //OR U413
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U413 (
    .O(n562),
    .I0(n558),
    .I1(n557)
  );
  //AND U413bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U413bar (
    .O(n562bar),
    .I0(n558bar),
    .I1(n557bar)
  );
  //OR U414
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U414 (
    .O(n557),
    .I0(in[176]),
    .I1(in[173])
  );
  //AND U414bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U414bar (
    .O(n557bar),
    .I0(inbar[176]),
    .I1(inbar[173])
  );
  //OR U415
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U415 (
    .O(n558),
    .I0(in[210]),
    .I1(in[181])
  );
  //AND U415bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U415bar (
    .O(n558bar),
    .I0(inbar[210]),
    .I1(inbar[181])
  );
  //OR U416
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U416 (
    .O(n564),
    .I0(n556),
    .I1(n555)
  );
  //AND U416bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U416bar (
    .O(n564bar),
    .I0(n556bar),
    .I1(n555bar)
  );
  //OR U417
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U417 (
    .O(n555),
    .I0(n554),
    .I1(n553)
  );
  //AND U417bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U417bar (
    .O(n555bar),
    .I0(n554bar),
    .I1(n553bar)
  );
  //OR U418
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U418 (
    .O(n553),
    .I0(in_13),
    .I1(in[234])
  );
  //AND U418bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U418bar (
    .O(n553bar),
    .I0(in_13bar),
    .I1(inbar[234])
  );
  //OR U419
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U419 (
    .O(n554),
    .I0(in_38),
    .I1(in_32)
  );
  //AND U419bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U419bar (
    .O(n554bar),
    .I0(in_38bar),
    .I1(in_32bar)
  );
  //OR U420
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U420 (
    .O(n556),
    .I0(n552),
    .I1(n551)
  );
  //AND U420bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U420bar (
    .O(n556bar),
    .I0(n552bar),
    .I1(n551bar)
  );
  //OR U421
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U421 (
    .O(n551),
    .I0(in_42),
    .I1(in_41)
  );
  //AND U421bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U421bar (
    .O(n551bar),
    .I0(in_42bar),
    .I1(in_41bar)
  );
  //OR U422
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U422 (
    .O(n552),
    .I0(in_7),
    .I1(in_49)
  );
  //AND U422bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U422bar (
    .O(n552bar),
    .I0(in_7bar),
    .I1(in_49bar)
  );
  //OR U423
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U423 (
    .O(n817),
    .I0(n550),
    .I1(n549)
  );
  //AND U423bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U423bar (
    .O(n817bar),
    .I0(n550bar),
    .I1(n549bar)
  );
  //OR U424
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U424 (
    .O(n549),
    .I0(n548),
    .I1(n547)
  );
  //AND U424bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U424bar (
    .O(n549bar),
    .I0(n548bar),
    .I1(n547bar)
  );
  //OR U425
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U425 (
    .O(n547),
    .I0(n546),
    .I1(n545)
  );
  //AND U425bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U425bar (
    .O(n547bar),
    .I0(n546bar),
    .I1(n545bar)
  );
  //OR U426
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U426 (
    .O(n545),
    .I0(in[159]),
    .I1(in[105])
  );
  //AND U426bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U426bar (
    .O(n545bar),
    .I0(inbar[159]),
    .I1(inbar[105])
  );
  //OR U427
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U427 (
    .O(n546),
    .I0(in[206]),
    .I1(in[183])
  );
  //AND U427bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U427bar (
    .O(n546bar),
    .I0(inbar[206]),
    .I1(inbar[183])
  );
  //OR U428
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U428 (
    .O(n548),
    .I0(n544),
    .I1(n543)
  );
  //AND U428bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U428bar (
    .O(n548bar),
    .I0(n544bar),
    .I1(n543bar)
  );
  //OR U429
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U429 (
    .O(n543),
    .I0(in[229]),
    .I1(in[219])
  );
  //AND U429bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U429bar (
    .O(n543bar),
    .I0(inbar[229]),
    .I1(inbar[219])
  );
  //OR U430
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U430 (
    .O(n544),
    .I0(in[235]),
    .I1(in[232])
  );
  //AND U430bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U430bar (
    .O(n544bar),
    .I0(inbar[235]),
    .I1(inbar[232])
  );
  //OR U431
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U431 (
    .O(n550),
    .I0(n542),
    .I1(n541)
  );
  //AND U431bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U431bar (
    .O(n550bar),
    .I0(n542bar),
    .I1(n541bar)
  );
  //OR U432
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U432 (
    .O(n541),
    .I0(n540),
    .I1(n539)
  );
  //AND U432bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U432bar (
    .O(n541bar),
    .I0(n540bar),
    .I1(n539bar)
  );
  //OR U433
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U433 (
    .O(n539),
    .I0(in[249]),
    .I1(in[242])
  );
  //AND U433bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U433bar (
    .O(n539bar),
    .I0(inbar[249]),
    .I1(inbar[242])
  );
  //OR U434
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U434 (
    .O(n540),
    .I0(in[89]),
    .I1(in[254])
  );
  //AND U434bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U434bar (
    .O(n540bar),
    .I0(inbar[89]),
    .I1(inbar[254])
  );
  //OR U435
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U435 (
    .O(n542),
    .I0(n538),
    .I1(n537)
  );
  //AND U435bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U435bar (
    .O(n542bar),
    .I0(n538bar),
    .I1(n537bar)
  );
  //OR U436
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U436 (
    .O(n537),
    .I0(in_14),
    .I1(in[99])
  );
  //AND U436bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U436bar (
    .O(n537bar),
    .I0(in_14bar),
    .I1(inbar[99])
  );
  //OR U437
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U437 (
    .O(n538),
    .I0(in_60),
    .I1(in_18)
  );
  //AND U437bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U437bar (
    .O(n538bar),
    .I0(in_60bar),
    .I1(in_18bar)
  );
  //OR U438
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U438 (
    .O(n566),
    .I0(in[113]),
    .I1(n763)
  );
  //AND U438bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U438bar (
    .O(n566bar),
    .I0(inbar[113]),
    .I1(n763bar)
  );
  //OR U439
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U439 (
    .O(n763),
    .I0(n536),
    .I1(n535)
  );
  //AND U439bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U439bar (
    .O(n763bar),
    .I0(n536bar),
    .I1(n535bar)
  );
  //OR U440
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U440 (
    .O(n535),
    .I0(n534),
    .I1(n533)
  );
  //AND U440bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U440bar (
    .O(n535bar),
    .I0(n534bar),
    .I1(n533bar)
  );
  //OR U441
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U441 (
    .O(n533),
    .I0(n532),
    .I1(n531)
  );
  //AND U441bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U441bar (
    .O(n533bar),
    .I0(n532bar),
    .I1(n531bar)
  );
  //OR U442
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U442 (
    .O(n531),
    .I0(in[115]),
    .I1(in[110])
  );
  //AND U442bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U442bar (
    .O(n531bar),
    .I0(inbar[115]),
    .I1(inbar[110])
  );
  //OR U443
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U443 (
    .O(n532),
    .I0(in[125]),
    .I1(in[117])
  );
  //AND U443bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U443bar (
    .O(n532bar),
    .I0(inbar[125]),
    .I1(inbar[117])
  );
  //OR U444
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U444 (
    .O(n534),
    .I0(n530),
    .I1(n529)
  );
  //AND U444bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U444bar (
    .O(n534bar),
    .I0(n530bar),
    .I1(n529bar)
  );
  //OR U445
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U445 (
    .O(n529),
    .I0(in[180]),
    .I1(in[128])
  );
  //AND U445bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U445bar (
    .O(n529bar),
    .I0(inbar[180]),
    .I1(inbar[128])
  );
  //OR U446
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U446 (
    .O(n530),
    .I0(in[205]),
    .I1(in[201])
  );
  //AND U446bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U446bar (
    .O(n530bar),
    .I0(inbar[205]),
    .I1(inbar[201])
  );
  //OR U447
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U447 (
    .O(n536),
    .I0(n528),
    .I1(n527)
  );
  //AND U447bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U447bar (
    .O(n536bar),
    .I0(n528bar),
    .I1(n527bar)
  );
  //OR U448
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U448 (
    .O(n527),
    .I0(n526),
    .I1(n525)
  );
  //AND U448bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U448bar (
    .O(n527bar),
    .I0(n526bar),
    .I1(n525bar)
  );
  //OR U449
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U449 (
    .O(n525),
    .I0(in[244]),
    .I1(in[239])
  );
  //AND U449bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U449bar (
    .O(n525bar),
    .I0(inbar[244]),
    .I1(inbar[239])
  );
  //OR U450
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U450 (
    .O(n526),
    .I0(in[95]),
    .I1(in[83])
  );
  //AND U450bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U450bar (
    .O(n526bar),
    .I0(inbar[95]),
    .I1(inbar[83])
  );
  //OR U451
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U451 (
    .O(n528),
    .I0(n524),
    .I1(n523)
  );
  //AND U451bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U451bar (
    .O(n528bar),
    .I0(n524bar),
    .I1(n523bar)
  );
  //OR U452
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U452 (
    .O(n523),
    .I0(in_24),
    .I1(in[97])
  );
  //AND U452bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U452bar (
    .O(n523bar),
    .I0(in_24bar),
    .I1(inbar[97])
  );
  //OR U453
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U453 (
    .O(n524),
    .I0(in_33),
    .I1(in_27)
  );
  //AND U453bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U453bar (
    .O(n524bar),
    .I0(in_33bar),
    .I1(in_27bar)
  );
  //OR U454
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U454 (
    .O(n568),
    .I0(n522),
    .I1(n521)
  );
  //AND U454bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U454bar (
    .O(n568bar),
    .I0(n522bar),
    .I1(n521bar)
  );
  //OR U455
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U455 (
    .O(n521),
    .I0(in[145]),
    .I1(in[126])
  );
  //AND U455bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U455bar (
    .O(n521bar),
    .I0(inbar[145]),
    .I1(inbar[126])
  );
  //OR U456
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U456 (
    .O(n522),
    .I0(in[169]),
    .I1(n520)
  );
  //AND U456bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U456bar (
    .O(n522bar),
    .I0(inbar[169]),
    .I1(n520bar)
  );
  //OR U457
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U457 (
    .O(n520),
    .I0(in[221]),
    .I1(in[172])
  );
  //AND U457bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U457bar (
    .O(n520bar),
    .I0(inbar[221]),
    .I1(inbar[172])
  );
  //OR U458
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U458 (
    .O(n570),
    .I0(n519),
    .I1(n518)
  );
  //AND U458bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U458bar (
    .O(n570bar),
    .I0(n519bar),
    .I1(n518bar)
  );
  //OR U459
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U459 (
    .O(n518),
    .I0(n517),
    .I1(n516)
  );
  //AND U459bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U459bar (
    .O(n518bar),
    .I0(n517bar),
    .I1(n516bar)
  );
  //OR U460
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U460 (
    .O(n516),
    .I0(in[241]),
    .I1(in[224])
  );
  //AND U460bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U460bar (
    .O(n516bar),
    .I0(inbar[241]),
    .I1(inbar[224])
  );
  //OR U461
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U461 (
    .O(n517),
    .I0(in[86]),
    .I1(n515)
  );
  //AND U461bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U461bar (
    .O(n517bar),
    .I0(inbar[86]),
    .I1(n515bar)
  );
  //OR U462
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U462 (
    .O(n515),
    .I0(in_43),
    .I1(in_34)
  );
  //AND U462bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U462bar (
    .O(n515bar),
    .I0(in_43bar),
    .I1(in_34bar)
  );
  //OR U463
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U463 (
    .O(n519),
    .I0(n514),
    .I1(n513)
  );
  //AND U463bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U463bar (
    .O(n519bar),
    .I0(n514bar),
    .I1(n513bar)
  );
  //OR U464
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U464 (
    .O(n513),
    .I0(in_65),
    .I1(in_51)
  );
  //AND U464bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U464bar (
    .O(n513bar),
    .I0(in_65bar),
    .I1(in_51bar)
  );
  //OR U465
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U465 (
    .O(n514),
    .I0(in_75),
    .I1(n512)
  );
  //AND U465bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U465bar (
    .O(n514bar),
    .I0(in_75bar),
    .I1(n512bar)
  );
  //OR U466
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U466 (
    .O(n512),
    .I0(in_81),
    .I1(in_77)
  );
  //AND U466bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U466bar (
    .O(n512bar),
    .I0(in_81bar),
    .I1(in_77bar)
  );
  //OR U467
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U467 (
    .O(n778),
    .I0(n511),
    .I1(n510)
  );
  //AND U467bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U467bar (
    .O(n778bar),
    .I0(n511bar),
    .I1(n510bar)
  );
  //OR U468
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U468 (
    .O(n510),
    .I0(n509),
    .I1(n508)
  );
  //AND U468bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U468bar (
    .O(n510bar),
    .I0(n509bar),
    .I1(n508bar)
  );
  //OR U469
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U469 (
    .O(n508),
    .I0(n507),
    .I1(n506)
  );
  //AND U469bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U469bar (
    .O(n508bar),
    .I0(n507bar),
    .I1(n506bar)
  );
  //OR U470
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U470 (
    .O(n506),
    .I0(in[107]),
    .I1(in[101])
  );
  //AND U470bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U470bar (
    .O(n506bar),
    .I0(inbar[107]),
    .I1(inbar[101])
  );
  //OR U471
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U471 (
    .O(n507),
    .I0(in[139]),
    .I1(in[132])
  );
  //AND U471bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U471bar (
    .O(n507bar),
    .I0(inbar[139]),
    .I1(inbar[132])
  );
  //OR U472
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U472 (
    .O(n509),
    .I0(n505),
    .I1(n504)
  );
  //AND U472bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U472bar (
    .O(n509bar),
    .I0(n505bar),
    .I1(n504bar)
  );
  //OR U473
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U473 (
    .O(n504),
    .I0(in[146]),
    .I1(in[141])
  );
  //AND U473bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U473bar (
    .O(n504bar),
    .I0(inbar[146]),
    .I1(inbar[141])
  );
  //OR U474
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U474 (
    .O(n505),
    .I0(in[203]),
    .I1(in[179])
  );
  //AND U474bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U474bar (
    .O(n505bar),
    .I0(inbar[203]),
    .I1(inbar[179])
  );
  //OR U475
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U475 (
    .O(n511),
    .I0(n503),
    .I1(n502)
  );
  //AND U475bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U475bar (
    .O(n511bar),
    .I0(n503bar),
    .I1(n502bar)
  );
  //OR U476
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U476 (
    .O(n502),
    .I0(n501),
    .I1(n500)
  );
  //AND U476bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U476bar (
    .O(n502bar),
    .I0(n501bar),
    .I1(n500bar)
  );
  //OR U477
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U477 (
    .O(n500),
    .I0(in[243]),
    .I1(in[222])
  );
  //AND U477bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U477bar (
    .O(n500bar),
    .I0(inbar[243]),
    .I1(inbar[222])
  );
  //OR U478
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U478 (
    .O(n501),
    .I0(in[251]),
    .I1(in[250])
  );
  //AND U478bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U478bar (
    .O(n501bar),
    .I0(inbar[251]),
    .I1(inbar[250])
  );
  //OR U479
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U479 (
    .O(n503),
    .I0(n499),
    .I1(n498)
  );
  //AND U479bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U479bar (
    .O(n503bar),
    .I0(n499bar),
    .I1(n498bar)
  );
  //OR U480
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U480 (
    .O(n498),
    .I0(in_37),
    .I1(in_19)
  );
  //AND U480bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U480bar (
    .O(n498bar),
    .I0(in_37bar),
    .I1(in_19bar)
  );
  //OR U481
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U481 (
    .O(n499),
    .I0(in_78),
    .I1(in_6)
  );
  //AND U481bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U481bar (
    .O(n499bar),
    .I0(in_78bar),
    .I1(in_6bar)
  );
  //OR U482
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U482 (
    .O(n603),
    .I0(n497),
    .I1(n496)
  );
  //AND U482bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U482bar (
    .O(n603bar),
    .I0(n497bar),
    .I1(n496bar)
  );
  //OR U483
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U483 (
    .O(n496),
    .I0(in[112]),
    .I1(in[102])
  );
  //AND U483bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U483bar (
    .O(n496bar),
    .I0(inbar[112]),
    .I1(inbar[102])
  );
  //OR U484
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U484 (
    .O(n497),
    .I0(in[123]),
    .I1(n495)
  );
  //AND U484bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U484bar (
    .O(n497bar),
    .I0(inbar[123]),
    .I1(n495bar)
  );
  //OR U485
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U485 (
    .O(n495),
    .I0(in[143]),
    .I1(in[130])
  );
  //AND U485bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U485bar (
    .O(n495bar),
    .I0(inbar[143]),
    .I1(inbar[130])
  );
  //OR U486
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U486 (
    .O(n605),
    .I0(n494),
    .I1(n493)
  );
  //AND U486bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U486bar (
    .O(n605bar),
    .I0(n494bar),
    .I1(n493bar)
  );
  //OR U487
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U487 (
    .O(n493),
    .I0(n492),
    .I1(n491)
  );
  //AND U487bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U487bar (
    .O(n493bar),
    .I0(n492bar),
    .I1(n491bar)
  );
  //OR U488
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U488 (
    .O(n491),
    .I0(in[216]),
    .I1(in[213])
  );
  //AND U488bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U488bar (
    .O(n491bar),
    .I0(inbar[216]),
    .I1(inbar[213])
  );
  //OR U489
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U489 (
    .O(n492),
    .I0(in[227]),
    .I1(n490)
  );
  //AND U489bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U489bar (
    .O(n492bar),
    .I0(inbar[227]),
    .I1(n490bar)
  );
  //OR U490
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U490 (
    .O(n490),
    .I0(in_0),
    .I1(in[248])
  );
  //AND U490bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U490bar (
    .O(n490bar),
    .I0(in_0bar),
    .I1(inbar[248])
  );
  //OR U491
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U491 (
    .O(n494),
    .I0(n489),
    .I1(n488)
  );
  //AND U491bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U491bar (
    .O(n494bar),
    .I0(n489bar),
    .I1(n488bar)
  );
  //OR U492
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U492 (
    .O(n488),
    .I0(in_46),
    .I1(in_44)
  );
  //AND U492bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U492bar (
    .O(n488bar),
    .I0(in_46bar),
    .I1(in_44bar)
  );
  //OR U493
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U493 (
    .O(n489),
    .I0(in_50),
    .I1(n487)
  );
  //AND U493bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U493bar (
    .O(n489bar),
    .I0(in_50bar),
    .I1(n487bar)
  );
  //OR U494
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U494 (
    .O(n487),
    .I0(in_9),
    .I1(in_80)
  );
  //AND U494bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U494bar (
    .O(n487bar),
    .I0(in_9bar),
    .I1(in_80bar)
  );
endmodule

module sBox_8 ( in, out );

  input wire [7:0] in;
//input_done

  output wire [7:0] out;
//output_done

  wire [255:0] decodeOut;
//wire_done

  decode_8 dec ( .in(in), .out(decodeOut) );
  encode_8 enc ( .in(decodeOut), .out(out) );
endmodule

module CD2_33 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD2_34 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD2_35 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD2_36 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD4_17 ( a, b, y );

  input wire [3:0] a;
  input wire [3:0] b;
  wire [3:0] abar;
  wire [3:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
//input_done

  output wire [15:0] y;
  wire [15:0] ybar;
//output_done

//wire_done

  //AND U1
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1 (
    .O(y[9]),
    .I0(b[1]),
    .I1(a[2])
  );
  //OR U1bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1bar (
    .O(ybar[9]),
    .I0(bbar[1]),
    .I1(abar[2])
  );
  //AND U2
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2 (
    .O(y[8]),
    .I0(b[0]),
    .I1(a[2])
  );
  //OR U2bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2bar (
    .O(ybar[8]),
    .I0(bbar[0]),
    .I1(abar[2])
  );
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[7]),
    .I0(b[3]),
    .I1(a[1])
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[7]),
    .I0(bbar[3]),
    .I1(abar[1])
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[6]),
    .I0(b[2]),
    .I1(a[1])
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[6]),
    .I0(bbar[2]),
    .I1(abar[1])
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[5]),
    .I0(a[1]),
    .I1(b[1])
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[5]),
    .I0(abar[1]),
    .I1(bbar[1])
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[4]),
    .I0(a[1]),
    .I1(b[0])
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[4]),
    .I0(abar[1]),
    .I1(bbar[0])
  );
  //AND U7
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7 (
    .O(y[3]),
    .I0(a[0]),
    .I1(b[3])
  );
  //OR U7bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7bar (
    .O(ybar[3]),
    .I0(abar[0]),
    .I1(bbar[3])
  );
  //AND U8
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8 (
    .O(y[2]),
    .I0(a[0]),
    .I1(b[2])
  );
  //OR U8bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8bar (
    .O(ybar[2]),
    .I0(abar[0]),
    .I1(bbar[2])
  );
  //AND U9
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9 (
    .O(y[1]),
    .I0(a[0]),
    .I1(b[1])
  );
  //OR U9bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9bar (
    .O(ybar[1]),
    .I0(abar[0]),
    .I1(bbar[1])
  );
  //AND U10
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10 (
    .O(y[15]),
    .I0(a[3]),
    .I1(b[3])
  );
  //OR U10bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10bar (
    .O(ybar[15]),
    .I0(abar[3]),
    .I1(bbar[3])
  );
  //AND U11
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11 (
    .O(y[14]),
    .I0(a[3]),
    .I1(b[2])
  );
  //OR U11bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11bar (
    .O(ybar[14]),
    .I0(abar[3]),
    .I1(bbar[2])
  );
  //AND U12
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12 (
    .O(y[13]),
    .I0(a[3]),
    .I1(b[1])
  );
  //OR U12bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12bar (
    .O(ybar[13]),
    .I0(abar[3]),
    .I1(bbar[1])
  );
  //AND U13
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13 (
    .O(y[12]),
    .I0(a[3]),
    .I1(b[0])
  );
  //OR U13bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13bar (
    .O(ybar[12]),
    .I0(abar[3]),
    .I1(bbar[0])
  );
  //AND U14
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14 (
    .O(y[11]),
    .I0(b[3]),
    .I1(a[2])
  );
  //OR U14bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14bar (
    .O(ybar[11]),
    .I0(bbar[3]),
    .I1(abar[2])
  );
  //AND U15
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15 (
    .O(y[10]),
    .I0(b[2]),
    .I1(a[2])
  );
  //OR U15bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15bar (
    .O(ybar[10]),
    .I0(bbar[2]),
    .I1(abar[2])
  );
  //AND U16
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16 (
    .O(y[0]),
    .I0(a[0]),
    .I1(b[0])
  );
  //OR U16bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16bar (
    .O(ybar[0]),
    .I0(abar[0]),
    .I1(bbar[0])
  );
endmodule

module CD4_18 ( a, b, y );

  input wire [3:0] a;
  input wire [3:0] b;
  wire [3:0] abar;
  wire [3:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
//input_done

  output wire [15:0] y;
  wire [15:0] ybar;
//output_done

//wire_done

  //AND U1
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1 (
    .O(y[9]),
    .I0(b[1]),
    .I1(a[2])
  );
  //OR U1bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1bar (
    .O(ybar[9]),
    .I0(bbar[1]),
    .I1(abar[2])
  );
  //AND U2
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2 (
    .O(y[8]),
    .I0(b[0]),
    .I1(a[2])
  );
  //OR U2bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2bar (
    .O(ybar[8]),
    .I0(bbar[0]),
    .I1(abar[2])
  );
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[7]),
    .I0(b[3]),
    .I1(a[1])
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[7]),
    .I0(bbar[3]),
    .I1(abar[1])
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[6]),
    .I0(b[2]),
    .I1(a[1])
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[6]),
    .I0(bbar[2]),
    .I1(abar[1])
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[5]),
    .I0(a[1]),
    .I1(b[1])
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[5]),
    .I0(abar[1]),
    .I1(bbar[1])
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[4]),
    .I0(a[1]),
    .I1(b[0])
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[4]),
    .I0(abar[1]),
    .I1(bbar[0])
  );
  //AND U7
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7 (
    .O(y[3]),
    .I0(a[0]),
    .I1(b[3])
  );
  //OR U7bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7bar (
    .O(ybar[3]),
    .I0(abar[0]),
    .I1(bbar[3])
  );
  //AND U8
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8 (
    .O(y[2]),
    .I0(a[0]),
    .I1(b[2])
  );
  //OR U8bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8bar (
    .O(ybar[2]),
    .I0(abar[0]),
    .I1(bbar[2])
  );
  //AND U9
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9 (
    .O(y[1]),
    .I0(a[0]),
    .I1(b[1])
  );
  //OR U9bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9bar (
    .O(ybar[1]),
    .I0(abar[0]),
    .I1(bbar[1])
  );
  //AND U10
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10 (
    .O(y[15]),
    .I0(a[3]),
    .I1(b[3])
  );
  //OR U10bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10bar (
    .O(ybar[15]),
    .I0(abar[3]),
    .I1(bbar[3])
  );
  //AND U11
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11 (
    .O(y[14]),
    .I0(a[3]),
    .I1(b[2])
  );
  //OR U11bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11bar (
    .O(ybar[14]),
    .I0(abar[3]),
    .I1(bbar[2])
  );
  //AND U12
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12 (
    .O(y[13]),
    .I0(a[3]),
    .I1(b[1])
  );
  //OR U12bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12bar (
    .O(ybar[13]),
    .I0(abar[3]),
    .I1(bbar[1])
  );
  //AND U13
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13 (
    .O(y[12]),
    .I0(a[3]),
    .I1(b[0])
  );
  //OR U13bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13bar (
    .O(ybar[12]),
    .I0(abar[3]),
    .I1(bbar[0])
  );
  //AND U14
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14 (
    .O(y[11]),
    .I0(b[3]),
    .I1(a[2])
  );
  //OR U14bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14bar (
    .O(ybar[11]),
    .I0(bbar[3]),
    .I1(abar[2])
  );
  //AND U15
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15 (
    .O(y[10]),
    .I0(b[2]),
    .I1(a[2])
  );
  //OR U15bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15bar (
    .O(ybar[10]),
    .I0(bbar[2]),
    .I1(abar[2])
  );
  //AND U16
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16 (
    .O(y[0]),
    .I0(a[0]),
    .I1(b[0])
  );
  //OR U16bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16bar (
    .O(ybar[0]),
    .I0(abar[0]),
    .I1(bbar[0])
  );
endmodule

module CD16_9 ( a, b, y );

  input wire [15:0] a;
  input wire [15:0] b;
  wire [15:0] abar;
  wire [15:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign abar[8] = ~a[8];
  assign abar[9] = ~a[9];
  assign abar[10] = ~a[10];
  assign abar[11] = ~a[11];
  assign abar[12] = ~a[12];
  assign abar[13] = ~a[13];
  assign abar[14] = ~a[14];
  assign abar[15] = ~a[15];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign bbar[8] = ~b[8];
  assign bbar[9] = ~b[9];
  assign bbar[10] = ~b[10];
  assign bbar[11] = ~b[11];
  assign bbar[12] = ~b[12];
  assign bbar[13] = ~b[13];
  assign bbar[14] = ~b[14];
  assign bbar[15] = ~b[15];
//input_done

  output wire [255:0] y;
  wire [255:0] ybar;
//output_done

//wire_done

  //AND U1
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1 (
    .O(y[9]),
    .I0(b[9]),
    .I1(a[0])
  );
  //OR U1bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1bar (
    .O(ybar[9]),
    .I0(bbar[9]),
    .I1(abar[0])
  );
  //AND U2
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2 (
    .O(y[99]),
    .I0(b[3]),
    .I1(a[6])
  );
  //OR U2bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2bar (
    .O(ybar[99]),
    .I0(bbar[3]),
    .I1(abar[6])
  );
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[98]),
    .I0(b[2]),
    .I1(a[6])
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[98]),
    .I0(bbar[2]),
    .I1(abar[6])
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[97]),
    .I0(b[1]),
    .I1(a[6])
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[97]),
    .I0(bbar[1]),
    .I1(abar[6])
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[96]),
    .I0(b[0]),
    .I1(a[6])
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[96]),
    .I0(bbar[0]),
    .I1(abar[6])
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[95]),
    .I0(b[15]),
    .I1(a[5])
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[95]),
    .I0(bbar[15]),
    .I1(abar[5])
  );
  //AND U7
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7 (
    .O(y[94]),
    .I0(b[14]),
    .I1(a[5])
  );
  //OR U7bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7bar (
    .O(ybar[94]),
    .I0(bbar[14]),
    .I1(abar[5])
  );
  //AND U8
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8 (
    .O(y[93]),
    .I0(b[13]),
    .I1(a[5])
  );
  //OR U8bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8bar (
    .O(ybar[93]),
    .I0(bbar[13]),
    .I1(abar[5])
  );
  //AND U9
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9 (
    .O(y[92]),
    .I0(b[12]),
    .I1(a[5])
  );
  //OR U9bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9bar (
    .O(ybar[92]),
    .I0(bbar[12]),
    .I1(abar[5])
  );
  //AND U10
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10 (
    .O(y[91]),
    .I0(b[11]),
    .I1(a[5])
  );
  //OR U10bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10bar (
    .O(ybar[91]),
    .I0(bbar[11]),
    .I1(abar[5])
  );
  //AND U11
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11 (
    .O(y[90]),
    .I0(b[10]),
    .I1(a[5])
  );
  //OR U11bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11bar (
    .O(ybar[90]),
    .I0(bbar[10]),
    .I1(abar[5])
  );
  //AND U12
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12 (
    .O(y[8]),
    .I0(b[8]),
    .I1(a[0])
  );
  //OR U12bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12bar (
    .O(ybar[8]),
    .I0(bbar[8]),
    .I1(abar[0])
  );
  //AND U13
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13 (
    .O(y[89]),
    .I0(a[5]),
    .I1(b[9])
  );
  //OR U13bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13bar (
    .O(ybar[89]),
    .I0(abar[5]),
    .I1(bbar[9])
  );
  //AND U14
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14 (
    .O(y[88]),
    .I0(b[8]),
    .I1(a[5])
  );
  //OR U14bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14bar (
    .O(ybar[88]),
    .I0(bbar[8]),
    .I1(abar[5])
  );
  //AND U15
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15 (
    .O(y[87]),
    .I0(b[7]),
    .I1(a[5])
  );
  //OR U15bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15bar (
    .O(ybar[87]),
    .I0(bbar[7]),
    .I1(abar[5])
  );
  //AND U16
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16 (
    .O(y[86]),
    .I0(b[6]),
    .I1(a[5])
  );
  //OR U16bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16bar (
    .O(ybar[86]),
    .I0(bbar[6]),
    .I1(abar[5])
  );
  //AND U17
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U17 (
    .O(y[85]),
    .I0(b[5]),
    .I1(a[5])
  );
  //OR U17bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U17bar (
    .O(ybar[85]),
    .I0(bbar[5]),
    .I1(abar[5])
  );
  //AND U18
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U18 (
    .O(y[84]),
    .I0(b[4]),
    .I1(a[5])
  );
  //OR U18bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U18bar (
    .O(ybar[84]),
    .I0(bbar[4]),
    .I1(abar[5])
  );
  //AND U19
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U19 (
    .O(y[83]),
    .I0(a[5]),
    .I1(b[3])
  );
  //OR U19bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U19bar (
    .O(ybar[83]),
    .I0(abar[5]),
    .I1(bbar[3])
  );
  //AND U20
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U20 (
    .O(y[82]),
    .I0(a[5]),
    .I1(b[2])
  );
  //OR U20bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U20bar (
    .O(ybar[82]),
    .I0(abar[5]),
    .I1(bbar[2])
  );
  //AND U21
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U21 (
    .O(y[81]),
    .I0(a[5]),
    .I1(b[1])
  );
  //OR U21bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U21bar (
    .O(ybar[81]),
    .I0(abar[5]),
    .I1(bbar[1])
  );
  //AND U22
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U22 (
    .O(y[80]),
    .I0(a[5]),
    .I1(b[0])
  );
  //OR U22bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U22bar (
    .O(ybar[80]),
    .I0(abar[5]),
    .I1(bbar[0])
  );
  //AND U23
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U23 (
    .O(y[7]),
    .I0(b[7]),
    .I1(a[0])
  );
  //OR U23bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U23bar (
    .O(ybar[7]),
    .I0(bbar[7]),
    .I1(abar[0])
  );
  //AND U24
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U24 (
    .O(y[79]),
    .I0(a[4]),
    .I1(b[15])
  );
  //OR U24bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U24bar (
    .O(ybar[79]),
    .I0(abar[4]),
    .I1(bbar[15])
  );
  //AND U25
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U25 (
    .O(y[78]),
    .I0(a[4]),
    .I1(b[14])
  );
  //OR U25bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U25bar (
    .O(ybar[78]),
    .I0(abar[4]),
    .I1(bbar[14])
  );
  //AND U26
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U26 (
    .O(y[77]),
    .I0(a[4]),
    .I1(b[13])
  );
  //OR U26bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U26bar (
    .O(ybar[77]),
    .I0(abar[4]),
    .I1(bbar[13])
  );
  //AND U27
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U27 (
    .O(y[76]),
    .I0(a[4]),
    .I1(b[12])
  );
  //OR U27bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U27bar (
    .O(ybar[76]),
    .I0(abar[4]),
    .I1(bbar[12])
  );
  //AND U28
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U28 (
    .O(y[75]),
    .I0(a[4]),
    .I1(b[11])
  );
  //OR U28bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U28bar (
    .O(ybar[75]),
    .I0(abar[4]),
    .I1(bbar[11])
  );
  //AND U29
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U29 (
    .O(y[74]),
    .I0(a[4]),
    .I1(b[10])
  );
  //OR U29bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U29bar (
    .O(ybar[74]),
    .I0(abar[4]),
    .I1(bbar[10])
  );
  //AND U30
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U30 (
    .O(y[73]),
    .I0(a[4]),
    .I1(b[9])
  );
  //OR U30bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U30bar (
    .O(ybar[73]),
    .I0(abar[4]),
    .I1(bbar[9])
  );
  //AND U31
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U31 (
    .O(y[72]),
    .I0(a[4]),
    .I1(b[8])
  );
  //OR U31bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U31bar (
    .O(ybar[72]),
    .I0(abar[4]),
    .I1(bbar[8])
  );
  //AND U32
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U32 (
    .O(y[71]),
    .I0(a[4]),
    .I1(b[7])
  );
  //OR U32bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U32bar (
    .O(ybar[71]),
    .I0(abar[4]),
    .I1(bbar[7])
  );
  //AND U33
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U33 (
    .O(y[70]),
    .I0(a[4]),
    .I1(b[6])
  );
  //OR U33bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U33bar (
    .O(ybar[70]),
    .I0(abar[4]),
    .I1(bbar[6])
  );
  //AND U34
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U34 (
    .O(y[6]),
    .I0(b[6]),
    .I1(a[0])
  );
  //OR U34bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U34bar (
    .O(ybar[6]),
    .I0(bbar[6]),
    .I1(abar[0])
  );
  //AND U35
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U35 (
    .O(y[69]),
    .I0(a[4]),
    .I1(b[5])
  );
  //OR U35bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U35bar (
    .O(ybar[69]),
    .I0(abar[4]),
    .I1(bbar[5])
  );
  //AND U36
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U36 (
    .O(y[68]),
    .I0(a[4]),
    .I1(b[4])
  );
  //OR U36bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U36bar (
    .O(ybar[68]),
    .I0(abar[4]),
    .I1(bbar[4])
  );
  //AND U37
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U37 (
    .O(y[67]),
    .I0(a[4]),
    .I1(b[3])
  );
  //OR U37bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U37bar (
    .O(ybar[67]),
    .I0(abar[4]),
    .I1(bbar[3])
  );
  //AND U38
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U38 (
    .O(y[66]),
    .I0(a[4]),
    .I1(b[2])
  );
  //OR U38bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U38bar (
    .O(ybar[66]),
    .I0(abar[4]),
    .I1(bbar[2])
  );
  //AND U39
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U39 (
    .O(y[65]),
    .I0(a[4]),
    .I1(b[1])
  );
  //OR U39bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U39bar (
    .O(ybar[65]),
    .I0(abar[4]),
    .I1(bbar[1])
  );
  //AND U40
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U40 (
    .O(y[64]),
    .I0(a[4]),
    .I1(b[0])
  );
  //OR U40bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U40bar (
    .O(ybar[64]),
    .I0(abar[4]),
    .I1(bbar[0])
  );
  //AND U41
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U41 (
    .O(y[63]),
    .I0(a[3]),
    .I1(b[15])
  );
  //OR U41bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U41bar (
    .O(ybar[63]),
    .I0(abar[3]),
    .I1(bbar[15])
  );
  //AND U42
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U42 (
    .O(y[62]),
    .I0(a[3]),
    .I1(b[14])
  );
  //OR U42bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U42bar (
    .O(ybar[62]),
    .I0(abar[3]),
    .I1(bbar[14])
  );
  //AND U43
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U43 (
    .O(y[61]),
    .I0(a[3]),
    .I1(b[13])
  );
  //OR U43bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U43bar (
    .O(ybar[61]),
    .I0(abar[3]),
    .I1(bbar[13])
  );
  //AND U44
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U44 (
    .O(y[60]),
    .I0(a[3]),
    .I1(b[12])
  );
  //OR U44bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U44bar (
    .O(ybar[60]),
    .I0(abar[3]),
    .I1(bbar[12])
  );
  //AND U45
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U45 (
    .O(y[5]),
    .I0(b[5]),
    .I1(a[0])
  );
  //OR U45bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U45bar (
    .O(ybar[5]),
    .I0(bbar[5]),
    .I1(abar[0])
  );
  //AND U46
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U46 (
    .O(y[59]),
    .I0(a[3]),
    .I1(b[11])
  );
  //OR U46bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U46bar (
    .O(ybar[59]),
    .I0(abar[3]),
    .I1(bbar[11])
  );
  //AND U47
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U47 (
    .O(y[58]),
    .I0(a[3]),
    .I1(b[10])
  );
  //OR U47bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U47bar (
    .O(ybar[58]),
    .I0(abar[3]),
    .I1(bbar[10])
  );
  //AND U48
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U48 (
    .O(y[57]),
    .I0(a[3]),
    .I1(b[9])
  );
  //OR U48bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U48bar (
    .O(ybar[57]),
    .I0(abar[3]),
    .I1(bbar[9])
  );
  //AND U49
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U49 (
    .O(y[56]),
    .I0(a[3]),
    .I1(b[8])
  );
  //OR U49bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U49bar (
    .O(ybar[56]),
    .I0(abar[3]),
    .I1(bbar[8])
  );
  //AND U50
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U50 (
    .O(y[55]),
    .I0(a[3]),
    .I1(b[7])
  );
  //OR U50bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U50bar (
    .O(ybar[55]),
    .I0(abar[3]),
    .I1(bbar[7])
  );
  //AND U51
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U51 (
    .O(y[54]),
    .I0(a[3]),
    .I1(b[6])
  );
  //OR U51bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U51bar (
    .O(ybar[54]),
    .I0(abar[3]),
    .I1(bbar[6])
  );
  //AND U52
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U52 (
    .O(y[53]),
    .I0(a[3]),
    .I1(b[5])
  );
  //OR U52bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U52bar (
    .O(ybar[53]),
    .I0(abar[3]),
    .I1(bbar[5])
  );
  //AND U53
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U53 (
    .O(y[52]),
    .I0(a[3]),
    .I1(b[4])
  );
  //OR U53bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U53bar (
    .O(ybar[52]),
    .I0(abar[3]),
    .I1(bbar[4])
  );
  //AND U54
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U54 (
    .O(y[51]),
    .I0(a[3]),
    .I1(b[3])
  );
  //OR U54bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U54bar (
    .O(ybar[51]),
    .I0(abar[3]),
    .I1(bbar[3])
  );
  //AND U55
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U55 (
    .O(y[50]),
    .I0(a[3]),
    .I1(b[2])
  );
  //OR U55bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U55bar (
    .O(ybar[50]),
    .I0(abar[3]),
    .I1(bbar[2])
  );
  //AND U56
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U56 (
    .O(y[4]),
    .I0(b[4]),
    .I1(a[0])
  );
  //OR U56bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U56bar (
    .O(ybar[4]),
    .I0(bbar[4]),
    .I1(abar[0])
  );
  //AND U57
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U57 (
    .O(y[49]),
    .I0(a[3]),
    .I1(b[1])
  );
  //OR U57bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U57bar (
    .O(ybar[49]),
    .I0(abar[3]),
    .I1(bbar[1])
  );
  //AND U58
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U58 (
    .O(y[48]),
    .I0(a[3]),
    .I1(b[0])
  );
  //OR U58bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U58bar (
    .O(ybar[48]),
    .I0(abar[3]),
    .I1(bbar[0])
  );
  //AND U59
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U59 (
    .O(y[47]),
    .I0(a[2]),
    .I1(b[15])
  );
  //OR U59bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U59bar (
    .O(ybar[47]),
    .I0(abar[2]),
    .I1(bbar[15])
  );
  //AND U60
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U60 (
    .O(y[46]),
    .I0(a[2]),
    .I1(b[14])
  );
  //OR U60bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U60bar (
    .O(ybar[46]),
    .I0(abar[2]),
    .I1(bbar[14])
  );
  //AND U61
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U61 (
    .O(y[45]),
    .I0(a[2]),
    .I1(b[13])
  );
  //OR U61bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U61bar (
    .O(ybar[45]),
    .I0(abar[2]),
    .I1(bbar[13])
  );
  //AND U62
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U62 (
    .O(y[44]),
    .I0(a[2]),
    .I1(b[12])
  );
  //OR U62bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U62bar (
    .O(ybar[44]),
    .I0(abar[2]),
    .I1(bbar[12])
  );
  //AND U63
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U63 (
    .O(y[43]),
    .I0(a[2]),
    .I1(b[11])
  );
  //OR U63bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U63bar (
    .O(ybar[43]),
    .I0(abar[2]),
    .I1(bbar[11])
  );
  //AND U64
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U64 (
    .O(y[42]),
    .I0(a[2]),
    .I1(b[10])
  );
  //OR U64bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U64bar (
    .O(ybar[42]),
    .I0(abar[2]),
    .I1(bbar[10])
  );
  //AND U65
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U65 (
    .O(y[41]),
    .I0(a[2]),
    .I1(b[9])
  );
  //OR U65bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U65bar (
    .O(ybar[41]),
    .I0(abar[2]),
    .I1(bbar[9])
  );
  //AND U66
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U66 (
    .O(y[40]),
    .I0(a[2]),
    .I1(b[8])
  );
  //OR U66bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U66bar (
    .O(ybar[40]),
    .I0(abar[2]),
    .I1(bbar[8])
  );
  //AND U67
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U67 (
    .O(y[3]),
    .I0(b[3]),
    .I1(a[0])
  );
  //OR U67bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U67bar (
    .O(ybar[3]),
    .I0(bbar[3]),
    .I1(abar[0])
  );
  //AND U68
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U68 (
    .O(y[39]),
    .I0(a[2]),
    .I1(b[7])
  );
  //OR U68bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U68bar (
    .O(ybar[39]),
    .I0(abar[2]),
    .I1(bbar[7])
  );
  //AND U69
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U69 (
    .O(y[38]),
    .I0(a[2]),
    .I1(b[6])
  );
  //OR U69bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U69bar (
    .O(ybar[38]),
    .I0(abar[2]),
    .I1(bbar[6])
  );
  //AND U70
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U70 (
    .O(y[37]),
    .I0(a[2]),
    .I1(b[5])
  );
  //OR U70bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U70bar (
    .O(ybar[37]),
    .I0(abar[2]),
    .I1(bbar[5])
  );
  //AND U71
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U71 (
    .O(y[36]),
    .I0(a[2]),
    .I1(b[4])
  );
  //OR U71bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U71bar (
    .O(ybar[36]),
    .I0(abar[2]),
    .I1(bbar[4])
  );
  //AND U72
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U72 (
    .O(y[35]),
    .I0(a[2]),
    .I1(b[3])
  );
  //OR U72bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U72bar (
    .O(ybar[35]),
    .I0(abar[2]),
    .I1(bbar[3])
  );
  //AND U73
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U73 (
    .O(y[34]),
    .I0(a[2]),
    .I1(b[2])
  );
  //OR U73bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U73bar (
    .O(ybar[34]),
    .I0(abar[2]),
    .I1(bbar[2])
  );
  //AND U74
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U74 (
    .O(y[33]),
    .I0(a[2]),
    .I1(b[1])
  );
  //OR U74bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U74bar (
    .O(ybar[33]),
    .I0(abar[2]),
    .I1(bbar[1])
  );
  //AND U75
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U75 (
    .O(y[32]),
    .I0(a[2]),
    .I1(b[0])
  );
  //OR U75bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U75bar (
    .O(ybar[32]),
    .I0(abar[2]),
    .I1(bbar[0])
  );
  //AND U76
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U76 (
    .O(y[31]),
    .I0(a[1]),
    .I1(b[15])
  );
  //OR U76bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U76bar (
    .O(ybar[31]),
    .I0(abar[1]),
    .I1(bbar[15])
  );
  //AND U77
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U77 (
    .O(y[30]),
    .I0(a[1]),
    .I1(b[14])
  );
  //OR U77bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U77bar (
    .O(ybar[30]),
    .I0(abar[1]),
    .I1(bbar[14])
  );
  //AND U78
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U78 (
    .O(y[2]),
    .I0(b[2]),
    .I1(a[0])
  );
  //OR U78bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U78bar (
    .O(ybar[2]),
    .I0(bbar[2]),
    .I1(abar[0])
  );
  //AND U79
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U79 (
    .O(y[29]),
    .I0(a[1]),
    .I1(b[13])
  );
  //OR U79bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U79bar (
    .O(ybar[29]),
    .I0(abar[1]),
    .I1(bbar[13])
  );
  //AND U80
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U80 (
    .O(y[28]),
    .I0(a[1]),
    .I1(b[12])
  );
  //OR U80bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U80bar (
    .O(ybar[28]),
    .I0(abar[1]),
    .I1(bbar[12])
  );
  //AND U81
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U81 (
    .O(y[27]),
    .I0(a[1]),
    .I1(b[11])
  );
  //OR U81bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U81bar (
    .O(ybar[27]),
    .I0(abar[1]),
    .I1(bbar[11])
  );
  //AND U82
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U82 (
    .O(y[26]),
    .I0(a[1]),
    .I1(b[10])
  );
  //OR U82bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U82bar (
    .O(ybar[26]),
    .I0(abar[1]),
    .I1(bbar[10])
  );
  //AND U83
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U83 (
    .O(y[25]),
    .I0(a[1]),
    .I1(b[9])
  );
  //OR U83bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U83bar (
    .O(ybar[25]),
    .I0(abar[1]),
    .I1(bbar[9])
  );
  //AND U84
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U84 (
    .O(y[255]),
    .I0(a[15]),
    .I1(b[15])
  );
  //OR U84bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U84bar (
    .O(ybar[255]),
    .I0(abar[15]),
    .I1(bbar[15])
  );
  //AND U85
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U85 (
    .O(y[254]),
    .I0(a[15]),
    .I1(b[14])
  );
  //OR U85bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U85bar (
    .O(ybar[254]),
    .I0(abar[15]),
    .I1(bbar[14])
  );
  //AND U86
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U86 (
    .O(y[253]),
    .I0(a[15]),
    .I1(b[13])
  );
  //OR U86bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U86bar (
    .O(ybar[253]),
    .I0(abar[15]),
    .I1(bbar[13])
  );
  //AND U87
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U87 (
    .O(y[252]),
    .I0(a[15]),
    .I1(b[12])
  );
  //OR U87bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U87bar (
    .O(ybar[252]),
    .I0(abar[15]),
    .I1(bbar[12])
  );
  //AND U88
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U88 (
    .O(y[251]),
    .I0(a[15]),
    .I1(b[11])
  );
  //OR U88bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U88bar (
    .O(ybar[251]),
    .I0(abar[15]),
    .I1(bbar[11])
  );
  //AND U89
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U89 (
    .O(y[250]),
    .I0(a[15]),
    .I1(b[10])
  );
  //OR U89bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U89bar (
    .O(ybar[250]),
    .I0(abar[15]),
    .I1(bbar[10])
  );
  //AND U90
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U90 (
    .O(y[24]),
    .I0(a[1]),
    .I1(b[8])
  );
  //OR U90bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U90bar (
    .O(ybar[24]),
    .I0(abar[1]),
    .I1(bbar[8])
  );
  //AND U91
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U91 (
    .O(y[249]),
    .I0(a[15]),
    .I1(b[9])
  );
  //OR U91bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U91bar (
    .O(ybar[249]),
    .I0(abar[15]),
    .I1(bbar[9])
  );
  //AND U92
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U92 (
    .O(y[248]),
    .I0(a[15]),
    .I1(b[8])
  );
  //OR U92bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U92bar (
    .O(ybar[248]),
    .I0(abar[15]),
    .I1(bbar[8])
  );
  //AND U93
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U93 (
    .O(y[247]),
    .I0(a[15]),
    .I1(b[7])
  );
  //OR U93bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U93bar (
    .O(ybar[247]),
    .I0(abar[15]),
    .I1(bbar[7])
  );
  //AND U94
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U94 (
    .O(y[246]),
    .I0(a[15]),
    .I1(b[6])
  );
  //OR U94bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U94bar (
    .O(ybar[246]),
    .I0(abar[15]),
    .I1(bbar[6])
  );
  //AND U95
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U95 (
    .O(y[245]),
    .I0(a[15]),
    .I1(b[5])
  );
  //OR U95bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U95bar (
    .O(ybar[245]),
    .I0(abar[15]),
    .I1(bbar[5])
  );
  //AND U96
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U96 (
    .O(y[244]),
    .I0(a[15]),
    .I1(b[4])
  );
  //OR U96bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U96bar (
    .O(ybar[244]),
    .I0(abar[15]),
    .I1(bbar[4])
  );
  //AND U97
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U97 (
    .O(y[243]),
    .I0(a[15]),
    .I1(b[3])
  );
  //OR U97bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U97bar (
    .O(ybar[243]),
    .I0(abar[15]),
    .I1(bbar[3])
  );
  //AND U98
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U98 (
    .O(y[242]),
    .I0(a[15]),
    .I1(b[2])
  );
  //OR U98bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U98bar (
    .O(ybar[242]),
    .I0(abar[15]),
    .I1(bbar[2])
  );
  //AND U99
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U99 (
    .O(y[241]),
    .I0(a[15]),
    .I1(b[1])
  );
  //OR U99bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U99bar (
    .O(ybar[241]),
    .I0(abar[15]),
    .I1(bbar[1])
  );
  //AND U100
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U100 (
    .O(y[240]),
    .I0(a[15]),
    .I1(b[0])
  );
  //OR U100bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U100bar (
    .O(ybar[240]),
    .I0(abar[15]),
    .I1(bbar[0])
  );
  //AND U101
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U101 (
    .O(y[23]),
    .I0(a[1]),
    .I1(b[7])
  );
  //OR U101bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U101bar (
    .O(ybar[23]),
    .I0(abar[1]),
    .I1(bbar[7])
  );
  //AND U102
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U102 (
    .O(y[239]),
    .I0(a[14]),
    .I1(b[15])
  );
  //OR U102bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U102bar (
    .O(ybar[239]),
    .I0(abar[14]),
    .I1(bbar[15])
  );
  //AND U103
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U103 (
    .O(y[238]),
    .I0(a[14]),
    .I1(b[14])
  );
  //OR U103bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U103bar (
    .O(ybar[238]),
    .I0(abar[14]),
    .I1(bbar[14])
  );
  //AND U104
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U104 (
    .O(y[237]),
    .I0(a[14]),
    .I1(b[13])
  );
  //OR U104bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U104bar (
    .O(ybar[237]),
    .I0(abar[14]),
    .I1(bbar[13])
  );
  //AND U105
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U105 (
    .O(y[236]),
    .I0(a[14]),
    .I1(b[12])
  );
  //OR U105bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U105bar (
    .O(ybar[236]),
    .I0(abar[14]),
    .I1(bbar[12])
  );
  //AND U106
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U106 (
    .O(y[235]),
    .I0(a[14]),
    .I1(b[11])
  );
  //OR U106bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U106bar (
    .O(ybar[235]),
    .I0(abar[14]),
    .I1(bbar[11])
  );
  //AND U107
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U107 (
    .O(y[234]),
    .I0(a[14]),
    .I1(b[10])
  );
  //OR U107bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U107bar (
    .O(ybar[234]),
    .I0(abar[14]),
    .I1(bbar[10])
  );
  //AND U108
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U108 (
    .O(y[233]),
    .I0(a[14]),
    .I1(b[9])
  );
  //OR U108bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U108bar (
    .O(ybar[233]),
    .I0(abar[14]),
    .I1(bbar[9])
  );
  //AND U109
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U109 (
    .O(y[232]),
    .I0(a[14]),
    .I1(b[8])
  );
  //OR U109bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U109bar (
    .O(ybar[232]),
    .I0(abar[14]),
    .I1(bbar[8])
  );
  //AND U110
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U110 (
    .O(y[231]),
    .I0(a[14]),
    .I1(b[7])
  );
  //OR U110bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U110bar (
    .O(ybar[231]),
    .I0(abar[14]),
    .I1(bbar[7])
  );
  //AND U111
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U111 (
    .O(y[230]),
    .I0(a[14]),
    .I1(b[6])
  );
  //OR U111bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U111bar (
    .O(ybar[230]),
    .I0(abar[14]),
    .I1(bbar[6])
  );
  //AND U112
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U112 (
    .O(y[22]),
    .I0(a[1]),
    .I1(b[6])
  );
  //OR U112bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U112bar (
    .O(ybar[22]),
    .I0(abar[1]),
    .I1(bbar[6])
  );
  //AND U113
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U113 (
    .O(y[229]),
    .I0(a[14]),
    .I1(b[5])
  );
  //OR U113bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U113bar (
    .O(ybar[229]),
    .I0(abar[14]),
    .I1(bbar[5])
  );
  //AND U114
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U114 (
    .O(y[228]),
    .I0(a[14]),
    .I1(b[4])
  );
  //OR U114bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U114bar (
    .O(ybar[228]),
    .I0(abar[14]),
    .I1(bbar[4])
  );
  //AND U115
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U115 (
    .O(y[227]),
    .I0(a[14]),
    .I1(b[3])
  );
  //OR U115bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U115bar (
    .O(ybar[227]),
    .I0(abar[14]),
    .I1(bbar[3])
  );
  //AND U116
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U116 (
    .O(y[226]),
    .I0(a[14]),
    .I1(b[2])
  );
  //OR U116bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U116bar (
    .O(ybar[226]),
    .I0(abar[14]),
    .I1(bbar[2])
  );
  //AND U117
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U117 (
    .O(y[225]),
    .I0(a[14]),
    .I1(b[1])
  );
  //OR U117bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U117bar (
    .O(ybar[225]),
    .I0(abar[14]),
    .I1(bbar[1])
  );
  //AND U118
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U118 (
    .O(y[224]),
    .I0(a[14]),
    .I1(b[0])
  );
  //OR U118bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U118bar (
    .O(ybar[224]),
    .I0(abar[14]),
    .I1(bbar[0])
  );
  //AND U119
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U119 (
    .O(y[223]),
    .I0(a[13]),
    .I1(b[15])
  );
  //OR U119bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U119bar (
    .O(ybar[223]),
    .I0(abar[13]),
    .I1(bbar[15])
  );
  //AND U120
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U120 (
    .O(y[222]),
    .I0(a[13]),
    .I1(b[14])
  );
  //OR U120bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U120bar (
    .O(ybar[222]),
    .I0(abar[13]),
    .I1(bbar[14])
  );
  //AND U121
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U121 (
    .O(y[221]),
    .I0(a[13]),
    .I1(b[13])
  );
  //OR U121bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U121bar (
    .O(ybar[221]),
    .I0(abar[13]),
    .I1(bbar[13])
  );
  //AND U122
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U122 (
    .O(y[220]),
    .I0(a[13]),
    .I1(b[12])
  );
  //OR U122bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U122bar (
    .O(ybar[220]),
    .I0(abar[13]),
    .I1(bbar[12])
  );
  //AND U123
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U123 (
    .O(y[21]),
    .I0(a[1]),
    .I1(b[5])
  );
  //OR U123bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U123bar (
    .O(ybar[21]),
    .I0(abar[1]),
    .I1(bbar[5])
  );
  //AND U124
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U124 (
    .O(y[219]),
    .I0(a[13]),
    .I1(b[11])
  );
  //OR U124bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U124bar (
    .O(ybar[219]),
    .I0(abar[13]),
    .I1(bbar[11])
  );
  //AND U125
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U125 (
    .O(y[218]),
    .I0(a[13]),
    .I1(b[10])
  );
  //OR U125bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U125bar (
    .O(ybar[218]),
    .I0(abar[13]),
    .I1(bbar[10])
  );
  //AND U126
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U126 (
    .O(y[217]),
    .I0(a[13]),
    .I1(b[9])
  );
  //OR U126bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U126bar (
    .O(ybar[217]),
    .I0(abar[13]),
    .I1(bbar[9])
  );
  //AND U127
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U127 (
    .O(y[216]),
    .I0(a[13]),
    .I1(b[8])
  );
  //OR U127bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U127bar (
    .O(ybar[216]),
    .I0(abar[13]),
    .I1(bbar[8])
  );
  //AND U128
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U128 (
    .O(y[215]),
    .I0(a[13]),
    .I1(b[7])
  );
  //OR U128bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U128bar (
    .O(ybar[215]),
    .I0(abar[13]),
    .I1(bbar[7])
  );
  //AND U129
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U129 (
    .O(y[214]),
    .I0(a[13]),
    .I1(b[6])
  );
  //OR U129bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U129bar (
    .O(ybar[214]),
    .I0(abar[13]),
    .I1(bbar[6])
  );
  //AND U130
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U130 (
    .O(y[213]),
    .I0(a[13]),
    .I1(b[5])
  );
  //OR U130bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U130bar (
    .O(ybar[213]),
    .I0(abar[13]),
    .I1(bbar[5])
  );
  //AND U131
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U131 (
    .O(y[212]),
    .I0(a[13]),
    .I1(b[4])
  );
  //OR U131bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U131bar (
    .O(ybar[212]),
    .I0(abar[13]),
    .I1(bbar[4])
  );
  //AND U132
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U132 (
    .O(y[211]),
    .I0(a[13]),
    .I1(b[3])
  );
  //OR U132bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U132bar (
    .O(ybar[211]),
    .I0(abar[13]),
    .I1(bbar[3])
  );
  //AND U133
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U133 (
    .O(y[210]),
    .I0(a[13]),
    .I1(b[2])
  );
  //OR U133bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U133bar (
    .O(ybar[210]),
    .I0(abar[13]),
    .I1(bbar[2])
  );
  //AND U134
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U134 (
    .O(y[20]),
    .I0(a[1]),
    .I1(b[4])
  );
  //OR U134bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U134bar (
    .O(ybar[20]),
    .I0(abar[1]),
    .I1(bbar[4])
  );
  //AND U135
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U135 (
    .O(y[209]),
    .I0(a[13]),
    .I1(b[1])
  );
  //OR U135bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U135bar (
    .O(ybar[209]),
    .I0(abar[13]),
    .I1(bbar[1])
  );
  //AND U136
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U136 (
    .O(y[208]),
    .I0(a[13]),
    .I1(b[0])
  );
  //OR U136bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U136bar (
    .O(ybar[208]),
    .I0(abar[13]),
    .I1(bbar[0])
  );
  //AND U137
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U137 (
    .O(y[207]),
    .I0(a[12]),
    .I1(b[15])
  );
  //OR U137bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U137bar (
    .O(ybar[207]),
    .I0(abar[12]),
    .I1(bbar[15])
  );
  //AND U138
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U138 (
    .O(y[206]),
    .I0(a[12]),
    .I1(b[14])
  );
  //OR U138bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U138bar (
    .O(ybar[206]),
    .I0(abar[12]),
    .I1(bbar[14])
  );
  //AND U139
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U139 (
    .O(y[205]),
    .I0(a[12]),
    .I1(b[13])
  );
  //OR U139bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U139bar (
    .O(ybar[205]),
    .I0(abar[12]),
    .I1(bbar[13])
  );
  //AND U140
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U140 (
    .O(y[204]),
    .I0(a[12]),
    .I1(b[12])
  );
  //OR U140bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U140bar (
    .O(ybar[204]),
    .I0(abar[12]),
    .I1(bbar[12])
  );
  //AND U141
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U141 (
    .O(y[203]),
    .I0(a[12]),
    .I1(b[11])
  );
  //OR U141bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U141bar (
    .O(ybar[203]),
    .I0(abar[12]),
    .I1(bbar[11])
  );
  //AND U142
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U142 (
    .O(y[202]),
    .I0(a[12]),
    .I1(b[10])
  );
  //OR U142bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U142bar (
    .O(ybar[202]),
    .I0(abar[12]),
    .I1(bbar[10])
  );
  //AND U143
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U143 (
    .O(y[201]),
    .I0(a[12]),
    .I1(b[9])
  );
  //OR U143bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U143bar (
    .O(ybar[201]),
    .I0(abar[12]),
    .I1(bbar[9])
  );
  //AND U144
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U144 (
    .O(y[200]),
    .I0(a[12]),
    .I1(b[8])
  );
  //OR U144bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U144bar (
    .O(ybar[200]),
    .I0(abar[12]),
    .I1(bbar[8])
  );
  //AND U145
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U145 (
    .O(y[1]),
    .I0(b[1]),
    .I1(a[0])
  );
  //OR U145bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U145bar (
    .O(ybar[1]),
    .I0(bbar[1]),
    .I1(abar[0])
  );
  //AND U146
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U146 (
    .O(y[19]),
    .I0(a[1]),
    .I1(b[3])
  );
  //OR U146bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U146bar (
    .O(ybar[19]),
    .I0(abar[1]),
    .I1(bbar[3])
  );
  //AND U147
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U147 (
    .O(y[199]),
    .I0(a[12]),
    .I1(b[7])
  );
  //OR U147bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U147bar (
    .O(ybar[199]),
    .I0(abar[12]),
    .I1(bbar[7])
  );
  //AND U148
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U148 (
    .O(y[198]),
    .I0(a[12]),
    .I1(b[6])
  );
  //OR U148bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U148bar (
    .O(ybar[198]),
    .I0(abar[12]),
    .I1(bbar[6])
  );
  //AND U149
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U149 (
    .O(y[197]),
    .I0(a[12]),
    .I1(b[5])
  );
  //OR U149bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U149bar (
    .O(ybar[197]),
    .I0(abar[12]),
    .I1(bbar[5])
  );
  //AND U150
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U150 (
    .O(y[196]),
    .I0(a[12]),
    .I1(b[4])
  );
  //OR U150bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U150bar (
    .O(ybar[196]),
    .I0(abar[12]),
    .I1(bbar[4])
  );
  //AND U151
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U151 (
    .O(y[195]),
    .I0(a[12]),
    .I1(b[3])
  );
  //OR U151bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U151bar (
    .O(ybar[195]),
    .I0(abar[12]),
    .I1(bbar[3])
  );
  //AND U152
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U152 (
    .O(y[194]),
    .I0(a[12]),
    .I1(b[2])
  );
  //OR U152bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U152bar (
    .O(ybar[194]),
    .I0(abar[12]),
    .I1(bbar[2])
  );
  //AND U153
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U153 (
    .O(y[193]),
    .I0(a[12]),
    .I1(b[1])
  );
  //OR U153bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U153bar (
    .O(ybar[193]),
    .I0(abar[12]),
    .I1(bbar[1])
  );
  //AND U154
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U154 (
    .O(y[192]),
    .I0(a[12]),
    .I1(b[0])
  );
  //OR U154bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U154bar (
    .O(ybar[192]),
    .I0(abar[12]),
    .I1(bbar[0])
  );
  //AND U155
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U155 (
    .O(y[191]),
    .I0(a[11]),
    .I1(b[15])
  );
  //OR U155bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U155bar (
    .O(ybar[191]),
    .I0(abar[11]),
    .I1(bbar[15])
  );
  //AND U156
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U156 (
    .O(y[190]),
    .I0(a[11]),
    .I1(b[14])
  );
  //OR U156bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U156bar (
    .O(ybar[190]),
    .I0(abar[11]),
    .I1(bbar[14])
  );
  //AND U157
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U157 (
    .O(y[18]),
    .I0(a[1]),
    .I1(b[2])
  );
  //OR U157bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U157bar (
    .O(ybar[18]),
    .I0(abar[1]),
    .I1(bbar[2])
  );
  //AND U158
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U158 (
    .O(y[189]),
    .I0(a[11]),
    .I1(b[13])
  );
  //OR U158bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U158bar (
    .O(ybar[189]),
    .I0(abar[11]),
    .I1(bbar[13])
  );
  //AND U159
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U159 (
    .O(y[188]),
    .I0(a[11]),
    .I1(b[12])
  );
  //OR U159bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U159bar (
    .O(ybar[188]),
    .I0(abar[11]),
    .I1(bbar[12])
  );
  //AND U160
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U160 (
    .O(y[187]),
    .I0(a[11]),
    .I1(b[11])
  );
  //OR U160bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U160bar (
    .O(ybar[187]),
    .I0(abar[11]),
    .I1(bbar[11])
  );
  //AND U161
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U161 (
    .O(y[186]),
    .I0(a[11]),
    .I1(b[10])
  );
  //OR U161bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U161bar (
    .O(ybar[186]),
    .I0(abar[11]),
    .I1(bbar[10])
  );
  //AND U162
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U162 (
    .O(y[185]),
    .I0(a[11]),
    .I1(b[9])
  );
  //OR U162bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U162bar (
    .O(ybar[185]),
    .I0(abar[11]),
    .I1(bbar[9])
  );
  //AND U163
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U163 (
    .O(y[184]),
    .I0(a[11]),
    .I1(b[8])
  );
  //OR U163bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U163bar (
    .O(ybar[184]),
    .I0(abar[11]),
    .I1(bbar[8])
  );
  //AND U164
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U164 (
    .O(y[183]),
    .I0(a[11]),
    .I1(b[7])
  );
  //OR U164bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U164bar (
    .O(ybar[183]),
    .I0(abar[11]),
    .I1(bbar[7])
  );
  //AND U165
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U165 (
    .O(y[182]),
    .I0(a[11]),
    .I1(b[6])
  );
  //OR U165bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U165bar (
    .O(ybar[182]),
    .I0(abar[11]),
    .I1(bbar[6])
  );
  //AND U166
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U166 (
    .O(y[181]),
    .I0(a[11]),
    .I1(b[5])
  );
  //OR U166bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U166bar (
    .O(ybar[181]),
    .I0(abar[11]),
    .I1(bbar[5])
  );
  //AND U167
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U167 (
    .O(y[180]),
    .I0(a[11]),
    .I1(b[4])
  );
  //OR U167bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U167bar (
    .O(ybar[180]),
    .I0(abar[11]),
    .I1(bbar[4])
  );
  //AND U168
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U168 (
    .O(y[17]),
    .I0(a[1]),
    .I1(b[1])
  );
  //OR U168bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U168bar (
    .O(ybar[17]),
    .I0(abar[1]),
    .I1(bbar[1])
  );
  //AND U169
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U169 (
    .O(y[179]),
    .I0(a[11]),
    .I1(b[3])
  );
  //OR U169bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U169bar (
    .O(ybar[179]),
    .I0(abar[11]),
    .I1(bbar[3])
  );
  //AND U170
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U170 (
    .O(y[178]),
    .I0(a[11]),
    .I1(b[2])
  );
  //OR U170bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U170bar (
    .O(ybar[178]),
    .I0(abar[11]),
    .I1(bbar[2])
  );
  //AND U171
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U171 (
    .O(y[177]),
    .I0(a[11]),
    .I1(b[1])
  );
  //OR U171bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U171bar (
    .O(ybar[177]),
    .I0(abar[11]),
    .I1(bbar[1])
  );
  //AND U172
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U172 (
    .O(y[176]),
    .I0(a[11]),
    .I1(b[0])
  );
  //OR U172bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U172bar (
    .O(ybar[176]),
    .I0(abar[11]),
    .I1(bbar[0])
  );
  //AND U173
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U173 (
    .O(y[175]),
    .I0(a[10]),
    .I1(b[15])
  );
  //OR U173bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U173bar (
    .O(ybar[175]),
    .I0(abar[10]),
    .I1(bbar[15])
  );
  //AND U174
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U174 (
    .O(y[174]),
    .I0(a[10]),
    .I1(b[14])
  );
  //OR U174bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U174bar (
    .O(ybar[174]),
    .I0(abar[10]),
    .I1(bbar[14])
  );
  //AND U175
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U175 (
    .O(y[173]),
    .I0(a[10]),
    .I1(b[13])
  );
  //OR U175bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U175bar (
    .O(ybar[173]),
    .I0(abar[10]),
    .I1(bbar[13])
  );
  //AND U176
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U176 (
    .O(y[172]),
    .I0(a[10]),
    .I1(b[12])
  );
  //OR U176bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U176bar (
    .O(ybar[172]),
    .I0(abar[10]),
    .I1(bbar[12])
  );
  //AND U177
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U177 (
    .O(y[171]),
    .I0(a[10]),
    .I1(b[11])
  );
  //OR U177bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U177bar (
    .O(ybar[171]),
    .I0(abar[10]),
    .I1(bbar[11])
  );
  //AND U178
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U178 (
    .O(y[170]),
    .I0(a[10]),
    .I1(b[10])
  );
  //OR U178bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U178bar (
    .O(ybar[170]),
    .I0(abar[10]),
    .I1(bbar[10])
  );
  //AND U179
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U179 (
    .O(y[16]),
    .I0(a[1]),
    .I1(b[0])
  );
  //OR U179bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U179bar (
    .O(ybar[16]),
    .I0(abar[1]),
    .I1(bbar[0])
  );
  //AND U180
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U180 (
    .O(y[169]),
    .I0(a[10]),
    .I1(b[9])
  );
  //OR U180bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U180bar (
    .O(ybar[169]),
    .I0(abar[10]),
    .I1(bbar[9])
  );
  //AND U181
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U181 (
    .O(y[168]),
    .I0(a[10]),
    .I1(b[8])
  );
  //OR U181bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U181bar (
    .O(ybar[168]),
    .I0(abar[10]),
    .I1(bbar[8])
  );
  //AND U182
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U182 (
    .O(y[167]),
    .I0(a[10]),
    .I1(b[7])
  );
  //OR U182bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U182bar (
    .O(ybar[167]),
    .I0(abar[10]),
    .I1(bbar[7])
  );
  //AND U183
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U183 (
    .O(y[166]),
    .I0(a[10]),
    .I1(b[6])
  );
  //OR U183bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U183bar (
    .O(ybar[166]),
    .I0(abar[10]),
    .I1(bbar[6])
  );
  //AND U184
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U184 (
    .O(y[165]),
    .I0(a[10]),
    .I1(b[5])
  );
  //OR U184bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U184bar (
    .O(ybar[165]),
    .I0(abar[10]),
    .I1(bbar[5])
  );
  //AND U185
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U185 (
    .O(y[164]),
    .I0(a[10]),
    .I1(b[4])
  );
  //OR U185bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U185bar (
    .O(ybar[164]),
    .I0(abar[10]),
    .I1(bbar[4])
  );
  //AND U186
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U186 (
    .O(y[163]),
    .I0(a[10]),
    .I1(b[3])
  );
  //OR U186bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U186bar (
    .O(ybar[163]),
    .I0(abar[10]),
    .I1(bbar[3])
  );
  //AND U187
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U187 (
    .O(y[162]),
    .I0(a[10]),
    .I1(b[2])
  );
  //OR U187bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U187bar (
    .O(ybar[162]),
    .I0(abar[10]),
    .I1(bbar[2])
  );
  //AND U188
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U188 (
    .O(y[161]),
    .I0(a[10]),
    .I1(b[1])
  );
  //OR U188bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U188bar (
    .O(ybar[161]),
    .I0(abar[10]),
    .I1(bbar[1])
  );
  //AND U189
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U189 (
    .O(y[160]),
    .I0(a[10]),
    .I1(b[0])
  );
  //OR U189bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U189bar (
    .O(ybar[160]),
    .I0(abar[10]),
    .I1(bbar[0])
  );
  //AND U190
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U190 (
    .O(y[15]),
    .I0(b[15]),
    .I1(a[0])
  );
  //OR U190bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U190bar (
    .O(ybar[15]),
    .I0(bbar[15]),
    .I1(abar[0])
  );
  //AND U191
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U191 (
    .O(y[159]),
    .I0(a[9]),
    .I1(b[15])
  );
  //OR U191bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U191bar (
    .O(ybar[159]),
    .I0(abar[9]),
    .I1(bbar[15])
  );
  //AND U192
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U192 (
    .O(y[158]),
    .I0(a[9]),
    .I1(b[14])
  );
  //OR U192bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U192bar (
    .O(ybar[158]),
    .I0(abar[9]),
    .I1(bbar[14])
  );
  //AND U193
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U193 (
    .O(y[157]),
    .I0(a[9]),
    .I1(b[13])
  );
  //OR U193bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U193bar (
    .O(ybar[157]),
    .I0(abar[9]),
    .I1(bbar[13])
  );
  //AND U194
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U194 (
    .O(y[156]),
    .I0(a[9]),
    .I1(b[12])
  );
  //OR U194bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U194bar (
    .O(ybar[156]),
    .I0(abar[9]),
    .I1(bbar[12])
  );
  //AND U195
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U195 (
    .O(y[155]),
    .I0(a[9]),
    .I1(b[11])
  );
  //OR U195bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U195bar (
    .O(ybar[155]),
    .I0(abar[9]),
    .I1(bbar[11])
  );
  //AND U196
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U196 (
    .O(y[154]),
    .I0(a[9]),
    .I1(b[10])
  );
  //OR U196bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U196bar (
    .O(ybar[154]),
    .I0(abar[9]),
    .I1(bbar[10])
  );
  //AND U197
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U197 (
    .O(y[153]),
    .I0(a[9]),
    .I1(b[9])
  );
  //OR U197bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U197bar (
    .O(ybar[153]),
    .I0(abar[9]),
    .I1(bbar[9])
  );
  //AND U198
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U198 (
    .O(y[152]),
    .I0(a[9]),
    .I1(b[8])
  );
  //OR U198bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U198bar (
    .O(ybar[152]),
    .I0(abar[9]),
    .I1(bbar[8])
  );
  //AND U199
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U199 (
    .O(y[151]),
    .I0(a[9]),
    .I1(b[7])
  );
  //OR U199bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U199bar (
    .O(ybar[151]),
    .I0(abar[9]),
    .I1(bbar[7])
  );
  //AND U200
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U200 (
    .O(y[150]),
    .I0(a[9]),
    .I1(b[6])
  );
  //OR U200bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U200bar (
    .O(ybar[150]),
    .I0(abar[9]),
    .I1(bbar[6])
  );
  //AND U201
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U201 (
    .O(y[14]),
    .I0(b[14]),
    .I1(a[0])
  );
  //OR U201bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U201bar (
    .O(ybar[14]),
    .I0(bbar[14]),
    .I1(abar[0])
  );
  //AND U202
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U202 (
    .O(y[149]),
    .I0(a[9]),
    .I1(b[5])
  );
  //OR U202bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U202bar (
    .O(ybar[149]),
    .I0(abar[9]),
    .I1(bbar[5])
  );
  //AND U203
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U203 (
    .O(y[148]),
    .I0(a[9]),
    .I1(b[4])
  );
  //OR U203bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U203bar (
    .O(ybar[148]),
    .I0(abar[9]),
    .I1(bbar[4])
  );
  //AND U204
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U204 (
    .O(y[147]),
    .I0(a[9]),
    .I1(b[3])
  );
  //OR U204bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U204bar (
    .O(ybar[147]),
    .I0(abar[9]),
    .I1(bbar[3])
  );
  //AND U205
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U205 (
    .O(y[146]),
    .I0(a[9]),
    .I1(b[2])
  );
  //OR U205bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U205bar (
    .O(ybar[146]),
    .I0(abar[9]),
    .I1(bbar[2])
  );
  //AND U206
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U206 (
    .O(y[145]),
    .I0(a[9]),
    .I1(b[1])
  );
  //OR U206bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U206bar (
    .O(ybar[145]),
    .I0(abar[9]),
    .I1(bbar[1])
  );
  //AND U207
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U207 (
    .O(y[144]),
    .I0(a[9]),
    .I1(b[0])
  );
  //OR U207bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U207bar (
    .O(ybar[144]),
    .I0(abar[9]),
    .I1(bbar[0])
  );
  //AND U208
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U208 (
    .O(y[143]),
    .I0(a[8]),
    .I1(b[15])
  );
  //OR U208bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U208bar (
    .O(ybar[143]),
    .I0(abar[8]),
    .I1(bbar[15])
  );
  //AND U209
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U209 (
    .O(y[142]),
    .I0(a[8]),
    .I1(b[14])
  );
  //OR U209bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U209bar (
    .O(ybar[142]),
    .I0(abar[8]),
    .I1(bbar[14])
  );
  //AND U210
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U210 (
    .O(y[141]),
    .I0(a[8]),
    .I1(b[13])
  );
  //OR U210bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U210bar (
    .O(ybar[141]),
    .I0(abar[8]),
    .I1(bbar[13])
  );
  //AND U211
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U211 (
    .O(y[140]),
    .I0(a[8]),
    .I1(b[12])
  );
  //OR U211bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U211bar (
    .O(ybar[140]),
    .I0(abar[8]),
    .I1(bbar[12])
  );
  //AND U212
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U212 (
    .O(y[13]),
    .I0(b[13]),
    .I1(a[0])
  );
  //OR U212bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U212bar (
    .O(ybar[13]),
    .I0(bbar[13]),
    .I1(abar[0])
  );
  //AND U213
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U213 (
    .O(y[139]),
    .I0(a[8]),
    .I1(b[11])
  );
  //OR U213bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U213bar (
    .O(ybar[139]),
    .I0(abar[8]),
    .I1(bbar[11])
  );
  //AND U214
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U214 (
    .O(y[138]),
    .I0(a[8]),
    .I1(b[10])
  );
  //OR U214bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U214bar (
    .O(ybar[138]),
    .I0(abar[8]),
    .I1(bbar[10])
  );
  //AND U215
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U215 (
    .O(y[137]),
    .I0(a[8]),
    .I1(b[9])
  );
  //OR U215bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U215bar (
    .O(ybar[137]),
    .I0(abar[8]),
    .I1(bbar[9])
  );
  //AND U216
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U216 (
    .O(y[136]),
    .I0(a[8]),
    .I1(b[8])
  );
  //OR U216bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U216bar (
    .O(ybar[136]),
    .I0(abar[8]),
    .I1(bbar[8])
  );
  //AND U217
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U217 (
    .O(y[135]),
    .I0(a[8]),
    .I1(b[7])
  );
  //OR U217bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U217bar (
    .O(ybar[135]),
    .I0(abar[8]),
    .I1(bbar[7])
  );
  //AND U218
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U218 (
    .O(y[134]),
    .I0(a[8]),
    .I1(b[6])
  );
  //OR U218bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U218bar (
    .O(ybar[134]),
    .I0(abar[8]),
    .I1(bbar[6])
  );
  //AND U219
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U219 (
    .O(y[133]),
    .I0(a[8]),
    .I1(b[5])
  );
  //OR U219bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U219bar (
    .O(ybar[133]),
    .I0(abar[8]),
    .I1(bbar[5])
  );
  //AND U220
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U220 (
    .O(y[132]),
    .I0(a[8]),
    .I1(b[4])
  );
  //OR U220bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U220bar (
    .O(ybar[132]),
    .I0(abar[8]),
    .I1(bbar[4])
  );
  //AND U221
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U221 (
    .O(y[131]),
    .I0(a[8]),
    .I1(b[3])
  );
  //OR U221bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U221bar (
    .O(ybar[131]),
    .I0(abar[8]),
    .I1(bbar[3])
  );
  //AND U222
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U222 (
    .O(y[130]),
    .I0(a[8]),
    .I1(b[2])
  );
  //OR U222bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U222bar (
    .O(ybar[130]),
    .I0(abar[8]),
    .I1(bbar[2])
  );
  //AND U223
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U223 (
    .O(y[12]),
    .I0(b[12]),
    .I1(a[0])
  );
  //OR U223bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U223bar (
    .O(ybar[12]),
    .I0(bbar[12]),
    .I1(abar[0])
  );
  //AND U224
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U224 (
    .O(y[129]),
    .I0(a[8]),
    .I1(b[1])
  );
  //OR U224bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U224bar (
    .O(ybar[129]),
    .I0(abar[8]),
    .I1(bbar[1])
  );
  //AND U225
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U225 (
    .O(y[128]),
    .I0(a[8]),
    .I1(b[0])
  );
  //OR U225bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U225bar (
    .O(ybar[128]),
    .I0(abar[8]),
    .I1(bbar[0])
  );
  //AND U226
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U226 (
    .O(y[127]),
    .I0(a[7]),
    .I1(b[15])
  );
  //OR U226bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U226bar (
    .O(ybar[127]),
    .I0(abar[7]),
    .I1(bbar[15])
  );
  //AND U227
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U227 (
    .O(y[126]),
    .I0(a[7]),
    .I1(b[14])
  );
  //OR U227bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U227bar (
    .O(ybar[126]),
    .I0(abar[7]),
    .I1(bbar[14])
  );
  //AND U228
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U228 (
    .O(y[125]),
    .I0(a[7]),
    .I1(b[13])
  );
  //OR U228bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U228bar (
    .O(ybar[125]),
    .I0(abar[7]),
    .I1(bbar[13])
  );
  //AND U229
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U229 (
    .O(y[124]),
    .I0(a[7]),
    .I1(b[12])
  );
  //OR U229bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U229bar (
    .O(ybar[124]),
    .I0(abar[7]),
    .I1(bbar[12])
  );
  //AND U230
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U230 (
    .O(y[123]),
    .I0(a[7]),
    .I1(b[11])
  );
  //OR U230bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U230bar (
    .O(ybar[123]),
    .I0(abar[7]),
    .I1(bbar[11])
  );
  //AND U231
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U231 (
    .O(y[122]),
    .I0(a[7]),
    .I1(b[10])
  );
  //OR U231bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U231bar (
    .O(ybar[122]),
    .I0(abar[7]),
    .I1(bbar[10])
  );
  //AND U232
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U232 (
    .O(y[121]),
    .I0(a[7]),
    .I1(b[9])
  );
  //OR U232bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U232bar (
    .O(ybar[121]),
    .I0(abar[7]),
    .I1(bbar[9])
  );
  //AND U233
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U233 (
    .O(y[120]),
    .I0(a[7]),
    .I1(b[8])
  );
  //OR U233bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U233bar (
    .O(ybar[120]),
    .I0(abar[7]),
    .I1(bbar[8])
  );
  //AND U234
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U234 (
    .O(y[11]),
    .I0(b[11]),
    .I1(a[0])
  );
  //OR U234bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U234bar (
    .O(ybar[11]),
    .I0(bbar[11]),
    .I1(abar[0])
  );
  //AND U235
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U235 (
    .O(y[119]),
    .I0(a[7]),
    .I1(b[7])
  );
  //OR U235bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U235bar (
    .O(ybar[119]),
    .I0(abar[7]),
    .I1(bbar[7])
  );
  //AND U236
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U236 (
    .O(y[118]),
    .I0(a[7]),
    .I1(b[6])
  );
  //OR U236bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U236bar (
    .O(ybar[118]),
    .I0(abar[7]),
    .I1(bbar[6])
  );
  //AND U237
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U237 (
    .O(y[117]),
    .I0(a[7]),
    .I1(b[5])
  );
  //OR U237bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U237bar (
    .O(ybar[117]),
    .I0(abar[7]),
    .I1(bbar[5])
  );
  //AND U238
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U238 (
    .O(y[116]),
    .I0(a[7]),
    .I1(b[4])
  );
  //OR U238bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U238bar (
    .O(ybar[116]),
    .I0(abar[7]),
    .I1(bbar[4])
  );
  //AND U239
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U239 (
    .O(y[115]),
    .I0(a[7]),
    .I1(b[3])
  );
  //OR U239bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U239bar (
    .O(ybar[115]),
    .I0(abar[7]),
    .I1(bbar[3])
  );
  //AND U240
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U240 (
    .O(y[114]),
    .I0(a[7]),
    .I1(b[2])
  );
  //OR U240bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U240bar (
    .O(ybar[114]),
    .I0(abar[7]),
    .I1(bbar[2])
  );
  //AND U241
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U241 (
    .O(y[113]),
    .I0(a[7]),
    .I1(b[1])
  );
  //OR U241bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U241bar (
    .O(ybar[113]),
    .I0(abar[7]),
    .I1(bbar[1])
  );
  //AND U242
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U242 (
    .O(y[112]),
    .I0(a[7]),
    .I1(b[0])
  );
  //OR U242bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U242bar (
    .O(ybar[112]),
    .I0(abar[7]),
    .I1(bbar[0])
  );
  //AND U243
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U243 (
    .O(y[111]),
    .I0(b[15]),
    .I1(a[6])
  );
  //OR U243bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U243bar (
    .O(ybar[111]),
    .I0(bbar[15]),
    .I1(abar[6])
  );
  //AND U244
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U244 (
    .O(y[110]),
    .I0(b[14]),
    .I1(a[6])
  );
  //OR U244bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U244bar (
    .O(ybar[110]),
    .I0(bbar[14]),
    .I1(abar[6])
  );
  //AND U245
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U245 (
    .O(y[10]),
    .I0(b[10]),
    .I1(a[0])
  );
  //OR U245bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U245bar (
    .O(ybar[10]),
    .I0(bbar[10]),
    .I1(abar[0])
  );
  //AND U246
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U246 (
    .O(y[109]),
    .I0(b[13]),
    .I1(a[6])
  );
  //OR U246bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U246bar (
    .O(ybar[109]),
    .I0(bbar[13]),
    .I1(abar[6])
  );
  //AND U247
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U247 (
    .O(y[108]),
    .I0(b[12]),
    .I1(a[6])
  );
  //OR U247bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U247bar (
    .O(ybar[108]),
    .I0(bbar[12]),
    .I1(abar[6])
  );
  //AND U248
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U248 (
    .O(y[107]),
    .I0(b[11]),
    .I1(a[6])
  );
  //OR U248bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U248bar (
    .O(ybar[107]),
    .I0(bbar[11]),
    .I1(abar[6])
  );
  //AND U249
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U249 (
    .O(y[106]),
    .I0(b[10]),
    .I1(a[6])
  );
  //OR U249bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U249bar (
    .O(ybar[106]),
    .I0(bbar[10]),
    .I1(abar[6])
  );
  //AND U250
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U250 (
    .O(y[105]),
    .I0(a[6]),
    .I1(b[9])
  );
  //OR U250bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U250bar (
    .O(ybar[105]),
    .I0(abar[6]),
    .I1(bbar[9])
  );
  //AND U251
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U251 (
    .O(y[104]),
    .I0(b[8]),
    .I1(a[6])
  );
  //OR U251bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U251bar (
    .O(ybar[104]),
    .I0(bbar[8]),
    .I1(abar[6])
  );
  //AND U252
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U252 (
    .O(y[103]),
    .I0(b[7]),
    .I1(a[6])
  );
  //OR U252bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U252bar (
    .O(ybar[103]),
    .I0(bbar[7]),
    .I1(abar[6])
  );
  //AND U253
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U253 (
    .O(y[102]),
    .I0(b[6]),
    .I1(a[6])
  );
  //OR U253bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U253bar (
    .O(ybar[102]),
    .I0(bbar[6]),
    .I1(abar[6])
  );
  //AND U254
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U254 (
    .O(y[101]),
    .I0(b[5]),
    .I1(a[6])
  );
  //OR U254bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U254bar (
    .O(ybar[101]),
    .I0(bbar[5]),
    .I1(abar[6])
  );
  //AND U255
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U255 (
    .O(y[100]),
    .I0(b[4]),
    .I1(a[6])
  );
  //OR U255bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U255bar (
    .O(ybar[100]),
    .I0(bbar[4]),
    .I1(abar[6])
  );
  //AND U256
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U256 (
    .O(y[0]),
    .I0(b[0]),
    .I1(a[0])
  );
  //OR U256bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U256bar (
    .O(ybar[0]),
    .I0(bbar[0]),
    .I1(abar[0])
  );
endmodule

module decode_9 ( in, out );

  input wire [7:0] in;
//input_done

  output wire [255:0] out;
//output_done

  wire [15:0] level1;
  wire [31:0] level2;
//wire_done

  CD2_36 cd_l1_1 ( .a(in[1]), .b(in[0]), .y(level1[3:0]) );
  CD2_35 cd_l1_2 ( .a(in[3]), .b(in[2]), .y(level1[7:4]) );
  CD2_34 cd_l1_3 ( .a(in[5]), .b(in[4]), .y(level1[11:8]) );
  CD2_33 cd_l1_4 ( .a(in[7]), .b(in[6]), .y(level1[15:12]) );
  CD4_18 cd_l2_1 ( .a(level1[7:4]), .b(level1[3:0]), .y(level2[15:0]) );
  CD4_17 cd_l2_2 ( .a(level1[15:12]), .b(level1[11:8]), .y(level2[31:16]) );
  CD16_9 cd_l3 ( .a(level2[31:16]), .b(level2[15:0]), .y(out) );
endmodule

module encode_9 ( in, out );

  input wire [255:0] in;
  wire [255:0] inbar;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
  assign inbar[8] = ~in[8];
  assign inbar[9] = ~in[9];
  assign inbar[10] = ~in[10];
  assign inbar[11] = ~in[11];
  assign inbar[12] = ~in[12];
  assign inbar[13] = ~in[13];
  assign inbar[14] = ~in[14];
  assign inbar[15] = ~in[15];
  assign inbar[16] = ~in[16];
  assign inbar[17] = ~in[17];
  assign inbar[18] = ~in[18];
  assign inbar[19] = ~in[19];
  assign inbar[20] = ~in[20];
  assign inbar[21] = ~in[21];
  assign inbar[22] = ~in[22];
  assign inbar[23] = ~in[23];
  assign inbar[24] = ~in[24];
  assign inbar[25] = ~in[25];
  assign inbar[26] = ~in[26];
  assign inbar[27] = ~in[27];
  assign inbar[28] = ~in[28];
  assign inbar[29] = ~in[29];
  assign inbar[30] = ~in[30];
  assign inbar[31] = ~in[31];
  assign inbar[32] = ~in[32];
  assign inbar[33] = ~in[33];
  assign inbar[34] = ~in[34];
  assign inbar[35] = ~in[35];
  assign inbar[36] = ~in[36];
  assign inbar[37] = ~in[37];
  assign inbar[38] = ~in[38];
  assign inbar[39] = ~in[39];
  assign inbar[40] = ~in[40];
  assign inbar[41] = ~in[41];
  assign inbar[42] = ~in[42];
  assign inbar[43] = ~in[43];
  assign inbar[44] = ~in[44];
  assign inbar[45] = ~in[45];
  assign inbar[46] = ~in[46];
  assign inbar[47] = ~in[47];
  assign inbar[48] = ~in[48];
  assign inbar[49] = ~in[49];
  assign inbar[50] = ~in[50];
  assign inbar[51] = ~in[51];
  assign inbar[52] = ~in[52];
  assign inbar[53] = ~in[53];
  assign inbar[54] = ~in[54];
  assign inbar[55] = ~in[55];
  assign inbar[56] = ~in[56];
  assign inbar[57] = ~in[57];
  assign inbar[58] = ~in[58];
  assign inbar[59] = ~in[59];
  assign inbar[60] = ~in[60];
  assign inbar[61] = ~in[61];
  assign inbar[62] = ~in[62];
  assign inbar[63] = ~in[63];
  assign inbar[64] = ~in[64];
  assign inbar[65] = ~in[65];
  assign inbar[66] = ~in[66];
  assign inbar[67] = ~in[67];
  assign inbar[68] = ~in[68];
  assign inbar[69] = ~in[69];
  assign inbar[70] = ~in[70];
  assign inbar[71] = ~in[71];
  assign inbar[72] = ~in[72];
  assign inbar[73] = ~in[73];
  assign inbar[74] = ~in[74];
  assign inbar[75] = ~in[75];
  assign inbar[76] = ~in[76];
  assign inbar[77] = ~in[77];
  assign inbar[78] = ~in[78];
  assign inbar[79] = ~in[79];
  assign inbar[80] = ~in[80];
  assign inbar[81] = ~in[81];
  assign inbar[82] = ~in[82];
  assign inbar[83] = ~in[83];
  assign inbar[84] = ~in[84];
  assign inbar[85] = ~in[85];
  assign inbar[86] = ~in[86];
  assign inbar[87] = ~in[87];
  assign inbar[88] = ~in[88];
  assign inbar[89] = ~in[89];
  assign inbar[90] = ~in[90];
  assign inbar[91] = ~in[91];
  assign inbar[92] = ~in[92];
  assign inbar[93] = ~in[93];
  assign inbar[94] = ~in[94];
  assign inbar[95] = ~in[95];
  assign inbar[96] = ~in[96];
  assign inbar[97] = ~in[97];
  assign inbar[98] = ~in[98];
  assign inbar[99] = ~in[99];
  assign inbar[100] = ~in[100];
  assign inbar[101] = ~in[101];
  assign inbar[102] = ~in[102];
  assign inbar[103] = ~in[103];
  assign inbar[104] = ~in[104];
  assign inbar[105] = ~in[105];
  assign inbar[106] = ~in[106];
  assign inbar[107] = ~in[107];
  assign inbar[108] = ~in[108];
  assign inbar[109] = ~in[109];
  assign inbar[110] = ~in[110];
  assign inbar[111] = ~in[111];
  assign inbar[112] = ~in[112];
  assign inbar[113] = ~in[113];
  assign inbar[114] = ~in[114];
  assign inbar[115] = ~in[115];
  assign inbar[116] = ~in[116];
  assign inbar[117] = ~in[117];
  assign inbar[118] = ~in[118];
  assign inbar[119] = ~in[119];
  assign inbar[120] = ~in[120];
  assign inbar[121] = ~in[121];
  assign inbar[122] = ~in[122];
  assign inbar[123] = ~in[123];
  assign inbar[124] = ~in[124];
  assign inbar[125] = ~in[125];
  assign inbar[126] = ~in[126];
  assign inbar[127] = ~in[127];
  assign inbar[128] = ~in[128];
  assign inbar[129] = ~in[129];
  assign inbar[130] = ~in[130];
  assign inbar[131] = ~in[131];
  assign inbar[132] = ~in[132];
  assign inbar[133] = ~in[133];
  assign inbar[134] = ~in[134];
  assign inbar[135] = ~in[135];
  assign inbar[136] = ~in[136];
  assign inbar[137] = ~in[137];
  assign inbar[138] = ~in[138];
  assign inbar[139] = ~in[139];
  assign inbar[140] = ~in[140];
  assign inbar[141] = ~in[141];
  assign inbar[142] = ~in[142];
  assign inbar[143] = ~in[143];
  assign inbar[144] = ~in[144];
  assign inbar[145] = ~in[145];
  assign inbar[146] = ~in[146];
  assign inbar[147] = ~in[147];
  assign inbar[148] = ~in[148];
  assign inbar[149] = ~in[149];
  assign inbar[150] = ~in[150];
  assign inbar[151] = ~in[151];
  assign inbar[152] = ~in[152];
  assign inbar[153] = ~in[153];
  assign inbar[154] = ~in[154];
  assign inbar[155] = ~in[155];
  assign inbar[156] = ~in[156];
  assign inbar[157] = ~in[157];
  assign inbar[158] = ~in[158];
  assign inbar[159] = ~in[159];
  assign inbar[160] = ~in[160];
  assign inbar[161] = ~in[161];
  assign inbar[162] = ~in[162];
  assign inbar[163] = ~in[163];
  assign inbar[164] = ~in[164];
  assign inbar[165] = ~in[165];
  assign inbar[166] = ~in[166];
  assign inbar[167] = ~in[167];
  assign inbar[168] = ~in[168];
  assign inbar[169] = ~in[169];
  assign inbar[170] = ~in[170];
  assign inbar[171] = ~in[171];
  assign inbar[172] = ~in[172];
  assign inbar[173] = ~in[173];
  assign inbar[174] = ~in[174];
  assign inbar[175] = ~in[175];
  assign inbar[176] = ~in[176];
  assign inbar[177] = ~in[177];
  assign inbar[178] = ~in[178];
  assign inbar[179] = ~in[179];
  assign inbar[180] = ~in[180];
  assign inbar[181] = ~in[181];
  assign inbar[182] = ~in[182];
  assign inbar[183] = ~in[183];
  assign inbar[184] = ~in[184];
  assign inbar[185] = ~in[185];
  assign inbar[186] = ~in[186];
  assign inbar[187] = ~in[187];
  assign inbar[188] = ~in[188];
  assign inbar[189] = ~in[189];
  assign inbar[190] = ~in[190];
  assign inbar[191] = ~in[191];
  assign inbar[192] = ~in[192];
  assign inbar[193] = ~in[193];
  assign inbar[194] = ~in[194];
  assign inbar[195] = ~in[195];
  assign inbar[196] = ~in[196];
  assign inbar[197] = ~in[197];
  assign inbar[198] = ~in[198];
  assign inbar[199] = ~in[199];
  assign inbar[200] = ~in[200];
  assign inbar[201] = ~in[201];
  assign inbar[202] = ~in[202];
  assign inbar[203] = ~in[203];
  assign inbar[204] = ~in[204];
  assign inbar[205] = ~in[205];
  assign inbar[206] = ~in[206];
  assign inbar[207] = ~in[207];
  assign inbar[208] = ~in[208];
  assign inbar[209] = ~in[209];
  assign inbar[210] = ~in[210];
  assign inbar[211] = ~in[211];
  assign inbar[212] = ~in[212];
  assign inbar[213] = ~in[213];
  assign inbar[214] = ~in[214];
  assign inbar[215] = ~in[215];
  assign inbar[216] = ~in[216];
  assign inbar[217] = ~in[217];
  assign inbar[218] = ~in[218];
  assign inbar[219] = ~in[219];
  assign inbar[220] = ~in[220];
  assign inbar[221] = ~in[221];
  assign inbar[222] = ~in[222];
  assign inbar[223] = ~in[223];
  assign inbar[224] = ~in[224];
  assign inbar[225] = ~in[225];
  assign inbar[226] = ~in[226];
  assign inbar[227] = ~in[227];
  assign inbar[228] = ~in[228];
  assign inbar[229] = ~in[229];
  assign inbar[230] = ~in[230];
  assign inbar[231] = ~in[231];
  assign inbar[232] = ~in[232];
  assign inbar[233] = ~in[233];
  assign inbar[234] = ~in[234];
  assign inbar[235] = ~in[235];
  assign inbar[236] = ~in[236];
  assign inbar[237] = ~in[237];
  assign inbar[238] = ~in[238];
  assign inbar[239] = ~in[239];
  assign inbar[240] = ~in[240];
  assign inbar[241] = ~in[241];
  assign inbar[242] = ~in[242];
  assign inbar[243] = ~in[243];
  assign inbar[244] = ~in[244];
  assign inbar[245] = ~in[245];
  assign inbar[246] = ~in[246];
  assign inbar[247] = ~in[247];
  assign inbar[248] = ~in[248];
  assign inbar[249] = ~in[249];
  assign inbar[250] = ~in[250];
  assign inbar[251] = ~in[251];
  assign inbar[252] = ~in[252];
  assign inbar[253] = ~in[253];
  assign inbar[254] = ~in[254];
  assign inbar[255] = ~in[255];
//input_done

  output wire [7:0] out;
  wire [7:0] outbar;
//output_done

  wire in_81;
  wire in_80;
  wire in_79;
  wire in_78;
  wire in_77;
  wire in_76;
  wire in_75;
  wire in_74;
  wire in_73;
  wire in_72;
  wire in_71;
  wire in_70;
  wire in_69;
  wire in_68;
  wire in_67;
  wire in_66;
  wire in_65;
  wire in_64;
  wire in_63;
  wire in_62;
  wire in_61;
  wire in_60;
  wire in_59;
  wire in_58;
  wire in_57;
  wire in_56;
  wire in_55;
  wire in_54;
  wire in_53;
  wire in_52;
  wire in_51;
  wire in_50;
  wire in_49;
  wire in_48;
  wire in_47;
  wire in_46;
  wire in_45;
  wire in_44;
  wire in_43;
  wire in_42;
  wire in_41;
  wire in_40;
  wire in_39;
  wire in_38;
  wire in_37;
  wire in_36;
  wire in_35;
  wire in_34;
  wire in_33;
  wire in_32;
  wire in_31;
  wire in_30;
  wire in_29;
  wire in_28;
  wire in_27;
  wire in_26;
  wire in_25;
  wire in_24;
  wire in_23;
  wire in_22;
  wire in_21;
  wire in_20;
  wire in_19;
  wire in_18;
  wire in_17;
  wire in_16;
  wire in_15;
  wire in_14;
  wire in_13;
  wire in_12;
  wire in_11;
  wire in_10;
  wire in_9;
  wire in_8;
  wire in_7;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_3;
  wire in_2;
  wire in_1;
  wire in_0;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire in_81bar;
  wire in_80bar;
  wire in_79bar;
  wire in_78bar;
  wire in_77bar;
  wire in_76bar;
  wire in_75bar;
  wire in_74bar;
  wire in_73bar;
  wire in_72bar;
  wire in_71bar;
  wire in_70bar;
  wire in_69bar;
  wire in_68bar;
  wire in_67bar;
  wire in_66bar;
  wire in_65bar;
  wire in_64bar;
  wire in_63bar;
  wire in_62bar;
  wire in_61bar;
  wire in_60bar;
  wire in_59bar;
  wire in_58bar;
  wire in_57bar;
  wire in_56bar;
  wire in_55bar;
  wire in_54bar;
  wire in_53bar;
  wire in_52bar;
  wire in_51bar;
  wire in_50bar;
  wire in_49bar;
  wire in_48bar;
  wire in_47bar;
  wire in_46bar;
  wire in_45bar;
  wire in_44bar;
  wire in_43bar;
  wire in_42bar;
  wire in_41bar;
  wire in_40bar;
  wire in_39bar;
  wire in_38bar;
  wire in_37bar;
  wire in_36bar;
  wire in_35bar;
  wire in_34bar;
  wire in_33bar;
  wire in_32bar;
  wire in_31bar;
  wire in_30bar;
  wire in_29bar;
  wire in_28bar;
  wire in_27bar;
  wire in_26bar;
  wire in_25bar;
  wire in_24bar;
  wire in_23bar;
  wire in_22bar;
  wire in_21bar;
  wire in_20bar;
  wire in_19bar;
  wire in_18bar;
  wire in_17bar;
  wire in_16bar;
  wire in_15bar;
  wire in_14bar;
  wire in_13bar;
  wire in_12bar;
  wire in_11bar;
  wire in_10bar;
  wire in_9bar;
  wire in_8bar;
  wire in_7bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_3bar;
  wire in_2bar;
  wire in_1bar;
  wire in_0bar;
  wire n487bar;
  wire n488bar;
  wire n489bar;
  wire n490bar;
  wire n491bar;
  wire n492bar;
  wire n493bar;
  wire n494bar;
  wire n495bar;
  wire n496bar;
  wire n497bar;
  wire n498bar;
  wire n499bar;
  wire n500bar;
  wire n501bar;
  wire n502bar;
  wire n503bar;
  wire n504bar;
  wire n505bar;
  wire n506bar;
  wire n507bar;
  wire n508bar;
  wire n509bar;
  wire n510bar;
  wire n511bar;
  wire n512bar;
  wire n513bar;
  wire n514bar;
  wire n515bar;
  wire n516bar;
  wire n517bar;
  wire n518bar;
  wire n519bar;
  wire n520bar;
  wire n521bar;
  wire n522bar;
  wire n523bar;
  wire n524bar;
  wire n525bar;
  wire n526bar;
  wire n527bar;
  wire n528bar;
  wire n529bar;
  wire n530bar;
  wire n531bar;
  wire n532bar;
  wire n533bar;
  wire n534bar;
  wire n535bar;
  wire n536bar;
  wire n537bar;
  wire n538bar;
  wire n539bar;
  wire n540bar;
  wire n541bar;
  wire n542bar;
  wire n543bar;
  wire n544bar;
  wire n545bar;
  wire n546bar;
  wire n547bar;
  wire n548bar;
  wire n549bar;
  wire n550bar;
  wire n551bar;
  wire n552bar;
  wire n553bar;
  wire n554bar;
  wire n555bar;
  wire n556bar;
  wire n557bar;
  wire n558bar;
  wire n559bar;
  wire n560bar;
  wire n561bar;
  wire n562bar;
  wire n563bar;
  wire n564bar;
  wire n565bar;
  wire n566bar;
  wire n567bar;
  wire n568bar;
  wire n569bar;
  wire n570bar;
  wire n571bar;
  wire n572bar;
  wire n573bar;
  wire n574bar;
  wire n575bar;
  wire n576bar;
  wire n577bar;
  wire n578bar;
  wire n579bar;
  wire n580bar;
  wire n581bar;
  wire n582bar;
  wire n583bar;
  wire n584bar;
  wire n585bar;
  wire n586bar;
  wire n587bar;
  wire n588bar;
  wire n589bar;
  wire n590bar;
  wire n591bar;
  wire n592bar;
  wire n593bar;
  wire n594bar;
  wire n595bar;
  wire n596bar;
  wire n597bar;
  wire n598bar;
  wire n599bar;
  wire n600bar;
  wire n601bar;
  wire n602bar;
  wire n603bar;
  wire n604bar;
  wire n605bar;
  wire n606bar;
  wire n607bar;
  wire n608bar;
  wire n609bar;
  wire n610bar;
  wire n611bar;
  wire n612bar;
  wire n613bar;
  wire n614bar;
  wire n615bar;
  wire n616bar;
  wire n617bar;
  wire n618bar;
  wire n619bar;
  wire n620bar;
  wire n621bar;
  wire n622bar;
  wire n623bar;
  wire n624bar;
  wire n625bar;
  wire n626bar;
  wire n627bar;
  wire n628bar;
  wire n629bar;
  wire n630bar;
  wire n631bar;
  wire n632bar;
  wire n633bar;
  wire n634bar;
  wire n635bar;
  wire n636bar;
  wire n637bar;
  wire n638bar;
  wire n639bar;
  wire n640bar;
  wire n641bar;
  wire n642bar;
  wire n643bar;
  wire n644bar;
  wire n645bar;
  wire n646bar;
  wire n647bar;
  wire n648bar;
  wire n649bar;
  wire n650bar;
  wire n651bar;
  wire n652bar;
  wire n653bar;
  wire n654bar;
  wire n655bar;
  wire n656bar;
  wire n657bar;
  wire n658bar;
  wire n659bar;
  wire n660bar;
  wire n661bar;
  wire n662bar;
  wire n663bar;
  wire n664bar;
  wire n665bar;
  wire n666bar;
  wire n667bar;
  wire n668bar;
  wire n669bar;
  wire n670bar;
  wire n671bar;
  wire n672bar;
  wire n673bar;
  wire n674bar;
  wire n675bar;
  wire n676bar;
  wire n677bar;
  wire n678bar;
  wire n679bar;
  wire n680bar;
  wire n681bar;
  wire n682bar;
  wire n683bar;
  wire n684bar;
  wire n685bar;
  wire n686bar;
  wire n687bar;
  wire n688bar;
  wire n689bar;
  wire n690bar;
  wire n691bar;
  wire n692bar;
  wire n693bar;
  wire n694bar;
  wire n695bar;
  wire n696bar;
  wire n697bar;
  wire n698bar;
  wire n699bar;
  wire n700bar;
  wire n701bar;
  wire n702bar;
  wire n703bar;
  wire n704bar;
  wire n705bar;
  wire n706bar;
  wire n707bar;
  wire n708bar;
  wire n709bar;
  wire n710bar;
  wire n711bar;
  wire n712bar;
  wire n713bar;
  wire n714bar;
  wire n715bar;
  wire n716bar;
  wire n717bar;
  wire n718bar;
  wire n719bar;
  wire n720bar;
  wire n721bar;
  wire n722bar;
  wire n723bar;
  wire n724bar;
  wire n725bar;
  wire n726bar;
  wire n727bar;
  wire n728bar;
  wire n729bar;
  wire n730bar;
  wire n731bar;
  wire n732bar;
  wire n733bar;
  wire n734bar;
  wire n735bar;
  wire n736bar;
  wire n737bar;
  wire n738bar;
  wire n739bar;
  wire n740bar;
  wire n741bar;
  wire n742bar;
  wire n743bar;
  wire n744bar;
  wire n745bar;
  wire n746bar;
  wire n747bar;
  wire n748bar;
  wire n749bar;
  wire n750bar;
  wire n751bar;
  wire n752bar;
  wire n753bar;
  wire n754bar;
  wire n755bar;
  wire n756bar;
  wire n757bar;
  wire n758bar;
  wire n759bar;
  wire n760bar;
  wire n761bar;
  wire n762bar;
  wire n763bar;
  wire n764bar;
  wire n765bar;
  wire n766bar;
  wire n767bar;
  wire n768bar;
  wire n769bar;
  wire n770bar;
  wire n771bar;
  wire n772bar;
  wire n773bar;
  wire n774bar;
  wire n775bar;
  wire n776bar;
  wire n777bar;
  wire n778bar;
  wire n779bar;
  wire n780bar;
  wire n781bar;
  wire n782bar;
  wire n783bar;
  wire n784bar;
  wire n785bar;
  wire n786bar;
  wire n787bar;
  wire n788bar;
  wire n789bar;
  wire n790bar;
  wire n791bar;
  wire n792bar;
  wire n793bar;
  wire n794bar;
  wire n795bar;
  wire n796bar;
  wire n797bar;
  wire n798bar;
  wire n799bar;
  wire n800bar;
  wire n801bar;
  wire n802bar;
  wire n803bar;
  wire n804bar;
  wire n805bar;
  wire n806bar;
  wire n807bar;
  wire n808bar;
  wire n809bar;
  wire n810bar;
  wire n811bar;
  wire n812bar;
  wire n813bar;
  wire n814bar;
  wire n815bar;
  wire n816bar;
  wire n817bar;
  wire n818bar;
  wire n819bar;
  wire n820bar;
  wire n821bar;
  wire n822bar;
  wire n823bar;
  wire n824bar;
  wire n825bar;
  wire n826bar;
  wire n827bar;
  wire n828bar;
  wire n829bar;
  wire n830bar;
  wire n831bar;
  wire n832bar;
  wire n833bar;
  wire n834bar;
  wire n835bar;
  wire n836bar;
  wire n837bar;
  wire n838bar;
  wire n839bar;
  wire n840bar;
  wire n841bar;
  wire n842bar;
  wire n843bar;
  wire n844bar;
  wire n845bar;
  wire n846bar;
  wire n847bar;
  wire n848bar;
  wire n849bar;
  wire n850bar;
  wire n851bar;
  wire n852bar;
  wire n853bar;
  wire n854bar;
  wire n855bar;
  wire n856bar;
  wire n857bar;
  wire n858bar;
  wire n859bar;
  wire n860bar;
  wire n861bar;
  wire n862bar;
  wire n863bar;
  wire n864bar;
  wire n865bar;
  wire n866bar;
  wire n867bar;
  wire n868bar;
  wire n869bar;
  wire n870bar;
  wire n871bar;
  wire n872bar;
  wire n873bar;
  wire n874bar;
  wire n875bar;
  wire n876bar;
  wire n877bar;
  wire n878bar;
  wire n879bar;
  wire n880bar;
  wire n881bar;
  wire n882bar;
  wire n883bar;
  wire n884bar;
  wire n885bar;
  wire n886bar;
  wire n887bar;
  wire n888bar;
  wire n889bar;
  wire n890bar;
  wire n891bar;
  wire n892bar;
  wire n893bar;
  wire n894bar;
  wire n895bar;
  wire n896bar;
  wire n897bar;
  wire n898bar;
  wire n899bar;
  wire n900bar;
  wire n901bar;
  wire n902bar;
  wire n903bar;
  wire n904bar;
  wire n905bar;
  wire n906bar;
  wire n907bar;
  wire n908bar;
  wire n909bar;
  wire n910bar;
  wire n911bar;
  wire n912bar;
  wire n913bar;
  wire n914bar;
  wire n915bar;
  wire n916bar;
  wire n917bar;
  wire n918bar;
  wire n919bar;
  wire n920bar;
  wire n921bar;
  wire n922bar;
  wire n923bar;
  wire n924bar;
  wire n925bar;
  wire n926bar;
  wire n927bar;
  wire n928bar;
  wire n929bar;
  wire n930bar;
  wire n931bar;
  wire n932bar;
  wire n933bar;
  wire n934bar;
  wire n935bar;
  wire n936bar;
  wire n937bar;
  wire n938bar;
  wire n939bar;
  wire n940bar;
  wire n941bar;
  wire n942bar;
  wire n943bar;
  wire n944bar;
  wire n945bar;
  wire n946bar;
  wire n947bar;
  wire n948bar;
  wire n949bar;
  wire n950bar;
  wire n951bar;
  wire n952bar;
  wire n953bar;
  wire n954bar;
  wire n955bar;
  wire n956bar;
  wire n957bar;
  wire n958bar;
  wire n959bar;
  wire n960bar;
  wire n961bar;
  wire n962bar;
  wire n963bar;
  wire n964bar;
  wire n965bar;
  wire n966bar;
  wire n967bar;
  wire n968bar;
  wire n969bar;
  wire n970bar;
  wire n971bar;
  wire n972bar;
//wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];
  //OR U1
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1 (
    .O(out[7]),
    .I0(n972),
    .I1(n971)
  );
  //AND U1bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1bar (
    .O(outbar[7]),
    .I0(n972bar),
    .I1(n971bar)
  );
  //OR U2
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2 (
    .O(n971),
    .I0(n970),
    .I1(n969)
  );
  //AND U2bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2bar (
    .O(n971bar),
    .I0(n970bar),
    .I1(n969bar)
  );
  //OR U3
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3 (
    .O(n969),
    .I0(n968),
    .I1(n967)
  );
  //AND U3bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3bar (
    .O(n969bar),
    .I0(n968bar),
    .I1(n967bar)
  );
  //OR U4
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4 (
    .O(n967),
    .I0(n966),
    .I1(n965)
  );
  //AND U4bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4bar (
    .O(n967bar),
    .I0(n966bar),
    .I1(n965bar)
  );
  //OR U5
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5 (
    .O(n968),
    .I0(n964),
    .I1(n963)
  );
  //AND U5bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5bar (
    .O(n968bar),
    .I0(n964bar),
    .I1(n963bar)
  );
  //OR U6
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6 (
    .O(n963),
    .I0(in[116]),
    .I1(n962)
  );
  //AND U6bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6bar (
    .O(n963bar),
    .I0(inbar[116]),
    .I1(n962bar)
  );
  //OR U7
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7 (
    .O(n970),
    .I0(n961),
    .I1(n960)
  );
  //AND U7bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7bar (
    .O(n970bar),
    .I0(n961bar),
    .I1(n960bar)
  );
  //OR U8
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8 (
    .O(n960),
    .I0(in[150]),
    .I1(in[127])
  );
  //AND U8bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8bar (
    .O(n960bar),
    .I0(inbar[150]),
    .I1(inbar[127])
  );
  //OR U9
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9 (
    .O(n961),
    .I0(in[160]),
    .I1(n959)
  );
  //AND U9bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9bar (
    .O(n961bar),
    .I0(inbar[160]),
    .I1(n959bar)
  );
  //OR U10
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10 (
    .O(n959),
    .I0(in[252]),
    .I1(in[168])
  );
  //AND U10bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10bar (
    .O(n959bar),
    .I0(inbar[252]),
    .I1(inbar[168])
  );
  //OR U11
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11 (
    .O(n972),
    .I0(n958),
    .I1(n957)
  );
  //AND U11bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11bar (
    .O(n972bar),
    .I0(n958bar),
    .I1(n957bar)
  );
  //OR U12
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12 (
    .O(n957),
    .I0(n956),
    .I1(n955)
  );
  //AND U12bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12bar (
    .O(n957bar),
    .I0(n956bar),
    .I1(n955bar)
  );
  //OR U13
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13 (
    .O(n955),
    .I0(in_17),
    .I1(in[96])
  );
  //AND U13bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13bar (
    .O(n955bar),
    .I0(in_17bar),
    .I1(inbar[96])
  );
  //OR U14
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14 (
    .O(n956),
    .I0(in_23),
    .I1(n954)
  );
  //AND U14bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14bar (
    .O(n956bar),
    .I0(in_23bar),
    .I1(n954bar)
  );
  //OR U15
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15 (
    .O(n954),
    .I0(in_31),
    .I1(in_26)
  );
  //AND U15bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15bar (
    .O(n954bar),
    .I0(in_31bar),
    .I1(in_26bar)
  );
  //OR U16
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16 (
    .O(n958),
    .I0(n953),
    .I1(n952)
  );
  //AND U16bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16bar (
    .O(n958bar),
    .I0(n953bar),
    .I1(n952bar)
  );
  //OR U17
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U17 (
    .O(n952),
    .I0(in_58),
    .I1(in_4)
  );
  //AND U17bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U17bar (
    .O(n952bar),
    .I0(in_58bar),
    .I1(in_4bar)
  );
  //OR U18
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U18 (
    .O(n953),
    .I0(in_59),
    .I1(n951)
  );
  //AND U18bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U18bar (
    .O(n953bar),
    .I0(in_59bar),
    .I1(n951bar)
  );
  //OR U19
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U19 (
    .O(n951),
    .I0(in_71),
    .I1(in_62)
  );
  //AND U19bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U19bar (
    .O(n951bar),
    .I0(in_71bar),
    .I1(in_62bar)
  );
  //OR U20
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U20 (
    .O(out[6]),
    .I0(n950),
    .I1(n949)
  );
  //AND U20bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U20bar (
    .O(outbar[6]),
    .I0(n950bar),
    .I1(n949bar)
  );
  //OR U21
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U21 (
    .O(n949),
    .I0(n948),
    .I1(n947)
  );
  //AND U21bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U21bar (
    .O(n949bar),
    .I0(n948bar),
    .I1(n947bar)
  );
  //OR U22
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U22 (
    .O(n947),
    .I0(n946),
    .I1(n945)
  );
  //AND U22bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U22bar (
    .O(n947bar),
    .I0(n946bar),
    .I1(n945bar)
  );
  //OR U23
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U23 (
    .O(n945),
    .I0(n944),
    .I1(n943)
  );
  //AND U23bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U23bar (
    .O(n945bar),
    .I0(n944bar),
    .I1(n943bar)
  );
  //OR U24
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U24 (
    .O(n946),
    .I0(n942),
    .I1(n941)
  );
  //AND U24bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U24bar (
    .O(n946bar),
    .I0(n942bar),
    .I1(n941bar)
  );
  //OR U25
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U25 (
    .O(n941),
    .I0(in[101]),
    .I1(n940)
  );
  //AND U25bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U25bar (
    .O(n941bar),
    .I0(inbar[101]),
    .I1(n940bar)
  );
  //OR U26
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U26 (
    .O(n948),
    .I0(n939),
    .I1(n938)
  );
  //AND U26bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U26bar (
    .O(n948bar),
    .I0(n939bar),
    .I1(n938bar)
  );
  //OR U27
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U27 (
    .O(n938),
    .I0(in[114]),
    .I1(in[104])
  );
  //AND U27bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U27bar (
    .O(n938bar),
    .I0(inbar[114]),
    .I1(inbar[104])
  );
  //OR U28
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U28 (
    .O(n939),
    .I0(in[128]),
    .I1(n937)
  );
  //AND U28bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U28bar (
    .O(n939bar),
    .I0(inbar[128]),
    .I1(n937bar)
  );
  //OR U29
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U29 (
    .O(n937),
    .I0(in[136]),
    .I1(in[134])
  );
  //AND U29bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U29bar (
    .O(n937bar),
    .I0(inbar[136]),
    .I1(inbar[134])
  );
  //OR U30
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U30 (
    .O(n950),
    .I0(n936),
    .I1(n935)
  );
  //AND U30bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U30bar (
    .O(n950bar),
    .I0(n936bar),
    .I1(n935bar)
  );
  //OR U31
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U31 (
    .O(n935),
    .I0(n934),
    .I1(n933)
  );
  //AND U31bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U31bar (
    .O(n935bar),
    .I0(n934bar),
    .I1(n933bar)
  );
  //OR U32
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U32 (
    .O(n933),
    .I0(in[177]),
    .I1(in[164])
  );
  //AND U32bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U32bar (
    .O(n933bar),
    .I0(inbar[177]),
    .I1(inbar[164])
  );
  //OR U33
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U33 (
    .O(n934),
    .I0(in[212]),
    .I1(n932)
  );
  //AND U33bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U33bar (
    .O(n934bar),
    .I0(inbar[212]),
    .I1(n932bar)
  );
  //OR U34
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U34 (
    .O(n932),
    .I0(in[248]),
    .I1(in[221])
  );
  //AND U34bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U34bar (
    .O(n932bar),
    .I0(inbar[248]),
    .I1(inbar[221])
  );
  //OR U35
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U35 (
    .O(n936),
    .I0(n931),
    .I1(n930)
  );
  //AND U35bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U35bar (
    .O(n936bar),
    .I0(n931bar),
    .I1(n930bar)
  );
  //OR U36
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U36 (
    .O(n930),
    .I0(in_18),
    .I1(in[93])
  );
  //AND U36bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U36bar (
    .O(n930bar),
    .I0(in_18bar),
    .I1(inbar[93])
  );
  //OR U37
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U37 (
    .O(n931),
    .I0(in_31),
    .I1(n929)
  );
  //AND U37bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U37bar (
    .O(n931bar),
    .I0(in_31bar),
    .I1(n929bar)
  );
  //OR U38
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U38 (
    .O(n929),
    .I0(in_7),
    .I1(in_39)
  );
  //AND U38bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U38bar (
    .O(n929bar),
    .I0(in_7bar),
    .I1(in_39bar)
  );
  //OR U39
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U39 (
    .O(out[5]),
    .I0(n928),
    .I1(n927)
  );
  //AND U39bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U39bar (
    .O(outbar[5]),
    .I0(n928bar),
    .I1(n927bar)
  );
  //OR U40
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U40 (
    .O(n927),
    .I0(n926),
    .I1(n925)
  );
  //AND U40bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U40bar (
    .O(n927bar),
    .I0(n926bar),
    .I1(n925bar)
  );
  //OR U41
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U41 (
    .O(n925),
    .I0(n924),
    .I1(n923)
  );
  //AND U41bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U41bar (
    .O(n925bar),
    .I0(n924bar),
    .I1(n923bar)
  );
  //OR U42
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U42 (
    .O(n923),
    .I0(n922),
    .I1(n921)
  );
  //AND U42bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U42bar (
    .O(n923bar),
    .I0(n922bar),
    .I1(n921bar)
  );
  //OR U43
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U43 (
    .O(n924),
    .I0(n940),
    .I1(n920)
  );
  //AND U43bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U43bar (
    .O(n924bar),
    .I0(n940bar),
    .I1(n920bar)
  );
  //OR U44
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U44 (
    .O(n920),
    .I0(in[111]),
    .I1(n919)
  );
  //AND U44bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U44bar (
    .O(n920bar),
    .I0(inbar[111]),
    .I1(n919bar)
  );
  //OR U45
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U45 (
    .O(n940),
    .I0(n918),
    .I1(n917)
  );
  //AND U45bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U45bar (
    .O(n940bar),
    .I0(n918bar),
    .I1(n917bar)
  );
  //OR U46
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U46 (
    .O(n917),
    .I0(n916),
    .I1(n915)
  );
  //AND U46bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U46bar (
    .O(n917bar),
    .I0(n916bar),
    .I1(n915bar)
  );
  //OR U47
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U47 (
    .O(n915),
    .I0(n914),
    .I1(n913)
  );
  //AND U47bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U47bar (
    .O(n915bar),
    .I0(n914bar),
    .I1(n913bar)
  );
  //OR U48
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U48 (
    .O(n913),
    .I0(in[140]),
    .I1(in[131])
  );
  //AND U48bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U48bar (
    .O(n913bar),
    .I0(inbar[140]),
    .I1(inbar[131])
  );
  //OR U49
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U49 (
    .O(n914),
    .I0(in[160]),
    .I1(in[144])
  );
  //AND U49bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U49bar (
    .O(n914bar),
    .I0(inbar[160]),
    .I1(inbar[144])
  );
  //OR U50
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U50 (
    .O(n916),
    .I0(n912),
    .I1(n911)
  );
  //AND U50bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U50bar (
    .O(n916bar),
    .I0(n912bar),
    .I1(n911bar)
  );
  //OR U51
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U51 (
    .O(n911),
    .I0(in[179]),
    .I1(in[174])
  );
  //AND U51bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U51bar (
    .O(n911bar),
    .I0(inbar[179]),
    .I1(inbar[174])
  );
  //OR U52
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U52 (
    .O(n912),
    .I0(in[188]),
    .I1(in[184])
  );
  //AND U52bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U52bar (
    .O(n912bar),
    .I0(inbar[188]),
    .I1(inbar[184])
  );
  //OR U53
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U53 (
    .O(n918),
    .I0(n910),
    .I1(n909)
  );
  //AND U53bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U53bar (
    .O(n918bar),
    .I0(n910bar),
    .I1(n909bar)
  );
  //OR U54
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U54 (
    .O(n909),
    .I0(n908),
    .I1(n907)
  );
  //AND U54bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U54bar (
    .O(n909bar),
    .I0(n908bar),
    .I1(n907bar)
  );
  //OR U55
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U55 (
    .O(n907),
    .I0(in[216]),
    .I1(in[200])
  );
  //AND U55bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U55bar (
    .O(n907bar),
    .I0(inbar[216]),
    .I1(inbar[200])
  );
  //OR U56
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U56 (
    .O(n908),
    .I0(in[228]),
    .I1(in[224])
  );
  //AND U56bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U56bar (
    .O(n908bar),
    .I0(inbar[228]),
    .I1(inbar[224])
  );
  //OR U57
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U57 (
    .O(n910),
    .I0(n906),
    .I1(n905)
  );
  //AND U57bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U57bar (
    .O(n910bar),
    .I0(n906bar),
    .I1(n905bar)
  );
  //OR U58
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U58 (
    .O(n905),
    .I0(in[247]),
    .I1(in[235])
  );
  //AND U58bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U58bar (
    .O(n905bar),
    .I0(inbar[247]),
    .I1(inbar[235])
  );
  //OR U59
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U59 (
    .O(n906),
    .I0(in_42),
    .I1(in[83])
  );
  //AND U59bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U59bar (
    .O(n906bar),
    .I0(in_42bar),
    .I1(inbar[83])
  );
  //OR U60
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U60 (
    .O(n926),
    .I0(n904),
    .I1(n903)
  );
  //AND U60bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U60bar (
    .O(n926bar),
    .I0(n904bar),
    .I1(n903bar)
  );
  //OR U61
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U61 (
    .O(n903),
    .I0(in[166]),
    .I1(in[123])
  );
  //AND U61bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U61bar (
    .O(n903bar),
    .I0(inbar[166]),
    .I1(inbar[123])
  );
  //OR U62
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U62 (
    .O(n904),
    .I0(in[170]),
    .I1(n902)
  );
  //AND U62bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U62bar (
    .O(n904bar),
    .I0(inbar[170]),
    .I1(n902bar)
  );
  //OR U63
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U63 (
    .O(n902),
    .I0(in[194]),
    .I1(in[183])
  );
  //AND U63bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U63bar (
    .O(n902bar),
    .I0(inbar[194]),
    .I1(inbar[183])
  );
  //OR U64
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U64 (
    .O(n928),
    .I0(n901),
    .I1(n900)
  );
  //AND U64bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U64bar (
    .O(n928bar),
    .I0(n901bar),
    .I1(n900bar)
  );
  //OR U65
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U65 (
    .O(n900),
    .I0(n899),
    .I1(n898)
  );
  //AND U65bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U65bar (
    .O(n900bar),
    .I0(n899bar),
    .I1(n898bar)
  );
  //OR U66
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U66 (
    .O(n898),
    .I0(in[241]),
    .I1(in[238])
  );
  //AND U66bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U66bar (
    .O(n898bar),
    .I0(inbar[241]),
    .I1(inbar[238])
  );
  //OR U67
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U67 (
    .O(n899),
    .I0(in[250]),
    .I1(n897)
  );
  //AND U67bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U67bar (
    .O(n899bar),
    .I0(inbar[250]),
    .I1(n897bar)
  );
  //OR U68
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U68 (
    .O(n897),
    .I0(in_24),
    .I1(in[84])
  );
  //AND U68bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U68bar (
    .O(n897bar),
    .I0(in_24bar),
    .I1(inbar[84])
  );
  //OR U69
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U69 (
    .O(n901),
    .I0(n896),
    .I1(n895)
  );
  //AND U69bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U69bar (
    .O(n901bar),
    .I0(n896bar),
    .I1(n895bar)
  );
  //OR U70
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U70 (
    .O(n895),
    .I0(in_41),
    .I1(in_29)
  );
  //AND U70bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U70bar (
    .O(n895bar),
    .I0(in_41bar),
    .I1(in_29bar)
  );
  //OR U71
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U71 (
    .O(n896),
    .I0(in_66),
    .I1(n894)
  );
  //AND U71bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U71bar (
    .O(n896bar),
    .I0(in_66bar),
    .I1(n894bar)
  );
  //OR U72
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U72 (
    .O(n894),
    .I0(in_76),
    .I1(in_71)
  );
  //AND U72bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U72bar (
    .O(n894bar),
    .I0(in_76bar),
    .I1(in_71bar)
  );
  //OR U73
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U73 (
    .O(out[4]),
    .I0(n893),
    .I1(n892)
  );
  //AND U73bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U73bar (
    .O(outbar[4]),
    .I0(n893bar),
    .I1(n892bar)
  );
  //OR U74
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U74 (
    .O(n892),
    .I0(n891),
    .I1(n890)
  );
  //AND U74bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U74bar (
    .O(n892bar),
    .I0(n891bar),
    .I1(n890bar)
  );
  //OR U75
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U75 (
    .O(n890),
    .I0(n889),
    .I1(n888)
  );
  //AND U75bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U75bar (
    .O(n890bar),
    .I0(n889bar),
    .I1(n888bar)
  );
  //OR U76
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U76 (
    .O(n888),
    .I0(n922),
    .I1(n887)
  );
  //AND U76bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U76bar (
    .O(n888bar),
    .I0(n922bar),
    .I1(n887bar)
  );
  //OR U77
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U77 (
    .O(n922),
    .I0(n886),
    .I1(n885)
  );
  //AND U77bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U77bar (
    .O(n922bar),
    .I0(n886bar),
    .I1(n885bar)
  );
  //OR U78
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U78 (
    .O(n885),
    .I0(n884),
    .I1(n883)
  );
  //AND U78bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U78bar (
    .O(n885bar),
    .I0(n884bar),
    .I1(n883bar)
  );
  //OR U79
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U79 (
    .O(n883),
    .I0(n882),
    .I1(n881)
  );
  //AND U79bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U79bar (
    .O(n883bar),
    .I0(n882bar),
    .I1(n881bar)
  );
  //OR U80
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U80 (
    .O(n881),
    .I0(in[118]),
    .I1(in[109])
  );
  //AND U80bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U80bar (
    .O(n881bar),
    .I0(inbar[118]),
    .I1(inbar[109])
  );
  //OR U81
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U81 (
    .O(n882),
    .I0(in[139]),
    .I1(in[120])
  );
  //AND U81bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U81bar (
    .O(n882bar),
    .I0(inbar[139]),
    .I1(inbar[120])
  );
  //OR U82
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U82 (
    .O(n884),
    .I0(n880),
    .I1(n879)
  );
  //AND U82bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U82bar (
    .O(n884bar),
    .I0(n880bar),
    .I1(n879bar)
  );
  //OR U83
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U83 (
    .O(n879),
    .I0(in[198]),
    .I1(in[154])
  );
  //AND U83bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U83bar (
    .O(n879bar),
    .I0(inbar[198]),
    .I1(inbar[154])
  );
  //OR U84
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U84 (
    .O(n880),
    .I0(in[210]),
    .I1(in[205])
  );
  //AND U84bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U84bar (
    .O(n880bar),
    .I0(inbar[210]),
    .I1(inbar[205])
  );
  //OR U85
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U85 (
    .O(n886),
    .I0(n878),
    .I1(n877)
  );
  //AND U85bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U85bar (
    .O(n886bar),
    .I0(n878bar),
    .I1(n877bar)
  );
  //OR U86
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U86 (
    .O(n877),
    .I0(n876),
    .I1(n875)
  );
  //AND U86bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U86bar (
    .O(n877bar),
    .I0(n876bar),
    .I1(n875bar)
  );
  //OR U87
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U87 (
    .O(n875),
    .I0(in[219]),
    .I1(in[217])
  );
  //AND U87bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U87bar (
    .O(n875bar),
    .I0(inbar[219]),
    .I1(inbar[217])
  );
  //OR U88
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U88 (
    .O(n876),
    .I0(in[86]),
    .I1(in[252])
  );
  //AND U88bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U88bar (
    .O(n876bar),
    .I0(inbar[86]),
    .I1(inbar[252])
  );
  //OR U89
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U89 (
    .O(n878),
    .I0(n874),
    .I1(n873)
  );
  //AND U89bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U89bar (
    .O(n878bar),
    .I0(n874bar),
    .I1(n873bar)
  );
  //OR U90
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U90 (
    .O(n873),
    .I0(in_40),
    .I1(in[91])
  );
  //AND U90bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U90bar (
    .O(n873bar),
    .I0(in_40bar),
    .I1(inbar[91])
  );
  //OR U91
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U91 (
    .O(n874),
    .I0(in_8),
    .I1(in_46)
  );
  //AND U91bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U91bar (
    .O(n874bar),
    .I0(in_8bar),
    .I1(in_46bar)
  );
  //OR U92
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U92 (
    .O(n889),
    .I0(n872),
    .I1(n871)
  );
  //AND U92bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U92bar (
    .O(n889bar),
    .I0(n872bar),
    .I1(n871bar)
  );
  //OR U93
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U93 (
    .O(n871),
    .I0(in[117]),
    .I1(n943)
  );
  //AND U93bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U93bar (
    .O(n871bar),
    .I0(inbar[117]),
    .I1(n943bar)
  );
  //OR U94
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U94 (
    .O(n943),
    .I0(n870),
    .I1(n869)
  );
  //AND U94bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U94bar (
    .O(n943bar),
    .I0(n870bar),
    .I1(n869bar)
  );
  //OR U95
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U95 (
    .O(n869),
    .I0(n868),
    .I1(n867)
  );
  //AND U95bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U95bar (
    .O(n869bar),
    .I0(n868bar),
    .I1(n867bar)
  );
  //OR U96
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U96 (
    .O(n867),
    .I0(n866),
    .I1(n865)
  );
  //AND U96bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U96bar (
    .O(n867bar),
    .I0(n866bar),
    .I1(n865bar)
  );
  //OR U97
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U97 (
    .O(n865),
    .I0(n864),
    .I1(n863)
  );
  //AND U97bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U97bar (
    .O(n865bar),
    .I0(n864bar),
    .I1(n863bar)
  );
  //OR U98
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U98 (
    .O(n866),
    .I0(in[108]),
    .I1(n919)
  );
  //AND U98bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U98bar (
    .O(n866bar),
    .I0(inbar[108]),
    .I1(n919bar)
  );
  //OR U99
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U99 (
    .O(n919),
    .I0(n862),
    .I1(n861)
  );
  //AND U99bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U99bar (
    .O(n919bar),
    .I0(n862bar),
    .I1(n861bar)
  );
  //OR U100
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U100 (
    .O(n861),
    .I0(n860),
    .I1(n859)
  );
  //AND U100bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U100bar (
    .O(n861bar),
    .I0(n860bar),
    .I1(n859bar)
  );
  //OR U101
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U101 (
    .O(n859),
    .I0(n858),
    .I1(n857)
  );
  //AND U101bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U101bar (
    .O(n859bar),
    .I0(n858bar),
    .I1(n857bar)
  );
  //OR U102
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U102 (
    .O(n857),
    .I0(in[119]),
    .I1(in[105])
  );
  //AND U102bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U102bar (
    .O(n857bar),
    .I0(inbar[119]),
    .I1(inbar[105])
  );
  //OR U103
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U103 (
    .O(n858),
    .I0(in[186]),
    .I1(in[175])
  );
  //AND U103bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U103bar (
    .O(n858bar),
    .I0(inbar[186]),
    .I1(inbar[175])
  );
  //OR U104
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U104 (
    .O(n860),
    .I0(n856),
    .I1(n855)
  );
  //AND U104bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U104bar (
    .O(n860bar),
    .I0(n856bar),
    .I1(n855bar)
  );
  //OR U105
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U105 (
    .O(n855),
    .I0(in[202]),
    .I1(in[193])
  );
  //AND U105bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U105bar (
    .O(n855bar),
    .I0(inbar[202]),
    .I1(inbar[193])
  );
  //OR U106
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U106 (
    .O(n856),
    .I0(in[225]),
    .I1(in[208])
  );
  //AND U106bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U106bar (
    .O(n856bar),
    .I0(inbar[225]),
    .I1(inbar[208])
  );
  //OR U107
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U107 (
    .O(n862),
    .I0(n854),
    .I1(n853)
  );
  //AND U107bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U107bar (
    .O(n862bar),
    .I0(n854bar),
    .I1(n853bar)
  );
  //OR U108
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U108 (
    .O(n853),
    .I0(n852),
    .I1(n851)
  );
  //AND U108bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U108bar (
    .O(n853bar),
    .I0(n852bar),
    .I1(n851bar)
  );
  //OR U109
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U109 (
    .O(n851),
    .I0(in_1),
    .I1(in[85])
  );
  //AND U109bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U109bar (
    .O(n851bar),
    .I0(in_1bar),
    .I1(inbar[85])
  );
  //OR U110
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U110 (
    .O(n852),
    .I0(in_23),
    .I1(in_19)
  );
  //AND U110bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U110bar (
    .O(n852bar),
    .I0(in_23bar),
    .I1(in_19bar)
  );
  //OR U111
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U111 (
    .O(n854),
    .I0(n850),
    .I1(n849)
  );
  //AND U111bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U111bar (
    .O(n854bar),
    .I0(n850bar),
    .I1(n849bar)
  );
  //OR U112
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U112 (
    .O(n849),
    .I0(in_43),
    .I1(in_33)
  );
  //AND U112bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U112bar (
    .O(n849bar),
    .I0(in_43bar),
    .I1(in_33bar)
  );
  //OR U113
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U113 (
    .O(n850),
    .I0(in_63),
    .I1(in_44)
  );
  //AND U113bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U113bar (
    .O(n850bar),
    .I0(in_63bar),
    .I1(in_44bar)
  );
  //OR U114
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U114 (
    .O(n868),
    .I0(n848),
    .I1(n847)
  );
  //AND U114bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U114bar (
    .O(n868bar),
    .I0(n848bar),
    .I1(n847bar)
  );
  //OR U115
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U115 (
    .O(n847),
    .I0(in[141]),
    .I1(in[112])
  );
  //AND U115bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U115bar (
    .O(n847bar),
    .I0(inbar[141]),
    .I1(inbar[112])
  );
  //OR U116
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U116 (
    .O(n848),
    .I0(in[147]),
    .I1(n846)
  );
  //AND U116bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U116bar (
    .O(n848bar),
    .I0(inbar[147]),
    .I1(n846bar)
  );
  //OR U117
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U117 (
    .O(n846),
    .I0(in[181]),
    .I1(in[167])
  );
  //AND U117bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U117bar (
    .O(n846bar),
    .I0(inbar[181]),
    .I1(inbar[167])
  );
  //OR U118
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U118 (
    .O(n870),
    .I0(n845),
    .I1(n844)
  );
  //AND U118bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U118bar (
    .O(n870bar),
    .I0(n845bar),
    .I1(n844bar)
  );
  //OR U119
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U119 (
    .O(n844),
    .I0(n843),
    .I1(n842)
  );
  //AND U119bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U119bar (
    .O(n844bar),
    .I0(n843bar),
    .I1(n842bar)
  );
  //OR U120
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U120 (
    .O(n842),
    .I0(in[229]),
    .I1(in[201])
  );
  //AND U120bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U120bar (
    .O(n842bar),
    .I0(inbar[229]),
    .I1(inbar[201])
  );
  //OR U121
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U121 (
    .O(n843),
    .I0(in[237]),
    .I1(n841)
  );
  //AND U121bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U121bar (
    .O(n843bar),
    .I0(inbar[237]),
    .I1(n841bar)
  );
  //OR U122
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U122 (
    .O(n841),
    .I0(in[94]),
    .I1(in[253])
  );
  //AND U122bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U122bar (
    .O(n841bar),
    .I0(inbar[94]),
    .I1(inbar[253])
  );
  //OR U123
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U123 (
    .O(n845),
    .I0(n840),
    .I1(n839)
  );
  //AND U123bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U123bar (
    .O(n845bar),
    .I0(n840bar),
    .I1(n839bar)
  );
  //OR U124
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U124 (
    .O(n839),
    .I0(in_21),
    .I1(in[96])
  );
  //AND U124bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U124bar (
    .O(n839bar),
    .I0(in_21bar),
    .I1(inbar[96])
  );
  //OR U125
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U125 (
    .O(n840),
    .I0(in_25),
    .I1(n838)
  );
  //AND U125bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U125bar (
    .O(n840bar),
    .I0(in_25bar),
    .I1(n838bar)
  );
  //OR U126
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U126 (
    .O(n838),
    .I0(in_81),
    .I1(in_45)
  );
  //AND U126bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U126bar (
    .O(n838bar),
    .I0(in_81bar),
    .I1(in_45bar)
  );
  //OR U127
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U127 (
    .O(n891),
    .I0(n837),
    .I1(n836)
  );
  //AND U127bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U127bar (
    .O(n891bar),
    .I0(n837bar),
    .I1(n836bar)
  );
  //OR U128
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U128 (
    .O(n836),
    .I0(in[142]),
    .I1(in[124])
  );
  //AND U128bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U128bar (
    .O(n836bar),
    .I0(inbar[142]),
    .I1(inbar[124])
  );
  //OR U129
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U129 (
    .O(n837),
    .I0(in[150]),
    .I1(n835)
  );
  //AND U129bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U129bar (
    .O(n837bar),
    .I0(inbar[150]),
    .I1(n835bar)
  );
  //OR U130
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U130 (
    .O(n835),
    .I0(in[172]),
    .I1(in[155])
  );
  //AND U130bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U130bar (
    .O(n835bar),
    .I0(inbar[172]),
    .I1(inbar[155])
  );
  //OR U131
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U131 (
    .O(n893),
    .I0(n834),
    .I1(n833)
  );
  //AND U131bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U131bar (
    .O(n893bar),
    .I0(n834bar),
    .I1(n833bar)
  );
  //OR U132
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U132 (
    .O(n833),
    .I0(n832),
    .I1(n831)
  );
  //AND U132bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U132bar (
    .O(n833bar),
    .I0(n832bar),
    .I1(n831bar)
  );
  //OR U133
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U133 (
    .O(n831),
    .I0(in[196]),
    .I1(in[173])
  );
  //AND U133bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U133bar (
    .O(n831bar),
    .I0(inbar[196]),
    .I1(inbar[173])
  );
  //OR U134
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U134 (
    .O(n832),
    .I0(in[222]),
    .I1(n830)
  );
  //AND U134bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U134bar (
    .O(n832bar),
    .I0(inbar[222]),
    .I1(n830bar)
  );
  //OR U135
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U135 (
    .O(n830),
    .I0(in[227]),
    .I1(in[226])
  );
  //AND U135bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U135bar (
    .O(n830bar),
    .I0(inbar[227]),
    .I1(inbar[226])
  );
  //OR U136
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U136 (
    .O(n834),
    .I0(n829),
    .I1(n828)
  );
  //AND U136bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U136bar (
    .O(n834bar),
    .I0(n829bar),
    .I1(n828bar)
  );
  //OR U137
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U137 (
    .O(n828),
    .I0(in[249]),
    .I1(in[231])
  );
  //AND U137bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U137bar (
    .O(n828bar),
    .I0(inbar[249]),
    .I1(inbar[231])
  );
  //OR U138
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U138 (
    .O(n829),
    .I0(in_28),
    .I1(n827)
  );
  //AND U138bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U138bar (
    .O(n829bar),
    .I0(in_28bar),
    .I1(n827bar)
  );
  //OR U139
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U139 (
    .O(n827),
    .I0(in_52),
    .I1(in_47)
  );
  //AND U139bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U139bar (
    .O(n827bar),
    .I0(in_52bar),
    .I1(in_47bar)
  );
  //OR U140
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U140 (
    .O(out[3]),
    .I0(n826),
    .I1(n825)
  );
  //AND U140bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U140bar (
    .O(outbar[3]),
    .I0(n826bar),
    .I1(n825bar)
  );
  //OR U141
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U141 (
    .O(n825),
    .I0(n824),
    .I1(n823)
  );
  //AND U141bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U141bar (
    .O(n825bar),
    .I0(n824bar),
    .I1(n823bar)
  );
  //OR U142
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U142 (
    .O(n823),
    .I0(n822),
    .I1(n821)
  );
  //AND U142bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U142bar (
    .O(n823bar),
    .I0(n822bar),
    .I1(n821bar)
  );
  //OR U143
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U143 (
    .O(n821),
    .I0(n820),
    .I1(n819)
  );
  //AND U143bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U143bar (
    .O(n821bar),
    .I0(n820bar),
    .I1(n819bar)
  );
  //OR U144
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U144 (
    .O(n822),
    .I0(n964),
    .I1(n818)
  );
  //AND U144bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U144bar (
    .O(n822bar),
    .I0(n964bar),
    .I1(n818bar)
  );
  //OR U145
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U145 (
    .O(n818),
    .I0(in[118]),
    .I1(n817)
  );
  //AND U145bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U145bar (
    .O(n818bar),
    .I0(inbar[118]),
    .I1(n817bar)
  );
  //OR U146
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U146 (
    .O(n964),
    .I0(n816),
    .I1(n815)
  );
  //AND U146bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U146bar (
    .O(n964bar),
    .I0(n816bar),
    .I1(n815bar)
  );
  //OR U147
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U147 (
    .O(n815),
    .I0(n814),
    .I1(n813)
  );
  //AND U147bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U147bar (
    .O(n815bar),
    .I0(n814bar),
    .I1(n813bar)
  );
  //OR U148
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U148 (
    .O(n813),
    .I0(n812),
    .I1(n811)
  );
  //AND U148bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U148bar (
    .O(n813bar),
    .I0(n812bar),
    .I1(n811bar)
  );
  //OR U149
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U149 (
    .O(n811),
    .I0(in[122]),
    .I1(in[111])
  );
  //AND U149bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U149bar (
    .O(n811bar),
    .I0(inbar[122]),
    .I1(inbar[111])
  );
  //OR U150
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U150 (
    .O(n812),
    .I0(in[154]),
    .I1(in[151])
  );
  //AND U150bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U150bar (
    .O(n812bar),
    .I0(inbar[154]),
    .I1(inbar[151])
  );
  //OR U151
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U151 (
    .O(n814),
    .I0(n810),
    .I1(n809)
  );
  //AND U151bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U151bar (
    .O(n814bar),
    .I0(n810bar),
    .I1(n809bar)
  );
  //OR U152
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U152 (
    .O(n809),
    .I0(in[187]),
    .I1(in[177])
  );
  //AND U152bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U152bar (
    .O(n809bar),
    .I0(inbar[187]),
    .I1(inbar[177])
  );
  //OR U153
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U153 (
    .O(n810),
    .I0(in[200]),
    .I1(in[192])
  );
  //AND U153bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U153bar (
    .O(n810bar),
    .I0(inbar[200]),
    .I1(inbar[192])
  );
  //OR U154
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U154 (
    .O(n816),
    .I0(n808),
    .I1(n807)
  );
  //AND U154bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U154bar (
    .O(n816bar),
    .I0(n808bar),
    .I1(n807bar)
  );
  //OR U155
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U155 (
    .O(n807),
    .I0(n806),
    .I1(n805)
  );
  //AND U155bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U155bar (
    .O(n807bar),
    .I0(n806bar),
    .I1(n805bar)
  );
  //OR U156
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U156 (
    .O(n805),
    .I0(in[225]),
    .I1(in[207])
  );
  //AND U156bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U156bar (
    .O(n805bar),
    .I0(inbar[225]),
    .I1(inbar[207])
  );
  //OR U157
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U157 (
    .O(n806),
    .I0(in[98]),
    .I1(in[226])
  );
  //AND U157bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U157bar (
    .O(n806bar),
    .I0(inbar[98]),
    .I1(inbar[226])
  );
  //OR U158
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U158 (
    .O(n808),
    .I0(n804),
    .I1(n803)
  );
  //AND U158bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U158bar (
    .O(n808bar),
    .I0(n804bar),
    .I1(n803bar)
  );
  //OR U159
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U159 (
    .O(n803),
    .I0(in_20),
    .I1(in_16)
  );
  //AND U159bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U159bar (
    .O(n803bar),
    .I0(in_20bar),
    .I1(in_16bar)
  );
  //OR U160
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U160 (
    .O(n804),
    .I0(in_55),
    .I1(in_45)
  );
  //AND U160bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U160bar (
    .O(n804bar),
    .I0(in_55bar),
    .I1(in_45bar)
  );
  //OR U161
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U161 (
    .O(n824),
    .I0(n802),
    .I1(n801)
  );
  //AND U161bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U161bar (
    .O(n824bar),
    .I0(n802bar),
    .I1(n801bar)
  );
  //OR U162
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U162 (
    .O(n801),
    .I0(in[162]),
    .I1(in[149])
  );
  //AND U162bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U162bar (
    .O(n801bar),
    .I0(inbar[162]),
    .I1(inbar[149])
  );
  //OR U163
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U163 (
    .O(n802),
    .I0(in[163]),
    .I1(n800)
  );
  //AND U163bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U163bar (
    .O(n802bar),
    .I0(inbar[163]),
    .I1(n800bar)
  );
  //OR U164
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U164 (
    .O(n800),
    .I0(in[191]),
    .I1(in[189])
  );
  //AND U164bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U164bar (
    .O(n800bar),
    .I0(inbar[191]),
    .I1(inbar[189])
  );
  //OR U165
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U165 (
    .O(n826),
    .I0(n799),
    .I1(n798)
  );
  //AND U165bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U165bar (
    .O(n826bar),
    .I0(n799bar),
    .I1(n798bar)
  );
  //OR U166
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U166 (
    .O(n798),
    .I0(n797),
    .I1(n796)
  );
  //AND U166bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U166bar (
    .O(n798bar),
    .I0(n797bar),
    .I1(n796bar)
  );
  //OR U167
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U167 (
    .O(n796),
    .I0(in[212]),
    .I1(in[193])
  );
  //AND U167bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U167bar (
    .O(n796bar),
    .I0(inbar[212]),
    .I1(inbar[193])
  );
  //OR U168
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U168 (
    .O(n797),
    .I0(in[238]),
    .I1(n795)
  );
  //AND U168bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U168bar (
    .O(n797bar),
    .I0(inbar[238]),
    .I1(n795bar)
  );
  //OR U169
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U169 (
    .O(n795),
    .I0(in[88]),
    .I1(in[247])
  );
  //AND U169bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U169bar (
    .O(n795bar),
    .I0(inbar[88]),
    .I1(inbar[247])
  );
  //OR U170
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U170 (
    .O(n799),
    .I0(n794),
    .I1(n793)
  );
  //AND U170bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U170bar (
    .O(n799bar),
    .I0(n794bar),
    .I1(n793bar)
  );
  //OR U171
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U171 (
    .O(n793),
    .I0(in[94]),
    .I1(in[92])
  );
  //AND U171bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U171bar (
    .O(n793bar),
    .I0(inbar[94]),
    .I1(inbar[92])
  );
  //OR U172
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U172 (
    .O(n794),
    .I0(in_52),
    .I1(n792)
  );
  //AND U172bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U172bar (
    .O(n794bar),
    .I0(in_52bar),
    .I1(n792bar)
  );
  //OR U173
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U173 (
    .O(n792),
    .I0(in_70),
    .I1(in_67)
  );
  //AND U173bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U173bar (
    .O(n792bar),
    .I0(in_70bar),
    .I1(in_67bar)
  );
  //OR U174
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U174 (
    .O(out[2]),
    .I0(n791),
    .I1(n790)
  );
  //AND U174bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U174bar (
    .O(outbar[2]),
    .I0(n791bar),
    .I1(n790bar)
  );
  //OR U175
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U175 (
    .O(n790),
    .I0(n789),
    .I1(n788)
  );
  //AND U175bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U175bar (
    .O(n790bar),
    .I0(n789bar),
    .I1(n788bar)
  );
  //OR U176
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U176 (
    .O(n788),
    .I0(n787),
    .I1(n786)
  );
  //AND U176bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U176bar (
    .O(n788bar),
    .I0(n787bar),
    .I1(n786bar)
  );
  //OR U177
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U177 (
    .O(n786),
    .I0(n819),
    .I1(n785)
  );
  //AND U177bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U177bar (
    .O(n786bar),
    .I0(n819bar),
    .I1(n785bar)
  );
  //OR U178
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U178 (
    .O(n819),
    .I0(n784),
    .I1(n783)
  );
  //AND U178bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U178bar (
    .O(n819bar),
    .I0(n784bar),
    .I1(n783bar)
  );
  //OR U179
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U179 (
    .O(n783),
    .I0(n782),
    .I1(n781)
  );
  //AND U179bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U179bar (
    .O(n783bar),
    .I0(n782bar),
    .I1(n781bar)
  );
  //OR U180
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U180 (
    .O(n781),
    .I0(n780),
    .I1(n779)
  );
  //AND U180bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U180bar (
    .O(n781bar),
    .I0(n780bar),
    .I1(n779bar)
  );
  //OR U181
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U181 (
    .O(n779),
    .I0(n962),
    .I1(n778)
  );
  //AND U181bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U181bar (
    .O(n779bar),
    .I0(n962bar),
    .I1(n778bar)
  );
  //OR U182
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U182 (
    .O(n962),
    .I0(n777),
    .I1(n776)
  );
  //AND U182bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U182bar (
    .O(n962bar),
    .I0(n777bar),
    .I1(n776bar)
  );
  //OR U183
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U183 (
    .O(n776),
    .I0(n775),
    .I1(n774)
  );
  //AND U183bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U183bar (
    .O(n776bar),
    .I0(n775bar),
    .I1(n774bar)
  );
  //OR U184
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U184 (
    .O(n774),
    .I0(n773),
    .I1(n772)
  );
  //AND U184bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U184bar (
    .O(n774bar),
    .I0(n773bar),
    .I1(n772bar)
  );
  //OR U185
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U185 (
    .O(n772),
    .I0(in[131]),
    .I1(in[120])
  );
  //AND U185bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U185bar (
    .O(n772bar),
    .I0(inbar[131]),
    .I1(inbar[120])
  );
  //OR U186
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U186 (
    .O(n773),
    .I0(in[153]),
    .I1(in[147])
  );
  //AND U186bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U186bar (
    .O(n773bar),
    .I0(inbar[153]),
    .I1(inbar[147])
  );
  //OR U187
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U187 (
    .O(n775),
    .I0(n771),
    .I1(n770)
  );
  //AND U187bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U187bar (
    .O(n775bar),
    .I0(n771bar),
    .I1(n770bar)
  );
  //OR U188
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U188 (
    .O(n770),
    .I0(in[170]),
    .I1(in[156])
  );
  //AND U188bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U188bar (
    .O(n770bar),
    .I0(inbar[170]),
    .I1(inbar[156])
  );
  //OR U189
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U189 (
    .O(n771),
    .I0(in[223]),
    .I1(in[190])
  );
  //AND U189bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U189bar (
    .O(n771bar),
    .I0(inbar[223]),
    .I1(inbar[190])
  );
  //OR U190
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U190 (
    .O(n777),
    .I0(n769),
    .I1(n768)
  );
  //AND U190bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U190bar (
    .O(n777bar),
    .I0(n769bar),
    .I1(n768bar)
  );
  //OR U191
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U191 (
    .O(n768),
    .I0(n767),
    .I1(n766)
  );
  //AND U191bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U191bar (
    .O(n768bar),
    .I0(n767bar),
    .I1(n766bar)
  );
  //OR U192
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U192 (
    .O(n766),
    .I0(in[236]),
    .I1(in[230])
  );
  //AND U192bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U192bar (
    .O(n766bar),
    .I0(inbar[236]),
    .I1(inbar[230])
  );
  //OR U193
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U193 (
    .O(n767),
    .I0(in[85]),
    .I1(in[240])
  );
  //AND U193bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U193bar (
    .O(n767bar),
    .I0(inbar[85]),
    .I1(inbar[240])
  );
  //OR U194
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U194 (
    .O(n769),
    .I0(n765),
    .I1(n764)
  );
  //AND U194bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U194bar (
    .O(n769bar),
    .I0(n765bar),
    .I1(n764bar)
  );
  //OR U195
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U195 (
    .O(n764),
    .I0(in_12),
    .I1(in[90])
  );
  //AND U195bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U195bar (
    .O(n764bar),
    .I0(in_12bar),
    .I1(inbar[90])
  );
  //OR U196
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U196 (
    .O(n765),
    .I0(in_39),
    .I1(in_28)
  );
  //AND U196bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U196bar (
    .O(n765bar),
    .I0(in_39bar),
    .I1(in_28bar)
  );
  //OR U197
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U197 (
    .O(n780),
    .I0(in[109]),
    .I1(n763)
  );
  //AND U197bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U197bar (
    .O(n780bar),
    .I0(inbar[109]),
    .I1(n763bar)
  );
  //OR U198
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U198 (
    .O(n782),
    .I0(n762),
    .I1(n761)
  );
  //AND U198bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U198bar (
    .O(n782bar),
    .I0(n762bar),
    .I1(n761bar)
  );
  //OR U199
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U199 (
    .O(n761),
    .I0(in[138]),
    .I1(in[129])
  );
  //AND U199bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U199bar (
    .O(n761bar),
    .I0(inbar[138]),
    .I1(inbar[129])
  );
  //OR U200
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U200 (
    .O(n762),
    .I0(in[157]),
    .I1(n760)
  );
  //AND U200bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U200bar (
    .O(n762bar),
    .I0(inbar[157]),
    .I1(n760bar)
  );
  //OR U201
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U201 (
    .O(n760),
    .I0(in[182]),
    .I1(in[167])
  );
  //AND U201bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U201bar (
    .O(n760bar),
    .I0(inbar[182]),
    .I1(inbar[167])
  );
  //OR U202
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U202 (
    .O(n784),
    .I0(n759),
    .I1(n758)
  );
  //AND U202bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U202bar (
    .O(n784bar),
    .I0(n759bar),
    .I1(n758bar)
  );
  //OR U203
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U203 (
    .O(n758),
    .I0(n757),
    .I1(n756)
  );
  //AND U203bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U203bar (
    .O(n758bar),
    .I0(n757bar),
    .I1(n756bar)
  );
  //OR U204
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U204 (
    .O(n756),
    .I0(in[195]),
    .I1(in[184])
  );
  //AND U204bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U204bar (
    .O(n756bar),
    .I0(inbar[195]),
    .I1(inbar[184])
  );
  //OR U205
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U205 (
    .O(n757),
    .I0(in[196]),
    .I1(n755)
  );
  //AND U205bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U205bar (
    .O(n757bar),
    .I0(inbar[196]),
    .I1(n755bar)
  );
  //OR U206
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U206 (
    .O(n755),
    .I0(in[215]),
    .I1(in[209])
  );
  //AND U206bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U206bar (
    .O(n755bar),
    .I0(inbar[215]),
    .I1(inbar[209])
  );
  //OR U207
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U207 (
    .O(n759),
    .I0(n754),
    .I1(n753)
  );
  //AND U207bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U207bar (
    .O(n759bar),
    .I0(n754bar),
    .I1(n753bar)
  );
  //OR U208
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U208 (
    .O(n753),
    .I0(in[93]),
    .I1(in[233])
  );
  //AND U208bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U208bar (
    .O(n753bar),
    .I0(inbar[93]),
    .I1(inbar[233])
  );
  //OR U209
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U209 (
    .O(n754),
    .I0(in_1),
    .I1(n752)
  );
  //AND U209bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U209bar (
    .O(n754bar),
    .I0(in_1bar),
    .I1(n752bar)
  );
  //OR U210
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U210 (
    .O(n752),
    .I0(in_69),
    .I1(in_66)
  );
  //AND U210bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U210bar (
    .O(n752bar),
    .I0(in_69bar),
    .I1(in_66bar)
  );
  //OR U211
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U211 (
    .O(n787),
    .I0(n966),
    .I1(n751)
  );
  //AND U211bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U211bar (
    .O(n787bar),
    .I0(n966bar),
    .I1(n751bar)
  );
  //OR U212
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U212 (
    .O(n751),
    .I0(in[134]),
    .I1(n750)
  );
  //AND U212bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U212bar (
    .O(n751bar),
    .I0(inbar[134]),
    .I1(n750bar)
  );
  //OR U213
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U213 (
    .O(n966),
    .I0(n749),
    .I1(n748)
  );
  //AND U213bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U213bar (
    .O(n966bar),
    .I0(n749bar),
    .I1(n748bar)
  );
  //OR U214
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U214 (
    .O(n748),
    .I0(n747),
    .I1(n746)
  );
  //AND U214bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U214bar (
    .O(n748bar),
    .I0(n747bar),
    .I1(n746bar)
  );
  //OR U215
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U215 (
    .O(n746),
    .I0(n745),
    .I1(n744)
  );
  //AND U215bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U215bar (
    .O(n746bar),
    .I0(n745bar),
    .I1(n744bar)
  );
  //OR U216
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U216 (
    .O(n744),
    .I0(in[136]),
    .I1(in[121])
  );
  //AND U216bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U216bar (
    .O(n744bar),
    .I0(inbar[136]),
    .I1(inbar[121])
  );
  //OR U217
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U217 (
    .O(n745),
    .I0(in[186]),
    .I1(in[174])
  );
  //AND U217bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U217bar (
    .O(n745bar),
    .I0(inbar[186]),
    .I1(inbar[174])
  );
  //OR U218
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U218 (
    .O(n747),
    .I0(n743),
    .I1(n742)
  );
  //AND U218bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U218bar (
    .O(n747bar),
    .I0(n743bar),
    .I1(n742bar)
  );
  //OR U219
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U219 (
    .O(n742),
    .I0(in[198]),
    .I1(in[197])
  );
  //AND U219bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U219bar (
    .O(n742bar),
    .I0(inbar[198]),
    .I1(inbar[197])
  );
  //OR U220
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U220 (
    .O(n743),
    .I0(in[214]),
    .I1(in[199])
  );
  //AND U220bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U220bar (
    .O(n743bar),
    .I0(inbar[214]),
    .I1(inbar[199])
  );
  //OR U221
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U221 (
    .O(n749),
    .I0(n741),
    .I1(n740)
  );
  //AND U221bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U221bar (
    .O(n749bar),
    .I0(n741bar),
    .I1(n740bar)
  );
  //OR U222
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U222 (
    .O(n740),
    .I0(n739),
    .I1(n738)
  );
  //AND U222bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U222bar (
    .O(n740bar),
    .I0(n739bar),
    .I1(n738bar)
  );
  //OR U223
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U223 (
    .O(n738),
    .I0(in[231]),
    .I1(in[220])
  );
  //AND U223bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U223bar (
    .O(n738bar),
    .I0(inbar[231]),
    .I1(inbar[220])
  );
  //OR U224
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U224 (
    .O(n739),
    .I0(in_25),
    .I1(in[245])
  );
  //AND U224bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U224bar (
    .O(n739bar),
    .I0(in_25bar),
    .I1(inbar[245])
  );
  //OR U225
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U225 (
    .O(n741),
    .I0(n737),
    .I1(n736)
  );
  //AND U225bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U225bar (
    .O(n741bar),
    .I0(n737bar),
    .I1(n736bar)
  );
  //OR U226
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U226 (
    .O(n736),
    .I0(in_53),
    .I1(in_29)
  );
  //AND U226bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U226bar (
    .O(n736bar),
    .I0(in_53bar),
    .I1(in_29bar)
  );
  //OR U227
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U227 (
    .O(n737),
    .I0(in_79),
    .I1(in_74)
  );
  //AND U227bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U227bar (
    .O(n737bar),
    .I0(in_79bar),
    .I1(in_74bar)
  );
  //OR U228
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U228 (
    .O(n789),
    .I0(n735),
    .I1(n734)
  );
  //AND U228bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U228bar (
    .O(n789bar),
    .I0(n735bar),
    .I1(n734bar)
  );
  //OR U229
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U229 (
    .O(n734),
    .I0(in[152]),
    .I1(in[140])
  );
  //AND U229bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U229bar (
    .O(n734bar),
    .I0(inbar[152]),
    .I1(inbar[140])
  );
  //OR U230
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U230 (
    .O(n735),
    .I0(in[155]),
    .I1(n733)
  );
  //AND U230bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U230bar (
    .O(n735bar),
    .I0(inbar[155]),
    .I1(n733bar)
  );
  //OR U231
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U231 (
    .O(n733),
    .I0(in[166]),
    .I1(in[165])
  );
  //AND U231bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U231bar (
    .O(n733bar),
    .I0(inbar[166]),
    .I1(inbar[165])
  );
  //OR U232
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U232 (
    .O(n791),
    .I0(n732),
    .I1(n731)
  );
  //AND U232bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U232bar (
    .O(n791bar),
    .I0(n732bar),
    .I1(n731bar)
  );
  //OR U233
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U233 (
    .O(n731),
    .I0(n730),
    .I1(n729)
  );
  //AND U233bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U233bar (
    .O(n731bar),
    .I0(n730bar),
    .I1(n729bar)
  );
  //OR U234
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U234 (
    .O(n729),
    .I0(in[202]),
    .I1(in[185])
  );
  //AND U234bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U234bar (
    .O(n729bar),
    .I0(inbar[202]),
    .I1(inbar[185])
  );
  //OR U235
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U235 (
    .O(n730),
    .I0(in[211]),
    .I1(n728)
  );
  //AND U235bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U235bar (
    .O(n730bar),
    .I0(inbar[211]),
    .I1(n728bar)
  );
  //OR U236
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U236 (
    .O(n728),
    .I0(in[255]),
    .I1(in[253])
  );
  //AND U236bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U236bar (
    .O(n728bar),
    .I0(inbar[255]),
    .I1(inbar[253])
  );
  //OR U237
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U237 (
    .O(n732),
    .I0(n727),
    .I1(n726)
  );
  //AND U237bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U237bar (
    .O(n732bar),
    .I0(n727bar),
    .I1(n726bar)
  );
  //OR U238
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U238 (
    .O(n726),
    .I0(in_35),
    .I1(in_15)
  );
  //AND U238bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U238bar (
    .O(n726bar),
    .I0(in_35bar),
    .I1(in_15bar)
  );
  //OR U239
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U239 (
    .O(n727),
    .I0(in_36),
    .I1(n725)
  );
  //AND U239bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U239bar (
    .O(n727bar),
    .I0(in_36bar),
    .I1(n725bar)
  );
  //OR U240
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U240 (
    .O(n725),
    .I0(in_48),
    .I1(in_40)
  );
  //AND U240bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U240bar (
    .O(n725bar),
    .I0(in_48bar),
    .I1(in_40bar)
  );
  //OR U241
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U241 (
    .O(out[1]),
    .I0(n724),
    .I1(n723)
  );
  //AND U241bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U241bar (
    .O(outbar[1]),
    .I0(n724bar),
    .I1(n723bar)
  );
  //OR U242
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U242 (
    .O(n723),
    .I0(n722),
    .I1(n721)
  );
  //AND U242bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U242bar (
    .O(n723bar),
    .I0(n722bar),
    .I1(n721bar)
  );
  //OR U243
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U243 (
    .O(n721),
    .I0(n720),
    .I1(n719)
  );
  //AND U243bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U243bar (
    .O(n721bar),
    .I0(n720bar),
    .I1(n719bar)
  );
  //OR U244
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U244 (
    .O(n719),
    .I0(n921),
    .I1(n887)
  );
  //AND U244bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U244bar (
    .O(n719bar),
    .I0(n921bar),
    .I1(n887bar)
  );
  //OR U245
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U245 (
    .O(n887),
    .I0(n718),
    .I1(n717)
  );
  //AND U245bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U245bar (
    .O(n887bar),
    .I0(n718bar),
    .I1(n717bar)
  );
  //OR U246
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U246 (
    .O(n717),
    .I0(n716),
    .I1(n715)
  );
  //AND U246bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U246bar (
    .O(n717bar),
    .I0(n716bar),
    .I1(n715bar)
  );
  //OR U247
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U247 (
    .O(n715),
    .I0(n714),
    .I1(n713)
  );
  //AND U247bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U247bar (
    .O(n715bar),
    .I0(n714bar),
    .I1(n713bar)
  );
  //OR U248
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U248 (
    .O(n713),
    .I0(in[116]),
    .I1(in[110])
  );
  //AND U248bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U248bar (
    .O(n713bar),
    .I0(inbar[116]),
    .I1(inbar[110])
  );
  //OR U249
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U249 (
    .O(n714),
    .I0(in[133]),
    .I1(in[130])
  );
  //AND U249bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U249bar (
    .O(n714bar),
    .I0(inbar[133]),
    .I1(inbar[130])
  );
  //OR U250
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U250 (
    .O(n716),
    .I0(n712),
    .I1(n711)
  );
  //AND U250bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U250bar (
    .O(n716bar),
    .I0(n712bar),
    .I1(n711bar)
  );
  //OR U251
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U251 (
    .O(n711),
    .I0(in[203]),
    .I1(in[135])
  );
  //AND U251bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U251bar (
    .O(n711bar),
    .I0(inbar[203]),
    .I1(inbar[135])
  );
  //OR U252
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U252 (
    .O(n712),
    .I0(in[232]),
    .I1(in[223])
  );
  //AND U252bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U252bar (
    .O(n712bar),
    .I0(inbar[232]),
    .I1(inbar[223])
  );
  //OR U253
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U253 (
    .O(n718),
    .I0(n710),
    .I1(n709)
  );
  //AND U253bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U253bar (
    .O(n718bar),
    .I0(n710bar),
    .I1(n709bar)
  );
  //OR U254
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U254 (
    .O(n709),
    .I0(n708),
    .I1(n707)
  );
  //AND U254bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U254bar (
    .O(n709bar),
    .I0(n708bar),
    .I1(n707bar)
  );
  //OR U255
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U255 (
    .O(n707),
    .I0(in[255]),
    .I1(in[233])
  );
  //AND U255bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U255bar (
    .O(n707bar),
    .I0(inbar[255]),
    .I1(inbar[233])
  );
  //OR U256
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U256 (
    .O(n708),
    .I0(in_53),
    .I1(in_34)
  );
  //AND U256bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U256bar (
    .O(n708bar),
    .I0(in_53bar),
    .I1(in_34bar)
  );
  //OR U257
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U257 (
    .O(n710),
    .I0(n706),
    .I1(n705)
  );
  //AND U257bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U257bar (
    .O(n710bar),
    .I0(n706bar),
    .I1(n705bar)
  );
  //OR U258
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U258 (
    .O(n705),
    .I0(in_57),
    .I1(in_55)
  );
  //AND U258bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U258bar (
    .O(n705bar),
    .I0(in_57bar),
    .I1(in_55bar)
  );
  //OR U259
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U259 (
    .O(n706),
    .I0(in_68),
    .I1(in_67)
  );
  //AND U259bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U259bar (
    .O(n706bar),
    .I0(in_68bar),
    .I1(in_67bar)
  );
  //OR U260
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U260 (
    .O(n921),
    .I0(n704),
    .I1(n703)
  );
  //AND U260bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U260bar (
    .O(n921bar),
    .I0(n704bar),
    .I1(n703bar)
  );
  //OR U261
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U261 (
    .O(n703),
    .I0(n702),
    .I1(n701)
  );
  //AND U261bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U261bar (
    .O(n703bar),
    .I0(n702bar),
    .I1(n701bar)
  );
  //OR U262
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U262 (
    .O(n701),
    .I0(n700),
    .I1(n699)
  );
  //AND U262bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U262bar (
    .O(n701bar),
    .I0(n700bar),
    .I1(n699bar)
  );
  //OR U263
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U263 (
    .O(n699),
    .I0(n944),
    .I1(n872)
  );
  //AND U263bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U263bar (
    .O(n699bar),
    .I0(n944bar),
    .I1(n872bar)
  );
  //OR U264
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U264 (
    .O(n872),
    .I0(n698),
    .I1(n697)
  );
  //AND U264bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U264bar (
    .O(n872bar),
    .I0(n698bar),
    .I1(n697bar)
  );
  //OR U265
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U265 (
    .O(n697),
    .I0(n696),
    .I1(n695)
  );
  //AND U265bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U265bar (
    .O(n697bar),
    .I0(n696bar),
    .I1(n695bar)
  );
  //OR U266
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U266 (
    .O(n695),
    .I0(n694),
    .I1(n693)
  );
  //AND U266bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U266bar (
    .O(n695bar),
    .I0(n694bar),
    .I1(n693bar)
  );
  //OR U267
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U267 (
    .O(n693),
    .I0(in[121]),
    .I1(in[102])
  );
  //AND U267bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U267bar (
    .O(n693bar),
    .I0(inbar[121]),
    .I1(inbar[102])
  );
  //OR U268
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U268 (
    .O(n694),
    .I0(in[162]),
    .I1(in[161])
  );
  //AND U268bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U268bar (
    .O(n694bar),
    .I0(inbar[162]),
    .I1(inbar[161])
  );
  //OR U269
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U269 (
    .O(n696),
    .I0(n692),
    .I1(n691)
  );
  //AND U269bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U269bar (
    .O(n696bar),
    .I0(n692bar),
    .I1(n691bar)
  );
  //OR U270
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U270 (
    .O(n691),
    .I0(in[192]),
    .I1(in[178])
  );
  //AND U270bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U270bar (
    .O(n691bar),
    .I0(inbar[192]),
    .I1(inbar[178])
  );
  //OR U271
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U271 (
    .O(n692),
    .I0(in[244]),
    .I1(in[209])
  );
  //AND U271bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U271bar (
    .O(n692bar),
    .I0(inbar[244]),
    .I1(inbar[209])
  );
  //OR U272
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U272 (
    .O(n698),
    .I0(n690),
    .I1(n689)
  );
  //AND U272bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U272bar (
    .O(n698bar),
    .I0(n690bar),
    .I1(n689bar)
  );
  //OR U273
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U273 (
    .O(n689),
    .I0(n688),
    .I1(n687)
  );
  //AND U273bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U273bar (
    .O(n689bar),
    .I0(n688bar),
    .I1(n687bar)
  );
  //OR U274
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U274 (
    .O(n687),
    .I0(in[90]),
    .I1(in[254])
  );
  //AND U274bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U274bar (
    .O(n687bar),
    .I0(inbar[90]),
    .I1(inbar[254])
  );
  //OR U275
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U275 (
    .O(n688),
    .I0(in_36),
    .I1(in_32)
  );
  //AND U275bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U275bar (
    .O(n688bar),
    .I0(in_36bar),
    .I1(in_32bar)
  );
  //OR U276
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U276 (
    .O(n690),
    .I0(n686),
    .I1(n685)
  );
  //AND U276bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U276bar (
    .O(n690bar),
    .I0(n686bar),
    .I1(n685bar)
  );
  //OR U277
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U277 (
    .O(n685),
    .I0(in_62),
    .I1(in_37)
  );
  //AND U277bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U277bar (
    .O(n685bar),
    .I0(in_62bar),
    .I1(in_37bar)
  );
  //OR U278
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U278 (
    .O(n686),
    .I0(in_75),
    .I1(in_73)
  );
  //AND U278bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U278bar (
    .O(n686bar),
    .I0(in_75bar),
    .I1(in_73bar)
  );
  //OR U279
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U279 (
    .O(n944),
    .I0(n684),
    .I1(n683)
  );
  //AND U279bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U279bar (
    .O(n944bar),
    .I0(n684bar),
    .I1(n683bar)
  );
  //OR U280
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U280 (
    .O(n683),
    .I0(n682),
    .I1(n681)
  );
  //AND U280bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U280bar (
    .O(n683bar),
    .I0(n682bar),
    .I1(n681bar)
  );
  //OR U281
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U281 (
    .O(n681),
    .I0(n680),
    .I1(n679)
  );
  //AND U281bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U281bar (
    .O(n681bar),
    .I0(n680bar),
    .I1(n679bar)
  );
  //OR U282
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U282 (
    .O(n679),
    .I0(in[171]),
    .I1(in[153])
  );
  //AND U282bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U282bar (
    .O(n679bar),
    .I0(inbar[171]),
    .I1(inbar[153])
  );
  //OR U283
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U283 (
    .O(n680),
    .I0(in[187]),
    .I1(in[176])
  );
  //AND U283bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U283bar (
    .O(n680bar),
    .I0(inbar[187]),
    .I1(inbar[176])
  );
  //OR U284
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U284 (
    .O(n682),
    .I0(n678),
    .I1(n677)
  );
  //AND U284bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U284bar (
    .O(n682bar),
    .I0(n678bar),
    .I1(n677bar)
  );
  //OR U285
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U285 (
    .O(n677),
    .I0(in[245]),
    .I1(in[211])
  );
  //AND U285bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U285bar (
    .O(n677bar),
    .I0(inbar[245]),
    .I1(inbar[211])
  );
  //OR U286
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U286 (
    .O(n678),
    .I0(in[97]),
    .I1(in[88])
  );
  //AND U286bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U286bar (
    .O(n678bar),
    .I0(inbar[97]),
    .I1(inbar[88])
  );
  //OR U287
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U287 (
    .O(n684),
    .I0(n676),
    .I1(n675)
  );
  //AND U287bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U287bar (
    .O(n684bar),
    .I0(n676bar),
    .I1(n675bar)
  );
  //OR U288
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U288 (
    .O(n675),
    .I0(n674),
    .I1(n673)
  );
  //AND U288bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U288bar (
    .O(n675bar),
    .I0(n674bar),
    .I1(n673bar)
  );
  //OR U289
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U289 (
    .O(n673),
    .I0(in_10),
    .I1(in_0)
  );
  //AND U289bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U289bar (
    .O(n673bar),
    .I0(in_10bar),
    .I1(in_0bar)
  );
  //OR U290
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U290 (
    .O(n674),
    .I0(in_59),
    .I1(in_5)
  );
  //AND U290bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U290bar (
    .O(n674bar),
    .I0(in_59bar),
    .I1(in_5bar)
  );
  //OR U291
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U291 (
    .O(n676),
    .I0(n672),
    .I1(n671)
  );
  //AND U291bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U291bar (
    .O(n676bar),
    .I0(n672bar),
    .I1(n671bar)
  );
  //OR U292
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U292 (
    .O(n671),
    .I0(in_60),
    .I1(in_6)
  );
  //AND U292bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U292bar (
    .O(n671bar),
    .I0(in_60bar),
    .I1(in_6bar)
  );
  //OR U293
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U293 (
    .O(n672),
    .I0(in_77),
    .I1(in_69)
  );
  //AND U293bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U293bar (
    .O(n672bar),
    .I0(in_77bar),
    .I1(in_69bar)
  );
  //OR U294
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U294 (
    .O(n700),
    .I0(in[113]),
    .I1(n864)
  );
  //AND U294bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U294bar (
    .O(n700bar),
    .I0(inbar[113]),
    .I1(n864bar)
  );
  //OR U295
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U295 (
    .O(n864),
    .I0(n670),
    .I1(n669)
  );
  //AND U295bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U295bar (
    .O(n864bar),
    .I0(n670bar),
    .I1(n669bar)
  );
  //OR U296
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U296 (
    .O(n669),
    .I0(n668),
    .I1(n667)
  );
  //AND U296bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U296bar (
    .O(n669bar),
    .I0(n668bar),
    .I1(n667bar)
  );
  //OR U297
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U297 (
    .O(n667),
    .I0(n666),
    .I1(n665)
  );
  //AND U297bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U297bar (
    .O(n667bar),
    .I0(n666bar),
    .I1(n665bar)
  );
  //OR U298
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U298 (
    .O(n665),
    .I0(in[125]),
    .I1(in[107])
  );
  //AND U298bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U298bar (
    .O(n665bar),
    .I0(inbar[125]),
    .I1(inbar[107])
  );
  //OR U299
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U299 (
    .O(n666),
    .I0(in[138]),
    .I1(in[126])
  );
  //AND U299bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U299bar (
    .O(n666bar),
    .I0(inbar[138]),
    .I1(inbar[126])
  );
  //OR U300
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U300 (
    .O(n668),
    .I0(n664),
    .I1(n663)
  );
  //AND U300bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U300bar (
    .O(n668bar),
    .I0(n664bar),
    .I1(n663bar)
  );
  //OR U301
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U301 (
    .O(n663),
    .I0(in[189]),
    .I1(in[143])
  );
  //AND U301bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U301bar (
    .O(n663bar),
    .I0(inbar[189]),
    .I1(inbar[143])
  );
  //OR U302
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U302 (
    .O(n664),
    .I0(in[99]),
    .I1(in[214])
  );
  //AND U302bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U302bar (
    .O(n664bar),
    .I0(inbar[99]),
    .I1(inbar[214])
  );
  //OR U303
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U303 (
    .O(n670),
    .I0(n662),
    .I1(n661)
  );
  //AND U303bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U303bar (
    .O(n670bar),
    .I0(n662bar),
    .I1(n661bar)
  );
  //OR U304
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U304 (
    .O(n661),
    .I0(n660),
    .I1(n659)
  );
  //AND U304bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U304bar (
    .O(n661bar),
    .I0(n660bar),
    .I1(n659bar)
  );
  //OR U305
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U305 (
    .O(n659),
    .I0(in_15),
    .I1(in_12)
  );
  //AND U305bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U305bar (
    .O(n659bar),
    .I0(in_15bar),
    .I1(in_12bar)
  );
  //OR U306
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U306 (
    .O(n660),
    .I0(in_20),
    .I1(in_2)
  );
  //AND U306bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U306bar (
    .O(n660bar),
    .I0(in_20bar),
    .I1(in_2bar)
  );
  //OR U307
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U307 (
    .O(n662),
    .I0(n658),
    .I1(n657)
  );
  //AND U307bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U307bar (
    .O(n662bar),
    .I0(n658bar),
    .I1(n657bar)
  );
  //OR U308
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U308 (
    .O(n657),
    .I0(in_30),
    .I1(in_3)
  );
  //AND U308bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U308bar (
    .O(n657bar),
    .I0(in_30bar),
    .I1(in_3bar)
  );
  //OR U309
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U309 (
    .O(n658),
    .I0(in_4),
    .I1(in_38)
  );
  //AND U309bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U309bar (
    .O(n658bar),
    .I0(in_4bar),
    .I1(in_38bar)
  );
  //OR U310
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U310 (
    .O(n702),
    .I0(n656),
    .I1(n655)
  );
  //AND U310bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U310bar (
    .O(n702bar),
    .I0(n656bar),
    .I1(n655bar)
  );
  //OR U311
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U311 (
    .O(n655),
    .I0(in[148]),
    .I1(in[137])
  );
  //AND U311bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U311bar (
    .O(n655bar),
    .I0(inbar[148]),
    .I1(inbar[137])
  );
  //OR U312
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U312 (
    .O(n656),
    .I0(in[149]),
    .I1(n654)
  );
  //AND U312bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U312bar (
    .O(n656bar),
    .I0(inbar[149]),
    .I1(n654bar)
  );
  //OR U313
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U313 (
    .O(n654),
    .I0(in[195]),
    .I1(in[190])
  );
  //AND U313bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U313bar (
    .O(n654bar),
    .I0(inbar[195]),
    .I1(inbar[190])
  );
  //OR U314
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U314 (
    .O(n704),
    .I0(n653),
    .I1(n652)
  );
  //AND U314bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U314bar (
    .O(n704bar),
    .I0(n653bar),
    .I1(n652bar)
  );
  //OR U315
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U315 (
    .O(n652),
    .I0(n651),
    .I1(n650)
  );
  //AND U315bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U315bar (
    .O(n652bar),
    .I0(n651bar),
    .I1(n650bar)
  );
  //OR U316
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U316 (
    .O(n650),
    .I0(in[98]),
    .I1(in[197])
  );
  //AND U316bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U316bar (
    .O(n650bar),
    .I0(inbar[98]),
    .I1(inbar[197])
  );
  //OR U317
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U317 (
    .O(n651),
    .I0(in_11),
    .I1(n649)
  );
  //AND U317bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U317bar (
    .O(n651bar),
    .I0(in_11bar),
    .I1(n649bar)
  );
  //OR U318
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U318 (
    .O(n649),
    .I0(in_26),
    .I1(in_14)
  );
  //AND U318bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U318bar (
    .O(n649bar),
    .I0(in_26bar),
    .I1(in_14bar)
  );
  //OR U319
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U319 (
    .O(n653),
    .I0(n648),
    .I1(n647)
  );
  //AND U319bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U319bar (
    .O(n653bar),
    .I0(n648bar),
    .I1(n647bar)
  );
  //OR U320
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U320 (
    .O(n647),
    .I0(in_35),
    .I1(in_27)
  );
  //AND U320bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U320bar (
    .O(n647bar),
    .I0(in_35bar),
    .I1(in_27bar)
  );
  //OR U321
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U321 (
    .O(n648),
    .I0(in_50),
    .I1(n646)
  );
  //AND U321bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U321bar (
    .O(n648bar),
    .I0(in_50bar),
    .I1(n646bar)
  );
  //OR U322
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U322 (
    .O(n646),
    .I0(in_78),
    .I1(in_61)
  );
  //AND U322bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U322bar (
    .O(n646bar),
    .I0(in_78bar),
    .I1(in_61bar)
  );
  //OR U323
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U323 (
    .O(n720),
    .I0(n942),
    .I1(n645)
  );
  //AND U323bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U323bar (
    .O(n720bar),
    .I0(n942bar),
    .I1(n645bar)
  );
  //OR U324
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U324 (
    .O(n645),
    .I0(in[106]),
    .I1(n863)
  );
  //AND U324bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U324bar (
    .O(n645bar),
    .I0(inbar[106]),
    .I1(n863bar)
  );
  //OR U325
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U325 (
    .O(n863),
    .I0(n644),
    .I1(n643)
  );
  //AND U325bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U325bar (
    .O(n863bar),
    .I0(n644bar),
    .I1(n643bar)
  );
  //OR U326
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U326 (
    .O(n643),
    .I0(n642),
    .I1(n641)
  );
  //AND U326bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U326bar (
    .O(n643bar),
    .I0(n642bar),
    .I1(n641bar)
  );
  //OR U327
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U327 (
    .O(n641),
    .I0(n640),
    .I1(n639)
  );
  //AND U327bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U327bar (
    .O(n641bar),
    .I0(n640bar),
    .I1(n639bar)
  );
  //OR U328
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U328 (
    .O(n639),
    .I0(in[127]),
    .I1(in[122])
  );
  //AND U328bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U328bar (
    .O(n639bar),
    .I0(inbar[127]),
    .I1(inbar[122])
  );
  //OR U329
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U329 (
    .O(n640),
    .I0(in[156]),
    .I1(in[132])
  );
  //AND U329bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U329bar (
    .O(n640bar),
    .I0(inbar[156]),
    .I1(inbar[132])
  );
  //OR U330
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U330 (
    .O(n642),
    .I0(n638),
    .I1(n637)
  );
  //AND U330bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U330bar (
    .O(n642bar),
    .I0(n638bar),
    .I1(n637bar)
  );
  //OR U331
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U331 (
    .O(n637),
    .I0(in[159]),
    .I1(in[157])
  );
  //AND U331bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U331bar (
    .O(n637bar),
    .I0(inbar[159]),
    .I1(inbar[157])
  );
  //OR U332
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U332 (
    .O(n638),
    .I0(in[185]),
    .I1(in[169])
  );
  //AND U332bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U332bar (
    .O(n638bar),
    .I0(inbar[185]),
    .I1(inbar[169])
  );
  //OR U333
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U333 (
    .O(n644),
    .I0(n636),
    .I1(n635)
  );
  //AND U333bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U333bar (
    .O(n644bar),
    .I0(n636bar),
    .I1(n635bar)
  );
  //OR U334
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U334 (
    .O(n635),
    .I0(n634),
    .I1(n633)
  );
  //AND U334bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U334bar (
    .O(n635bar),
    .I0(n634bar),
    .I1(n633bar)
  );
  //OR U335
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U335 (
    .O(n633),
    .I0(in[239]),
    .I1(in[218])
  );
  //AND U335bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U335bar (
    .O(n633bar),
    .I0(inbar[239]),
    .I1(inbar[218])
  );
  //OR U336
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U336 (
    .O(n634),
    .I0(in_13),
    .I1(in[87])
  );
  //AND U336bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U336bar (
    .O(n634bar),
    .I0(in_13bar),
    .I1(inbar[87])
  );
  //OR U337
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U337 (
    .O(n636),
    .I0(n632),
    .I1(n631)
  );
  //AND U337bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U337bar (
    .O(n636bar),
    .I0(n632bar),
    .I1(n631bar)
  );
  //OR U338
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U338 (
    .O(n631),
    .I0(in_72),
    .I1(in_70)
  );
  //AND U338bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U338bar (
    .O(n631bar),
    .I0(in_72bar),
    .I1(in_70bar)
  );
  //OR U339
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U339 (
    .O(n632),
    .I0(in_80),
    .I1(in_74)
  );
  //AND U339bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U339bar (
    .O(n632bar),
    .I0(in_80bar),
    .I1(in_74bar)
  );
  //OR U340
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U340 (
    .O(n942),
    .I0(n630),
    .I1(n629)
  );
  //AND U340bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U340bar (
    .O(n942bar),
    .I0(n630bar),
    .I1(n629bar)
  );
  //OR U341
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U341 (
    .O(n629),
    .I0(n628),
    .I1(n627)
  );
  //AND U341bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U341bar (
    .O(n629bar),
    .I0(n628bar),
    .I1(n627bar)
  );
  //OR U342
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U342 (
    .O(n627),
    .I0(n626),
    .I1(n625)
  );
  //AND U342bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U342bar (
    .O(n627bar),
    .I0(n626bar),
    .I1(n625bar)
  );
  //OR U343
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U343 (
    .O(n625),
    .I0(in[146]),
    .I1(in[100])
  );
  //AND U343bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U343bar (
    .O(n625bar),
    .I0(inbar[146]),
    .I1(inbar[100])
  );
  //OR U344
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U344 (
    .O(n626),
    .I0(in[168]),
    .I1(in[152])
  );
  //AND U344bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U344bar (
    .O(n626bar),
    .I0(inbar[168]),
    .I1(inbar[152])
  );
  //OR U345
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U345 (
    .O(n628),
    .I0(n624),
    .I1(n623)
  );
  //AND U345bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U345bar (
    .O(n628bar),
    .I0(n624bar),
    .I1(n623bar)
  );
  //OR U346
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U346 (
    .O(n623),
    .I0(in[199]),
    .I1(in[182])
  );
  //AND U346bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U346bar (
    .O(n623bar),
    .I0(inbar[199]),
    .I1(inbar[182])
  );
  //OR U347
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U347 (
    .O(n624),
    .I0(in[236]),
    .I1(in[204])
  );
  //AND U347bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U347bar (
    .O(n624bar),
    .I0(inbar[236]),
    .I1(inbar[204])
  );
  //OR U348
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U348 (
    .O(n630),
    .I0(n622),
    .I1(n621)
  );
  //AND U348bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U348bar (
    .O(n630bar),
    .I0(n622bar),
    .I1(n621bar)
  );
  //OR U349
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U349 (
    .O(n621),
    .I0(n620),
    .I1(n619)
  );
  //AND U349bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U349bar (
    .O(n621bar),
    .I0(n620bar),
    .I1(n619bar)
  );
  //OR U350
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U350 (
    .O(n619),
    .I0(in[89]),
    .I1(in[246])
  );
  //AND U350bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U350bar (
    .O(n619bar),
    .I0(inbar[89]),
    .I1(inbar[246])
  );
  //OR U351
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U351 (
    .O(n620),
    .I0(in[95]),
    .I1(in[92])
  );
  //AND U351bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U351bar (
    .O(n620bar),
    .I0(inbar[95]),
    .I1(inbar[92])
  );
  //OR U352
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U352 (
    .O(n622),
    .I0(n618),
    .I1(n617)
  );
  //AND U352bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U352bar (
    .O(n622bar),
    .I0(n618bar),
    .I1(n617bar)
  );
  //OR U353
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U353 (
    .O(n617),
    .I0(in_22),
    .I1(in_16)
  );
  //AND U353bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U353bar (
    .O(n617bar),
    .I0(in_22bar),
    .I1(in_16bar)
  );
  //OR U354
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U354 (
    .O(n618),
    .I0(in_51),
    .I1(in_49)
  );
  //AND U354bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U354bar (
    .O(n618bar),
    .I0(in_51bar),
    .I1(in_49bar)
  );
  //OR U355
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U355 (
    .O(n722),
    .I0(n616),
    .I1(n615)
  );
  //AND U355bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U355bar (
    .O(n722bar),
    .I0(n616bar),
    .I1(n615bar)
  );
  //OR U356
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U356 (
    .O(n615),
    .I0(in[158]),
    .I1(in[115])
  );
  //AND U356bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U356bar (
    .O(n615bar),
    .I0(inbar[158]),
    .I1(inbar[115])
  );
  //OR U357
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U357 (
    .O(n616),
    .I0(in[163]),
    .I1(n614)
  );
  //AND U357bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U357bar (
    .O(n616bar),
    .I0(inbar[163]),
    .I1(n614bar)
  );
  //OR U358
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U358 (
    .O(n614),
    .I0(in[206]),
    .I1(in[165])
  );
  //AND U358bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U358bar (
    .O(n614bar),
    .I0(inbar[206]),
    .I1(inbar[165])
  );
  //OR U359
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U359 (
    .O(n724),
    .I0(n613),
    .I1(n612)
  );
  //AND U359bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U359bar (
    .O(n724bar),
    .I0(n613bar),
    .I1(n612bar)
  );
  //OR U360
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U360 (
    .O(n612),
    .I0(n611),
    .I1(n610)
  );
  //AND U360bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U360bar (
    .O(n612bar),
    .I0(n611bar),
    .I1(n610bar)
  );
  //OR U361
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U361 (
    .O(n610),
    .I0(in[213]),
    .I1(in[207])
  );
  //AND U361bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U361bar (
    .O(n610bar),
    .I0(inbar[213]),
    .I1(inbar[207])
  );
  //OR U362
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U362 (
    .O(n611),
    .I0(in[215]),
    .I1(n609)
  );
  //AND U362bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U362bar (
    .O(n611bar),
    .I0(inbar[215]),
    .I1(n609bar)
  );
  //OR U363
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U363 (
    .O(n609),
    .I0(in[230]),
    .I1(in[220])
  );
  //AND U363bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U363bar (
    .O(n609bar),
    .I0(inbar[230]),
    .I1(inbar[220])
  );
  //OR U364
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U364 (
    .O(n613),
    .I0(n608),
    .I1(n607)
  );
  //AND U364bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U364bar (
    .O(n613bar),
    .I0(n608bar),
    .I1(n607bar)
  );
  //OR U365
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U365 (
    .O(n607),
    .I0(in[251]),
    .I1(in[234])
  );
  //AND U365bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U365bar (
    .O(n607bar),
    .I0(inbar[251]),
    .I1(inbar[234])
  );
  //OR U366
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U366 (
    .O(n608),
    .I0(in_17),
    .I1(n606)
  );
  //AND U366bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U366bar (
    .O(n608bar),
    .I0(in_17bar),
    .I1(n606bar)
  );
  //OR U367
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U367 (
    .O(n606),
    .I0(in_65),
    .I1(in_56)
  );
  //AND U367bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U367bar (
    .O(n606bar),
    .I0(in_65bar),
    .I1(in_56bar)
  );
  //OR U368
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U368 (
    .O(out[0]),
    .I0(n605),
    .I1(n604)
  );
  //AND U368bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U368bar (
    .O(outbar[0]),
    .I0(n605bar),
    .I1(n604bar)
  );
  //OR U369
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U369 (
    .O(n604),
    .I0(n603),
    .I1(n602)
  );
  //AND U369bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U369bar (
    .O(n604bar),
    .I0(n603bar),
    .I1(n602bar)
  );
  //OR U370
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U370 (
    .O(n602),
    .I0(n601),
    .I1(n600)
  );
  //AND U370bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U370bar (
    .O(n602bar),
    .I0(n601bar),
    .I1(n600bar)
  );
  //OR U371
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U371 (
    .O(n600),
    .I0(n820),
    .I1(n785)
  );
  //AND U371bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U371bar (
    .O(n600bar),
    .I0(n820bar),
    .I1(n785bar)
  );
  //OR U372
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U372 (
    .O(n785),
    .I0(n599),
    .I1(n598)
  );
  //AND U372bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U372bar (
    .O(n785bar),
    .I0(n599bar),
    .I1(n598bar)
  );
  //OR U373
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U373 (
    .O(n598),
    .I0(n597),
    .I1(n596)
  );
  //AND U373bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U373bar (
    .O(n598bar),
    .I0(n597bar),
    .I1(n596bar)
  );
  //OR U374
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U374 (
    .O(n596),
    .I0(n595),
    .I1(n594)
  );
  //AND U374bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U374bar (
    .O(n596bar),
    .I0(n595bar),
    .I1(n594bar)
  );
  //OR U375
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U375 (
    .O(n594),
    .I0(in[135]),
    .I1(in[104])
  );
  //AND U375bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U375bar (
    .O(n594bar),
    .I0(inbar[135]),
    .I1(inbar[104])
  );
  //OR U376
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U376 (
    .O(n595),
    .I0(in[188]),
    .I1(in[178])
  );
  //AND U376bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U376bar (
    .O(n595bar),
    .I0(inbar[188]),
    .I1(inbar[178])
  );
  //OR U377
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U377 (
    .O(n597),
    .I0(n593),
    .I1(n592)
  );
  //AND U377bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U377bar (
    .O(n597bar),
    .I0(n593bar),
    .I1(n592bar)
  );
  //OR U378
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U378 (
    .O(n592),
    .I0(in[217]),
    .I1(in[194])
  );
  //AND U378bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U378bar (
    .O(n592bar),
    .I0(inbar[217]),
    .I1(inbar[194])
  );
  //OR U379
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U379 (
    .O(n593),
    .I0(in[237]),
    .I1(in[218])
  );
  //AND U379bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U379bar (
    .O(n593bar),
    .I0(inbar[237]),
    .I1(inbar[218])
  );
  //OR U380
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U380 (
    .O(n599),
    .I0(n591),
    .I1(n590)
  );
  //AND U380bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U380bar (
    .O(n599bar),
    .I0(n591bar),
    .I1(n590bar)
  );
  //OR U381
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U381 (
    .O(n590),
    .I0(n589),
    .I1(n588)
  );
  //AND U381bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U381bar (
    .O(n590bar),
    .I0(n589bar),
    .I1(n588bar)
  );
  //OR U382
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U382 (
    .O(n588),
    .I0(in_2),
    .I1(in_10)
  );
  //AND U382bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U382bar (
    .O(n588bar),
    .I0(in_2bar),
    .I1(in_10bar)
  );
  //OR U383
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U383 (
    .O(n589),
    .I0(in_47),
    .I1(in_22)
  );
  //AND U383bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U383bar (
    .O(n589bar),
    .I0(in_47bar),
    .I1(in_22bar)
  );
  //OR U384
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U384 (
    .O(n591),
    .I0(n587),
    .I1(n586)
  );
  //AND U384bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U384bar (
    .O(n591bar),
    .I0(n587bar),
    .I1(n586bar)
  );
  //OR U385
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U385 (
    .O(n586),
    .I0(in_56),
    .I1(in_54)
  );
  //AND U385bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U385bar (
    .O(n586bar),
    .I0(in_56bar),
    .I1(in_54bar)
  );
  //OR U386
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U386 (
    .O(n587),
    .I0(in_63),
    .I1(in_61)
  );
  //AND U386bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U386bar (
    .O(n587bar),
    .I0(in_63bar),
    .I1(in_61bar)
  );
  //OR U387
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U387 (
    .O(n820),
    .I0(n585),
    .I1(n584)
  );
  //AND U387bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U387bar (
    .O(n820bar),
    .I0(n585bar),
    .I1(n584bar)
  );
  //OR U388
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U388 (
    .O(n584),
    .I0(n583),
    .I1(n582)
  );
  //AND U388bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U388bar (
    .O(n584bar),
    .I0(n583bar),
    .I1(n582bar)
  );
  //OR U389
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U389 (
    .O(n582),
    .I0(n581),
    .I1(n580)
  );
  //AND U389bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U389bar (
    .O(n582bar),
    .I0(n581bar),
    .I1(n580bar)
  );
  //OR U390
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U390 (
    .O(n580),
    .I0(in[158]),
    .I1(in[142])
  );
  //AND U390bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U390bar (
    .O(n580bar),
    .I0(inbar[158]),
    .I1(inbar[142])
  );
  //OR U391
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U391 (
    .O(n581),
    .I0(in[175]),
    .I1(in[164])
  );
  //AND U391bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U391bar (
    .O(n581bar),
    .I0(inbar[175]),
    .I1(inbar[164])
  );
  //OR U392
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U392 (
    .O(n583),
    .I0(n579),
    .I1(n578)
  );
  //AND U392bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U392bar (
    .O(n583bar),
    .I0(n579bar),
    .I1(n578bar)
  );
  //OR U393
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U393 (
    .O(n578),
    .I0(in[228]),
    .I1(in[204])
  );
  //AND U393bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U393bar (
    .O(n578bar),
    .I0(inbar[228]),
    .I1(inbar[204])
  );
  //OR U394
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U394 (
    .O(n579),
    .I0(in[91]),
    .I1(in[87])
  );
  //AND U394bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U394bar (
    .O(n579bar),
    .I0(inbar[91]),
    .I1(inbar[87])
  );
  //OR U395
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U395 (
    .O(n585),
    .I0(n577),
    .I1(n576)
  );
  //AND U395bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U395bar (
    .O(n585bar),
    .I0(n577bar),
    .I1(n576bar)
  );
  //OR U396
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U396 (
    .O(n576),
    .I0(n575),
    .I1(n574)
  );
  //AND U396bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U396bar (
    .O(n576bar),
    .I0(n575bar),
    .I1(n574bar)
  );
  //OR U397
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U397 (
    .O(n574),
    .I0(in_21),
    .I1(in_11)
  );
  //AND U397bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U397bar (
    .O(n574bar),
    .I0(in_21bar),
    .I1(in_11bar)
  );
  //OR U398
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U398 (
    .O(n575),
    .I0(in_5),
    .I1(in_3)
  );
  //AND U398bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U398bar (
    .O(n575bar),
    .I0(in_5bar),
    .I1(in_3bar)
  );
  //OR U399
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U399 (
    .O(n577),
    .I0(n573),
    .I1(n572)
  );
  //AND U399bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U399bar (
    .O(n577bar),
    .I0(n573bar),
    .I1(n572bar)
  );
  //OR U400
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U400 (
    .O(n572),
    .I0(in_68),
    .I1(in_64)
  );
  //AND U400bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U400bar (
    .O(n572bar),
    .I0(in_68bar),
    .I1(in_64bar)
  );
  //OR U401
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U401 (
    .O(n573),
    .I0(in_76),
    .I1(in_73)
  );
  //AND U401bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U401bar (
    .O(n573bar),
    .I0(in_76bar),
    .I1(in_73bar)
  );
  //OR U402
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U402 (
    .O(n601),
    .I0(n778),
    .I1(n571)
  );
  //AND U402bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U402bar (
    .O(n601bar),
    .I0(n778bar),
    .I1(n571bar)
  );
  //OR U403
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U403 (
    .O(n571),
    .I0(in[100]),
    .I1(n965)
  );
  //AND U403bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U403bar (
    .O(n571bar),
    .I0(inbar[100]),
    .I1(n965bar)
  );
  //OR U404
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U404 (
    .O(n965),
    .I0(n570),
    .I1(n569)
  );
  //AND U404bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U404bar (
    .O(n965bar),
    .I0(n570bar),
    .I1(n569bar)
  );
  //OR U405
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U405 (
    .O(n569),
    .I0(n568),
    .I1(n567)
  );
  //AND U405bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U405bar (
    .O(n569bar),
    .I0(n568bar),
    .I1(n567bar)
  );
  //OR U406
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U406 (
    .O(n567),
    .I0(n566),
    .I1(n565)
  );
  //AND U406bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U406bar (
    .O(n567bar),
    .I0(n566bar),
    .I1(n565bar)
  );
  //OR U407
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U407 (
    .O(n565),
    .I0(n817),
    .I1(n750)
  );
  //AND U407bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U407bar (
    .O(n565bar),
    .I0(n817bar),
    .I1(n750bar)
  );
  //OR U408
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U408 (
    .O(n750),
    .I0(n564),
    .I1(n563)
  );
  //AND U408bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U408bar (
    .O(n750bar),
    .I0(n564bar),
    .I1(n563bar)
  );
  //OR U409
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U409 (
    .O(n563),
    .I0(n562),
    .I1(n561)
  );
  //AND U409bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U409bar (
    .O(n563bar),
    .I0(n562bar),
    .I1(n561bar)
  );
  //OR U410
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U410 (
    .O(n561),
    .I0(n560),
    .I1(n559)
  );
  //AND U410bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U410bar (
    .O(n561bar),
    .I0(n560bar),
    .I1(n559bar)
  );
  //OR U411
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U411 (
    .O(n559),
    .I0(in[119]),
    .I1(in[103])
  );
  //AND U411bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U411bar (
    .O(n559bar),
    .I0(inbar[119]),
    .I1(inbar[103])
  );
  //OR U412
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U412 (
    .O(n560),
    .I0(in[137]),
    .I1(in[133])
  );
  //AND U412bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U412bar (
    .O(n560bar),
    .I0(inbar[137]),
    .I1(inbar[133])
  );
  //OR U413
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U413 (
    .O(n562),
    .I0(n558),
    .I1(n557)
  );
  //AND U413bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U413bar (
    .O(n562bar),
    .I0(n558bar),
    .I1(n557bar)
  );
  //OR U414
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U414 (
    .O(n557),
    .I0(in[176]),
    .I1(in[173])
  );
  //AND U414bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U414bar (
    .O(n557bar),
    .I0(inbar[176]),
    .I1(inbar[173])
  );
  //OR U415
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U415 (
    .O(n558),
    .I0(in[210]),
    .I1(in[181])
  );
  //AND U415bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U415bar (
    .O(n558bar),
    .I0(inbar[210]),
    .I1(inbar[181])
  );
  //OR U416
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U416 (
    .O(n564),
    .I0(n556),
    .I1(n555)
  );
  //AND U416bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U416bar (
    .O(n564bar),
    .I0(n556bar),
    .I1(n555bar)
  );
  //OR U417
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U417 (
    .O(n555),
    .I0(n554),
    .I1(n553)
  );
  //AND U417bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U417bar (
    .O(n555bar),
    .I0(n554bar),
    .I1(n553bar)
  );
  //OR U418
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U418 (
    .O(n553),
    .I0(in_13),
    .I1(in[234])
  );
  //AND U418bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U418bar (
    .O(n553bar),
    .I0(in_13bar),
    .I1(inbar[234])
  );
  //OR U419
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U419 (
    .O(n554),
    .I0(in_38),
    .I1(in_32)
  );
  //AND U419bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U419bar (
    .O(n554bar),
    .I0(in_38bar),
    .I1(in_32bar)
  );
  //OR U420
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U420 (
    .O(n556),
    .I0(n552),
    .I1(n551)
  );
  //AND U420bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U420bar (
    .O(n556bar),
    .I0(n552bar),
    .I1(n551bar)
  );
  //OR U421
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U421 (
    .O(n551),
    .I0(in_42),
    .I1(in_41)
  );
  //AND U421bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U421bar (
    .O(n551bar),
    .I0(in_42bar),
    .I1(in_41bar)
  );
  //OR U422
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U422 (
    .O(n552),
    .I0(in_7),
    .I1(in_49)
  );
  //AND U422bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U422bar (
    .O(n552bar),
    .I0(in_7bar),
    .I1(in_49bar)
  );
  //OR U423
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U423 (
    .O(n817),
    .I0(n550),
    .I1(n549)
  );
  //AND U423bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U423bar (
    .O(n817bar),
    .I0(n550bar),
    .I1(n549bar)
  );
  //OR U424
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U424 (
    .O(n549),
    .I0(n548),
    .I1(n547)
  );
  //AND U424bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U424bar (
    .O(n549bar),
    .I0(n548bar),
    .I1(n547bar)
  );
  //OR U425
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U425 (
    .O(n547),
    .I0(n546),
    .I1(n545)
  );
  //AND U425bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U425bar (
    .O(n547bar),
    .I0(n546bar),
    .I1(n545bar)
  );
  //OR U426
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U426 (
    .O(n545),
    .I0(in[159]),
    .I1(in[105])
  );
  //AND U426bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U426bar (
    .O(n545bar),
    .I0(inbar[159]),
    .I1(inbar[105])
  );
  //OR U427
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U427 (
    .O(n546),
    .I0(in[206]),
    .I1(in[183])
  );
  //AND U427bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U427bar (
    .O(n546bar),
    .I0(inbar[206]),
    .I1(inbar[183])
  );
  //OR U428
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U428 (
    .O(n548),
    .I0(n544),
    .I1(n543)
  );
  //AND U428bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U428bar (
    .O(n548bar),
    .I0(n544bar),
    .I1(n543bar)
  );
  //OR U429
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U429 (
    .O(n543),
    .I0(in[229]),
    .I1(in[219])
  );
  //AND U429bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U429bar (
    .O(n543bar),
    .I0(inbar[229]),
    .I1(inbar[219])
  );
  //OR U430
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U430 (
    .O(n544),
    .I0(in[235]),
    .I1(in[232])
  );
  //AND U430bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U430bar (
    .O(n544bar),
    .I0(inbar[235]),
    .I1(inbar[232])
  );
  //OR U431
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U431 (
    .O(n550),
    .I0(n542),
    .I1(n541)
  );
  //AND U431bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U431bar (
    .O(n550bar),
    .I0(n542bar),
    .I1(n541bar)
  );
  //OR U432
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U432 (
    .O(n541),
    .I0(n540),
    .I1(n539)
  );
  //AND U432bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U432bar (
    .O(n541bar),
    .I0(n540bar),
    .I1(n539bar)
  );
  //OR U433
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U433 (
    .O(n539),
    .I0(in[249]),
    .I1(in[242])
  );
  //AND U433bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U433bar (
    .O(n539bar),
    .I0(inbar[249]),
    .I1(inbar[242])
  );
  //OR U434
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U434 (
    .O(n540),
    .I0(in[89]),
    .I1(in[254])
  );
  //AND U434bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U434bar (
    .O(n540bar),
    .I0(inbar[89]),
    .I1(inbar[254])
  );
  //OR U435
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U435 (
    .O(n542),
    .I0(n538),
    .I1(n537)
  );
  //AND U435bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U435bar (
    .O(n542bar),
    .I0(n538bar),
    .I1(n537bar)
  );
  //OR U436
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U436 (
    .O(n537),
    .I0(in_14),
    .I1(in[99])
  );
  //AND U436bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U436bar (
    .O(n537bar),
    .I0(in_14bar),
    .I1(inbar[99])
  );
  //OR U437
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U437 (
    .O(n538),
    .I0(in_60),
    .I1(in_18)
  );
  //AND U437bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U437bar (
    .O(n538bar),
    .I0(in_60bar),
    .I1(in_18bar)
  );
  //OR U438
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U438 (
    .O(n566),
    .I0(in[113]),
    .I1(n763)
  );
  //AND U438bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U438bar (
    .O(n566bar),
    .I0(inbar[113]),
    .I1(n763bar)
  );
  //OR U439
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U439 (
    .O(n763),
    .I0(n536),
    .I1(n535)
  );
  //AND U439bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U439bar (
    .O(n763bar),
    .I0(n536bar),
    .I1(n535bar)
  );
  //OR U440
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U440 (
    .O(n535),
    .I0(n534),
    .I1(n533)
  );
  //AND U440bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U440bar (
    .O(n535bar),
    .I0(n534bar),
    .I1(n533bar)
  );
  //OR U441
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U441 (
    .O(n533),
    .I0(n532),
    .I1(n531)
  );
  //AND U441bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U441bar (
    .O(n533bar),
    .I0(n532bar),
    .I1(n531bar)
  );
  //OR U442
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U442 (
    .O(n531),
    .I0(in[115]),
    .I1(in[110])
  );
  //AND U442bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U442bar (
    .O(n531bar),
    .I0(inbar[115]),
    .I1(inbar[110])
  );
  //OR U443
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U443 (
    .O(n532),
    .I0(in[125]),
    .I1(in[117])
  );
  //AND U443bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U443bar (
    .O(n532bar),
    .I0(inbar[125]),
    .I1(inbar[117])
  );
  //OR U444
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U444 (
    .O(n534),
    .I0(n530),
    .I1(n529)
  );
  //AND U444bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U444bar (
    .O(n534bar),
    .I0(n530bar),
    .I1(n529bar)
  );
  //OR U445
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U445 (
    .O(n529),
    .I0(in[180]),
    .I1(in[128])
  );
  //AND U445bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U445bar (
    .O(n529bar),
    .I0(inbar[180]),
    .I1(inbar[128])
  );
  //OR U446
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U446 (
    .O(n530),
    .I0(in[205]),
    .I1(in[201])
  );
  //AND U446bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U446bar (
    .O(n530bar),
    .I0(inbar[205]),
    .I1(inbar[201])
  );
  //OR U447
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U447 (
    .O(n536),
    .I0(n528),
    .I1(n527)
  );
  //AND U447bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U447bar (
    .O(n536bar),
    .I0(n528bar),
    .I1(n527bar)
  );
  //OR U448
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U448 (
    .O(n527),
    .I0(n526),
    .I1(n525)
  );
  //AND U448bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U448bar (
    .O(n527bar),
    .I0(n526bar),
    .I1(n525bar)
  );
  //OR U449
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U449 (
    .O(n525),
    .I0(in[244]),
    .I1(in[239])
  );
  //AND U449bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U449bar (
    .O(n525bar),
    .I0(inbar[244]),
    .I1(inbar[239])
  );
  //OR U450
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U450 (
    .O(n526),
    .I0(in[95]),
    .I1(in[83])
  );
  //AND U450bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U450bar (
    .O(n526bar),
    .I0(inbar[95]),
    .I1(inbar[83])
  );
  //OR U451
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U451 (
    .O(n528),
    .I0(n524),
    .I1(n523)
  );
  //AND U451bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U451bar (
    .O(n528bar),
    .I0(n524bar),
    .I1(n523bar)
  );
  //OR U452
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U452 (
    .O(n523),
    .I0(in_24),
    .I1(in[97])
  );
  //AND U452bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U452bar (
    .O(n523bar),
    .I0(in_24bar),
    .I1(inbar[97])
  );
  //OR U453
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U453 (
    .O(n524),
    .I0(in_33),
    .I1(in_27)
  );
  //AND U453bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U453bar (
    .O(n524bar),
    .I0(in_33bar),
    .I1(in_27bar)
  );
  //OR U454
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U454 (
    .O(n568),
    .I0(n522),
    .I1(n521)
  );
  //AND U454bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U454bar (
    .O(n568bar),
    .I0(n522bar),
    .I1(n521bar)
  );
  //OR U455
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U455 (
    .O(n521),
    .I0(in[145]),
    .I1(in[126])
  );
  //AND U455bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U455bar (
    .O(n521bar),
    .I0(inbar[145]),
    .I1(inbar[126])
  );
  //OR U456
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U456 (
    .O(n522),
    .I0(in[169]),
    .I1(n520)
  );
  //AND U456bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U456bar (
    .O(n522bar),
    .I0(inbar[169]),
    .I1(n520bar)
  );
  //OR U457
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U457 (
    .O(n520),
    .I0(in[221]),
    .I1(in[172])
  );
  //AND U457bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U457bar (
    .O(n520bar),
    .I0(inbar[221]),
    .I1(inbar[172])
  );
  //OR U458
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U458 (
    .O(n570),
    .I0(n519),
    .I1(n518)
  );
  //AND U458bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U458bar (
    .O(n570bar),
    .I0(n519bar),
    .I1(n518bar)
  );
  //OR U459
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U459 (
    .O(n518),
    .I0(n517),
    .I1(n516)
  );
  //AND U459bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U459bar (
    .O(n518bar),
    .I0(n517bar),
    .I1(n516bar)
  );
  //OR U460
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U460 (
    .O(n516),
    .I0(in[241]),
    .I1(in[224])
  );
  //AND U460bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U460bar (
    .O(n516bar),
    .I0(inbar[241]),
    .I1(inbar[224])
  );
  //OR U461
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U461 (
    .O(n517),
    .I0(in[86]),
    .I1(n515)
  );
  //AND U461bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U461bar (
    .O(n517bar),
    .I0(inbar[86]),
    .I1(n515bar)
  );
  //OR U462
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U462 (
    .O(n515),
    .I0(in_43),
    .I1(in_34)
  );
  //AND U462bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U462bar (
    .O(n515bar),
    .I0(in_43bar),
    .I1(in_34bar)
  );
  //OR U463
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U463 (
    .O(n519),
    .I0(n514),
    .I1(n513)
  );
  //AND U463bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U463bar (
    .O(n519bar),
    .I0(n514bar),
    .I1(n513bar)
  );
  //OR U464
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U464 (
    .O(n513),
    .I0(in_65),
    .I1(in_51)
  );
  //AND U464bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U464bar (
    .O(n513bar),
    .I0(in_65bar),
    .I1(in_51bar)
  );
  //OR U465
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U465 (
    .O(n514),
    .I0(in_75),
    .I1(n512)
  );
  //AND U465bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U465bar (
    .O(n514bar),
    .I0(in_75bar),
    .I1(n512bar)
  );
  //OR U466
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U466 (
    .O(n512),
    .I0(in_81),
    .I1(in_77)
  );
  //AND U466bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U466bar (
    .O(n512bar),
    .I0(in_81bar),
    .I1(in_77bar)
  );
  //OR U467
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U467 (
    .O(n778),
    .I0(n511),
    .I1(n510)
  );
  //AND U467bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U467bar (
    .O(n778bar),
    .I0(n511bar),
    .I1(n510bar)
  );
  //OR U468
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U468 (
    .O(n510),
    .I0(n509),
    .I1(n508)
  );
  //AND U468bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U468bar (
    .O(n510bar),
    .I0(n509bar),
    .I1(n508bar)
  );
  //OR U469
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U469 (
    .O(n508),
    .I0(n507),
    .I1(n506)
  );
  //AND U469bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U469bar (
    .O(n508bar),
    .I0(n507bar),
    .I1(n506bar)
  );
  //OR U470
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U470 (
    .O(n506),
    .I0(in[107]),
    .I1(in[101])
  );
  //AND U470bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U470bar (
    .O(n506bar),
    .I0(inbar[107]),
    .I1(inbar[101])
  );
  //OR U471
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U471 (
    .O(n507),
    .I0(in[139]),
    .I1(in[132])
  );
  //AND U471bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U471bar (
    .O(n507bar),
    .I0(inbar[139]),
    .I1(inbar[132])
  );
  //OR U472
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U472 (
    .O(n509),
    .I0(n505),
    .I1(n504)
  );
  //AND U472bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U472bar (
    .O(n509bar),
    .I0(n505bar),
    .I1(n504bar)
  );
  //OR U473
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U473 (
    .O(n504),
    .I0(in[146]),
    .I1(in[141])
  );
  //AND U473bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U473bar (
    .O(n504bar),
    .I0(inbar[146]),
    .I1(inbar[141])
  );
  //OR U474
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U474 (
    .O(n505),
    .I0(in[203]),
    .I1(in[179])
  );
  //AND U474bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U474bar (
    .O(n505bar),
    .I0(inbar[203]),
    .I1(inbar[179])
  );
  //OR U475
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U475 (
    .O(n511),
    .I0(n503),
    .I1(n502)
  );
  //AND U475bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U475bar (
    .O(n511bar),
    .I0(n503bar),
    .I1(n502bar)
  );
  //OR U476
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U476 (
    .O(n502),
    .I0(n501),
    .I1(n500)
  );
  //AND U476bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U476bar (
    .O(n502bar),
    .I0(n501bar),
    .I1(n500bar)
  );
  //OR U477
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U477 (
    .O(n500),
    .I0(in[243]),
    .I1(in[222])
  );
  //AND U477bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U477bar (
    .O(n500bar),
    .I0(inbar[243]),
    .I1(inbar[222])
  );
  //OR U478
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U478 (
    .O(n501),
    .I0(in[251]),
    .I1(in[250])
  );
  //AND U478bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U478bar (
    .O(n501bar),
    .I0(inbar[251]),
    .I1(inbar[250])
  );
  //OR U479
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U479 (
    .O(n503),
    .I0(n499),
    .I1(n498)
  );
  //AND U479bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U479bar (
    .O(n503bar),
    .I0(n499bar),
    .I1(n498bar)
  );
  //OR U480
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U480 (
    .O(n498),
    .I0(in_37),
    .I1(in_19)
  );
  //AND U480bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U480bar (
    .O(n498bar),
    .I0(in_37bar),
    .I1(in_19bar)
  );
  //OR U481
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U481 (
    .O(n499),
    .I0(in_78),
    .I1(in_6)
  );
  //AND U481bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U481bar (
    .O(n499bar),
    .I0(in_78bar),
    .I1(in_6bar)
  );
  //OR U482
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U482 (
    .O(n603),
    .I0(n497),
    .I1(n496)
  );
  //AND U482bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U482bar (
    .O(n603bar),
    .I0(n497bar),
    .I1(n496bar)
  );
  //OR U483
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U483 (
    .O(n496),
    .I0(in[112]),
    .I1(in[102])
  );
  //AND U483bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U483bar (
    .O(n496bar),
    .I0(inbar[112]),
    .I1(inbar[102])
  );
  //OR U484
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U484 (
    .O(n497),
    .I0(in[123]),
    .I1(n495)
  );
  //AND U484bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U484bar (
    .O(n497bar),
    .I0(inbar[123]),
    .I1(n495bar)
  );
  //OR U485
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U485 (
    .O(n495),
    .I0(in[143]),
    .I1(in[130])
  );
  //AND U485bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U485bar (
    .O(n495bar),
    .I0(inbar[143]),
    .I1(inbar[130])
  );
  //OR U486
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U486 (
    .O(n605),
    .I0(n494),
    .I1(n493)
  );
  //AND U486bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U486bar (
    .O(n605bar),
    .I0(n494bar),
    .I1(n493bar)
  );
  //OR U487
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U487 (
    .O(n493),
    .I0(n492),
    .I1(n491)
  );
  //AND U487bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U487bar (
    .O(n493bar),
    .I0(n492bar),
    .I1(n491bar)
  );
  //OR U488
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U488 (
    .O(n491),
    .I0(in[216]),
    .I1(in[213])
  );
  //AND U488bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U488bar (
    .O(n491bar),
    .I0(inbar[216]),
    .I1(inbar[213])
  );
  //OR U489
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U489 (
    .O(n492),
    .I0(in[227]),
    .I1(n490)
  );
  //AND U489bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U489bar (
    .O(n492bar),
    .I0(inbar[227]),
    .I1(n490bar)
  );
  //OR U490
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U490 (
    .O(n490),
    .I0(in_0),
    .I1(in[248])
  );
  //AND U490bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U490bar (
    .O(n490bar),
    .I0(in_0bar),
    .I1(inbar[248])
  );
  //OR U491
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U491 (
    .O(n494),
    .I0(n489),
    .I1(n488)
  );
  //AND U491bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U491bar (
    .O(n494bar),
    .I0(n489bar),
    .I1(n488bar)
  );
  //OR U492
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U492 (
    .O(n488),
    .I0(in_46),
    .I1(in_44)
  );
  //AND U492bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U492bar (
    .O(n488bar),
    .I0(in_46bar),
    .I1(in_44bar)
  );
  //OR U493
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U493 (
    .O(n489),
    .I0(in_50),
    .I1(n487)
  );
  //AND U493bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U493bar (
    .O(n489bar),
    .I0(in_50bar),
    .I1(n487bar)
  );
  //OR U494
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U494 (
    .O(n487),
    .I0(in_9),
    .I1(in_80)
  );
  //AND U494bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U494bar (
    .O(n487bar),
    .I0(in_9bar),
    .I1(in_80bar)
  );
endmodule

module sBox_9 ( in, out );

  input wire [7:0] in;
//input_done

  output wire [7:0] out;
//output_done

  wire [255:0] decodeOut;
//wire_done

  decode_9 dec ( .in(in), .out(decodeOut) );
  encode_9 enc ( .in(decodeOut), .out(out) );
endmodule

module CD2_37 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD2_38 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD2_39 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD2_40 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD4_19 ( a, b, y );

  input wire [3:0] a;
  input wire [3:0] b;
  wire [3:0] abar;
  wire [3:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
//input_done

  output wire [15:0] y;
  wire [15:0] ybar;
//output_done

//wire_done

  //AND U1
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1 (
    .O(y[9]),
    .I0(b[1]),
    .I1(a[2])
  );
  //OR U1bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1bar (
    .O(ybar[9]),
    .I0(bbar[1]),
    .I1(abar[2])
  );
  //AND U2
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2 (
    .O(y[8]),
    .I0(b[0]),
    .I1(a[2])
  );
  //OR U2bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2bar (
    .O(ybar[8]),
    .I0(bbar[0]),
    .I1(abar[2])
  );
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[7]),
    .I0(b[3]),
    .I1(a[1])
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[7]),
    .I0(bbar[3]),
    .I1(abar[1])
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[6]),
    .I0(b[2]),
    .I1(a[1])
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[6]),
    .I0(bbar[2]),
    .I1(abar[1])
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[5]),
    .I0(a[1]),
    .I1(b[1])
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[5]),
    .I0(abar[1]),
    .I1(bbar[1])
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[4]),
    .I0(a[1]),
    .I1(b[0])
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[4]),
    .I0(abar[1]),
    .I1(bbar[0])
  );
  //AND U7
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7 (
    .O(y[3]),
    .I0(a[0]),
    .I1(b[3])
  );
  //OR U7bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7bar (
    .O(ybar[3]),
    .I0(abar[0]),
    .I1(bbar[3])
  );
  //AND U8
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8 (
    .O(y[2]),
    .I0(a[0]),
    .I1(b[2])
  );
  //OR U8bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8bar (
    .O(ybar[2]),
    .I0(abar[0]),
    .I1(bbar[2])
  );
  //AND U9
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9 (
    .O(y[1]),
    .I0(a[0]),
    .I1(b[1])
  );
  //OR U9bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9bar (
    .O(ybar[1]),
    .I0(abar[0]),
    .I1(bbar[1])
  );
  //AND U10
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10 (
    .O(y[15]),
    .I0(a[3]),
    .I1(b[3])
  );
  //OR U10bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10bar (
    .O(ybar[15]),
    .I0(abar[3]),
    .I1(bbar[3])
  );
  //AND U11
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11 (
    .O(y[14]),
    .I0(a[3]),
    .I1(b[2])
  );
  //OR U11bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11bar (
    .O(ybar[14]),
    .I0(abar[3]),
    .I1(bbar[2])
  );
  //AND U12
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12 (
    .O(y[13]),
    .I0(a[3]),
    .I1(b[1])
  );
  //OR U12bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12bar (
    .O(ybar[13]),
    .I0(abar[3]),
    .I1(bbar[1])
  );
  //AND U13
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13 (
    .O(y[12]),
    .I0(a[3]),
    .I1(b[0])
  );
  //OR U13bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13bar (
    .O(ybar[12]),
    .I0(abar[3]),
    .I1(bbar[0])
  );
  //AND U14
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14 (
    .O(y[11]),
    .I0(b[3]),
    .I1(a[2])
  );
  //OR U14bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14bar (
    .O(ybar[11]),
    .I0(bbar[3]),
    .I1(abar[2])
  );
  //AND U15
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15 (
    .O(y[10]),
    .I0(b[2]),
    .I1(a[2])
  );
  //OR U15bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15bar (
    .O(ybar[10]),
    .I0(bbar[2]),
    .I1(abar[2])
  );
  //AND U16
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16 (
    .O(y[0]),
    .I0(a[0]),
    .I1(b[0])
  );
  //OR U16bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16bar (
    .O(ybar[0]),
    .I0(abar[0]),
    .I1(bbar[0])
  );
endmodule

module CD4_20 ( a, b, y );

  input wire [3:0] a;
  input wire [3:0] b;
  wire [3:0] abar;
  wire [3:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
//input_done

  output wire [15:0] y;
  wire [15:0] ybar;
//output_done

//wire_done

  //AND U1
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1 (
    .O(y[9]),
    .I0(b[1]),
    .I1(a[2])
  );
  //OR U1bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1bar (
    .O(ybar[9]),
    .I0(bbar[1]),
    .I1(abar[2])
  );
  //AND U2
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2 (
    .O(y[8]),
    .I0(b[0]),
    .I1(a[2])
  );
  //OR U2bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2bar (
    .O(ybar[8]),
    .I0(bbar[0]),
    .I1(abar[2])
  );
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[7]),
    .I0(b[3]),
    .I1(a[1])
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[7]),
    .I0(bbar[3]),
    .I1(abar[1])
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[6]),
    .I0(b[2]),
    .I1(a[1])
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[6]),
    .I0(bbar[2]),
    .I1(abar[1])
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[5]),
    .I0(a[1]),
    .I1(b[1])
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[5]),
    .I0(abar[1]),
    .I1(bbar[1])
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[4]),
    .I0(a[1]),
    .I1(b[0])
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[4]),
    .I0(abar[1]),
    .I1(bbar[0])
  );
  //AND U7
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7 (
    .O(y[3]),
    .I0(a[0]),
    .I1(b[3])
  );
  //OR U7bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7bar (
    .O(ybar[3]),
    .I0(abar[0]),
    .I1(bbar[3])
  );
  //AND U8
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8 (
    .O(y[2]),
    .I0(a[0]),
    .I1(b[2])
  );
  //OR U8bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8bar (
    .O(ybar[2]),
    .I0(abar[0]),
    .I1(bbar[2])
  );
  //AND U9
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9 (
    .O(y[1]),
    .I0(a[0]),
    .I1(b[1])
  );
  //OR U9bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9bar (
    .O(ybar[1]),
    .I0(abar[0]),
    .I1(bbar[1])
  );
  //AND U10
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10 (
    .O(y[15]),
    .I0(a[3]),
    .I1(b[3])
  );
  //OR U10bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10bar (
    .O(ybar[15]),
    .I0(abar[3]),
    .I1(bbar[3])
  );
  //AND U11
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11 (
    .O(y[14]),
    .I0(a[3]),
    .I1(b[2])
  );
  //OR U11bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11bar (
    .O(ybar[14]),
    .I0(abar[3]),
    .I1(bbar[2])
  );
  //AND U12
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12 (
    .O(y[13]),
    .I0(a[3]),
    .I1(b[1])
  );
  //OR U12bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12bar (
    .O(ybar[13]),
    .I0(abar[3]),
    .I1(bbar[1])
  );
  //AND U13
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13 (
    .O(y[12]),
    .I0(a[3]),
    .I1(b[0])
  );
  //OR U13bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13bar (
    .O(ybar[12]),
    .I0(abar[3]),
    .I1(bbar[0])
  );
  //AND U14
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14 (
    .O(y[11]),
    .I0(b[3]),
    .I1(a[2])
  );
  //OR U14bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14bar (
    .O(ybar[11]),
    .I0(bbar[3]),
    .I1(abar[2])
  );
  //AND U15
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15 (
    .O(y[10]),
    .I0(b[2]),
    .I1(a[2])
  );
  //OR U15bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15bar (
    .O(ybar[10]),
    .I0(bbar[2]),
    .I1(abar[2])
  );
  //AND U16
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16 (
    .O(y[0]),
    .I0(a[0]),
    .I1(b[0])
  );
  //OR U16bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16bar (
    .O(ybar[0]),
    .I0(abar[0]),
    .I1(bbar[0])
  );
endmodule

module CD16_10 ( a, b, y );

  input wire [15:0] a;
  input wire [15:0] b;
  wire [15:0] abar;
  wire [15:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign abar[8] = ~a[8];
  assign abar[9] = ~a[9];
  assign abar[10] = ~a[10];
  assign abar[11] = ~a[11];
  assign abar[12] = ~a[12];
  assign abar[13] = ~a[13];
  assign abar[14] = ~a[14];
  assign abar[15] = ~a[15];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign bbar[8] = ~b[8];
  assign bbar[9] = ~b[9];
  assign bbar[10] = ~b[10];
  assign bbar[11] = ~b[11];
  assign bbar[12] = ~b[12];
  assign bbar[13] = ~b[13];
  assign bbar[14] = ~b[14];
  assign bbar[15] = ~b[15];
//input_done

  output wire [255:0] y;
  wire [255:0] ybar;
//output_done

//wire_done

  //AND U1
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1 (
    .O(y[9]),
    .I0(b[9]),
    .I1(a[0])
  );
  //OR U1bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1bar (
    .O(ybar[9]),
    .I0(bbar[9]),
    .I1(abar[0])
  );
  //AND U2
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2 (
    .O(y[99]),
    .I0(b[3]),
    .I1(a[6])
  );
  //OR U2bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2bar (
    .O(ybar[99]),
    .I0(bbar[3]),
    .I1(abar[6])
  );
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[98]),
    .I0(b[2]),
    .I1(a[6])
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[98]),
    .I0(bbar[2]),
    .I1(abar[6])
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[97]),
    .I0(b[1]),
    .I1(a[6])
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[97]),
    .I0(bbar[1]),
    .I1(abar[6])
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[96]),
    .I0(b[0]),
    .I1(a[6])
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[96]),
    .I0(bbar[0]),
    .I1(abar[6])
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[95]),
    .I0(b[15]),
    .I1(a[5])
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[95]),
    .I0(bbar[15]),
    .I1(abar[5])
  );
  //AND U7
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7 (
    .O(y[94]),
    .I0(b[14]),
    .I1(a[5])
  );
  //OR U7bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7bar (
    .O(ybar[94]),
    .I0(bbar[14]),
    .I1(abar[5])
  );
  //AND U8
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8 (
    .O(y[93]),
    .I0(b[13]),
    .I1(a[5])
  );
  //OR U8bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8bar (
    .O(ybar[93]),
    .I0(bbar[13]),
    .I1(abar[5])
  );
  //AND U9
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9 (
    .O(y[92]),
    .I0(b[12]),
    .I1(a[5])
  );
  //OR U9bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9bar (
    .O(ybar[92]),
    .I0(bbar[12]),
    .I1(abar[5])
  );
  //AND U10
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10 (
    .O(y[91]),
    .I0(b[11]),
    .I1(a[5])
  );
  //OR U10bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10bar (
    .O(ybar[91]),
    .I0(bbar[11]),
    .I1(abar[5])
  );
  //AND U11
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11 (
    .O(y[90]),
    .I0(b[10]),
    .I1(a[5])
  );
  //OR U11bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11bar (
    .O(ybar[90]),
    .I0(bbar[10]),
    .I1(abar[5])
  );
  //AND U12
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12 (
    .O(y[8]),
    .I0(b[8]),
    .I1(a[0])
  );
  //OR U12bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12bar (
    .O(ybar[8]),
    .I0(bbar[8]),
    .I1(abar[0])
  );
  //AND U13
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13 (
    .O(y[89]),
    .I0(a[5]),
    .I1(b[9])
  );
  //OR U13bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13bar (
    .O(ybar[89]),
    .I0(abar[5]),
    .I1(bbar[9])
  );
  //AND U14
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14 (
    .O(y[88]),
    .I0(b[8]),
    .I1(a[5])
  );
  //OR U14bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14bar (
    .O(ybar[88]),
    .I0(bbar[8]),
    .I1(abar[5])
  );
  //AND U15
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15 (
    .O(y[87]),
    .I0(b[7]),
    .I1(a[5])
  );
  //OR U15bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15bar (
    .O(ybar[87]),
    .I0(bbar[7]),
    .I1(abar[5])
  );
  //AND U16
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16 (
    .O(y[86]),
    .I0(b[6]),
    .I1(a[5])
  );
  //OR U16bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16bar (
    .O(ybar[86]),
    .I0(bbar[6]),
    .I1(abar[5])
  );
  //AND U17
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U17 (
    .O(y[85]),
    .I0(b[5]),
    .I1(a[5])
  );
  //OR U17bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U17bar (
    .O(ybar[85]),
    .I0(bbar[5]),
    .I1(abar[5])
  );
  //AND U18
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U18 (
    .O(y[84]),
    .I0(b[4]),
    .I1(a[5])
  );
  //OR U18bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U18bar (
    .O(ybar[84]),
    .I0(bbar[4]),
    .I1(abar[5])
  );
  //AND U19
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U19 (
    .O(y[83]),
    .I0(a[5]),
    .I1(b[3])
  );
  //OR U19bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U19bar (
    .O(ybar[83]),
    .I0(abar[5]),
    .I1(bbar[3])
  );
  //AND U20
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U20 (
    .O(y[82]),
    .I0(a[5]),
    .I1(b[2])
  );
  //OR U20bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U20bar (
    .O(ybar[82]),
    .I0(abar[5]),
    .I1(bbar[2])
  );
  //AND U21
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U21 (
    .O(y[81]),
    .I0(a[5]),
    .I1(b[1])
  );
  //OR U21bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U21bar (
    .O(ybar[81]),
    .I0(abar[5]),
    .I1(bbar[1])
  );
  //AND U22
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U22 (
    .O(y[80]),
    .I0(a[5]),
    .I1(b[0])
  );
  //OR U22bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U22bar (
    .O(ybar[80]),
    .I0(abar[5]),
    .I1(bbar[0])
  );
  //AND U23
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U23 (
    .O(y[7]),
    .I0(b[7]),
    .I1(a[0])
  );
  //OR U23bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U23bar (
    .O(ybar[7]),
    .I0(bbar[7]),
    .I1(abar[0])
  );
  //AND U24
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U24 (
    .O(y[79]),
    .I0(a[4]),
    .I1(b[15])
  );
  //OR U24bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U24bar (
    .O(ybar[79]),
    .I0(abar[4]),
    .I1(bbar[15])
  );
  //AND U25
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U25 (
    .O(y[78]),
    .I0(a[4]),
    .I1(b[14])
  );
  //OR U25bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U25bar (
    .O(ybar[78]),
    .I0(abar[4]),
    .I1(bbar[14])
  );
  //AND U26
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U26 (
    .O(y[77]),
    .I0(a[4]),
    .I1(b[13])
  );
  //OR U26bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U26bar (
    .O(ybar[77]),
    .I0(abar[4]),
    .I1(bbar[13])
  );
  //AND U27
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U27 (
    .O(y[76]),
    .I0(a[4]),
    .I1(b[12])
  );
  //OR U27bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U27bar (
    .O(ybar[76]),
    .I0(abar[4]),
    .I1(bbar[12])
  );
  //AND U28
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U28 (
    .O(y[75]),
    .I0(a[4]),
    .I1(b[11])
  );
  //OR U28bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U28bar (
    .O(ybar[75]),
    .I0(abar[4]),
    .I1(bbar[11])
  );
  //AND U29
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U29 (
    .O(y[74]),
    .I0(a[4]),
    .I1(b[10])
  );
  //OR U29bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U29bar (
    .O(ybar[74]),
    .I0(abar[4]),
    .I1(bbar[10])
  );
  //AND U30
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U30 (
    .O(y[73]),
    .I0(a[4]),
    .I1(b[9])
  );
  //OR U30bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U30bar (
    .O(ybar[73]),
    .I0(abar[4]),
    .I1(bbar[9])
  );
  //AND U31
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U31 (
    .O(y[72]),
    .I0(a[4]),
    .I1(b[8])
  );
  //OR U31bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U31bar (
    .O(ybar[72]),
    .I0(abar[4]),
    .I1(bbar[8])
  );
  //AND U32
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U32 (
    .O(y[71]),
    .I0(a[4]),
    .I1(b[7])
  );
  //OR U32bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U32bar (
    .O(ybar[71]),
    .I0(abar[4]),
    .I1(bbar[7])
  );
  //AND U33
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U33 (
    .O(y[70]),
    .I0(a[4]),
    .I1(b[6])
  );
  //OR U33bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U33bar (
    .O(ybar[70]),
    .I0(abar[4]),
    .I1(bbar[6])
  );
  //AND U34
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U34 (
    .O(y[6]),
    .I0(b[6]),
    .I1(a[0])
  );
  //OR U34bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U34bar (
    .O(ybar[6]),
    .I0(bbar[6]),
    .I1(abar[0])
  );
  //AND U35
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U35 (
    .O(y[69]),
    .I0(a[4]),
    .I1(b[5])
  );
  //OR U35bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U35bar (
    .O(ybar[69]),
    .I0(abar[4]),
    .I1(bbar[5])
  );
  //AND U36
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U36 (
    .O(y[68]),
    .I0(a[4]),
    .I1(b[4])
  );
  //OR U36bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U36bar (
    .O(ybar[68]),
    .I0(abar[4]),
    .I1(bbar[4])
  );
  //AND U37
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U37 (
    .O(y[67]),
    .I0(a[4]),
    .I1(b[3])
  );
  //OR U37bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U37bar (
    .O(ybar[67]),
    .I0(abar[4]),
    .I1(bbar[3])
  );
  //AND U38
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U38 (
    .O(y[66]),
    .I0(a[4]),
    .I1(b[2])
  );
  //OR U38bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U38bar (
    .O(ybar[66]),
    .I0(abar[4]),
    .I1(bbar[2])
  );
  //AND U39
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U39 (
    .O(y[65]),
    .I0(a[4]),
    .I1(b[1])
  );
  //OR U39bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U39bar (
    .O(ybar[65]),
    .I0(abar[4]),
    .I1(bbar[1])
  );
  //AND U40
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U40 (
    .O(y[64]),
    .I0(a[4]),
    .I1(b[0])
  );
  //OR U40bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U40bar (
    .O(ybar[64]),
    .I0(abar[4]),
    .I1(bbar[0])
  );
  //AND U41
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U41 (
    .O(y[63]),
    .I0(a[3]),
    .I1(b[15])
  );
  //OR U41bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U41bar (
    .O(ybar[63]),
    .I0(abar[3]),
    .I1(bbar[15])
  );
  //AND U42
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U42 (
    .O(y[62]),
    .I0(a[3]),
    .I1(b[14])
  );
  //OR U42bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U42bar (
    .O(ybar[62]),
    .I0(abar[3]),
    .I1(bbar[14])
  );
  //AND U43
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U43 (
    .O(y[61]),
    .I0(a[3]),
    .I1(b[13])
  );
  //OR U43bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U43bar (
    .O(ybar[61]),
    .I0(abar[3]),
    .I1(bbar[13])
  );
  //AND U44
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U44 (
    .O(y[60]),
    .I0(a[3]),
    .I1(b[12])
  );
  //OR U44bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U44bar (
    .O(ybar[60]),
    .I0(abar[3]),
    .I1(bbar[12])
  );
  //AND U45
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U45 (
    .O(y[5]),
    .I0(b[5]),
    .I1(a[0])
  );
  //OR U45bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U45bar (
    .O(ybar[5]),
    .I0(bbar[5]),
    .I1(abar[0])
  );
  //AND U46
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U46 (
    .O(y[59]),
    .I0(a[3]),
    .I1(b[11])
  );
  //OR U46bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U46bar (
    .O(ybar[59]),
    .I0(abar[3]),
    .I1(bbar[11])
  );
  //AND U47
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U47 (
    .O(y[58]),
    .I0(a[3]),
    .I1(b[10])
  );
  //OR U47bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U47bar (
    .O(ybar[58]),
    .I0(abar[3]),
    .I1(bbar[10])
  );
  //AND U48
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U48 (
    .O(y[57]),
    .I0(a[3]),
    .I1(b[9])
  );
  //OR U48bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U48bar (
    .O(ybar[57]),
    .I0(abar[3]),
    .I1(bbar[9])
  );
  //AND U49
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U49 (
    .O(y[56]),
    .I0(a[3]),
    .I1(b[8])
  );
  //OR U49bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U49bar (
    .O(ybar[56]),
    .I0(abar[3]),
    .I1(bbar[8])
  );
  //AND U50
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U50 (
    .O(y[55]),
    .I0(a[3]),
    .I1(b[7])
  );
  //OR U50bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U50bar (
    .O(ybar[55]),
    .I0(abar[3]),
    .I1(bbar[7])
  );
  //AND U51
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U51 (
    .O(y[54]),
    .I0(a[3]),
    .I1(b[6])
  );
  //OR U51bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U51bar (
    .O(ybar[54]),
    .I0(abar[3]),
    .I1(bbar[6])
  );
  //AND U52
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U52 (
    .O(y[53]),
    .I0(a[3]),
    .I1(b[5])
  );
  //OR U52bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U52bar (
    .O(ybar[53]),
    .I0(abar[3]),
    .I1(bbar[5])
  );
  //AND U53
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U53 (
    .O(y[52]),
    .I0(a[3]),
    .I1(b[4])
  );
  //OR U53bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U53bar (
    .O(ybar[52]),
    .I0(abar[3]),
    .I1(bbar[4])
  );
  //AND U54
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U54 (
    .O(y[51]),
    .I0(a[3]),
    .I1(b[3])
  );
  //OR U54bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U54bar (
    .O(ybar[51]),
    .I0(abar[3]),
    .I1(bbar[3])
  );
  //AND U55
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U55 (
    .O(y[50]),
    .I0(a[3]),
    .I1(b[2])
  );
  //OR U55bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U55bar (
    .O(ybar[50]),
    .I0(abar[3]),
    .I1(bbar[2])
  );
  //AND U56
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U56 (
    .O(y[4]),
    .I0(b[4]),
    .I1(a[0])
  );
  //OR U56bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U56bar (
    .O(ybar[4]),
    .I0(bbar[4]),
    .I1(abar[0])
  );
  //AND U57
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U57 (
    .O(y[49]),
    .I0(a[3]),
    .I1(b[1])
  );
  //OR U57bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U57bar (
    .O(ybar[49]),
    .I0(abar[3]),
    .I1(bbar[1])
  );
  //AND U58
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U58 (
    .O(y[48]),
    .I0(a[3]),
    .I1(b[0])
  );
  //OR U58bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U58bar (
    .O(ybar[48]),
    .I0(abar[3]),
    .I1(bbar[0])
  );
  //AND U59
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U59 (
    .O(y[47]),
    .I0(a[2]),
    .I1(b[15])
  );
  //OR U59bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U59bar (
    .O(ybar[47]),
    .I0(abar[2]),
    .I1(bbar[15])
  );
  //AND U60
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U60 (
    .O(y[46]),
    .I0(a[2]),
    .I1(b[14])
  );
  //OR U60bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U60bar (
    .O(ybar[46]),
    .I0(abar[2]),
    .I1(bbar[14])
  );
  //AND U61
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U61 (
    .O(y[45]),
    .I0(a[2]),
    .I1(b[13])
  );
  //OR U61bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U61bar (
    .O(ybar[45]),
    .I0(abar[2]),
    .I1(bbar[13])
  );
  //AND U62
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U62 (
    .O(y[44]),
    .I0(a[2]),
    .I1(b[12])
  );
  //OR U62bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U62bar (
    .O(ybar[44]),
    .I0(abar[2]),
    .I1(bbar[12])
  );
  //AND U63
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U63 (
    .O(y[43]),
    .I0(a[2]),
    .I1(b[11])
  );
  //OR U63bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U63bar (
    .O(ybar[43]),
    .I0(abar[2]),
    .I1(bbar[11])
  );
  //AND U64
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U64 (
    .O(y[42]),
    .I0(a[2]),
    .I1(b[10])
  );
  //OR U64bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U64bar (
    .O(ybar[42]),
    .I0(abar[2]),
    .I1(bbar[10])
  );
  //AND U65
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U65 (
    .O(y[41]),
    .I0(a[2]),
    .I1(b[9])
  );
  //OR U65bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U65bar (
    .O(ybar[41]),
    .I0(abar[2]),
    .I1(bbar[9])
  );
  //AND U66
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U66 (
    .O(y[40]),
    .I0(a[2]),
    .I1(b[8])
  );
  //OR U66bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U66bar (
    .O(ybar[40]),
    .I0(abar[2]),
    .I1(bbar[8])
  );
  //AND U67
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U67 (
    .O(y[3]),
    .I0(b[3]),
    .I1(a[0])
  );
  //OR U67bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U67bar (
    .O(ybar[3]),
    .I0(bbar[3]),
    .I1(abar[0])
  );
  //AND U68
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U68 (
    .O(y[39]),
    .I0(a[2]),
    .I1(b[7])
  );
  //OR U68bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U68bar (
    .O(ybar[39]),
    .I0(abar[2]),
    .I1(bbar[7])
  );
  //AND U69
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U69 (
    .O(y[38]),
    .I0(a[2]),
    .I1(b[6])
  );
  //OR U69bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U69bar (
    .O(ybar[38]),
    .I0(abar[2]),
    .I1(bbar[6])
  );
  //AND U70
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U70 (
    .O(y[37]),
    .I0(a[2]),
    .I1(b[5])
  );
  //OR U70bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U70bar (
    .O(ybar[37]),
    .I0(abar[2]),
    .I1(bbar[5])
  );
  //AND U71
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U71 (
    .O(y[36]),
    .I0(a[2]),
    .I1(b[4])
  );
  //OR U71bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U71bar (
    .O(ybar[36]),
    .I0(abar[2]),
    .I1(bbar[4])
  );
  //AND U72
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U72 (
    .O(y[35]),
    .I0(a[2]),
    .I1(b[3])
  );
  //OR U72bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U72bar (
    .O(ybar[35]),
    .I0(abar[2]),
    .I1(bbar[3])
  );
  //AND U73
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U73 (
    .O(y[34]),
    .I0(a[2]),
    .I1(b[2])
  );
  //OR U73bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U73bar (
    .O(ybar[34]),
    .I0(abar[2]),
    .I1(bbar[2])
  );
  //AND U74
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U74 (
    .O(y[33]),
    .I0(a[2]),
    .I1(b[1])
  );
  //OR U74bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U74bar (
    .O(ybar[33]),
    .I0(abar[2]),
    .I1(bbar[1])
  );
  //AND U75
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U75 (
    .O(y[32]),
    .I0(a[2]),
    .I1(b[0])
  );
  //OR U75bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U75bar (
    .O(ybar[32]),
    .I0(abar[2]),
    .I1(bbar[0])
  );
  //AND U76
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U76 (
    .O(y[31]),
    .I0(a[1]),
    .I1(b[15])
  );
  //OR U76bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U76bar (
    .O(ybar[31]),
    .I0(abar[1]),
    .I1(bbar[15])
  );
  //AND U77
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U77 (
    .O(y[30]),
    .I0(a[1]),
    .I1(b[14])
  );
  //OR U77bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U77bar (
    .O(ybar[30]),
    .I0(abar[1]),
    .I1(bbar[14])
  );
  //AND U78
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U78 (
    .O(y[2]),
    .I0(b[2]),
    .I1(a[0])
  );
  //OR U78bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U78bar (
    .O(ybar[2]),
    .I0(bbar[2]),
    .I1(abar[0])
  );
  //AND U79
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U79 (
    .O(y[29]),
    .I0(a[1]),
    .I1(b[13])
  );
  //OR U79bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U79bar (
    .O(ybar[29]),
    .I0(abar[1]),
    .I1(bbar[13])
  );
  //AND U80
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U80 (
    .O(y[28]),
    .I0(a[1]),
    .I1(b[12])
  );
  //OR U80bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U80bar (
    .O(ybar[28]),
    .I0(abar[1]),
    .I1(bbar[12])
  );
  //AND U81
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U81 (
    .O(y[27]),
    .I0(a[1]),
    .I1(b[11])
  );
  //OR U81bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U81bar (
    .O(ybar[27]),
    .I0(abar[1]),
    .I1(bbar[11])
  );
  //AND U82
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U82 (
    .O(y[26]),
    .I0(a[1]),
    .I1(b[10])
  );
  //OR U82bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U82bar (
    .O(ybar[26]),
    .I0(abar[1]),
    .I1(bbar[10])
  );
  //AND U83
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U83 (
    .O(y[25]),
    .I0(a[1]),
    .I1(b[9])
  );
  //OR U83bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U83bar (
    .O(ybar[25]),
    .I0(abar[1]),
    .I1(bbar[9])
  );
  //AND U84
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U84 (
    .O(y[255]),
    .I0(a[15]),
    .I1(b[15])
  );
  //OR U84bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U84bar (
    .O(ybar[255]),
    .I0(abar[15]),
    .I1(bbar[15])
  );
  //AND U85
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U85 (
    .O(y[254]),
    .I0(a[15]),
    .I1(b[14])
  );
  //OR U85bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U85bar (
    .O(ybar[254]),
    .I0(abar[15]),
    .I1(bbar[14])
  );
  //AND U86
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U86 (
    .O(y[253]),
    .I0(a[15]),
    .I1(b[13])
  );
  //OR U86bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U86bar (
    .O(ybar[253]),
    .I0(abar[15]),
    .I1(bbar[13])
  );
  //AND U87
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U87 (
    .O(y[252]),
    .I0(a[15]),
    .I1(b[12])
  );
  //OR U87bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U87bar (
    .O(ybar[252]),
    .I0(abar[15]),
    .I1(bbar[12])
  );
  //AND U88
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U88 (
    .O(y[251]),
    .I0(a[15]),
    .I1(b[11])
  );
  //OR U88bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U88bar (
    .O(ybar[251]),
    .I0(abar[15]),
    .I1(bbar[11])
  );
  //AND U89
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U89 (
    .O(y[250]),
    .I0(a[15]),
    .I1(b[10])
  );
  //OR U89bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U89bar (
    .O(ybar[250]),
    .I0(abar[15]),
    .I1(bbar[10])
  );
  //AND U90
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U90 (
    .O(y[24]),
    .I0(a[1]),
    .I1(b[8])
  );
  //OR U90bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U90bar (
    .O(ybar[24]),
    .I0(abar[1]),
    .I1(bbar[8])
  );
  //AND U91
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U91 (
    .O(y[249]),
    .I0(a[15]),
    .I1(b[9])
  );
  //OR U91bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U91bar (
    .O(ybar[249]),
    .I0(abar[15]),
    .I1(bbar[9])
  );
  //AND U92
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U92 (
    .O(y[248]),
    .I0(a[15]),
    .I1(b[8])
  );
  //OR U92bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U92bar (
    .O(ybar[248]),
    .I0(abar[15]),
    .I1(bbar[8])
  );
  //AND U93
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U93 (
    .O(y[247]),
    .I0(a[15]),
    .I1(b[7])
  );
  //OR U93bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U93bar (
    .O(ybar[247]),
    .I0(abar[15]),
    .I1(bbar[7])
  );
  //AND U94
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U94 (
    .O(y[246]),
    .I0(a[15]),
    .I1(b[6])
  );
  //OR U94bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U94bar (
    .O(ybar[246]),
    .I0(abar[15]),
    .I1(bbar[6])
  );
  //AND U95
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U95 (
    .O(y[245]),
    .I0(a[15]),
    .I1(b[5])
  );
  //OR U95bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U95bar (
    .O(ybar[245]),
    .I0(abar[15]),
    .I1(bbar[5])
  );
  //AND U96
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U96 (
    .O(y[244]),
    .I0(a[15]),
    .I1(b[4])
  );
  //OR U96bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U96bar (
    .O(ybar[244]),
    .I0(abar[15]),
    .I1(bbar[4])
  );
  //AND U97
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U97 (
    .O(y[243]),
    .I0(a[15]),
    .I1(b[3])
  );
  //OR U97bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U97bar (
    .O(ybar[243]),
    .I0(abar[15]),
    .I1(bbar[3])
  );
  //AND U98
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U98 (
    .O(y[242]),
    .I0(a[15]),
    .I1(b[2])
  );
  //OR U98bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U98bar (
    .O(ybar[242]),
    .I0(abar[15]),
    .I1(bbar[2])
  );
  //AND U99
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U99 (
    .O(y[241]),
    .I0(a[15]),
    .I1(b[1])
  );
  //OR U99bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U99bar (
    .O(ybar[241]),
    .I0(abar[15]),
    .I1(bbar[1])
  );
  //AND U100
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U100 (
    .O(y[240]),
    .I0(a[15]),
    .I1(b[0])
  );
  //OR U100bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U100bar (
    .O(ybar[240]),
    .I0(abar[15]),
    .I1(bbar[0])
  );
  //AND U101
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U101 (
    .O(y[23]),
    .I0(a[1]),
    .I1(b[7])
  );
  //OR U101bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U101bar (
    .O(ybar[23]),
    .I0(abar[1]),
    .I1(bbar[7])
  );
  //AND U102
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U102 (
    .O(y[239]),
    .I0(a[14]),
    .I1(b[15])
  );
  //OR U102bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U102bar (
    .O(ybar[239]),
    .I0(abar[14]),
    .I1(bbar[15])
  );
  //AND U103
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U103 (
    .O(y[238]),
    .I0(a[14]),
    .I1(b[14])
  );
  //OR U103bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U103bar (
    .O(ybar[238]),
    .I0(abar[14]),
    .I1(bbar[14])
  );
  //AND U104
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U104 (
    .O(y[237]),
    .I0(a[14]),
    .I1(b[13])
  );
  //OR U104bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U104bar (
    .O(ybar[237]),
    .I0(abar[14]),
    .I1(bbar[13])
  );
  //AND U105
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U105 (
    .O(y[236]),
    .I0(a[14]),
    .I1(b[12])
  );
  //OR U105bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U105bar (
    .O(ybar[236]),
    .I0(abar[14]),
    .I1(bbar[12])
  );
  //AND U106
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U106 (
    .O(y[235]),
    .I0(a[14]),
    .I1(b[11])
  );
  //OR U106bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U106bar (
    .O(ybar[235]),
    .I0(abar[14]),
    .I1(bbar[11])
  );
  //AND U107
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U107 (
    .O(y[234]),
    .I0(a[14]),
    .I1(b[10])
  );
  //OR U107bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U107bar (
    .O(ybar[234]),
    .I0(abar[14]),
    .I1(bbar[10])
  );
  //AND U108
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U108 (
    .O(y[233]),
    .I0(a[14]),
    .I1(b[9])
  );
  //OR U108bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U108bar (
    .O(ybar[233]),
    .I0(abar[14]),
    .I1(bbar[9])
  );
  //AND U109
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U109 (
    .O(y[232]),
    .I0(a[14]),
    .I1(b[8])
  );
  //OR U109bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U109bar (
    .O(ybar[232]),
    .I0(abar[14]),
    .I1(bbar[8])
  );
  //AND U110
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U110 (
    .O(y[231]),
    .I0(a[14]),
    .I1(b[7])
  );
  //OR U110bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U110bar (
    .O(ybar[231]),
    .I0(abar[14]),
    .I1(bbar[7])
  );
  //AND U111
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U111 (
    .O(y[230]),
    .I0(a[14]),
    .I1(b[6])
  );
  //OR U111bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U111bar (
    .O(ybar[230]),
    .I0(abar[14]),
    .I1(bbar[6])
  );
  //AND U112
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U112 (
    .O(y[22]),
    .I0(a[1]),
    .I1(b[6])
  );
  //OR U112bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U112bar (
    .O(ybar[22]),
    .I0(abar[1]),
    .I1(bbar[6])
  );
  //AND U113
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U113 (
    .O(y[229]),
    .I0(a[14]),
    .I1(b[5])
  );
  //OR U113bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U113bar (
    .O(ybar[229]),
    .I0(abar[14]),
    .I1(bbar[5])
  );
  //AND U114
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U114 (
    .O(y[228]),
    .I0(a[14]),
    .I1(b[4])
  );
  //OR U114bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U114bar (
    .O(ybar[228]),
    .I0(abar[14]),
    .I1(bbar[4])
  );
  //AND U115
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U115 (
    .O(y[227]),
    .I0(a[14]),
    .I1(b[3])
  );
  //OR U115bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U115bar (
    .O(ybar[227]),
    .I0(abar[14]),
    .I1(bbar[3])
  );
  //AND U116
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U116 (
    .O(y[226]),
    .I0(a[14]),
    .I1(b[2])
  );
  //OR U116bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U116bar (
    .O(ybar[226]),
    .I0(abar[14]),
    .I1(bbar[2])
  );
  //AND U117
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U117 (
    .O(y[225]),
    .I0(a[14]),
    .I1(b[1])
  );
  //OR U117bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U117bar (
    .O(ybar[225]),
    .I0(abar[14]),
    .I1(bbar[1])
  );
  //AND U118
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U118 (
    .O(y[224]),
    .I0(a[14]),
    .I1(b[0])
  );
  //OR U118bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U118bar (
    .O(ybar[224]),
    .I0(abar[14]),
    .I1(bbar[0])
  );
  //AND U119
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U119 (
    .O(y[223]),
    .I0(a[13]),
    .I1(b[15])
  );
  //OR U119bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U119bar (
    .O(ybar[223]),
    .I0(abar[13]),
    .I1(bbar[15])
  );
  //AND U120
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U120 (
    .O(y[222]),
    .I0(a[13]),
    .I1(b[14])
  );
  //OR U120bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U120bar (
    .O(ybar[222]),
    .I0(abar[13]),
    .I1(bbar[14])
  );
  //AND U121
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U121 (
    .O(y[221]),
    .I0(a[13]),
    .I1(b[13])
  );
  //OR U121bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U121bar (
    .O(ybar[221]),
    .I0(abar[13]),
    .I1(bbar[13])
  );
  //AND U122
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U122 (
    .O(y[220]),
    .I0(a[13]),
    .I1(b[12])
  );
  //OR U122bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U122bar (
    .O(ybar[220]),
    .I0(abar[13]),
    .I1(bbar[12])
  );
  //AND U123
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U123 (
    .O(y[21]),
    .I0(a[1]),
    .I1(b[5])
  );
  //OR U123bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U123bar (
    .O(ybar[21]),
    .I0(abar[1]),
    .I1(bbar[5])
  );
  //AND U124
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U124 (
    .O(y[219]),
    .I0(a[13]),
    .I1(b[11])
  );
  //OR U124bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U124bar (
    .O(ybar[219]),
    .I0(abar[13]),
    .I1(bbar[11])
  );
  //AND U125
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U125 (
    .O(y[218]),
    .I0(a[13]),
    .I1(b[10])
  );
  //OR U125bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U125bar (
    .O(ybar[218]),
    .I0(abar[13]),
    .I1(bbar[10])
  );
  //AND U126
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U126 (
    .O(y[217]),
    .I0(a[13]),
    .I1(b[9])
  );
  //OR U126bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U126bar (
    .O(ybar[217]),
    .I0(abar[13]),
    .I1(bbar[9])
  );
  //AND U127
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U127 (
    .O(y[216]),
    .I0(a[13]),
    .I1(b[8])
  );
  //OR U127bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U127bar (
    .O(ybar[216]),
    .I0(abar[13]),
    .I1(bbar[8])
  );
  //AND U128
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U128 (
    .O(y[215]),
    .I0(a[13]),
    .I1(b[7])
  );
  //OR U128bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U128bar (
    .O(ybar[215]),
    .I0(abar[13]),
    .I1(bbar[7])
  );
  //AND U129
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U129 (
    .O(y[214]),
    .I0(a[13]),
    .I1(b[6])
  );
  //OR U129bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U129bar (
    .O(ybar[214]),
    .I0(abar[13]),
    .I1(bbar[6])
  );
  //AND U130
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U130 (
    .O(y[213]),
    .I0(a[13]),
    .I1(b[5])
  );
  //OR U130bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U130bar (
    .O(ybar[213]),
    .I0(abar[13]),
    .I1(bbar[5])
  );
  //AND U131
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U131 (
    .O(y[212]),
    .I0(a[13]),
    .I1(b[4])
  );
  //OR U131bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U131bar (
    .O(ybar[212]),
    .I0(abar[13]),
    .I1(bbar[4])
  );
  //AND U132
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U132 (
    .O(y[211]),
    .I0(a[13]),
    .I1(b[3])
  );
  //OR U132bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U132bar (
    .O(ybar[211]),
    .I0(abar[13]),
    .I1(bbar[3])
  );
  //AND U133
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U133 (
    .O(y[210]),
    .I0(a[13]),
    .I1(b[2])
  );
  //OR U133bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U133bar (
    .O(ybar[210]),
    .I0(abar[13]),
    .I1(bbar[2])
  );
  //AND U134
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U134 (
    .O(y[20]),
    .I0(a[1]),
    .I1(b[4])
  );
  //OR U134bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U134bar (
    .O(ybar[20]),
    .I0(abar[1]),
    .I1(bbar[4])
  );
  //AND U135
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U135 (
    .O(y[209]),
    .I0(a[13]),
    .I1(b[1])
  );
  //OR U135bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U135bar (
    .O(ybar[209]),
    .I0(abar[13]),
    .I1(bbar[1])
  );
  //AND U136
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U136 (
    .O(y[208]),
    .I0(a[13]),
    .I1(b[0])
  );
  //OR U136bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U136bar (
    .O(ybar[208]),
    .I0(abar[13]),
    .I1(bbar[0])
  );
  //AND U137
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U137 (
    .O(y[207]),
    .I0(a[12]),
    .I1(b[15])
  );
  //OR U137bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U137bar (
    .O(ybar[207]),
    .I0(abar[12]),
    .I1(bbar[15])
  );
  //AND U138
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U138 (
    .O(y[206]),
    .I0(a[12]),
    .I1(b[14])
  );
  //OR U138bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U138bar (
    .O(ybar[206]),
    .I0(abar[12]),
    .I1(bbar[14])
  );
  //AND U139
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U139 (
    .O(y[205]),
    .I0(a[12]),
    .I1(b[13])
  );
  //OR U139bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U139bar (
    .O(ybar[205]),
    .I0(abar[12]),
    .I1(bbar[13])
  );
  //AND U140
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U140 (
    .O(y[204]),
    .I0(a[12]),
    .I1(b[12])
  );
  //OR U140bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U140bar (
    .O(ybar[204]),
    .I0(abar[12]),
    .I1(bbar[12])
  );
  //AND U141
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U141 (
    .O(y[203]),
    .I0(a[12]),
    .I1(b[11])
  );
  //OR U141bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U141bar (
    .O(ybar[203]),
    .I0(abar[12]),
    .I1(bbar[11])
  );
  //AND U142
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U142 (
    .O(y[202]),
    .I0(a[12]),
    .I1(b[10])
  );
  //OR U142bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U142bar (
    .O(ybar[202]),
    .I0(abar[12]),
    .I1(bbar[10])
  );
  //AND U143
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U143 (
    .O(y[201]),
    .I0(a[12]),
    .I1(b[9])
  );
  //OR U143bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U143bar (
    .O(ybar[201]),
    .I0(abar[12]),
    .I1(bbar[9])
  );
  //AND U144
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U144 (
    .O(y[200]),
    .I0(a[12]),
    .I1(b[8])
  );
  //OR U144bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U144bar (
    .O(ybar[200]),
    .I0(abar[12]),
    .I1(bbar[8])
  );
  //AND U145
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U145 (
    .O(y[1]),
    .I0(b[1]),
    .I1(a[0])
  );
  //OR U145bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U145bar (
    .O(ybar[1]),
    .I0(bbar[1]),
    .I1(abar[0])
  );
  //AND U146
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U146 (
    .O(y[19]),
    .I0(a[1]),
    .I1(b[3])
  );
  //OR U146bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U146bar (
    .O(ybar[19]),
    .I0(abar[1]),
    .I1(bbar[3])
  );
  //AND U147
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U147 (
    .O(y[199]),
    .I0(a[12]),
    .I1(b[7])
  );
  //OR U147bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U147bar (
    .O(ybar[199]),
    .I0(abar[12]),
    .I1(bbar[7])
  );
  //AND U148
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U148 (
    .O(y[198]),
    .I0(a[12]),
    .I1(b[6])
  );
  //OR U148bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U148bar (
    .O(ybar[198]),
    .I0(abar[12]),
    .I1(bbar[6])
  );
  //AND U149
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U149 (
    .O(y[197]),
    .I0(a[12]),
    .I1(b[5])
  );
  //OR U149bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U149bar (
    .O(ybar[197]),
    .I0(abar[12]),
    .I1(bbar[5])
  );
  //AND U150
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U150 (
    .O(y[196]),
    .I0(a[12]),
    .I1(b[4])
  );
  //OR U150bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U150bar (
    .O(ybar[196]),
    .I0(abar[12]),
    .I1(bbar[4])
  );
  //AND U151
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U151 (
    .O(y[195]),
    .I0(a[12]),
    .I1(b[3])
  );
  //OR U151bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U151bar (
    .O(ybar[195]),
    .I0(abar[12]),
    .I1(bbar[3])
  );
  //AND U152
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U152 (
    .O(y[194]),
    .I0(a[12]),
    .I1(b[2])
  );
  //OR U152bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U152bar (
    .O(ybar[194]),
    .I0(abar[12]),
    .I1(bbar[2])
  );
  //AND U153
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U153 (
    .O(y[193]),
    .I0(a[12]),
    .I1(b[1])
  );
  //OR U153bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U153bar (
    .O(ybar[193]),
    .I0(abar[12]),
    .I1(bbar[1])
  );
  //AND U154
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U154 (
    .O(y[192]),
    .I0(a[12]),
    .I1(b[0])
  );
  //OR U154bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U154bar (
    .O(ybar[192]),
    .I0(abar[12]),
    .I1(bbar[0])
  );
  //AND U155
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U155 (
    .O(y[191]),
    .I0(a[11]),
    .I1(b[15])
  );
  //OR U155bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U155bar (
    .O(ybar[191]),
    .I0(abar[11]),
    .I1(bbar[15])
  );
  //AND U156
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U156 (
    .O(y[190]),
    .I0(a[11]),
    .I1(b[14])
  );
  //OR U156bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U156bar (
    .O(ybar[190]),
    .I0(abar[11]),
    .I1(bbar[14])
  );
  //AND U157
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U157 (
    .O(y[18]),
    .I0(a[1]),
    .I1(b[2])
  );
  //OR U157bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U157bar (
    .O(ybar[18]),
    .I0(abar[1]),
    .I1(bbar[2])
  );
  //AND U158
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U158 (
    .O(y[189]),
    .I0(a[11]),
    .I1(b[13])
  );
  //OR U158bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U158bar (
    .O(ybar[189]),
    .I0(abar[11]),
    .I1(bbar[13])
  );
  //AND U159
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U159 (
    .O(y[188]),
    .I0(a[11]),
    .I1(b[12])
  );
  //OR U159bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U159bar (
    .O(ybar[188]),
    .I0(abar[11]),
    .I1(bbar[12])
  );
  //AND U160
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U160 (
    .O(y[187]),
    .I0(a[11]),
    .I1(b[11])
  );
  //OR U160bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U160bar (
    .O(ybar[187]),
    .I0(abar[11]),
    .I1(bbar[11])
  );
  //AND U161
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U161 (
    .O(y[186]),
    .I0(a[11]),
    .I1(b[10])
  );
  //OR U161bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U161bar (
    .O(ybar[186]),
    .I0(abar[11]),
    .I1(bbar[10])
  );
  //AND U162
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U162 (
    .O(y[185]),
    .I0(a[11]),
    .I1(b[9])
  );
  //OR U162bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U162bar (
    .O(ybar[185]),
    .I0(abar[11]),
    .I1(bbar[9])
  );
  //AND U163
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U163 (
    .O(y[184]),
    .I0(a[11]),
    .I1(b[8])
  );
  //OR U163bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U163bar (
    .O(ybar[184]),
    .I0(abar[11]),
    .I1(bbar[8])
  );
  //AND U164
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U164 (
    .O(y[183]),
    .I0(a[11]),
    .I1(b[7])
  );
  //OR U164bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U164bar (
    .O(ybar[183]),
    .I0(abar[11]),
    .I1(bbar[7])
  );
  //AND U165
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U165 (
    .O(y[182]),
    .I0(a[11]),
    .I1(b[6])
  );
  //OR U165bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U165bar (
    .O(ybar[182]),
    .I0(abar[11]),
    .I1(bbar[6])
  );
  //AND U166
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U166 (
    .O(y[181]),
    .I0(a[11]),
    .I1(b[5])
  );
  //OR U166bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U166bar (
    .O(ybar[181]),
    .I0(abar[11]),
    .I1(bbar[5])
  );
  //AND U167
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U167 (
    .O(y[180]),
    .I0(a[11]),
    .I1(b[4])
  );
  //OR U167bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U167bar (
    .O(ybar[180]),
    .I0(abar[11]),
    .I1(bbar[4])
  );
  //AND U168
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U168 (
    .O(y[17]),
    .I0(a[1]),
    .I1(b[1])
  );
  //OR U168bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U168bar (
    .O(ybar[17]),
    .I0(abar[1]),
    .I1(bbar[1])
  );
  //AND U169
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U169 (
    .O(y[179]),
    .I0(a[11]),
    .I1(b[3])
  );
  //OR U169bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U169bar (
    .O(ybar[179]),
    .I0(abar[11]),
    .I1(bbar[3])
  );
  //AND U170
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U170 (
    .O(y[178]),
    .I0(a[11]),
    .I1(b[2])
  );
  //OR U170bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U170bar (
    .O(ybar[178]),
    .I0(abar[11]),
    .I1(bbar[2])
  );
  //AND U171
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U171 (
    .O(y[177]),
    .I0(a[11]),
    .I1(b[1])
  );
  //OR U171bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U171bar (
    .O(ybar[177]),
    .I0(abar[11]),
    .I1(bbar[1])
  );
  //AND U172
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U172 (
    .O(y[176]),
    .I0(a[11]),
    .I1(b[0])
  );
  //OR U172bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U172bar (
    .O(ybar[176]),
    .I0(abar[11]),
    .I1(bbar[0])
  );
  //AND U173
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U173 (
    .O(y[175]),
    .I0(a[10]),
    .I1(b[15])
  );
  //OR U173bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U173bar (
    .O(ybar[175]),
    .I0(abar[10]),
    .I1(bbar[15])
  );
  //AND U174
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U174 (
    .O(y[174]),
    .I0(a[10]),
    .I1(b[14])
  );
  //OR U174bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U174bar (
    .O(ybar[174]),
    .I0(abar[10]),
    .I1(bbar[14])
  );
  //AND U175
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U175 (
    .O(y[173]),
    .I0(a[10]),
    .I1(b[13])
  );
  //OR U175bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U175bar (
    .O(ybar[173]),
    .I0(abar[10]),
    .I1(bbar[13])
  );
  //AND U176
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U176 (
    .O(y[172]),
    .I0(a[10]),
    .I1(b[12])
  );
  //OR U176bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U176bar (
    .O(ybar[172]),
    .I0(abar[10]),
    .I1(bbar[12])
  );
  //AND U177
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U177 (
    .O(y[171]),
    .I0(a[10]),
    .I1(b[11])
  );
  //OR U177bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U177bar (
    .O(ybar[171]),
    .I0(abar[10]),
    .I1(bbar[11])
  );
  //AND U178
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U178 (
    .O(y[170]),
    .I0(a[10]),
    .I1(b[10])
  );
  //OR U178bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U178bar (
    .O(ybar[170]),
    .I0(abar[10]),
    .I1(bbar[10])
  );
  //AND U179
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U179 (
    .O(y[16]),
    .I0(a[1]),
    .I1(b[0])
  );
  //OR U179bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U179bar (
    .O(ybar[16]),
    .I0(abar[1]),
    .I1(bbar[0])
  );
  //AND U180
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U180 (
    .O(y[169]),
    .I0(a[10]),
    .I1(b[9])
  );
  //OR U180bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U180bar (
    .O(ybar[169]),
    .I0(abar[10]),
    .I1(bbar[9])
  );
  //AND U181
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U181 (
    .O(y[168]),
    .I0(a[10]),
    .I1(b[8])
  );
  //OR U181bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U181bar (
    .O(ybar[168]),
    .I0(abar[10]),
    .I1(bbar[8])
  );
  //AND U182
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U182 (
    .O(y[167]),
    .I0(a[10]),
    .I1(b[7])
  );
  //OR U182bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U182bar (
    .O(ybar[167]),
    .I0(abar[10]),
    .I1(bbar[7])
  );
  //AND U183
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U183 (
    .O(y[166]),
    .I0(a[10]),
    .I1(b[6])
  );
  //OR U183bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U183bar (
    .O(ybar[166]),
    .I0(abar[10]),
    .I1(bbar[6])
  );
  //AND U184
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U184 (
    .O(y[165]),
    .I0(a[10]),
    .I1(b[5])
  );
  //OR U184bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U184bar (
    .O(ybar[165]),
    .I0(abar[10]),
    .I1(bbar[5])
  );
  //AND U185
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U185 (
    .O(y[164]),
    .I0(a[10]),
    .I1(b[4])
  );
  //OR U185bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U185bar (
    .O(ybar[164]),
    .I0(abar[10]),
    .I1(bbar[4])
  );
  //AND U186
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U186 (
    .O(y[163]),
    .I0(a[10]),
    .I1(b[3])
  );
  //OR U186bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U186bar (
    .O(ybar[163]),
    .I0(abar[10]),
    .I1(bbar[3])
  );
  //AND U187
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U187 (
    .O(y[162]),
    .I0(a[10]),
    .I1(b[2])
  );
  //OR U187bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U187bar (
    .O(ybar[162]),
    .I0(abar[10]),
    .I1(bbar[2])
  );
  //AND U188
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U188 (
    .O(y[161]),
    .I0(a[10]),
    .I1(b[1])
  );
  //OR U188bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U188bar (
    .O(ybar[161]),
    .I0(abar[10]),
    .I1(bbar[1])
  );
  //AND U189
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U189 (
    .O(y[160]),
    .I0(a[10]),
    .I1(b[0])
  );
  //OR U189bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U189bar (
    .O(ybar[160]),
    .I0(abar[10]),
    .I1(bbar[0])
  );
  //AND U190
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U190 (
    .O(y[15]),
    .I0(b[15]),
    .I1(a[0])
  );
  //OR U190bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U190bar (
    .O(ybar[15]),
    .I0(bbar[15]),
    .I1(abar[0])
  );
  //AND U191
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U191 (
    .O(y[159]),
    .I0(a[9]),
    .I1(b[15])
  );
  //OR U191bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U191bar (
    .O(ybar[159]),
    .I0(abar[9]),
    .I1(bbar[15])
  );
  //AND U192
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U192 (
    .O(y[158]),
    .I0(a[9]),
    .I1(b[14])
  );
  //OR U192bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U192bar (
    .O(ybar[158]),
    .I0(abar[9]),
    .I1(bbar[14])
  );
  //AND U193
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U193 (
    .O(y[157]),
    .I0(a[9]),
    .I1(b[13])
  );
  //OR U193bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U193bar (
    .O(ybar[157]),
    .I0(abar[9]),
    .I1(bbar[13])
  );
  //AND U194
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U194 (
    .O(y[156]),
    .I0(a[9]),
    .I1(b[12])
  );
  //OR U194bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U194bar (
    .O(ybar[156]),
    .I0(abar[9]),
    .I1(bbar[12])
  );
  //AND U195
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U195 (
    .O(y[155]),
    .I0(a[9]),
    .I1(b[11])
  );
  //OR U195bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U195bar (
    .O(ybar[155]),
    .I0(abar[9]),
    .I1(bbar[11])
  );
  //AND U196
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U196 (
    .O(y[154]),
    .I0(a[9]),
    .I1(b[10])
  );
  //OR U196bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U196bar (
    .O(ybar[154]),
    .I0(abar[9]),
    .I1(bbar[10])
  );
  //AND U197
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U197 (
    .O(y[153]),
    .I0(a[9]),
    .I1(b[9])
  );
  //OR U197bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U197bar (
    .O(ybar[153]),
    .I0(abar[9]),
    .I1(bbar[9])
  );
  //AND U198
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U198 (
    .O(y[152]),
    .I0(a[9]),
    .I1(b[8])
  );
  //OR U198bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U198bar (
    .O(ybar[152]),
    .I0(abar[9]),
    .I1(bbar[8])
  );
  //AND U199
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U199 (
    .O(y[151]),
    .I0(a[9]),
    .I1(b[7])
  );
  //OR U199bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U199bar (
    .O(ybar[151]),
    .I0(abar[9]),
    .I1(bbar[7])
  );
  //AND U200
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U200 (
    .O(y[150]),
    .I0(a[9]),
    .I1(b[6])
  );
  //OR U200bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U200bar (
    .O(ybar[150]),
    .I0(abar[9]),
    .I1(bbar[6])
  );
  //AND U201
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U201 (
    .O(y[14]),
    .I0(b[14]),
    .I1(a[0])
  );
  //OR U201bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U201bar (
    .O(ybar[14]),
    .I0(bbar[14]),
    .I1(abar[0])
  );
  //AND U202
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U202 (
    .O(y[149]),
    .I0(a[9]),
    .I1(b[5])
  );
  //OR U202bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U202bar (
    .O(ybar[149]),
    .I0(abar[9]),
    .I1(bbar[5])
  );
  //AND U203
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U203 (
    .O(y[148]),
    .I0(a[9]),
    .I1(b[4])
  );
  //OR U203bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U203bar (
    .O(ybar[148]),
    .I0(abar[9]),
    .I1(bbar[4])
  );
  //AND U204
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U204 (
    .O(y[147]),
    .I0(a[9]),
    .I1(b[3])
  );
  //OR U204bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U204bar (
    .O(ybar[147]),
    .I0(abar[9]),
    .I1(bbar[3])
  );
  //AND U205
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U205 (
    .O(y[146]),
    .I0(a[9]),
    .I1(b[2])
  );
  //OR U205bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U205bar (
    .O(ybar[146]),
    .I0(abar[9]),
    .I1(bbar[2])
  );
  //AND U206
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U206 (
    .O(y[145]),
    .I0(a[9]),
    .I1(b[1])
  );
  //OR U206bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U206bar (
    .O(ybar[145]),
    .I0(abar[9]),
    .I1(bbar[1])
  );
  //AND U207
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U207 (
    .O(y[144]),
    .I0(a[9]),
    .I1(b[0])
  );
  //OR U207bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U207bar (
    .O(ybar[144]),
    .I0(abar[9]),
    .I1(bbar[0])
  );
  //AND U208
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U208 (
    .O(y[143]),
    .I0(a[8]),
    .I1(b[15])
  );
  //OR U208bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U208bar (
    .O(ybar[143]),
    .I0(abar[8]),
    .I1(bbar[15])
  );
  //AND U209
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U209 (
    .O(y[142]),
    .I0(a[8]),
    .I1(b[14])
  );
  //OR U209bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U209bar (
    .O(ybar[142]),
    .I0(abar[8]),
    .I1(bbar[14])
  );
  //AND U210
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U210 (
    .O(y[141]),
    .I0(a[8]),
    .I1(b[13])
  );
  //OR U210bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U210bar (
    .O(ybar[141]),
    .I0(abar[8]),
    .I1(bbar[13])
  );
  //AND U211
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U211 (
    .O(y[140]),
    .I0(a[8]),
    .I1(b[12])
  );
  //OR U211bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U211bar (
    .O(ybar[140]),
    .I0(abar[8]),
    .I1(bbar[12])
  );
  //AND U212
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U212 (
    .O(y[13]),
    .I0(b[13]),
    .I1(a[0])
  );
  //OR U212bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U212bar (
    .O(ybar[13]),
    .I0(bbar[13]),
    .I1(abar[0])
  );
  //AND U213
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U213 (
    .O(y[139]),
    .I0(a[8]),
    .I1(b[11])
  );
  //OR U213bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U213bar (
    .O(ybar[139]),
    .I0(abar[8]),
    .I1(bbar[11])
  );
  //AND U214
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U214 (
    .O(y[138]),
    .I0(a[8]),
    .I1(b[10])
  );
  //OR U214bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U214bar (
    .O(ybar[138]),
    .I0(abar[8]),
    .I1(bbar[10])
  );
  //AND U215
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U215 (
    .O(y[137]),
    .I0(a[8]),
    .I1(b[9])
  );
  //OR U215bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U215bar (
    .O(ybar[137]),
    .I0(abar[8]),
    .I1(bbar[9])
  );
  //AND U216
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U216 (
    .O(y[136]),
    .I0(a[8]),
    .I1(b[8])
  );
  //OR U216bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U216bar (
    .O(ybar[136]),
    .I0(abar[8]),
    .I1(bbar[8])
  );
  //AND U217
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U217 (
    .O(y[135]),
    .I0(a[8]),
    .I1(b[7])
  );
  //OR U217bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U217bar (
    .O(ybar[135]),
    .I0(abar[8]),
    .I1(bbar[7])
  );
  //AND U218
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U218 (
    .O(y[134]),
    .I0(a[8]),
    .I1(b[6])
  );
  //OR U218bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U218bar (
    .O(ybar[134]),
    .I0(abar[8]),
    .I1(bbar[6])
  );
  //AND U219
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U219 (
    .O(y[133]),
    .I0(a[8]),
    .I1(b[5])
  );
  //OR U219bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U219bar (
    .O(ybar[133]),
    .I0(abar[8]),
    .I1(bbar[5])
  );
  //AND U220
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U220 (
    .O(y[132]),
    .I0(a[8]),
    .I1(b[4])
  );
  //OR U220bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U220bar (
    .O(ybar[132]),
    .I0(abar[8]),
    .I1(bbar[4])
  );
  //AND U221
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U221 (
    .O(y[131]),
    .I0(a[8]),
    .I1(b[3])
  );
  //OR U221bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U221bar (
    .O(ybar[131]),
    .I0(abar[8]),
    .I1(bbar[3])
  );
  //AND U222
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U222 (
    .O(y[130]),
    .I0(a[8]),
    .I1(b[2])
  );
  //OR U222bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U222bar (
    .O(ybar[130]),
    .I0(abar[8]),
    .I1(bbar[2])
  );
  //AND U223
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U223 (
    .O(y[12]),
    .I0(b[12]),
    .I1(a[0])
  );
  //OR U223bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U223bar (
    .O(ybar[12]),
    .I0(bbar[12]),
    .I1(abar[0])
  );
  //AND U224
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U224 (
    .O(y[129]),
    .I0(a[8]),
    .I1(b[1])
  );
  //OR U224bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U224bar (
    .O(ybar[129]),
    .I0(abar[8]),
    .I1(bbar[1])
  );
  //AND U225
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U225 (
    .O(y[128]),
    .I0(a[8]),
    .I1(b[0])
  );
  //OR U225bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U225bar (
    .O(ybar[128]),
    .I0(abar[8]),
    .I1(bbar[0])
  );
  //AND U226
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U226 (
    .O(y[127]),
    .I0(a[7]),
    .I1(b[15])
  );
  //OR U226bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U226bar (
    .O(ybar[127]),
    .I0(abar[7]),
    .I1(bbar[15])
  );
  //AND U227
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U227 (
    .O(y[126]),
    .I0(a[7]),
    .I1(b[14])
  );
  //OR U227bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U227bar (
    .O(ybar[126]),
    .I0(abar[7]),
    .I1(bbar[14])
  );
  //AND U228
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U228 (
    .O(y[125]),
    .I0(a[7]),
    .I1(b[13])
  );
  //OR U228bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U228bar (
    .O(ybar[125]),
    .I0(abar[7]),
    .I1(bbar[13])
  );
  //AND U229
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U229 (
    .O(y[124]),
    .I0(a[7]),
    .I1(b[12])
  );
  //OR U229bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U229bar (
    .O(ybar[124]),
    .I0(abar[7]),
    .I1(bbar[12])
  );
  //AND U230
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U230 (
    .O(y[123]),
    .I0(a[7]),
    .I1(b[11])
  );
  //OR U230bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U230bar (
    .O(ybar[123]),
    .I0(abar[7]),
    .I1(bbar[11])
  );
  //AND U231
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U231 (
    .O(y[122]),
    .I0(a[7]),
    .I1(b[10])
  );
  //OR U231bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U231bar (
    .O(ybar[122]),
    .I0(abar[7]),
    .I1(bbar[10])
  );
  //AND U232
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U232 (
    .O(y[121]),
    .I0(a[7]),
    .I1(b[9])
  );
  //OR U232bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U232bar (
    .O(ybar[121]),
    .I0(abar[7]),
    .I1(bbar[9])
  );
  //AND U233
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U233 (
    .O(y[120]),
    .I0(a[7]),
    .I1(b[8])
  );
  //OR U233bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U233bar (
    .O(ybar[120]),
    .I0(abar[7]),
    .I1(bbar[8])
  );
  //AND U234
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U234 (
    .O(y[11]),
    .I0(b[11]),
    .I1(a[0])
  );
  //OR U234bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U234bar (
    .O(ybar[11]),
    .I0(bbar[11]),
    .I1(abar[0])
  );
  //AND U235
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U235 (
    .O(y[119]),
    .I0(a[7]),
    .I1(b[7])
  );
  //OR U235bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U235bar (
    .O(ybar[119]),
    .I0(abar[7]),
    .I1(bbar[7])
  );
  //AND U236
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U236 (
    .O(y[118]),
    .I0(a[7]),
    .I1(b[6])
  );
  //OR U236bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U236bar (
    .O(ybar[118]),
    .I0(abar[7]),
    .I1(bbar[6])
  );
  //AND U237
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U237 (
    .O(y[117]),
    .I0(a[7]),
    .I1(b[5])
  );
  //OR U237bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U237bar (
    .O(ybar[117]),
    .I0(abar[7]),
    .I1(bbar[5])
  );
  //AND U238
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U238 (
    .O(y[116]),
    .I0(a[7]),
    .I1(b[4])
  );
  //OR U238bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U238bar (
    .O(ybar[116]),
    .I0(abar[7]),
    .I1(bbar[4])
  );
  //AND U239
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U239 (
    .O(y[115]),
    .I0(a[7]),
    .I1(b[3])
  );
  //OR U239bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U239bar (
    .O(ybar[115]),
    .I0(abar[7]),
    .I1(bbar[3])
  );
  //AND U240
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U240 (
    .O(y[114]),
    .I0(a[7]),
    .I1(b[2])
  );
  //OR U240bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U240bar (
    .O(ybar[114]),
    .I0(abar[7]),
    .I1(bbar[2])
  );
  //AND U241
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U241 (
    .O(y[113]),
    .I0(a[7]),
    .I1(b[1])
  );
  //OR U241bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U241bar (
    .O(ybar[113]),
    .I0(abar[7]),
    .I1(bbar[1])
  );
  //AND U242
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U242 (
    .O(y[112]),
    .I0(a[7]),
    .I1(b[0])
  );
  //OR U242bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U242bar (
    .O(ybar[112]),
    .I0(abar[7]),
    .I1(bbar[0])
  );
  //AND U243
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U243 (
    .O(y[111]),
    .I0(b[15]),
    .I1(a[6])
  );
  //OR U243bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U243bar (
    .O(ybar[111]),
    .I0(bbar[15]),
    .I1(abar[6])
  );
  //AND U244
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U244 (
    .O(y[110]),
    .I0(b[14]),
    .I1(a[6])
  );
  //OR U244bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U244bar (
    .O(ybar[110]),
    .I0(bbar[14]),
    .I1(abar[6])
  );
  //AND U245
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U245 (
    .O(y[10]),
    .I0(b[10]),
    .I1(a[0])
  );
  //OR U245bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U245bar (
    .O(ybar[10]),
    .I0(bbar[10]),
    .I1(abar[0])
  );
  //AND U246
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U246 (
    .O(y[109]),
    .I0(b[13]),
    .I1(a[6])
  );
  //OR U246bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U246bar (
    .O(ybar[109]),
    .I0(bbar[13]),
    .I1(abar[6])
  );
  //AND U247
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U247 (
    .O(y[108]),
    .I0(b[12]),
    .I1(a[6])
  );
  //OR U247bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U247bar (
    .O(ybar[108]),
    .I0(bbar[12]),
    .I1(abar[6])
  );
  //AND U248
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U248 (
    .O(y[107]),
    .I0(b[11]),
    .I1(a[6])
  );
  //OR U248bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U248bar (
    .O(ybar[107]),
    .I0(bbar[11]),
    .I1(abar[6])
  );
  //AND U249
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U249 (
    .O(y[106]),
    .I0(b[10]),
    .I1(a[6])
  );
  //OR U249bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U249bar (
    .O(ybar[106]),
    .I0(bbar[10]),
    .I1(abar[6])
  );
  //AND U250
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U250 (
    .O(y[105]),
    .I0(a[6]),
    .I1(b[9])
  );
  //OR U250bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U250bar (
    .O(ybar[105]),
    .I0(abar[6]),
    .I1(bbar[9])
  );
  //AND U251
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U251 (
    .O(y[104]),
    .I0(b[8]),
    .I1(a[6])
  );
  //OR U251bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U251bar (
    .O(ybar[104]),
    .I0(bbar[8]),
    .I1(abar[6])
  );
  //AND U252
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U252 (
    .O(y[103]),
    .I0(b[7]),
    .I1(a[6])
  );
  //OR U252bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U252bar (
    .O(ybar[103]),
    .I0(bbar[7]),
    .I1(abar[6])
  );
  //AND U253
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U253 (
    .O(y[102]),
    .I0(b[6]),
    .I1(a[6])
  );
  //OR U253bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U253bar (
    .O(ybar[102]),
    .I0(bbar[6]),
    .I1(abar[6])
  );
  //AND U254
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U254 (
    .O(y[101]),
    .I0(b[5]),
    .I1(a[6])
  );
  //OR U254bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U254bar (
    .O(ybar[101]),
    .I0(bbar[5]),
    .I1(abar[6])
  );
  //AND U255
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U255 (
    .O(y[100]),
    .I0(b[4]),
    .I1(a[6])
  );
  //OR U255bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U255bar (
    .O(ybar[100]),
    .I0(bbar[4]),
    .I1(abar[6])
  );
  //AND U256
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U256 (
    .O(y[0]),
    .I0(b[0]),
    .I1(a[0])
  );
  //OR U256bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U256bar (
    .O(ybar[0]),
    .I0(bbar[0]),
    .I1(abar[0])
  );
endmodule

module decode_10 ( in, out );

  input wire [7:0] in;
//input_done

  output wire [255:0] out;
//output_done

  wire [15:0] level1;
  wire [31:0] level2;
//wire_done

  CD2_40 cd_l1_1 ( .a(in[1]), .b(in[0]), .y(level1[3:0]) );
  CD2_39 cd_l1_2 ( .a(in[3]), .b(in[2]), .y(level1[7:4]) );
  CD2_38 cd_l1_3 ( .a(in[5]), .b(in[4]), .y(level1[11:8]) );
  CD2_37 cd_l1_4 ( .a(in[7]), .b(in[6]), .y(level1[15:12]) );
  CD4_20 cd_l2_1 ( .a(level1[7:4]), .b(level1[3:0]), .y(level2[15:0]) );
  CD4_19 cd_l2_2 ( .a(level1[15:12]), .b(level1[11:8]), .y(level2[31:16]) );
  CD16_10 cd_l3 ( .a(level2[31:16]), .b(level2[15:0]), .y(out) );
endmodule

module encode_10 ( in, out );

  input wire [255:0] in;
  wire [255:0] inbar;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
  assign inbar[8] = ~in[8];
  assign inbar[9] = ~in[9];
  assign inbar[10] = ~in[10];
  assign inbar[11] = ~in[11];
  assign inbar[12] = ~in[12];
  assign inbar[13] = ~in[13];
  assign inbar[14] = ~in[14];
  assign inbar[15] = ~in[15];
  assign inbar[16] = ~in[16];
  assign inbar[17] = ~in[17];
  assign inbar[18] = ~in[18];
  assign inbar[19] = ~in[19];
  assign inbar[20] = ~in[20];
  assign inbar[21] = ~in[21];
  assign inbar[22] = ~in[22];
  assign inbar[23] = ~in[23];
  assign inbar[24] = ~in[24];
  assign inbar[25] = ~in[25];
  assign inbar[26] = ~in[26];
  assign inbar[27] = ~in[27];
  assign inbar[28] = ~in[28];
  assign inbar[29] = ~in[29];
  assign inbar[30] = ~in[30];
  assign inbar[31] = ~in[31];
  assign inbar[32] = ~in[32];
  assign inbar[33] = ~in[33];
  assign inbar[34] = ~in[34];
  assign inbar[35] = ~in[35];
  assign inbar[36] = ~in[36];
  assign inbar[37] = ~in[37];
  assign inbar[38] = ~in[38];
  assign inbar[39] = ~in[39];
  assign inbar[40] = ~in[40];
  assign inbar[41] = ~in[41];
  assign inbar[42] = ~in[42];
  assign inbar[43] = ~in[43];
  assign inbar[44] = ~in[44];
  assign inbar[45] = ~in[45];
  assign inbar[46] = ~in[46];
  assign inbar[47] = ~in[47];
  assign inbar[48] = ~in[48];
  assign inbar[49] = ~in[49];
  assign inbar[50] = ~in[50];
  assign inbar[51] = ~in[51];
  assign inbar[52] = ~in[52];
  assign inbar[53] = ~in[53];
  assign inbar[54] = ~in[54];
  assign inbar[55] = ~in[55];
  assign inbar[56] = ~in[56];
  assign inbar[57] = ~in[57];
  assign inbar[58] = ~in[58];
  assign inbar[59] = ~in[59];
  assign inbar[60] = ~in[60];
  assign inbar[61] = ~in[61];
  assign inbar[62] = ~in[62];
  assign inbar[63] = ~in[63];
  assign inbar[64] = ~in[64];
  assign inbar[65] = ~in[65];
  assign inbar[66] = ~in[66];
  assign inbar[67] = ~in[67];
  assign inbar[68] = ~in[68];
  assign inbar[69] = ~in[69];
  assign inbar[70] = ~in[70];
  assign inbar[71] = ~in[71];
  assign inbar[72] = ~in[72];
  assign inbar[73] = ~in[73];
  assign inbar[74] = ~in[74];
  assign inbar[75] = ~in[75];
  assign inbar[76] = ~in[76];
  assign inbar[77] = ~in[77];
  assign inbar[78] = ~in[78];
  assign inbar[79] = ~in[79];
  assign inbar[80] = ~in[80];
  assign inbar[81] = ~in[81];
  assign inbar[82] = ~in[82];
  assign inbar[83] = ~in[83];
  assign inbar[84] = ~in[84];
  assign inbar[85] = ~in[85];
  assign inbar[86] = ~in[86];
  assign inbar[87] = ~in[87];
  assign inbar[88] = ~in[88];
  assign inbar[89] = ~in[89];
  assign inbar[90] = ~in[90];
  assign inbar[91] = ~in[91];
  assign inbar[92] = ~in[92];
  assign inbar[93] = ~in[93];
  assign inbar[94] = ~in[94];
  assign inbar[95] = ~in[95];
  assign inbar[96] = ~in[96];
  assign inbar[97] = ~in[97];
  assign inbar[98] = ~in[98];
  assign inbar[99] = ~in[99];
  assign inbar[100] = ~in[100];
  assign inbar[101] = ~in[101];
  assign inbar[102] = ~in[102];
  assign inbar[103] = ~in[103];
  assign inbar[104] = ~in[104];
  assign inbar[105] = ~in[105];
  assign inbar[106] = ~in[106];
  assign inbar[107] = ~in[107];
  assign inbar[108] = ~in[108];
  assign inbar[109] = ~in[109];
  assign inbar[110] = ~in[110];
  assign inbar[111] = ~in[111];
  assign inbar[112] = ~in[112];
  assign inbar[113] = ~in[113];
  assign inbar[114] = ~in[114];
  assign inbar[115] = ~in[115];
  assign inbar[116] = ~in[116];
  assign inbar[117] = ~in[117];
  assign inbar[118] = ~in[118];
  assign inbar[119] = ~in[119];
  assign inbar[120] = ~in[120];
  assign inbar[121] = ~in[121];
  assign inbar[122] = ~in[122];
  assign inbar[123] = ~in[123];
  assign inbar[124] = ~in[124];
  assign inbar[125] = ~in[125];
  assign inbar[126] = ~in[126];
  assign inbar[127] = ~in[127];
  assign inbar[128] = ~in[128];
  assign inbar[129] = ~in[129];
  assign inbar[130] = ~in[130];
  assign inbar[131] = ~in[131];
  assign inbar[132] = ~in[132];
  assign inbar[133] = ~in[133];
  assign inbar[134] = ~in[134];
  assign inbar[135] = ~in[135];
  assign inbar[136] = ~in[136];
  assign inbar[137] = ~in[137];
  assign inbar[138] = ~in[138];
  assign inbar[139] = ~in[139];
  assign inbar[140] = ~in[140];
  assign inbar[141] = ~in[141];
  assign inbar[142] = ~in[142];
  assign inbar[143] = ~in[143];
  assign inbar[144] = ~in[144];
  assign inbar[145] = ~in[145];
  assign inbar[146] = ~in[146];
  assign inbar[147] = ~in[147];
  assign inbar[148] = ~in[148];
  assign inbar[149] = ~in[149];
  assign inbar[150] = ~in[150];
  assign inbar[151] = ~in[151];
  assign inbar[152] = ~in[152];
  assign inbar[153] = ~in[153];
  assign inbar[154] = ~in[154];
  assign inbar[155] = ~in[155];
  assign inbar[156] = ~in[156];
  assign inbar[157] = ~in[157];
  assign inbar[158] = ~in[158];
  assign inbar[159] = ~in[159];
  assign inbar[160] = ~in[160];
  assign inbar[161] = ~in[161];
  assign inbar[162] = ~in[162];
  assign inbar[163] = ~in[163];
  assign inbar[164] = ~in[164];
  assign inbar[165] = ~in[165];
  assign inbar[166] = ~in[166];
  assign inbar[167] = ~in[167];
  assign inbar[168] = ~in[168];
  assign inbar[169] = ~in[169];
  assign inbar[170] = ~in[170];
  assign inbar[171] = ~in[171];
  assign inbar[172] = ~in[172];
  assign inbar[173] = ~in[173];
  assign inbar[174] = ~in[174];
  assign inbar[175] = ~in[175];
  assign inbar[176] = ~in[176];
  assign inbar[177] = ~in[177];
  assign inbar[178] = ~in[178];
  assign inbar[179] = ~in[179];
  assign inbar[180] = ~in[180];
  assign inbar[181] = ~in[181];
  assign inbar[182] = ~in[182];
  assign inbar[183] = ~in[183];
  assign inbar[184] = ~in[184];
  assign inbar[185] = ~in[185];
  assign inbar[186] = ~in[186];
  assign inbar[187] = ~in[187];
  assign inbar[188] = ~in[188];
  assign inbar[189] = ~in[189];
  assign inbar[190] = ~in[190];
  assign inbar[191] = ~in[191];
  assign inbar[192] = ~in[192];
  assign inbar[193] = ~in[193];
  assign inbar[194] = ~in[194];
  assign inbar[195] = ~in[195];
  assign inbar[196] = ~in[196];
  assign inbar[197] = ~in[197];
  assign inbar[198] = ~in[198];
  assign inbar[199] = ~in[199];
  assign inbar[200] = ~in[200];
  assign inbar[201] = ~in[201];
  assign inbar[202] = ~in[202];
  assign inbar[203] = ~in[203];
  assign inbar[204] = ~in[204];
  assign inbar[205] = ~in[205];
  assign inbar[206] = ~in[206];
  assign inbar[207] = ~in[207];
  assign inbar[208] = ~in[208];
  assign inbar[209] = ~in[209];
  assign inbar[210] = ~in[210];
  assign inbar[211] = ~in[211];
  assign inbar[212] = ~in[212];
  assign inbar[213] = ~in[213];
  assign inbar[214] = ~in[214];
  assign inbar[215] = ~in[215];
  assign inbar[216] = ~in[216];
  assign inbar[217] = ~in[217];
  assign inbar[218] = ~in[218];
  assign inbar[219] = ~in[219];
  assign inbar[220] = ~in[220];
  assign inbar[221] = ~in[221];
  assign inbar[222] = ~in[222];
  assign inbar[223] = ~in[223];
  assign inbar[224] = ~in[224];
  assign inbar[225] = ~in[225];
  assign inbar[226] = ~in[226];
  assign inbar[227] = ~in[227];
  assign inbar[228] = ~in[228];
  assign inbar[229] = ~in[229];
  assign inbar[230] = ~in[230];
  assign inbar[231] = ~in[231];
  assign inbar[232] = ~in[232];
  assign inbar[233] = ~in[233];
  assign inbar[234] = ~in[234];
  assign inbar[235] = ~in[235];
  assign inbar[236] = ~in[236];
  assign inbar[237] = ~in[237];
  assign inbar[238] = ~in[238];
  assign inbar[239] = ~in[239];
  assign inbar[240] = ~in[240];
  assign inbar[241] = ~in[241];
  assign inbar[242] = ~in[242];
  assign inbar[243] = ~in[243];
  assign inbar[244] = ~in[244];
  assign inbar[245] = ~in[245];
  assign inbar[246] = ~in[246];
  assign inbar[247] = ~in[247];
  assign inbar[248] = ~in[248];
  assign inbar[249] = ~in[249];
  assign inbar[250] = ~in[250];
  assign inbar[251] = ~in[251];
  assign inbar[252] = ~in[252];
  assign inbar[253] = ~in[253];
  assign inbar[254] = ~in[254];
  assign inbar[255] = ~in[255];
//input_done

  output wire [7:0] out;
  wire [7:0] outbar;
//output_done

  wire in_81;
  wire in_80;
  wire in_79;
  wire in_78;
  wire in_77;
  wire in_76;
  wire in_75;
  wire in_74;
  wire in_73;
  wire in_72;
  wire in_71;
  wire in_70;
  wire in_69;
  wire in_68;
  wire in_67;
  wire in_66;
  wire in_65;
  wire in_64;
  wire in_63;
  wire in_62;
  wire in_61;
  wire in_60;
  wire in_59;
  wire in_58;
  wire in_57;
  wire in_56;
  wire in_55;
  wire in_54;
  wire in_53;
  wire in_52;
  wire in_51;
  wire in_50;
  wire in_49;
  wire in_48;
  wire in_47;
  wire in_46;
  wire in_45;
  wire in_44;
  wire in_43;
  wire in_42;
  wire in_41;
  wire in_40;
  wire in_39;
  wire in_38;
  wire in_37;
  wire in_36;
  wire in_35;
  wire in_34;
  wire in_33;
  wire in_32;
  wire in_31;
  wire in_30;
  wire in_29;
  wire in_28;
  wire in_27;
  wire in_26;
  wire in_25;
  wire in_24;
  wire in_23;
  wire in_22;
  wire in_21;
  wire in_20;
  wire in_19;
  wire in_18;
  wire in_17;
  wire in_16;
  wire in_15;
  wire in_14;
  wire in_13;
  wire in_12;
  wire in_11;
  wire in_10;
  wire in_9;
  wire in_8;
  wire in_7;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_3;
  wire in_2;
  wire in_1;
  wire in_0;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire in_81bar;
  wire in_80bar;
  wire in_79bar;
  wire in_78bar;
  wire in_77bar;
  wire in_76bar;
  wire in_75bar;
  wire in_74bar;
  wire in_73bar;
  wire in_72bar;
  wire in_71bar;
  wire in_70bar;
  wire in_69bar;
  wire in_68bar;
  wire in_67bar;
  wire in_66bar;
  wire in_65bar;
  wire in_64bar;
  wire in_63bar;
  wire in_62bar;
  wire in_61bar;
  wire in_60bar;
  wire in_59bar;
  wire in_58bar;
  wire in_57bar;
  wire in_56bar;
  wire in_55bar;
  wire in_54bar;
  wire in_53bar;
  wire in_52bar;
  wire in_51bar;
  wire in_50bar;
  wire in_49bar;
  wire in_48bar;
  wire in_47bar;
  wire in_46bar;
  wire in_45bar;
  wire in_44bar;
  wire in_43bar;
  wire in_42bar;
  wire in_41bar;
  wire in_40bar;
  wire in_39bar;
  wire in_38bar;
  wire in_37bar;
  wire in_36bar;
  wire in_35bar;
  wire in_34bar;
  wire in_33bar;
  wire in_32bar;
  wire in_31bar;
  wire in_30bar;
  wire in_29bar;
  wire in_28bar;
  wire in_27bar;
  wire in_26bar;
  wire in_25bar;
  wire in_24bar;
  wire in_23bar;
  wire in_22bar;
  wire in_21bar;
  wire in_20bar;
  wire in_19bar;
  wire in_18bar;
  wire in_17bar;
  wire in_16bar;
  wire in_15bar;
  wire in_14bar;
  wire in_13bar;
  wire in_12bar;
  wire in_11bar;
  wire in_10bar;
  wire in_9bar;
  wire in_8bar;
  wire in_7bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_3bar;
  wire in_2bar;
  wire in_1bar;
  wire in_0bar;
  wire n487bar;
  wire n488bar;
  wire n489bar;
  wire n490bar;
  wire n491bar;
  wire n492bar;
  wire n493bar;
  wire n494bar;
  wire n495bar;
  wire n496bar;
  wire n497bar;
  wire n498bar;
  wire n499bar;
  wire n500bar;
  wire n501bar;
  wire n502bar;
  wire n503bar;
  wire n504bar;
  wire n505bar;
  wire n506bar;
  wire n507bar;
  wire n508bar;
  wire n509bar;
  wire n510bar;
  wire n511bar;
  wire n512bar;
  wire n513bar;
  wire n514bar;
  wire n515bar;
  wire n516bar;
  wire n517bar;
  wire n518bar;
  wire n519bar;
  wire n520bar;
  wire n521bar;
  wire n522bar;
  wire n523bar;
  wire n524bar;
  wire n525bar;
  wire n526bar;
  wire n527bar;
  wire n528bar;
  wire n529bar;
  wire n530bar;
  wire n531bar;
  wire n532bar;
  wire n533bar;
  wire n534bar;
  wire n535bar;
  wire n536bar;
  wire n537bar;
  wire n538bar;
  wire n539bar;
  wire n540bar;
  wire n541bar;
  wire n542bar;
  wire n543bar;
  wire n544bar;
  wire n545bar;
  wire n546bar;
  wire n547bar;
  wire n548bar;
  wire n549bar;
  wire n550bar;
  wire n551bar;
  wire n552bar;
  wire n553bar;
  wire n554bar;
  wire n555bar;
  wire n556bar;
  wire n557bar;
  wire n558bar;
  wire n559bar;
  wire n560bar;
  wire n561bar;
  wire n562bar;
  wire n563bar;
  wire n564bar;
  wire n565bar;
  wire n566bar;
  wire n567bar;
  wire n568bar;
  wire n569bar;
  wire n570bar;
  wire n571bar;
  wire n572bar;
  wire n573bar;
  wire n574bar;
  wire n575bar;
  wire n576bar;
  wire n577bar;
  wire n578bar;
  wire n579bar;
  wire n580bar;
  wire n581bar;
  wire n582bar;
  wire n583bar;
  wire n584bar;
  wire n585bar;
  wire n586bar;
  wire n587bar;
  wire n588bar;
  wire n589bar;
  wire n590bar;
  wire n591bar;
  wire n592bar;
  wire n593bar;
  wire n594bar;
  wire n595bar;
  wire n596bar;
  wire n597bar;
  wire n598bar;
  wire n599bar;
  wire n600bar;
  wire n601bar;
  wire n602bar;
  wire n603bar;
  wire n604bar;
  wire n605bar;
  wire n606bar;
  wire n607bar;
  wire n608bar;
  wire n609bar;
  wire n610bar;
  wire n611bar;
  wire n612bar;
  wire n613bar;
  wire n614bar;
  wire n615bar;
  wire n616bar;
  wire n617bar;
  wire n618bar;
  wire n619bar;
  wire n620bar;
  wire n621bar;
  wire n622bar;
  wire n623bar;
  wire n624bar;
  wire n625bar;
  wire n626bar;
  wire n627bar;
  wire n628bar;
  wire n629bar;
  wire n630bar;
  wire n631bar;
  wire n632bar;
  wire n633bar;
  wire n634bar;
  wire n635bar;
  wire n636bar;
  wire n637bar;
  wire n638bar;
  wire n639bar;
  wire n640bar;
  wire n641bar;
  wire n642bar;
  wire n643bar;
  wire n644bar;
  wire n645bar;
  wire n646bar;
  wire n647bar;
  wire n648bar;
  wire n649bar;
  wire n650bar;
  wire n651bar;
  wire n652bar;
  wire n653bar;
  wire n654bar;
  wire n655bar;
  wire n656bar;
  wire n657bar;
  wire n658bar;
  wire n659bar;
  wire n660bar;
  wire n661bar;
  wire n662bar;
  wire n663bar;
  wire n664bar;
  wire n665bar;
  wire n666bar;
  wire n667bar;
  wire n668bar;
  wire n669bar;
  wire n670bar;
  wire n671bar;
  wire n672bar;
  wire n673bar;
  wire n674bar;
  wire n675bar;
  wire n676bar;
  wire n677bar;
  wire n678bar;
  wire n679bar;
  wire n680bar;
  wire n681bar;
  wire n682bar;
  wire n683bar;
  wire n684bar;
  wire n685bar;
  wire n686bar;
  wire n687bar;
  wire n688bar;
  wire n689bar;
  wire n690bar;
  wire n691bar;
  wire n692bar;
  wire n693bar;
  wire n694bar;
  wire n695bar;
  wire n696bar;
  wire n697bar;
  wire n698bar;
  wire n699bar;
  wire n700bar;
  wire n701bar;
  wire n702bar;
  wire n703bar;
  wire n704bar;
  wire n705bar;
  wire n706bar;
  wire n707bar;
  wire n708bar;
  wire n709bar;
  wire n710bar;
  wire n711bar;
  wire n712bar;
  wire n713bar;
  wire n714bar;
  wire n715bar;
  wire n716bar;
  wire n717bar;
  wire n718bar;
  wire n719bar;
  wire n720bar;
  wire n721bar;
  wire n722bar;
  wire n723bar;
  wire n724bar;
  wire n725bar;
  wire n726bar;
  wire n727bar;
  wire n728bar;
  wire n729bar;
  wire n730bar;
  wire n731bar;
  wire n732bar;
  wire n733bar;
  wire n734bar;
  wire n735bar;
  wire n736bar;
  wire n737bar;
  wire n738bar;
  wire n739bar;
  wire n740bar;
  wire n741bar;
  wire n742bar;
  wire n743bar;
  wire n744bar;
  wire n745bar;
  wire n746bar;
  wire n747bar;
  wire n748bar;
  wire n749bar;
  wire n750bar;
  wire n751bar;
  wire n752bar;
  wire n753bar;
  wire n754bar;
  wire n755bar;
  wire n756bar;
  wire n757bar;
  wire n758bar;
  wire n759bar;
  wire n760bar;
  wire n761bar;
  wire n762bar;
  wire n763bar;
  wire n764bar;
  wire n765bar;
  wire n766bar;
  wire n767bar;
  wire n768bar;
  wire n769bar;
  wire n770bar;
  wire n771bar;
  wire n772bar;
  wire n773bar;
  wire n774bar;
  wire n775bar;
  wire n776bar;
  wire n777bar;
  wire n778bar;
  wire n779bar;
  wire n780bar;
  wire n781bar;
  wire n782bar;
  wire n783bar;
  wire n784bar;
  wire n785bar;
  wire n786bar;
  wire n787bar;
  wire n788bar;
  wire n789bar;
  wire n790bar;
  wire n791bar;
  wire n792bar;
  wire n793bar;
  wire n794bar;
  wire n795bar;
  wire n796bar;
  wire n797bar;
  wire n798bar;
  wire n799bar;
  wire n800bar;
  wire n801bar;
  wire n802bar;
  wire n803bar;
  wire n804bar;
  wire n805bar;
  wire n806bar;
  wire n807bar;
  wire n808bar;
  wire n809bar;
  wire n810bar;
  wire n811bar;
  wire n812bar;
  wire n813bar;
  wire n814bar;
  wire n815bar;
  wire n816bar;
  wire n817bar;
  wire n818bar;
  wire n819bar;
  wire n820bar;
  wire n821bar;
  wire n822bar;
  wire n823bar;
  wire n824bar;
  wire n825bar;
  wire n826bar;
  wire n827bar;
  wire n828bar;
  wire n829bar;
  wire n830bar;
  wire n831bar;
  wire n832bar;
  wire n833bar;
  wire n834bar;
  wire n835bar;
  wire n836bar;
  wire n837bar;
  wire n838bar;
  wire n839bar;
  wire n840bar;
  wire n841bar;
  wire n842bar;
  wire n843bar;
  wire n844bar;
  wire n845bar;
  wire n846bar;
  wire n847bar;
  wire n848bar;
  wire n849bar;
  wire n850bar;
  wire n851bar;
  wire n852bar;
  wire n853bar;
  wire n854bar;
  wire n855bar;
  wire n856bar;
  wire n857bar;
  wire n858bar;
  wire n859bar;
  wire n860bar;
  wire n861bar;
  wire n862bar;
  wire n863bar;
  wire n864bar;
  wire n865bar;
  wire n866bar;
  wire n867bar;
  wire n868bar;
  wire n869bar;
  wire n870bar;
  wire n871bar;
  wire n872bar;
  wire n873bar;
  wire n874bar;
  wire n875bar;
  wire n876bar;
  wire n877bar;
  wire n878bar;
  wire n879bar;
  wire n880bar;
  wire n881bar;
  wire n882bar;
  wire n883bar;
  wire n884bar;
  wire n885bar;
  wire n886bar;
  wire n887bar;
  wire n888bar;
  wire n889bar;
  wire n890bar;
  wire n891bar;
  wire n892bar;
  wire n893bar;
  wire n894bar;
  wire n895bar;
  wire n896bar;
  wire n897bar;
  wire n898bar;
  wire n899bar;
  wire n900bar;
  wire n901bar;
  wire n902bar;
  wire n903bar;
  wire n904bar;
  wire n905bar;
  wire n906bar;
  wire n907bar;
  wire n908bar;
  wire n909bar;
  wire n910bar;
  wire n911bar;
  wire n912bar;
  wire n913bar;
  wire n914bar;
  wire n915bar;
  wire n916bar;
  wire n917bar;
  wire n918bar;
  wire n919bar;
  wire n920bar;
  wire n921bar;
  wire n922bar;
  wire n923bar;
  wire n924bar;
  wire n925bar;
  wire n926bar;
  wire n927bar;
  wire n928bar;
  wire n929bar;
  wire n930bar;
  wire n931bar;
  wire n932bar;
  wire n933bar;
  wire n934bar;
  wire n935bar;
  wire n936bar;
  wire n937bar;
  wire n938bar;
  wire n939bar;
  wire n940bar;
  wire n941bar;
  wire n942bar;
  wire n943bar;
  wire n944bar;
  wire n945bar;
  wire n946bar;
  wire n947bar;
  wire n948bar;
  wire n949bar;
  wire n950bar;
  wire n951bar;
  wire n952bar;
  wire n953bar;
  wire n954bar;
  wire n955bar;
  wire n956bar;
  wire n957bar;
  wire n958bar;
  wire n959bar;
  wire n960bar;
  wire n961bar;
  wire n962bar;
  wire n963bar;
  wire n964bar;
  wire n965bar;
  wire n966bar;
  wire n967bar;
  wire n968bar;
  wire n969bar;
  wire n970bar;
  wire n971bar;
  wire n972bar;
//wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];
  //OR U1
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1 (
    .O(out[7]),
    .I0(n972),
    .I1(n971)
  );
  //AND U1bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1bar (
    .O(outbar[7]),
    .I0(n972bar),
    .I1(n971bar)
  );
  //OR U2
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2 (
    .O(n971),
    .I0(n970),
    .I1(n969)
  );
  //AND U2bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2bar (
    .O(n971bar),
    .I0(n970bar),
    .I1(n969bar)
  );
  //OR U3
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3 (
    .O(n969),
    .I0(n968),
    .I1(n967)
  );
  //AND U3bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3bar (
    .O(n969bar),
    .I0(n968bar),
    .I1(n967bar)
  );
  //OR U4
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4 (
    .O(n967),
    .I0(n966),
    .I1(n965)
  );
  //AND U4bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4bar (
    .O(n967bar),
    .I0(n966bar),
    .I1(n965bar)
  );
  //OR U5
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5 (
    .O(n968),
    .I0(n964),
    .I1(n963)
  );
  //AND U5bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5bar (
    .O(n968bar),
    .I0(n964bar),
    .I1(n963bar)
  );
  //OR U6
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6 (
    .O(n963),
    .I0(in[116]),
    .I1(n962)
  );
  //AND U6bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6bar (
    .O(n963bar),
    .I0(inbar[116]),
    .I1(n962bar)
  );
  //OR U7
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7 (
    .O(n970),
    .I0(n961),
    .I1(n960)
  );
  //AND U7bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7bar (
    .O(n970bar),
    .I0(n961bar),
    .I1(n960bar)
  );
  //OR U8
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8 (
    .O(n960),
    .I0(in[150]),
    .I1(in[127])
  );
  //AND U8bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8bar (
    .O(n960bar),
    .I0(inbar[150]),
    .I1(inbar[127])
  );
  //OR U9
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9 (
    .O(n961),
    .I0(in[160]),
    .I1(n959)
  );
  //AND U9bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9bar (
    .O(n961bar),
    .I0(inbar[160]),
    .I1(n959bar)
  );
  //OR U10
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10 (
    .O(n959),
    .I0(in[252]),
    .I1(in[168])
  );
  //AND U10bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10bar (
    .O(n959bar),
    .I0(inbar[252]),
    .I1(inbar[168])
  );
  //OR U11
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11 (
    .O(n972),
    .I0(n958),
    .I1(n957)
  );
  //AND U11bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11bar (
    .O(n972bar),
    .I0(n958bar),
    .I1(n957bar)
  );
  //OR U12
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12 (
    .O(n957),
    .I0(n956),
    .I1(n955)
  );
  //AND U12bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12bar (
    .O(n957bar),
    .I0(n956bar),
    .I1(n955bar)
  );
  //OR U13
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13 (
    .O(n955),
    .I0(in_17),
    .I1(in[96])
  );
  //AND U13bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13bar (
    .O(n955bar),
    .I0(in_17bar),
    .I1(inbar[96])
  );
  //OR U14
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14 (
    .O(n956),
    .I0(in_23),
    .I1(n954)
  );
  //AND U14bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14bar (
    .O(n956bar),
    .I0(in_23bar),
    .I1(n954bar)
  );
  //OR U15
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15 (
    .O(n954),
    .I0(in_31),
    .I1(in_26)
  );
  //AND U15bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15bar (
    .O(n954bar),
    .I0(in_31bar),
    .I1(in_26bar)
  );
  //OR U16
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16 (
    .O(n958),
    .I0(n953),
    .I1(n952)
  );
  //AND U16bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16bar (
    .O(n958bar),
    .I0(n953bar),
    .I1(n952bar)
  );
  //OR U17
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U17 (
    .O(n952),
    .I0(in_58),
    .I1(in_4)
  );
  //AND U17bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U17bar (
    .O(n952bar),
    .I0(in_58bar),
    .I1(in_4bar)
  );
  //OR U18
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U18 (
    .O(n953),
    .I0(in_59),
    .I1(n951)
  );
  //AND U18bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U18bar (
    .O(n953bar),
    .I0(in_59bar),
    .I1(n951bar)
  );
  //OR U19
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U19 (
    .O(n951),
    .I0(in_71),
    .I1(in_62)
  );
  //AND U19bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U19bar (
    .O(n951bar),
    .I0(in_71bar),
    .I1(in_62bar)
  );
  //OR U20
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U20 (
    .O(out[6]),
    .I0(n950),
    .I1(n949)
  );
  //AND U20bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U20bar (
    .O(outbar[6]),
    .I0(n950bar),
    .I1(n949bar)
  );
  //OR U21
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U21 (
    .O(n949),
    .I0(n948),
    .I1(n947)
  );
  //AND U21bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U21bar (
    .O(n949bar),
    .I0(n948bar),
    .I1(n947bar)
  );
  //OR U22
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U22 (
    .O(n947),
    .I0(n946),
    .I1(n945)
  );
  //AND U22bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U22bar (
    .O(n947bar),
    .I0(n946bar),
    .I1(n945bar)
  );
  //OR U23
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U23 (
    .O(n945),
    .I0(n944),
    .I1(n943)
  );
  //AND U23bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U23bar (
    .O(n945bar),
    .I0(n944bar),
    .I1(n943bar)
  );
  //OR U24
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U24 (
    .O(n946),
    .I0(n942),
    .I1(n941)
  );
  //AND U24bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U24bar (
    .O(n946bar),
    .I0(n942bar),
    .I1(n941bar)
  );
  //OR U25
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U25 (
    .O(n941),
    .I0(in[101]),
    .I1(n940)
  );
  //AND U25bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U25bar (
    .O(n941bar),
    .I0(inbar[101]),
    .I1(n940bar)
  );
  //OR U26
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U26 (
    .O(n948),
    .I0(n939),
    .I1(n938)
  );
  //AND U26bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U26bar (
    .O(n948bar),
    .I0(n939bar),
    .I1(n938bar)
  );
  //OR U27
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U27 (
    .O(n938),
    .I0(in[114]),
    .I1(in[104])
  );
  //AND U27bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U27bar (
    .O(n938bar),
    .I0(inbar[114]),
    .I1(inbar[104])
  );
  //OR U28
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U28 (
    .O(n939),
    .I0(in[128]),
    .I1(n937)
  );
  //AND U28bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U28bar (
    .O(n939bar),
    .I0(inbar[128]),
    .I1(n937bar)
  );
  //OR U29
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U29 (
    .O(n937),
    .I0(in[136]),
    .I1(in[134])
  );
  //AND U29bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U29bar (
    .O(n937bar),
    .I0(inbar[136]),
    .I1(inbar[134])
  );
  //OR U30
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U30 (
    .O(n950),
    .I0(n936),
    .I1(n935)
  );
  //AND U30bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U30bar (
    .O(n950bar),
    .I0(n936bar),
    .I1(n935bar)
  );
  //OR U31
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U31 (
    .O(n935),
    .I0(n934),
    .I1(n933)
  );
  //AND U31bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U31bar (
    .O(n935bar),
    .I0(n934bar),
    .I1(n933bar)
  );
  //OR U32
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U32 (
    .O(n933),
    .I0(in[177]),
    .I1(in[164])
  );
  //AND U32bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U32bar (
    .O(n933bar),
    .I0(inbar[177]),
    .I1(inbar[164])
  );
  //OR U33
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U33 (
    .O(n934),
    .I0(in[212]),
    .I1(n932)
  );
  //AND U33bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U33bar (
    .O(n934bar),
    .I0(inbar[212]),
    .I1(n932bar)
  );
  //OR U34
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U34 (
    .O(n932),
    .I0(in[248]),
    .I1(in[221])
  );
  //AND U34bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U34bar (
    .O(n932bar),
    .I0(inbar[248]),
    .I1(inbar[221])
  );
  //OR U35
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U35 (
    .O(n936),
    .I0(n931),
    .I1(n930)
  );
  //AND U35bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U35bar (
    .O(n936bar),
    .I0(n931bar),
    .I1(n930bar)
  );
  //OR U36
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U36 (
    .O(n930),
    .I0(in_18),
    .I1(in[93])
  );
  //AND U36bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U36bar (
    .O(n930bar),
    .I0(in_18bar),
    .I1(inbar[93])
  );
  //OR U37
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U37 (
    .O(n931),
    .I0(in_31),
    .I1(n929)
  );
  //AND U37bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U37bar (
    .O(n931bar),
    .I0(in_31bar),
    .I1(n929bar)
  );
  //OR U38
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U38 (
    .O(n929),
    .I0(in_7),
    .I1(in_39)
  );
  //AND U38bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U38bar (
    .O(n929bar),
    .I0(in_7bar),
    .I1(in_39bar)
  );
  //OR U39
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U39 (
    .O(out[5]),
    .I0(n928),
    .I1(n927)
  );
  //AND U39bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U39bar (
    .O(outbar[5]),
    .I0(n928bar),
    .I1(n927bar)
  );
  //OR U40
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U40 (
    .O(n927),
    .I0(n926),
    .I1(n925)
  );
  //AND U40bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U40bar (
    .O(n927bar),
    .I0(n926bar),
    .I1(n925bar)
  );
  //OR U41
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U41 (
    .O(n925),
    .I0(n924),
    .I1(n923)
  );
  //AND U41bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U41bar (
    .O(n925bar),
    .I0(n924bar),
    .I1(n923bar)
  );
  //OR U42
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U42 (
    .O(n923),
    .I0(n922),
    .I1(n921)
  );
  //AND U42bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U42bar (
    .O(n923bar),
    .I0(n922bar),
    .I1(n921bar)
  );
  //OR U43
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U43 (
    .O(n924),
    .I0(n940),
    .I1(n920)
  );
  //AND U43bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U43bar (
    .O(n924bar),
    .I0(n940bar),
    .I1(n920bar)
  );
  //OR U44
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U44 (
    .O(n920),
    .I0(in[111]),
    .I1(n919)
  );
  //AND U44bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U44bar (
    .O(n920bar),
    .I0(inbar[111]),
    .I1(n919bar)
  );
  //OR U45
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U45 (
    .O(n940),
    .I0(n918),
    .I1(n917)
  );
  //AND U45bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U45bar (
    .O(n940bar),
    .I0(n918bar),
    .I1(n917bar)
  );
  //OR U46
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U46 (
    .O(n917),
    .I0(n916),
    .I1(n915)
  );
  //AND U46bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U46bar (
    .O(n917bar),
    .I0(n916bar),
    .I1(n915bar)
  );
  //OR U47
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U47 (
    .O(n915),
    .I0(n914),
    .I1(n913)
  );
  //AND U47bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U47bar (
    .O(n915bar),
    .I0(n914bar),
    .I1(n913bar)
  );
  //OR U48
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U48 (
    .O(n913),
    .I0(in[140]),
    .I1(in[131])
  );
  //AND U48bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U48bar (
    .O(n913bar),
    .I0(inbar[140]),
    .I1(inbar[131])
  );
  //OR U49
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U49 (
    .O(n914),
    .I0(in[160]),
    .I1(in[144])
  );
  //AND U49bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U49bar (
    .O(n914bar),
    .I0(inbar[160]),
    .I1(inbar[144])
  );
  //OR U50
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U50 (
    .O(n916),
    .I0(n912),
    .I1(n911)
  );
  //AND U50bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U50bar (
    .O(n916bar),
    .I0(n912bar),
    .I1(n911bar)
  );
  //OR U51
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U51 (
    .O(n911),
    .I0(in[179]),
    .I1(in[174])
  );
  //AND U51bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U51bar (
    .O(n911bar),
    .I0(inbar[179]),
    .I1(inbar[174])
  );
  //OR U52
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U52 (
    .O(n912),
    .I0(in[188]),
    .I1(in[184])
  );
  //AND U52bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U52bar (
    .O(n912bar),
    .I0(inbar[188]),
    .I1(inbar[184])
  );
  //OR U53
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U53 (
    .O(n918),
    .I0(n910),
    .I1(n909)
  );
  //AND U53bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U53bar (
    .O(n918bar),
    .I0(n910bar),
    .I1(n909bar)
  );
  //OR U54
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U54 (
    .O(n909),
    .I0(n908),
    .I1(n907)
  );
  //AND U54bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U54bar (
    .O(n909bar),
    .I0(n908bar),
    .I1(n907bar)
  );
  //OR U55
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U55 (
    .O(n907),
    .I0(in[216]),
    .I1(in[200])
  );
  //AND U55bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U55bar (
    .O(n907bar),
    .I0(inbar[216]),
    .I1(inbar[200])
  );
  //OR U56
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U56 (
    .O(n908),
    .I0(in[228]),
    .I1(in[224])
  );
  //AND U56bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U56bar (
    .O(n908bar),
    .I0(inbar[228]),
    .I1(inbar[224])
  );
  //OR U57
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U57 (
    .O(n910),
    .I0(n906),
    .I1(n905)
  );
  //AND U57bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U57bar (
    .O(n910bar),
    .I0(n906bar),
    .I1(n905bar)
  );
  //OR U58
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U58 (
    .O(n905),
    .I0(in[247]),
    .I1(in[235])
  );
  //AND U58bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U58bar (
    .O(n905bar),
    .I0(inbar[247]),
    .I1(inbar[235])
  );
  //OR U59
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U59 (
    .O(n906),
    .I0(in_42),
    .I1(in[83])
  );
  //AND U59bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U59bar (
    .O(n906bar),
    .I0(in_42bar),
    .I1(inbar[83])
  );
  //OR U60
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U60 (
    .O(n926),
    .I0(n904),
    .I1(n903)
  );
  //AND U60bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U60bar (
    .O(n926bar),
    .I0(n904bar),
    .I1(n903bar)
  );
  //OR U61
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U61 (
    .O(n903),
    .I0(in[166]),
    .I1(in[123])
  );
  //AND U61bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U61bar (
    .O(n903bar),
    .I0(inbar[166]),
    .I1(inbar[123])
  );
  //OR U62
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U62 (
    .O(n904),
    .I0(in[170]),
    .I1(n902)
  );
  //AND U62bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U62bar (
    .O(n904bar),
    .I0(inbar[170]),
    .I1(n902bar)
  );
  //OR U63
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U63 (
    .O(n902),
    .I0(in[194]),
    .I1(in[183])
  );
  //AND U63bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U63bar (
    .O(n902bar),
    .I0(inbar[194]),
    .I1(inbar[183])
  );
  //OR U64
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U64 (
    .O(n928),
    .I0(n901),
    .I1(n900)
  );
  //AND U64bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U64bar (
    .O(n928bar),
    .I0(n901bar),
    .I1(n900bar)
  );
  //OR U65
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U65 (
    .O(n900),
    .I0(n899),
    .I1(n898)
  );
  //AND U65bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U65bar (
    .O(n900bar),
    .I0(n899bar),
    .I1(n898bar)
  );
  //OR U66
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U66 (
    .O(n898),
    .I0(in[241]),
    .I1(in[238])
  );
  //AND U66bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U66bar (
    .O(n898bar),
    .I0(inbar[241]),
    .I1(inbar[238])
  );
  //OR U67
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U67 (
    .O(n899),
    .I0(in[250]),
    .I1(n897)
  );
  //AND U67bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U67bar (
    .O(n899bar),
    .I0(inbar[250]),
    .I1(n897bar)
  );
  //OR U68
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U68 (
    .O(n897),
    .I0(in_24),
    .I1(in[84])
  );
  //AND U68bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U68bar (
    .O(n897bar),
    .I0(in_24bar),
    .I1(inbar[84])
  );
  //OR U69
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U69 (
    .O(n901),
    .I0(n896),
    .I1(n895)
  );
  //AND U69bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U69bar (
    .O(n901bar),
    .I0(n896bar),
    .I1(n895bar)
  );
  //OR U70
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U70 (
    .O(n895),
    .I0(in_41),
    .I1(in_29)
  );
  //AND U70bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U70bar (
    .O(n895bar),
    .I0(in_41bar),
    .I1(in_29bar)
  );
  //OR U71
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U71 (
    .O(n896),
    .I0(in_66),
    .I1(n894)
  );
  //AND U71bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U71bar (
    .O(n896bar),
    .I0(in_66bar),
    .I1(n894bar)
  );
  //OR U72
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U72 (
    .O(n894),
    .I0(in_76),
    .I1(in_71)
  );
  //AND U72bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U72bar (
    .O(n894bar),
    .I0(in_76bar),
    .I1(in_71bar)
  );
  //OR U73
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U73 (
    .O(out[4]),
    .I0(n893),
    .I1(n892)
  );
  //AND U73bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U73bar (
    .O(outbar[4]),
    .I0(n893bar),
    .I1(n892bar)
  );
  //OR U74
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U74 (
    .O(n892),
    .I0(n891),
    .I1(n890)
  );
  //AND U74bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U74bar (
    .O(n892bar),
    .I0(n891bar),
    .I1(n890bar)
  );
  //OR U75
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U75 (
    .O(n890),
    .I0(n889),
    .I1(n888)
  );
  //AND U75bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U75bar (
    .O(n890bar),
    .I0(n889bar),
    .I1(n888bar)
  );
  //OR U76
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U76 (
    .O(n888),
    .I0(n922),
    .I1(n887)
  );
  //AND U76bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U76bar (
    .O(n888bar),
    .I0(n922bar),
    .I1(n887bar)
  );
  //OR U77
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U77 (
    .O(n922),
    .I0(n886),
    .I1(n885)
  );
  //AND U77bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U77bar (
    .O(n922bar),
    .I0(n886bar),
    .I1(n885bar)
  );
  //OR U78
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U78 (
    .O(n885),
    .I0(n884),
    .I1(n883)
  );
  //AND U78bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U78bar (
    .O(n885bar),
    .I0(n884bar),
    .I1(n883bar)
  );
  //OR U79
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U79 (
    .O(n883),
    .I0(n882),
    .I1(n881)
  );
  //AND U79bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U79bar (
    .O(n883bar),
    .I0(n882bar),
    .I1(n881bar)
  );
  //OR U80
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U80 (
    .O(n881),
    .I0(in[118]),
    .I1(in[109])
  );
  //AND U80bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U80bar (
    .O(n881bar),
    .I0(inbar[118]),
    .I1(inbar[109])
  );
  //OR U81
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U81 (
    .O(n882),
    .I0(in[139]),
    .I1(in[120])
  );
  //AND U81bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U81bar (
    .O(n882bar),
    .I0(inbar[139]),
    .I1(inbar[120])
  );
  //OR U82
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U82 (
    .O(n884),
    .I0(n880),
    .I1(n879)
  );
  //AND U82bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U82bar (
    .O(n884bar),
    .I0(n880bar),
    .I1(n879bar)
  );
  //OR U83
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U83 (
    .O(n879),
    .I0(in[198]),
    .I1(in[154])
  );
  //AND U83bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U83bar (
    .O(n879bar),
    .I0(inbar[198]),
    .I1(inbar[154])
  );
  //OR U84
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U84 (
    .O(n880),
    .I0(in[210]),
    .I1(in[205])
  );
  //AND U84bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U84bar (
    .O(n880bar),
    .I0(inbar[210]),
    .I1(inbar[205])
  );
  //OR U85
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U85 (
    .O(n886),
    .I0(n878),
    .I1(n877)
  );
  //AND U85bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U85bar (
    .O(n886bar),
    .I0(n878bar),
    .I1(n877bar)
  );
  //OR U86
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U86 (
    .O(n877),
    .I0(n876),
    .I1(n875)
  );
  //AND U86bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U86bar (
    .O(n877bar),
    .I0(n876bar),
    .I1(n875bar)
  );
  //OR U87
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U87 (
    .O(n875),
    .I0(in[219]),
    .I1(in[217])
  );
  //AND U87bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U87bar (
    .O(n875bar),
    .I0(inbar[219]),
    .I1(inbar[217])
  );
  //OR U88
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U88 (
    .O(n876),
    .I0(in[86]),
    .I1(in[252])
  );
  //AND U88bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U88bar (
    .O(n876bar),
    .I0(inbar[86]),
    .I1(inbar[252])
  );
  //OR U89
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U89 (
    .O(n878),
    .I0(n874),
    .I1(n873)
  );
  //AND U89bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U89bar (
    .O(n878bar),
    .I0(n874bar),
    .I1(n873bar)
  );
  //OR U90
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U90 (
    .O(n873),
    .I0(in_40),
    .I1(in[91])
  );
  //AND U90bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U90bar (
    .O(n873bar),
    .I0(in_40bar),
    .I1(inbar[91])
  );
  //OR U91
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U91 (
    .O(n874),
    .I0(in_8),
    .I1(in_46)
  );
  //AND U91bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U91bar (
    .O(n874bar),
    .I0(in_8bar),
    .I1(in_46bar)
  );
  //OR U92
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U92 (
    .O(n889),
    .I0(n872),
    .I1(n871)
  );
  //AND U92bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U92bar (
    .O(n889bar),
    .I0(n872bar),
    .I1(n871bar)
  );
  //OR U93
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U93 (
    .O(n871),
    .I0(in[117]),
    .I1(n943)
  );
  //AND U93bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U93bar (
    .O(n871bar),
    .I0(inbar[117]),
    .I1(n943bar)
  );
  //OR U94
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U94 (
    .O(n943),
    .I0(n870),
    .I1(n869)
  );
  //AND U94bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U94bar (
    .O(n943bar),
    .I0(n870bar),
    .I1(n869bar)
  );
  //OR U95
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U95 (
    .O(n869),
    .I0(n868),
    .I1(n867)
  );
  //AND U95bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U95bar (
    .O(n869bar),
    .I0(n868bar),
    .I1(n867bar)
  );
  //OR U96
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U96 (
    .O(n867),
    .I0(n866),
    .I1(n865)
  );
  //AND U96bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U96bar (
    .O(n867bar),
    .I0(n866bar),
    .I1(n865bar)
  );
  //OR U97
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U97 (
    .O(n865),
    .I0(n864),
    .I1(n863)
  );
  //AND U97bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U97bar (
    .O(n865bar),
    .I0(n864bar),
    .I1(n863bar)
  );
  //OR U98
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U98 (
    .O(n866),
    .I0(in[108]),
    .I1(n919)
  );
  //AND U98bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U98bar (
    .O(n866bar),
    .I0(inbar[108]),
    .I1(n919bar)
  );
  //OR U99
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U99 (
    .O(n919),
    .I0(n862),
    .I1(n861)
  );
  //AND U99bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U99bar (
    .O(n919bar),
    .I0(n862bar),
    .I1(n861bar)
  );
  //OR U100
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U100 (
    .O(n861),
    .I0(n860),
    .I1(n859)
  );
  //AND U100bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U100bar (
    .O(n861bar),
    .I0(n860bar),
    .I1(n859bar)
  );
  //OR U101
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U101 (
    .O(n859),
    .I0(n858),
    .I1(n857)
  );
  //AND U101bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U101bar (
    .O(n859bar),
    .I0(n858bar),
    .I1(n857bar)
  );
  //OR U102
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U102 (
    .O(n857),
    .I0(in[119]),
    .I1(in[105])
  );
  //AND U102bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U102bar (
    .O(n857bar),
    .I0(inbar[119]),
    .I1(inbar[105])
  );
  //OR U103
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U103 (
    .O(n858),
    .I0(in[186]),
    .I1(in[175])
  );
  //AND U103bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U103bar (
    .O(n858bar),
    .I0(inbar[186]),
    .I1(inbar[175])
  );
  //OR U104
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U104 (
    .O(n860),
    .I0(n856),
    .I1(n855)
  );
  //AND U104bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U104bar (
    .O(n860bar),
    .I0(n856bar),
    .I1(n855bar)
  );
  //OR U105
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U105 (
    .O(n855),
    .I0(in[202]),
    .I1(in[193])
  );
  //AND U105bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U105bar (
    .O(n855bar),
    .I0(inbar[202]),
    .I1(inbar[193])
  );
  //OR U106
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U106 (
    .O(n856),
    .I0(in[225]),
    .I1(in[208])
  );
  //AND U106bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U106bar (
    .O(n856bar),
    .I0(inbar[225]),
    .I1(inbar[208])
  );
  //OR U107
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U107 (
    .O(n862),
    .I0(n854),
    .I1(n853)
  );
  //AND U107bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U107bar (
    .O(n862bar),
    .I0(n854bar),
    .I1(n853bar)
  );
  //OR U108
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U108 (
    .O(n853),
    .I0(n852),
    .I1(n851)
  );
  //AND U108bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U108bar (
    .O(n853bar),
    .I0(n852bar),
    .I1(n851bar)
  );
  //OR U109
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U109 (
    .O(n851),
    .I0(in_1),
    .I1(in[85])
  );
  //AND U109bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U109bar (
    .O(n851bar),
    .I0(in_1bar),
    .I1(inbar[85])
  );
  //OR U110
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U110 (
    .O(n852),
    .I0(in_23),
    .I1(in_19)
  );
  //AND U110bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U110bar (
    .O(n852bar),
    .I0(in_23bar),
    .I1(in_19bar)
  );
  //OR U111
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U111 (
    .O(n854),
    .I0(n850),
    .I1(n849)
  );
  //AND U111bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U111bar (
    .O(n854bar),
    .I0(n850bar),
    .I1(n849bar)
  );
  //OR U112
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U112 (
    .O(n849),
    .I0(in_43),
    .I1(in_33)
  );
  //AND U112bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U112bar (
    .O(n849bar),
    .I0(in_43bar),
    .I1(in_33bar)
  );
  //OR U113
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U113 (
    .O(n850),
    .I0(in_63),
    .I1(in_44)
  );
  //AND U113bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U113bar (
    .O(n850bar),
    .I0(in_63bar),
    .I1(in_44bar)
  );
  //OR U114
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U114 (
    .O(n868),
    .I0(n848),
    .I1(n847)
  );
  //AND U114bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U114bar (
    .O(n868bar),
    .I0(n848bar),
    .I1(n847bar)
  );
  //OR U115
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U115 (
    .O(n847),
    .I0(in[141]),
    .I1(in[112])
  );
  //AND U115bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U115bar (
    .O(n847bar),
    .I0(inbar[141]),
    .I1(inbar[112])
  );
  //OR U116
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U116 (
    .O(n848),
    .I0(in[147]),
    .I1(n846)
  );
  //AND U116bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U116bar (
    .O(n848bar),
    .I0(inbar[147]),
    .I1(n846bar)
  );
  //OR U117
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U117 (
    .O(n846),
    .I0(in[181]),
    .I1(in[167])
  );
  //AND U117bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U117bar (
    .O(n846bar),
    .I0(inbar[181]),
    .I1(inbar[167])
  );
  //OR U118
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U118 (
    .O(n870),
    .I0(n845),
    .I1(n844)
  );
  //AND U118bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U118bar (
    .O(n870bar),
    .I0(n845bar),
    .I1(n844bar)
  );
  //OR U119
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U119 (
    .O(n844),
    .I0(n843),
    .I1(n842)
  );
  //AND U119bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U119bar (
    .O(n844bar),
    .I0(n843bar),
    .I1(n842bar)
  );
  //OR U120
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U120 (
    .O(n842),
    .I0(in[229]),
    .I1(in[201])
  );
  //AND U120bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U120bar (
    .O(n842bar),
    .I0(inbar[229]),
    .I1(inbar[201])
  );
  //OR U121
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U121 (
    .O(n843),
    .I0(in[237]),
    .I1(n841)
  );
  //AND U121bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U121bar (
    .O(n843bar),
    .I0(inbar[237]),
    .I1(n841bar)
  );
  //OR U122
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U122 (
    .O(n841),
    .I0(in[94]),
    .I1(in[253])
  );
  //AND U122bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U122bar (
    .O(n841bar),
    .I0(inbar[94]),
    .I1(inbar[253])
  );
  //OR U123
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U123 (
    .O(n845),
    .I0(n840),
    .I1(n839)
  );
  //AND U123bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U123bar (
    .O(n845bar),
    .I0(n840bar),
    .I1(n839bar)
  );
  //OR U124
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U124 (
    .O(n839),
    .I0(in_21),
    .I1(in[96])
  );
  //AND U124bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U124bar (
    .O(n839bar),
    .I0(in_21bar),
    .I1(inbar[96])
  );
  //OR U125
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U125 (
    .O(n840),
    .I0(in_25),
    .I1(n838)
  );
  //AND U125bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U125bar (
    .O(n840bar),
    .I0(in_25bar),
    .I1(n838bar)
  );
  //OR U126
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U126 (
    .O(n838),
    .I0(in_81),
    .I1(in_45)
  );
  //AND U126bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U126bar (
    .O(n838bar),
    .I0(in_81bar),
    .I1(in_45bar)
  );
  //OR U127
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U127 (
    .O(n891),
    .I0(n837),
    .I1(n836)
  );
  //AND U127bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U127bar (
    .O(n891bar),
    .I0(n837bar),
    .I1(n836bar)
  );
  //OR U128
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U128 (
    .O(n836),
    .I0(in[142]),
    .I1(in[124])
  );
  //AND U128bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U128bar (
    .O(n836bar),
    .I0(inbar[142]),
    .I1(inbar[124])
  );
  //OR U129
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U129 (
    .O(n837),
    .I0(in[150]),
    .I1(n835)
  );
  //AND U129bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U129bar (
    .O(n837bar),
    .I0(inbar[150]),
    .I1(n835bar)
  );
  //OR U130
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U130 (
    .O(n835),
    .I0(in[172]),
    .I1(in[155])
  );
  //AND U130bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U130bar (
    .O(n835bar),
    .I0(inbar[172]),
    .I1(inbar[155])
  );
  //OR U131
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U131 (
    .O(n893),
    .I0(n834),
    .I1(n833)
  );
  //AND U131bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U131bar (
    .O(n893bar),
    .I0(n834bar),
    .I1(n833bar)
  );
  //OR U132
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U132 (
    .O(n833),
    .I0(n832),
    .I1(n831)
  );
  //AND U132bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U132bar (
    .O(n833bar),
    .I0(n832bar),
    .I1(n831bar)
  );
  //OR U133
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U133 (
    .O(n831),
    .I0(in[196]),
    .I1(in[173])
  );
  //AND U133bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U133bar (
    .O(n831bar),
    .I0(inbar[196]),
    .I1(inbar[173])
  );
  //OR U134
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U134 (
    .O(n832),
    .I0(in[222]),
    .I1(n830)
  );
  //AND U134bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U134bar (
    .O(n832bar),
    .I0(inbar[222]),
    .I1(n830bar)
  );
  //OR U135
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U135 (
    .O(n830),
    .I0(in[227]),
    .I1(in[226])
  );
  //AND U135bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U135bar (
    .O(n830bar),
    .I0(inbar[227]),
    .I1(inbar[226])
  );
  //OR U136
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U136 (
    .O(n834),
    .I0(n829),
    .I1(n828)
  );
  //AND U136bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U136bar (
    .O(n834bar),
    .I0(n829bar),
    .I1(n828bar)
  );
  //OR U137
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U137 (
    .O(n828),
    .I0(in[249]),
    .I1(in[231])
  );
  //AND U137bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U137bar (
    .O(n828bar),
    .I0(inbar[249]),
    .I1(inbar[231])
  );
  //OR U138
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U138 (
    .O(n829),
    .I0(in_28),
    .I1(n827)
  );
  //AND U138bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U138bar (
    .O(n829bar),
    .I0(in_28bar),
    .I1(n827bar)
  );
  //OR U139
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U139 (
    .O(n827),
    .I0(in_52),
    .I1(in_47)
  );
  //AND U139bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U139bar (
    .O(n827bar),
    .I0(in_52bar),
    .I1(in_47bar)
  );
  //OR U140
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U140 (
    .O(out[3]),
    .I0(n826),
    .I1(n825)
  );
  //AND U140bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U140bar (
    .O(outbar[3]),
    .I0(n826bar),
    .I1(n825bar)
  );
  //OR U141
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U141 (
    .O(n825),
    .I0(n824),
    .I1(n823)
  );
  //AND U141bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U141bar (
    .O(n825bar),
    .I0(n824bar),
    .I1(n823bar)
  );
  //OR U142
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U142 (
    .O(n823),
    .I0(n822),
    .I1(n821)
  );
  //AND U142bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U142bar (
    .O(n823bar),
    .I0(n822bar),
    .I1(n821bar)
  );
  //OR U143
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U143 (
    .O(n821),
    .I0(n820),
    .I1(n819)
  );
  //AND U143bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U143bar (
    .O(n821bar),
    .I0(n820bar),
    .I1(n819bar)
  );
  //OR U144
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U144 (
    .O(n822),
    .I0(n964),
    .I1(n818)
  );
  //AND U144bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U144bar (
    .O(n822bar),
    .I0(n964bar),
    .I1(n818bar)
  );
  //OR U145
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U145 (
    .O(n818),
    .I0(in[118]),
    .I1(n817)
  );
  //AND U145bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U145bar (
    .O(n818bar),
    .I0(inbar[118]),
    .I1(n817bar)
  );
  //OR U146
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U146 (
    .O(n964),
    .I0(n816),
    .I1(n815)
  );
  //AND U146bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U146bar (
    .O(n964bar),
    .I0(n816bar),
    .I1(n815bar)
  );
  //OR U147
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U147 (
    .O(n815),
    .I0(n814),
    .I1(n813)
  );
  //AND U147bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U147bar (
    .O(n815bar),
    .I0(n814bar),
    .I1(n813bar)
  );
  //OR U148
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U148 (
    .O(n813),
    .I0(n812),
    .I1(n811)
  );
  //AND U148bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U148bar (
    .O(n813bar),
    .I0(n812bar),
    .I1(n811bar)
  );
  //OR U149
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U149 (
    .O(n811),
    .I0(in[122]),
    .I1(in[111])
  );
  //AND U149bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U149bar (
    .O(n811bar),
    .I0(inbar[122]),
    .I1(inbar[111])
  );
  //OR U150
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U150 (
    .O(n812),
    .I0(in[154]),
    .I1(in[151])
  );
  //AND U150bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U150bar (
    .O(n812bar),
    .I0(inbar[154]),
    .I1(inbar[151])
  );
  //OR U151
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U151 (
    .O(n814),
    .I0(n810),
    .I1(n809)
  );
  //AND U151bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U151bar (
    .O(n814bar),
    .I0(n810bar),
    .I1(n809bar)
  );
  //OR U152
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U152 (
    .O(n809),
    .I0(in[187]),
    .I1(in[177])
  );
  //AND U152bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U152bar (
    .O(n809bar),
    .I0(inbar[187]),
    .I1(inbar[177])
  );
  //OR U153
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U153 (
    .O(n810),
    .I0(in[200]),
    .I1(in[192])
  );
  //AND U153bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U153bar (
    .O(n810bar),
    .I0(inbar[200]),
    .I1(inbar[192])
  );
  //OR U154
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U154 (
    .O(n816),
    .I0(n808),
    .I1(n807)
  );
  //AND U154bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U154bar (
    .O(n816bar),
    .I0(n808bar),
    .I1(n807bar)
  );
  //OR U155
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U155 (
    .O(n807),
    .I0(n806),
    .I1(n805)
  );
  //AND U155bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U155bar (
    .O(n807bar),
    .I0(n806bar),
    .I1(n805bar)
  );
  //OR U156
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U156 (
    .O(n805),
    .I0(in[225]),
    .I1(in[207])
  );
  //AND U156bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U156bar (
    .O(n805bar),
    .I0(inbar[225]),
    .I1(inbar[207])
  );
  //OR U157
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U157 (
    .O(n806),
    .I0(in[98]),
    .I1(in[226])
  );
  //AND U157bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U157bar (
    .O(n806bar),
    .I0(inbar[98]),
    .I1(inbar[226])
  );
  //OR U158
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U158 (
    .O(n808),
    .I0(n804),
    .I1(n803)
  );
  //AND U158bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U158bar (
    .O(n808bar),
    .I0(n804bar),
    .I1(n803bar)
  );
  //OR U159
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U159 (
    .O(n803),
    .I0(in_20),
    .I1(in_16)
  );
  //AND U159bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U159bar (
    .O(n803bar),
    .I0(in_20bar),
    .I1(in_16bar)
  );
  //OR U160
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U160 (
    .O(n804),
    .I0(in_55),
    .I1(in_45)
  );
  //AND U160bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U160bar (
    .O(n804bar),
    .I0(in_55bar),
    .I1(in_45bar)
  );
  //OR U161
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U161 (
    .O(n824),
    .I0(n802),
    .I1(n801)
  );
  //AND U161bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U161bar (
    .O(n824bar),
    .I0(n802bar),
    .I1(n801bar)
  );
  //OR U162
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U162 (
    .O(n801),
    .I0(in[162]),
    .I1(in[149])
  );
  //AND U162bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U162bar (
    .O(n801bar),
    .I0(inbar[162]),
    .I1(inbar[149])
  );
  //OR U163
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U163 (
    .O(n802),
    .I0(in[163]),
    .I1(n800)
  );
  //AND U163bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U163bar (
    .O(n802bar),
    .I0(inbar[163]),
    .I1(n800bar)
  );
  //OR U164
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U164 (
    .O(n800),
    .I0(in[191]),
    .I1(in[189])
  );
  //AND U164bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U164bar (
    .O(n800bar),
    .I0(inbar[191]),
    .I1(inbar[189])
  );
  //OR U165
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U165 (
    .O(n826),
    .I0(n799),
    .I1(n798)
  );
  //AND U165bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U165bar (
    .O(n826bar),
    .I0(n799bar),
    .I1(n798bar)
  );
  //OR U166
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U166 (
    .O(n798),
    .I0(n797),
    .I1(n796)
  );
  //AND U166bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U166bar (
    .O(n798bar),
    .I0(n797bar),
    .I1(n796bar)
  );
  //OR U167
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U167 (
    .O(n796),
    .I0(in[212]),
    .I1(in[193])
  );
  //AND U167bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U167bar (
    .O(n796bar),
    .I0(inbar[212]),
    .I1(inbar[193])
  );
  //OR U168
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U168 (
    .O(n797),
    .I0(in[238]),
    .I1(n795)
  );
  //AND U168bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U168bar (
    .O(n797bar),
    .I0(inbar[238]),
    .I1(n795bar)
  );
  //OR U169
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U169 (
    .O(n795),
    .I0(in[88]),
    .I1(in[247])
  );
  //AND U169bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U169bar (
    .O(n795bar),
    .I0(inbar[88]),
    .I1(inbar[247])
  );
  //OR U170
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U170 (
    .O(n799),
    .I0(n794),
    .I1(n793)
  );
  //AND U170bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U170bar (
    .O(n799bar),
    .I0(n794bar),
    .I1(n793bar)
  );
  //OR U171
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U171 (
    .O(n793),
    .I0(in[94]),
    .I1(in[92])
  );
  //AND U171bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U171bar (
    .O(n793bar),
    .I0(inbar[94]),
    .I1(inbar[92])
  );
  //OR U172
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U172 (
    .O(n794),
    .I0(in_52),
    .I1(n792)
  );
  //AND U172bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U172bar (
    .O(n794bar),
    .I0(in_52bar),
    .I1(n792bar)
  );
  //OR U173
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U173 (
    .O(n792),
    .I0(in_70),
    .I1(in_67)
  );
  //AND U173bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U173bar (
    .O(n792bar),
    .I0(in_70bar),
    .I1(in_67bar)
  );
  //OR U174
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U174 (
    .O(out[2]),
    .I0(n791),
    .I1(n790)
  );
  //AND U174bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U174bar (
    .O(outbar[2]),
    .I0(n791bar),
    .I1(n790bar)
  );
  //OR U175
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U175 (
    .O(n790),
    .I0(n789),
    .I1(n788)
  );
  //AND U175bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U175bar (
    .O(n790bar),
    .I0(n789bar),
    .I1(n788bar)
  );
  //OR U176
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U176 (
    .O(n788),
    .I0(n787),
    .I1(n786)
  );
  //AND U176bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U176bar (
    .O(n788bar),
    .I0(n787bar),
    .I1(n786bar)
  );
  //OR U177
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U177 (
    .O(n786),
    .I0(n819),
    .I1(n785)
  );
  //AND U177bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U177bar (
    .O(n786bar),
    .I0(n819bar),
    .I1(n785bar)
  );
  //OR U178
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U178 (
    .O(n819),
    .I0(n784),
    .I1(n783)
  );
  //AND U178bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U178bar (
    .O(n819bar),
    .I0(n784bar),
    .I1(n783bar)
  );
  //OR U179
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U179 (
    .O(n783),
    .I0(n782),
    .I1(n781)
  );
  //AND U179bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U179bar (
    .O(n783bar),
    .I0(n782bar),
    .I1(n781bar)
  );
  //OR U180
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U180 (
    .O(n781),
    .I0(n780),
    .I1(n779)
  );
  //AND U180bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U180bar (
    .O(n781bar),
    .I0(n780bar),
    .I1(n779bar)
  );
  //OR U181
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U181 (
    .O(n779),
    .I0(n962),
    .I1(n778)
  );
  //AND U181bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U181bar (
    .O(n779bar),
    .I0(n962bar),
    .I1(n778bar)
  );
  //OR U182
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U182 (
    .O(n962),
    .I0(n777),
    .I1(n776)
  );
  //AND U182bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U182bar (
    .O(n962bar),
    .I0(n777bar),
    .I1(n776bar)
  );
  //OR U183
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U183 (
    .O(n776),
    .I0(n775),
    .I1(n774)
  );
  //AND U183bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U183bar (
    .O(n776bar),
    .I0(n775bar),
    .I1(n774bar)
  );
  //OR U184
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U184 (
    .O(n774),
    .I0(n773),
    .I1(n772)
  );
  //AND U184bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U184bar (
    .O(n774bar),
    .I0(n773bar),
    .I1(n772bar)
  );
  //OR U185
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U185 (
    .O(n772),
    .I0(in[131]),
    .I1(in[120])
  );
  //AND U185bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U185bar (
    .O(n772bar),
    .I0(inbar[131]),
    .I1(inbar[120])
  );
  //OR U186
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U186 (
    .O(n773),
    .I0(in[153]),
    .I1(in[147])
  );
  //AND U186bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U186bar (
    .O(n773bar),
    .I0(inbar[153]),
    .I1(inbar[147])
  );
  //OR U187
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U187 (
    .O(n775),
    .I0(n771),
    .I1(n770)
  );
  //AND U187bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U187bar (
    .O(n775bar),
    .I0(n771bar),
    .I1(n770bar)
  );
  //OR U188
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U188 (
    .O(n770),
    .I0(in[170]),
    .I1(in[156])
  );
  //AND U188bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U188bar (
    .O(n770bar),
    .I0(inbar[170]),
    .I1(inbar[156])
  );
  //OR U189
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U189 (
    .O(n771),
    .I0(in[223]),
    .I1(in[190])
  );
  //AND U189bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U189bar (
    .O(n771bar),
    .I0(inbar[223]),
    .I1(inbar[190])
  );
  //OR U190
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U190 (
    .O(n777),
    .I0(n769),
    .I1(n768)
  );
  //AND U190bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U190bar (
    .O(n777bar),
    .I0(n769bar),
    .I1(n768bar)
  );
  //OR U191
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U191 (
    .O(n768),
    .I0(n767),
    .I1(n766)
  );
  //AND U191bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U191bar (
    .O(n768bar),
    .I0(n767bar),
    .I1(n766bar)
  );
  //OR U192
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U192 (
    .O(n766),
    .I0(in[236]),
    .I1(in[230])
  );
  //AND U192bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U192bar (
    .O(n766bar),
    .I0(inbar[236]),
    .I1(inbar[230])
  );
  //OR U193
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U193 (
    .O(n767),
    .I0(in[85]),
    .I1(in[240])
  );
  //AND U193bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U193bar (
    .O(n767bar),
    .I0(inbar[85]),
    .I1(inbar[240])
  );
  //OR U194
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U194 (
    .O(n769),
    .I0(n765),
    .I1(n764)
  );
  //AND U194bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U194bar (
    .O(n769bar),
    .I0(n765bar),
    .I1(n764bar)
  );
  //OR U195
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U195 (
    .O(n764),
    .I0(in_12),
    .I1(in[90])
  );
  //AND U195bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U195bar (
    .O(n764bar),
    .I0(in_12bar),
    .I1(inbar[90])
  );
  //OR U196
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U196 (
    .O(n765),
    .I0(in_39),
    .I1(in_28)
  );
  //AND U196bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U196bar (
    .O(n765bar),
    .I0(in_39bar),
    .I1(in_28bar)
  );
  //OR U197
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U197 (
    .O(n780),
    .I0(in[109]),
    .I1(n763)
  );
  //AND U197bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U197bar (
    .O(n780bar),
    .I0(inbar[109]),
    .I1(n763bar)
  );
  //OR U198
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U198 (
    .O(n782),
    .I0(n762),
    .I1(n761)
  );
  //AND U198bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U198bar (
    .O(n782bar),
    .I0(n762bar),
    .I1(n761bar)
  );
  //OR U199
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U199 (
    .O(n761),
    .I0(in[138]),
    .I1(in[129])
  );
  //AND U199bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U199bar (
    .O(n761bar),
    .I0(inbar[138]),
    .I1(inbar[129])
  );
  //OR U200
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U200 (
    .O(n762),
    .I0(in[157]),
    .I1(n760)
  );
  //AND U200bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U200bar (
    .O(n762bar),
    .I0(inbar[157]),
    .I1(n760bar)
  );
  //OR U201
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U201 (
    .O(n760),
    .I0(in[182]),
    .I1(in[167])
  );
  //AND U201bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U201bar (
    .O(n760bar),
    .I0(inbar[182]),
    .I1(inbar[167])
  );
  //OR U202
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U202 (
    .O(n784),
    .I0(n759),
    .I1(n758)
  );
  //AND U202bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U202bar (
    .O(n784bar),
    .I0(n759bar),
    .I1(n758bar)
  );
  //OR U203
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U203 (
    .O(n758),
    .I0(n757),
    .I1(n756)
  );
  //AND U203bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U203bar (
    .O(n758bar),
    .I0(n757bar),
    .I1(n756bar)
  );
  //OR U204
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U204 (
    .O(n756),
    .I0(in[195]),
    .I1(in[184])
  );
  //AND U204bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U204bar (
    .O(n756bar),
    .I0(inbar[195]),
    .I1(inbar[184])
  );
  //OR U205
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U205 (
    .O(n757),
    .I0(in[196]),
    .I1(n755)
  );
  //AND U205bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U205bar (
    .O(n757bar),
    .I0(inbar[196]),
    .I1(n755bar)
  );
  //OR U206
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U206 (
    .O(n755),
    .I0(in[215]),
    .I1(in[209])
  );
  //AND U206bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U206bar (
    .O(n755bar),
    .I0(inbar[215]),
    .I1(inbar[209])
  );
  //OR U207
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U207 (
    .O(n759),
    .I0(n754),
    .I1(n753)
  );
  //AND U207bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U207bar (
    .O(n759bar),
    .I0(n754bar),
    .I1(n753bar)
  );
  //OR U208
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U208 (
    .O(n753),
    .I0(in[93]),
    .I1(in[233])
  );
  //AND U208bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U208bar (
    .O(n753bar),
    .I0(inbar[93]),
    .I1(inbar[233])
  );
  //OR U209
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U209 (
    .O(n754),
    .I0(in_1),
    .I1(n752)
  );
  //AND U209bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U209bar (
    .O(n754bar),
    .I0(in_1bar),
    .I1(n752bar)
  );
  //OR U210
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U210 (
    .O(n752),
    .I0(in_69),
    .I1(in_66)
  );
  //AND U210bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U210bar (
    .O(n752bar),
    .I0(in_69bar),
    .I1(in_66bar)
  );
  //OR U211
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U211 (
    .O(n787),
    .I0(n966),
    .I1(n751)
  );
  //AND U211bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U211bar (
    .O(n787bar),
    .I0(n966bar),
    .I1(n751bar)
  );
  //OR U212
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U212 (
    .O(n751),
    .I0(in[134]),
    .I1(n750)
  );
  //AND U212bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U212bar (
    .O(n751bar),
    .I0(inbar[134]),
    .I1(n750bar)
  );
  //OR U213
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U213 (
    .O(n966),
    .I0(n749),
    .I1(n748)
  );
  //AND U213bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U213bar (
    .O(n966bar),
    .I0(n749bar),
    .I1(n748bar)
  );
  //OR U214
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U214 (
    .O(n748),
    .I0(n747),
    .I1(n746)
  );
  //AND U214bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U214bar (
    .O(n748bar),
    .I0(n747bar),
    .I1(n746bar)
  );
  //OR U215
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U215 (
    .O(n746),
    .I0(n745),
    .I1(n744)
  );
  //AND U215bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U215bar (
    .O(n746bar),
    .I0(n745bar),
    .I1(n744bar)
  );
  //OR U216
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U216 (
    .O(n744),
    .I0(in[136]),
    .I1(in[121])
  );
  //AND U216bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U216bar (
    .O(n744bar),
    .I0(inbar[136]),
    .I1(inbar[121])
  );
  //OR U217
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U217 (
    .O(n745),
    .I0(in[186]),
    .I1(in[174])
  );
  //AND U217bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U217bar (
    .O(n745bar),
    .I0(inbar[186]),
    .I1(inbar[174])
  );
  //OR U218
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U218 (
    .O(n747),
    .I0(n743),
    .I1(n742)
  );
  //AND U218bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U218bar (
    .O(n747bar),
    .I0(n743bar),
    .I1(n742bar)
  );
  //OR U219
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U219 (
    .O(n742),
    .I0(in[198]),
    .I1(in[197])
  );
  //AND U219bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U219bar (
    .O(n742bar),
    .I0(inbar[198]),
    .I1(inbar[197])
  );
  //OR U220
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U220 (
    .O(n743),
    .I0(in[214]),
    .I1(in[199])
  );
  //AND U220bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U220bar (
    .O(n743bar),
    .I0(inbar[214]),
    .I1(inbar[199])
  );
  //OR U221
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U221 (
    .O(n749),
    .I0(n741),
    .I1(n740)
  );
  //AND U221bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U221bar (
    .O(n749bar),
    .I0(n741bar),
    .I1(n740bar)
  );
  //OR U222
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U222 (
    .O(n740),
    .I0(n739),
    .I1(n738)
  );
  //AND U222bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U222bar (
    .O(n740bar),
    .I0(n739bar),
    .I1(n738bar)
  );
  //OR U223
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U223 (
    .O(n738),
    .I0(in[231]),
    .I1(in[220])
  );
  //AND U223bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U223bar (
    .O(n738bar),
    .I0(inbar[231]),
    .I1(inbar[220])
  );
  //OR U224
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U224 (
    .O(n739),
    .I0(in_25),
    .I1(in[245])
  );
  //AND U224bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U224bar (
    .O(n739bar),
    .I0(in_25bar),
    .I1(inbar[245])
  );
  //OR U225
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U225 (
    .O(n741),
    .I0(n737),
    .I1(n736)
  );
  //AND U225bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U225bar (
    .O(n741bar),
    .I0(n737bar),
    .I1(n736bar)
  );
  //OR U226
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U226 (
    .O(n736),
    .I0(in_53),
    .I1(in_29)
  );
  //AND U226bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U226bar (
    .O(n736bar),
    .I0(in_53bar),
    .I1(in_29bar)
  );
  //OR U227
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U227 (
    .O(n737),
    .I0(in_79),
    .I1(in_74)
  );
  //AND U227bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U227bar (
    .O(n737bar),
    .I0(in_79bar),
    .I1(in_74bar)
  );
  //OR U228
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U228 (
    .O(n789),
    .I0(n735),
    .I1(n734)
  );
  //AND U228bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U228bar (
    .O(n789bar),
    .I0(n735bar),
    .I1(n734bar)
  );
  //OR U229
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U229 (
    .O(n734),
    .I0(in[152]),
    .I1(in[140])
  );
  //AND U229bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U229bar (
    .O(n734bar),
    .I0(inbar[152]),
    .I1(inbar[140])
  );
  //OR U230
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U230 (
    .O(n735),
    .I0(in[155]),
    .I1(n733)
  );
  //AND U230bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U230bar (
    .O(n735bar),
    .I0(inbar[155]),
    .I1(n733bar)
  );
  //OR U231
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U231 (
    .O(n733),
    .I0(in[166]),
    .I1(in[165])
  );
  //AND U231bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U231bar (
    .O(n733bar),
    .I0(inbar[166]),
    .I1(inbar[165])
  );
  //OR U232
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U232 (
    .O(n791),
    .I0(n732),
    .I1(n731)
  );
  //AND U232bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U232bar (
    .O(n791bar),
    .I0(n732bar),
    .I1(n731bar)
  );
  //OR U233
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U233 (
    .O(n731),
    .I0(n730),
    .I1(n729)
  );
  //AND U233bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U233bar (
    .O(n731bar),
    .I0(n730bar),
    .I1(n729bar)
  );
  //OR U234
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U234 (
    .O(n729),
    .I0(in[202]),
    .I1(in[185])
  );
  //AND U234bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U234bar (
    .O(n729bar),
    .I0(inbar[202]),
    .I1(inbar[185])
  );
  //OR U235
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U235 (
    .O(n730),
    .I0(in[211]),
    .I1(n728)
  );
  //AND U235bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U235bar (
    .O(n730bar),
    .I0(inbar[211]),
    .I1(n728bar)
  );
  //OR U236
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U236 (
    .O(n728),
    .I0(in[255]),
    .I1(in[253])
  );
  //AND U236bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U236bar (
    .O(n728bar),
    .I0(inbar[255]),
    .I1(inbar[253])
  );
  //OR U237
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U237 (
    .O(n732),
    .I0(n727),
    .I1(n726)
  );
  //AND U237bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U237bar (
    .O(n732bar),
    .I0(n727bar),
    .I1(n726bar)
  );
  //OR U238
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U238 (
    .O(n726),
    .I0(in_35),
    .I1(in_15)
  );
  //AND U238bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U238bar (
    .O(n726bar),
    .I0(in_35bar),
    .I1(in_15bar)
  );
  //OR U239
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U239 (
    .O(n727),
    .I0(in_36),
    .I1(n725)
  );
  //AND U239bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U239bar (
    .O(n727bar),
    .I0(in_36bar),
    .I1(n725bar)
  );
  //OR U240
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U240 (
    .O(n725),
    .I0(in_48),
    .I1(in_40)
  );
  //AND U240bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U240bar (
    .O(n725bar),
    .I0(in_48bar),
    .I1(in_40bar)
  );
  //OR U241
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U241 (
    .O(out[1]),
    .I0(n724),
    .I1(n723)
  );
  //AND U241bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U241bar (
    .O(outbar[1]),
    .I0(n724bar),
    .I1(n723bar)
  );
  //OR U242
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U242 (
    .O(n723),
    .I0(n722),
    .I1(n721)
  );
  //AND U242bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U242bar (
    .O(n723bar),
    .I0(n722bar),
    .I1(n721bar)
  );
  //OR U243
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U243 (
    .O(n721),
    .I0(n720),
    .I1(n719)
  );
  //AND U243bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U243bar (
    .O(n721bar),
    .I0(n720bar),
    .I1(n719bar)
  );
  //OR U244
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U244 (
    .O(n719),
    .I0(n921),
    .I1(n887)
  );
  //AND U244bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U244bar (
    .O(n719bar),
    .I0(n921bar),
    .I1(n887bar)
  );
  //OR U245
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U245 (
    .O(n887),
    .I0(n718),
    .I1(n717)
  );
  //AND U245bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U245bar (
    .O(n887bar),
    .I0(n718bar),
    .I1(n717bar)
  );
  //OR U246
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U246 (
    .O(n717),
    .I0(n716),
    .I1(n715)
  );
  //AND U246bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U246bar (
    .O(n717bar),
    .I0(n716bar),
    .I1(n715bar)
  );
  //OR U247
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U247 (
    .O(n715),
    .I0(n714),
    .I1(n713)
  );
  //AND U247bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U247bar (
    .O(n715bar),
    .I0(n714bar),
    .I1(n713bar)
  );
  //OR U248
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U248 (
    .O(n713),
    .I0(in[116]),
    .I1(in[110])
  );
  //AND U248bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U248bar (
    .O(n713bar),
    .I0(inbar[116]),
    .I1(inbar[110])
  );
  //OR U249
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U249 (
    .O(n714),
    .I0(in[133]),
    .I1(in[130])
  );
  //AND U249bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U249bar (
    .O(n714bar),
    .I0(inbar[133]),
    .I1(inbar[130])
  );
  //OR U250
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U250 (
    .O(n716),
    .I0(n712),
    .I1(n711)
  );
  //AND U250bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U250bar (
    .O(n716bar),
    .I0(n712bar),
    .I1(n711bar)
  );
  //OR U251
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U251 (
    .O(n711),
    .I0(in[203]),
    .I1(in[135])
  );
  //AND U251bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U251bar (
    .O(n711bar),
    .I0(inbar[203]),
    .I1(inbar[135])
  );
  //OR U252
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U252 (
    .O(n712),
    .I0(in[232]),
    .I1(in[223])
  );
  //AND U252bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U252bar (
    .O(n712bar),
    .I0(inbar[232]),
    .I1(inbar[223])
  );
  //OR U253
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U253 (
    .O(n718),
    .I0(n710),
    .I1(n709)
  );
  //AND U253bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U253bar (
    .O(n718bar),
    .I0(n710bar),
    .I1(n709bar)
  );
  //OR U254
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U254 (
    .O(n709),
    .I0(n708),
    .I1(n707)
  );
  //AND U254bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U254bar (
    .O(n709bar),
    .I0(n708bar),
    .I1(n707bar)
  );
  //OR U255
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U255 (
    .O(n707),
    .I0(in[255]),
    .I1(in[233])
  );
  //AND U255bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U255bar (
    .O(n707bar),
    .I0(inbar[255]),
    .I1(inbar[233])
  );
  //OR U256
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U256 (
    .O(n708),
    .I0(in_53),
    .I1(in_34)
  );
  //AND U256bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U256bar (
    .O(n708bar),
    .I0(in_53bar),
    .I1(in_34bar)
  );
  //OR U257
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U257 (
    .O(n710),
    .I0(n706),
    .I1(n705)
  );
  //AND U257bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U257bar (
    .O(n710bar),
    .I0(n706bar),
    .I1(n705bar)
  );
  //OR U258
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U258 (
    .O(n705),
    .I0(in_57),
    .I1(in_55)
  );
  //AND U258bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U258bar (
    .O(n705bar),
    .I0(in_57bar),
    .I1(in_55bar)
  );
  //OR U259
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U259 (
    .O(n706),
    .I0(in_68),
    .I1(in_67)
  );
  //AND U259bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U259bar (
    .O(n706bar),
    .I0(in_68bar),
    .I1(in_67bar)
  );
  //OR U260
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U260 (
    .O(n921),
    .I0(n704),
    .I1(n703)
  );
  //AND U260bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U260bar (
    .O(n921bar),
    .I0(n704bar),
    .I1(n703bar)
  );
  //OR U261
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U261 (
    .O(n703),
    .I0(n702),
    .I1(n701)
  );
  //AND U261bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U261bar (
    .O(n703bar),
    .I0(n702bar),
    .I1(n701bar)
  );
  //OR U262
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U262 (
    .O(n701),
    .I0(n700),
    .I1(n699)
  );
  //AND U262bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U262bar (
    .O(n701bar),
    .I0(n700bar),
    .I1(n699bar)
  );
  //OR U263
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U263 (
    .O(n699),
    .I0(n944),
    .I1(n872)
  );
  //AND U263bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U263bar (
    .O(n699bar),
    .I0(n944bar),
    .I1(n872bar)
  );
  //OR U264
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U264 (
    .O(n872),
    .I0(n698),
    .I1(n697)
  );
  //AND U264bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U264bar (
    .O(n872bar),
    .I0(n698bar),
    .I1(n697bar)
  );
  //OR U265
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U265 (
    .O(n697),
    .I0(n696),
    .I1(n695)
  );
  //AND U265bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U265bar (
    .O(n697bar),
    .I0(n696bar),
    .I1(n695bar)
  );
  //OR U266
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U266 (
    .O(n695),
    .I0(n694),
    .I1(n693)
  );
  //AND U266bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U266bar (
    .O(n695bar),
    .I0(n694bar),
    .I1(n693bar)
  );
  //OR U267
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U267 (
    .O(n693),
    .I0(in[121]),
    .I1(in[102])
  );
  //AND U267bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U267bar (
    .O(n693bar),
    .I0(inbar[121]),
    .I1(inbar[102])
  );
  //OR U268
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U268 (
    .O(n694),
    .I0(in[162]),
    .I1(in[161])
  );
  //AND U268bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U268bar (
    .O(n694bar),
    .I0(inbar[162]),
    .I1(inbar[161])
  );
  //OR U269
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U269 (
    .O(n696),
    .I0(n692),
    .I1(n691)
  );
  //AND U269bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U269bar (
    .O(n696bar),
    .I0(n692bar),
    .I1(n691bar)
  );
  //OR U270
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U270 (
    .O(n691),
    .I0(in[192]),
    .I1(in[178])
  );
  //AND U270bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U270bar (
    .O(n691bar),
    .I0(inbar[192]),
    .I1(inbar[178])
  );
  //OR U271
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U271 (
    .O(n692),
    .I0(in[244]),
    .I1(in[209])
  );
  //AND U271bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U271bar (
    .O(n692bar),
    .I0(inbar[244]),
    .I1(inbar[209])
  );
  //OR U272
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U272 (
    .O(n698),
    .I0(n690),
    .I1(n689)
  );
  //AND U272bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U272bar (
    .O(n698bar),
    .I0(n690bar),
    .I1(n689bar)
  );
  //OR U273
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U273 (
    .O(n689),
    .I0(n688),
    .I1(n687)
  );
  //AND U273bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U273bar (
    .O(n689bar),
    .I0(n688bar),
    .I1(n687bar)
  );
  //OR U274
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U274 (
    .O(n687),
    .I0(in[90]),
    .I1(in[254])
  );
  //AND U274bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U274bar (
    .O(n687bar),
    .I0(inbar[90]),
    .I1(inbar[254])
  );
  //OR U275
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U275 (
    .O(n688),
    .I0(in_36),
    .I1(in_32)
  );
  //AND U275bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U275bar (
    .O(n688bar),
    .I0(in_36bar),
    .I1(in_32bar)
  );
  //OR U276
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U276 (
    .O(n690),
    .I0(n686),
    .I1(n685)
  );
  //AND U276bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U276bar (
    .O(n690bar),
    .I0(n686bar),
    .I1(n685bar)
  );
  //OR U277
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U277 (
    .O(n685),
    .I0(in_62),
    .I1(in_37)
  );
  //AND U277bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U277bar (
    .O(n685bar),
    .I0(in_62bar),
    .I1(in_37bar)
  );
  //OR U278
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U278 (
    .O(n686),
    .I0(in_75),
    .I1(in_73)
  );
  //AND U278bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U278bar (
    .O(n686bar),
    .I0(in_75bar),
    .I1(in_73bar)
  );
  //OR U279
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U279 (
    .O(n944),
    .I0(n684),
    .I1(n683)
  );
  //AND U279bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U279bar (
    .O(n944bar),
    .I0(n684bar),
    .I1(n683bar)
  );
  //OR U280
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U280 (
    .O(n683),
    .I0(n682),
    .I1(n681)
  );
  //AND U280bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U280bar (
    .O(n683bar),
    .I0(n682bar),
    .I1(n681bar)
  );
  //OR U281
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U281 (
    .O(n681),
    .I0(n680),
    .I1(n679)
  );
  //AND U281bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U281bar (
    .O(n681bar),
    .I0(n680bar),
    .I1(n679bar)
  );
  //OR U282
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U282 (
    .O(n679),
    .I0(in[171]),
    .I1(in[153])
  );
  //AND U282bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U282bar (
    .O(n679bar),
    .I0(inbar[171]),
    .I1(inbar[153])
  );
  //OR U283
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U283 (
    .O(n680),
    .I0(in[187]),
    .I1(in[176])
  );
  //AND U283bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U283bar (
    .O(n680bar),
    .I0(inbar[187]),
    .I1(inbar[176])
  );
  //OR U284
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U284 (
    .O(n682),
    .I0(n678),
    .I1(n677)
  );
  //AND U284bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U284bar (
    .O(n682bar),
    .I0(n678bar),
    .I1(n677bar)
  );
  //OR U285
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U285 (
    .O(n677),
    .I0(in[245]),
    .I1(in[211])
  );
  //AND U285bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U285bar (
    .O(n677bar),
    .I0(inbar[245]),
    .I1(inbar[211])
  );
  //OR U286
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U286 (
    .O(n678),
    .I0(in[97]),
    .I1(in[88])
  );
  //AND U286bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U286bar (
    .O(n678bar),
    .I0(inbar[97]),
    .I1(inbar[88])
  );
  //OR U287
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U287 (
    .O(n684),
    .I0(n676),
    .I1(n675)
  );
  //AND U287bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U287bar (
    .O(n684bar),
    .I0(n676bar),
    .I1(n675bar)
  );
  //OR U288
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U288 (
    .O(n675),
    .I0(n674),
    .I1(n673)
  );
  //AND U288bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U288bar (
    .O(n675bar),
    .I0(n674bar),
    .I1(n673bar)
  );
  //OR U289
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U289 (
    .O(n673),
    .I0(in_10),
    .I1(in_0)
  );
  //AND U289bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U289bar (
    .O(n673bar),
    .I0(in_10bar),
    .I1(in_0bar)
  );
  //OR U290
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U290 (
    .O(n674),
    .I0(in_59),
    .I1(in_5)
  );
  //AND U290bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U290bar (
    .O(n674bar),
    .I0(in_59bar),
    .I1(in_5bar)
  );
  //OR U291
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U291 (
    .O(n676),
    .I0(n672),
    .I1(n671)
  );
  //AND U291bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U291bar (
    .O(n676bar),
    .I0(n672bar),
    .I1(n671bar)
  );
  //OR U292
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U292 (
    .O(n671),
    .I0(in_60),
    .I1(in_6)
  );
  //AND U292bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U292bar (
    .O(n671bar),
    .I0(in_60bar),
    .I1(in_6bar)
  );
  //OR U293
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U293 (
    .O(n672),
    .I0(in_77),
    .I1(in_69)
  );
  //AND U293bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U293bar (
    .O(n672bar),
    .I0(in_77bar),
    .I1(in_69bar)
  );
  //OR U294
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U294 (
    .O(n700),
    .I0(in[113]),
    .I1(n864)
  );
  //AND U294bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U294bar (
    .O(n700bar),
    .I0(inbar[113]),
    .I1(n864bar)
  );
  //OR U295
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U295 (
    .O(n864),
    .I0(n670),
    .I1(n669)
  );
  //AND U295bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U295bar (
    .O(n864bar),
    .I0(n670bar),
    .I1(n669bar)
  );
  //OR U296
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U296 (
    .O(n669),
    .I0(n668),
    .I1(n667)
  );
  //AND U296bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U296bar (
    .O(n669bar),
    .I0(n668bar),
    .I1(n667bar)
  );
  //OR U297
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U297 (
    .O(n667),
    .I0(n666),
    .I1(n665)
  );
  //AND U297bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U297bar (
    .O(n667bar),
    .I0(n666bar),
    .I1(n665bar)
  );
  //OR U298
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U298 (
    .O(n665),
    .I0(in[125]),
    .I1(in[107])
  );
  //AND U298bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U298bar (
    .O(n665bar),
    .I0(inbar[125]),
    .I1(inbar[107])
  );
  //OR U299
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U299 (
    .O(n666),
    .I0(in[138]),
    .I1(in[126])
  );
  //AND U299bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U299bar (
    .O(n666bar),
    .I0(inbar[138]),
    .I1(inbar[126])
  );
  //OR U300
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U300 (
    .O(n668),
    .I0(n664),
    .I1(n663)
  );
  //AND U300bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U300bar (
    .O(n668bar),
    .I0(n664bar),
    .I1(n663bar)
  );
  //OR U301
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U301 (
    .O(n663),
    .I0(in[189]),
    .I1(in[143])
  );
  //AND U301bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U301bar (
    .O(n663bar),
    .I0(inbar[189]),
    .I1(inbar[143])
  );
  //OR U302
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U302 (
    .O(n664),
    .I0(in[99]),
    .I1(in[214])
  );
  //AND U302bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U302bar (
    .O(n664bar),
    .I0(inbar[99]),
    .I1(inbar[214])
  );
  //OR U303
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U303 (
    .O(n670),
    .I0(n662),
    .I1(n661)
  );
  //AND U303bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U303bar (
    .O(n670bar),
    .I0(n662bar),
    .I1(n661bar)
  );
  //OR U304
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U304 (
    .O(n661),
    .I0(n660),
    .I1(n659)
  );
  //AND U304bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U304bar (
    .O(n661bar),
    .I0(n660bar),
    .I1(n659bar)
  );
  //OR U305
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U305 (
    .O(n659),
    .I0(in_15),
    .I1(in_12)
  );
  //AND U305bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U305bar (
    .O(n659bar),
    .I0(in_15bar),
    .I1(in_12bar)
  );
  //OR U306
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U306 (
    .O(n660),
    .I0(in_20),
    .I1(in_2)
  );
  //AND U306bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U306bar (
    .O(n660bar),
    .I0(in_20bar),
    .I1(in_2bar)
  );
  //OR U307
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U307 (
    .O(n662),
    .I0(n658),
    .I1(n657)
  );
  //AND U307bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U307bar (
    .O(n662bar),
    .I0(n658bar),
    .I1(n657bar)
  );
  //OR U308
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U308 (
    .O(n657),
    .I0(in_30),
    .I1(in_3)
  );
  //AND U308bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U308bar (
    .O(n657bar),
    .I0(in_30bar),
    .I1(in_3bar)
  );
  //OR U309
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U309 (
    .O(n658),
    .I0(in_4),
    .I1(in_38)
  );
  //AND U309bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U309bar (
    .O(n658bar),
    .I0(in_4bar),
    .I1(in_38bar)
  );
  //OR U310
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U310 (
    .O(n702),
    .I0(n656),
    .I1(n655)
  );
  //AND U310bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U310bar (
    .O(n702bar),
    .I0(n656bar),
    .I1(n655bar)
  );
  //OR U311
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U311 (
    .O(n655),
    .I0(in[148]),
    .I1(in[137])
  );
  //AND U311bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U311bar (
    .O(n655bar),
    .I0(inbar[148]),
    .I1(inbar[137])
  );
  //OR U312
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U312 (
    .O(n656),
    .I0(in[149]),
    .I1(n654)
  );
  //AND U312bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U312bar (
    .O(n656bar),
    .I0(inbar[149]),
    .I1(n654bar)
  );
  //OR U313
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U313 (
    .O(n654),
    .I0(in[195]),
    .I1(in[190])
  );
  //AND U313bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U313bar (
    .O(n654bar),
    .I0(inbar[195]),
    .I1(inbar[190])
  );
  //OR U314
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U314 (
    .O(n704),
    .I0(n653),
    .I1(n652)
  );
  //AND U314bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U314bar (
    .O(n704bar),
    .I0(n653bar),
    .I1(n652bar)
  );
  //OR U315
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U315 (
    .O(n652),
    .I0(n651),
    .I1(n650)
  );
  //AND U315bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U315bar (
    .O(n652bar),
    .I0(n651bar),
    .I1(n650bar)
  );
  //OR U316
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U316 (
    .O(n650),
    .I0(in[98]),
    .I1(in[197])
  );
  //AND U316bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U316bar (
    .O(n650bar),
    .I0(inbar[98]),
    .I1(inbar[197])
  );
  //OR U317
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U317 (
    .O(n651),
    .I0(in_11),
    .I1(n649)
  );
  //AND U317bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U317bar (
    .O(n651bar),
    .I0(in_11bar),
    .I1(n649bar)
  );
  //OR U318
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U318 (
    .O(n649),
    .I0(in_26),
    .I1(in_14)
  );
  //AND U318bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U318bar (
    .O(n649bar),
    .I0(in_26bar),
    .I1(in_14bar)
  );
  //OR U319
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U319 (
    .O(n653),
    .I0(n648),
    .I1(n647)
  );
  //AND U319bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U319bar (
    .O(n653bar),
    .I0(n648bar),
    .I1(n647bar)
  );
  //OR U320
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U320 (
    .O(n647),
    .I0(in_35),
    .I1(in_27)
  );
  //AND U320bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U320bar (
    .O(n647bar),
    .I0(in_35bar),
    .I1(in_27bar)
  );
  //OR U321
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U321 (
    .O(n648),
    .I0(in_50),
    .I1(n646)
  );
  //AND U321bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U321bar (
    .O(n648bar),
    .I0(in_50bar),
    .I1(n646bar)
  );
  //OR U322
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U322 (
    .O(n646),
    .I0(in_78),
    .I1(in_61)
  );
  //AND U322bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U322bar (
    .O(n646bar),
    .I0(in_78bar),
    .I1(in_61bar)
  );
  //OR U323
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U323 (
    .O(n720),
    .I0(n942),
    .I1(n645)
  );
  //AND U323bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U323bar (
    .O(n720bar),
    .I0(n942bar),
    .I1(n645bar)
  );
  //OR U324
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U324 (
    .O(n645),
    .I0(in[106]),
    .I1(n863)
  );
  //AND U324bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U324bar (
    .O(n645bar),
    .I0(inbar[106]),
    .I1(n863bar)
  );
  //OR U325
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U325 (
    .O(n863),
    .I0(n644),
    .I1(n643)
  );
  //AND U325bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U325bar (
    .O(n863bar),
    .I0(n644bar),
    .I1(n643bar)
  );
  //OR U326
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U326 (
    .O(n643),
    .I0(n642),
    .I1(n641)
  );
  //AND U326bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U326bar (
    .O(n643bar),
    .I0(n642bar),
    .I1(n641bar)
  );
  //OR U327
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U327 (
    .O(n641),
    .I0(n640),
    .I1(n639)
  );
  //AND U327bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U327bar (
    .O(n641bar),
    .I0(n640bar),
    .I1(n639bar)
  );
  //OR U328
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U328 (
    .O(n639),
    .I0(in[127]),
    .I1(in[122])
  );
  //AND U328bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U328bar (
    .O(n639bar),
    .I0(inbar[127]),
    .I1(inbar[122])
  );
  //OR U329
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U329 (
    .O(n640),
    .I0(in[156]),
    .I1(in[132])
  );
  //AND U329bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U329bar (
    .O(n640bar),
    .I0(inbar[156]),
    .I1(inbar[132])
  );
  //OR U330
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U330 (
    .O(n642),
    .I0(n638),
    .I1(n637)
  );
  //AND U330bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U330bar (
    .O(n642bar),
    .I0(n638bar),
    .I1(n637bar)
  );
  //OR U331
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U331 (
    .O(n637),
    .I0(in[159]),
    .I1(in[157])
  );
  //AND U331bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U331bar (
    .O(n637bar),
    .I0(inbar[159]),
    .I1(inbar[157])
  );
  //OR U332
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U332 (
    .O(n638),
    .I0(in[185]),
    .I1(in[169])
  );
  //AND U332bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U332bar (
    .O(n638bar),
    .I0(inbar[185]),
    .I1(inbar[169])
  );
  //OR U333
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U333 (
    .O(n644),
    .I0(n636),
    .I1(n635)
  );
  //AND U333bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U333bar (
    .O(n644bar),
    .I0(n636bar),
    .I1(n635bar)
  );
  //OR U334
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U334 (
    .O(n635),
    .I0(n634),
    .I1(n633)
  );
  //AND U334bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U334bar (
    .O(n635bar),
    .I0(n634bar),
    .I1(n633bar)
  );
  //OR U335
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U335 (
    .O(n633),
    .I0(in[239]),
    .I1(in[218])
  );
  //AND U335bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U335bar (
    .O(n633bar),
    .I0(inbar[239]),
    .I1(inbar[218])
  );
  //OR U336
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U336 (
    .O(n634),
    .I0(in_13),
    .I1(in[87])
  );
  //AND U336bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U336bar (
    .O(n634bar),
    .I0(in_13bar),
    .I1(inbar[87])
  );
  //OR U337
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U337 (
    .O(n636),
    .I0(n632),
    .I1(n631)
  );
  //AND U337bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U337bar (
    .O(n636bar),
    .I0(n632bar),
    .I1(n631bar)
  );
  //OR U338
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U338 (
    .O(n631),
    .I0(in_72),
    .I1(in_70)
  );
  //AND U338bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U338bar (
    .O(n631bar),
    .I0(in_72bar),
    .I1(in_70bar)
  );
  //OR U339
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U339 (
    .O(n632),
    .I0(in_80),
    .I1(in_74)
  );
  //AND U339bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U339bar (
    .O(n632bar),
    .I0(in_80bar),
    .I1(in_74bar)
  );
  //OR U340
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U340 (
    .O(n942),
    .I0(n630),
    .I1(n629)
  );
  //AND U340bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U340bar (
    .O(n942bar),
    .I0(n630bar),
    .I1(n629bar)
  );
  //OR U341
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U341 (
    .O(n629),
    .I0(n628),
    .I1(n627)
  );
  //AND U341bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U341bar (
    .O(n629bar),
    .I0(n628bar),
    .I1(n627bar)
  );
  //OR U342
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U342 (
    .O(n627),
    .I0(n626),
    .I1(n625)
  );
  //AND U342bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U342bar (
    .O(n627bar),
    .I0(n626bar),
    .I1(n625bar)
  );
  //OR U343
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U343 (
    .O(n625),
    .I0(in[146]),
    .I1(in[100])
  );
  //AND U343bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U343bar (
    .O(n625bar),
    .I0(inbar[146]),
    .I1(inbar[100])
  );
  //OR U344
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U344 (
    .O(n626),
    .I0(in[168]),
    .I1(in[152])
  );
  //AND U344bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U344bar (
    .O(n626bar),
    .I0(inbar[168]),
    .I1(inbar[152])
  );
  //OR U345
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U345 (
    .O(n628),
    .I0(n624),
    .I1(n623)
  );
  //AND U345bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U345bar (
    .O(n628bar),
    .I0(n624bar),
    .I1(n623bar)
  );
  //OR U346
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U346 (
    .O(n623),
    .I0(in[199]),
    .I1(in[182])
  );
  //AND U346bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U346bar (
    .O(n623bar),
    .I0(inbar[199]),
    .I1(inbar[182])
  );
  //OR U347
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U347 (
    .O(n624),
    .I0(in[236]),
    .I1(in[204])
  );
  //AND U347bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U347bar (
    .O(n624bar),
    .I0(inbar[236]),
    .I1(inbar[204])
  );
  //OR U348
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U348 (
    .O(n630),
    .I0(n622),
    .I1(n621)
  );
  //AND U348bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U348bar (
    .O(n630bar),
    .I0(n622bar),
    .I1(n621bar)
  );
  //OR U349
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U349 (
    .O(n621),
    .I0(n620),
    .I1(n619)
  );
  //AND U349bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U349bar (
    .O(n621bar),
    .I0(n620bar),
    .I1(n619bar)
  );
  //OR U350
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U350 (
    .O(n619),
    .I0(in[89]),
    .I1(in[246])
  );
  //AND U350bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U350bar (
    .O(n619bar),
    .I0(inbar[89]),
    .I1(inbar[246])
  );
  //OR U351
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U351 (
    .O(n620),
    .I0(in[95]),
    .I1(in[92])
  );
  //AND U351bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U351bar (
    .O(n620bar),
    .I0(inbar[95]),
    .I1(inbar[92])
  );
  //OR U352
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U352 (
    .O(n622),
    .I0(n618),
    .I1(n617)
  );
  //AND U352bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U352bar (
    .O(n622bar),
    .I0(n618bar),
    .I1(n617bar)
  );
  //OR U353
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U353 (
    .O(n617),
    .I0(in_22),
    .I1(in_16)
  );
  //AND U353bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U353bar (
    .O(n617bar),
    .I0(in_22bar),
    .I1(in_16bar)
  );
  //OR U354
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U354 (
    .O(n618),
    .I0(in_51),
    .I1(in_49)
  );
  //AND U354bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U354bar (
    .O(n618bar),
    .I0(in_51bar),
    .I1(in_49bar)
  );
  //OR U355
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U355 (
    .O(n722),
    .I0(n616),
    .I1(n615)
  );
  //AND U355bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U355bar (
    .O(n722bar),
    .I0(n616bar),
    .I1(n615bar)
  );
  //OR U356
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U356 (
    .O(n615),
    .I0(in[158]),
    .I1(in[115])
  );
  //AND U356bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U356bar (
    .O(n615bar),
    .I0(inbar[158]),
    .I1(inbar[115])
  );
  //OR U357
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U357 (
    .O(n616),
    .I0(in[163]),
    .I1(n614)
  );
  //AND U357bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U357bar (
    .O(n616bar),
    .I0(inbar[163]),
    .I1(n614bar)
  );
  //OR U358
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U358 (
    .O(n614),
    .I0(in[206]),
    .I1(in[165])
  );
  //AND U358bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U358bar (
    .O(n614bar),
    .I0(inbar[206]),
    .I1(inbar[165])
  );
  //OR U359
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U359 (
    .O(n724),
    .I0(n613),
    .I1(n612)
  );
  //AND U359bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U359bar (
    .O(n724bar),
    .I0(n613bar),
    .I1(n612bar)
  );
  //OR U360
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U360 (
    .O(n612),
    .I0(n611),
    .I1(n610)
  );
  //AND U360bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U360bar (
    .O(n612bar),
    .I0(n611bar),
    .I1(n610bar)
  );
  //OR U361
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U361 (
    .O(n610),
    .I0(in[213]),
    .I1(in[207])
  );
  //AND U361bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U361bar (
    .O(n610bar),
    .I0(inbar[213]),
    .I1(inbar[207])
  );
  //OR U362
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U362 (
    .O(n611),
    .I0(in[215]),
    .I1(n609)
  );
  //AND U362bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U362bar (
    .O(n611bar),
    .I0(inbar[215]),
    .I1(n609bar)
  );
  //OR U363
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U363 (
    .O(n609),
    .I0(in[230]),
    .I1(in[220])
  );
  //AND U363bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U363bar (
    .O(n609bar),
    .I0(inbar[230]),
    .I1(inbar[220])
  );
  //OR U364
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U364 (
    .O(n613),
    .I0(n608),
    .I1(n607)
  );
  //AND U364bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U364bar (
    .O(n613bar),
    .I0(n608bar),
    .I1(n607bar)
  );
  //OR U365
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U365 (
    .O(n607),
    .I0(in[251]),
    .I1(in[234])
  );
  //AND U365bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U365bar (
    .O(n607bar),
    .I0(inbar[251]),
    .I1(inbar[234])
  );
  //OR U366
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U366 (
    .O(n608),
    .I0(in_17),
    .I1(n606)
  );
  //AND U366bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U366bar (
    .O(n608bar),
    .I0(in_17bar),
    .I1(n606bar)
  );
  //OR U367
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U367 (
    .O(n606),
    .I0(in_65),
    .I1(in_56)
  );
  //AND U367bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U367bar (
    .O(n606bar),
    .I0(in_65bar),
    .I1(in_56bar)
  );
  //OR U368
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U368 (
    .O(out[0]),
    .I0(n605),
    .I1(n604)
  );
  //AND U368bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U368bar (
    .O(outbar[0]),
    .I0(n605bar),
    .I1(n604bar)
  );
  //OR U369
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U369 (
    .O(n604),
    .I0(n603),
    .I1(n602)
  );
  //AND U369bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U369bar (
    .O(n604bar),
    .I0(n603bar),
    .I1(n602bar)
  );
  //OR U370
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U370 (
    .O(n602),
    .I0(n601),
    .I1(n600)
  );
  //AND U370bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U370bar (
    .O(n602bar),
    .I0(n601bar),
    .I1(n600bar)
  );
  //OR U371
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U371 (
    .O(n600),
    .I0(n820),
    .I1(n785)
  );
  //AND U371bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U371bar (
    .O(n600bar),
    .I0(n820bar),
    .I1(n785bar)
  );
  //OR U372
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U372 (
    .O(n785),
    .I0(n599),
    .I1(n598)
  );
  //AND U372bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U372bar (
    .O(n785bar),
    .I0(n599bar),
    .I1(n598bar)
  );
  //OR U373
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U373 (
    .O(n598),
    .I0(n597),
    .I1(n596)
  );
  //AND U373bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U373bar (
    .O(n598bar),
    .I0(n597bar),
    .I1(n596bar)
  );
  //OR U374
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U374 (
    .O(n596),
    .I0(n595),
    .I1(n594)
  );
  //AND U374bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U374bar (
    .O(n596bar),
    .I0(n595bar),
    .I1(n594bar)
  );
  //OR U375
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U375 (
    .O(n594),
    .I0(in[135]),
    .I1(in[104])
  );
  //AND U375bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U375bar (
    .O(n594bar),
    .I0(inbar[135]),
    .I1(inbar[104])
  );
  //OR U376
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U376 (
    .O(n595),
    .I0(in[188]),
    .I1(in[178])
  );
  //AND U376bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U376bar (
    .O(n595bar),
    .I0(inbar[188]),
    .I1(inbar[178])
  );
  //OR U377
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U377 (
    .O(n597),
    .I0(n593),
    .I1(n592)
  );
  //AND U377bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U377bar (
    .O(n597bar),
    .I0(n593bar),
    .I1(n592bar)
  );
  //OR U378
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U378 (
    .O(n592),
    .I0(in[217]),
    .I1(in[194])
  );
  //AND U378bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U378bar (
    .O(n592bar),
    .I0(inbar[217]),
    .I1(inbar[194])
  );
  //OR U379
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U379 (
    .O(n593),
    .I0(in[237]),
    .I1(in[218])
  );
  //AND U379bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U379bar (
    .O(n593bar),
    .I0(inbar[237]),
    .I1(inbar[218])
  );
  //OR U380
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U380 (
    .O(n599),
    .I0(n591),
    .I1(n590)
  );
  //AND U380bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U380bar (
    .O(n599bar),
    .I0(n591bar),
    .I1(n590bar)
  );
  //OR U381
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U381 (
    .O(n590),
    .I0(n589),
    .I1(n588)
  );
  //AND U381bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U381bar (
    .O(n590bar),
    .I0(n589bar),
    .I1(n588bar)
  );
  //OR U382
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U382 (
    .O(n588),
    .I0(in_2),
    .I1(in_10)
  );
  //AND U382bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U382bar (
    .O(n588bar),
    .I0(in_2bar),
    .I1(in_10bar)
  );
  //OR U383
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U383 (
    .O(n589),
    .I0(in_47),
    .I1(in_22)
  );
  //AND U383bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U383bar (
    .O(n589bar),
    .I0(in_47bar),
    .I1(in_22bar)
  );
  //OR U384
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U384 (
    .O(n591),
    .I0(n587),
    .I1(n586)
  );
  //AND U384bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U384bar (
    .O(n591bar),
    .I0(n587bar),
    .I1(n586bar)
  );
  //OR U385
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U385 (
    .O(n586),
    .I0(in_56),
    .I1(in_54)
  );
  //AND U385bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U385bar (
    .O(n586bar),
    .I0(in_56bar),
    .I1(in_54bar)
  );
  //OR U386
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U386 (
    .O(n587),
    .I0(in_63),
    .I1(in_61)
  );
  //AND U386bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U386bar (
    .O(n587bar),
    .I0(in_63bar),
    .I1(in_61bar)
  );
  //OR U387
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U387 (
    .O(n820),
    .I0(n585),
    .I1(n584)
  );
  //AND U387bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U387bar (
    .O(n820bar),
    .I0(n585bar),
    .I1(n584bar)
  );
  //OR U388
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U388 (
    .O(n584),
    .I0(n583),
    .I1(n582)
  );
  //AND U388bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U388bar (
    .O(n584bar),
    .I0(n583bar),
    .I1(n582bar)
  );
  //OR U389
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U389 (
    .O(n582),
    .I0(n581),
    .I1(n580)
  );
  //AND U389bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U389bar (
    .O(n582bar),
    .I0(n581bar),
    .I1(n580bar)
  );
  //OR U390
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U390 (
    .O(n580),
    .I0(in[158]),
    .I1(in[142])
  );
  //AND U390bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U390bar (
    .O(n580bar),
    .I0(inbar[158]),
    .I1(inbar[142])
  );
  //OR U391
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U391 (
    .O(n581),
    .I0(in[175]),
    .I1(in[164])
  );
  //AND U391bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U391bar (
    .O(n581bar),
    .I0(inbar[175]),
    .I1(inbar[164])
  );
  //OR U392
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U392 (
    .O(n583),
    .I0(n579),
    .I1(n578)
  );
  //AND U392bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U392bar (
    .O(n583bar),
    .I0(n579bar),
    .I1(n578bar)
  );
  //OR U393
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U393 (
    .O(n578),
    .I0(in[228]),
    .I1(in[204])
  );
  //AND U393bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U393bar (
    .O(n578bar),
    .I0(inbar[228]),
    .I1(inbar[204])
  );
  //OR U394
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U394 (
    .O(n579),
    .I0(in[91]),
    .I1(in[87])
  );
  //AND U394bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U394bar (
    .O(n579bar),
    .I0(inbar[91]),
    .I1(inbar[87])
  );
  //OR U395
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U395 (
    .O(n585),
    .I0(n577),
    .I1(n576)
  );
  //AND U395bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U395bar (
    .O(n585bar),
    .I0(n577bar),
    .I1(n576bar)
  );
  //OR U396
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U396 (
    .O(n576),
    .I0(n575),
    .I1(n574)
  );
  //AND U396bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U396bar (
    .O(n576bar),
    .I0(n575bar),
    .I1(n574bar)
  );
  //OR U397
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U397 (
    .O(n574),
    .I0(in_21),
    .I1(in_11)
  );
  //AND U397bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U397bar (
    .O(n574bar),
    .I0(in_21bar),
    .I1(in_11bar)
  );
  //OR U398
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U398 (
    .O(n575),
    .I0(in_5),
    .I1(in_3)
  );
  //AND U398bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U398bar (
    .O(n575bar),
    .I0(in_5bar),
    .I1(in_3bar)
  );
  //OR U399
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U399 (
    .O(n577),
    .I0(n573),
    .I1(n572)
  );
  //AND U399bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U399bar (
    .O(n577bar),
    .I0(n573bar),
    .I1(n572bar)
  );
  //OR U400
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U400 (
    .O(n572),
    .I0(in_68),
    .I1(in_64)
  );
  //AND U400bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U400bar (
    .O(n572bar),
    .I0(in_68bar),
    .I1(in_64bar)
  );
  //OR U401
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U401 (
    .O(n573),
    .I0(in_76),
    .I1(in_73)
  );
  //AND U401bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U401bar (
    .O(n573bar),
    .I0(in_76bar),
    .I1(in_73bar)
  );
  //OR U402
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U402 (
    .O(n601),
    .I0(n778),
    .I1(n571)
  );
  //AND U402bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U402bar (
    .O(n601bar),
    .I0(n778bar),
    .I1(n571bar)
  );
  //OR U403
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U403 (
    .O(n571),
    .I0(in[100]),
    .I1(n965)
  );
  //AND U403bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U403bar (
    .O(n571bar),
    .I0(inbar[100]),
    .I1(n965bar)
  );
  //OR U404
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U404 (
    .O(n965),
    .I0(n570),
    .I1(n569)
  );
  //AND U404bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U404bar (
    .O(n965bar),
    .I0(n570bar),
    .I1(n569bar)
  );
  //OR U405
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U405 (
    .O(n569),
    .I0(n568),
    .I1(n567)
  );
  //AND U405bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U405bar (
    .O(n569bar),
    .I0(n568bar),
    .I1(n567bar)
  );
  //OR U406
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U406 (
    .O(n567),
    .I0(n566),
    .I1(n565)
  );
  //AND U406bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U406bar (
    .O(n567bar),
    .I0(n566bar),
    .I1(n565bar)
  );
  //OR U407
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U407 (
    .O(n565),
    .I0(n817),
    .I1(n750)
  );
  //AND U407bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U407bar (
    .O(n565bar),
    .I0(n817bar),
    .I1(n750bar)
  );
  //OR U408
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U408 (
    .O(n750),
    .I0(n564),
    .I1(n563)
  );
  //AND U408bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U408bar (
    .O(n750bar),
    .I0(n564bar),
    .I1(n563bar)
  );
  //OR U409
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U409 (
    .O(n563),
    .I0(n562),
    .I1(n561)
  );
  //AND U409bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U409bar (
    .O(n563bar),
    .I0(n562bar),
    .I1(n561bar)
  );
  //OR U410
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U410 (
    .O(n561),
    .I0(n560),
    .I1(n559)
  );
  //AND U410bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U410bar (
    .O(n561bar),
    .I0(n560bar),
    .I1(n559bar)
  );
  //OR U411
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U411 (
    .O(n559),
    .I0(in[119]),
    .I1(in[103])
  );
  //AND U411bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U411bar (
    .O(n559bar),
    .I0(inbar[119]),
    .I1(inbar[103])
  );
  //OR U412
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U412 (
    .O(n560),
    .I0(in[137]),
    .I1(in[133])
  );
  //AND U412bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U412bar (
    .O(n560bar),
    .I0(inbar[137]),
    .I1(inbar[133])
  );
  //OR U413
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U413 (
    .O(n562),
    .I0(n558),
    .I1(n557)
  );
  //AND U413bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U413bar (
    .O(n562bar),
    .I0(n558bar),
    .I1(n557bar)
  );
  //OR U414
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U414 (
    .O(n557),
    .I0(in[176]),
    .I1(in[173])
  );
  //AND U414bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U414bar (
    .O(n557bar),
    .I0(inbar[176]),
    .I1(inbar[173])
  );
  //OR U415
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U415 (
    .O(n558),
    .I0(in[210]),
    .I1(in[181])
  );
  //AND U415bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U415bar (
    .O(n558bar),
    .I0(inbar[210]),
    .I1(inbar[181])
  );
  //OR U416
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U416 (
    .O(n564),
    .I0(n556),
    .I1(n555)
  );
  //AND U416bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U416bar (
    .O(n564bar),
    .I0(n556bar),
    .I1(n555bar)
  );
  //OR U417
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U417 (
    .O(n555),
    .I0(n554),
    .I1(n553)
  );
  //AND U417bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U417bar (
    .O(n555bar),
    .I0(n554bar),
    .I1(n553bar)
  );
  //OR U418
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U418 (
    .O(n553),
    .I0(in_13),
    .I1(in[234])
  );
  //AND U418bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U418bar (
    .O(n553bar),
    .I0(in_13bar),
    .I1(inbar[234])
  );
  //OR U419
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U419 (
    .O(n554),
    .I0(in_38),
    .I1(in_32)
  );
  //AND U419bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U419bar (
    .O(n554bar),
    .I0(in_38bar),
    .I1(in_32bar)
  );
  //OR U420
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U420 (
    .O(n556),
    .I0(n552),
    .I1(n551)
  );
  //AND U420bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U420bar (
    .O(n556bar),
    .I0(n552bar),
    .I1(n551bar)
  );
  //OR U421
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U421 (
    .O(n551),
    .I0(in_42),
    .I1(in_41)
  );
  //AND U421bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U421bar (
    .O(n551bar),
    .I0(in_42bar),
    .I1(in_41bar)
  );
  //OR U422
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U422 (
    .O(n552),
    .I0(in_7),
    .I1(in_49)
  );
  //AND U422bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U422bar (
    .O(n552bar),
    .I0(in_7bar),
    .I1(in_49bar)
  );
  //OR U423
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U423 (
    .O(n817),
    .I0(n550),
    .I1(n549)
  );
  //AND U423bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U423bar (
    .O(n817bar),
    .I0(n550bar),
    .I1(n549bar)
  );
  //OR U424
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U424 (
    .O(n549),
    .I0(n548),
    .I1(n547)
  );
  //AND U424bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U424bar (
    .O(n549bar),
    .I0(n548bar),
    .I1(n547bar)
  );
  //OR U425
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U425 (
    .O(n547),
    .I0(n546),
    .I1(n545)
  );
  //AND U425bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U425bar (
    .O(n547bar),
    .I0(n546bar),
    .I1(n545bar)
  );
  //OR U426
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U426 (
    .O(n545),
    .I0(in[159]),
    .I1(in[105])
  );
  //AND U426bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U426bar (
    .O(n545bar),
    .I0(inbar[159]),
    .I1(inbar[105])
  );
  //OR U427
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U427 (
    .O(n546),
    .I0(in[206]),
    .I1(in[183])
  );
  //AND U427bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U427bar (
    .O(n546bar),
    .I0(inbar[206]),
    .I1(inbar[183])
  );
  //OR U428
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U428 (
    .O(n548),
    .I0(n544),
    .I1(n543)
  );
  //AND U428bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U428bar (
    .O(n548bar),
    .I0(n544bar),
    .I1(n543bar)
  );
  //OR U429
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U429 (
    .O(n543),
    .I0(in[229]),
    .I1(in[219])
  );
  //AND U429bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U429bar (
    .O(n543bar),
    .I0(inbar[229]),
    .I1(inbar[219])
  );
  //OR U430
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U430 (
    .O(n544),
    .I0(in[235]),
    .I1(in[232])
  );
  //AND U430bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U430bar (
    .O(n544bar),
    .I0(inbar[235]),
    .I1(inbar[232])
  );
  //OR U431
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U431 (
    .O(n550),
    .I0(n542),
    .I1(n541)
  );
  //AND U431bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U431bar (
    .O(n550bar),
    .I0(n542bar),
    .I1(n541bar)
  );
  //OR U432
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U432 (
    .O(n541),
    .I0(n540),
    .I1(n539)
  );
  //AND U432bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U432bar (
    .O(n541bar),
    .I0(n540bar),
    .I1(n539bar)
  );
  //OR U433
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U433 (
    .O(n539),
    .I0(in[249]),
    .I1(in[242])
  );
  //AND U433bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U433bar (
    .O(n539bar),
    .I0(inbar[249]),
    .I1(inbar[242])
  );
  //OR U434
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U434 (
    .O(n540),
    .I0(in[89]),
    .I1(in[254])
  );
  //AND U434bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U434bar (
    .O(n540bar),
    .I0(inbar[89]),
    .I1(inbar[254])
  );
  //OR U435
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U435 (
    .O(n542),
    .I0(n538),
    .I1(n537)
  );
  //AND U435bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U435bar (
    .O(n542bar),
    .I0(n538bar),
    .I1(n537bar)
  );
  //OR U436
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U436 (
    .O(n537),
    .I0(in_14),
    .I1(in[99])
  );
  //AND U436bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U436bar (
    .O(n537bar),
    .I0(in_14bar),
    .I1(inbar[99])
  );
  //OR U437
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U437 (
    .O(n538),
    .I0(in_60),
    .I1(in_18)
  );
  //AND U437bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U437bar (
    .O(n538bar),
    .I0(in_60bar),
    .I1(in_18bar)
  );
  //OR U438
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U438 (
    .O(n566),
    .I0(in[113]),
    .I1(n763)
  );
  //AND U438bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U438bar (
    .O(n566bar),
    .I0(inbar[113]),
    .I1(n763bar)
  );
  //OR U439
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U439 (
    .O(n763),
    .I0(n536),
    .I1(n535)
  );
  //AND U439bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U439bar (
    .O(n763bar),
    .I0(n536bar),
    .I1(n535bar)
  );
  //OR U440
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U440 (
    .O(n535),
    .I0(n534),
    .I1(n533)
  );
  //AND U440bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U440bar (
    .O(n535bar),
    .I0(n534bar),
    .I1(n533bar)
  );
  //OR U441
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U441 (
    .O(n533),
    .I0(n532),
    .I1(n531)
  );
  //AND U441bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U441bar (
    .O(n533bar),
    .I0(n532bar),
    .I1(n531bar)
  );
  //OR U442
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U442 (
    .O(n531),
    .I0(in[115]),
    .I1(in[110])
  );
  //AND U442bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U442bar (
    .O(n531bar),
    .I0(inbar[115]),
    .I1(inbar[110])
  );
  //OR U443
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U443 (
    .O(n532),
    .I0(in[125]),
    .I1(in[117])
  );
  //AND U443bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U443bar (
    .O(n532bar),
    .I0(inbar[125]),
    .I1(inbar[117])
  );
  //OR U444
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U444 (
    .O(n534),
    .I0(n530),
    .I1(n529)
  );
  //AND U444bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U444bar (
    .O(n534bar),
    .I0(n530bar),
    .I1(n529bar)
  );
  //OR U445
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U445 (
    .O(n529),
    .I0(in[180]),
    .I1(in[128])
  );
  //AND U445bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U445bar (
    .O(n529bar),
    .I0(inbar[180]),
    .I1(inbar[128])
  );
  //OR U446
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U446 (
    .O(n530),
    .I0(in[205]),
    .I1(in[201])
  );
  //AND U446bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U446bar (
    .O(n530bar),
    .I0(inbar[205]),
    .I1(inbar[201])
  );
  //OR U447
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U447 (
    .O(n536),
    .I0(n528),
    .I1(n527)
  );
  //AND U447bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U447bar (
    .O(n536bar),
    .I0(n528bar),
    .I1(n527bar)
  );
  //OR U448
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U448 (
    .O(n527),
    .I0(n526),
    .I1(n525)
  );
  //AND U448bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U448bar (
    .O(n527bar),
    .I0(n526bar),
    .I1(n525bar)
  );
  //OR U449
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U449 (
    .O(n525),
    .I0(in[244]),
    .I1(in[239])
  );
  //AND U449bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U449bar (
    .O(n525bar),
    .I0(inbar[244]),
    .I1(inbar[239])
  );
  //OR U450
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U450 (
    .O(n526),
    .I0(in[95]),
    .I1(in[83])
  );
  //AND U450bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U450bar (
    .O(n526bar),
    .I0(inbar[95]),
    .I1(inbar[83])
  );
  //OR U451
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U451 (
    .O(n528),
    .I0(n524),
    .I1(n523)
  );
  //AND U451bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U451bar (
    .O(n528bar),
    .I0(n524bar),
    .I1(n523bar)
  );
  //OR U452
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U452 (
    .O(n523),
    .I0(in_24),
    .I1(in[97])
  );
  //AND U452bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U452bar (
    .O(n523bar),
    .I0(in_24bar),
    .I1(inbar[97])
  );
  //OR U453
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U453 (
    .O(n524),
    .I0(in_33),
    .I1(in_27)
  );
  //AND U453bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U453bar (
    .O(n524bar),
    .I0(in_33bar),
    .I1(in_27bar)
  );
  //OR U454
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U454 (
    .O(n568),
    .I0(n522),
    .I1(n521)
  );
  //AND U454bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U454bar (
    .O(n568bar),
    .I0(n522bar),
    .I1(n521bar)
  );
  //OR U455
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U455 (
    .O(n521),
    .I0(in[145]),
    .I1(in[126])
  );
  //AND U455bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U455bar (
    .O(n521bar),
    .I0(inbar[145]),
    .I1(inbar[126])
  );
  //OR U456
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U456 (
    .O(n522),
    .I0(in[169]),
    .I1(n520)
  );
  //AND U456bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U456bar (
    .O(n522bar),
    .I0(inbar[169]),
    .I1(n520bar)
  );
  //OR U457
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U457 (
    .O(n520),
    .I0(in[221]),
    .I1(in[172])
  );
  //AND U457bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U457bar (
    .O(n520bar),
    .I0(inbar[221]),
    .I1(inbar[172])
  );
  //OR U458
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U458 (
    .O(n570),
    .I0(n519),
    .I1(n518)
  );
  //AND U458bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U458bar (
    .O(n570bar),
    .I0(n519bar),
    .I1(n518bar)
  );
  //OR U459
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U459 (
    .O(n518),
    .I0(n517),
    .I1(n516)
  );
  //AND U459bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U459bar (
    .O(n518bar),
    .I0(n517bar),
    .I1(n516bar)
  );
  //OR U460
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U460 (
    .O(n516),
    .I0(in[241]),
    .I1(in[224])
  );
  //AND U460bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U460bar (
    .O(n516bar),
    .I0(inbar[241]),
    .I1(inbar[224])
  );
  //OR U461
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U461 (
    .O(n517),
    .I0(in[86]),
    .I1(n515)
  );
  //AND U461bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U461bar (
    .O(n517bar),
    .I0(inbar[86]),
    .I1(n515bar)
  );
  //OR U462
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U462 (
    .O(n515),
    .I0(in_43),
    .I1(in_34)
  );
  //AND U462bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U462bar (
    .O(n515bar),
    .I0(in_43bar),
    .I1(in_34bar)
  );
  //OR U463
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U463 (
    .O(n519),
    .I0(n514),
    .I1(n513)
  );
  //AND U463bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U463bar (
    .O(n519bar),
    .I0(n514bar),
    .I1(n513bar)
  );
  //OR U464
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U464 (
    .O(n513),
    .I0(in_65),
    .I1(in_51)
  );
  //AND U464bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U464bar (
    .O(n513bar),
    .I0(in_65bar),
    .I1(in_51bar)
  );
  //OR U465
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U465 (
    .O(n514),
    .I0(in_75),
    .I1(n512)
  );
  //AND U465bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U465bar (
    .O(n514bar),
    .I0(in_75bar),
    .I1(n512bar)
  );
  //OR U466
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U466 (
    .O(n512),
    .I0(in_81),
    .I1(in_77)
  );
  //AND U466bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U466bar (
    .O(n512bar),
    .I0(in_81bar),
    .I1(in_77bar)
  );
  //OR U467
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U467 (
    .O(n778),
    .I0(n511),
    .I1(n510)
  );
  //AND U467bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U467bar (
    .O(n778bar),
    .I0(n511bar),
    .I1(n510bar)
  );
  //OR U468
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U468 (
    .O(n510),
    .I0(n509),
    .I1(n508)
  );
  //AND U468bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U468bar (
    .O(n510bar),
    .I0(n509bar),
    .I1(n508bar)
  );
  //OR U469
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U469 (
    .O(n508),
    .I0(n507),
    .I1(n506)
  );
  //AND U469bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U469bar (
    .O(n508bar),
    .I0(n507bar),
    .I1(n506bar)
  );
  //OR U470
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U470 (
    .O(n506),
    .I0(in[107]),
    .I1(in[101])
  );
  //AND U470bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U470bar (
    .O(n506bar),
    .I0(inbar[107]),
    .I1(inbar[101])
  );
  //OR U471
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U471 (
    .O(n507),
    .I0(in[139]),
    .I1(in[132])
  );
  //AND U471bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U471bar (
    .O(n507bar),
    .I0(inbar[139]),
    .I1(inbar[132])
  );
  //OR U472
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U472 (
    .O(n509),
    .I0(n505),
    .I1(n504)
  );
  //AND U472bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U472bar (
    .O(n509bar),
    .I0(n505bar),
    .I1(n504bar)
  );
  //OR U473
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U473 (
    .O(n504),
    .I0(in[146]),
    .I1(in[141])
  );
  //AND U473bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U473bar (
    .O(n504bar),
    .I0(inbar[146]),
    .I1(inbar[141])
  );
  //OR U474
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U474 (
    .O(n505),
    .I0(in[203]),
    .I1(in[179])
  );
  //AND U474bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U474bar (
    .O(n505bar),
    .I0(inbar[203]),
    .I1(inbar[179])
  );
  //OR U475
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U475 (
    .O(n511),
    .I0(n503),
    .I1(n502)
  );
  //AND U475bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U475bar (
    .O(n511bar),
    .I0(n503bar),
    .I1(n502bar)
  );
  //OR U476
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U476 (
    .O(n502),
    .I0(n501),
    .I1(n500)
  );
  //AND U476bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U476bar (
    .O(n502bar),
    .I0(n501bar),
    .I1(n500bar)
  );
  //OR U477
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U477 (
    .O(n500),
    .I0(in[243]),
    .I1(in[222])
  );
  //AND U477bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U477bar (
    .O(n500bar),
    .I0(inbar[243]),
    .I1(inbar[222])
  );
  //OR U478
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U478 (
    .O(n501),
    .I0(in[251]),
    .I1(in[250])
  );
  //AND U478bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U478bar (
    .O(n501bar),
    .I0(inbar[251]),
    .I1(inbar[250])
  );
  //OR U479
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U479 (
    .O(n503),
    .I0(n499),
    .I1(n498)
  );
  //AND U479bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U479bar (
    .O(n503bar),
    .I0(n499bar),
    .I1(n498bar)
  );
  //OR U480
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U480 (
    .O(n498),
    .I0(in_37),
    .I1(in_19)
  );
  //AND U480bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U480bar (
    .O(n498bar),
    .I0(in_37bar),
    .I1(in_19bar)
  );
  //OR U481
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U481 (
    .O(n499),
    .I0(in_78),
    .I1(in_6)
  );
  //AND U481bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U481bar (
    .O(n499bar),
    .I0(in_78bar),
    .I1(in_6bar)
  );
  //OR U482
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U482 (
    .O(n603),
    .I0(n497),
    .I1(n496)
  );
  //AND U482bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U482bar (
    .O(n603bar),
    .I0(n497bar),
    .I1(n496bar)
  );
  //OR U483
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U483 (
    .O(n496),
    .I0(in[112]),
    .I1(in[102])
  );
  //AND U483bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U483bar (
    .O(n496bar),
    .I0(inbar[112]),
    .I1(inbar[102])
  );
  //OR U484
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U484 (
    .O(n497),
    .I0(in[123]),
    .I1(n495)
  );
  //AND U484bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U484bar (
    .O(n497bar),
    .I0(inbar[123]),
    .I1(n495bar)
  );
  //OR U485
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U485 (
    .O(n495),
    .I0(in[143]),
    .I1(in[130])
  );
  //AND U485bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U485bar (
    .O(n495bar),
    .I0(inbar[143]),
    .I1(inbar[130])
  );
  //OR U486
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U486 (
    .O(n605),
    .I0(n494),
    .I1(n493)
  );
  //AND U486bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U486bar (
    .O(n605bar),
    .I0(n494bar),
    .I1(n493bar)
  );
  //OR U487
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U487 (
    .O(n493),
    .I0(n492),
    .I1(n491)
  );
  //AND U487bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U487bar (
    .O(n493bar),
    .I0(n492bar),
    .I1(n491bar)
  );
  //OR U488
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U488 (
    .O(n491),
    .I0(in[216]),
    .I1(in[213])
  );
  //AND U488bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U488bar (
    .O(n491bar),
    .I0(inbar[216]),
    .I1(inbar[213])
  );
  //OR U489
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U489 (
    .O(n492),
    .I0(in[227]),
    .I1(n490)
  );
  //AND U489bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U489bar (
    .O(n492bar),
    .I0(inbar[227]),
    .I1(n490bar)
  );
  //OR U490
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U490 (
    .O(n490),
    .I0(in_0),
    .I1(in[248])
  );
  //AND U490bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U490bar (
    .O(n490bar),
    .I0(in_0bar),
    .I1(inbar[248])
  );
  //OR U491
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U491 (
    .O(n494),
    .I0(n489),
    .I1(n488)
  );
  //AND U491bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U491bar (
    .O(n494bar),
    .I0(n489bar),
    .I1(n488bar)
  );
  //OR U492
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U492 (
    .O(n488),
    .I0(in_46),
    .I1(in_44)
  );
  //AND U492bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U492bar (
    .O(n488bar),
    .I0(in_46bar),
    .I1(in_44bar)
  );
  //OR U493
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U493 (
    .O(n489),
    .I0(in_50),
    .I1(n487)
  );
  //AND U493bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U493bar (
    .O(n489bar),
    .I0(in_50bar),
    .I1(n487bar)
  );
  //OR U494
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U494 (
    .O(n487),
    .I0(in_9),
    .I1(in_80)
  );
  //AND U494bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U494bar (
    .O(n487bar),
    .I0(in_9bar),
    .I1(in_80bar)
  );
endmodule

module sBox_10 ( in, out );

  input wire [7:0] in;
//input_done

  output wire [7:0] out;
//output_done

  wire [255:0] decodeOut;
//wire_done

  decode_10 dec ( .in(in), .out(decodeOut) );
  encode_10 enc ( .in(decodeOut), .out(out) );
endmodule

module CD2_41 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD2_42 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD2_43 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD2_44 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD4_21 ( a, b, y );

  input wire [3:0] a;
  input wire [3:0] b;
  wire [3:0] abar;
  wire [3:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
//input_done

  output wire [15:0] y;
  wire [15:0] ybar;
//output_done

//wire_done

  //AND U1
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1 (
    .O(y[9]),
    .I0(b[1]),
    .I1(a[2])
  );
  //OR U1bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1bar (
    .O(ybar[9]),
    .I0(bbar[1]),
    .I1(abar[2])
  );
  //AND U2
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2 (
    .O(y[8]),
    .I0(b[0]),
    .I1(a[2])
  );
  //OR U2bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2bar (
    .O(ybar[8]),
    .I0(bbar[0]),
    .I1(abar[2])
  );
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[7]),
    .I0(b[3]),
    .I1(a[1])
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[7]),
    .I0(bbar[3]),
    .I1(abar[1])
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[6]),
    .I0(b[2]),
    .I1(a[1])
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[6]),
    .I0(bbar[2]),
    .I1(abar[1])
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[5]),
    .I0(a[1]),
    .I1(b[1])
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[5]),
    .I0(abar[1]),
    .I1(bbar[1])
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[4]),
    .I0(a[1]),
    .I1(b[0])
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[4]),
    .I0(abar[1]),
    .I1(bbar[0])
  );
  //AND U7
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7 (
    .O(y[3]),
    .I0(a[0]),
    .I1(b[3])
  );
  //OR U7bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7bar (
    .O(ybar[3]),
    .I0(abar[0]),
    .I1(bbar[3])
  );
  //AND U8
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8 (
    .O(y[2]),
    .I0(a[0]),
    .I1(b[2])
  );
  //OR U8bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8bar (
    .O(ybar[2]),
    .I0(abar[0]),
    .I1(bbar[2])
  );
  //AND U9
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9 (
    .O(y[1]),
    .I0(a[0]),
    .I1(b[1])
  );
  //OR U9bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9bar (
    .O(ybar[1]),
    .I0(abar[0]),
    .I1(bbar[1])
  );
  //AND U10
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10 (
    .O(y[15]),
    .I0(a[3]),
    .I1(b[3])
  );
  //OR U10bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10bar (
    .O(ybar[15]),
    .I0(abar[3]),
    .I1(bbar[3])
  );
  //AND U11
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11 (
    .O(y[14]),
    .I0(a[3]),
    .I1(b[2])
  );
  //OR U11bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11bar (
    .O(ybar[14]),
    .I0(abar[3]),
    .I1(bbar[2])
  );
  //AND U12
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12 (
    .O(y[13]),
    .I0(a[3]),
    .I1(b[1])
  );
  //OR U12bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12bar (
    .O(ybar[13]),
    .I0(abar[3]),
    .I1(bbar[1])
  );
  //AND U13
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13 (
    .O(y[12]),
    .I0(a[3]),
    .I1(b[0])
  );
  //OR U13bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13bar (
    .O(ybar[12]),
    .I0(abar[3]),
    .I1(bbar[0])
  );
  //AND U14
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14 (
    .O(y[11]),
    .I0(b[3]),
    .I1(a[2])
  );
  //OR U14bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14bar (
    .O(ybar[11]),
    .I0(bbar[3]),
    .I1(abar[2])
  );
  //AND U15
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15 (
    .O(y[10]),
    .I0(b[2]),
    .I1(a[2])
  );
  //OR U15bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15bar (
    .O(ybar[10]),
    .I0(bbar[2]),
    .I1(abar[2])
  );
  //AND U16
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16 (
    .O(y[0]),
    .I0(a[0]),
    .I1(b[0])
  );
  //OR U16bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16bar (
    .O(ybar[0]),
    .I0(abar[0]),
    .I1(bbar[0])
  );
endmodule

module CD4_22 ( a, b, y );

  input wire [3:0] a;
  input wire [3:0] b;
  wire [3:0] abar;
  wire [3:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
//input_done

  output wire [15:0] y;
  wire [15:0] ybar;
//output_done

//wire_done

  //AND U1
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1 (
    .O(y[9]),
    .I0(b[1]),
    .I1(a[2])
  );
  //OR U1bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1bar (
    .O(ybar[9]),
    .I0(bbar[1]),
    .I1(abar[2])
  );
  //AND U2
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2 (
    .O(y[8]),
    .I0(b[0]),
    .I1(a[2])
  );
  //OR U2bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2bar (
    .O(ybar[8]),
    .I0(bbar[0]),
    .I1(abar[2])
  );
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[7]),
    .I0(b[3]),
    .I1(a[1])
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[7]),
    .I0(bbar[3]),
    .I1(abar[1])
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[6]),
    .I0(b[2]),
    .I1(a[1])
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[6]),
    .I0(bbar[2]),
    .I1(abar[1])
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[5]),
    .I0(a[1]),
    .I1(b[1])
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[5]),
    .I0(abar[1]),
    .I1(bbar[1])
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[4]),
    .I0(a[1]),
    .I1(b[0])
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[4]),
    .I0(abar[1]),
    .I1(bbar[0])
  );
  //AND U7
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7 (
    .O(y[3]),
    .I0(a[0]),
    .I1(b[3])
  );
  //OR U7bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7bar (
    .O(ybar[3]),
    .I0(abar[0]),
    .I1(bbar[3])
  );
  //AND U8
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8 (
    .O(y[2]),
    .I0(a[0]),
    .I1(b[2])
  );
  //OR U8bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8bar (
    .O(ybar[2]),
    .I0(abar[0]),
    .I1(bbar[2])
  );
  //AND U9
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9 (
    .O(y[1]),
    .I0(a[0]),
    .I1(b[1])
  );
  //OR U9bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9bar (
    .O(ybar[1]),
    .I0(abar[0]),
    .I1(bbar[1])
  );
  //AND U10
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10 (
    .O(y[15]),
    .I0(a[3]),
    .I1(b[3])
  );
  //OR U10bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10bar (
    .O(ybar[15]),
    .I0(abar[3]),
    .I1(bbar[3])
  );
  //AND U11
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11 (
    .O(y[14]),
    .I0(a[3]),
    .I1(b[2])
  );
  //OR U11bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11bar (
    .O(ybar[14]),
    .I0(abar[3]),
    .I1(bbar[2])
  );
  //AND U12
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12 (
    .O(y[13]),
    .I0(a[3]),
    .I1(b[1])
  );
  //OR U12bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12bar (
    .O(ybar[13]),
    .I0(abar[3]),
    .I1(bbar[1])
  );
  //AND U13
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13 (
    .O(y[12]),
    .I0(a[3]),
    .I1(b[0])
  );
  //OR U13bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13bar (
    .O(ybar[12]),
    .I0(abar[3]),
    .I1(bbar[0])
  );
  //AND U14
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14 (
    .O(y[11]),
    .I0(b[3]),
    .I1(a[2])
  );
  //OR U14bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14bar (
    .O(ybar[11]),
    .I0(bbar[3]),
    .I1(abar[2])
  );
  //AND U15
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15 (
    .O(y[10]),
    .I0(b[2]),
    .I1(a[2])
  );
  //OR U15bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15bar (
    .O(ybar[10]),
    .I0(bbar[2]),
    .I1(abar[2])
  );
  //AND U16
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16 (
    .O(y[0]),
    .I0(a[0]),
    .I1(b[0])
  );
  //OR U16bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16bar (
    .O(ybar[0]),
    .I0(abar[0]),
    .I1(bbar[0])
  );
endmodule

module CD16_11 ( a, b, y );

  input wire [15:0] a;
  input wire [15:0] b;
  wire [15:0] abar;
  wire [15:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign abar[8] = ~a[8];
  assign abar[9] = ~a[9];
  assign abar[10] = ~a[10];
  assign abar[11] = ~a[11];
  assign abar[12] = ~a[12];
  assign abar[13] = ~a[13];
  assign abar[14] = ~a[14];
  assign abar[15] = ~a[15];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign bbar[8] = ~b[8];
  assign bbar[9] = ~b[9];
  assign bbar[10] = ~b[10];
  assign bbar[11] = ~b[11];
  assign bbar[12] = ~b[12];
  assign bbar[13] = ~b[13];
  assign bbar[14] = ~b[14];
  assign bbar[15] = ~b[15];
//input_done

  output wire [255:0] y;
  wire [255:0] ybar;
//output_done

//wire_done

  //AND U1
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1 (
    .O(y[9]),
    .I0(b[9]),
    .I1(a[0])
  );
  //OR U1bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1bar (
    .O(ybar[9]),
    .I0(bbar[9]),
    .I1(abar[0])
  );
  //AND U2
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2 (
    .O(y[99]),
    .I0(b[3]),
    .I1(a[6])
  );
  //OR U2bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2bar (
    .O(ybar[99]),
    .I0(bbar[3]),
    .I1(abar[6])
  );
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[98]),
    .I0(b[2]),
    .I1(a[6])
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[98]),
    .I0(bbar[2]),
    .I1(abar[6])
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[97]),
    .I0(b[1]),
    .I1(a[6])
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[97]),
    .I0(bbar[1]),
    .I1(abar[6])
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[96]),
    .I0(b[0]),
    .I1(a[6])
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[96]),
    .I0(bbar[0]),
    .I1(abar[6])
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[95]),
    .I0(b[15]),
    .I1(a[5])
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[95]),
    .I0(bbar[15]),
    .I1(abar[5])
  );
  //AND U7
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7 (
    .O(y[94]),
    .I0(b[14]),
    .I1(a[5])
  );
  //OR U7bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7bar (
    .O(ybar[94]),
    .I0(bbar[14]),
    .I1(abar[5])
  );
  //AND U8
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8 (
    .O(y[93]),
    .I0(b[13]),
    .I1(a[5])
  );
  //OR U8bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8bar (
    .O(ybar[93]),
    .I0(bbar[13]),
    .I1(abar[5])
  );
  //AND U9
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9 (
    .O(y[92]),
    .I0(b[12]),
    .I1(a[5])
  );
  //OR U9bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9bar (
    .O(ybar[92]),
    .I0(bbar[12]),
    .I1(abar[5])
  );
  //AND U10
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10 (
    .O(y[91]),
    .I0(b[11]),
    .I1(a[5])
  );
  //OR U10bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10bar (
    .O(ybar[91]),
    .I0(bbar[11]),
    .I1(abar[5])
  );
  //AND U11
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11 (
    .O(y[90]),
    .I0(b[10]),
    .I1(a[5])
  );
  //OR U11bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11bar (
    .O(ybar[90]),
    .I0(bbar[10]),
    .I1(abar[5])
  );
  //AND U12
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12 (
    .O(y[8]),
    .I0(b[8]),
    .I1(a[0])
  );
  //OR U12bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12bar (
    .O(ybar[8]),
    .I0(bbar[8]),
    .I1(abar[0])
  );
  //AND U13
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13 (
    .O(y[89]),
    .I0(a[5]),
    .I1(b[9])
  );
  //OR U13bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13bar (
    .O(ybar[89]),
    .I0(abar[5]),
    .I1(bbar[9])
  );
  //AND U14
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14 (
    .O(y[88]),
    .I0(b[8]),
    .I1(a[5])
  );
  //OR U14bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14bar (
    .O(ybar[88]),
    .I0(bbar[8]),
    .I1(abar[5])
  );
  //AND U15
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15 (
    .O(y[87]),
    .I0(b[7]),
    .I1(a[5])
  );
  //OR U15bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15bar (
    .O(ybar[87]),
    .I0(bbar[7]),
    .I1(abar[5])
  );
  //AND U16
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16 (
    .O(y[86]),
    .I0(b[6]),
    .I1(a[5])
  );
  //OR U16bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16bar (
    .O(ybar[86]),
    .I0(bbar[6]),
    .I1(abar[5])
  );
  //AND U17
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U17 (
    .O(y[85]),
    .I0(b[5]),
    .I1(a[5])
  );
  //OR U17bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U17bar (
    .O(ybar[85]),
    .I0(bbar[5]),
    .I1(abar[5])
  );
  //AND U18
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U18 (
    .O(y[84]),
    .I0(b[4]),
    .I1(a[5])
  );
  //OR U18bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U18bar (
    .O(ybar[84]),
    .I0(bbar[4]),
    .I1(abar[5])
  );
  //AND U19
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U19 (
    .O(y[83]),
    .I0(a[5]),
    .I1(b[3])
  );
  //OR U19bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U19bar (
    .O(ybar[83]),
    .I0(abar[5]),
    .I1(bbar[3])
  );
  //AND U20
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U20 (
    .O(y[82]),
    .I0(a[5]),
    .I1(b[2])
  );
  //OR U20bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U20bar (
    .O(ybar[82]),
    .I0(abar[5]),
    .I1(bbar[2])
  );
  //AND U21
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U21 (
    .O(y[81]),
    .I0(a[5]),
    .I1(b[1])
  );
  //OR U21bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U21bar (
    .O(ybar[81]),
    .I0(abar[5]),
    .I1(bbar[1])
  );
  //AND U22
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U22 (
    .O(y[80]),
    .I0(a[5]),
    .I1(b[0])
  );
  //OR U22bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U22bar (
    .O(ybar[80]),
    .I0(abar[5]),
    .I1(bbar[0])
  );
  //AND U23
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U23 (
    .O(y[7]),
    .I0(b[7]),
    .I1(a[0])
  );
  //OR U23bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U23bar (
    .O(ybar[7]),
    .I0(bbar[7]),
    .I1(abar[0])
  );
  //AND U24
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U24 (
    .O(y[79]),
    .I0(a[4]),
    .I1(b[15])
  );
  //OR U24bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U24bar (
    .O(ybar[79]),
    .I0(abar[4]),
    .I1(bbar[15])
  );
  //AND U25
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U25 (
    .O(y[78]),
    .I0(a[4]),
    .I1(b[14])
  );
  //OR U25bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U25bar (
    .O(ybar[78]),
    .I0(abar[4]),
    .I1(bbar[14])
  );
  //AND U26
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U26 (
    .O(y[77]),
    .I0(a[4]),
    .I1(b[13])
  );
  //OR U26bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U26bar (
    .O(ybar[77]),
    .I0(abar[4]),
    .I1(bbar[13])
  );
  //AND U27
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U27 (
    .O(y[76]),
    .I0(a[4]),
    .I1(b[12])
  );
  //OR U27bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U27bar (
    .O(ybar[76]),
    .I0(abar[4]),
    .I1(bbar[12])
  );
  //AND U28
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U28 (
    .O(y[75]),
    .I0(a[4]),
    .I1(b[11])
  );
  //OR U28bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U28bar (
    .O(ybar[75]),
    .I0(abar[4]),
    .I1(bbar[11])
  );
  //AND U29
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U29 (
    .O(y[74]),
    .I0(a[4]),
    .I1(b[10])
  );
  //OR U29bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U29bar (
    .O(ybar[74]),
    .I0(abar[4]),
    .I1(bbar[10])
  );
  //AND U30
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U30 (
    .O(y[73]),
    .I0(a[4]),
    .I1(b[9])
  );
  //OR U30bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U30bar (
    .O(ybar[73]),
    .I0(abar[4]),
    .I1(bbar[9])
  );
  //AND U31
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U31 (
    .O(y[72]),
    .I0(a[4]),
    .I1(b[8])
  );
  //OR U31bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U31bar (
    .O(ybar[72]),
    .I0(abar[4]),
    .I1(bbar[8])
  );
  //AND U32
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U32 (
    .O(y[71]),
    .I0(a[4]),
    .I1(b[7])
  );
  //OR U32bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U32bar (
    .O(ybar[71]),
    .I0(abar[4]),
    .I1(bbar[7])
  );
  //AND U33
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U33 (
    .O(y[70]),
    .I0(a[4]),
    .I1(b[6])
  );
  //OR U33bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U33bar (
    .O(ybar[70]),
    .I0(abar[4]),
    .I1(bbar[6])
  );
  //AND U34
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U34 (
    .O(y[6]),
    .I0(b[6]),
    .I1(a[0])
  );
  //OR U34bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U34bar (
    .O(ybar[6]),
    .I0(bbar[6]),
    .I1(abar[0])
  );
  //AND U35
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U35 (
    .O(y[69]),
    .I0(a[4]),
    .I1(b[5])
  );
  //OR U35bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U35bar (
    .O(ybar[69]),
    .I0(abar[4]),
    .I1(bbar[5])
  );
  //AND U36
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U36 (
    .O(y[68]),
    .I0(a[4]),
    .I1(b[4])
  );
  //OR U36bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U36bar (
    .O(ybar[68]),
    .I0(abar[4]),
    .I1(bbar[4])
  );
  //AND U37
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U37 (
    .O(y[67]),
    .I0(a[4]),
    .I1(b[3])
  );
  //OR U37bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U37bar (
    .O(ybar[67]),
    .I0(abar[4]),
    .I1(bbar[3])
  );
  //AND U38
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U38 (
    .O(y[66]),
    .I0(a[4]),
    .I1(b[2])
  );
  //OR U38bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U38bar (
    .O(ybar[66]),
    .I0(abar[4]),
    .I1(bbar[2])
  );
  //AND U39
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U39 (
    .O(y[65]),
    .I0(a[4]),
    .I1(b[1])
  );
  //OR U39bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U39bar (
    .O(ybar[65]),
    .I0(abar[4]),
    .I1(bbar[1])
  );
  //AND U40
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U40 (
    .O(y[64]),
    .I0(a[4]),
    .I1(b[0])
  );
  //OR U40bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U40bar (
    .O(ybar[64]),
    .I0(abar[4]),
    .I1(bbar[0])
  );
  //AND U41
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U41 (
    .O(y[63]),
    .I0(a[3]),
    .I1(b[15])
  );
  //OR U41bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U41bar (
    .O(ybar[63]),
    .I0(abar[3]),
    .I1(bbar[15])
  );
  //AND U42
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U42 (
    .O(y[62]),
    .I0(a[3]),
    .I1(b[14])
  );
  //OR U42bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U42bar (
    .O(ybar[62]),
    .I0(abar[3]),
    .I1(bbar[14])
  );
  //AND U43
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U43 (
    .O(y[61]),
    .I0(a[3]),
    .I1(b[13])
  );
  //OR U43bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U43bar (
    .O(ybar[61]),
    .I0(abar[3]),
    .I1(bbar[13])
  );
  //AND U44
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U44 (
    .O(y[60]),
    .I0(a[3]),
    .I1(b[12])
  );
  //OR U44bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U44bar (
    .O(ybar[60]),
    .I0(abar[3]),
    .I1(bbar[12])
  );
  //AND U45
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U45 (
    .O(y[5]),
    .I0(b[5]),
    .I1(a[0])
  );
  //OR U45bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U45bar (
    .O(ybar[5]),
    .I0(bbar[5]),
    .I1(abar[0])
  );
  //AND U46
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U46 (
    .O(y[59]),
    .I0(a[3]),
    .I1(b[11])
  );
  //OR U46bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U46bar (
    .O(ybar[59]),
    .I0(abar[3]),
    .I1(bbar[11])
  );
  //AND U47
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U47 (
    .O(y[58]),
    .I0(a[3]),
    .I1(b[10])
  );
  //OR U47bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U47bar (
    .O(ybar[58]),
    .I0(abar[3]),
    .I1(bbar[10])
  );
  //AND U48
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U48 (
    .O(y[57]),
    .I0(a[3]),
    .I1(b[9])
  );
  //OR U48bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U48bar (
    .O(ybar[57]),
    .I0(abar[3]),
    .I1(bbar[9])
  );
  //AND U49
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U49 (
    .O(y[56]),
    .I0(a[3]),
    .I1(b[8])
  );
  //OR U49bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U49bar (
    .O(ybar[56]),
    .I0(abar[3]),
    .I1(bbar[8])
  );
  //AND U50
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U50 (
    .O(y[55]),
    .I0(a[3]),
    .I1(b[7])
  );
  //OR U50bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U50bar (
    .O(ybar[55]),
    .I0(abar[3]),
    .I1(bbar[7])
  );
  //AND U51
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U51 (
    .O(y[54]),
    .I0(a[3]),
    .I1(b[6])
  );
  //OR U51bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U51bar (
    .O(ybar[54]),
    .I0(abar[3]),
    .I1(bbar[6])
  );
  //AND U52
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U52 (
    .O(y[53]),
    .I0(a[3]),
    .I1(b[5])
  );
  //OR U52bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U52bar (
    .O(ybar[53]),
    .I0(abar[3]),
    .I1(bbar[5])
  );
  //AND U53
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U53 (
    .O(y[52]),
    .I0(a[3]),
    .I1(b[4])
  );
  //OR U53bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U53bar (
    .O(ybar[52]),
    .I0(abar[3]),
    .I1(bbar[4])
  );
  //AND U54
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U54 (
    .O(y[51]),
    .I0(a[3]),
    .I1(b[3])
  );
  //OR U54bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U54bar (
    .O(ybar[51]),
    .I0(abar[3]),
    .I1(bbar[3])
  );
  //AND U55
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U55 (
    .O(y[50]),
    .I0(a[3]),
    .I1(b[2])
  );
  //OR U55bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U55bar (
    .O(ybar[50]),
    .I0(abar[3]),
    .I1(bbar[2])
  );
  //AND U56
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U56 (
    .O(y[4]),
    .I0(b[4]),
    .I1(a[0])
  );
  //OR U56bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U56bar (
    .O(ybar[4]),
    .I0(bbar[4]),
    .I1(abar[0])
  );
  //AND U57
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U57 (
    .O(y[49]),
    .I0(a[3]),
    .I1(b[1])
  );
  //OR U57bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U57bar (
    .O(ybar[49]),
    .I0(abar[3]),
    .I1(bbar[1])
  );
  //AND U58
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U58 (
    .O(y[48]),
    .I0(a[3]),
    .I1(b[0])
  );
  //OR U58bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U58bar (
    .O(ybar[48]),
    .I0(abar[3]),
    .I1(bbar[0])
  );
  //AND U59
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U59 (
    .O(y[47]),
    .I0(a[2]),
    .I1(b[15])
  );
  //OR U59bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U59bar (
    .O(ybar[47]),
    .I0(abar[2]),
    .I1(bbar[15])
  );
  //AND U60
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U60 (
    .O(y[46]),
    .I0(a[2]),
    .I1(b[14])
  );
  //OR U60bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U60bar (
    .O(ybar[46]),
    .I0(abar[2]),
    .I1(bbar[14])
  );
  //AND U61
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U61 (
    .O(y[45]),
    .I0(a[2]),
    .I1(b[13])
  );
  //OR U61bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U61bar (
    .O(ybar[45]),
    .I0(abar[2]),
    .I1(bbar[13])
  );
  //AND U62
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U62 (
    .O(y[44]),
    .I0(a[2]),
    .I1(b[12])
  );
  //OR U62bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U62bar (
    .O(ybar[44]),
    .I0(abar[2]),
    .I1(bbar[12])
  );
  //AND U63
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U63 (
    .O(y[43]),
    .I0(a[2]),
    .I1(b[11])
  );
  //OR U63bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U63bar (
    .O(ybar[43]),
    .I0(abar[2]),
    .I1(bbar[11])
  );
  //AND U64
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U64 (
    .O(y[42]),
    .I0(a[2]),
    .I1(b[10])
  );
  //OR U64bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U64bar (
    .O(ybar[42]),
    .I0(abar[2]),
    .I1(bbar[10])
  );
  //AND U65
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U65 (
    .O(y[41]),
    .I0(a[2]),
    .I1(b[9])
  );
  //OR U65bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U65bar (
    .O(ybar[41]),
    .I0(abar[2]),
    .I1(bbar[9])
  );
  //AND U66
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U66 (
    .O(y[40]),
    .I0(a[2]),
    .I1(b[8])
  );
  //OR U66bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U66bar (
    .O(ybar[40]),
    .I0(abar[2]),
    .I1(bbar[8])
  );
  //AND U67
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U67 (
    .O(y[3]),
    .I0(b[3]),
    .I1(a[0])
  );
  //OR U67bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U67bar (
    .O(ybar[3]),
    .I0(bbar[3]),
    .I1(abar[0])
  );
  //AND U68
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U68 (
    .O(y[39]),
    .I0(a[2]),
    .I1(b[7])
  );
  //OR U68bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U68bar (
    .O(ybar[39]),
    .I0(abar[2]),
    .I1(bbar[7])
  );
  //AND U69
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U69 (
    .O(y[38]),
    .I0(a[2]),
    .I1(b[6])
  );
  //OR U69bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U69bar (
    .O(ybar[38]),
    .I0(abar[2]),
    .I1(bbar[6])
  );
  //AND U70
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U70 (
    .O(y[37]),
    .I0(a[2]),
    .I1(b[5])
  );
  //OR U70bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U70bar (
    .O(ybar[37]),
    .I0(abar[2]),
    .I1(bbar[5])
  );
  //AND U71
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U71 (
    .O(y[36]),
    .I0(a[2]),
    .I1(b[4])
  );
  //OR U71bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U71bar (
    .O(ybar[36]),
    .I0(abar[2]),
    .I1(bbar[4])
  );
  //AND U72
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U72 (
    .O(y[35]),
    .I0(a[2]),
    .I1(b[3])
  );
  //OR U72bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U72bar (
    .O(ybar[35]),
    .I0(abar[2]),
    .I1(bbar[3])
  );
  //AND U73
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U73 (
    .O(y[34]),
    .I0(a[2]),
    .I1(b[2])
  );
  //OR U73bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U73bar (
    .O(ybar[34]),
    .I0(abar[2]),
    .I1(bbar[2])
  );
  //AND U74
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U74 (
    .O(y[33]),
    .I0(a[2]),
    .I1(b[1])
  );
  //OR U74bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U74bar (
    .O(ybar[33]),
    .I0(abar[2]),
    .I1(bbar[1])
  );
  //AND U75
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U75 (
    .O(y[32]),
    .I0(a[2]),
    .I1(b[0])
  );
  //OR U75bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U75bar (
    .O(ybar[32]),
    .I0(abar[2]),
    .I1(bbar[0])
  );
  //AND U76
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U76 (
    .O(y[31]),
    .I0(a[1]),
    .I1(b[15])
  );
  //OR U76bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U76bar (
    .O(ybar[31]),
    .I0(abar[1]),
    .I1(bbar[15])
  );
  //AND U77
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U77 (
    .O(y[30]),
    .I0(a[1]),
    .I1(b[14])
  );
  //OR U77bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U77bar (
    .O(ybar[30]),
    .I0(abar[1]),
    .I1(bbar[14])
  );
  //AND U78
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U78 (
    .O(y[2]),
    .I0(b[2]),
    .I1(a[0])
  );
  //OR U78bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U78bar (
    .O(ybar[2]),
    .I0(bbar[2]),
    .I1(abar[0])
  );
  //AND U79
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U79 (
    .O(y[29]),
    .I0(a[1]),
    .I1(b[13])
  );
  //OR U79bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U79bar (
    .O(ybar[29]),
    .I0(abar[1]),
    .I1(bbar[13])
  );
  //AND U80
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U80 (
    .O(y[28]),
    .I0(a[1]),
    .I1(b[12])
  );
  //OR U80bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U80bar (
    .O(ybar[28]),
    .I0(abar[1]),
    .I1(bbar[12])
  );
  //AND U81
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U81 (
    .O(y[27]),
    .I0(a[1]),
    .I1(b[11])
  );
  //OR U81bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U81bar (
    .O(ybar[27]),
    .I0(abar[1]),
    .I1(bbar[11])
  );
  //AND U82
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U82 (
    .O(y[26]),
    .I0(a[1]),
    .I1(b[10])
  );
  //OR U82bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U82bar (
    .O(ybar[26]),
    .I0(abar[1]),
    .I1(bbar[10])
  );
  //AND U83
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U83 (
    .O(y[25]),
    .I0(a[1]),
    .I1(b[9])
  );
  //OR U83bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U83bar (
    .O(ybar[25]),
    .I0(abar[1]),
    .I1(bbar[9])
  );
  //AND U84
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U84 (
    .O(y[255]),
    .I0(a[15]),
    .I1(b[15])
  );
  //OR U84bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U84bar (
    .O(ybar[255]),
    .I0(abar[15]),
    .I1(bbar[15])
  );
  //AND U85
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U85 (
    .O(y[254]),
    .I0(a[15]),
    .I1(b[14])
  );
  //OR U85bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U85bar (
    .O(ybar[254]),
    .I0(abar[15]),
    .I1(bbar[14])
  );
  //AND U86
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U86 (
    .O(y[253]),
    .I0(a[15]),
    .I1(b[13])
  );
  //OR U86bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U86bar (
    .O(ybar[253]),
    .I0(abar[15]),
    .I1(bbar[13])
  );
  //AND U87
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U87 (
    .O(y[252]),
    .I0(a[15]),
    .I1(b[12])
  );
  //OR U87bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U87bar (
    .O(ybar[252]),
    .I0(abar[15]),
    .I1(bbar[12])
  );
  //AND U88
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U88 (
    .O(y[251]),
    .I0(a[15]),
    .I1(b[11])
  );
  //OR U88bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U88bar (
    .O(ybar[251]),
    .I0(abar[15]),
    .I1(bbar[11])
  );
  //AND U89
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U89 (
    .O(y[250]),
    .I0(a[15]),
    .I1(b[10])
  );
  //OR U89bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U89bar (
    .O(ybar[250]),
    .I0(abar[15]),
    .I1(bbar[10])
  );
  //AND U90
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U90 (
    .O(y[24]),
    .I0(a[1]),
    .I1(b[8])
  );
  //OR U90bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U90bar (
    .O(ybar[24]),
    .I0(abar[1]),
    .I1(bbar[8])
  );
  //AND U91
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U91 (
    .O(y[249]),
    .I0(a[15]),
    .I1(b[9])
  );
  //OR U91bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U91bar (
    .O(ybar[249]),
    .I0(abar[15]),
    .I1(bbar[9])
  );
  //AND U92
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U92 (
    .O(y[248]),
    .I0(a[15]),
    .I1(b[8])
  );
  //OR U92bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U92bar (
    .O(ybar[248]),
    .I0(abar[15]),
    .I1(bbar[8])
  );
  //AND U93
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U93 (
    .O(y[247]),
    .I0(a[15]),
    .I1(b[7])
  );
  //OR U93bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U93bar (
    .O(ybar[247]),
    .I0(abar[15]),
    .I1(bbar[7])
  );
  //AND U94
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U94 (
    .O(y[246]),
    .I0(a[15]),
    .I1(b[6])
  );
  //OR U94bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U94bar (
    .O(ybar[246]),
    .I0(abar[15]),
    .I1(bbar[6])
  );
  //AND U95
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U95 (
    .O(y[245]),
    .I0(a[15]),
    .I1(b[5])
  );
  //OR U95bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U95bar (
    .O(ybar[245]),
    .I0(abar[15]),
    .I1(bbar[5])
  );
  //AND U96
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U96 (
    .O(y[244]),
    .I0(a[15]),
    .I1(b[4])
  );
  //OR U96bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U96bar (
    .O(ybar[244]),
    .I0(abar[15]),
    .I1(bbar[4])
  );
  //AND U97
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U97 (
    .O(y[243]),
    .I0(a[15]),
    .I1(b[3])
  );
  //OR U97bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U97bar (
    .O(ybar[243]),
    .I0(abar[15]),
    .I1(bbar[3])
  );
  //AND U98
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U98 (
    .O(y[242]),
    .I0(a[15]),
    .I1(b[2])
  );
  //OR U98bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U98bar (
    .O(ybar[242]),
    .I0(abar[15]),
    .I1(bbar[2])
  );
  //AND U99
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U99 (
    .O(y[241]),
    .I0(a[15]),
    .I1(b[1])
  );
  //OR U99bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U99bar (
    .O(ybar[241]),
    .I0(abar[15]),
    .I1(bbar[1])
  );
  //AND U100
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U100 (
    .O(y[240]),
    .I0(a[15]),
    .I1(b[0])
  );
  //OR U100bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U100bar (
    .O(ybar[240]),
    .I0(abar[15]),
    .I1(bbar[0])
  );
  //AND U101
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U101 (
    .O(y[23]),
    .I0(a[1]),
    .I1(b[7])
  );
  //OR U101bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U101bar (
    .O(ybar[23]),
    .I0(abar[1]),
    .I1(bbar[7])
  );
  //AND U102
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U102 (
    .O(y[239]),
    .I0(a[14]),
    .I1(b[15])
  );
  //OR U102bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U102bar (
    .O(ybar[239]),
    .I0(abar[14]),
    .I1(bbar[15])
  );
  //AND U103
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U103 (
    .O(y[238]),
    .I0(a[14]),
    .I1(b[14])
  );
  //OR U103bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U103bar (
    .O(ybar[238]),
    .I0(abar[14]),
    .I1(bbar[14])
  );
  //AND U104
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U104 (
    .O(y[237]),
    .I0(a[14]),
    .I1(b[13])
  );
  //OR U104bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U104bar (
    .O(ybar[237]),
    .I0(abar[14]),
    .I1(bbar[13])
  );
  //AND U105
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U105 (
    .O(y[236]),
    .I0(a[14]),
    .I1(b[12])
  );
  //OR U105bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U105bar (
    .O(ybar[236]),
    .I0(abar[14]),
    .I1(bbar[12])
  );
  //AND U106
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U106 (
    .O(y[235]),
    .I0(a[14]),
    .I1(b[11])
  );
  //OR U106bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U106bar (
    .O(ybar[235]),
    .I0(abar[14]),
    .I1(bbar[11])
  );
  //AND U107
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U107 (
    .O(y[234]),
    .I0(a[14]),
    .I1(b[10])
  );
  //OR U107bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U107bar (
    .O(ybar[234]),
    .I0(abar[14]),
    .I1(bbar[10])
  );
  //AND U108
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U108 (
    .O(y[233]),
    .I0(a[14]),
    .I1(b[9])
  );
  //OR U108bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U108bar (
    .O(ybar[233]),
    .I0(abar[14]),
    .I1(bbar[9])
  );
  //AND U109
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U109 (
    .O(y[232]),
    .I0(a[14]),
    .I1(b[8])
  );
  //OR U109bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U109bar (
    .O(ybar[232]),
    .I0(abar[14]),
    .I1(bbar[8])
  );
  //AND U110
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U110 (
    .O(y[231]),
    .I0(a[14]),
    .I1(b[7])
  );
  //OR U110bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U110bar (
    .O(ybar[231]),
    .I0(abar[14]),
    .I1(bbar[7])
  );
  //AND U111
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U111 (
    .O(y[230]),
    .I0(a[14]),
    .I1(b[6])
  );
  //OR U111bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U111bar (
    .O(ybar[230]),
    .I0(abar[14]),
    .I1(bbar[6])
  );
  //AND U112
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U112 (
    .O(y[22]),
    .I0(a[1]),
    .I1(b[6])
  );
  //OR U112bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U112bar (
    .O(ybar[22]),
    .I0(abar[1]),
    .I1(bbar[6])
  );
  //AND U113
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U113 (
    .O(y[229]),
    .I0(a[14]),
    .I1(b[5])
  );
  //OR U113bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U113bar (
    .O(ybar[229]),
    .I0(abar[14]),
    .I1(bbar[5])
  );
  //AND U114
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U114 (
    .O(y[228]),
    .I0(a[14]),
    .I1(b[4])
  );
  //OR U114bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U114bar (
    .O(ybar[228]),
    .I0(abar[14]),
    .I1(bbar[4])
  );
  //AND U115
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U115 (
    .O(y[227]),
    .I0(a[14]),
    .I1(b[3])
  );
  //OR U115bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U115bar (
    .O(ybar[227]),
    .I0(abar[14]),
    .I1(bbar[3])
  );
  //AND U116
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U116 (
    .O(y[226]),
    .I0(a[14]),
    .I1(b[2])
  );
  //OR U116bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U116bar (
    .O(ybar[226]),
    .I0(abar[14]),
    .I1(bbar[2])
  );
  //AND U117
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U117 (
    .O(y[225]),
    .I0(a[14]),
    .I1(b[1])
  );
  //OR U117bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U117bar (
    .O(ybar[225]),
    .I0(abar[14]),
    .I1(bbar[1])
  );
  //AND U118
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U118 (
    .O(y[224]),
    .I0(a[14]),
    .I1(b[0])
  );
  //OR U118bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U118bar (
    .O(ybar[224]),
    .I0(abar[14]),
    .I1(bbar[0])
  );
  //AND U119
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U119 (
    .O(y[223]),
    .I0(a[13]),
    .I1(b[15])
  );
  //OR U119bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U119bar (
    .O(ybar[223]),
    .I0(abar[13]),
    .I1(bbar[15])
  );
  //AND U120
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U120 (
    .O(y[222]),
    .I0(a[13]),
    .I1(b[14])
  );
  //OR U120bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U120bar (
    .O(ybar[222]),
    .I0(abar[13]),
    .I1(bbar[14])
  );
  //AND U121
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U121 (
    .O(y[221]),
    .I0(a[13]),
    .I1(b[13])
  );
  //OR U121bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U121bar (
    .O(ybar[221]),
    .I0(abar[13]),
    .I1(bbar[13])
  );
  //AND U122
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U122 (
    .O(y[220]),
    .I0(a[13]),
    .I1(b[12])
  );
  //OR U122bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U122bar (
    .O(ybar[220]),
    .I0(abar[13]),
    .I1(bbar[12])
  );
  //AND U123
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U123 (
    .O(y[21]),
    .I0(a[1]),
    .I1(b[5])
  );
  //OR U123bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U123bar (
    .O(ybar[21]),
    .I0(abar[1]),
    .I1(bbar[5])
  );
  //AND U124
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U124 (
    .O(y[219]),
    .I0(a[13]),
    .I1(b[11])
  );
  //OR U124bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U124bar (
    .O(ybar[219]),
    .I0(abar[13]),
    .I1(bbar[11])
  );
  //AND U125
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U125 (
    .O(y[218]),
    .I0(a[13]),
    .I1(b[10])
  );
  //OR U125bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U125bar (
    .O(ybar[218]),
    .I0(abar[13]),
    .I1(bbar[10])
  );
  //AND U126
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U126 (
    .O(y[217]),
    .I0(a[13]),
    .I1(b[9])
  );
  //OR U126bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U126bar (
    .O(ybar[217]),
    .I0(abar[13]),
    .I1(bbar[9])
  );
  //AND U127
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U127 (
    .O(y[216]),
    .I0(a[13]),
    .I1(b[8])
  );
  //OR U127bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U127bar (
    .O(ybar[216]),
    .I0(abar[13]),
    .I1(bbar[8])
  );
  //AND U128
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U128 (
    .O(y[215]),
    .I0(a[13]),
    .I1(b[7])
  );
  //OR U128bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U128bar (
    .O(ybar[215]),
    .I0(abar[13]),
    .I1(bbar[7])
  );
  //AND U129
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U129 (
    .O(y[214]),
    .I0(a[13]),
    .I1(b[6])
  );
  //OR U129bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U129bar (
    .O(ybar[214]),
    .I0(abar[13]),
    .I1(bbar[6])
  );
  //AND U130
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U130 (
    .O(y[213]),
    .I0(a[13]),
    .I1(b[5])
  );
  //OR U130bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U130bar (
    .O(ybar[213]),
    .I0(abar[13]),
    .I1(bbar[5])
  );
  //AND U131
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U131 (
    .O(y[212]),
    .I0(a[13]),
    .I1(b[4])
  );
  //OR U131bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U131bar (
    .O(ybar[212]),
    .I0(abar[13]),
    .I1(bbar[4])
  );
  //AND U132
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U132 (
    .O(y[211]),
    .I0(a[13]),
    .I1(b[3])
  );
  //OR U132bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U132bar (
    .O(ybar[211]),
    .I0(abar[13]),
    .I1(bbar[3])
  );
  //AND U133
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U133 (
    .O(y[210]),
    .I0(a[13]),
    .I1(b[2])
  );
  //OR U133bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U133bar (
    .O(ybar[210]),
    .I0(abar[13]),
    .I1(bbar[2])
  );
  //AND U134
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U134 (
    .O(y[20]),
    .I0(a[1]),
    .I1(b[4])
  );
  //OR U134bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U134bar (
    .O(ybar[20]),
    .I0(abar[1]),
    .I1(bbar[4])
  );
  //AND U135
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U135 (
    .O(y[209]),
    .I0(a[13]),
    .I1(b[1])
  );
  //OR U135bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U135bar (
    .O(ybar[209]),
    .I0(abar[13]),
    .I1(bbar[1])
  );
  //AND U136
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U136 (
    .O(y[208]),
    .I0(a[13]),
    .I1(b[0])
  );
  //OR U136bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U136bar (
    .O(ybar[208]),
    .I0(abar[13]),
    .I1(bbar[0])
  );
  //AND U137
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U137 (
    .O(y[207]),
    .I0(a[12]),
    .I1(b[15])
  );
  //OR U137bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U137bar (
    .O(ybar[207]),
    .I0(abar[12]),
    .I1(bbar[15])
  );
  //AND U138
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U138 (
    .O(y[206]),
    .I0(a[12]),
    .I1(b[14])
  );
  //OR U138bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U138bar (
    .O(ybar[206]),
    .I0(abar[12]),
    .I1(bbar[14])
  );
  //AND U139
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U139 (
    .O(y[205]),
    .I0(a[12]),
    .I1(b[13])
  );
  //OR U139bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U139bar (
    .O(ybar[205]),
    .I0(abar[12]),
    .I1(bbar[13])
  );
  //AND U140
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U140 (
    .O(y[204]),
    .I0(a[12]),
    .I1(b[12])
  );
  //OR U140bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U140bar (
    .O(ybar[204]),
    .I0(abar[12]),
    .I1(bbar[12])
  );
  //AND U141
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U141 (
    .O(y[203]),
    .I0(a[12]),
    .I1(b[11])
  );
  //OR U141bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U141bar (
    .O(ybar[203]),
    .I0(abar[12]),
    .I1(bbar[11])
  );
  //AND U142
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U142 (
    .O(y[202]),
    .I0(a[12]),
    .I1(b[10])
  );
  //OR U142bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U142bar (
    .O(ybar[202]),
    .I0(abar[12]),
    .I1(bbar[10])
  );
  //AND U143
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U143 (
    .O(y[201]),
    .I0(a[12]),
    .I1(b[9])
  );
  //OR U143bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U143bar (
    .O(ybar[201]),
    .I0(abar[12]),
    .I1(bbar[9])
  );
  //AND U144
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U144 (
    .O(y[200]),
    .I0(a[12]),
    .I1(b[8])
  );
  //OR U144bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U144bar (
    .O(ybar[200]),
    .I0(abar[12]),
    .I1(bbar[8])
  );
  //AND U145
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U145 (
    .O(y[1]),
    .I0(b[1]),
    .I1(a[0])
  );
  //OR U145bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U145bar (
    .O(ybar[1]),
    .I0(bbar[1]),
    .I1(abar[0])
  );
  //AND U146
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U146 (
    .O(y[19]),
    .I0(a[1]),
    .I1(b[3])
  );
  //OR U146bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U146bar (
    .O(ybar[19]),
    .I0(abar[1]),
    .I1(bbar[3])
  );
  //AND U147
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U147 (
    .O(y[199]),
    .I0(a[12]),
    .I1(b[7])
  );
  //OR U147bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U147bar (
    .O(ybar[199]),
    .I0(abar[12]),
    .I1(bbar[7])
  );
  //AND U148
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U148 (
    .O(y[198]),
    .I0(a[12]),
    .I1(b[6])
  );
  //OR U148bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U148bar (
    .O(ybar[198]),
    .I0(abar[12]),
    .I1(bbar[6])
  );
  //AND U149
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U149 (
    .O(y[197]),
    .I0(a[12]),
    .I1(b[5])
  );
  //OR U149bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U149bar (
    .O(ybar[197]),
    .I0(abar[12]),
    .I1(bbar[5])
  );
  //AND U150
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U150 (
    .O(y[196]),
    .I0(a[12]),
    .I1(b[4])
  );
  //OR U150bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U150bar (
    .O(ybar[196]),
    .I0(abar[12]),
    .I1(bbar[4])
  );
  //AND U151
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U151 (
    .O(y[195]),
    .I0(a[12]),
    .I1(b[3])
  );
  //OR U151bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U151bar (
    .O(ybar[195]),
    .I0(abar[12]),
    .I1(bbar[3])
  );
  //AND U152
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U152 (
    .O(y[194]),
    .I0(a[12]),
    .I1(b[2])
  );
  //OR U152bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U152bar (
    .O(ybar[194]),
    .I0(abar[12]),
    .I1(bbar[2])
  );
  //AND U153
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U153 (
    .O(y[193]),
    .I0(a[12]),
    .I1(b[1])
  );
  //OR U153bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U153bar (
    .O(ybar[193]),
    .I0(abar[12]),
    .I1(bbar[1])
  );
  //AND U154
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U154 (
    .O(y[192]),
    .I0(a[12]),
    .I1(b[0])
  );
  //OR U154bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U154bar (
    .O(ybar[192]),
    .I0(abar[12]),
    .I1(bbar[0])
  );
  //AND U155
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U155 (
    .O(y[191]),
    .I0(a[11]),
    .I1(b[15])
  );
  //OR U155bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U155bar (
    .O(ybar[191]),
    .I0(abar[11]),
    .I1(bbar[15])
  );
  //AND U156
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U156 (
    .O(y[190]),
    .I0(a[11]),
    .I1(b[14])
  );
  //OR U156bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U156bar (
    .O(ybar[190]),
    .I0(abar[11]),
    .I1(bbar[14])
  );
  //AND U157
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U157 (
    .O(y[18]),
    .I0(a[1]),
    .I1(b[2])
  );
  //OR U157bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U157bar (
    .O(ybar[18]),
    .I0(abar[1]),
    .I1(bbar[2])
  );
  //AND U158
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U158 (
    .O(y[189]),
    .I0(a[11]),
    .I1(b[13])
  );
  //OR U158bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U158bar (
    .O(ybar[189]),
    .I0(abar[11]),
    .I1(bbar[13])
  );
  //AND U159
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U159 (
    .O(y[188]),
    .I0(a[11]),
    .I1(b[12])
  );
  //OR U159bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U159bar (
    .O(ybar[188]),
    .I0(abar[11]),
    .I1(bbar[12])
  );
  //AND U160
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U160 (
    .O(y[187]),
    .I0(a[11]),
    .I1(b[11])
  );
  //OR U160bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U160bar (
    .O(ybar[187]),
    .I0(abar[11]),
    .I1(bbar[11])
  );
  //AND U161
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U161 (
    .O(y[186]),
    .I0(a[11]),
    .I1(b[10])
  );
  //OR U161bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U161bar (
    .O(ybar[186]),
    .I0(abar[11]),
    .I1(bbar[10])
  );
  //AND U162
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U162 (
    .O(y[185]),
    .I0(a[11]),
    .I1(b[9])
  );
  //OR U162bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U162bar (
    .O(ybar[185]),
    .I0(abar[11]),
    .I1(bbar[9])
  );
  //AND U163
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U163 (
    .O(y[184]),
    .I0(a[11]),
    .I1(b[8])
  );
  //OR U163bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U163bar (
    .O(ybar[184]),
    .I0(abar[11]),
    .I1(bbar[8])
  );
  //AND U164
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U164 (
    .O(y[183]),
    .I0(a[11]),
    .I1(b[7])
  );
  //OR U164bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U164bar (
    .O(ybar[183]),
    .I0(abar[11]),
    .I1(bbar[7])
  );
  //AND U165
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U165 (
    .O(y[182]),
    .I0(a[11]),
    .I1(b[6])
  );
  //OR U165bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U165bar (
    .O(ybar[182]),
    .I0(abar[11]),
    .I1(bbar[6])
  );
  //AND U166
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U166 (
    .O(y[181]),
    .I0(a[11]),
    .I1(b[5])
  );
  //OR U166bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U166bar (
    .O(ybar[181]),
    .I0(abar[11]),
    .I1(bbar[5])
  );
  //AND U167
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U167 (
    .O(y[180]),
    .I0(a[11]),
    .I1(b[4])
  );
  //OR U167bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U167bar (
    .O(ybar[180]),
    .I0(abar[11]),
    .I1(bbar[4])
  );
  //AND U168
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U168 (
    .O(y[17]),
    .I0(a[1]),
    .I1(b[1])
  );
  //OR U168bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U168bar (
    .O(ybar[17]),
    .I0(abar[1]),
    .I1(bbar[1])
  );
  //AND U169
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U169 (
    .O(y[179]),
    .I0(a[11]),
    .I1(b[3])
  );
  //OR U169bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U169bar (
    .O(ybar[179]),
    .I0(abar[11]),
    .I1(bbar[3])
  );
  //AND U170
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U170 (
    .O(y[178]),
    .I0(a[11]),
    .I1(b[2])
  );
  //OR U170bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U170bar (
    .O(ybar[178]),
    .I0(abar[11]),
    .I1(bbar[2])
  );
  //AND U171
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U171 (
    .O(y[177]),
    .I0(a[11]),
    .I1(b[1])
  );
  //OR U171bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U171bar (
    .O(ybar[177]),
    .I0(abar[11]),
    .I1(bbar[1])
  );
  //AND U172
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U172 (
    .O(y[176]),
    .I0(a[11]),
    .I1(b[0])
  );
  //OR U172bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U172bar (
    .O(ybar[176]),
    .I0(abar[11]),
    .I1(bbar[0])
  );
  //AND U173
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U173 (
    .O(y[175]),
    .I0(a[10]),
    .I1(b[15])
  );
  //OR U173bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U173bar (
    .O(ybar[175]),
    .I0(abar[10]),
    .I1(bbar[15])
  );
  //AND U174
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U174 (
    .O(y[174]),
    .I0(a[10]),
    .I1(b[14])
  );
  //OR U174bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U174bar (
    .O(ybar[174]),
    .I0(abar[10]),
    .I1(bbar[14])
  );
  //AND U175
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U175 (
    .O(y[173]),
    .I0(a[10]),
    .I1(b[13])
  );
  //OR U175bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U175bar (
    .O(ybar[173]),
    .I0(abar[10]),
    .I1(bbar[13])
  );
  //AND U176
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U176 (
    .O(y[172]),
    .I0(a[10]),
    .I1(b[12])
  );
  //OR U176bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U176bar (
    .O(ybar[172]),
    .I0(abar[10]),
    .I1(bbar[12])
  );
  //AND U177
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U177 (
    .O(y[171]),
    .I0(a[10]),
    .I1(b[11])
  );
  //OR U177bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U177bar (
    .O(ybar[171]),
    .I0(abar[10]),
    .I1(bbar[11])
  );
  //AND U178
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U178 (
    .O(y[170]),
    .I0(a[10]),
    .I1(b[10])
  );
  //OR U178bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U178bar (
    .O(ybar[170]),
    .I0(abar[10]),
    .I1(bbar[10])
  );
  //AND U179
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U179 (
    .O(y[16]),
    .I0(a[1]),
    .I1(b[0])
  );
  //OR U179bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U179bar (
    .O(ybar[16]),
    .I0(abar[1]),
    .I1(bbar[0])
  );
  //AND U180
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U180 (
    .O(y[169]),
    .I0(a[10]),
    .I1(b[9])
  );
  //OR U180bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U180bar (
    .O(ybar[169]),
    .I0(abar[10]),
    .I1(bbar[9])
  );
  //AND U181
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U181 (
    .O(y[168]),
    .I0(a[10]),
    .I1(b[8])
  );
  //OR U181bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U181bar (
    .O(ybar[168]),
    .I0(abar[10]),
    .I1(bbar[8])
  );
  //AND U182
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U182 (
    .O(y[167]),
    .I0(a[10]),
    .I1(b[7])
  );
  //OR U182bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U182bar (
    .O(ybar[167]),
    .I0(abar[10]),
    .I1(bbar[7])
  );
  //AND U183
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U183 (
    .O(y[166]),
    .I0(a[10]),
    .I1(b[6])
  );
  //OR U183bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U183bar (
    .O(ybar[166]),
    .I0(abar[10]),
    .I1(bbar[6])
  );
  //AND U184
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U184 (
    .O(y[165]),
    .I0(a[10]),
    .I1(b[5])
  );
  //OR U184bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U184bar (
    .O(ybar[165]),
    .I0(abar[10]),
    .I1(bbar[5])
  );
  //AND U185
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U185 (
    .O(y[164]),
    .I0(a[10]),
    .I1(b[4])
  );
  //OR U185bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U185bar (
    .O(ybar[164]),
    .I0(abar[10]),
    .I1(bbar[4])
  );
  //AND U186
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U186 (
    .O(y[163]),
    .I0(a[10]),
    .I1(b[3])
  );
  //OR U186bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U186bar (
    .O(ybar[163]),
    .I0(abar[10]),
    .I1(bbar[3])
  );
  //AND U187
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U187 (
    .O(y[162]),
    .I0(a[10]),
    .I1(b[2])
  );
  //OR U187bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U187bar (
    .O(ybar[162]),
    .I0(abar[10]),
    .I1(bbar[2])
  );
  //AND U188
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U188 (
    .O(y[161]),
    .I0(a[10]),
    .I1(b[1])
  );
  //OR U188bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U188bar (
    .O(ybar[161]),
    .I0(abar[10]),
    .I1(bbar[1])
  );
  //AND U189
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U189 (
    .O(y[160]),
    .I0(a[10]),
    .I1(b[0])
  );
  //OR U189bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U189bar (
    .O(ybar[160]),
    .I0(abar[10]),
    .I1(bbar[0])
  );
  //AND U190
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U190 (
    .O(y[15]),
    .I0(b[15]),
    .I1(a[0])
  );
  //OR U190bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U190bar (
    .O(ybar[15]),
    .I0(bbar[15]),
    .I1(abar[0])
  );
  //AND U191
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U191 (
    .O(y[159]),
    .I0(a[9]),
    .I1(b[15])
  );
  //OR U191bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U191bar (
    .O(ybar[159]),
    .I0(abar[9]),
    .I1(bbar[15])
  );
  //AND U192
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U192 (
    .O(y[158]),
    .I0(a[9]),
    .I1(b[14])
  );
  //OR U192bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U192bar (
    .O(ybar[158]),
    .I0(abar[9]),
    .I1(bbar[14])
  );
  //AND U193
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U193 (
    .O(y[157]),
    .I0(a[9]),
    .I1(b[13])
  );
  //OR U193bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U193bar (
    .O(ybar[157]),
    .I0(abar[9]),
    .I1(bbar[13])
  );
  //AND U194
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U194 (
    .O(y[156]),
    .I0(a[9]),
    .I1(b[12])
  );
  //OR U194bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U194bar (
    .O(ybar[156]),
    .I0(abar[9]),
    .I1(bbar[12])
  );
  //AND U195
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U195 (
    .O(y[155]),
    .I0(a[9]),
    .I1(b[11])
  );
  //OR U195bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U195bar (
    .O(ybar[155]),
    .I0(abar[9]),
    .I1(bbar[11])
  );
  //AND U196
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U196 (
    .O(y[154]),
    .I0(a[9]),
    .I1(b[10])
  );
  //OR U196bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U196bar (
    .O(ybar[154]),
    .I0(abar[9]),
    .I1(bbar[10])
  );
  //AND U197
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U197 (
    .O(y[153]),
    .I0(a[9]),
    .I1(b[9])
  );
  //OR U197bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U197bar (
    .O(ybar[153]),
    .I0(abar[9]),
    .I1(bbar[9])
  );
  //AND U198
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U198 (
    .O(y[152]),
    .I0(a[9]),
    .I1(b[8])
  );
  //OR U198bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U198bar (
    .O(ybar[152]),
    .I0(abar[9]),
    .I1(bbar[8])
  );
  //AND U199
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U199 (
    .O(y[151]),
    .I0(a[9]),
    .I1(b[7])
  );
  //OR U199bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U199bar (
    .O(ybar[151]),
    .I0(abar[9]),
    .I1(bbar[7])
  );
  //AND U200
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U200 (
    .O(y[150]),
    .I0(a[9]),
    .I1(b[6])
  );
  //OR U200bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U200bar (
    .O(ybar[150]),
    .I0(abar[9]),
    .I1(bbar[6])
  );
  //AND U201
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U201 (
    .O(y[14]),
    .I0(b[14]),
    .I1(a[0])
  );
  //OR U201bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U201bar (
    .O(ybar[14]),
    .I0(bbar[14]),
    .I1(abar[0])
  );
  //AND U202
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U202 (
    .O(y[149]),
    .I0(a[9]),
    .I1(b[5])
  );
  //OR U202bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U202bar (
    .O(ybar[149]),
    .I0(abar[9]),
    .I1(bbar[5])
  );
  //AND U203
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U203 (
    .O(y[148]),
    .I0(a[9]),
    .I1(b[4])
  );
  //OR U203bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U203bar (
    .O(ybar[148]),
    .I0(abar[9]),
    .I1(bbar[4])
  );
  //AND U204
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U204 (
    .O(y[147]),
    .I0(a[9]),
    .I1(b[3])
  );
  //OR U204bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U204bar (
    .O(ybar[147]),
    .I0(abar[9]),
    .I1(bbar[3])
  );
  //AND U205
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U205 (
    .O(y[146]),
    .I0(a[9]),
    .I1(b[2])
  );
  //OR U205bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U205bar (
    .O(ybar[146]),
    .I0(abar[9]),
    .I1(bbar[2])
  );
  //AND U206
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U206 (
    .O(y[145]),
    .I0(a[9]),
    .I1(b[1])
  );
  //OR U206bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U206bar (
    .O(ybar[145]),
    .I0(abar[9]),
    .I1(bbar[1])
  );
  //AND U207
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U207 (
    .O(y[144]),
    .I0(a[9]),
    .I1(b[0])
  );
  //OR U207bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U207bar (
    .O(ybar[144]),
    .I0(abar[9]),
    .I1(bbar[0])
  );
  //AND U208
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U208 (
    .O(y[143]),
    .I0(a[8]),
    .I1(b[15])
  );
  //OR U208bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U208bar (
    .O(ybar[143]),
    .I0(abar[8]),
    .I1(bbar[15])
  );
  //AND U209
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U209 (
    .O(y[142]),
    .I0(a[8]),
    .I1(b[14])
  );
  //OR U209bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U209bar (
    .O(ybar[142]),
    .I0(abar[8]),
    .I1(bbar[14])
  );
  //AND U210
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U210 (
    .O(y[141]),
    .I0(a[8]),
    .I1(b[13])
  );
  //OR U210bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U210bar (
    .O(ybar[141]),
    .I0(abar[8]),
    .I1(bbar[13])
  );
  //AND U211
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U211 (
    .O(y[140]),
    .I0(a[8]),
    .I1(b[12])
  );
  //OR U211bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U211bar (
    .O(ybar[140]),
    .I0(abar[8]),
    .I1(bbar[12])
  );
  //AND U212
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U212 (
    .O(y[13]),
    .I0(b[13]),
    .I1(a[0])
  );
  //OR U212bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U212bar (
    .O(ybar[13]),
    .I0(bbar[13]),
    .I1(abar[0])
  );
  //AND U213
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U213 (
    .O(y[139]),
    .I0(a[8]),
    .I1(b[11])
  );
  //OR U213bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U213bar (
    .O(ybar[139]),
    .I0(abar[8]),
    .I1(bbar[11])
  );
  //AND U214
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U214 (
    .O(y[138]),
    .I0(a[8]),
    .I1(b[10])
  );
  //OR U214bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U214bar (
    .O(ybar[138]),
    .I0(abar[8]),
    .I1(bbar[10])
  );
  //AND U215
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U215 (
    .O(y[137]),
    .I0(a[8]),
    .I1(b[9])
  );
  //OR U215bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U215bar (
    .O(ybar[137]),
    .I0(abar[8]),
    .I1(bbar[9])
  );
  //AND U216
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U216 (
    .O(y[136]),
    .I0(a[8]),
    .I1(b[8])
  );
  //OR U216bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U216bar (
    .O(ybar[136]),
    .I0(abar[8]),
    .I1(bbar[8])
  );
  //AND U217
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U217 (
    .O(y[135]),
    .I0(a[8]),
    .I1(b[7])
  );
  //OR U217bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U217bar (
    .O(ybar[135]),
    .I0(abar[8]),
    .I1(bbar[7])
  );
  //AND U218
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U218 (
    .O(y[134]),
    .I0(a[8]),
    .I1(b[6])
  );
  //OR U218bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U218bar (
    .O(ybar[134]),
    .I0(abar[8]),
    .I1(bbar[6])
  );
  //AND U219
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U219 (
    .O(y[133]),
    .I0(a[8]),
    .I1(b[5])
  );
  //OR U219bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U219bar (
    .O(ybar[133]),
    .I0(abar[8]),
    .I1(bbar[5])
  );
  //AND U220
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U220 (
    .O(y[132]),
    .I0(a[8]),
    .I1(b[4])
  );
  //OR U220bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U220bar (
    .O(ybar[132]),
    .I0(abar[8]),
    .I1(bbar[4])
  );
  //AND U221
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U221 (
    .O(y[131]),
    .I0(a[8]),
    .I1(b[3])
  );
  //OR U221bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U221bar (
    .O(ybar[131]),
    .I0(abar[8]),
    .I1(bbar[3])
  );
  //AND U222
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U222 (
    .O(y[130]),
    .I0(a[8]),
    .I1(b[2])
  );
  //OR U222bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U222bar (
    .O(ybar[130]),
    .I0(abar[8]),
    .I1(bbar[2])
  );
  //AND U223
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U223 (
    .O(y[12]),
    .I0(b[12]),
    .I1(a[0])
  );
  //OR U223bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U223bar (
    .O(ybar[12]),
    .I0(bbar[12]),
    .I1(abar[0])
  );
  //AND U224
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U224 (
    .O(y[129]),
    .I0(a[8]),
    .I1(b[1])
  );
  //OR U224bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U224bar (
    .O(ybar[129]),
    .I0(abar[8]),
    .I1(bbar[1])
  );
  //AND U225
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U225 (
    .O(y[128]),
    .I0(a[8]),
    .I1(b[0])
  );
  //OR U225bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U225bar (
    .O(ybar[128]),
    .I0(abar[8]),
    .I1(bbar[0])
  );
  //AND U226
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U226 (
    .O(y[127]),
    .I0(a[7]),
    .I1(b[15])
  );
  //OR U226bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U226bar (
    .O(ybar[127]),
    .I0(abar[7]),
    .I1(bbar[15])
  );
  //AND U227
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U227 (
    .O(y[126]),
    .I0(a[7]),
    .I1(b[14])
  );
  //OR U227bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U227bar (
    .O(ybar[126]),
    .I0(abar[7]),
    .I1(bbar[14])
  );
  //AND U228
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U228 (
    .O(y[125]),
    .I0(a[7]),
    .I1(b[13])
  );
  //OR U228bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U228bar (
    .O(ybar[125]),
    .I0(abar[7]),
    .I1(bbar[13])
  );
  //AND U229
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U229 (
    .O(y[124]),
    .I0(a[7]),
    .I1(b[12])
  );
  //OR U229bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U229bar (
    .O(ybar[124]),
    .I0(abar[7]),
    .I1(bbar[12])
  );
  //AND U230
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U230 (
    .O(y[123]),
    .I0(a[7]),
    .I1(b[11])
  );
  //OR U230bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U230bar (
    .O(ybar[123]),
    .I0(abar[7]),
    .I1(bbar[11])
  );
  //AND U231
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U231 (
    .O(y[122]),
    .I0(a[7]),
    .I1(b[10])
  );
  //OR U231bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U231bar (
    .O(ybar[122]),
    .I0(abar[7]),
    .I1(bbar[10])
  );
  //AND U232
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U232 (
    .O(y[121]),
    .I0(a[7]),
    .I1(b[9])
  );
  //OR U232bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U232bar (
    .O(ybar[121]),
    .I0(abar[7]),
    .I1(bbar[9])
  );
  //AND U233
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U233 (
    .O(y[120]),
    .I0(a[7]),
    .I1(b[8])
  );
  //OR U233bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U233bar (
    .O(ybar[120]),
    .I0(abar[7]),
    .I1(bbar[8])
  );
  //AND U234
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U234 (
    .O(y[11]),
    .I0(b[11]),
    .I1(a[0])
  );
  //OR U234bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U234bar (
    .O(ybar[11]),
    .I0(bbar[11]),
    .I1(abar[0])
  );
  //AND U235
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U235 (
    .O(y[119]),
    .I0(a[7]),
    .I1(b[7])
  );
  //OR U235bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U235bar (
    .O(ybar[119]),
    .I0(abar[7]),
    .I1(bbar[7])
  );
  //AND U236
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U236 (
    .O(y[118]),
    .I0(a[7]),
    .I1(b[6])
  );
  //OR U236bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U236bar (
    .O(ybar[118]),
    .I0(abar[7]),
    .I1(bbar[6])
  );
  //AND U237
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U237 (
    .O(y[117]),
    .I0(a[7]),
    .I1(b[5])
  );
  //OR U237bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U237bar (
    .O(ybar[117]),
    .I0(abar[7]),
    .I1(bbar[5])
  );
  //AND U238
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U238 (
    .O(y[116]),
    .I0(a[7]),
    .I1(b[4])
  );
  //OR U238bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U238bar (
    .O(ybar[116]),
    .I0(abar[7]),
    .I1(bbar[4])
  );
  //AND U239
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U239 (
    .O(y[115]),
    .I0(a[7]),
    .I1(b[3])
  );
  //OR U239bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U239bar (
    .O(ybar[115]),
    .I0(abar[7]),
    .I1(bbar[3])
  );
  //AND U240
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U240 (
    .O(y[114]),
    .I0(a[7]),
    .I1(b[2])
  );
  //OR U240bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U240bar (
    .O(ybar[114]),
    .I0(abar[7]),
    .I1(bbar[2])
  );
  //AND U241
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U241 (
    .O(y[113]),
    .I0(a[7]),
    .I1(b[1])
  );
  //OR U241bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U241bar (
    .O(ybar[113]),
    .I0(abar[7]),
    .I1(bbar[1])
  );
  //AND U242
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U242 (
    .O(y[112]),
    .I0(a[7]),
    .I1(b[0])
  );
  //OR U242bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U242bar (
    .O(ybar[112]),
    .I0(abar[7]),
    .I1(bbar[0])
  );
  //AND U243
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U243 (
    .O(y[111]),
    .I0(b[15]),
    .I1(a[6])
  );
  //OR U243bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U243bar (
    .O(ybar[111]),
    .I0(bbar[15]),
    .I1(abar[6])
  );
  //AND U244
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U244 (
    .O(y[110]),
    .I0(b[14]),
    .I1(a[6])
  );
  //OR U244bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U244bar (
    .O(ybar[110]),
    .I0(bbar[14]),
    .I1(abar[6])
  );
  //AND U245
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U245 (
    .O(y[10]),
    .I0(b[10]),
    .I1(a[0])
  );
  //OR U245bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U245bar (
    .O(ybar[10]),
    .I0(bbar[10]),
    .I1(abar[0])
  );
  //AND U246
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U246 (
    .O(y[109]),
    .I0(b[13]),
    .I1(a[6])
  );
  //OR U246bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U246bar (
    .O(ybar[109]),
    .I0(bbar[13]),
    .I1(abar[6])
  );
  //AND U247
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U247 (
    .O(y[108]),
    .I0(b[12]),
    .I1(a[6])
  );
  //OR U247bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U247bar (
    .O(ybar[108]),
    .I0(bbar[12]),
    .I1(abar[6])
  );
  //AND U248
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U248 (
    .O(y[107]),
    .I0(b[11]),
    .I1(a[6])
  );
  //OR U248bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U248bar (
    .O(ybar[107]),
    .I0(bbar[11]),
    .I1(abar[6])
  );
  //AND U249
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U249 (
    .O(y[106]),
    .I0(b[10]),
    .I1(a[6])
  );
  //OR U249bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U249bar (
    .O(ybar[106]),
    .I0(bbar[10]),
    .I1(abar[6])
  );
  //AND U250
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U250 (
    .O(y[105]),
    .I0(a[6]),
    .I1(b[9])
  );
  //OR U250bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U250bar (
    .O(ybar[105]),
    .I0(abar[6]),
    .I1(bbar[9])
  );
  //AND U251
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U251 (
    .O(y[104]),
    .I0(b[8]),
    .I1(a[6])
  );
  //OR U251bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U251bar (
    .O(ybar[104]),
    .I0(bbar[8]),
    .I1(abar[6])
  );
  //AND U252
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U252 (
    .O(y[103]),
    .I0(b[7]),
    .I1(a[6])
  );
  //OR U252bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U252bar (
    .O(ybar[103]),
    .I0(bbar[7]),
    .I1(abar[6])
  );
  //AND U253
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U253 (
    .O(y[102]),
    .I0(b[6]),
    .I1(a[6])
  );
  //OR U253bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U253bar (
    .O(ybar[102]),
    .I0(bbar[6]),
    .I1(abar[6])
  );
  //AND U254
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U254 (
    .O(y[101]),
    .I0(b[5]),
    .I1(a[6])
  );
  //OR U254bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U254bar (
    .O(ybar[101]),
    .I0(bbar[5]),
    .I1(abar[6])
  );
  //AND U255
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U255 (
    .O(y[100]),
    .I0(b[4]),
    .I1(a[6])
  );
  //OR U255bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U255bar (
    .O(ybar[100]),
    .I0(bbar[4]),
    .I1(abar[6])
  );
  //AND U256
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U256 (
    .O(y[0]),
    .I0(b[0]),
    .I1(a[0])
  );
  //OR U256bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U256bar (
    .O(ybar[0]),
    .I0(bbar[0]),
    .I1(abar[0])
  );
endmodule

module decode_11 ( in, out );

  input wire [7:0] in;
//input_done

  output wire [255:0] out;
//output_done

  wire [15:0] level1;
  wire [31:0] level2;
//wire_done

  CD2_44 cd_l1_1 ( .a(in[1]), .b(in[0]), .y(level1[3:0]) );
  CD2_43 cd_l1_2 ( .a(in[3]), .b(in[2]), .y(level1[7:4]) );
  CD2_42 cd_l1_3 ( .a(in[5]), .b(in[4]), .y(level1[11:8]) );
  CD2_41 cd_l1_4 ( .a(in[7]), .b(in[6]), .y(level1[15:12]) );
  CD4_22 cd_l2_1 ( .a(level1[7:4]), .b(level1[3:0]), .y(level2[15:0]) );
  CD4_21 cd_l2_2 ( .a(level1[15:12]), .b(level1[11:8]), .y(level2[31:16]) );
  CD16_11 cd_l3 ( .a(level2[31:16]), .b(level2[15:0]), .y(out) );
endmodule

module encode_11 ( in, out );

  input wire [255:0] in;
  wire [255:0] inbar;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
  assign inbar[8] = ~in[8];
  assign inbar[9] = ~in[9];
  assign inbar[10] = ~in[10];
  assign inbar[11] = ~in[11];
  assign inbar[12] = ~in[12];
  assign inbar[13] = ~in[13];
  assign inbar[14] = ~in[14];
  assign inbar[15] = ~in[15];
  assign inbar[16] = ~in[16];
  assign inbar[17] = ~in[17];
  assign inbar[18] = ~in[18];
  assign inbar[19] = ~in[19];
  assign inbar[20] = ~in[20];
  assign inbar[21] = ~in[21];
  assign inbar[22] = ~in[22];
  assign inbar[23] = ~in[23];
  assign inbar[24] = ~in[24];
  assign inbar[25] = ~in[25];
  assign inbar[26] = ~in[26];
  assign inbar[27] = ~in[27];
  assign inbar[28] = ~in[28];
  assign inbar[29] = ~in[29];
  assign inbar[30] = ~in[30];
  assign inbar[31] = ~in[31];
  assign inbar[32] = ~in[32];
  assign inbar[33] = ~in[33];
  assign inbar[34] = ~in[34];
  assign inbar[35] = ~in[35];
  assign inbar[36] = ~in[36];
  assign inbar[37] = ~in[37];
  assign inbar[38] = ~in[38];
  assign inbar[39] = ~in[39];
  assign inbar[40] = ~in[40];
  assign inbar[41] = ~in[41];
  assign inbar[42] = ~in[42];
  assign inbar[43] = ~in[43];
  assign inbar[44] = ~in[44];
  assign inbar[45] = ~in[45];
  assign inbar[46] = ~in[46];
  assign inbar[47] = ~in[47];
  assign inbar[48] = ~in[48];
  assign inbar[49] = ~in[49];
  assign inbar[50] = ~in[50];
  assign inbar[51] = ~in[51];
  assign inbar[52] = ~in[52];
  assign inbar[53] = ~in[53];
  assign inbar[54] = ~in[54];
  assign inbar[55] = ~in[55];
  assign inbar[56] = ~in[56];
  assign inbar[57] = ~in[57];
  assign inbar[58] = ~in[58];
  assign inbar[59] = ~in[59];
  assign inbar[60] = ~in[60];
  assign inbar[61] = ~in[61];
  assign inbar[62] = ~in[62];
  assign inbar[63] = ~in[63];
  assign inbar[64] = ~in[64];
  assign inbar[65] = ~in[65];
  assign inbar[66] = ~in[66];
  assign inbar[67] = ~in[67];
  assign inbar[68] = ~in[68];
  assign inbar[69] = ~in[69];
  assign inbar[70] = ~in[70];
  assign inbar[71] = ~in[71];
  assign inbar[72] = ~in[72];
  assign inbar[73] = ~in[73];
  assign inbar[74] = ~in[74];
  assign inbar[75] = ~in[75];
  assign inbar[76] = ~in[76];
  assign inbar[77] = ~in[77];
  assign inbar[78] = ~in[78];
  assign inbar[79] = ~in[79];
  assign inbar[80] = ~in[80];
  assign inbar[81] = ~in[81];
  assign inbar[82] = ~in[82];
  assign inbar[83] = ~in[83];
  assign inbar[84] = ~in[84];
  assign inbar[85] = ~in[85];
  assign inbar[86] = ~in[86];
  assign inbar[87] = ~in[87];
  assign inbar[88] = ~in[88];
  assign inbar[89] = ~in[89];
  assign inbar[90] = ~in[90];
  assign inbar[91] = ~in[91];
  assign inbar[92] = ~in[92];
  assign inbar[93] = ~in[93];
  assign inbar[94] = ~in[94];
  assign inbar[95] = ~in[95];
  assign inbar[96] = ~in[96];
  assign inbar[97] = ~in[97];
  assign inbar[98] = ~in[98];
  assign inbar[99] = ~in[99];
  assign inbar[100] = ~in[100];
  assign inbar[101] = ~in[101];
  assign inbar[102] = ~in[102];
  assign inbar[103] = ~in[103];
  assign inbar[104] = ~in[104];
  assign inbar[105] = ~in[105];
  assign inbar[106] = ~in[106];
  assign inbar[107] = ~in[107];
  assign inbar[108] = ~in[108];
  assign inbar[109] = ~in[109];
  assign inbar[110] = ~in[110];
  assign inbar[111] = ~in[111];
  assign inbar[112] = ~in[112];
  assign inbar[113] = ~in[113];
  assign inbar[114] = ~in[114];
  assign inbar[115] = ~in[115];
  assign inbar[116] = ~in[116];
  assign inbar[117] = ~in[117];
  assign inbar[118] = ~in[118];
  assign inbar[119] = ~in[119];
  assign inbar[120] = ~in[120];
  assign inbar[121] = ~in[121];
  assign inbar[122] = ~in[122];
  assign inbar[123] = ~in[123];
  assign inbar[124] = ~in[124];
  assign inbar[125] = ~in[125];
  assign inbar[126] = ~in[126];
  assign inbar[127] = ~in[127];
  assign inbar[128] = ~in[128];
  assign inbar[129] = ~in[129];
  assign inbar[130] = ~in[130];
  assign inbar[131] = ~in[131];
  assign inbar[132] = ~in[132];
  assign inbar[133] = ~in[133];
  assign inbar[134] = ~in[134];
  assign inbar[135] = ~in[135];
  assign inbar[136] = ~in[136];
  assign inbar[137] = ~in[137];
  assign inbar[138] = ~in[138];
  assign inbar[139] = ~in[139];
  assign inbar[140] = ~in[140];
  assign inbar[141] = ~in[141];
  assign inbar[142] = ~in[142];
  assign inbar[143] = ~in[143];
  assign inbar[144] = ~in[144];
  assign inbar[145] = ~in[145];
  assign inbar[146] = ~in[146];
  assign inbar[147] = ~in[147];
  assign inbar[148] = ~in[148];
  assign inbar[149] = ~in[149];
  assign inbar[150] = ~in[150];
  assign inbar[151] = ~in[151];
  assign inbar[152] = ~in[152];
  assign inbar[153] = ~in[153];
  assign inbar[154] = ~in[154];
  assign inbar[155] = ~in[155];
  assign inbar[156] = ~in[156];
  assign inbar[157] = ~in[157];
  assign inbar[158] = ~in[158];
  assign inbar[159] = ~in[159];
  assign inbar[160] = ~in[160];
  assign inbar[161] = ~in[161];
  assign inbar[162] = ~in[162];
  assign inbar[163] = ~in[163];
  assign inbar[164] = ~in[164];
  assign inbar[165] = ~in[165];
  assign inbar[166] = ~in[166];
  assign inbar[167] = ~in[167];
  assign inbar[168] = ~in[168];
  assign inbar[169] = ~in[169];
  assign inbar[170] = ~in[170];
  assign inbar[171] = ~in[171];
  assign inbar[172] = ~in[172];
  assign inbar[173] = ~in[173];
  assign inbar[174] = ~in[174];
  assign inbar[175] = ~in[175];
  assign inbar[176] = ~in[176];
  assign inbar[177] = ~in[177];
  assign inbar[178] = ~in[178];
  assign inbar[179] = ~in[179];
  assign inbar[180] = ~in[180];
  assign inbar[181] = ~in[181];
  assign inbar[182] = ~in[182];
  assign inbar[183] = ~in[183];
  assign inbar[184] = ~in[184];
  assign inbar[185] = ~in[185];
  assign inbar[186] = ~in[186];
  assign inbar[187] = ~in[187];
  assign inbar[188] = ~in[188];
  assign inbar[189] = ~in[189];
  assign inbar[190] = ~in[190];
  assign inbar[191] = ~in[191];
  assign inbar[192] = ~in[192];
  assign inbar[193] = ~in[193];
  assign inbar[194] = ~in[194];
  assign inbar[195] = ~in[195];
  assign inbar[196] = ~in[196];
  assign inbar[197] = ~in[197];
  assign inbar[198] = ~in[198];
  assign inbar[199] = ~in[199];
  assign inbar[200] = ~in[200];
  assign inbar[201] = ~in[201];
  assign inbar[202] = ~in[202];
  assign inbar[203] = ~in[203];
  assign inbar[204] = ~in[204];
  assign inbar[205] = ~in[205];
  assign inbar[206] = ~in[206];
  assign inbar[207] = ~in[207];
  assign inbar[208] = ~in[208];
  assign inbar[209] = ~in[209];
  assign inbar[210] = ~in[210];
  assign inbar[211] = ~in[211];
  assign inbar[212] = ~in[212];
  assign inbar[213] = ~in[213];
  assign inbar[214] = ~in[214];
  assign inbar[215] = ~in[215];
  assign inbar[216] = ~in[216];
  assign inbar[217] = ~in[217];
  assign inbar[218] = ~in[218];
  assign inbar[219] = ~in[219];
  assign inbar[220] = ~in[220];
  assign inbar[221] = ~in[221];
  assign inbar[222] = ~in[222];
  assign inbar[223] = ~in[223];
  assign inbar[224] = ~in[224];
  assign inbar[225] = ~in[225];
  assign inbar[226] = ~in[226];
  assign inbar[227] = ~in[227];
  assign inbar[228] = ~in[228];
  assign inbar[229] = ~in[229];
  assign inbar[230] = ~in[230];
  assign inbar[231] = ~in[231];
  assign inbar[232] = ~in[232];
  assign inbar[233] = ~in[233];
  assign inbar[234] = ~in[234];
  assign inbar[235] = ~in[235];
  assign inbar[236] = ~in[236];
  assign inbar[237] = ~in[237];
  assign inbar[238] = ~in[238];
  assign inbar[239] = ~in[239];
  assign inbar[240] = ~in[240];
  assign inbar[241] = ~in[241];
  assign inbar[242] = ~in[242];
  assign inbar[243] = ~in[243];
  assign inbar[244] = ~in[244];
  assign inbar[245] = ~in[245];
  assign inbar[246] = ~in[246];
  assign inbar[247] = ~in[247];
  assign inbar[248] = ~in[248];
  assign inbar[249] = ~in[249];
  assign inbar[250] = ~in[250];
  assign inbar[251] = ~in[251];
  assign inbar[252] = ~in[252];
  assign inbar[253] = ~in[253];
  assign inbar[254] = ~in[254];
  assign inbar[255] = ~in[255];
//input_done

  output wire [7:0] out;
  wire [7:0] outbar;
//output_done

  wire in_81;
  wire in_80;
  wire in_79;
  wire in_78;
  wire in_77;
  wire in_76;
  wire in_75;
  wire in_74;
  wire in_73;
  wire in_72;
  wire in_71;
  wire in_70;
  wire in_69;
  wire in_68;
  wire in_67;
  wire in_66;
  wire in_65;
  wire in_64;
  wire in_63;
  wire in_62;
  wire in_61;
  wire in_60;
  wire in_59;
  wire in_58;
  wire in_57;
  wire in_56;
  wire in_55;
  wire in_54;
  wire in_53;
  wire in_52;
  wire in_51;
  wire in_50;
  wire in_49;
  wire in_48;
  wire in_47;
  wire in_46;
  wire in_45;
  wire in_44;
  wire in_43;
  wire in_42;
  wire in_41;
  wire in_40;
  wire in_39;
  wire in_38;
  wire in_37;
  wire in_36;
  wire in_35;
  wire in_34;
  wire in_33;
  wire in_32;
  wire in_31;
  wire in_30;
  wire in_29;
  wire in_28;
  wire in_27;
  wire in_26;
  wire in_25;
  wire in_24;
  wire in_23;
  wire in_22;
  wire in_21;
  wire in_20;
  wire in_19;
  wire in_18;
  wire in_17;
  wire in_16;
  wire in_15;
  wire in_14;
  wire in_13;
  wire in_12;
  wire in_11;
  wire in_10;
  wire in_9;
  wire in_8;
  wire in_7;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_3;
  wire in_2;
  wire in_1;
  wire in_0;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire in_81bar;
  wire in_80bar;
  wire in_79bar;
  wire in_78bar;
  wire in_77bar;
  wire in_76bar;
  wire in_75bar;
  wire in_74bar;
  wire in_73bar;
  wire in_72bar;
  wire in_71bar;
  wire in_70bar;
  wire in_69bar;
  wire in_68bar;
  wire in_67bar;
  wire in_66bar;
  wire in_65bar;
  wire in_64bar;
  wire in_63bar;
  wire in_62bar;
  wire in_61bar;
  wire in_60bar;
  wire in_59bar;
  wire in_58bar;
  wire in_57bar;
  wire in_56bar;
  wire in_55bar;
  wire in_54bar;
  wire in_53bar;
  wire in_52bar;
  wire in_51bar;
  wire in_50bar;
  wire in_49bar;
  wire in_48bar;
  wire in_47bar;
  wire in_46bar;
  wire in_45bar;
  wire in_44bar;
  wire in_43bar;
  wire in_42bar;
  wire in_41bar;
  wire in_40bar;
  wire in_39bar;
  wire in_38bar;
  wire in_37bar;
  wire in_36bar;
  wire in_35bar;
  wire in_34bar;
  wire in_33bar;
  wire in_32bar;
  wire in_31bar;
  wire in_30bar;
  wire in_29bar;
  wire in_28bar;
  wire in_27bar;
  wire in_26bar;
  wire in_25bar;
  wire in_24bar;
  wire in_23bar;
  wire in_22bar;
  wire in_21bar;
  wire in_20bar;
  wire in_19bar;
  wire in_18bar;
  wire in_17bar;
  wire in_16bar;
  wire in_15bar;
  wire in_14bar;
  wire in_13bar;
  wire in_12bar;
  wire in_11bar;
  wire in_10bar;
  wire in_9bar;
  wire in_8bar;
  wire in_7bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_3bar;
  wire in_2bar;
  wire in_1bar;
  wire in_0bar;
  wire n487bar;
  wire n488bar;
  wire n489bar;
  wire n490bar;
  wire n491bar;
  wire n492bar;
  wire n493bar;
  wire n494bar;
  wire n495bar;
  wire n496bar;
  wire n497bar;
  wire n498bar;
  wire n499bar;
  wire n500bar;
  wire n501bar;
  wire n502bar;
  wire n503bar;
  wire n504bar;
  wire n505bar;
  wire n506bar;
  wire n507bar;
  wire n508bar;
  wire n509bar;
  wire n510bar;
  wire n511bar;
  wire n512bar;
  wire n513bar;
  wire n514bar;
  wire n515bar;
  wire n516bar;
  wire n517bar;
  wire n518bar;
  wire n519bar;
  wire n520bar;
  wire n521bar;
  wire n522bar;
  wire n523bar;
  wire n524bar;
  wire n525bar;
  wire n526bar;
  wire n527bar;
  wire n528bar;
  wire n529bar;
  wire n530bar;
  wire n531bar;
  wire n532bar;
  wire n533bar;
  wire n534bar;
  wire n535bar;
  wire n536bar;
  wire n537bar;
  wire n538bar;
  wire n539bar;
  wire n540bar;
  wire n541bar;
  wire n542bar;
  wire n543bar;
  wire n544bar;
  wire n545bar;
  wire n546bar;
  wire n547bar;
  wire n548bar;
  wire n549bar;
  wire n550bar;
  wire n551bar;
  wire n552bar;
  wire n553bar;
  wire n554bar;
  wire n555bar;
  wire n556bar;
  wire n557bar;
  wire n558bar;
  wire n559bar;
  wire n560bar;
  wire n561bar;
  wire n562bar;
  wire n563bar;
  wire n564bar;
  wire n565bar;
  wire n566bar;
  wire n567bar;
  wire n568bar;
  wire n569bar;
  wire n570bar;
  wire n571bar;
  wire n572bar;
  wire n573bar;
  wire n574bar;
  wire n575bar;
  wire n576bar;
  wire n577bar;
  wire n578bar;
  wire n579bar;
  wire n580bar;
  wire n581bar;
  wire n582bar;
  wire n583bar;
  wire n584bar;
  wire n585bar;
  wire n586bar;
  wire n587bar;
  wire n588bar;
  wire n589bar;
  wire n590bar;
  wire n591bar;
  wire n592bar;
  wire n593bar;
  wire n594bar;
  wire n595bar;
  wire n596bar;
  wire n597bar;
  wire n598bar;
  wire n599bar;
  wire n600bar;
  wire n601bar;
  wire n602bar;
  wire n603bar;
  wire n604bar;
  wire n605bar;
  wire n606bar;
  wire n607bar;
  wire n608bar;
  wire n609bar;
  wire n610bar;
  wire n611bar;
  wire n612bar;
  wire n613bar;
  wire n614bar;
  wire n615bar;
  wire n616bar;
  wire n617bar;
  wire n618bar;
  wire n619bar;
  wire n620bar;
  wire n621bar;
  wire n622bar;
  wire n623bar;
  wire n624bar;
  wire n625bar;
  wire n626bar;
  wire n627bar;
  wire n628bar;
  wire n629bar;
  wire n630bar;
  wire n631bar;
  wire n632bar;
  wire n633bar;
  wire n634bar;
  wire n635bar;
  wire n636bar;
  wire n637bar;
  wire n638bar;
  wire n639bar;
  wire n640bar;
  wire n641bar;
  wire n642bar;
  wire n643bar;
  wire n644bar;
  wire n645bar;
  wire n646bar;
  wire n647bar;
  wire n648bar;
  wire n649bar;
  wire n650bar;
  wire n651bar;
  wire n652bar;
  wire n653bar;
  wire n654bar;
  wire n655bar;
  wire n656bar;
  wire n657bar;
  wire n658bar;
  wire n659bar;
  wire n660bar;
  wire n661bar;
  wire n662bar;
  wire n663bar;
  wire n664bar;
  wire n665bar;
  wire n666bar;
  wire n667bar;
  wire n668bar;
  wire n669bar;
  wire n670bar;
  wire n671bar;
  wire n672bar;
  wire n673bar;
  wire n674bar;
  wire n675bar;
  wire n676bar;
  wire n677bar;
  wire n678bar;
  wire n679bar;
  wire n680bar;
  wire n681bar;
  wire n682bar;
  wire n683bar;
  wire n684bar;
  wire n685bar;
  wire n686bar;
  wire n687bar;
  wire n688bar;
  wire n689bar;
  wire n690bar;
  wire n691bar;
  wire n692bar;
  wire n693bar;
  wire n694bar;
  wire n695bar;
  wire n696bar;
  wire n697bar;
  wire n698bar;
  wire n699bar;
  wire n700bar;
  wire n701bar;
  wire n702bar;
  wire n703bar;
  wire n704bar;
  wire n705bar;
  wire n706bar;
  wire n707bar;
  wire n708bar;
  wire n709bar;
  wire n710bar;
  wire n711bar;
  wire n712bar;
  wire n713bar;
  wire n714bar;
  wire n715bar;
  wire n716bar;
  wire n717bar;
  wire n718bar;
  wire n719bar;
  wire n720bar;
  wire n721bar;
  wire n722bar;
  wire n723bar;
  wire n724bar;
  wire n725bar;
  wire n726bar;
  wire n727bar;
  wire n728bar;
  wire n729bar;
  wire n730bar;
  wire n731bar;
  wire n732bar;
  wire n733bar;
  wire n734bar;
  wire n735bar;
  wire n736bar;
  wire n737bar;
  wire n738bar;
  wire n739bar;
  wire n740bar;
  wire n741bar;
  wire n742bar;
  wire n743bar;
  wire n744bar;
  wire n745bar;
  wire n746bar;
  wire n747bar;
  wire n748bar;
  wire n749bar;
  wire n750bar;
  wire n751bar;
  wire n752bar;
  wire n753bar;
  wire n754bar;
  wire n755bar;
  wire n756bar;
  wire n757bar;
  wire n758bar;
  wire n759bar;
  wire n760bar;
  wire n761bar;
  wire n762bar;
  wire n763bar;
  wire n764bar;
  wire n765bar;
  wire n766bar;
  wire n767bar;
  wire n768bar;
  wire n769bar;
  wire n770bar;
  wire n771bar;
  wire n772bar;
  wire n773bar;
  wire n774bar;
  wire n775bar;
  wire n776bar;
  wire n777bar;
  wire n778bar;
  wire n779bar;
  wire n780bar;
  wire n781bar;
  wire n782bar;
  wire n783bar;
  wire n784bar;
  wire n785bar;
  wire n786bar;
  wire n787bar;
  wire n788bar;
  wire n789bar;
  wire n790bar;
  wire n791bar;
  wire n792bar;
  wire n793bar;
  wire n794bar;
  wire n795bar;
  wire n796bar;
  wire n797bar;
  wire n798bar;
  wire n799bar;
  wire n800bar;
  wire n801bar;
  wire n802bar;
  wire n803bar;
  wire n804bar;
  wire n805bar;
  wire n806bar;
  wire n807bar;
  wire n808bar;
  wire n809bar;
  wire n810bar;
  wire n811bar;
  wire n812bar;
  wire n813bar;
  wire n814bar;
  wire n815bar;
  wire n816bar;
  wire n817bar;
  wire n818bar;
  wire n819bar;
  wire n820bar;
  wire n821bar;
  wire n822bar;
  wire n823bar;
  wire n824bar;
  wire n825bar;
  wire n826bar;
  wire n827bar;
  wire n828bar;
  wire n829bar;
  wire n830bar;
  wire n831bar;
  wire n832bar;
  wire n833bar;
  wire n834bar;
  wire n835bar;
  wire n836bar;
  wire n837bar;
  wire n838bar;
  wire n839bar;
  wire n840bar;
  wire n841bar;
  wire n842bar;
  wire n843bar;
  wire n844bar;
  wire n845bar;
  wire n846bar;
  wire n847bar;
  wire n848bar;
  wire n849bar;
  wire n850bar;
  wire n851bar;
  wire n852bar;
  wire n853bar;
  wire n854bar;
  wire n855bar;
  wire n856bar;
  wire n857bar;
  wire n858bar;
  wire n859bar;
  wire n860bar;
  wire n861bar;
  wire n862bar;
  wire n863bar;
  wire n864bar;
  wire n865bar;
  wire n866bar;
  wire n867bar;
  wire n868bar;
  wire n869bar;
  wire n870bar;
  wire n871bar;
  wire n872bar;
  wire n873bar;
  wire n874bar;
  wire n875bar;
  wire n876bar;
  wire n877bar;
  wire n878bar;
  wire n879bar;
  wire n880bar;
  wire n881bar;
  wire n882bar;
  wire n883bar;
  wire n884bar;
  wire n885bar;
  wire n886bar;
  wire n887bar;
  wire n888bar;
  wire n889bar;
  wire n890bar;
  wire n891bar;
  wire n892bar;
  wire n893bar;
  wire n894bar;
  wire n895bar;
  wire n896bar;
  wire n897bar;
  wire n898bar;
  wire n899bar;
  wire n900bar;
  wire n901bar;
  wire n902bar;
  wire n903bar;
  wire n904bar;
  wire n905bar;
  wire n906bar;
  wire n907bar;
  wire n908bar;
  wire n909bar;
  wire n910bar;
  wire n911bar;
  wire n912bar;
  wire n913bar;
  wire n914bar;
  wire n915bar;
  wire n916bar;
  wire n917bar;
  wire n918bar;
  wire n919bar;
  wire n920bar;
  wire n921bar;
  wire n922bar;
  wire n923bar;
  wire n924bar;
  wire n925bar;
  wire n926bar;
  wire n927bar;
  wire n928bar;
  wire n929bar;
  wire n930bar;
  wire n931bar;
  wire n932bar;
  wire n933bar;
  wire n934bar;
  wire n935bar;
  wire n936bar;
  wire n937bar;
  wire n938bar;
  wire n939bar;
  wire n940bar;
  wire n941bar;
  wire n942bar;
  wire n943bar;
  wire n944bar;
  wire n945bar;
  wire n946bar;
  wire n947bar;
  wire n948bar;
  wire n949bar;
  wire n950bar;
  wire n951bar;
  wire n952bar;
  wire n953bar;
  wire n954bar;
  wire n955bar;
  wire n956bar;
  wire n957bar;
  wire n958bar;
  wire n959bar;
  wire n960bar;
  wire n961bar;
  wire n962bar;
  wire n963bar;
  wire n964bar;
  wire n965bar;
  wire n966bar;
  wire n967bar;
  wire n968bar;
  wire n969bar;
  wire n970bar;
  wire n971bar;
  wire n972bar;
//wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];
  //OR U1
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1 (
    .O(out[7]),
    .I0(n972),
    .I1(n971)
  );
  //AND U1bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1bar (
    .O(outbar[7]),
    .I0(n972bar),
    .I1(n971bar)
  );
  //OR U2
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2 (
    .O(n971),
    .I0(n970),
    .I1(n969)
  );
  //AND U2bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2bar (
    .O(n971bar),
    .I0(n970bar),
    .I1(n969bar)
  );
  //OR U3
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3 (
    .O(n969),
    .I0(n968),
    .I1(n967)
  );
  //AND U3bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3bar (
    .O(n969bar),
    .I0(n968bar),
    .I1(n967bar)
  );
  //OR U4
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4 (
    .O(n967),
    .I0(n966),
    .I1(n965)
  );
  //AND U4bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4bar (
    .O(n967bar),
    .I0(n966bar),
    .I1(n965bar)
  );
  //OR U5
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5 (
    .O(n968),
    .I0(n964),
    .I1(n963)
  );
  //AND U5bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5bar (
    .O(n968bar),
    .I0(n964bar),
    .I1(n963bar)
  );
  //OR U6
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6 (
    .O(n963),
    .I0(in[116]),
    .I1(n962)
  );
  //AND U6bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6bar (
    .O(n963bar),
    .I0(inbar[116]),
    .I1(n962bar)
  );
  //OR U7
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7 (
    .O(n970),
    .I0(n961),
    .I1(n960)
  );
  //AND U7bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7bar (
    .O(n970bar),
    .I0(n961bar),
    .I1(n960bar)
  );
  //OR U8
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8 (
    .O(n960),
    .I0(in[150]),
    .I1(in[127])
  );
  //AND U8bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8bar (
    .O(n960bar),
    .I0(inbar[150]),
    .I1(inbar[127])
  );
  //OR U9
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9 (
    .O(n961),
    .I0(in[160]),
    .I1(n959)
  );
  //AND U9bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9bar (
    .O(n961bar),
    .I0(inbar[160]),
    .I1(n959bar)
  );
  //OR U10
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10 (
    .O(n959),
    .I0(in[252]),
    .I1(in[168])
  );
  //AND U10bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10bar (
    .O(n959bar),
    .I0(inbar[252]),
    .I1(inbar[168])
  );
  //OR U11
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11 (
    .O(n972),
    .I0(n958),
    .I1(n957)
  );
  //AND U11bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11bar (
    .O(n972bar),
    .I0(n958bar),
    .I1(n957bar)
  );
  //OR U12
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12 (
    .O(n957),
    .I0(n956),
    .I1(n955)
  );
  //AND U12bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12bar (
    .O(n957bar),
    .I0(n956bar),
    .I1(n955bar)
  );
  //OR U13
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13 (
    .O(n955),
    .I0(in_17),
    .I1(in[96])
  );
  //AND U13bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13bar (
    .O(n955bar),
    .I0(in_17bar),
    .I1(inbar[96])
  );
  //OR U14
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14 (
    .O(n956),
    .I0(in_23),
    .I1(n954)
  );
  //AND U14bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14bar (
    .O(n956bar),
    .I0(in_23bar),
    .I1(n954bar)
  );
  //OR U15
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15 (
    .O(n954),
    .I0(in_31),
    .I1(in_26)
  );
  //AND U15bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15bar (
    .O(n954bar),
    .I0(in_31bar),
    .I1(in_26bar)
  );
  //OR U16
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16 (
    .O(n958),
    .I0(n953),
    .I1(n952)
  );
  //AND U16bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16bar (
    .O(n958bar),
    .I0(n953bar),
    .I1(n952bar)
  );
  //OR U17
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U17 (
    .O(n952),
    .I0(in_58),
    .I1(in_4)
  );
  //AND U17bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U17bar (
    .O(n952bar),
    .I0(in_58bar),
    .I1(in_4bar)
  );
  //OR U18
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U18 (
    .O(n953),
    .I0(in_59),
    .I1(n951)
  );
  //AND U18bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U18bar (
    .O(n953bar),
    .I0(in_59bar),
    .I1(n951bar)
  );
  //OR U19
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U19 (
    .O(n951),
    .I0(in_71),
    .I1(in_62)
  );
  //AND U19bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U19bar (
    .O(n951bar),
    .I0(in_71bar),
    .I1(in_62bar)
  );
  //OR U20
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U20 (
    .O(out[6]),
    .I0(n950),
    .I1(n949)
  );
  //AND U20bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U20bar (
    .O(outbar[6]),
    .I0(n950bar),
    .I1(n949bar)
  );
  //OR U21
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U21 (
    .O(n949),
    .I0(n948),
    .I1(n947)
  );
  //AND U21bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U21bar (
    .O(n949bar),
    .I0(n948bar),
    .I1(n947bar)
  );
  //OR U22
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U22 (
    .O(n947),
    .I0(n946),
    .I1(n945)
  );
  //AND U22bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U22bar (
    .O(n947bar),
    .I0(n946bar),
    .I1(n945bar)
  );
  //OR U23
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U23 (
    .O(n945),
    .I0(n944),
    .I1(n943)
  );
  //AND U23bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U23bar (
    .O(n945bar),
    .I0(n944bar),
    .I1(n943bar)
  );
  //OR U24
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U24 (
    .O(n946),
    .I0(n942),
    .I1(n941)
  );
  //AND U24bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U24bar (
    .O(n946bar),
    .I0(n942bar),
    .I1(n941bar)
  );
  //OR U25
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U25 (
    .O(n941),
    .I0(in[101]),
    .I1(n940)
  );
  //AND U25bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U25bar (
    .O(n941bar),
    .I0(inbar[101]),
    .I1(n940bar)
  );
  //OR U26
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U26 (
    .O(n948),
    .I0(n939),
    .I1(n938)
  );
  //AND U26bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U26bar (
    .O(n948bar),
    .I0(n939bar),
    .I1(n938bar)
  );
  //OR U27
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U27 (
    .O(n938),
    .I0(in[114]),
    .I1(in[104])
  );
  //AND U27bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U27bar (
    .O(n938bar),
    .I0(inbar[114]),
    .I1(inbar[104])
  );
  //OR U28
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U28 (
    .O(n939),
    .I0(in[128]),
    .I1(n937)
  );
  //AND U28bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U28bar (
    .O(n939bar),
    .I0(inbar[128]),
    .I1(n937bar)
  );
  //OR U29
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U29 (
    .O(n937),
    .I0(in[136]),
    .I1(in[134])
  );
  //AND U29bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U29bar (
    .O(n937bar),
    .I0(inbar[136]),
    .I1(inbar[134])
  );
  //OR U30
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U30 (
    .O(n950),
    .I0(n936),
    .I1(n935)
  );
  //AND U30bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U30bar (
    .O(n950bar),
    .I0(n936bar),
    .I1(n935bar)
  );
  //OR U31
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U31 (
    .O(n935),
    .I0(n934),
    .I1(n933)
  );
  //AND U31bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U31bar (
    .O(n935bar),
    .I0(n934bar),
    .I1(n933bar)
  );
  //OR U32
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U32 (
    .O(n933),
    .I0(in[177]),
    .I1(in[164])
  );
  //AND U32bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U32bar (
    .O(n933bar),
    .I0(inbar[177]),
    .I1(inbar[164])
  );
  //OR U33
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U33 (
    .O(n934),
    .I0(in[212]),
    .I1(n932)
  );
  //AND U33bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U33bar (
    .O(n934bar),
    .I0(inbar[212]),
    .I1(n932bar)
  );
  //OR U34
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U34 (
    .O(n932),
    .I0(in[248]),
    .I1(in[221])
  );
  //AND U34bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U34bar (
    .O(n932bar),
    .I0(inbar[248]),
    .I1(inbar[221])
  );
  //OR U35
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U35 (
    .O(n936),
    .I0(n931),
    .I1(n930)
  );
  //AND U35bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U35bar (
    .O(n936bar),
    .I0(n931bar),
    .I1(n930bar)
  );
  //OR U36
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U36 (
    .O(n930),
    .I0(in_18),
    .I1(in[93])
  );
  //AND U36bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U36bar (
    .O(n930bar),
    .I0(in_18bar),
    .I1(inbar[93])
  );
  //OR U37
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U37 (
    .O(n931),
    .I0(in_31),
    .I1(n929)
  );
  //AND U37bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U37bar (
    .O(n931bar),
    .I0(in_31bar),
    .I1(n929bar)
  );
  //OR U38
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U38 (
    .O(n929),
    .I0(in_7),
    .I1(in_39)
  );
  //AND U38bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U38bar (
    .O(n929bar),
    .I0(in_7bar),
    .I1(in_39bar)
  );
  //OR U39
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U39 (
    .O(out[5]),
    .I0(n928),
    .I1(n927)
  );
  //AND U39bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U39bar (
    .O(outbar[5]),
    .I0(n928bar),
    .I1(n927bar)
  );
  //OR U40
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U40 (
    .O(n927),
    .I0(n926),
    .I1(n925)
  );
  //AND U40bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U40bar (
    .O(n927bar),
    .I0(n926bar),
    .I1(n925bar)
  );
  //OR U41
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U41 (
    .O(n925),
    .I0(n924),
    .I1(n923)
  );
  //AND U41bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U41bar (
    .O(n925bar),
    .I0(n924bar),
    .I1(n923bar)
  );
  //OR U42
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U42 (
    .O(n923),
    .I0(n922),
    .I1(n921)
  );
  //AND U42bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U42bar (
    .O(n923bar),
    .I0(n922bar),
    .I1(n921bar)
  );
  //OR U43
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U43 (
    .O(n924),
    .I0(n940),
    .I1(n920)
  );
  //AND U43bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U43bar (
    .O(n924bar),
    .I0(n940bar),
    .I1(n920bar)
  );
  //OR U44
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U44 (
    .O(n920),
    .I0(in[111]),
    .I1(n919)
  );
  //AND U44bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U44bar (
    .O(n920bar),
    .I0(inbar[111]),
    .I1(n919bar)
  );
  //OR U45
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U45 (
    .O(n940),
    .I0(n918),
    .I1(n917)
  );
  //AND U45bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U45bar (
    .O(n940bar),
    .I0(n918bar),
    .I1(n917bar)
  );
  //OR U46
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U46 (
    .O(n917),
    .I0(n916),
    .I1(n915)
  );
  //AND U46bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U46bar (
    .O(n917bar),
    .I0(n916bar),
    .I1(n915bar)
  );
  //OR U47
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U47 (
    .O(n915),
    .I0(n914),
    .I1(n913)
  );
  //AND U47bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U47bar (
    .O(n915bar),
    .I0(n914bar),
    .I1(n913bar)
  );
  //OR U48
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U48 (
    .O(n913),
    .I0(in[140]),
    .I1(in[131])
  );
  //AND U48bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U48bar (
    .O(n913bar),
    .I0(inbar[140]),
    .I1(inbar[131])
  );
  //OR U49
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U49 (
    .O(n914),
    .I0(in[160]),
    .I1(in[144])
  );
  //AND U49bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U49bar (
    .O(n914bar),
    .I0(inbar[160]),
    .I1(inbar[144])
  );
  //OR U50
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U50 (
    .O(n916),
    .I0(n912),
    .I1(n911)
  );
  //AND U50bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U50bar (
    .O(n916bar),
    .I0(n912bar),
    .I1(n911bar)
  );
  //OR U51
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U51 (
    .O(n911),
    .I0(in[179]),
    .I1(in[174])
  );
  //AND U51bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U51bar (
    .O(n911bar),
    .I0(inbar[179]),
    .I1(inbar[174])
  );
  //OR U52
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U52 (
    .O(n912),
    .I0(in[188]),
    .I1(in[184])
  );
  //AND U52bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U52bar (
    .O(n912bar),
    .I0(inbar[188]),
    .I1(inbar[184])
  );
  //OR U53
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U53 (
    .O(n918),
    .I0(n910),
    .I1(n909)
  );
  //AND U53bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U53bar (
    .O(n918bar),
    .I0(n910bar),
    .I1(n909bar)
  );
  //OR U54
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U54 (
    .O(n909),
    .I0(n908),
    .I1(n907)
  );
  //AND U54bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U54bar (
    .O(n909bar),
    .I0(n908bar),
    .I1(n907bar)
  );
  //OR U55
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U55 (
    .O(n907),
    .I0(in[216]),
    .I1(in[200])
  );
  //AND U55bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U55bar (
    .O(n907bar),
    .I0(inbar[216]),
    .I1(inbar[200])
  );
  //OR U56
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U56 (
    .O(n908),
    .I0(in[228]),
    .I1(in[224])
  );
  //AND U56bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U56bar (
    .O(n908bar),
    .I0(inbar[228]),
    .I1(inbar[224])
  );
  //OR U57
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U57 (
    .O(n910),
    .I0(n906),
    .I1(n905)
  );
  //AND U57bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U57bar (
    .O(n910bar),
    .I0(n906bar),
    .I1(n905bar)
  );
  //OR U58
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U58 (
    .O(n905),
    .I0(in[247]),
    .I1(in[235])
  );
  //AND U58bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U58bar (
    .O(n905bar),
    .I0(inbar[247]),
    .I1(inbar[235])
  );
  //OR U59
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U59 (
    .O(n906),
    .I0(in_42),
    .I1(in[83])
  );
  //AND U59bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U59bar (
    .O(n906bar),
    .I0(in_42bar),
    .I1(inbar[83])
  );
  //OR U60
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U60 (
    .O(n926),
    .I0(n904),
    .I1(n903)
  );
  //AND U60bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U60bar (
    .O(n926bar),
    .I0(n904bar),
    .I1(n903bar)
  );
  //OR U61
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U61 (
    .O(n903),
    .I0(in[166]),
    .I1(in[123])
  );
  //AND U61bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U61bar (
    .O(n903bar),
    .I0(inbar[166]),
    .I1(inbar[123])
  );
  //OR U62
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U62 (
    .O(n904),
    .I0(in[170]),
    .I1(n902)
  );
  //AND U62bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U62bar (
    .O(n904bar),
    .I0(inbar[170]),
    .I1(n902bar)
  );
  //OR U63
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U63 (
    .O(n902),
    .I0(in[194]),
    .I1(in[183])
  );
  //AND U63bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U63bar (
    .O(n902bar),
    .I0(inbar[194]),
    .I1(inbar[183])
  );
  //OR U64
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U64 (
    .O(n928),
    .I0(n901),
    .I1(n900)
  );
  //AND U64bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U64bar (
    .O(n928bar),
    .I0(n901bar),
    .I1(n900bar)
  );
  //OR U65
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U65 (
    .O(n900),
    .I0(n899),
    .I1(n898)
  );
  //AND U65bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U65bar (
    .O(n900bar),
    .I0(n899bar),
    .I1(n898bar)
  );
  //OR U66
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U66 (
    .O(n898),
    .I0(in[241]),
    .I1(in[238])
  );
  //AND U66bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U66bar (
    .O(n898bar),
    .I0(inbar[241]),
    .I1(inbar[238])
  );
  //OR U67
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U67 (
    .O(n899),
    .I0(in[250]),
    .I1(n897)
  );
  //AND U67bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U67bar (
    .O(n899bar),
    .I0(inbar[250]),
    .I1(n897bar)
  );
  //OR U68
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U68 (
    .O(n897),
    .I0(in_24),
    .I1(in[84])
  );
  //AND U68bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U68bar (
    .O(n897bar),
    .I0(in_24bar),
    .I1(inbar[84])
  );
  //OR U69
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U69 (
    .O(n901),
    .I0(n896),
    .I1(n895)
  );
  //AND U69bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U69bar (
    .O(n901bar),
    .I0(n896bar),
    .I1(n895bar)
  );
  //OR U70
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U70 (
    .O(n895),
    .I0(in_41),
    .I1(in_29)
  );
  //AND U70bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U70bar (
    .O(n895bar),
    .I0(in_41bar),
    .I1(in_29bar)
  );
  //OR U71
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U71 (
    .O(n896),
    .I0(in_66),
    .I1(n894)
  );
  //AND U71bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U71bar (
    .O(n896bar),
    .I0(in_66bar),
    .I1(n894bar)
  );
  //OR U72
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U72 (
    .O(n894),
    .I0(in_76),
    .I1(in_71)
  );
  //AND U72bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U72bar (
    .O(n894bar),
    .I0(in_76bar),
    .I1(in_71bar)
  );
  //OR U73
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U73 (
    .O(out[4]),
    .I0(n893),
    .I1(n892)
  );
  //AND U73bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U73bar (
    .O(outbar[4]),
    .I0(n893bar),
    .I1(n892bar)
  );
  //OR U74
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U74 (
    .O(n892),
    .I0(n891),
    .I1(n890)
  );
  //AND U74bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U74bar (
    .O(n892bar),
    .I0(n891bar),
    .I1(n890bar)
  );
  //OR U75
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U75 (
    .O(n890),
    .I0(n889),
    .I1(n888)
  );
  //AND U75bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U75bar (
    .O(n890bar),
    .I0(n889bar),
    .I1(n888bar)
  );
  //OR U76
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U76 (
    .O(n888),
    .I0(n922),
    .I1(n887)
  );
  //AND U76bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U76bar (
    .O(n888bar),
    .I0(n922bar),
    .I1(n887bar)
  );
  //OR U77
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U77 (
    .O(n922),
    .I0(n886),
    .I1(n885)
  );
  //AND U77bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U77bar (
    .O(n922bar),
    .I0(n886bar),
    .I1(n885bar)
  );
  //OR U78
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U78 (
    .O(n885),
    .I0(n884),
    .I1(n883)
  );
  //AND U78bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U78bar (
    .O(n885bar),
    .I0(n884bar),
    .I1(n883bar)
  );
  //OR U79
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U79 (
    .O(n883),
    .I0(n882),
    .I1(n881)
  );
  //AND U79bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U79bar (
    .O(n883bar),
    .I0(n882bar),
    .I1(n881bar)
  );
  //OR U80
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U80 (
    .O(n881),
    .I0(in[118]),
    .I1(in[109])
  );
  //AND U80bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U80bar (
    .O(n881bar),
    .I0(inbar[118]),
    .I1(inbar[109])
  );
  //OR U81
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U81 (
    .O(n882),
    .I0(in[139]),
    .I1(in[120])
  );
  //AND U81bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U81bar (
    .O(n882bar),
    .I0(inbar[139]),
    .I1(inbar[120])
  );
  //OR U82
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U82 (
    .O(n884),
    .I0(n880),
    .I1(n879)
  );
  //AND U82bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U82bar (
    .O(n884bar),
    .I0(n880bar),
    .I1(n879bar)
  );
  //OR U83
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U83 (
    .O(n879),
    .I0(in[198]),
    .I1(in[154])
  );
  //AND U83bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U83bar (
    .O(n879bar),
    .I0(inbar[198]),
    .I1(inbar[154])
  );
  //OR U84
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U84 (
    .O(n880),
    .I0(in[210]),
    .I1(in[205])
  );
  //AND U84bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U84bar (
    .O(n880bar),
    .I0(inbar[210]),
    .I1(inbar[205])
  );
  //OR U85
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U85 (
    .O(n886),
    .I0(n878),
    .I1(n877)
  );
  //AND U85bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U85bar (
    .O(n886bar),
    .I0(n878bar),
    .I1(n877bar)
  );
  //OR U86
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U86 (
    .O(n877),
    .I0(n876),
    .I1(n875)
  );
  //AND U86bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U86bar (
    .O(n877bar),
    .I0(n876bar),
    .I1(n875bar)
  );
  //OR U87
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U87 (
    .O(n875),
    .I0(in[219]),
    .I1(in[217])
  );
  //AND U87bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U87bar (
    .O(n875bar),
    .I0(inbar[219]),
    .I1(inbar[217])
  );
  //OR U88
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U88 (
    .O(n876),
    .I0(in[86]),
    .I1(in[252])
  );
  //AND U88bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U88bar (
    .O(n876bar),
    .I0(inbar[86]),
    .I1(inbar[252])
  );
  //OR U89
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U89 (
    .O(n878),
    .I0(n874),
    .I1(n873)
  );
  //AND U89bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U89bar (
    .O(n878bar),
    .I0(n874bar),
    .I1(n873bar)
  );
  //OR U90
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U90 (
    .O(n873),
    .I0(in_40),
    .I1(in[91])
  );
  //AND U90bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U90bar (
    .O(n873bar),
    .I0(in_40bar),
    .I1(inbar[91])
  );
  //OR U91
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U91 (
    .O(n874),
    .I0(in_8),
    .I1(in_46)
  );
  //AND U91bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U91bar (
    .O(n874bar),
    .I0(in_8bar),
    .I1(in_46bar)
  );
  //OR U92
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U92 (
    .O(n889),
    .I0(n872),
    .I1(n871)
  );
  //AND U92bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U92bar (
    .O(n889bar),
    .I0(n872bar),
    .I1(n871bar)
  );
  //OR U93
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U93 (
    .O(n871),
    .I0(in[117]),
    .I1(n943)
  );
  //AND U93bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U93bar (
    .O(n871bar),
    .I0(inbar[117]),
    .I1(n943bar)
  );
  //OR U94
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U94 (
    .O(n943),
    .I0(n870),
    .I1(n869)
  );
  //AND U94bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U94bar (
    .O(n943bar),
    .I0(n870bar),
    .I1(n869bar)
  );
  //OR U95
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U95 (
    .O(n869),
    .I0(n868),
    .I1(n867)
  );
  //AND U95bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U95bar (
    .O(n869bar),
    .I0(n868bar),
    .I1(n867bar)
  );
  //OR U96
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U96 (
    .O(n867),
    .I0(n866),
    .I1(n865)
  );
  //AND U96bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U96bar (
    .O(n867bar),
    .I0(n866bar),
    .I1(n865bar)
  );
  //OR U97
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U97 (
    .O(n865),
    .I0(n864),
    .I1(n863)
  );
  //AND U97bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U97bar (
    .O(n865bar),
    .I0(n864bar),
    .I1(n863bar)
  );
  //OR U98
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U98 (
    .O(n866),
    .I0(in[108]),
    .I1(n919)
  );
  //AND U98bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U98bar (
    .O(n866bar),
    .I0(inbar[108]),
    .I1(n919bar)
  );
  //OR U99
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U99 (
    .O(n919),
    .I0(n862),
    .I1(n861)
  );
  //AND U99bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U99bar (
    .O(n919bar),
    .I0(n862bar),
    .I1(n861bar)
  );
  //OR U100
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U100 (
    .O(n861),
    .I0(n860),
    .I1(n859)
  );
  //AND U100bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U100bar (
    .O(n861bar),
    .I0(n860bar),
    .I1(n859bar)
  );
  //OR U101
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U101 (
    .O(n859),
    .I0(n858),
    .I1(n857)
  );
  //AND U101bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U101bar (
    .O(n859bar),
    .I0(n858bar),
    .I1(n857bar)
  );
  //OR U102
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U102 (
    .O(n857),
    .I0(in[119]),
    .I1(in[105])
  );
  //AND U102bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U102bar (
    .O(n857bar),
    .I0(inbar[119]),
    .I1(inbar[105])
  );
  //OR U103
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U103 (
    .O(n858),
    .I0(in[186]),
    .I1(in[175])
  );
  //AND U103bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U103bar (
    .O(n858bar),
    .I0(inbar[186]),
    .I1(inbar[175])
  );
  //OR U104
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U104 (
    .O(n860),
    .I0(n856),
    .I1(n855)
  );
  //AND U104bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U104bar (
    .O(n860bar),
    .I0(n856bar),
    .I1(n855bar)
  );
  //OR U105
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U105 (
    .O(n855),
    .I0(in[202]),
    .I1(in[193])
  );
  //AND U105bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U105bar (
    .O(n855bar),
    .I0(inbar[202]),
    .I1(inbar[193])
  );
  //OR U106
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U106 (
    .O(n856),
    .I0(in[225]),
    .I1(in[208])
  );
  //AND U106bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U106bar (
    .O(n856bar),
    .I0(inbar[225]),
    .I1(inbar[208])
  );
  //OR U107
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U107 (
    .O(n862),
    .I0(n854),
    .I1(n853)
  );
  //AND U107bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U107bar (
    .O(n862bar),
    .I0(n854bar),
    .I1(n853bar)
  );
  //OR U108
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U108 (
    .O(n853),
    .I0(n852),
    .I1(n851)
  );
  //AND U108bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U108bar (
    .O(n853bar),
    .I0(n852bar),
    .I1(n851bar)
  );
  //OR U109
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U109 (
    .O(n851),
    .I0(in_1),
    .I1(in[85])
  );
  //AND U109bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U109bar (
    .O(n851bar),
    .I0(in_1bar),
    .I1(inbar[85])
  );
  //OR U110
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U110 (
    .O(n852),
    .I0(in_23),
    .I1(in_19)
  );
  //AND U110bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U110bar (
    .O(n852bar),
    .I0(in_23bar),
    .I1(in_19bar)
  );
  //OR U111
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U111 (
    .O(n854),
    .I0(n850),
    .I1(n849)
  );
  //AND U111bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U111bar (
    .O(n854bar),
    .I0(n850bar),
    .I1(n849bar)
  );
  //OR U112
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U112 (
    .O(n849),
    .I0(in_43),
    .I1(in_33)
  );
  //AND U112bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U112bar (
    .O(n849bar),
    .I0(in_43bar),
    .I1(in_33bar)
  );
  //OR U113
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U113 (
    .O(n850),
    .I0(in_63),
    .I1(in_44)
  );
  //AND U113bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U113bar (
    .O(n850bar),
    .I0(in_63bar),
    .I1(in_44bar)
  );
  //OR U114
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U114 (
    .O(n868),
    .I0(n848),
    .I1(n847)
  );
  //AND U114bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U114bar (
    .O(n868bar),
    .I0(n848bar),
    .I1(n847bar)
  );
  //OR U115
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U115 (
    .O(n847),
    .I0(in[141]),
    .I1(in[112])
  );
  //AND U115bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U115bar (
    .O(n847bar),
    .I0(inbar[141]),
    .I1(inbar[112])
  );
  //OR U116
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U116 (
    .O(n848),
    .I0(in[147]),
    .I1(n846)
  );
  //AND U116bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U116bar (
    .O(n848bar),
    .I0(inbar[147]),
    .I1(n846bar)
  );
  //OR U117
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U117 (
    .O(n846),
    .I0(in[181]),
    .I1(in[167])
  );
  //AND U117bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U117bar (
    .O(n846bar),
    .I0(inbar[181]),
    .I1(inbar[167])
  );
  //OR U118
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U118 (
    .O(n870),
    .I0(n845),
    .I1(n844)
  );
  //AND U118bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U118bar (
    .O(n870bar),
    .I0(n845bar),
    .I1(n844bar)
  );
  //OR U119
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U119 (
    .O(n844),
    .I0(n843),
    .I1(n842)
  );
  //AND U119bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U119bar (
    .O(n844bar),
    .I0(n843bar),
    .I1(n842bar)
  );
  //OR U120
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U120 (
    .O(n842),
    .I0(in[229]),
    .I1(in[201])
  );
  //AND U120bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U120bar (
    .O(n842bar),
    .I0(inbar[229]),
    .I1(inbar[201])
  );
  //OR U121
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U121 (
    .O(n843),
    .I0(in[237]),
    .I1(n841)
  );
  //AND U121bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U121bar (
    .O(n843bar),
    .I0(inbar[237]),
    .I1(n841bar)
  );
  //OR U122
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U122 (
    .O(n841),
    .I0(in[94]),
    .I1(in[253])
  );
  //AND U122bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U122bar (
    .O(n841bar),
    .I0(inbar[94]),
    .I1(inbar[253])
  );
  //OR U123
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U123 (
    .O(n845),
    .I0(n840),
    .I1(n839)
  );
  //AND U123bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U123bar (
    .O(n845bar),
    .I0(n840bar),
    .I1(n839bar)
  );
  //OR U124
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U124 (
    .O(n839),
    .I0(in_21),
    .I1(in[96])
  );
  //AND U124bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U124bar (
    .O(n839bar),
    .I0(in_21bar),
    .I1(inbar[96])
  );
  //OR U125
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U125 (
    .O(n840),
    .I0(in_25),
    .I1(n838)
  );
  //AND U125bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U125bar (
    .O(n840bar),
    .I0(in_25bar),
    .I1(n838bar)
  );
  //OR U126
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U126 (
    .O(n838),
    .I0(in_81),
    .I1(in_45)
  );
  //AND U126bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U126bar (
    .O(n838bar),
    .I0(in_81bar),
    .I1(in_45bar)
  );
  //OR U127
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U127 (
    .O(n891),
    .I0(n837),
    .I1(n836)
  );
  //AND U127bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U127bar (
    .O(n891bar),
    .I0(n837bar),
    .I1(n836bar)
  );
  //OR U128
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U128 (
    .O(n836),
    .I0(in[142]),
    .I1(in[124])
  );
  //AND U128bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U128bar (
    .O(n836bar),
    .I0(inbar[142]),
    .I1(inbar[124])
  );
  //OR U129
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U129 (
    .O(n837),
    .I0(in[150]),
    .I1(n835)
  );
  //AND U129bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U129bar (
    .O(n837bar),
    .I0(inbar[150]),
    .I1(n835bar)
  );
  //OR U130
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U130 (
    .O(n835),
    .I0(in[172]),
    .I1(in[155])
  );
  //AND U130bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U130bar (
    .O(n835bar),
    .I0(inbar[172]),
    .I1(inbar[155])
  );
  //OR U131
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U131 (
    .O(n893),
    .I0(n834),
    .I1(n833)
  );
  //AND U131bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U131bar (
    .O(n893bar),
    .I0(n834bar),
    .I1(n833bar)
  );
  //OR U132
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U132 (
    .O(n833),
    .I0(n832),
    .I1(n831)
  );
  //AND U132bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U132bar (
    .O(n833bar),
    .I0(n832bar),
    .I1(n831bar)
  );
  //OR U133
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U133 (
    .O(n831),
    .I0(in[196]),
    .I1(in[173])
  );
  //AND U133bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U133bar (
    .O(n831bar),
    .I0(inbar[196]),
    .I1(inbar[173])
  );
  //OR U134
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U134 (
    .O(n832),
    .I0(in[222]),
    .I1(n830)
  );
  //AND U134bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U134bar (
    .O(n832bar),
    .I0(inbar[222]),
    .I1(n830bar)
  );
  //OR U135
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U135 (
    .O(n830),
    .I0(in[227]),
    .I1(in[226])
  );
  //AND U135bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U135bar (
    .O(n830bar),
    .I0(inbar[227]),
    .I1(inbar[226])
  );
  //OR U136
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U136 (
    .O(n834),
    .I0(n829),
    .I1(n828)
  );
  //AND U136bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U136bar (
    .O(n834bar),
    .I0(n829bar),
    .I1(n828bar)
  );
  //OR U137
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U137 (
    .O(n828),
    .I0(in[249]),
    .I1(in[231])
  );
  //AND U137bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U137bar (
    .O(n828bar),
    .I0(inbar[249]),
    .I1(inbar[231])
  );
  //OR U138
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U138 (
    .O(n829),
    .I0(in_28),
    .I1(n827)
  );
  //AND U138bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U138bar (
    .O(n829bar),
    .I0(in_28bar),
    .I1(n827bar)
  );
  //OR U139
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U139 (
    .O(n827),
    .I0(in_52),
    .I1(in_47)
  );
  //AND U139bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U139bar (
    .O(n827bar),
    .I0(in_52bar),
    .I1(in_47bar)
  );
  //OR U140
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U140 (
    .O(out[3]),
    .I0(n826),
    .I1(n825)
  );
  //AND U140bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U140bar (
    .O(outbar[3]),
    .I0(n826bar),
    .I1(n825bar)
  );
  //OR U141
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U141 (
    .O(n825),
    .I0(n824),
    .I1(n823)
  );
  //AND U141bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U141bar (
    .O(n825bar),
    .I0(n824bar),
    .I1(n823bar)
  );
  //OR U142
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U142 (
    .O(n823),
    .I0(n822),
    .I1(n821)
  );
  //AND U142bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U142bar (
    .O(n823bar),
    .I0(n822bar),
    .I1(n821bar)
  );
  //OR U143
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U143 (
    .O(n821),
    .I0(n820),
    .I1(n819)
  );
  //AND U143bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U143bar (
    .O(n821bar),
    .I0(n820bar),
    .I1(n819bar)
  );
  //OR U144
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U144 (
    .O(n822),
    .I0(n964),
    .I1(n818)
  );
  //AND U144bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U144bar (
    .O(n822bar),
    .I0(n964bar),
    .I1(n818bar)
  );
  //OR U145
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U145 (
    .O(n818),
    .I0(in[118]),
    .I1(n817)
  );
  //AND U145bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U145bar (
    .O(n818bar),
    .I0(inbar[118]),
    .I1(n817bar)
  );
  //OR U146
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U146 (
    .O(n964),
    .I0(n816),
    .I1(n815)
  );
  //AND U146bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U146bar (
    .O(n964bar),
    .I0(n816bar),
    .I1(n815bar)
  );
  //OR U147
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U147 (
    .O(n815),
    .I0(n814),
    .I1(n813)
  );
  //AND U147bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U147bar (
    .O(n815bar),
    .I0(n814bar),
    .I1(n813bar)
  );
  //OR U148
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U148 (
    .O(n813),
    .I0(n812),
    .I1(n811)
  );
  //AND U148bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U148bar (
    .O(n813bar),
    .I0(n812bar),
    .I1(n811bar)
  );
  //OR U149
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U149 (
    .O(n811),
    .I0(in[122]),
    .I1(in[111])
  );
  //AND U149bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U149bar (
    .O(n811bar),
    .I0(inbar[122]),
    .I1(inbar[111])
  );
  //OR U150
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U150 (
    .O(n812),
    .I0(in[154]),
    .I1(in[151])
  );
  //AND U150bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U150bar (
    .O(n812bar),
    .I0(inbar[154]),
    .I1(inbar[151])
  );
  //OR U151
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U151 (
    .O(n814),
    .I0(n810),
    .I1(n809)
  );
  //AND U151bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U151bar (
    .O(n814bar),
    .I0(n810bar),
    .I1(n809bar)
  );
  //OR U152
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U152 (
    .O(n809),
    .I0(in[187]),
    .I1(in[177])
  );
  //AND U152bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U152bar (
    .O(n809bar),
    .I0(inbar[187]),
    .I1(inbar[177])
  );
  //OR U153
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U153 (
    .O(n810),
    .I0(in[200]),
    .I1(in[192])
  );
  //AND U153bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U153bar (
    .O(n810bar),
    .I0(inbar[200]),
    .I1(inbar[192])
  );
  //OR U154
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U154 (
    .O(n816),
    .I0(n808),
    .I1(n807)
  );
  //AND U154bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U154bar (
    .O(n816bar),
    .I0(n808bar),
    .I1(n807bar)
  );
  //OR U155
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U155 (
    .O(n807),
    .I0(n806),
    .I1(n805)
  );
  //AND U155bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U155bar (
    .O(n807bar),
    .I0(n806bar),
    .I1(n805bar)
  );
  //OR U156
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U156 (
    .O(n805),
    .I0(in[225]),
    .I1(in[207])
  );
  //AND U156bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U156bar (
    .O(n805bar),
    .I0(inbar[225]),
    .I1(inbar[207])
  );
  //OR U157
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U157 (
    .O(n806),
    .I0(in[98]),
    .I1(in[226])
  );
  //AND U157bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U157bar (
    .O(n806bar),
    .I0(inbar[98]),
    .I1(inbar[226])
  );
  //OR U158
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U158 (
    .O(n808),
    .I0(n804),
    .I1(n803)
  );
  //AND U158bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U158bar (
    .O(n808bar),
    .I0(n804bar),
    .I1(n803bar)
  );
  //OR U159
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U159 (
    .O(n803),
    .I0(in_20),
    .I1(in_16)
  );
  //AND U159bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U159bar (
    .O(n803bar),
    .I0(in_20bar),
    .I1(in_16bar)
  );
  //OR U160
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U160 (
    .O(n804),
    .I0(in_55),
    .I1(in_45)
  );
  //AND U160bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U160bar (
    .O(n804bar),
    .I0(in_55bar),
    .I1(in_45bar)
  );
  //OR U161
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U161 (
    .O(n824),
    .I0(n802),
    .I1(n801)
  );
  //AND U161bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U161bar (
    .O(n824bar),
    .I0(n802bar),
    .I1(n801bar)
  );
  //OR U162
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U162 (
    .O(n801),
    .I0(in[162]),
    .I1(in[149])
  );
  //AND U162bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U162bar (
    .O(n801bar),
    .I0(inbar[162]),
    .I1(inbar[149])
  );
  //OR U163
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U163 (
    .O(n802),
    .I0(in[163]),
    .I1(n800)
  );
  //AND U163bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U163bar (
    .O(n802bar),
    .I0(inbar[163]),
    .I1(n800bar)
  );
  //OR U164
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U164 (
    .O(n800),
    .I0(in[191]),
    .I1(in[189])
  );
  //AND U164bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U164bar (
    .O(n800bar),
    .I0(inbar[191]),
    .I1(inbar[189])
  );
  //OR U165
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U165 (
    .O(n826),
    .I0(n799),
    .I1(n798)
  );
  //AND U165bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U165bar (
    .O(n826bar),
    .I0(n799bar),
    .I1(n798bar)
  );
  //OR U166
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U166 (
    .O(n798),
    .I0(n797),
    .I1(n796)
  );
  //AND U166bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U166bar (
    .O(n798bar),
    .I0(n797bar),
    .I1(n796bar)
  );
  //OR U167
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U167 (
    .O(n796),
    .I0(in[212]),
    .I1(in[193])
  );
  //AND U167bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U167bar (
    .O(n796bar),
    .I0(inbar[212]),
    .I1(inbar[193])
  );
  //OR U168
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U168 (
    .O(n797),
    .I0(in[238]),
    .I1(n795)
  );
  //AND U168bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U168bar (
    .O(n797bar),
    .I0(inbar[238]),
    .I1(n795bar)
  );
  //OR U169
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U169 (
    .O(n795),
    .I0(in[88]),
    .I1(in[247])
  );
  //AND U169bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U169bar (
    .O(n795bar),
    .I0(inbar[88]),
    .I1(inbar[247])
  );
  //OR U170
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U170 (
    .O(n799),
    .I0(n794),
    .I1(n793)
  );
  //AND U170bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U170bar (
    .O(n799bar),
    .I0(n794bar),
    .I1(n793bar)
  );
  //OR U171
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U171 (
    .O(n793),
    .I0(in[94]),
    .I1(in[92])
  );
  //AND U171bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U171bar (
    .O(n793bar),
    .I0(inbar[94]),
    .I1(inbar[92])
  );
  //OR U172
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U172 (
    .O(n794),
    .I0(in_52),
    .I1(n792)
  );
  //AND U172bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U172bar (
    .O(n794bar),
    .I0(in_52bar),
    .I1(n792bar)
  );
  //OR U173
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U173 (
    .O(n792),
    .I0(in_70),
    .I1(in_67)
  );
  //AND U173bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U173bar (
    .O(n792bar),
    .I0(in_70bar),
    .I1(in_67bar)
  );
  //OR U174
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U174 (
    .O(out[2]),
    .I0(n791),
    .I1(n790)
  );
  //AND U174bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U174bar (
    .O(outbar[2]),
    .I0(n791bar),
    .I1(n790bar)
  );
  //OR U175
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U175 (
    .O(n790),
    .I0(n789),
    .I1(n788)
  );
  //AND U175bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U175bar (
    .O(n790bar),
    .I0(n789bar),
    .I1(n788bar)
  );
  //OR U176
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U176 (
    .O(n788),
    .I0(n787),
    .I1(n786)
  );
  //AND U176bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U176bar (
    .O(n788bar),
    .I0(n787bar),
    .I1(n786bar)
  );
  //OR U177
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U177 (
    .O(n786),
    .I0(n819),
    .I1(n785)
  );
  //AND U177bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U177bar (
    .O(n786bar),
    .I0(n819bar),
    .I1(n785bar)
  );
  //OR U178
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U178 (
    .O(n819),
    .I0(n784),
    .I1(n783)
  );
  //AND U178bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U178bar (
    .O(n819bar),
    .I0(n784bar),
    .I1(n783bar)
  );
  //OR U179
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U179 (
    .O(n783),
    .I0(n782),
    .I1(n781)
  );
  //AND U179bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U179bar (
    .O(n783bar),
    .I0(n782bar),
    .I1(n781bar)
  );
  //OR U180
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U180 (
    .O(n781),
    .I0(n780),
    .I1(n779)
  );
  //AND U180bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U180bar (
    .O(n781bar),
    .I0(n780bar),
    .I1(n779bar)
  );
  //OR U181
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U181 (
    .O(n779),
    .I0(n962),
    .I1(n778)
  );
  //AND U181bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U181bar (
    .O(n779bar),
    .I0(n962bar),
    .I1(n778bar)
  );
  //OR U182
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U182 (
    .O(n962),
    .I0(n777),
    .I1(n776)
  );
  //AND U182bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U182bar (
    .O(n962bar),
    .I0(n777bar),
    .I1(n776bar)
  );
  //OR U183
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U183 (
    .O(n776),
    .I0(n775),
    .I1(n774)
  );
  //AND U183bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U183bar (
    .O(n776bar),
    .I0(n775bar),
    .I1(n774bar)
  );
  //OR U184
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U184 (
    .O(n774),
    .I0(n773),
    .I1(n772)
  );
  //AND U184bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U184bar (
    .O(n774bar),
    .I0(n773bar),
    .I1(n772bar)
  );
  //OR U185
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U185 (
    .O(n772),
    .I0(in[131]),
    .I1(in[120])
  );
  //AND U185bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U185bar (
    .O(n772bar),
    .I0(inbar[131]),
    .I1(inbar[120])
  );
  //OR U186
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U186 (
    .O(n773),
    .I0(in[153]),
    .I1(in[147])
  );
  //AND U186bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U186bar (
    .O(n773bar),
    .I0(inbar[153]),
    .I1(inbar[147])
  );
  //OR U187
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U187 (
    .O(n775),
    .I0(n771),
    .I1(n770)
  );
  //AND U187bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U187bar (
    .O(n775bar),
    .I0(n771bar),
    .I1(n770bar)
  );
  //OR U188
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U188 (
    .O(n770),
    .I0(in[170]),
    .I1(in[156])
  );
  //AND U188bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U188bar (
    .O(n770bar),
    .I0(inbar[170]),
    .I1(inbar[156])
  );
  //OR U189
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U189 (
    .O(n771),
    .I0(in[223]),
    .I1(in[190])
  );
  //AND U189bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U189bar (
    .O(n771bar),
    .I0(inbar[223]),
    .I1(inbar[190])
  );
  //OR U190
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U190 (
    .O(n777),
    .I0(n769),
    .I1(n768)
  );
  //AND U190bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U190bar (
    .O(n777bar),
    .I0(n769bar),
    .I1(n768bar)
  );
  //OR U191
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U191 (
    .O(n768),
    .I0(n767),
    .I1(n766)
  );
  //AND U191bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U191bar (
    .O(n768bar),
    .I0(n767bar),
    .I1(n766bar)
  );
  //OR U192
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U192 (
    .O(n766),
    .I0(in[236]),
    .I1(in[230])
  );
  //AND U192bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U192bar (
    .O(n766bar),
    .I0(inbar[236]),
    .I1(inbar[230])
  );
  //OR U193
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U193 (
    .O(n767),
    .I0(in[85]),
    .I1(in[240])
  );
  //AND U193bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U193bar (
    .O(n767bar),
    .I0(inbar[85]),
    .I1(inbar[240])
  );
  //OR U194
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U194 (
    .O(n769),
    .I0(n765),
    .I1(n764)
  );
  //AND U194bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U194bar (
    .O(n769bar),
    .I0(n765bar),
    .I1(n764bar)
  );
  //OR U195
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U195 (
    .O(n764),
    .I0(in_12),
    .I1(in[90])
  );
  //AND U195bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U195bar (
    .O(n764bar),
    .I0(in_12bar),
    .I1(inbar[90])
  );
  //OR U196
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U196 (
    .O(n765),
    .I0(in_39),
    .I1(in_28)
  );
  //AND U196bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U196bar (
    .O(n765bar),
    .I0(in_39bar),
    .I1(in_28bar)
  );
  //OR U197
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U197 (
    .O(n780),
    .I0(in[109]),
    .I1(n763)
  );
  //AND U197bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U197bar (
    .O(n780bar),
    .I0(inbar[109]),
    .I1(n763bar)
  );
  //OR U198
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U198 (
    .O(n782),
    .I0(n762),
    .I1(n761)
  );
  //AND U198bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U198bar (
    .O(n782bar),
    .I0(n762bar),
    .I1(n761bar)
  );
  //OR U199
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U199 (
    .O(n761),
    .I0(in[138]),
    .I1(in[129])
  );
  //AND U199bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U199bar (
    .O(n761bar),
    .I0(inbar[138]),
    .I1(inbar[129])
  );
  //OR U200
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U200 (
    .O(n762),
    .I0(in[157]),
    .I1(n760)
  );
  //AND U200bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U200bar (
    .O(n762bar),
    .I0(inbar[157]),
    .I1(n760bar)
  );
  //OR U201
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U201 (
    .O(n760),
    .I0(in[182]),
    .I1(in[167])
  );
  //AND U201bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U201bar (
    .O(n760bar),
    .I0(inbar[182]),
    .I1(inbar[167])
  );
  //OR U202
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U202 (
    .O(n784),
    .I0(n759),
    .I1(n758)
  );
  //AND U202bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U202bar (
    .O(n784bar),
    .I0(n759bar),
    .I1(n758bar)
  );
  //OR U203
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U203 (
    .O(n758),
    .I0(n757),
    .I1(n756)
  );
  //AND U203bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U203bar (
    .O(n758bar),
    .I0(n757bar),
    .I1(n756bar)
  );
  //OR U204
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U204 (
    .O(n756),
    .I0(in[195]),
    .I1(in[184])
  );
  //AND U204bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U204bar (
    .O(n756bar),
    .I0(inbar[195]),
    .I1(inbar[184])
  );
  //OR U205
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U205 (
    .O(n757),
    .I0(in[196]),
    .I1(n755)
  );
  //AND U205bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U205bar (
    .O(n757bar),
    .I0(inbar[196]),
    .I1(n755bar)
  );
  //OR U206
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U206 (
    .O(n755),
    .I0(in[215]),
    .I1(in[209])
  );
  //AND U206bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U206bar (
    .O(n755bar),
    .I0(inbar[215]),
    .I1(inbar[209])
  );
  //OR U207
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U207 (
    .O(n759),
    .I0(n754),
    .I1(n753)
  );
  //AND U207bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U207bar (
    .O(n759bar),
    .I0(n754bar),
    .I1(n753bar)
  );
  //OR U208
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U208 (
    .O(n753),
    .I0(in[93]),
    .I1(in[233])
  );
  //AND U208bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U208bar (
    .O(n753bar),
    .I0(inbar[93]),
    .I1(inbar[233])
  );
  //OR U209
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U209 (
    .O(n754),
    .I0(in_1),
    .I1(n752)
  );
  //AND U209bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U209bar (
    .O(n754bar),
    .I0(in_1bar),
    .I1(n752bar)
  );
  //OR U210
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U210 (
    .O(n752),
    .I0(in_69),
    .I1(in_66)
  );
  //AND U210bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U210bar (
    .O(n752bar),
    .I0(in_69bar),
    .I1(in_66bar)
  );
  //OR U211
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U211 (
    .O(n787),
    .I0(n966),
    .I1(n751)
  );
  //AND U211bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U211bar (
    .O(n787bar),
    .I0(n966bar),
    .I1(n751bar)
  );
  //OR U212
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U212 (
    .O(n751),
    .I0(in[134]),
    .I1(n750)
  );
  //AND U212bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U212bar (
    .O(n751bar),
    .I0(inbar[134]),
    .I1(n750bar)
  );
  //OR U213
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U213 (
    .O(n966),
    .I0(n749),
    .I1(n748)
  );
  //AND U213bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U213bar (
    .O(n966bar),
    .I0(n749bar),
    .I1(n748bar)
  );
  //OR U214
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U214 (
    .O(n748),
    .I0(n747),
    .I1(n746)
  );
  //AND U214bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U214bar (
    .O(n748bar),
    .I0(n747bar),
    .I1(n746bar)
  );
  //OR U215
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U215 (
    .O(n746),
    .I0(n745),
    .I1(n744)
  );
  //AND U215bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U215bar (
    .O(n746bar),
    .I0(n745bar),
    .I1(n744bar)
  );
  //OR U216
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U216 (
    .O(n744),
    .I0(in[136]),
    .I1(in[121])
  );
  //AND U216bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U216bar (
    .O(n744bar),
    .I0(inbar[136]),
    .I1(inbar[121])
  );
  //OR U217
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U217 (
    .O(n745),
    .I0(in[186]),
    .I1(in[174])
  );
  //AND U217bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U217bar (
    .O(n745bar),
    .I0(inbar[186]),
    .I1(inbar[174])
  );
  //OR U218
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U218 (
    .O(n747),
    .I0(n743),
    .I1(n742)
  );
  //AND U218bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U218bar (
    .O(n747bar),
    .I0(n743bar),
    .I1(n742bar)
  );
  //OR U219
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U219 (
    .O(n742),
    .I0(in[198]),
    .I1(in[197])
  );
  //AND U219bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U219bar (
    .O(n742bar),
    .I0(inbar[198]),
    .I1(inbar[197])
  );
  //OR U220
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U220 (
    .O(n743),
    .I0(in[214]),
    .I1(in[199])
  );
  //AND U220bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U220bar (
    .O(n743bar),
    .I0(inbar[214]),
    .I1(inbar[199])
  );
  //OR U221
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U221 (
    .O(n749),
    .I0(n741),
    .I1(n740)
  );
  //AND U221bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U221bar (
    .O(n749bar),
    .I0(n741bar),
    .I1(n740bar)
  );
  //OR U222
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U222 (
    .O(n740),
    .I0(n739),
    .I1(n738)
  );
  //AND U222bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U222bar (
    .O(n740bar),
    .I0(n739bar),
    .I1(n738bar)
  );
  //OR U223
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U223 (
    .O(n738),
    .I0(in[231]),
    .I1(in[220])
  );
  //AND U223bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U223bar (
    .O(n738bar),
    .I0(inbar[231]),
    .I1(inbar[220])
  );
  //OR U224
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U224 (
    .O(n739),
    .I0(in_25),
    .I1(in[245])
  );
  //AND U224bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U224bar (
    .O(n739bar),
    .I0(in_25bar),
    .I1(inbar[245])
  );
  //OR U225
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U225 (
    .O(n741),
    .I0(n737),
    .I1(n736)
  );
  //AND U225bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U225bar (
    .O(n741bar),
    .I0(n737bar),
    .I1(n736bar)
  );
  //OR U226
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U226 (
    .O(n736),
    .I0(in_53),
    .I1(in_29)
  );
  //AND U226bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U226bar (
    .O(n736bar),
    .I0(in_53bar),
    .I1(in_29bar)
  );
  //OR U227
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U227 (
    .O(n737),
    .I0(in_79),
    .I1(in_74)
  );
  //AND U227bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U227bar (
    .O(n737bar),
    .I0(in_79bar),
    .I1(in_74bar)
  );
  //OR U228
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U228 (
    .O(n789),
    .I0(n735),
    .I1(n734)
  );
  //AND U228bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U228bar (
    .O(n789bar),
    .I0(n735bar),
    .I1(n734bar)
  );
  //OR U229
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U229 (
    .O(n734),
    .I0(in[152]),
    .I1(in[140])
  );
  //AND U229bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U229bar (
    .O(n734bar),
    .I0(inbar[152]),
    .I1(inbar[140])
  );
  //OR U230
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U230 (
    .O(n735),
    .I0(in[155]),
    .I1(n733)
  );
  //AND U230bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U230bar (
    .O(n735bar),
    .I0(inbar[155]),
    .I1(n733bar)
  );
  //OR U231
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U231 (
    .O(n733),
    .I0(in[166]),
    .I1(in[165])
  );
  //AND U231bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U231bar (
    .O(n733bar),
    .I0(inbar[166]),
    .I1(inbar[165])
  );
  //OR U232
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U232 (
    .O(n791),
    .I0(n732),
    .I1(n731)
  );
  //AND U232bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U232bar (
    .O(n791bar),
    .I0(n732bar),
    .I1(n731bar)
  );
  //OR U233
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U233 (
    .O(n731),
    .I0(n730),
    .I1(n729)
  );
  //AND U233bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U233bar (
    .O(n731bar),
    .I0(n730bar),
    .I1(n729bar)
  );
  //OR U234
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U234 (
    .O(n729),
    .I0(in[202]),
    .I1(in[185])
  );
  //AND U234bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U234bar (
    .O(n729bar),
    .I0(inbar[202]),
    .I1(inbar[185])
  );
  //OR U235
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U235 (
    .O(n730),
    .I0(in[211]),
    .I1(n728)
  );
  //AND U235bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U235bar (
    .O(n730bar),
    .I0(inbar[211]),
    .I1(n728bar)
  );
  //OR U236
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U236 (
    .O(n728),
    .I0(in[255]),
    .I1(in[253])
  );
  //AND U236bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U236bar (
    .O(n728bar),
    .I0(inbar[255]),
    .I1(inbar[253])
  );
  //OR U237
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U237 (
    .O(n732),
    .I0(n727),
    .I1(n726)
  );
  //AND U237bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U237bar (
    .O(n732bar),
    .I0(n727bar),
    .I1(n726bar)
  );
  //OR U238
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U238 (
    .O(n726),
    .I0(in_35),
    .I1(in_15)
  );
  //AND U238bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U238bar (
    .O(n726bar),
    .I0(in_35bar),
    .I1(in_15bar)
  );
  //OR U239
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U239 (
    .O(n727),
    .I0(in_36),
    .I1(n725)
  );
  //AND U239bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U239bar (
    .O(n727bar),
    .I0(in_36bar),
    .I1(n725bar)
  );
  //OR U240
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U240 (
    .O(n725),
    .I0(in_48),
    .I1(in_40)
  );
  //AND U240bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U240bar (
    .O(n725bar),
    .I0(in_48bar),
    .I1(in_40bar)
  );
  //OR U241
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U241 (
    .O(out[1]),
    .I0(n724),
    .I1(n723)
  );
  //AND U241bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U241bar (
    .O(outbar[1]),
    .I0(n724bar),
    .I1(n723bar)
  );
  //OR U242
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U242 (
    .O(n723),
    .I0(n722),
    .I1(n721)
  );
  //AND U242bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U242bar (
    .O(n723bar),
    .I0(n722bar),
    .I1(n721bar)
  );
  //OR U243
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U243 (
    .O(n721),
    .I0(n720),
    .I1(n719)
  );
  //AND U243bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U243bar (
    .O(n721bar),
    .I0(n720bar),
    .I1(n719bar)
  );
  //OR U244
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U244 (
    .O(n719),
    .I0(n921),
    .I1(n887)
  );
  //AND U244bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U244bar (
    .O(n719bar),
    .I0(n921bar),
    .I1(n887bar)
  );
  //OR U245
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U245 (
    .O(n887),
    .I0(n718),
    .I1(n717)
  );
  //AND U245bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U245bar (
    .O(n887bar),
    .I0(n718bar),
    .I1(n717bar)
  );
  //OR U246
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U246 (
    .O(n717),
    .I0(n716),
    .I1(n715)
  );
  //AND U246bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U246bar (
    .O(n717bar),
    .I0(n716bar),
    .I1(n715bar)
  );
  //OR U247
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U247 (
    .O(n715),
    .I0(n714),
    .I1(n713)
  );
  //AND U247bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U247bar (
    .O(n715bar),
    .I0(n714bar),
    .I1(n713bar)
  );
  //OR U248
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U248 (
    .O(n713),
    .I0(in[116]),
    .I1(in[110])
  );
  //AND U248bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U248bar (
    .O(n713bar),
    .I0(inbar[116]),
    .I1(inbar[110])
  );
  //OR U249
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U249 (
    .O(n714),
    .I0(in[133]),
    .I1(in[130])
  );
  //AND U249bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U249bar (
    .O(n714bar),
    .I0(inbar[133]),
    .I1(inbar[130])
  );
  //OR U250
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U250 (
    .O(n716),
    .I0(n712),
    .I1(n711)
  );
  //AND U250bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U250bar (
    .O(n716bar),
    .I0(n712bar),
    .I1(n711bar)
  );
  //OR U251
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U251 (
    .O(n711),
    .I0(in[203]),
    .I1(in[135])
  );
  //AND U251bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U251bar (
    .O(n711bar),
    .I0(inbar[203]),
    .I1(inbar[135])
  );
  //OR U252
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U252 (
    .O(n712),
    .I0(in[232]),
    .I1(in[223])
  );
  //AND U252bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U252bar (
    .O(n712bar),
    .I0(inbar[232]),
    .I1(inbar[223])
  );
  //OR U253
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U253 (
    .O(n718),
    .I0(n710),
    .I1(n709)
  );
  //AND U253bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U253bar (
    .O(n718bar),
    .I0(n710bar),
    .I1(n709bar)
  );
  //OR U254
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U254 (
    .O(n709),
    .I0(n708),
    .I1(n707)
  );
  //AND U254bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U254bar (
    .O(n709bar),
    .I0(n708bar),
    .I1(n707bar)
  );
  //OR U255
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U255 (
    .O(n707),
    .I0(in[255]),
    .I1(in[233])
  );
  //AND U255bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U255bar (
    .O(n707bar),
    .I0(inbar[255]),
    .I1(inbar[233])
  );
  //OR U256
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U256 (
    .O(n708),
    .I0(in_53),
    .I1(in_34)
  );
  //AND U256bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U256bar (
    .O(n708bar),
    .I0(in_53bar),
    .I1(in_34bar)
  );
  //OR U257
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U257 (
    .O(n710),
    .I0(n706),
    .I1(n705)
  );
  //AND U257bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U257bar (
    .O(n710bar),
    .I0(n706bar),
    .I1(n705bar)
  );
  //OR U258
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U258 (
    .O(n705),
    .I0(in_57),
    .I1(in_55)
  );
  //AND U258bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U258bar (
    .O(n705bar),
    .I0(in_57bar),
    .I1(in_55bar)
  );
  //OR U259
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U259 (
    .O(n706),
    .I0(in_68),
    .I1(in_67)
  );
  //AND U259bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U259bar (
    .O(n706bar),
    .I0(in_68bar),
    .I1(in_67bar)
  );
  //OR U260
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U260 (
    .O(n921),
    .I0(n704),
    .I1(n703)
  );
  //AND U260bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U260bar (
    .O(n921bar),
    .I0(n704bar),
    .I1(n703bar)
  );
  //OR U261
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U261 (
    .O(n703),
    .I0(n702),
    .I1(n701)
  );
  //AND U261bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U261bar (
    .O(n703bar),
    .I0(n702bar),
    .I1(n701bar)
  );
  //OR U262
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U262 (
    .O(n701),
    .I0(n700),
    .I1(n699)
  );
  //AND U262bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U262bar (
    .O(n701bar),
    .I0(n700bar),
    .I1(n699bar)
  );
  //OR U263
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U263 (
    .O(n699),
    .I0(n944),
    .I1(n872)
  );
  //AND U263bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U263bar (
    .O(n699bar),
    .I0(n944bar),
    .I1(n872bar)
  );
  //OR U264
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U264 (
    .O(n872),
    .I0(n698),
    .I1(n697)
  );
  //AND U264bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U264bar (
    .O(n872bar),
    .I0(n698bar),
    .I1(n697bar)
  );
  //OR U265
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U265 (
    .O(n697),
    .I0(n696),
    .I1(n695)
  );
  //AND U265bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U265bar (
    .O(n697bar),
    .I0(n696bar),
    .I1(n695bar)
  );
  //OR U266
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U266 (
    .O(n695),
    .I0(n694),
    .I1(n693)
  );
  //AND U266bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U266bar (
    .O(n695bar),
    .I0(n694bar),
    .I1(n693bar)
  );
  //OR U267
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U267 (
    .O(n693),
    .I0(in[121]),
    .I1(in[102])
  );
  //AND U267bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U267bar (
    .O(n693bar),
    .I0(inbar[121]),
    .I1(inbar[102])
  );
  //OR U268
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U268 (
    .O(n694),
    .I0(in[162]),
    .I1(in[161])
  );
  //AND U268bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U268bar (
    .O(n694bar),
    .I0(inbar[162]),
    .I1(inbar[161])
  );
  //OR U269
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U269 (
    .O(n696),
    .I0(n692),
    .I1(n691)
  );
  //AND U269bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U269bar (
    .O(n696bar),
    .I0(n692bar),
    .I1(n691bar)
  );
  //OR U270
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U270 (
    .O(n691),
    .I0(in[192]),
    .I1(in[178])
  );
  //AND U270bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U270bar (
    .O(n691bar),
    .I0(inbar[192]),
    .I1(inbar[178])
  );
  //OR U271
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U271 (
    .O(n692),
    .I0(in[244]),
    .I1(in[209])
  );
  //AND U271bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U271bar (
    .O(n692bar),
    .I0(inbar[244]),
    .I1(inbar[209])
  );
  //OR U272
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U272 (
    .O(n698),
    .I0(n690),
    .I1(n689)
  );
  //AND U272bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U272bar (
    .O(n698bar),
    .I0(n690bar),
    .I1(n689bar)
  );
  //OR U273
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U273 (
    .O(n689),
    .I0(n688),
    .I1(n687)
  );
  //AND U273bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U273bar (
    .O(n689bar),
    .I0(n688bar),
    .I1(n687bar)
  );
  //OR U274
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U274 (
    .O(n687),
    .I0(in[90]),
    .I1(in[254])
  );
  //AND U274bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U274bar (
    .O(n687bar),
    .I0(inbar[90]),
    .I1(inbar[254])
  );
  //OR U275
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U275 (
    .O(n688),
    .I0(in_36),
    .I1(in_32)
  );
  //AND U275bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U275bar (
    .O(n688bar),
    .I0(in_36bar),
    .I1(in_32bar)
  );
  //OR U276
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U276 (
    .O(n690),
    .I0(n686),
    .I1(n685)
  );
  //AND U276bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U276bar (
    .O(n690bar),
    .I0(n686bar),
    .I1(n685bar)
  );
  //OR U277
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U277 (
    .O(n685),
    .I0(in_62),
    .I1(in_37)
  );
  //AND U277bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U277bar (
    .O(n685bar),
    .I0(in_62bar),
    .I1(in_37bar)
  );
  //OR U278
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U278 (
    .O(n686),
    .I0(in_75),
    .I1(in_73)
  );
  //AND U278bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U278bar (
    .O(n686bar),
    .I0(in_75bar),
    .I1(in_73bar)
  );
  //OR U279
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U279 (
    .O(n944),
    .I0(n684),
    .I1(n683)
  );
  //AND U279bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U279bar (
    .O(n944bar),
    .I0(n684bar),
    .I1(n683bar)
  );
  //OR U280
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U280 (
    .O(n683),
    .I0(n682),
    .I1(n681)
  );
  //AND U280bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U280bar (
    .O(n683bar),
    .I0(n682bar),
    .I1(n681bar)
  );
  //OR U281
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U281 (
    .O(n681),
    .I0(n680),
    .I1(n679)
  );
  //AND U281bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U281bar (
    .O(n681bar),
    .I0(n680bar),
    .I1(n679bar)
  );
  //OR U282
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U282 (
    .O(n679),
    .I0(in[171]),
    .I1(in[153])
  );
  //AND U282bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U282bar (
    .O(n679bar),
    .I0(inbar[171]),
    .I1(inbar[153])
  );
  //OR U283
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U283 (
    .O(n680),
    .I0(in[187]),
    .I1(in[176])
  );
  //AND U283bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U283bar (
    .O(n680bar),
    .I0(inbar[187]),
    .I1(inbar[176])
  );
  //OR U284
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U284 (
    .O(n682),
    .I0(n678),
    .I1(n677)
  );
  //AND U284bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U284bar (
    .O(n682bar),
    .I0(n678bar),
    .I1(n677bar)
  );
  //OR U285
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U285 (
    .O(n677),
    .I0(in[245]),
    .I1(in[211])
  );
  //AND U285bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U285bar (
    .O(n677bar),
    .I0(inbar[245]),
    .I1(inbar[211])
  );
  //OR U286
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U286 (
    .O(n678),
    .I0(in[97]),
    .I1(in[88])
  );
  //AND U286bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U286bar (
    .O(n678bar),
    .I0(inbar[97]),
    .I1(inbar[88])
  );
  //OR U287
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U287 (
    .O(n684),
    .I0(n676),
    .I1(n675)
  );
  //AND U287bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U287bar (
    .O(n684bar),
    .I0(n676bar),
    .I1(n675bar)
  );
  //OR U288
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U288 (
    .O(n675),
    .I0(n674),
    .I1(n673)
  );
  //AND U288bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U288bar (
    .O(n675bar),
    .I0(n674bar),
    .I1(n673bar)
  );
  //OR U289
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U289 (
    .O(n673),
    .I0(in_10),
    .I1(in_0)
  );
  //AND U289bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U289bar (
    .O(n673bar),
    .I0(in_10bar),
    .I1(in_0bar)
  );
  //OR U290
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U290 (
    .O(n674),
    .I0(in_59),
    .I1(in_5)
  );
  //AND U290bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U290bar (
    .O(n674bar),
    .I0(in_59bar),
    .I1(in_5bar)
  );
  //OR U291
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U291 (
    .O(n676),
    .I0(n672),
    .I1(n671)
  );
  //AND U291bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U291bar (
    .O(n676bar),
    .I0(n672bar),
    .I1(n671bar)
  );
  //OR U292
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U292 (
    .O(n671),
    .I0(in_60),
    .I1(in_6)
  );
  //AND U292bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U292bar (
    .O(n671bar),
    .I0(in_60bar),
    .I1(in_6bar)
  );
  //OR U293
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U293 (
    .O(n672),
    .I0(in_77),
    .I1(in_69)
  );
  //AND U293bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U293bar (
    .O(n672bar),
    .I0(in_77bar),
    .I1(in_69bar)
  );
  //OR U294
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U294 (
    .O(n700),
    .I0(in[113]),
    .I1(n864)
  );
  //AND U294bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U294bar (
    .O(n700bar),
    .I0(inbar[113]),
    .I1(n864bar)
  );
  //OR U295
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U295 (
    .O(n864),
    .I0(n670),
    .I1(n669)
  );
  //AND U295bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U295bar (
    .O(n864bar),
    .I0(n670bar),
    .I1(n669bar)
  );
  //OR U296
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U296 (
    .O(n669),
    .I0(n668),
    .I1(n667)
  );
  //AND U296bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U296bar (
    .O(n669bar),
    .I0(n668bar),
    .I1(n667bar)
  );
  //OR U297
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U297 (
    .O(n667),
    .I0(n666),
    .I1(n665)
  );
  //AND U297bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U297bar (
    .O(n667bar),
    .I0(n666bar),
    .I1(n665bar)
  );
  //OR U298
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U298 (
    .O(n665),
    .I0(in[125]),
    .I1(in[107])
  );
  //AND U298bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U298bar (
    .O(n665bar),
    .I0(inbar[125]),
    .I1(inbar[107])
  );
  //OR U299
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U299 (
    .O(n666),
    .I0(in[138]),
    .I1(in[126])
  );
  //AND U299bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U299bar (
    .O(n666bar),
    .I0(inbar[138]),
    .I1(inbar[126])
  );
  //OR U300
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U300 (
    .O(n668),
    .I0(n664),
    .I1(n663)
  );
  //AND U300bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U300bar (
    .O(n668bar),
    .I0(n664bar),
    .I1(n663bar)
  );
  //OR U301
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U301 (
    .O(n663),
    .I0(in[189]),
    .I1(in[143])
  );
  //AND U301bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U301bar (
    .O(n663bar),
    .I0(inbar[189]),
    .I1(inbar[143])
  );
  //OR U302
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U302 (
    .O(n664),
    .I0(in[99]),
    .I1(in[214])
  );
  //AND U302bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U302bar (
    .O(n664bar),
    .I0(inbar[99]),
    .I1(inbar[214])
  );
  //OR U303
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U303 (
    .O(n670),
    .I0(n662),
    .I1(n661)
  );
  //AND U303bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U303bar (
    .O(n670bar),
    .I0(n662bar),
    .I1(n661bar)
  );
  //OR U304
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U304 (
    .O(n661),
    .I0(n660),
    .I1(n659)
  );
  //AND U304bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U304bar (
    .O(n661bar),
    .I0(n660bar),
    .I1(n659bar)
  );
  //OR U305
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U305 (
    .O(n659),
    .I0(in_15),
    .I1(in_12)
  );
  //AND U305bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U305bar (
    .O(n659bar),
    .I0(in_15bar),
    .I1(in_12bar)
  );
  //OR U306
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U306 (
    .O(n660),
    .I0(in_20),
    .I1(in_2)
  );
  //AND U306bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U306bar (
    .O(n660bar),
    .I0(in_20bar),
    .I1(in_2bar)
  );
  //OR U307
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U307 (
    .O(n662),
    .I0(n658),
    .I1(n657)
  );
  //AND U307bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U307bar (
    .O(n662bar),
    .I0(n658bar),
    .I1(n657bar)
  );
  //OR U308
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U308 (
    .O(n657),
    .I0(in_30),
    .I1(in_3)
  );
  //AND U308bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U308bar (
    .O(n657bar),
    .I0(in_30bar),
    .I1(in_3bar)
  );
  //OR U309
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U309 (
    .O(n658),
    .I0(in_4),
    .I1(in_38)
  );
  //AND U309bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U309bar (
    .O(n658bar),
    .I0(in_4bar),
    .I1(in_38bar)
  );
  //OR U310
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U310 (
    .O(n702),
    .I0(n656),
    .I1(n655)
  );
  //AND U310bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U310bar (
    .O(n702bar),
    .I0(n656bar),
    .I1(n655bar)
  );
  //OR U311
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U311 (
    .O(n655),
    .I0(in[148]),
    .I1(in[137])
  );
  //AND U311bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U311bar (
    .O(n655bar),
    .I0(inbar[148]),
    .I1(inbar[137])
  );
  //OR U312
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U312 (
    .O(n656),
    .I0(in[149]),
    .I1(n654)
  );
  //AND U312bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U312bar (
    .O(n656bar),
    .I0(inbar[149]),
    .I1(n654bar)
  );
  //OR U313
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U313 (
    .O(n654),
    .I0(in[195]),
    .I1(in[190])
  );
  //AND U313bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U313bar (
    .O(n654bar),
    .I0(inbar[195]),
    .I1(inbar[190])
  );
  //OR U314
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U314 (
    .O(n704),
    .I0(n653),
    .I1(n652)
  );
  //AND U314bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U314bar (
    .O(n704bar),
    .I0(n653bar),
    .I1(n652bar)
  );
  //OR U315
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U315 (
    .O(n652),
    .I0(n651),
    .I1(n650)
  );
  //AND U315bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U315bar (
    .O(n652bar),
    .I0(n651bar),
    .I1(n650bar)
  );
  //OR U316
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U316 (
    .O(n650),
    .I0(in[98]),
    .I1(in[197])
  );
  //AND U316bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U316bar (
    .O(n650bar),
    .I0(inbar[98]),
    .I1(inbar[197])
  );
  //OR U317
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U317 (
    .O(n651),
    .I0(in_11),
    .I1(n649)
  );
  //AND U317bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U317bar (
    .O(n651bar),
    .I0(in_11bar),
    .I1(n649bar)
  );
  //OR U318
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U318 (
    .O(n649),
    .I0(in_26),
    .I1(in_14)
  );
  //AND U318bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U318bar (
    .O(n649bar),
    .I0(in_26bar),
    .I1(in_14bar)
  );
  //OR U319
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U319 (
    .O(n653),
    .I0(n648),
    .I1(n647)
  );
  //AND U319bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U319bar (
    .O(n653bar),
    .I0(n648bar),
    .I1(n647bar)
  );
  //OR U320
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U320 (
    .O(n647),
    .I0(in_35),
    .I1(in_27)
  );
  //AND U320bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U320bar (
    .O(n647bar),
    .I0(in_35bar),
    .I1(in_27bar)
  );
  //OR U321
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U321 (
    .O(n648),
    .I0(in_50),
    .I1(n646)
  );
  //AND U321bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U321bar (
    .O(n648bar),
    .I0(in_50bar),
    .I1(n646bar)
  );
  //OR U322
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U322 (
    .O(n646),
    .I0(in_78),
    .I1(in_61)
  );
  //AND U322bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U322bar (
    .O(n646bar),
    .I0(in_78bar),
    .I1(in_61bar)
  );
  //OR U323
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U323 (
    .O(n720),
    .I0(n942),
    .I1(n645)
  );
  //AND U323bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U323bar (
    .O(n720bar),
    .I0(n942bar),
    .I1(n645bar)
  );
  //OR U324
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U324 (
    .O(n645),
    .I0(in[106]),
    .I1(n863)
  );
  //AND U324bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U324bar (
    .O(n645bar),
    .I0(inbar[106]),
    .I1(n863bar)
  );
  //OR U325
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U325 (
    .O(n863),
    .I0(n644),
    .I1(n643)
  );
  //AND U325bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U325bar (
    .O(n863bar),
    .I0(n644bar),
    .I1(n643bar)
  );
  //OR U326
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U326 (
    .O(n643),
    .I0(n642),
    .I1(n641)
  );
  //AND U326bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U326bar (
    .O(n643bar),
    .I0(n642bar),
    .I1(n641bar)
  );
  //OR U327
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U327 (
    .O(n641),
    .I0(n640),
    .I1(n639)
  );
  //AND U327bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U327bar (
    .O(n641bar),
    .I0(n640bar),
    .I1(n639bar)
  );
  //OR U328
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U328 (
    .O(n639),
    .I0(in[127]),
    .I1(in[122])
  );
  //AND U328bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U328bar (
    .O(n639bar),
    .I0(inbar[127]),
    .I1(inbar[122])
  );
  //OR U329
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U329 (
    .O(n640),
    .I0(in[156]),
    .I1(in[132])
  );
  //AND U329bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U329bar (
    .O(n640bar),
    .I0(inbar[156]),
    .I1(inbar[132])
  );
  //OR U330
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U330 (
    .O(n642),
    .I0(n638),
    .I1(n637)
  );
  //AND U330bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U330bar (
    .O(n642bar),
    .I0(n638bar),
    .I1(n637bar)
  );
  //OR U331
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U331 (
    .O(n637),
    .I0(in[159]),
    .I1(in[157])
  );
  //AND U331bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U331bar (
    .O(n637bar),
    .I0(inbar[159]),
    .I1(inbar[157])
  );
  //OR U332
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U332 (
    .O(n638),
    .I0(in[185]),
    .I1(in[169])
  );
  //AND U332bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U332bar (
    .O(n638bar),
    .I0(inbar[185]),
    .I1(inbar[169])
  );
  //OR U333
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U333 (
    .O(n644),
    .I0(n636),
    .I1(n635)
  );
  //AND U333bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U333bar (
    .O(n644bar),
    .I0(n636bar),
    .I1(n635bar)
  );
  //OR U334
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U334 (
    .O(n635),
    .I0(n634),
    .I1(n633)
  );
  //AND U334bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U334bar (
    .O(n635bar),
    .I0(n634bar),
    .I1(n633bar)
  );
  //OR U335
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U335 (
    .O(n633),
    .I0(in[239]),
    .I1(in[218])
  );
  //AND U335bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U335bar (
    .O(n633bar),
    .I0(inbar[239]),
    .I1(inbar[218])
  );
  //OR U336
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U336 (
    .O(n634),
    .I0(in_13),
    .I1(in[87])
  );
  //AND U336bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U336bar (
    .O(n634bar),
    .I0(in_13bar),
    .I1(inbar[87])
  );
  //OR U337
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U337 (
    .O(n636),
    .I0(n632),
    .I1(n631)
  );
  //AND U337bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U337bar (
    .O(n636bar),
    .I0(n632bar),
    .I1(n631bar)
  );
  //OR U338
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U338 (
    .O(n631),
    .I0(in_72),
    .I1(in_70)
  );
  //AND U338bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U338bar (
    .O(n631bar),
    .I0(in_72bar),
    .I1(in_70bar)
  );
  //OR U339
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U339 (
    .O(n632),
    .I0(in_80),
    .I1(in_74)
  );
  //AND U339bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U339bar (
    .O(n632bar),
    .I0(in_80bar),
    .I1(in_74bar)
  );
  //OR U340
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U340 (
    .O(n942),
    .I0(n630),
    .I1(n629)
  );
  //AND U340bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U340bar (
    .O(n942bar),
    .I0(n630bar),
    .I1(n629bar)
  );
  //OR U341
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U341 (
    .O(n629),
    .I0(n628),
    .I1(n627)
  );
  //AND U341bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U341bar (
    .O(n629bar),
    .I0(n628bar),
    .I1(n627bar)
  );
  //OR U342
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U342 (
    .O(n627),
    .I0(n626),
    .I1(n625)
  );
  //AND U342bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U342bar (
    .O(n627bar),
    .I0(n626bar),
    .I1(n625bar)
  );
  //OR U343
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U343 (
    .O(n625),
    .I0(in[146]),
    .I1(in[100])
  );
  //AND U343bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U343bar (
    .O(n625bar),
    .I0(inbar[146]),
    .I1(inbar[100])
  );
  //OR U344
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U344 (
    .O(n626),
    .I0(in[168]),
    .I1(in[152])
  );
  //AND U344bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U344bar (
    .O(n626bar),
    .I0(inbar[168]),
    .I1(inbar[152])
  );
  //OR U345
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U345 (
    .O(n628),
    .I0(n624),
    .I1(n623)
  );
  //AND U345bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U345bar (
    .O(n628bar),
    .I0(n624bar),
    .I1(n623bar)
  );
  //OR U346
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U346 (
    .O(n623),
    .I0(in[199]),
    .I1(in[182])
  );
  //AND U346bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U346bar (
    .O(n623bar),
    .I0(inbar[199]),
    .I1(inbar[182])
  );
  //OR U347
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U347 (
    .O(n624),
    .I0(in[236]),
    .I1(in[204])
  );
  //AND U347bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U347bar (
    .O(n624bar),
    .I0(inbar[236]),
    .I1(inbar[204])
  );
  //OR U348
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U348 (
    .O(n630),
    .I0(n622),
    .I1(n621)
  );
  //AND U348bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U348bar (
    .O(n630bar),
    .I0(n622bar),
    .I1(n621bar)
  );
  //OR U349
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U349 (
    .O(n621),
    .I0(n620),
    .I1(n619)
  );
  //AND U349bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U349bar (
    .O(n621bar),
    .I0(n620bar),
    .I1(n619bar)
  );
  //OR U350
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U350 (
    .O(n619),
    .I0(in[89]),
    .I1(in[246])
  );
  //AND U350bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U350bar (
    .O(n619bar),
    .I0(inbar[89]),
    .I1(inbar[246])
  );
  //OR U351
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U351 (
    .O(n620),
    .I0(in[95]),
    .I1(in[92])
  );
  //AND U351bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U351bar (
    .O(n620bar),
    .I0(inbar[95]),
    .I1(inbar[92])
  );
  //OR U352
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U352 (
    .O(n622),
    .I0(n618),
    .I1(n617)
  );
  //AND U352bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U352bar (
    .O(n622bar),
    .I0(n618bar),
    .I1(n617bar)
  );
  //OR U353
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U353 (
    .O(n617),
    .I0(in_22),
    .I1(in_16)
  );
  //AND U353bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U353bar (
    .O(n617bar),
    .I0(in_22bar),
    .I1(in_16bar)
  );
  //OR U354
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U354 (
    .O(n618),
    .I0(in_51),
    .I1(in_49)
  );
  //AND U354bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U354bar (
    .O(n618bar),
    .I0(in_51bar),
    .I1(in_49bar)
  );
  //OR U355
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U355 (
    .O(n722),
    .I0(n616),
    .I1(n615)
  );
  //AND U355bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U355bar (
    .O(n722bar),
    .I0(n616bar),
    .I1(n615bar)
  );
  //OR U356
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U356 (
    .O(n615),
    .I0(in[158]),
    .I1(in[115])
  );
  //AND U356bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U356bar (
    .O(n615bar),
    .I0(inbar[158]),
    .I1(inbar[115])
  );
  //OR U357
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U357 (
    .O(n616),
    .I0(in[163]),
    .I1(n614)
  );
  //AND U357bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U357bar (
    .O(n616bar),
    .I0(inbar[163]),
    .I1(n614bar)
  );
  //OR U358
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U358 (
    .O(n614),
    .I0(in[206]),
    .I1(in[165])
  );
  //AND U358bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U358bar (
    .O(n614bar),
    .I0(inbar[206]),
    .I1(inbar[165])
  );
  //OR U359
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U359 (
    .O(n724),
    .I0(n613),
    .I1(n612)
  );
  //AND U359bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U359bar (
    .O(n724bar),
    .I0(n613bar),
    .I1(n612bar)
  );
  //OR U360
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U360 (
    .O(n612),
    .I0(n611),
    .I1(n610)
  );
  //AND U360bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U360bar (
    .O(n612bar),
    .I0(n611bar),
    .I1(n610bar)
  );
  //OR U361
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U361 (
    .O(n610),
    .I0(in[213]),
    .I1(in[207])
  );
  //AND U361bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U361bar (
    .O(n610bar),
    .I0(inbar[213]),
    .I1(inbar[207])
  );
  //OR U362
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U362 (
    .O(n611),
    .I0(in[215]),
    .I1(n609)
  );
  //AND U362bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U362bar (
    .O(n611bar),
    .I0(inbar[215]),
    .I1(n609bar)
  );
  //OR U363
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U363 (
    .O(n609),
    .I0(in[230]),
    .I1(in[220])
  );
  //AND U363bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U363bar (
    .O(n609bar),
    .I0(inbar[230]),
    .I1(inbar[220])
  );
  //OR U364
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U364 (
    .O(n613),
    .I0(n608),
    .I1(n607)
  );
  //AND U364bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U364bar (
    .O(n613bar),
    .I0(n608bar),
    .I1(n607bar)
  );
  //OR U365
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U365 (
    .O(n607),
    .I0(in[251]),
    .I1(in[234])
  );
  //AND U365bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U365bar (
    .O(n607bar),
    .I0(inbar[251]),
    .I1(inbar[234])
  );
  //OR U366
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U366 (
    .O(n608),
    .I0(in_17),
    .I1(n606)
  );
  //AND U366bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U366bar (
    .O(n608bar),
    .I0(in_17bar),
    .I1(n606bar)
  );
  //OR U367
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U367 (
    .O(n606),
    .I0(in_65),
    .I1(in_56)
  );
  //AND U367bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U367bar (
    .O(n606bar),
    .I0(in_65bar),
    .I1(in_56bar)
  );
  //OR U368
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U368 (
    .O(out[0]),
    .I0(n605),
    .I1(n604)
  );
  //AND U368bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U368bar (
    .O(outbar[0]),
    .I0(n605bar),
    .I1(n604bar)
  );
  //OR U369
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U369 (
    .O(n604),
    .I0(n603),
    .I1(n602)
  );
  //AND U369bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U369bar (
    .O(n604bar),
    .I0(n603bar),
    .I1(n602bar)
  );
  //OR U370
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U370 (
    .O(n602),
    .I0(n601),
    .I1(n600)
  );
  //AND U370bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U370bar (
    .O(n602bar),
    .I0(n601bar),
    .I1(n600bar)
  );
  //OR U371
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U371 (
    .O(n600),
    .I0(n820),
    .I1(n785)
  );
  //AND U371bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U371bar (
    .O(n600bar),
    .I0(n820bar),
    .I1(n785bar)
  );
  //OR U372
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U372 (
    .O(n785),
    .I0(n599),
    .I1(n598)
  );
  //AND U372bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U372bar (
    .O(n785bar),
    .I0(n599bar),
    .I1(n598bar)
  );
  //OR U373
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U373 (
    .O(n598),
    .I0(n597),
    .I1(n596)
  );
  //AND U373bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U373bar (
    .O(n598bar),
    .I0(n597bar),
    .I1(n596bar)
  );
  //OR U374
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U374 (
    .O(n596),
    .I0(n595),
    .I1(n594)
  );
  //AND U374bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U374bar (
    .O(n596bar),
    .I0(n595bar),
    .I1(n594bar)
  );
  //OR U375
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U375 (
    .O(n594),
    .I0(in[135]),
    .I1(in[104])
  );
  //AND U375bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U375bar (
    .O(n594bar),
    .I0(inbar[135]),
    .I1(inbar[104])
  );
  //OR U376
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U376 (
    .O(n595),
    .I0(in[188]),
    .I1(in[178])
  );
  //AND U376bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U376bar (
    .O(n595bar),
    .I0(inbar[188]),
    .I1(inbar[178])
  );
  //OR U377
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U377 (
    .O(n597),
    .I0(n593),
    .I1(n592)
  );
  //AND U377bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U377bar (
    .O(n597bar),
    .I0(n593bar),
    .I1(n592bar)
  );
  //OR U378
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U378 (
    .O(n592),
    .I0(in[217]),
    .I1(in[194])
  );
  //AND U378bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U378bar (
    .O(n592bar),
    .I0(inbar[217]),
    .I1(inbar[194])
  );
  //OR U379
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U379 (
    .O(n593),
    .I0(in[237]),
    .I1(in[218])
  );
  //AND U379bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U379bar (
    .O(n593bar),
    .I0(inbar[237]),
    .I1(inbar[218])
  );
  //OR U380
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U380 (
    .O(n599),
    .I0(n591),
    .I1(n590)
  );
  //AND U380bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U380bar (
    .O(n599bar),
    .I0(n591bar),
    .I1(n590bar)
  );
  //OR U381
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U381 (
    .O(n590),
    .I0(n589),
    .I1(n588)
  );
  //AND U381bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U381bar (
    .O(n590bar),
    .I0(n589bar),
    .I1(n588bar)
  );
  //OR U382
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U382 (
    .O(n588),
    .I0(in_2),
    .I1(in_10)
  );
  //AND U382bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U382bar (
    .O(n588bar),
    .I0(in_2bar),
    .I1(in_10bar)
  );
  //OR U383
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U383 (
    .O(n589),
    .I0(in_47),
    .I1(in_22)
  );
  //AND U383bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U383bar (
    .O(n589bar),
    .I0(in_47bar),
    .I1(in_22bar)
  );
  //OR U384
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U384 (
    .O(n591),
    .I0(n587),
    .I1(n586)
  );
  //AND U384bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U384bar (
    .O(n591bar),
    .I0(n587bar),
    .I1(n586bar)
  );
  //OR U385
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U385 (
    .O(n586),
    .I0(in_56),
    .I1(in_54)
  );
  //AND U385bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U385bar (
    .O(n586bar),
    .I0(in_56bar),
    .I1(in_54bar)
  );
  //OR U386
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U386 (
    .O(n587),
    .I0(in_63),
    .I1(in_61)
  );
  //AND U386bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U386bar (
    .O(n587bar),
    .I0(in_63bar),
    .I1(in_61bar)
  );
  //OR U387
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U387 (
    .O(n820),
    .I0(n585),
    .I1(n584)
  );
  //AND U387bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U387bar (
    .O(n820bar),
    .I0(n585bar),
    .I1(n584bar)
  );
  //OR U388
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U388 (
    .O(n584),
    .I0(n583),
    .I1(n582)
  );
  //AND U388bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U388bar (
    .O(n584bar),
    .I0(n583bar),
    .I1(n582bar)
  );
  //OR U389
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U389 (
    .O(n582),
    .I0(n581),
    .I1(n580)
  );
  //AND U389bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U389bar (
    .O(n582bar),
    .I0(n581bar),
    .I1(n580bar)
  );
  //OR U390
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U390 (
    .O(n580),
    .I0(in[158]),
    .I1(in[142])
  );
  //AND U390bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U390bar (
    .O(n580bar),
    .I0(inbar[158]),
    .I1(inbar[142])
  );
  //OR U391
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U391 (
    .O(n581),
    .I0(in[175]),
    .I1(in[164])
  );
  //AND U391bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U391bar (
    .O(n581bar),
    .I0(inbar[175]),
    .I1(inbar[164])
  );
  //OR U392
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U392 (
    .O(n583),
    .I0(n579),
    .I1(n578)
  );
  //AND U392bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U392bar (
    .O(n583bar),
    .I0(n579bar),
    .I1(n578bar)
  );
  //OR U393
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U393 (
    .O(n578),
    .I0(in[228]),
    .I1(in[204])
  );
  //AND U393bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U393bar (
    .O(n578bar),
    .I0(inbar[228]),
    .I1(inbar[204])
  );
  //OR U394
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U394 (
    .O(n579),
    .I0(in[91]),
    .I1(in[87])
  );
  //AND U394bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U394bar (
    .O(n579bar),
    .I0(inbar[91]),
    .I1(inbar[87])
  );
  //OR U395
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U395 (
    .O(n585),
    .I0(n577),
    .I1(n576)
  );
  //AND U395bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U395bar (
    .O(n585bar),
    .I0(n577bar),
    .I1(n576bar)
  );
  //OR U396
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U396 (
    .O(n576),
    .I0(n575),
    .I1(n574)
  );
  //AND U396bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U396bar (
    .O(n576bar),
    .I0(n575bar),
    .I1(n574bar)
  );
  //OR U397
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U397 (
    .O(n574),
    .I0(in_21),
    .I1(in_11)
  );
  //AND U397bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U397bar (
    .O(n574bar),
    .I0(in_21bar),
    .I1(in_11bar)
  );
  //OR U398
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U398 (
    .O(n575),
    .I0(in_5),
    .I1(in_3)
  );
  //AND U398bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U398bar (
    .O(n575bar),
    .I0(in_5bar),
    .I1(in_3bar)
  );
  //OR U399
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U399 (
    .O(n577),
    .I0(n573),
    .I1(n572)
  );
  //AND U399bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U399bar (
    .O(n577bar),
    .I0(n573bar),
    .I1(n572bar)
  );
  //OR U400
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U400 (
    .O(n572),
    .I0(in_68),
    .I1(in_64)
  );
  //AND U400bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U400bar (
    .O(n572bar),
    .I0(in_68bar),
    .I1(in_64bar)
  );
  //OR U401
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U401 (
    .O(n573),
    .I0(in_76),
    .I1(in_73)
  );
  //AND U401bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U401bar (
    .O(n573bar),
    .I0(in_76bar),
    .I1(in_73bar)
  );
  //OR U402
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U402 (
    .O(n601),
    .I0(n778),
    .I1(n571)
  );
  //AND U402bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U402bar (
    .O(n601bar),
    .I0(n778bar),
    .I1(n571bar)
  );
  //OR U403
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U403 (
    .O(n571),
    .I0(in[100]),
    .I1(n965)
  );
  //AND U403bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U403bar (
    .O(n571bar),
    .I0(inbar[100]),
    .I1(n965bar)
  );
  //OR U404
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U404 (
    .O(n965),
    .I0(n570),
    .I1(n569)
  );
  //AND U404bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U404bar (
    .O(n965bar),
    .I0(n570bar),
    .I1(n569bar)
  );
  //OR U405
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U405 (
    .O(n569),
    .I0(n568),
    .I1(n567)
  );
  //AND U405bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U405bar (
    .O(n569bar),
    .I0(n568bar),
    .I1(n567bar)
  );
  //OR U406
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U406 (
    .O(n567),
    .I0(n566),
    .I1(n565)
  );
  //AND U406bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U406bar (
    .O(n567bar),
    .I0(n566bar),
    .I1(n565bar)
  );
  //OR U407
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U407 (
    .O(n565),
    .I0(n817),
    .I1(n750)
  );
  //AND U407bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U407bar (
    .O(n565bar),
    .I0(n817bar),
    .I1(n750bar)
  );
  //OR U408
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U408 (
    .O(n750),
    .I0(n564),
    .I1(n563)
  );
  //AND U408bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U408bar (
    .O(n750bar),
    .I0(n564bar),
    .I1(n563bar)
  );
  //OR U409
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U409 (
    .O(n563),
    .I0(n562),
    .I1(n561)
  );
  //AND U409bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U409bar (
    .O(n563bar),
    .I0(n562bar),
    .I1(n561bar)
  );
  //OR U410
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U410 (
    .O(n561),
    .I0(n560),
    .I1(n559)
  );
  //AND U410bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U410bar (
    .O(n561bar),
    .I0(n560bar),
    .I1(n559bar)
  );
  //OR U411
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U411 (
    .O(n559),
    .I0(in[119]),
    .I1(in[103])
  );
  //AND U411bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U411bar (
    .O(n559bar),
    .I0(inbar[119]),
    .I1(inbar[103])
  );
  //OR U412
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U412 (
    .O(n560),
    .I0(in[137]),
    .I1(in[133])
  );
  //AND U412bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U412bar (
    .O(n560bar),
    .I0(inbar[137]),
    .I1(inbar[133])
  );
  //OR U413
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U413 (
    .O(n562),
    .I0(n558),
    .I1(n557)
  );
  //AND U413bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U413bar (
    .O(n562bar),
    .I0(n558bar),
    .I1(n557bar)
  );
  //OR U414
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U414 (
    .O(n557),
    .I0(in[176]),
    .I1(in[173])
  );
  //AND U414bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U414bar (
    .O(n557bar),
    .I0(inbar[176]),
    .I1(inbar[173])
  );
  //OR U415
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U415 (
    .O(n558),
    .I0(in[210]),
    .I1(in[181])
  );
  //AND U415bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U415bar (
    .O(n558bar),
    .I0(inbar[210]),
    .I1(inbar[181])
  );
  //OR U416
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U416 (
    .O(n564),
    .I0(n556),
    .I1(n555)
  );
  //AND U416bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U416bar (
    .O(n564bar),
    .I0(n556bar),
    .I1(n555bar)
  );
  //OR U417
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U417 (
    .O(n555),
    .I0(n554),
    .I1(n553)
  );
  //AND U417bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U417bar (
    .O(n555bar),
    .I0(n554bar),
    .I1(n553bar)
  );
  //OR U418
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U418 (
    .O(n553),
    .I0(in_13),
    .I1(in[234])
  );
  //AND U418bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U418bar (
    .O(n553bar),
    .I0(in_13bar),
    .I1(inbar[234])
  );
  //OR U419
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U419 (
    .O(n554),
    .I0(in_38),
    .I1(in_32)
  );
  //AND U419bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U419bar (
    .O(n554bar),
    .I0(in_38bar),
    .I1(in_32bar)
  );
  //OR U420
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U420 (
    .O(n556),
    .I0(n552),
    .I1(n551)
  );
  //AND U420bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U420bar (
    .O(n556bar),
    .I0(n552bar),
    .I1(n551bar)
  );
  //OR U421
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U421 (
    .O(n551),
    .I0(in_42),
    .I1(in_41)
  );
  //AND U421bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U421bar (
    .O(n551bar),
    .I0(in_42bar),
    .I1(in_41bar)
  );
  //OR U422
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U422 (
    .O(n552),
    .I0(in_7),
    .I1(in_49)
  );
  //AND U422bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U422bar (
    .O(n552bar),
    .I0(in_7bar),
    .I1(in_49bar)
  );
  //OR U423
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U423 (
    .O(n817),
    .I0(n550),
    .I1(n549)
  );
  //AND U423bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U423bar (
    .O(n817bar),
    .I0(n550bar),
    .I1(n549bar)
  );
  //OR U424
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U424 (
    .O(n549),
    .I0(n548),
    .I1(n547)
  );
  //AND U424bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U424bar (
    .O(n549bar),
    .I0(n548bar),
    .I1(n547bar)
  );
  //OR U425
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U425 (
    .O(n547),
    .I0(n546),
    .I1(n545)
  );
  //AND U425bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U425bar (
    .O(n547bar),
    .I0(n546bar),
    .I1(n545bar)
  );
  //OR U426
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U426 (
    .O(n545),
    .I0(in[159]),
    .I1(in[105])
  );
  //AND U426bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U426bar (
    .O(n545bar),
    .I0(inbar[159]),
    .I1(inbar[105])
  );
  //OR U427
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U427 (
    .O(n546),
    .I0(in[206]),
    .I1(in[183])
  );
  //AND U427bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U427bar (
    .O(n546bar),
    .I0(inbar[206]),
    .I1(inbar[183])
  );
  //OR U428
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U428 (
    .O(n548),
    .I0(n544),
    .I1(n543)
  );
  //AND U428bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U428bar (
    .O(n548bar),
    .I0(n544bar),
    .I1(n543bar)
  );
  //OR U429
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U429 (
    .O(n543),
    .I0(in[229]),
    .I1(in[219])
  );
  //AND U429bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U429bar (
    .O(n543bar),
    .I0(inbar[229]),
    .I1(inbar[219])
  );
  //OR U430
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U430 (
    .O(n544),
    .I0(in[235]),
    .I1(in[232])
  );
  //AND U430bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U430bar (
    .O(n544bar),
    .I0(inbar[235]),
    .I1(inbar[232])
  );
  //OR U431
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U431 (
    .O(n550),
    .I0(n542),
    .I1(n541)
  );
  //AND U431bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U431bar (
    .O(n550bar),
    .I0(n542bar),
    .I1(n541bar)
  );
  //OR U432
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U432 (
    .O(n541),
    .I0(n540),
    .I1(n539)
  );
  //AND U432bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U432bar (
    .O(n541bar),
    .I0(n540bar),
    .I1(n539bar)
  );
  //OR U433
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U433 (
    .O(n539),
    .I0(in[249]),
    .I1(in[242])
  );
  //AND U433bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U433bar (
    .O(n539bar),
    .I0(inbar[249]),
    .I1(inbar[242])
  );
  //OR U434
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U434 (
    .O(n540),
    .I0(in[89]),
    .I1(in[254])
  );
  //AND U434bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U434bar (
    .O(n540bar),
    .I0(inbar[89]),
    .I1(inbar[254])
  );
  //OR U435
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U435 (
    .O(n542),
    .I0(n538),
    .I1(n537)
  );
  //AND U435bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U435bar (
    .O(n542bar),
    .I0(n538bar),
    .I1(n537bar)
  );
  //OR U436
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U436 (
    .O(n537),
    .I0(in_14),
    .I1(in[99])
  );
  //AND U436bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U436bar (
    .O(n537bar),
    .I0(in_14bar),
    .I1(inbar[99])
  );
  //OR U437
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U437 (
    .O(n538),
    .I0(in_60),
    .I1(in_18)
  );
  //AND U437bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U437bar (
    .O(n538bar),
    .I0(in_60bar),
    .I1(in_18bar)
  );
  //OR U438
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U438 (
    .O(n566),
    .I0(in[113]),
    .I1(n763)
  );
  //AND U438bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U438bar (
    .O(n566bar),
    .I0(inbar[113]),
    .I1(n763bar)
  );
  //OR U439
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U439 (
    .O(n763),
    .I0(n536),
    .I1(n535)
  );
  //AND U439bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U439bar (
    .O(n763bar),
    .I0(n536bar),
    .I1(n535bar)
  );
  //OR U440
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U440 (
    .O(n535),
    .I0(n534),
    .I1(n533)
  );
  //AND U440bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U440bar (
    .O(n535bar),
    .I0(n534bar),
    .I1(n533bar)
  );
  //OR U441
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U441 (
    .O(n533),
    .I0(n532),
    .I1(n531)
  );
  //AND U441bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U441bar (
    .O(n533bar),
    .I0(n532bar),
    .I1(n531bar)
  );
  //OR U442
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U442 (
    .O(n531),
    .I0(in[115]),
    .I1(in[110])
  );
  //AND U442bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U442bar (
    .O(n531bar),
    .I0(inbar[115]),
    .I1(inbar[110])
  );
  //OR U443
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U443 (
    .O(n532),
    .I0(in[125]),
    .I1(in[117])
  );
  //AND U443bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U443bar (
    .O(n532bar),
    .I0(inbar[125]),
    .I1(inbar[117])
  );
  //OR U444
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U444 (
    .O(n534),
    .I0(n530),
    .I1(n529)
  );
  //AND U444bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U444bar (
    .O(n534bar),
    .I0(n530bar),
    .I1(n529bar)
  );
  //OR U445
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U445 (
    .O(n529),
    .I0(in[180]),
    .I1(in[128])
  );
  //AND U445bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U445bar (
    .O(n529bar),
    .I0(inbar[180]),
    .I1(inbar[128])
  );
  //OR U446
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U446 (
    .O(n530),
    .I0(in[205]),
    .I1(in[201])
  );
  //AND U446bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U446bar (
    .O(n530bar),
    .I0(inbar[205]),
    .I1(inbar[201])
  );
  //OR U447
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U447 (
    .O(n536),
    .I0(n528),
    .I1(n527)
  );
  //AND U447bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U447bar (
    .O(n536bar),
    .I0(n528bar),
    .I1(n527bar)
  );
  //OR U448
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U448 (
    .O(n527),
    .I0(n526),
    .I1(n525)
  );
  //AND U448bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U448bar (
    .O(n527bar),
    .I0(n526bar),
    .I1(n525bar)
  );
  //OR U449
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U449 (
    .O(n525),
    .I0(in[244]),
    .I1(in[239])
  );
  //AND U449bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U449bar (
    .O(n525bar),
    .I0(inbar[244]),
    .I1(inbar[239])
  );
  //OR U450
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U450 (
    .O(n526),
    .I0(in[95]),
    .I1(in[83])
  );
  //AND U450bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U450bar (
    .O(n526bar),
    .I0(inbar[95]),
    .I1(inbar[83])
  );
  //OR U451
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U451 (
    .O(n528),
    .I0(n524),
    .I1(n523)
  );
  //AND U451bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U451bar (
    .O(n528bar),
    .I0(n524bar),
    .I1(n523bar)
  );
  //OR U452
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U452 (
    .O(n523),
    .I0(in_24),
    .I1(in[97])
  );
  //AND U452bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U452bar (
    .O(n523bar),
    .I0(in_24bar),
    .I1(inbar[97])
  );
  //OR U453
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U453 (
    .O(n524),
    .I0(in_33),
    .I1(in_27)
  );
  //AND U453bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U453bar (
    .O(n524bar),
    .I0(in_33bar),
    .I1(in_27bar)
  );
  //OR U454
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U454 (
    .O(n568),
    .I0(n522),
    .I1(n521)
  );
  //AND U454bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U454bar (
    .O(n568bar),
    .I0(n522bar),
    .I1(n521bar)
  );
  //OR U455
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U455 (
    .O(n521),
    .I0(in[145]),
    .I1(in[126])
  );
  //AND U455bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U455bar (
    .O(n521bar),
    .I0(inbar[145]),
    .I1(inbar[126])
  );
  //OR U456
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U456 (
    .O(n522),
    .I0(in[169]),
    .I1(n520)
  );
  //AND U456bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U456bar (
    .O(n522bar),
    .I0(inbar[169]),
    .I1(n520bar)
  );
  //OR U457
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U457 (
    .O(n520),
    .I0(in[221]),
    .I1(in[172])
  );
  //AND U457bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U457bar (
    .O(n520bar),
    .I0(inbar[221]),
    .I1(inbar[172])
  );
  //OR U458
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U458 (
    .O(n570),
    .I0(n519),
    .I1(n518)
  );
  //AND U458bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U458bar (
    .O(n570bar),
    .I0(n519bar),
    .I1(n518bar)
  );
  //OR U459
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U459 (
    .O(n518),
    .I0(n517),
    .I1(n516)
  );
  //AND U459bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U459bar (
    .O(n518bar),
    .I0(n517bar),
    .I1(n516bar)
  );
  //OR U460
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U460 (
    .O(n516),
    .I0(in[241]),
    .I1(in[224])
  );
  //AND U460bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U460bar (
    .O(n516bar),
    .I0(inbar[241]),
    .I1(inbar[224])
  );
  //OR U461
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U461 (
    .O(n517),
    .I0(in[86]),
    .I1(n515)
  );
  //AND U461bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U461bar (
    .O(n517bar),
    .I0(inbar[86]),
    .I1(n515bar)
  );
  //OR U462
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U462 (
    .O(n515),
    .I0(in_43),
    .I1(in_34)
  );
  //AND U462bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U462bar (
    .O(n515bar),
    .I0(in_43bar),
    .I1(in_34bar)
  );
  //OR U463
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U463 (
    .O(n519),
    .I0(n514),
    .I1(n513)
  );
  //AND U463bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U463bar (
    .O(n519bar),
    .I0(n514bar),
    .I1(n513bar)
  );
  //OR U464
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U464 (
    .O(n513),
    .I0(in_65),
    .I1(in_51)
  );
  //AND U464bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U464bar (
    .O(n513bar),
    .I0(in_65bar),
    .I1(in_51bar)
  );
  //OR U465
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U465 (
    .O(n514),
    .I0(in_75),
    .I1(n512)
  );
  //AND U465bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U465bar (
    .O(n514bar),
    .I0(in_75bar),
    .I1(n512bar)
  );
  //OR U466
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U466 (
    .O(n512),
    .I0(in_81),
    .I1(in_77)
  );
  //AND U466bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U466bar (
    .O(n512bar),
    .I0(in_81bar),
    .I1(in_77bar)
  );
  //OR U467
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U467 (
    .O(n778),
    .I0(n511),
    .I1(n510)
  );
  //AND U467bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U467bar (
    .O(n778bar),
    .I0(n511bar),
    .I1(n510bar)
  );
  //OR U468
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U468 (
    .O(n510),
    .I0(n509),
    .I1(n508)
  );
  //AND U468bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U468bar (
    .O(n510bar),
    .I0(n509bar),
    .I1(n508bar)
  );
  //OR U469
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U469 (
    .O(n508),
    .I0(n507),
    .I1(n506)
  );
  //AND U469bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U469bar (
    .O(n508bar),
    .I0(n507bar),
    .I1(n506bar)
  );
  //OR U470
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U470 (
    .O(n506),
    .I0(in[107]),
    .I1(in[101])
  );
  //AND U470bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U470bar (
    .O(n506bar),
    .I0(inbar[107]),
    .I1(inbar[101])
  );
  //OR U471
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U471 (
    .O(n507),
    .I0(in[139]),
    .I1(in[132])
  );
  //AND U471bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U471bar (
    .O(n507bar),
    .I0(inbar[139]),
    .I1(inbar[132])
  );
  //OR U472
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U472 (
    .O(n509),
    .I0(n505),
    .I1(n504)
  );
  //AND U472bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U472bar (
    .O(n509bar),
    .I0(n505bar),
    .I1(n504bar)
  );
  //OR U473
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U473 (
    .O(n504),
    .I0(in[146]),
    .I1(in[141])
  );
  //AND U473bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U473bar (
    .O(n504bar),
    .I0(inbar[146]),
    .I1(inbar[141])
  );
  //OR U474
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U474 (
    .O(n505),
    .I0(in[203]),
    .I1(in[179])
  );
  //AND U474bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U474bar (
    .O(n505bar),
    .I0(inbar[203]),
    .I1(inbar[179])
  );
  //OR U475
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U475 (
    .O(n511),
    .I0(n503),
    .I1(n502)
  );
  //AND U475bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U475bar (
    .O(n511bar),
    .I0(n503bar),
    .I1(n502bar)
  );
  //OR U476
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U476 (
    .O(n502),
    .I0(n501),
    .I1(n500)
  );
  //AND U476bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U476bar (
    .O(n502bar),
    .I0(n501bar),
    .I1(n500bar)
  );
  //OR U477
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U477 (
    .O(n500),
    .I0(in[243]),
    .I1(in[222])
  );
  //AND U477bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U477bar (
    .O(n500bar),
    .I0(inbar[243]),
    .I1(inbar[222])
  );
  //OR U478
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U478 (
    .O(n501),
    .I0(in[251]),
    .I1(in[250])
  );
  //AND U478bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U478bar (
    .O(n501bar),
    .I0(inbar[251]),
    .I1(inbar[250])
  );
  //OR U479
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U479 (
    .O(n503),
    .I0(n499),
    .I1(n498)
  );
  //AND U479bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U479bar (
    .O(n503bar),
    .I0(n499bar),
    .I1(n498bar)
  );
  //OR U480
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U480 (
    .O(n498),
    .I0(in_37),
    .I1(in_19)
  );
  //AND U480bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U480bar (
    .O(n498bar),
    .I0(in_37bar),
    .I1(in_19bar)
  );
  //OR U481
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U481 (
    .O(n499),
    .I0(in_78),
    .I1(in_6)
  );
  //AND U481bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U481bar (
    .O(n499bar),
    .I0(in_78bar),
    .I1(in_6bar)
  );
  //OR U482
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U482 (
    .O(n603),
    .I0(n497),
    .I1(n496)
  );
  //AND U482bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U482bar (
    .O(n603bar),
    .I0(n497bar),
    .I1(n496bar)
  );
  //OR U483
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U483 (
    .O(n496),
    .I0(in[112]),
    .I1(in[102])
  );
  //AND U483bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U483bar (
    .O(n496bar),
    .I0(inbar[112]),
    .I1(inbar[102])
  );
  //OR U484
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U484 (
    .O(n497),
    .I0(in[123]),
    .I1(n495)
  );
  //AND U484bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U484bar (
    .O(n497bar),
    .I0(inbar[123]),
    .I1(n495bar)
  );
  //OR U485
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U485 (
    .O(n495),
    .I0(in[143]),
    .I1(in[130])
  );
  //AND U485bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U485bar (
    .O(n495bar),
    .I0(inbar[143]),
    .I1(inbar[130])
  );
  //OR U486
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U486 (
    .O(n605),
    .I0(n494),
    .I1(n493)
  );
  //AND U486bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U486bar (
    .O(n605bar),
    .I0(n494bar),
    .I1(n493bar)
  );
  //OR U487
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U487 (
    .O(n493),
    .I0(n492),
    .I1(n491)
  );
  //AND U487bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U487bar (
    .O(n493bar),
    .I0(n492bar),
    .I1(n491bar)
  );
  //OR U488
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U488 (
    .O(n491),
    .I0(in[216]),
    .I1(in[213])
  );
  //AND U488bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U488bar (
    .O(n491bar),
    .I0(inbar[216]),
    .I1(inbar[213])
  );
  //OR U489
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U489 (
    .O(n492),
    .I0(in[227]),
    .I1(n490)
  );
  //AND U489bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U489bar (
    .O(n492bar),
    .I0(inbar[227]),
    .I1(n490bar)
  );
  //OR U490
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U490 (
    .O(n490),
    .I0(in_0),
    .I1(in[248])
  );
  //AND U490bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U490bar (
    .O(n490bar),
    .I0(in_0bar),
    .I1(inbar[248])
  );
  //OR U491
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U491 (
    .O(n494),
    .I0(n489),
    .I1(n488)
  );
  //AND U491bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U491bar (
    .O(n494bar),
    .I0(n489bar),
    .I1(n488bar)
  );
  //OR U492
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U492 (
    .O(n488),
    .I0(in_46),
    .I1(in_44)
  );
  //AND U492bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U492bar (
    .O(n488bar),
    .I0(in_46bar),
    .I1(in_44bar)
  );
  //OR U493
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U493 (
    .O(n489),
    .I0(in_50),
    .I1(n487)
  );
  //AND U493bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U493bar (
    .O(n489bar),
    .I0(in_50bar),
    .I1(n487bar)
  );
  //OR U494
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U494 (
    .O(n487),
    .I0(in_9),
    .I1(in_80)
  );
  //AND U494bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U494bar (
    .O(n487bar),
    .I0(in_9bar),
    .I1(in_80bar)
  );
endmodule

module sBox_11 ( in, out );

  input wire [7:0] in;
//input_done

  output wire [7:0] out;
//output_done

  wire [255:0] decodeOut;
//wire_done

  decode_11 dec ( .in(in), .out(decodeOut) );
  encode_11 enc ( .in(decodeOut), .out(out) );
endmodule

module CD2_45 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD2_46 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD2_47 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD2_48 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD4_23 ( a, b, y );

  input wire [3:0] a;
  input wire [3:0] b;
  wire [3:0] abar;
  wire [3:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
//input_done

  output wire [15:0] y;
  wire [15:0] ybar;
//output_done

//wire_done

  //AND U1
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1 (
    .O(y[9]),
    .I0(b[1]),
    .I1(a[2])
  );
  //OR U1bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1bar (
    .O(ybar[9]),
    .I0(bbar[1]),
    .I1(abar[2])
  );
  //AND U2
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2 (
    .O(y[8]),
    .I0(b[0]),
    .I1(a[2])
  );
  //OR U2bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2bar (
    .O(ybar[8]),
    .I0(bbar[0]),
    .I1(abar[2])
  );
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[7]),
    .I0(b[3]),
    .I1(a[1])
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[7]),
    .I0(bbar[3]),
    .I1(abar[1])
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[6]),
    .I0(b[2]),
    .I1(a[1])
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[6]),
    .I0(bbar[2]),
    .I1(abar[1])
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[5]),
    .I0(a[1]),
    .I1(b[1])
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[5]),
    .I0(abar[1]),
    .I1(bbar[1])
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[4]),
    .I0(a[1]),
    .I1(b[0])
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[4]),
    .I0(abar[1]),
    .I1(bbar[0])
  );
  //AND U7
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7 (
    .O(y[3]),
    .I0(a[0]),
    .I1(b[3])
  );
  //OR U7bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7bar (
    .O(ybar[3]),
    .I0(abar[0]),
    .I1(bbar[3])
  );
  //AND U8
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8 (
    .O(y[2]),
    .I0(a[0]),
    .I1(b[2])
  );
  //OR U8bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8bar (
    .O(ybar[2]),
    .I0(abar[0]),
    .I1(bbar[2])
  );
  //AND U9
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9 (
    .O(y[1]),
    .I0(a[0]),
    .I1(b[1])
  );
  //OR U9bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9bar (
    .O(ybar[1]),
    .I0(abar[0]),
    .I1(bbar[1])
  );
  //AND U10
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10 (
    .O(y[15]),
    .I0(a[3]),
    .I1(b[3])
  );
  //OR U10bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10bar (
    .O(ybar[15]),
    .I0(abar[3]),
    .I1(bbar[3])
  );
  //AND U11
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11 (
    .O(y[14]),
    .I0(a[3]),
    .I1(b[2])
  );
  //OR U11bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11bar (
    .O(ybar[14]),
    .I0(abar[3]),
    .I1(bbar[2])
  );
  //AND U12
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12 (
    .O(y[13]),
    .I0(a[3]),
    .I1(b[1])
  );
  //OR U12bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12bar (
    .O(ybar[13]),
    .I0(abar[3]),
    .I1(bbar[1])
  );
  //AND U13
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13 (
    .O(y[12]),
    .I0(a[3]),
    .I1(b[0])
  );
  //OR U13bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13bar (
    .O(ybar[12]),
    .I0(abar[3]),
    .I1(bbar[0])
  );
  //AND U14
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14 (
    .O(y[11]),
    .I0(b[3]),
    .I1(a[2])
  );
  //OR U14bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14bar (
    .O(ybar[11]),
    .I0(bbar[3]),
    .I1(abar[2])
  );
  //AND U15
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15 (
    .O(y[10]),
    .I0(b[2]),
    .I1(a[2])
  );
  //OR U15bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15bar (
    .O(ybar[10]),
    .I0(bbar[2]),
    .I1(abar[2])
  );
  //AND U16
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16 (
    .O(y[0]),
    .I0(a[0]),
    .I1(b[0])
  );
  //OR U16bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16bar (
    .O(ybar[0]),
    .I0(abar[0]),
    .I1(bbar[0])
  );
endmodule

module CD4_24 ( a, b, y );

  input wire [3:0] a;
  input wire [3:0] b;
  wire [3:0] abar;
  wire [3:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
//input_done

  output wire [15:0] y;
  wire [15:0] ybar;
//output_done

//wire_done

  //AND U1
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1 (
    .O(y[9]),
    .I0(b[1]),
    .I1(a[2])
  );
  //OR U1bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1bar (
    .O(ybar[9]),
    .I0(bbar[1]),
    .I1(abar[2])
  );
  //AND U2
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2 (
    .O(y[8]),
    .I0(b[0]),
    .I1(a[2])
  );
  //OR U2bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2bar (
    .O(ybar[8]),
    .I0(bbar[0]),
    .I1(abar[2])
  );
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[7]),
    .I0(b[3]),
    .I1(a[1])
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[7]),
    .I0(bbar[3]),
    .I1(abar[1])
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[6]),
    .I0(b[2]),
    .I1(a[1])
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[6]),
    .I0(bbar[2]),
    .I1(abar[1])
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[5]),
    .I0(a[1]),
    .I1(b[1])
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[5]),
    .I0(abar[1]),
    .I1(bbar[1])
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[4]),
    .I0(a[1]),
    .I1(b[0])
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[4]),
    .I0(abar[1]),
    .I1(bbar[0])
  );
  //AND U7
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7 (
    .O(y[3]),
    .I0(a[0]),
    .I1(b[3])
  );
  //OR U7bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7bar (
    .O(ybar[3]),
    .I0(abar[0]),
    .I1(bbar[3])
  );
  //AND U8
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8 (
    .O(y[2]),
    .I0(a[0]),
    .I1(b[2])
  );
  //OR U8bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8bar (
    .O(ybar[2]),
    .I0(abar[0]),
    .I1(bbar[2])
  );
  //AND U9
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9 (
    .O(y[1]),
    .I0(a[0]),
    .I1(b[1])
  );
  //OR U9bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9bar (
    .O(ybar[1]),
    .I0(abar[0]),
    .I1(bbar[1])
  );
  //AND U10
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10 (
    .O(y[15]),
    .I0(a[3]),
    .I1(b[3])
  );
  //OR U10bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10bar (
    .O(ybar[15]),
    .I0(abar[3]),
    .I1(bbar[3])
  );
  //AND U11
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11 (
    .O(y[14]),
    .I0(a[3]),
    .I1(b[2])
  );
  //OR U11bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11bar (
    .O(ybar[14]),
    .I0(abar[3]),
    .I1(bbar[2])
  );
  //AND U12
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12 (
    .O(y[13]),
    .I0(a[3]),
    .I1(b[1])
  );
  //OR U12bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12bar (
    .O(ybar[13]),
    .I0(abar[3]),
    .I1(bbar[1])
  );
  //AND U13
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13 (
    .O(y[12]),
    .I0(a[3]),
    .I1(b[0])
  );
  //OR U13bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13bar (
    .O(ybar[12]),
    .I0(abar[3]),
    .I1(bbar[0])
  );
  //AND U14
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14 (
    .O(y[11]),
    .I0(b[3]),
    .I1(a[2])
  );
  //OR U14bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14bar (
    .O(ybar[11]),
    .I0(bbar[3]),
    .I1(abar[2])
  );
  //AND U15
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15 (
    .O(y[10]),
    .I0(b[2]),
    .I1(a[2])
  );
  //OR U15bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15bar (
    .O(ybar[10]),
    .I0(bbar[2]),
    .I1(abar[2])
  );
  //AND U16
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16 (
    .O(y[0]),
    .I0(a[0]),
    .I1(b[0])
  );
  //OR U16bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16bar (
    .O(ybar[0]),
    .I0(abar[0]),
    .I1(bbar[0])
  );
endmodule

module CD16_12 ( a, b, y );

  input wire [15:0] a;
  input wire [15:0] b;
  wire [15:0] abar;
  wire [15:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign abar[8] = ~a[8];
  assign abar[9] = ~a[9];
  assign abar[10] = ~a[10];
  assign abar[11] = ~a[11];
  assign abar[12] = ~a[12];
  assign abar[13] = ~a[13];
  assign abar[14] = ~a[14];
  assign abar[15] = ~a[15];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign bbar[8] = ~b[8];
  assign bbar[9] = ~b[9];
  assign bbar[10] = ~b[10];
  assign bbar[11] = ~b[11];
  assign bbar[12] = ~b[12];
  assign bbar[13] = ~b[13];
  assign bbar[14] = ~b[14];
  assign bbar[15] = ~b[15];
//input_done

  output wire [255:0] y;
  wire [255:0] ybar;
//output_done

//wire_done

  //AND U1
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1 (
    .O(y[9]),
    .I0(b[9]),
    .I1(a[0])
  );
  //OR U1bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1bar (
    .O(ybar[9]),
    .I0(bbar[9]),
    .I1(abar[0])
  );
  //AND U2
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2 (
    .O(y[99]),
    .I0(b[3]),
    .I1(a[6])
  );
  //OR U2bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2bar (
    .O(ybar[99]),
    .I0(bbar[3]),
    .I1(abar[6])
  );
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[98]),
    .I0(b[2]),
    .I1(a[6])
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[98]),
    .I0(bbar[2]),
    .I1(abar[6])
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[97]),
    .I0(b[1]),
    .I1(a[6])
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[97]),
    .I0(bbar[1]),
    .I1(abar[6])
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[96]),
    .I0(b[0]),
    .I1(a[6])
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[96]),
    .I0(bbar[0]),
    .I1(abar[6])
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[95]),
    .I0(b[15]),
    .I1(a[5])
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[95]),
    .I0(bbar[15]),
    .I1(abar[5])
  );
  //AND U7
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7 (
    .O(y[94]),
    .I0(b[14]),
    .I1(a[5])
  );
  //OR U7bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7bar (
    .O(ybar[94]),
    .I0(bbar[14]),
    .I1(abar[5])
  );
  //AND U8
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8 (
    .O(y[93]),
    .I0(b[13]),
    .I1(a[5])
  );
  //OR U8bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8bar (
    .O(ybar[93]),
    .I0(bbar[13]),
    .I1(abar[5])
  );
  //AND U9
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9 (
    .O(y[92]),
    .I0(b[12]),
    .I1(a[5])
  );
  //OR U9bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9bar (
    .O(ybar[92]),
    .I0(bbar[12]),
    .I1(abar[5])
  );
  //AND U10
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10 (
    .O(y[91]),
    .I0(b[11]),
    .I1(a[5])
  );
  //OR U10bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10bar (
    .O(ybar[91]),
    .I0(bbar[11]),
    .I1(abar[5])
  );
  //AND U11
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11 (
    .O(y[90]),
    .I0(b[10]),
    .I1(a[5])
  );
  //OR U11bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11bar (
    .O(ybar[90]),
    .I0(bbar[10]),
    .I1(abar[5])
  );
  //AND U12
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12 (
    .O(y[8]),
    .I0(b[8]),
    .I1(a[0])
  );
  //OR U12bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12bar (
    .O(ybar[8]),
    .I0(bbar[8]),
    .I1(abar[0])
  );
  //AND U13
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13 (
    .O(y[89]),
    .I0(a[5]),
    .I1(b[9])
  );
  //OR U13bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13bar (
    .O(ybar[89]),
    .I0(abar[5]),
    .I1(bbar[9])
  );
  //AND U14
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14 (
    .O(y[88]),
    .I0(b[8]),
    .I1(a[5])
  );
  //OR U14bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14bar (
    .O(ybar[88]),
    .I0(bbar[8]),
    .I1(abar[5])
  );
  //AND U15
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15 (
    .O(y[87]),
    .I0(b[7]),
    .I1(a[5])
  );
  //OR U15bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15bar (
    .O(ybar[87]),
    .I0(bbar[7]),
    .I1(abar[5])
  );
  //AND U16
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16 (
    .O(y[86]),
    .I0(b[6]),
    .I1(a[5])
  );
  //OR U16bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16bar (
    .O(ybar[86]),
    .I0(bbar[6]),
    .I1(abar[5])
  );
  //AND U17
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U17 (
    .O(y[85]),
    .I0(b[5]),
    .I1(a[5])
  );
  //OR U17bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U17bar (
    .O(ybar[85]),
    .I0(bbar[5]),
    .I1(abar[5])
  );
  //AND U18
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U18 (
    .O(y[84]),
    .I0(b[4]),
    .I1(a[5])
  );
  //OR U18bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U18bar (
    .O(ybar[84]),
    .I0(bbar[4]),
    .I1(abar[5])
  );
  //AND U19
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U19 (
    .O(y[83]),
    .I0(a[5]),
    .I1(b[3])
  );
  //OR U19bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U19bar (
    .O(ybar[83]),
    .I0(abar[5]),
    .I1(bbar[3])
  );
  //AND U20
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U20 (
    .O(y[82]),
    .I0(a[5]),
    .I1(b[2])
  );
  //OR U20bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U20bar (
    .O(ybar[82]),
    .I0(abar[5]),
    .I1(bbar[2])
  );
  //AND U21
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U21 (
    .O(y[81]),
    .I0(a[5]),
    .I1(b[1])
  );
  //OR U21bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U21bar (
    .O(ybar[81]),
    .I0(abar[5]),
    .I1(bbar[1])
  );
  //AND U22
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U22 (
    .O(y[80]),
    .I0(a[5]),
    .I1(b[0])
  );
  //OR U22bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U22bar (
    .O(ybar[80]),
    .I0(abar[5]),
    .I1(bbar[0])
  );
  //AND U23
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U23 (
    .O(y[7]),
    .I0(b[7]),
    .I1(a[0])
  );
  //OR U23bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U23bar (
    .O(ybar[7]),
    .I0(bbar[7]),
    .I1(abar[0])
  );
  //AND U24
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U24 (
    .O(y[79]),
    .I0(a[4]),
    .I1(b[15])
  );
  //OR U24bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U24bar (
    .O(ybar[79]),
    .I0(abar[4]),
    .I1(bbar[15])
  );
  //AND U25
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U25 (
    .O(y[78]),
    .I0(a[4]),
    .I1(b[14])
  );
  //OR U25bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U25bar (
    .O(ybar[78]),
    .I0(abar[4]),
    .I1(bbar[14])
  );
  //AND U26
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U26 (
    .O(y[77]),
    .I0(a[4]),
    .I1(b[13])
  );
  //OR U26bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U26bar (
    .O(ybar[77]),
    .I0(abar[4]),
    .I1(bbar[13])
  );
  //AND U27
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U27 (
    .O(y[76]),
    .I0(a[4]),
    .I1(b[12])
  );
  //OR U27bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U27bar (
    .O(ybar[76]),
    .I0(abar[4]),
    .I1(bbar[12])
  );
  //AND U28
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U28 (
    .O(y[75]),
    .I0(a[4]),
    .I1(b[11])
  );
  //OR U28bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U28bar (
    .O(ybar[75]),
    .I0(abar[4]),
    .I1(bbar[11])
  );
  //AND U29
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U29 (
    .O(y[74]),
    .I0(a[4]),
    .I1(b[10])
  );
  //OR U29bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U29bar (
    .O(ybar[74]),
    .I0(abar[4]),
    .I1(bbar[10])
  );
  //AND U30
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U30 (
    .O(y[73]),
    .I0(a[4]),
    .I1(b[9])
  );
  //OR U30bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U30bar (
    .O(ybar[73]),
    .I0(abar[4]),
    .I1(bbar[9])
  );
  //AND U31
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U31 (
    .O(y[72]),
    .I0(a[4]),
    .I1(b[8])
  );
  //OR U31bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U31bar (
    .O(ybar[72]),
    .I0(abar[4]),
    .I1(bbar[8])
  );
  //AND U32
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U32 (
    .O(y[71]),
    .I0(a[4]),
    .I1(b[7])
  );
  //OR U32bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U32bar (
    .O(ybar[71]),
    .I0(abar[4]),
    .I1(bbar[7])
  );
  //AND U33
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U33 (
    .O(y[70]),
    .I0(a[4]),
    .I1(b[6])
  );
  //OR U33bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U33bar (
    .O(ybar[70]),
    .I0(abar[4]),
    .I1(bbar[6])
  );
  //AND U34
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U34 (
    .O(y[6]),
    .I0(b[6]),
    .I1(a[0])
  );
  //OR U34bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U34bar (
    .O(ybar[6]),
    .I0(bbar[6]),
    .I1(abar[0])
  );
  //AND U35
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U35 (
    .O(y[69]),
    .I0(a[4]),
    .I1(b[5])
  );
  //OR U35bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U35bar (
    .O(ybar[69]),
    .I0(abar[4]),
    .I1(bbar[5])
  );
  //AND U36
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U36 (
    .O(y[68]),
    .I0(a[4]),
    .I1(b[4])
  );
  //OR U36bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U36bar (
    .O(ybar[68]),
    .I0(abar[4]),
    .I1(bbar[4])
  );
  //AND U37
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U37 (
    .O(y[67]),
    .I0(a[4]),
    .I1(b[3])
  );
  //OR U37bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U37bar (
    .O(ybar[67]),
    .I0(abar[4]),
    .I1(bbar[3])
  );
  //AND U38
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U38 (
    .O(y[66]),
    .I0(a[4]),
    .I1(b[2])
  );
  //OR U38bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U38bar (
    .O(ybar[66]),
    .I0(abar[4]),
    .I1(bbar[2])
  );
  //AND U39
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U39 (
    .O(y[65]),
    .I0(a[4]),
    .I1(b[1])
  );
  //OR U39bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U39bar (
    .O(ybar[65]),
    .I0(abar[4]),
    .I1(bbar[1])
  );
  //AND U40
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U40 (
    .O(y[64]),
    .I0(a[4]),
    .I1(b[0])
  );
  //OR U40bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U40bar (
    .O(ybar[64]),
    .I0(abar[4]),
    .I1(bbar[0])
  );
  //AND U41
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U41 (
    .O(y[63]),
    .I0(a[3]),
    .I1(b[15])
  );
  //OR U41bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U41bar (
    .O(ybar[63]),
    .I0(abar[3]),
    .I1(bbar[15])
  );
  //AND U42
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U42 (
    .O(y[62]),
    .I0(a[3]),
    .I1(b[14])
  );
  //OR U42bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U42bar (
    .O(ybar[62]),
    .I0(abar[3]),
    .I1(bbar[14])
  );
  //AND U43
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U43 (
    .O(y[61]),
    .I0(a[3]),
    .I1(b[13])
  );
  //OR U43bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U43bar (
    .O(ybar[61]),
    .I0(abar[3]),
    .I1(bbar[13])
  );
  //AND U44
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U44 (
    .O(y[60]),
    .I0(a[3]),
    .I1(b[12])
  );
  //OR U44bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U44bar (
    .O(ybar[60]),
    .I0(abar[3]),
    .I1(bbar[12])
  );
  //AND U45
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U45 (
    .O(y[5]),
    .I0(b[5]),
    .I1(a[0])
  );
  //OR U45bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U45bar (
    .O(ybar[5]),
    .I0(bbar[5]),
    .I1(abar[0])
  );
  //AND U46
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U46 (
    .O(y[59]),
    .I0(a[3]),
    .I1(b[11])
  );
  //OR U46bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U46bar (
    .O(ybar[59]),
    .I0(abar[3]),
    .I1(bbar[11])
  );
  //AND U47
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U47 (
    .O(y[58]),
    .I0(a[3]),
    .I1(b[10])
  );
  //OR U47bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U47bar (
    .O(ybar[58]),
    .I0(abar[3]),
    .I1(bbar[10])
  );
  //AND U48
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U48 (
    .O(y[57]),
    .I0(a[3]),
    .I1(b[9])
  );
  //OR U48bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U48bar (
    .O(ybar[57]),
    .I0(abar[3]),
    .I1(bbar[9])
  );
  //AND U49
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U49 (
    .O(y[56]),
    .I0(a[3]),
    .I1(b[8])
  );
  //OR U49bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U49bar (
    .O(ybar[56]),
    .I0(abar[3]),
    .I1(bbar[8])
  );
  //AND U50
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U50 (
    .O(y[55]),
    .I0(a[3]),
    .I1(b[7])
  );
  //OR U50bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U50bar (
    .O(ybar[55]),
    .I0(abar[3]),
    .I1(bbar[7])
  );
  //AND U51
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U51 (
    .O(y[54]),
    .I0(a[3]),
    .I1(b[6])
  );
  //OR U51bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U51bar (
    .O(ybar[54]),
    .I0(abar[3]),
    .I1(bbar[6])
  );
  //AND U52
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U52 (
    .O(y[53]),
    .I0(a[3]),
    .I1(b[5])
  );
  //OR U52bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U52bar (
    .O(ybar[53]),
    .I0(abar[3]),
    .I1(bbar[5])
  );
  //AND U53
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U53 (
    .O(y[52]),
    .I0(a[3]),
    .I1(b[4])
  );
  //OR U53bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U53bar (
    .O(ybar[52]),
    .I0(abar[3]),
    .I1(bbar[4])
  );
  //AND U54
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U54 (
    .O(y[51]),
    .I0(a[3]),
    .I1(b[3])
  );
  //OR U54bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U54bar (
    .O(ybar[51]),
    .I0(abar[3]),
    .I1(bbar[3])
  );
  //AND U55
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U55 (
    .O(y[50]),
    .I0(a[3]),
    .I1(b[2])
  );
  //OR U55bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U55bar (
    .O(ybar[50]),
    .I0(abar[3]),
    .I1(bbar[2])
  );
  //AND U56
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U56 (
    .O(y[4]),
    .I0(b[4]),
    .I1(a[0])
  );
  //OR U56bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U56bar (
    .O(ybar[4]),
    .I0(bbar[4]),
    .I1(abar[0])
  );
  //AND U57
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U57 (
    .O(y[49]),
    .I0(a[3]),
    .I1(b[1])
  );
  //OR U57bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U57bar (
    .O(ybar[49]),
    .I0(abar[3]),
    .I1(bbar[1])
  );
  //AND U58
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U58 (
    .O(y[48]),
    .I0(a[3]),
    .I1(b[0])
  );
  //OR U58bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U58bar (
    .O(ybar[48]),
    .I0(abar[3]),
    .I1(bbar[0])
  );
  //AND U59
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U59 (
    .O(y[47]),
    .I0(a[2]),
    .I1(b[15])
  );
  //OR U59bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U59bar (
    .O(ybar[47]),
    .I0(abar[2]),
    .I1(bbar[15])
  );
  //AND U60
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U60 (
    .O(y[46]),
    .I0(a[2]),
    .I1(b[14])
  );
  //OR U60bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U60bar (
    .O(ybar[46]),
    .I0(abar[2]),
    .I1(bbar[14])
  );
  //AND U61
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U61 (
    .O(y[45]),
    .I0(a[2]),
    .I1(b[13])
  );
  //OR U61bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U61bar (
    .O(ybar[45]),
    .I0(abar[2]),
    .I1(bbar[13])
  );
  //AND U62
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U62 (
    .O(y[44]),
    .I0(a[2]),
    .I1(b[12])
  );
  //OR U62bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U62bar (
    .O(ybar[44]),
    .I0(abar[2]),
    .I1(bbar[12])
  );
  //AND U63
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U63 (
    .O(y[43]),
    .I0(a[2]),
    .I1(b[11])
  );
  //OR U63bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U63bar (
    .O(ybar[43]),
    .I0(abar[2]),
    .I1(bbar[11])
  );
  //AND U64
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U64 (
    .O(y[42]),
    .I0(a[2]),
    .I1(b[10])
  );
  //OR U64bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U64bar (
    .O(ybar[42]),
    .I0(abar[2]),
    .I1(bbar[10])
  );
  //AND U65
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U65 (
    .O(y[41]),
    .I0(a[2]),
    .I1(b[9])
  );
  //OR U65bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U65bar (
    .O(ybar[41]),
    .I0(abar[2]),
    .I1(bbar[9])
  );
  //AND U66
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U66 (
    .O(y[40]),
    .I0(a[2]),
    .I1(b[8])
  );
  //OR U66bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U66bar (
    .O(ybar[40]),
    .I0(abar[2]),
    .I1(bbar[8])
  );
  //AND U67
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U67 (
    .O(y[3]),
    .I0(b[3]),
    .I1(a[0])
  );
  //OR U67bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U67bar (
    .O(ybar[3]),
    .I0(bbar[3]),
    .I1(abar[0])
  );
  //AND U68
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U68 (
    .O(y[39]),
    .I0(a[2]),
    .I1(b[7])
  );
  //OR U68bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U68bar (
    .O(ybar[39]),
    .I0(abar[2]),
    .I1(bbar[7])
  );
  //AND U69
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U69 (
    .O(y[38]),
    .I0(a[2]),
    .I1(b[6])
  );
  //OR U69bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U69bar (
    .O(ybar[38]),
    .I0(abar[2]),
    .I1(bbar[6])
  );
  //AND U70
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U70 (
    .O(y[37]),
    .I0(a[2]),
    .I1(b[5])
  );
  //OR U70bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U70bar (
    .O(ybar[37]),
    .I0(abar[2]),
    .I1(bbar[5])
  );
  //AND U71
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U71 (
    .O(y[36]),
    .I0(a[2]),
    .I1(b[4])
  );
  //OR U71bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U71bar (
    .O(ybar[36]),
    .I0(abar[2]),
    .I1(bbar[4])
  );
  //AND U72
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U72 (
    .O(y[35]),
    .I0(a[2]),
    .I1(b[3])
  );
  //OR U72bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U72bar (
    .O(ybar[35]),
    .I0(abar[2]),
    .I1(bbar[3])
  );
  //AND U73
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U73 (
    .O(y[34]),
    .I0(a[2]),
    .I1(b[2])
  );
  //OR U73bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U73bar (
    .O(ybar[34]),
    .I0(abar[2]),
    .I1(bbar[2])
  );
  //AND U74
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U74 (
    .O(y[33]),
    .I0(a[2]),
    .I1(b[1])
  );
  //OR U74bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U74bar (
    .O(ybar[33]),
    .I0(abar[2]),
    .I1(bbar[1])
  );
  //AND U75
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U75 (
    .O(y[32]),
    .I0(a[2]),
    .I1(b[0])
  );
  //OR U75bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U75bar (
    .O(ybar[32]),
    .I0(abar[2]),
    .I1(bbar[0])
  );
  //AND U76
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U76 (
    .O(y[31]),
    .I0(a[1]),
    .I1(b[15])
  );
  //OR U76bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U76bar (
    .O(ybar[31]),
    .I0(abar[1]),
    .I1(bbar[15])
  );
  //AND U77
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U77 (
    .O(y[30]),
    .I0(a[1]),
    .I1(b[14])
  );
  //OR U77bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U77bar (
    .O(ybar[30]),
    .I0(abar[1]),
    .I1(bbar[14])
  );
  //AND U78
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U78 (
    .O(y[2]),
    .I0(b[2]),
    .I1(a[0])
  );
  //OR U78bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U78bar (
    .O(ybar[2]),
    .I0(bbar[2]),
    .I1(abar[0])
  );
  //AND U79
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U79 (
    .O(y[29]),
    .I0(a[1]),
    .I1(b[13])
  );
  //OR U79bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U79bar (
    .O(ybar[29]),
    .I0(abar[1]),
    .I1(bbar[13])
  );
  //AND U80
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U80 (
    .O(y[28]),
    .I0(a[1]),
    .I1(b[12])
  );
  //OR U80bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U80bar (
    .O(ybar[28]),
    .I0(abar[1]),
    .I1(bbar[12])
  );
  //AND U81
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U81 (
    .O(y[27]),
    .I0(a[1]),
    .I1(b[11])
  );
  //OR U81bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U81bar (
    .O(ybar[27]),
    .I0(abar[1]),
    .I1(bbar[11])
  );
  //AND U82
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U82 (
    .O(y[26]),
    .I0(a[1]),
    .I1(b[10])
  );
  //OR U82bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U82bar (
    .O(ybar[26]),
    .I0(abar[1]),
    .I1(bbar[10])
  );
  //AND U83
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U83 (
    .O(y[25]),
    .I0(a[1]),
    .I1(b[9])
  );
  //OR U83bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U83bar (
    .O(ybar[25]),
    .I0(abar[1]),
    .I1(bbar[9])
  );
  //AND U84
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U84 (
    .O(y[255]),
    .I0(a[15]),
    .I1(b[15])
  );
  //OR U84bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U84bar (
    .O(ybar[255]),
    .I0(abar[15]),
    .I1(bbar[15])
  );
  //AND U85
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U85 (
    .O(y[254]),
    .I0(a[15]),
    .I1(b[14])
  );
  //OR U85bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U85bar (
    .O(ybar[254]),
    .I0(abar[15]),
    .I1(bbar[14])
  );
  //AND U86
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U86 (
    .O(y[253]),
    .I0(a[15]),
    .I1(b[13])
  );
  //OR U86bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U86bar (
    .O(ybar[253]),
    .I0(abar[15]),
    .I1(bbar[13])
  );
  //AND U87
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U87 (
    .O(y[252]),
    .I0(a[15]),
    .I1(b[12])
  );
  //OR U87bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U87bar (
    .O(ybar[252]),
    .I0(abar[15]),
    .I1(bbar[12])
  );
  //AND U88
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U88 (
    .O(y[251]),
    .I0(a[15]),
    .I1(b[11])
  );
  //OR U88bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U88bar (
    .O(ybar[251]),
    .I0(abar[15]),
    .I1(bbar[11])
  );
  //AND U89
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U89 (
    .O(y[250]),
    .I0(a[15]),
    .I1(b[10])
  );
  //OR U89bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U89bar (
    .O(ybar[250]),
    .I0(abar[15]),
    .I1(bbar[10])
  );
  //AND U90
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U90 (
    .O(y[24]),
    .I0(a[1]),
    .I1(b[8])
  );
  //OR U90bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U90bar (
    .O(ybar[24]),
    .I0(abar[1]),
    .I1(bbar[8])
  );
  //AND U91
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U91 (
    .O(y[249]),
    .I0(a[15]),
    .I1(b[9])
  );
  //OR U91bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U91bar (
    .O(ybar[249]),
    .I0(abar[15]),
    .I1(bbar[9])
  );
  //AND U92
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U92 (
    .O(y[248]),
    .I0(a[15]),
    .I1(b[8])
  );
  //OR U92bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U92bar (
    .O(ybar[248]),
    .I0(abar[15]),
    .I1(bbar[8])
  );
  //AND U93
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U93 (
    .O(y[247]),
    .I0(a[15]),
    .I1(b[7])
  );
  //OR U93bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U93bar (
    .O(ybar[247]),
    .I0(abar[15]),
    .I1(bbar[7])
  );
  //AND U94
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U94 (
    .O(y[246]),
    .I0(a[15]),
    .I1(b[6])
  );
  //OR U94bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U94bar (
    .O(ybar[246]),
    .I0(abar[15]),
    .I1(bbar[6])
  );
  //AND U95
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U95 (
    .O(y[245]),
    .I0(a[15]),
    .I1(b[5])
  );
  //OR U95bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U95bar (
    .O(ybar[245]),
    .I0(abar[15]),
    .I1(bbar[5])
  );
  //AND U96
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U96 (
    .O(y[244]),
    .I0(a[15]),
    .I1(b[4])
  );
  //OR U96bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U96bar (
    .O(ybar[244]),
    .I0(abar[15]),
    .I1(bbar[4])
  );
  //AND U97
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U97 (
    .O(y[243]),
    .I0(a[15]),
    .I1(b[3])
  );
  //OR U97bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U97bar (
    .O(ybar[243]),
    .I0(abar[15]),
    .I1(bbar[3])
  );
  //AND U98
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U98 (
    .O(y[242]),
    .I0(a[15]),
    .I1(b[2])
  );
  //OR U98bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U98bar (
    .O(ybar[242]),
    .I0(abar[15]),
    .I1(bbar[2])
  );
  //AND U99
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U99 (
    .O(y[241]),
    .I0(a[15]),
    .I1(b[1])
  );
  //OR U99bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U99bar (
    .O(ybar[241]),
    .I0(abar[15]),
    .I1(bbar[1])
  );
  //AND U100
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U100 (
    .O(y[240]),
    .I0(a[15]),
    .I1(b[0])
  );
  //OR U100bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U100bar (
    .O(ybar[240]),
    .I0(abar[15]),
    .I1(bbar[0])
  );
  //AND U101
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U101 (
    .O(y[23]),
    .I0(a[1]),
    .I1(b[7])
  );
  //OR U101bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U101bar (
    .O(ybar[23]),
    .I0(abar[1]),
    .I1(bbar[7])
  );
  //AND U102
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U102 (
    .O(y[239]),
    .I0(a[14]),
    .I1(b[15])
  );
  //OR U102bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U102bar (
    .O(ybar[239]),
    .I0(abar[14]),
    .I1(bbar[15])
  );
  //AND U103
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U103 (
    .O(y[238]),
    .I0(a[14]),
    .I1(b[14])
  );
  //OR U103bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U103bar (
    .O(ybar[238]),
    .I0(abar[14]),
    .I1(bbar[14])
  );
  //AND U104
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U104 (
    .O(y[237]),
    .I0(a[14]),
    .I1(b[13])
  );
  //OR U104bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U104bar (
    .O(ybar[237]),
    .I0(abar[14]),
    .I1(bbar[13])
  );
  //AND U105
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U105 (
    .O(y[236]),
    .I0(a[14]),
    .I1(b[12])
  );
  //OR U105bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U105bar (
    .O(ybar[236]),
    .I0(abar[14]),
    .I1(bbar[12])
  );
  //AND U106
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U106 (
    .O(y[235]),
    .I0(a[14]),
    .I1(b[11])
  );
  //OR U106bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U106bar (
    .O(ybar[235]),
    .I0(abar[14]),
    .I1(bbar[11])
  );
  //AND U107
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U107 (
    .O(y[234]),
    .I0(a[14]),
    .I1(b[10])
  );
  //OR U107bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U107bar (
    .O(ybar[234]),
    .I0(abar[14]),
    .I1(bbar[10])
  );
  //AND U108
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U108 (
    .O(y[233]),
    .I0(a[14]),
    .I1(b[9])
  );
  //OR U108bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U108bar (
    .O(ybar[233]),
    .I0(abar[14]),
    .I1(bbar[9])
  );
  //AND U109
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U109 (
    .O(y[232]),
    .I0(a[14]),
    .I1(b[8])
  );
  //OR U109bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U109bar (
    .O(ybar[232]),
    .I0(abar[14]),
    .I1(bbar[8])
  );
  //AND U110
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U110 (
    .O(y[231]),
    .I0(a[14]),
    .I1(b[7])
  );
  //OR U110bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U110bar (
    .O(ybar[231]),
    .I0(abar[14]),
    .I1(bbar[7])
  );
  //AND U111
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U111 (
    .O(y[230]),
    .I0(a[14]),
    .I1(b[6])
  );
  //OR U111bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U111bar (
    .O(ybar[230]),
    .I0(abar[14]),
    .I1(bbar[6])
  );
  //AND U112
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U112 (
    .O(y[22]),
    .I0(a[1]),
    .I1(b[6])
  );
  //OR U112bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U112bar (
    .O(ybar[22]),
    .I0(abar[1]),
    .I1(bbar[6])
  );
  //AND U113
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U113 (
    .O(y[229]),
    .I0(a[14]),
    .I1(b[5])
  );
  //OR U113bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U113bar (
    .O(ybar[229]),
    .I0(abar[14]),
    .I1(bbar[5])
  );
  //AND U114
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U114 (
    .O(y[228]),
    .I0(a[14]),
    .I1(b[4])
  );
  //OR U114bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U114bar (
    .O(ybar[228]),
    .I0(abar[14]),
    .I1(bbar[4])
  );
  //AND U115
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U115 (
    .O(y[227]),
    .I0(a[14]),
    .I1(b[3])
  );
  //OR U115bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U115bar (
    .O(ybar[227]),
    .I0(abar[14]),
    .I1(bbar[3])
  );
  //AND U116
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U116 (
    .O(y[226]),
    .I0(a[14]),
    .I1(b[2])
  );
  //OR U116bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U116bar (
    .O(ybar[226]),
    .I0(abar[14]),
    .I1(bbar[2])
  );
  //AND U117
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U117 (
    .O(y[225]),
    .I0(a[14]),
    .I1(b[1])
  );
  //OR U117bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U117bar (
    .O(ybar[225]),
    .I0(abar[14]),
    .I1(bbar[1])
  );
  //AND U118
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U118 (
    .O(y[224]),
    .I0(a[14]),
    .I1(b[0])
  );
  //OR U118bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U118bar (
    .O(ybar[224]),
    .I0(abar[14]),
    .I1(bbar[0])
  );
  //AND U119
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U119 (
    .O(y[223]),
    .I0(a[13]),
    .I1(b[15])
  );
  //OR U119bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U119bar (
    .O(ybar[223]),
    .I0(abar[13]),
    .I1(bbar[15])
  );
  //AND U120
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U120 (
    .O(y[222]),
    .I0(a[13]),
    .I1(b[14])
  );
  //OR U120bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U120bar (
    .O(ybar[222]),
    .I0(abar[13]),
    .I1(bbar[14])
  );
  //AND U121
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U121 (
    .O(y[221]),
    .I0(a[13]),
    .I1(b[13])
  );
  //OR U121bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U121bar (
    .O(ybar[221]),
    .I0(abar[13]),
    .I1(bbar[13])
  );
  //AND U122
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U122 (
    .O(y[220]),
    .I0(a[13]),
    .I1(b[12])
  );
  //OR U122bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U122bar (
    .O(ybar[220]),
    .I0(abar[13]),
    .I1(bbar[12])
  );
  //AND U123
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U123 (
    .O(y[21]),
    .I0(a[1]),
    .I1(b[5])
  );
  //OR U123bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U123bar (
    .O(ybar[21]),
    .I0(abar[1]),
    .I1(bbar[5])
  );
  //AND U124
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U124 (
    .O(y[219]),
    .I0(a[13]),
    .I1(b[11])
  );
  //OR U124bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U124bar (
    .O(ybar[219]),
    .I0(abar[13]),
    .I1(bbar[11])
  );
  //AND U125
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U125 (
    .O(y[218]),
    .I0(a[13]),
    .I1(b[10])
  );
  //OR U125bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U125bar (
    .O(ybar[218]),
    .I0(abar[13]),
    .I1(bbar[10])
  );
  //AND U126
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U126 (
    .O(y[217]),
    .I0(a[13]),
    .I1(b[9])
  );
  //OR U126bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U126bar (
    .O(ybar[217]),
    .I0(abar[13]),
    .I1(bbar[9])
  );
  //AND U127
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U127 (
    .O(y[216]),
    .I0(a[13]),
    .I1(b[8])
  );
  //OR U127bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U127bar (
    .O(ybar[216]),
    .I0(abar[13]),
    .I1(bbar[8])
  );
  //AND U128
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U128 (
    .O(y[215]),
    .I0(a[13]),
    .I1(b[7])
  );
  //OR U128bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U128bar (
    .O(ybar[215]),
    .I0(abar[13]),
    .I1(bbar[7])
  );
  //AND U129
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U129 (
    .O(y[214]),
    .I0(a[13]),
    .I1(b[6])
  );
  //OR U129bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U129bar (
    .O(ybar[214]),
    .I0(abar[13]),
    .I1(bbar[6])
  );
  //AND U130
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U130 (
    .O(y[213]),
    .I0(a[13]),
    .I1(b[5])
  );
  //OR U130bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U130bar (
    .O(ybar[213]),
    .I0(abar[13]),
    .I1(bbar[5])
  );
  //AND U131
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U131 (
    .O(y[212]),
    .I0(a[13]),
    .I1(b[4])
  );
  //OR U131bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U131bar (
    .O(ybar[212]),
    .I0(abar[13]),
    .I1(bbar[4])
  );
  //AND U132
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U132 (
    .O(y[211]),
    .I0(a[13]),
    .I1(b[3])
  );
  //OR U132bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U132bar (
    .O(ybar[211]),
    .I0(abar[13]),
    .I1(bbar[3])
  );
  //AND U133
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U133 (
    .O(y[210]),
    .I0(a[13]),
    .I1(b[2])
  );
  //OR U133bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U133bar (
    .O(ybar[210]),
    .I0(abar[13]),
    .I1(bbar[2])
  );
  //AND U134
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U134 (
    .O(y[20]),
    .I0(a[1]),
    .I1(b[4])
  );
  //OR U134bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U134bar (
    .O(ybar[20]),
    .I0(abar[1]),
    .I1(bbar[4])
  );
  //AND U135
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U135 (
    .O(y[209]),
    .I0(a[13]),
    .I1(b[1])
  );
  //OR U135bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U135bar (
    .O(ybar[209]),
    .I0(abar[13]),
    .I1(bbar[1])
  );
  //AND U136
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U136 (
    .O(y[208]),
    .I0(a[13]),
    .I1(b[0])
  );
  //OR U136bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U136bar (
    .O(ybar[208]),
    .I0(abar[13]),
    .I1(bbar[0])
  );
  //AND U137
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U137 (
    .O(y[207]),
    .I0(a[12]),
    .I1(b[15])
  );
  //OR U137bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U137bar (
    .O(ybar[207]),
    .I0(abar[12]),
    .I1(bbar[15])
  );
  //AND U138
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U138 (
    .O(y[206]),
    .I0(a[12]),
    .I1(b[14])
  );
  //OR U138bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U138bar (
    .O(ybar[206]),
    .I0(abar[12]),
    .I1(bbar[14])
  );
  //AND U139
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U139 (
    .O(y[205]),
    .I0(a[12]),
    .I1(b[13])
  );
  //OR U139bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U139bar (
    .O(ybar[205]),
    .I0(abar[12]),
    .I1(bbar[13])
  );
  //AND U140
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U140 (
    .O(y[204]),
    .I0(a[12]),
    .I1(b[12])
  );
  //OR U140bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U140bar (
    .O(ybar[204]),
    .I0(abar[12]),
    .I1(bbar[12])
  );
  //AND U141
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U141 (
    .O(y[203]),
    .I0(a[12]),
    .I1(b[11])
  );
  //OR U141bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U141bar (
    .O(ybar[203]),
    .I0(abar[12]),
    .I1(bbar[11])
  );
  //AND U142
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U142 (
    .O(y[202]),
    .I0(a[12]),
    .I1(b[10])
  );
  //OR U142bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U142bar (
    .O(ybar[202]),
    .I0(abar[12]),
    .I1(bbar[10])
  );
  //AND U143
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U143 (
    .O(y[201]),
    .I0(a[12]),
    .I1(b[9])
  );
  //OR U143bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U143bar (
    .O(ybar[201]),
    .I0(abar[12]),
    .I1(bbar[9])
  );
  //AND U144
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U144 (
    .O(y[200]),
    .I0(a[12]),
    .I1(b[8])
  );
  //OR U144bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U144bar (
    .O(ybar[200]),
    .I0(abar[12]),
    .I1(bbar[8])
  );
  //AND U145
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U145 (
    .O(y[1]),
    .I0(b[1]),
    .I1(a[0])
  );
  //OR U145bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U145bar (
    .O(ybar[1]),
    .I0(bbar[1]),
    .I1(abar[0])
  );
  //AND U146
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U146 (
    .O(y[19]),
    .I0(a[1]),
    .I1(b[3])
  );
  //OR U146bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U146bar (
    .O(ybar[19]),
    .I0(abar[1]),
    .I1(bbar[3])
  );
  //AND U147
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U147 (
    .O(y[199]),
    .I0(a[12]),
    .I1(b[7])
  );
  //OR U147bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U147bar (
    .O(ybar[199]),
    .I0(abar[12]),
    .I1(bbar[7])
  );
  //AND U148
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U148 (
    .O(y[198]),
    .I0(a[12]),
    .I1(b[6])
  );
  //OR U148bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U148bar (
    .O(ybar[198]),
    .I0(abar[12]),
    .I1(bbar[6])
  );
  //AND U149
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U149 (
    .O(y[197]),
    .I0(a[12]),
    .I1(b[5])
  );
  //OR U149bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U149bar (
    .O(ybar[197]),
    .I0(abar[12]),
    .I1(bbar[5])
  );
  //AND U150
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U150 (
    .O(y[196]),
    .I0(a[12]),
    .I1(b[4])
  );
  //OR U150bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U150bar (
    .O(ybar[196]),
    .I0(abar[12]),
    .I1(bbar[4])
  );
  //AND U151
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U151 (
    .O(y[195]),
    .I0(a[12]),
    .I1(b[3])
  );
  //OR U151bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U151bar (
    .O(ybar[195]),
    .I0(abar[12]),
    .I1(bbar[3])
  );
  //AND U152
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U152 (
    .O(y[194]),
    .I0(a[12]),
    .I1(b[2])
  );
  //OR U152bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U152bar (
    .O(ybar[194]),
    .I0(abar[12]),
    .I1(bbar[2])
  );
  //AND U153
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U153 (
    .O(y[193]),
    .I0(a[12]),
    .I1(b[1])
  );
  //OR U153bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U153bar (
    .O(ybar[193]),
    .I0(abar[12]),
    .I1(bbar[1])
  );
  //AND U154
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U154 (
    .O(y[192]),
    .I0(a[12]),
    .I1(b[0])
  );
  //OR U154bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U154bar (
    .O(ybar[192]),
    .I0(abar[12]),
    .I1(bbar[0])
  );
  //AND U155
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U155 (
    .O(y[191]),
    .I0(a[11]),
    .I1(b[15])
  );
  //OR U155bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U155bar (
    .O(ybar[191]),
    .I0(abar[11]),
    .I1(bbar[15])
  );
  //AND U156
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U156 (
    .O(y[190]),
    .I0(a[11]),
    .I1(b[14])
  );
  //OR U156bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U156bar (
    .O(ybar[190]),
    .I0(abar[11]),
    .I1(bbar[14])
  );
  //AND U157
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U157 (
    .O(y[18]),
    .I0(a[1]),
    .I1(b[2])
  );
  //OR U157bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U157bar (
    .O(ybar[18]),
    .I0(abar[1]),
    .I1(bbar[2])
  );
  //AND U158
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U158 (
    .O(y[189]),
    .I0(a[11]),
    .I1(b[13])
  );
  //OR U158bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U158bar (
    .O(ybar[189]),
    .I0(abar[11]),
    .I1(bbar[13])
  );
  //AND U159
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U159 (
    .O(y[188]),
    .I0(a[11]),
    .I1(b[12])
  );
  //OR U159bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U159bar (
    .O(ybar[188]),
    .I0(abar[11]),
    .I1(bbar[12])
  );
  //AND U160
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U160 (
    .O(y[187]),
    .I0(a[11]),
    .I1(b[11])
  );
  //OR U160bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U160bar (
    .O(ybar[187]),
    .I0(abar[11]),
    .I1(bbar[11])
  );
  //AND U161
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U161 (
    .O(y[186]),
    .I0(a[11]),
    .I1(b[10])
  );
  //OR U161bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U161bar (
    .O(ybar[186]),
    .I0(abar[11]),
    .I1(bbar[10])
  );
  //AND U162
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U162 (
    .O(y[185]),
    .I0(a[11]),
    .I1(b[9])
  );
  //OR U162bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U162bar (
    .O(ybar[185]),
    .I0(abar[11]),
    .I1(bbar[9])
  );
  //AND U163
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U163 (
    .O(y[184]),
    .I0(a[11]),
    .I1(b[8])
  );
  //OR U163bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U163bar (
    .O(ybar[184]),
    .I0(abar[11]),
    .I1(bbar[8])
  );
  //AND U164
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U164 (
    .O(y[183]),
    .I0(a[11]),
    .I1(b[7])
  );
  //OR U164bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U164bar (
    .O(ybar[183]),
    .I0(abar[11]),
    .I1(bbar[7])
  );
  //AND U165
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U165 (
    .O(y[182]),
    .I0(a[11]),
    .I1(b[6])
  );
  //OR U165bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U165bar (
    .O(ybar[182]),
    .I0(abar[11]),
    .I1(bbar[6])
  );
  //AND U166
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U166 (
    .O(y[181]),
    .I0(a[11]),
    .I1(b[5])
  );
  //OR U166bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U166bar (
    .O(ybar[181]),
    .I0(abar[11]),
    .I1(bbar[5])
  );
  //AND U167
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U167 (
    .O(y[180]),
    .I0(a[11]),
    .I1(b[4])
  );
  //OR U167bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U167bar (
    .O(ybar[180]),
    .I0(abar[11]),
    .I1(bbar[4])
  );
  //AND U168
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U168 (
    .O(y[17]),
    .I0(a[1]),
    .I1(b[1])
  );
  //OR U168bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U168bar (
    .O(ybar[17]),
    .I0(abar[1]),
    .I1(bbar[1])
  );
  //AND U169
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U169 (
    .O(y[179]),
    .I0(a[11]),
    .I1(b[3])
  );
  //OR U169bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U169bar (
    .O(ybar[179]),
    .I0(abar[11]),
    .I1(bbar[3])
  );
  //AND U170
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U170 (
    .O(y[178]),
    .I0(a[11]),
    .I1(b[2])
  );
  //OR U170bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U170bar (
    .O(ybar[178]),
    .I0(abar[11]),
    .I1(bbar[2])
  );
  //AND U171
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U171 (
    .O(y[177]),
    .I0(a[11]),
    .I1(b[1])
  );
  //OR U171bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U171bar (
    .O(ybar[177]),
    .I0(abar[11]),
    .I1(bbar[1])
  );
  //AND U172
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U172 (
    .O(y[176]),
    .I0(a[11]),
    .I1(b[0])
  );
  //OR U172bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U172bar (
    .O(ybar[176]),
    .I0(abar[11]),
    .I1(bbar[0])
  );
  //AND U173
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U173 (
    .O(y[175]),
    .I0(a[10]),
    .I1(b[15])
  );
  //OR U173bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U173bar (
    .O(ybar[175]),
    .I0(abar[10]),
    .I1(bbar[15])
  );
  //AND U174
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U174 (
    .O(y[174]),
    .I0(a[10]),
    .I1(b[14])
  );
  //OR U174bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U174bar (
    .O(ybar[174]),
    .I0(abar[10]),
    .I1(bbar[14])
  );
  //AND U175
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U175 (
    .O(y[173]),
    .I0(a[10]),
    .I1(b[13])
  );
  //OR U175bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U175bar (
    .O(ybar[173]),
    .I0(abar[10]),
    .I1(bbar[13])
  );
  //AND U176
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U176 (
    .O(y[172]),
    .I0(a[10]),
    .I1(b[12])
  );
  //OR U176bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U176bar (
    .O(ybar[172]),
    .I0(abar[10]),
    .I1(bbar[12])
  );
  //AND U177
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U177 (
    .O(y[171]),
    .I0(a[10]),
    .I1(b[11])
  );
  //OR U177bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U177bar (
    .O(ybar[171]),
    .I0(abar[10]),
    .I1(bbar[11])
  );
  //AND U178
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U178 (
    .O(y[170]),
    .I0(a[10]),
    .I1(b[10])
  );
  //OR U178bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U178bar (
    .O(ybar[170]),
    .I0(abar[10]),
    .I1(bbar[10])
  );
  //AND U179
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U179 (
    .O(y[16]),
    .I0(a[1]),
    .I1(b[0])
  );
  //OR U179bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U179bar (
    .O(ybar[16]),
    .I0(abar[1]),
    .I1(bbar[0])
  );
  //AND U180
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U180 (
    .O(y[169]),
    .I0(a[10]),
    .I1(b[9])
  );
  //OR U180bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U180bar (
    .O(ybar[169]),
    .I0(abar[10]),
    .I1(bbar[9])
  );
  //AND U181
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U181 (
    .O(y[168]),
    .I0(a[10]),
    .I1(b[8])
  );
  //OR U181bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U181bar (
    .O(ybar[168]),
    .I0(abar[10]),
    .I1(bbar[8])
  );
  //AND U182
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U182 (
    .O(y[167]),
    .I0(a[10]),
    .I1(b[7])
  );
  //OR U182bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U182bar (
    .O(ybar[167]),
    .I0(abar[10]),
    .I1(bbar[7])
  );
  //AND U183
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U183 (
    .O(y[166]),
    .I0(a[10]),
    .I1(b[6])
  );
  //OR U183bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U183bar (
    .O(ybar[166]),
    .I0(abar[10]),
    .I1(bbar[6])
  );
  //AND U184
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U184 (
    .O(y[165]),
    .I0(a[10]),
    .I1(b[5])
  );
  //OR U184bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U184bar (
    .O(ybar[165]),
    .I0(abar[10]),
    .I1(bbar[5])
  );
  //AND U185
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U185 (
    .O(y[164]),
    .I0(a[10]),
    .I1(b[4])
  );
  //OR U185bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U185bar (
    .O(ybar[164]),
    .I0(abar[10]),
    .I1(bbar[4])
  );
  //AND U186
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U186 (
    .O(y[163]),
    .I0(a[10]),
    .I1(b[3])
  );
  //OR U186bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U186bar (
    .O(ybar[163]),
    .I0(abar[10]),
    .I1(bbar[3])
  );
  //AND U187
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U187 (
    .O(y[162]),
    .I0(a[10]),
    .I1(b[2])
  );
  //OR U187bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U187bar (
    .O(ybar[162]),
    .I0(abar[10]),
    .I1(bbar[2])
  );
  //AND U188
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U188 (
    .O(y[161]),
    .I0(a[10]),
    .I1(b[1])
  );
  //OR U188bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U188bar (
    .O(ybar[161]),
    .I0(abar[10]),
    .I1(bbar[1])
  );
  //AND U189
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U189 (
    .O(y[160]),
    .I0(a[10]),
    .I1(b[0])
  );
  //OR U189bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U189bar (
    .O(ybar[160]),
    .I0(abar[10]),
    .I1(bbar[0])
  );
  //AND U190
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U190 (
    .O(y[15]),
    .I0(b[15]),
    .I1(a[0])
  );
  //OR U190bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U190bar (
    .O(ybar[15]),
    .I0(bbar[15]),
    .I1(abar[0])
  );
  //AND U191
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U191 (
    .O(y[159]),
    .I0(a[9]),
    .I1(b[15])
  );
  //OR U191bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U191bar (
    .O(ybar[159]),
    .I0(abar[9]),
    .I1(bbar[15])
  );
  //AND U192
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U192 (
    .O(y[158]),
    .I0(a[9]),
    .I1(b[14])
  );
  //OR U192bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U192bar (
    .O(ybar[158]),
    .I0(abar[9]),
    .I1(bbar[14])
  );
  //AND U193
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U193 (
    .O(y[157]),
    .I0(a[9]),
    .I1(b[13])
  );
  //OR U193bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U193bar (
    .O(ybar[157]),
    .I0(abar[9]),
    .I1(bbar[13])
  );
  //AND U194
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U194 (
    .O(y[156]),
    .I0(a[9]),
    .I1(b[12])
  );
  //OR U194bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U194bar (
    .O(ybar[156]),
    .I0(abar[9]),
    .I1(bbar[12])
  );
  //AND U195
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U195 (
    .O(y[155]),
    .I0(a[9]),
    .I1(b[11])
  );
  //OR U195bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U195bar (
    .O(ybar[155]),
    .I0(abar[9]),
    .I1(bbar[11])
  );
  //AND U196
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U196 (
    .O(y[154]),
    .I0(a[9]),
    .I1(b[10])
  );
  //OR U196bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U196bar (
    .O(ybar[154]),
    .I0(abar[9]),
    .I1(bbar[10])
  );
  //AND U197
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U197 (
    .O(y[153]),
    .I0(a[9]),
    .I1(b[9])
  );
  //OR U197bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U197bar (
    .O(ybar[153]),
    .I0(abar[9]),
    .I1(bbar[9])
  );
  //AND U198
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U198 (
    .O(y[152]),
    .I0(a[9]),
    .I1(b[8])
  );
  //OR U198bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U198bar (
    .O(ybar[152]),
    .I0(abar[9]),
    .I1(bbar[8])
  );
  //AND U199
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U199 (
    .O(y[151]),
    .I0(a[9]),
    .I1(b[7])
  );
  //OR U199bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U199bar (
    .O(ybar[151]),
    .I0(abar[9]),
    .I1(bbar[7])
  );
  //AND U200
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U200 (
    .O(y[150]),
    .I0(a[9]),
    .I1(b[6])
  );
  //OR U200bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U200bar (
    .O(ybar[150]),
    .I0(abar[9]),
    .I1(bbar[6])
  );
  //AND U201
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U201 (
    .O(y[14]),
    .I0(b[14]),
    .I1(a[0])
  );
  //OR U201bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U201bar (
    .O(ybar[14]),
    .I0(bbar[14]),
    .I1(abar[0])
  );
  //AND U202
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U202 (
    .O(y[149]),
    .I0(a[9]),
    .I1(b[5])
  );
  //OR U202bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U202bar (
    .O(ybar[149]),
    .I0(abar[9]),
    .I1(bbar[5])
  );
  //AND U203
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U203 (
    .O(y[148]),
    .I0(a[9]),
    .I1(b[4])
  );
  //OR U203bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U203bar (
    .O(ybar[148]),
    .I0(abar[9]),
    .I1(bbar[4])
  );
  //AND U204
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U204 (
    .O(y[147]),
    .I0(a[9]),
    .I1(b[3])
  );
  //OR U204bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U204bar (
    .O(ybar[147]),
    .I0(abar[9]),
    .I1(bbar[3])
  );
  //AND U205
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U205 (
    .O(y[146]),
    .I0(a[9]),
    .I1(b[2])
  );
  //OR U205bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U205bar (
    .O(ybar[146]),
    .I0(abar[9]),
    .I1(bbar[2])
  );
  //AND U206
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U206 (
    .O(y[145]),
    .I0(a[9]),
    .I1(b[1])
  );
  //OR U206bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U206bar (
    .O(ybar[145]),
    .I0(abar[9]),
    .I1(bbar[1])
  );
  //AND U207
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U207 (
    .O(y[144]),
    .I0(a[9]),
    .I1(b[0])
  );
  //OR U207bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U207bar (
    .O(ybar[144]),
    .I0(abar[9]),
    .I1(bbar[0])
  );
  //AND U208
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U208 (
    .O(y[143]),
    .I0(a[8]),
    .I1(b[15])
  );
  //OR U208bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U208bar (
    .O(ybar[143]),
    .I0(abar[8]),
    .I1(bbar[15])
  );
  //AND U209
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U209 (
    .O(y[142]),
    .I0(a[8]),
    .I1(b[14])
  );
  //OR U209bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U209bar (
    .O(ybar[142]),
    .I0(abar[8]),
    .I1(bbar[14])
  );
  //AND U210
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U210 (
    .O(y[141]),
    .I0(a[8]),
    .I1(b[13])
  );
  //OR U210bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U210bar (
    .O(ybar[141]),
    .I0(abar[8]),
    .I1(bbar[13])
  );
  //AND U211
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U211 (
    .O(y[140]),
    .I0(a[8]),
    .I1(b[12])
  );
  //OR U211bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U211bar (
    .O(ybar[140]),
    .I0(abar[8]),
    .I1(bbar[12])
  );
  //AND U212
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U212 (
    .O(y[13]),
    .I0(b[13]),
    .I1(a[0])
  );
  //OR U212bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U212bar (
    .O(ybar[13]),
    .I0(bbar[13]),
    .I1(abar[0])
  );
  //AND U213
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U213 (
    .O(y[139]),
    .I0(a[8]),
    .I1(b[11])
  );
  //OR U213bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U213bar (
    .O(ybar[139]),
    .I0(abar[8]),
    .I1(bbar[11])
  );
  //AND U214
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U214 (
    .O(y[138]),
    .I0(a[8]),
    .I1(b[10])
  );
  //OR U214bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U214bar (
    .O(ybar[138]),
    .I0(abar[8]),
    .I1(bbar[10])
  );
  //AND U215
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U215 (
    .O(y[137]),
    .I0(a[8]),
    .I1(b[9])
  );
  //OR U215bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U215bar (
    .O(ybar[137]),
    .I0(abar[8]),
    .I1(bbar[9])
  );
  //AND U216
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U216 (
    .O(y[136]),
    .I0(a[8]),
    .I1(b[8])
  );
  //OR U216bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U216bar (
    .O(ybar[136]),
    .I0(abar[8]),
    .I1(bbar[8])
  );
  //AND U217
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U217 (
    .O(y[135]),
    .I0(a[8]),
    .I1(b[7])
  );
  //OR U217bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U217bar (
    .O(ybar[135]),
    .I0(abar[8]),
    .I1(bbar[7])
  );
  //AND U218
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U218 (
    .O(y[134]),
    .I0(a[8]),
    .I1(b[6])
  );
  //OR U218bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U218bar (
    .O(ybar[134]),
    .I0(abar[8]),
    .I1(bbar[6])
  );
  //AND U219
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U219 (
    .O(y[133]),
    .I0(a[8]),
    .I1(b[5])
  );
  //OR U219bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U219bar (
    .O(ybar[133]),
    .I0(abar[8]),
    .I1(bbar[5])
  );
  //AND U220
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U220 (
    .O(y[132]),
    .I0(a[8]),
    .I1(b[4])
  );
  //OR U220bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U220bar (
    .O(ybar[132]),
    .I0(abar[8]),
    .I1(bbar[4])
  );
  //AND U221
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U221 (
    .O(y[131]),
    .I0(a[8]),
    .I1(b[3])
  );
  //OR U221bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U221bar (
    .O(ybar[131]),
    .I0(abar[8]),
    .I1(bbar[3])
  );
  //AND U222
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U222 (
    .O(y[130]),
    .I0(a[8]),
    .I1(b[2])
  );
  //OR U222bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U222bar (
    .O(ybar[130]),
    .I0(abar[8]),
    .I1(bbar[2])
  );
  //AND U223
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U223 (
    .O(y[12]),
    .I0(b[12]),
    .I1(a[0])
  );
  //OR U223bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U223bar (
    .O(ybar[12]),
    .I0(bbar[12]),
    .I1(abar[0])
  );
  //AND U224
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U224 (
    .O(y[129]),
    .I0(a[8]),
    .I1(b[1])
  );
  //OR U224bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U224bar (
    .O(ybar[129]),
    .I0(abar[8]),
    .I1(bbar[1])
  );
  //AND U225
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U225 (
    .O(y[128]),
    .I0(a[8]),
    .I1(b[0])
  );
  //OR U225bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U225bar (
    .O(ybar[128]),
    .I0(abar[8]),
    .I1(bbar[0])
  );
  //AND U226
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U226 (
    .O(y[127]),
    .I0(a[7]),
    .I1(b[15])
  );
  //OR U226bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U226bar (
    .O(ybar[127]),
    .I0(abar[7]),
    .I1(bbar[15])
  );
  //AND U227
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U227 (
    .O(y[126]),
    .I0(a[7]),
    .I1(b[14])
  );
  //OR U227bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U227bar (
    .O(ybar[126]),
    .I0(abar[7]),
    .I1(bbar[14])
  );
  //AND U228
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U228 (
    .O(y[125]),
    .I0(a[7]),
    .I1(b[13])
  );
  //OR U228bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U228bar (
    .O(ybar[125]),
    .I0(abar[7]),
    .I1(bbar[13])
  );
  //AND U229
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U229 (
    .O(y[124]),
    .I0(a[7]),
    .I1(b[12])
  );
  //OR U229bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U229bar (
    .O(ybar[124]),
    .I0(abar[7]),
    .I1(bbar[12])
  );
  //AND U230
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U230 (
    .O(y[123]),
    .I0(a[7]),
    .I1(b[11])
  );
  //OR U230bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U230bar (
    .O(ybar[123]),
    .I0(abar[7]),
    .I1(bbar[11])
  );
  //AND U231
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U231 (
    .O(y[122]),
    .I0(a[7]),
    .I1(b[10])
  );
  //OR U231bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U231bar (
    .O(ybar[122]),
    .I0(abar[7]),
    .I1(bbar[10])
  );
  //AND U232
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U232 (
    .O(y[121]),
    .I0(a[7]),
    .I1(b[9])
  );
  //OR U232bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U232bar (
    .O(ybar[121]),
    .I0(abar[7]),
    .I1(bbar[9])
  );
  //AND U233
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U233 (
    .O(y[120]),
    .I0(a[7]),
    .I1(b[8])
  );
  //OR U233bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U233bar (
    .O(ybar[120]),
    .I0(abar[7]),
    .I1(bbar[8])
  );
  //AND U234
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U234 (
    .O(y[11]),
    .I0(b[11]),
    .I1(a[0])
  );
  //OR U234bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U234bar (
    .O(ybar[11]),
    .I0(bbar[11]),
    .I1(abar[0])
  );
  //AND U235
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U235 (
    .O(y[119]),
    .I0(a[7]),
    .I1(b[7])
  );
  //OR U235bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U235bar (
    .O(ybar[119]),
    .I0(abar[7]),
    .I1(bbar[7])
  );
  //AND U236
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U236 (
    .O(y[118]),
    .I0(a[7]),
    .I1(b[6])
  );
  //OR U236bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U236bar (
    .O(ybar[118]),
    .I0(abar[7]),
    .I1(bbar[6])
  );
  //AND U237
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U237 (
    .O(y[117]),
    .I0(a[7]),
    .I1(b[5])
  );
  //OR U237bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U237bar (
    .O(ybar[117]),
    .I0(abar[7]),
    .I1(bbar[5])
  );
  //AND U238
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U238 (
    .O(y[116]),
    .I0(a[7]),
    .I1(b[4])
  );
  //OR U238bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U238bar (
    .O(ybar[116]),
    .I0(abar[7]),
    .I1(bbar[4])
  );
  //AND U239
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U239 (
    .O(y[115]),
    .I0(a[7]),
    .I1(b[3])
  );
  //OR U239bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U239bar (
    .O(ybar[115]),
    .I0(abar[7]),
    .I1(bbar[3])
  );
  //AND U240
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U240 (
    .O(y[114]),
    .I0(a[7]),
    .I1(b[2])
  );
  //OR U240bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U240bar (
    .O(ybar[114]),
    .I0(abar[7]),
    .I1(bbar[2])
  );
  //AND U241
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U241 (
    .O(y[113]),
    .I0(a[7]),
    .I1(b[1])
  );
  //OR U241bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U241bar (
    .O(ybar[113]),
    .I0(abar[7]),
    .I1(bbar[1])
  );
  //AND U242
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U242 (
    .O(y[112]),
    .I0(a[7]),
    .I1(b[0])
  );
  //OR U242bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U242bar (
    .O(ybar[112]),
    .I0(abar[7]),
    .I1(bbar[0])
  );
  //AND U243
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U243 (
    .O(y[111]),
    .I0(b[15]),
    .I1(a[6])
  );
  //OR U243bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U243bar (
    .O(ybar[111]),
    .I0(bbar[15]),
    .I1(abar[6])
  );
  //AND U244
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U244 (
    .O(y[110]),
    .I0(b[14]),
    .I1(a[6])
  );
  //OR U244bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U244bar (
    .O(ybar[110]),
    .I0(bbar[14]),
    .I1(abar[6])
  );
  //AND U245
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U245 (
    .O(y[10]),
    .I0(b[10]),
    .I1(a[0])
  );
  //OR U245bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U245bar (
    .O(ybar[10]),
    .I0(bbar[10]),
    .I1(abar[0])
  );
  //AND U246
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U246 (
    .O(y[109]),
    .I0(b[13]),
    .I1(a[6])
  );
  //OR U246bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U246bar (
    .O(ybar[109]),
    .I0(bbar[13]),
    .I1(abar[6])
  );
  //AND U247
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U247 (
    .O(y[108]),
    .I0(b[12]),
    .I1(a[6])
  );
  //OR U247bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U247bar (
    .O(ybar[108]),
    .I0(bbar[12]),
    .I1(abar[6])
  );
  //AND U248
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U248 (
    .O(y[107]),
    .I0(b[11]),
    .I1(a[6])
  );
  //OR U248bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U248bar (
    .O(ybar[107]),
    .I0(bbar[11]),
    .I1(abar[6])
  );
  //AND U249
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U249 (
    .O(y[106]),
    .I0(b[10]),
    .I1(a[6])
  );
  //OR U249bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U249bar (
    .O(ybar[106]),
    .I0(bbar[10]),
    .I1(abar[6])
  );
  //AND U250
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U250 (
    .O(y[105]),
    .I0(a[6]),
    .I1(b[9])
  );
  //OR U250bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U250bar (
    .O(ybar[105]),
    .I0(abar[6]),
    .I1(bbar[9])
  );
  //AND U251
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U251 (
    .O(y[104]),
    .I0(b[8]),
    .I1(a[6])
  );
  //OR U251bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U251bar (
    .O(ybar[104]),
    .I0(bbar[8]),
    .I1(abar[6])
  );
  //AND U252
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U252 (
    .O(y[103]),
    .I0(b[7]),
    .I1(a[6])
  );
  //OR U252bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U252bar (
    .O(ybar[103]),
    .I0(bbar[7]),
    .I1(abar[6])
  );
  //AND U253
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U253 (
    .O(y[102]),
    .I0(b[6]),
    .I1(a[6])
  );
  //OR U253bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U253bar (
    .O(ybar[102]),
    .I0(bbar[6]),
    .I1(abar[6])
  );
  //AND U254
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U254 (
    .O(y[101]),
    .I0(b[5]),
    .I1(a[6])
  );
  //OR U254bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U254bar (
    .O(ybar[101]),
    .I0(bbar[5]),
    .I1(abar[6])
  );
  //AND U255
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U255 (
    .O(y[100]),
    .I0(b[4]),
    .I1(a[6])
  );
  //OR U255bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U255bar (
    .O(ybar[100]),
    .I0(bbar[4]),
    .I1(abar[6])
  );
  //AND U256
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U256 (
    .O(y[0]),
    .I0(b[0]),
    .I1(a[0])
  );
  //OR U256bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U256bar (
    .O(ybar[0]),
    .I0(bbar[0]),
    .I1(abar[0])
  );
endmodule

module decode_12 ( in, out );

  input wire [7:0] in;
//input_done

  output wire [255:0] out;
//output_done

  wire [15:0] level1;
  wire [31:0] level2;
//wire_done

  CD2_48 cd_l1_1 ( .a(in[1]), .b(in[0]), .y(level1[3:0]) );
  CD2_47 cd_l1_2 ( .a(in[3]), .b(in[2]), .y(level1[7:4]) );
  CD2_46 cd_l1_3 ( .a(in[5]), .b(in[4]), .y(level1[11:8]) );
  CD2_45 cd_l1_4 ( .a(in[7]), .b(in[6]), .y(level1[15:12]) );
  CD4_24 cd_l2_1 ( .a(level1[7:4]), .b(level1[3:0]), .y(level2[15:0]) );
  CD4_23 cd_l2_2 ( .a(level1[15:12]), .b(level1[11:8]), .y(level2[31:16]) );
  CD16_12 cd_l3 ( .a(level2[31:16]), .b(level2[15:0]), .y(out) );
endmodule

module encode_12 ( in, out );

  input wire [255:0] in;
  wire [255:0] inbar;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
  assign inbar[8] = ~in[8];
  assign inbar[9] = ~in[9];
  assign inbar[10] = ~in[10];
  assign inbar[11] = ~in[11];
  assign inbar[12] = ~in[12];
  assign inbar[13] = ~in[13];
  assign inbar[14] = ~in[14];
  assign inbar[15] = ~in[15];
  assign inbar[16] = ~in[16];
  assign inbar[17] = ~in[17];
  assign inbar[18] = ~in[18];
  assign inbar[19] = ~in[19];
  assign inbar[20] = ~in[20];
  assign inbar[21] = ~in[21];
  assign inbar[22] = ~in[22];
  assign inbar[23] = ~in[23];
  assign inbar[24] = ~in[24];
  assign inbar[25] = ~in[25];
  assign inbar[26] = ~in[26];
  assign inbar[27] = ~in[27];
  assign inbar[28] = ~in[28];
  assign inbar[29] = ~in[29];
  assign inbar[30] = ~in[30];
  assign inbar[31] = ~in[31];
  assign inbar[32] = ~in[32];
  assign inbar[33] = ~in[33];
  assign inbar[34] = ~in[34];
  assign inbar[35] = ~in[35];
  assign inbar[36] = ~in[36];
  assign inbar[37] = ~in[37];
  assign inbar[38] = ~in[38];
  assign inbar[39] = ~in[39];
  assign inbar[40] = ~in[40];
  assign inbar[41] = ~in[41];
  assign inbar[42] = ~in[42];
  assign inbar[43] = ~in[43];
  assign inbar[44] = ~in[44];
  assign inbar[45] = ~in[45];
  assign inbar[46] = ~in[46];
  assign inbar[47] = ~in[47];
  assign inbar[48] = ~in[48];
  assign inbar[49] = ~in[49];
  assign inbar[50] = ~in[50];
  assign inbar[51] = ~in[51];
  assign inbar[52] = ~in[52];
  assign inbar[53] = ~in[53];
  assign inbar[54] = ~in[54];
  assign inbar[55] = ~in[55];
  assign inbar[56] = ~in[56];
  assign inbar[57] = ~in[57];
  assign inbar[58] = ~in[58];
  assign inbar[59] = ~in[59];
  assign inbar[60] = ~in[60];
  assign inbar[61] = ~in[61];
  assign inbar[62] = ~in[62];
  assign inbar[63] = ~in[63];
  assign inbar[64] = ~in[64];
  assign inbar[65] = ~in[65];
  assign inbar[66] = ~in[66];
  assign inbar[67] = ~in[67];
  assign inbar[68] = ~in[68];
  assign inbar[69] = ~in[69];
  assign inbar[70] = ~in[70];
  assign inbar[71] = ~in[71];
  assign inbar[72] = ~in[72];
  assign inbar[73] = ~in[73];
  assign inbar[74] = ~in[74];
  assign inbar[75] = ~in[75];
  assign inbar[76] = ~in[76];
  assign inbar[77] = ~in[77];
  assign inbar[78] = ~in[78];
  assign inbar[79] = ~in[79];
  assign inbar[80] = ~in[80];
  assign inbar[81] = ~in[81];
  assign inbar[82] = ~in[82];
  assign inbar[83] = ~in[83];
  assign inbar[84] = ~in[84];
  assign inbar[85] = ~in[85];
  assign inbar[86] = ~in[86];
  assign inbar[87] = ~in[87];
  assign inbar[88] = ~in[88];
  assign inbar[89] = ~in[89];
  assign inbar[90] = ~in[90];
  assign inbar[91] = ~in[91];
  assign inbar[92] = ~in[92];
  assign inbar[93] = ~in[93];
  assign inbar[94] = ~in[94];
  assign inbar[95] = ~in[95];
  assign inbar[96] = ~in[96];
  assign inbar[97] = ~in[97];
  assign inbar[98] = ~in[98];
  assign inbar[99] = ~in[99];
  assign inbar[100] = ~in[100];
  assign inbar[101] = ~in[101];
  assign inbar[102] = ~in[102];
  assign inbar[103] = ~in[103];
  assign inbar[104] = ~in[104];
  assign inbar[105] = ~in[105];
  assign inbar[106] = ~in[106];
  assign inbar[107] = ~in[107];
  assign inbar[108] = ~in[108];
  assign inbar[109] = ~in[109];
  assign inbar[110] = ~in[110];
  assign inbar[111] = ~in[111];
  assign inbar[112] = ~in[112];
  assign inbar[113] = ~in[113];
  assign inbar[114] = ~in[114];
  assign inbar[115] = ~in[115];
  assign inbar[116] = ~in[116];
  assign inbar[117] = ~in[117];
  assign inbar[118] = ~in[118];
  assign inbar[119] = ~in[119];
  assign inbar[120] = ~in[120];
  assign inbar[121] = ~in[121];
  assign inbar[122] = ~in[122];
  assign inbar[123] = ~in[123];
  assign inbar[124] = ~in[124];
  assign inbar[125] = ~in[125];
  assign inbar[126] = ~in[126];
  assign inbar[127] = ~in[127];
  assign inbar[128] = ~in[128];
  assign inbar[129] = ~in[129];
  assign inbar[130] = ~in[130];
  assign inbar[131] = ~in[131];
  assign inbar[132] = ~in[132];
  assign inbar[133] = ~in[133];
  assign inbar[134] = ~in[134];
  assign inbar[135] = ~in[135];
  assign inbar[136] = ~in[136];
  assign inbar[137] = ~in[137];
  assign inbar[138] = ~in[138];
  assign inbar[139] = ~in[139];
  assign inbar[140] = ~in[140];
  assign inbar[141] = ~in[141];
  assign inbar[142] = ~in[142];
  assign inbar[143] = ~in[143];
  assign inbar[144] = ~in[144];
  assign inbar[145] = ~in[145];
  assign inbar[146] = ~in[146];
  assign inbar[147] = ~in[147];
  assign inbar[148] = ~in[148];
  assign inbar[149] = ~in[149];
  assign inbar[150] = ~in[150];
  assign inbar[151] = ~in[151];
  assign inbar[152] = ~in[152];
  assign inbar[153] = ~in[153];
  assign inbar[154] = ~in[154];
  assign inbar[155] = ~in[155];
  assign inbar[156] = ~in[156];
  assign inbar[157] = ~in[157];
  assign inbar[158] = ~in[158];
  assign inbar[159] = ~in[159];
  assign inbar[160] = ~in[160];
  assign inbar[161] = ~in[161];
  assign inbar[162] = ~in[162];
  assign inbar[163] = ~in[163];
  assign inbar[164] = ~in[164];
  assign inbar[165] = ~in[165];
  assign inbar[166] = ~in[166];
  assign inbar[167] = ~in[167];
  assign inbar[168] = ~in[168];
  assign inbar[169] = ~in[169];
  assign inbar[170] = ~in[170];
  assign inbar[171] = ~in[171];
  assign inbar[172] = ~in[172];
  assign inbar[173] = ~in[173];
  assign inbar[174] = ~in[174];
  assign inbar[175] = ~in[175];
  assign inbar[176] = ~in[176];
  assign inbar[177] = ~in[177];
  assign inbar[178] = ~in[178];
  assign inbar[179] = ~in[179];
  assign inbar[180] = ~in[180];
  assign inbar[181] = ~in[181];
  assign inbar[182] = ~in[182];
  assign inbar[183] = ~in[183];
  assign inbar[184] = ~in[184];
  assign inbar[185] = ~in[185];
  assign inbar[186] = ~in[186];
  assign inbar[187] = ~in[187];
  assign inbar[188] = ~in[188];
  assign inbar[189] = ~in[189];
  assign inbar[190] = ~in[190];
  assign inbar[191] = ~in[191];
  assign inbar[192] = ~in[192];
  assign inbar[193] = ~in[193];
  assign inbar[194] = ~in[194];
  assign inbar[195] = ~in[195];
  assign inbar[196] = ~in[196];
  assign inbar[197] = ~in[197];
  assign inbar[198] = ~in[198];
  assign inbar[199] = ~in[199];
  assign inbar[200] = ~in[200];
  assign inbar[201] = ~in[201];
  assign inbar[202] = ~in[202];
  assign inbar[203] = ~in[203];
  assign inbar[204] = ~in[204];
  assign inbar[205] = ~in[205];
  assign inbar[206] = ~in[206];
  assign inbar[207] = ~in[207];
  assign inbar[208] = ~in[208];
  assign inbar[209] = ~in[209];
  assign inbar[210] = ~in[210];
  assign inbar[211] = ~in[211];
  assign inbar[212] = ~in[212];
  assign inbar[213] = ~in[213];
  assign inbar[214] = ~in[214];
  assign inbar[215] = ~in[215];
  assign inbar[216] = ~in[216];
  assign inbar[217] = ~in[217];
  assign inbar[218] = ~in[218];
  assign inbar[219] = ~in[219];
  assign inbar[220] = ~in[220];
  assign inbar[221] = ~in[221];
  assign inbar[222] = ~in[222];
  assign inbar[223] = ~in[223];
  assign inbar[224] = ~in[224];
  assign inbar[225] = ~in[225];
  assign inbar[226] = ~in[226];
  assign inbar[227] = ~in[227];
  assign inbar[228] = ~in[228];
  assign inbar[229] = ~in[229];
  assign inbar[230] = ~in[230];
  assign inbar[231] = ~in[231];
  assign inbar[232] = ~in[232];
  assign inbar[233] = ~in[233];
  assign inbar[234] = ~in[234];
  assign inbar[235] = ~in[235];
  assign inbar[236] = ~in[236];
  assign inbar[237] = ~in[237];
  assign inbar[238] = ~in[238];
  assign inbar[239] = ~in[239];
  assign inbar[240] = ~in[240];
  assign inbar[241] = ~in[241];
  assign inbar[242] = ~in[242];
  assign inbar[243] = ~in[243];
  assign inbar[244] = ~in[244];
  assign inbar[245] = ~in[245];
  assign inbar[246] = ~in[246];
  assign inbar[247] = ~in[247];
  assign inbar[248] = ~in[248];
  assign inbar[249] = ~in[249];
  assign inbar[250] = ~in[250];
  assign inbar[251] = ~in[251];
  assign inbar[252] = ~in[252];
  assign inbar[253] = ~in[253];
  assign inbar[254] = ~in[254];
  assign inbar[255] = ~in[255];
//input_done

  output wire [7:0] out;
  wire [7:0] outbar;
//output_done

  wire in_81;
  wire in_80;
  wire in_79;
  wire in_78;
  wire in_77;
  wire in_76;
  wire in_75;
  wire in_74;
  wire in_73;
  wire in_72;
  wire in_71;
  wire in_70;
  wire in_69;
  wire in_68;
  wire in_67;
  wire in_66;
  wire in_65;
  wire in_64;
  wire in_63;
  wire in_62;
  wire in_61;
  wire in_60;
  wire in_59;
  wire in_58;
  wire in_57;
  wire in_56;
  wire in_55;
  wire in_54;
  wire in_53;
  wire in_52;
  wire in_51;
  wire in_50;
  wire in_49;
  wire in_48;
  wire in_47;
  wire in_46;
  wire in_45;
  wire in_44;
  wire in_43;
  wire in_42;
  wire in_41;
  wire in_40;
  wire in_39;
  wire in_38;
  wire in_37;
  wire in_36;
  wire in_35;
  wire in_34;
  wire in_33;
  wire in_32;
  wire in_31;
  wire in_30;
  wire in_29;
  wire in_28;
  wire in_27;
  wire in_26;
  wire in_25;
  wire in_24;
  wire in_23;
  wire in_22;
  wire in_21;
  wire in_20;
  wire in_19;
  wire in_18;
  wire in_17;
  wire in_16;
  wire in_15;
  wire in_14;
  wire in_13;
  wire in_12;
  wire in_11;
  wire in_10;
  wire in_9;
  wire in_8;
  wire in_7;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_3;
  wire in_2;
  wire in_1;
  wire in_0;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire in_81bar;
  wire in_80bar;
  wire in_79bar;
  wire in_78bar;
  wire in_77bar;
  wire in_76bar;
  wire in_75bar;
  wire in_74bar;
  wire in_73bar;
  wire in_72bar;
  wire in_71bar;
  wire in_70bar;
  wire in_69bar;
  wire in_68bar;
  wire in_67bar;
  wire in_66bar;
  wire in_65bar;
  wire in_64bar;
  wire in_63bar;
  wire in_62bar;
  wire in_61bar;
  wire in_60bar;
  wire in_59bar;
  wire in_58bar;
  wire in_57bar;
  wire in_56bar;
  wire in_55bar;
  wire in_54bar;
  wire in_53bar;
  wire in_52bar;
  wire in_51bar;
  wire in_50bar;
  wire in_49bar;
  wire in_48bar;
  wire in_47bar;
  wire in_46bar;
  wire in_45bar;
  wire in_44bar;
  wire in_43bar;
  wire in_42bar;
  wire in_41bar;
  wire in_40bar;
  wire in_39bar;
  wire in_38bar;
  wire in_37bar;
  wire in_36bar;
  wire in_35bar;
  wire in_34bar;
  wire in_33bar;
  wire in_32bar;
  wire in_31bar;
  wire in_30bar;
  wire in_29bar;
  wire in_28bar;
  wire in_27bar;
  wire in_26bar;
  wire in_25bar;
  wire in_24bar;
  wire in_23bar;
  wire in_22bar;
  wire in_21bar;
  wire in_20bar;
  wire in_19bar;
  wire in_18bar;
  wire in_17bar;
  wire in_16bar;
  wire in_15bar;
  wire in_14bar;
  wire in_13bar;
  wire in_12bar;
  wire in_11bar;
  wire in_10bar;
  wire in_9bar;
  wire in_8bar;
  wire in_7bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_3bar;
  wire in_2bar;
  wire in_1bar;
  wire in_0bar;
  wire n487bar;
  wire n488bar;
  wire n489bar;
  wire n490bar;
  wire n491bar;
  wire n492bar;
  wire n493bar;
  wire n494bar;
  wire n495bar;
  wire n496bar;
  wire n497bar;
  wire n498bar;
  wire n499bar;
  wire n500bar;
  wire n501bar;
  wire n502bar;
  wire n503bar;
  wire n504bar;
  wire n505bar;
  wire n506bar;
  wire n507bar;
  wire n508bar;
  wire n509bar;
  wire n510bar;
  wire n511bar;
  wire n512bar;
  wire n513bar;
  wire n514bar;
  wire n515bar;
  wire n516bar;
  wire n517bar;
  wire n518bar;
  wire n519bar;
  wire n520bar;
  wire n521bar;
  wire n522bar;
  wire n523bar;
  wire n524bar;
  wire n525bar;
  wire n526bar;
  wire n527bar;
  wire n528bar;
  wire n529bar;
  wire n530bar;
  wire n531bar;
  wire n532bar;
  wire n533bar;
  wire n534bar;
  wire n535bar;
  wire n536bar;
  wire n537bar;
  wire n538bar;
  wire n539bar;
  wire n540bar;
  wire n541bar;
  wire n542bar;
  wire n543bar;
  wire n544bar;
  wire n545bar;
  wire n546bar;
  wire n547bar;
  wire n548bar;
  wire n549bar;
  wire n550bar;
  wire n551bar;
  wire n552bar;
  wire n553bar;
  wire n554bar;
  wire n555bar;
  wire n556bar;
  wire n557bar;
  wire n558bar;
  wire n559bar;
  wire n560bar;
  wire n561bar;
  wire n562bar;
  wire n563bar;
  wire n564bar;
  wire n565bar;
  wire n566bar;
  wire n567bar;
  wire n568bar;
  wire n569bar;
  wire n570bar;
  wire n571bar;
  wire n572bar;
  wire n573bar;
  wire n574bar;
  wire n575bar;
  wire n576bar;
  wire n577bar;
  wire n578bar;
  wire n579bar;
  wire n580bar;
  wire n581bar;
  wire n582bar;
  wire n583bar;
  wire n584bar;
  wire n585bar;
  wire n586bar;
  wire n587bar;
  wire n588bar;
  wire n589bar;
  wire n590bar;
  wire n591bar;
  wire n592bar;
  wire n593bar;
  wire n594bar;
  wire n595bar;
  wire n596bar;
  wire n597bar;
  wire n598bar;
  wire n599bar;
  wire n600bar;
  wire n601bar;
  wire n602bar;
  wire n603bar;
  wire n604bar;
  wire n605bar;
  wire n606bar;
  wire n607bar;
  wire n608bar;
  wire n609bar;
  wire n610bar;
  wire n611bar;
  wire n612bar;
  wire n613bar;
  wire n614bar;
  wire n615bar;
  wire n616bar;
  wire n617bar;
  wire n618bar;
  wire n619bar;
  wire n620bar;
  wire n621bar;
  wire n622bar;
  wire n623bar;
  wire n624bar;
  wire n625bar;
  wire n626bar;
  wire n627bar;
  wire n628bar;
  wire n629bar;
  wire n630bar;
  wire n631bar;
  wire n632bar;
  wire n633bar;
  wire n634bar;
  wire n635bar;
  wire n636bar;
  wire n637bar;
  wire n638bar;
  wire n639bar;
  wire n640bar;
  wire n641bar;
  wire n642bar;
  wire n643bar;
  wire n644bar;
  wire n645bar;
  wire n646bar;
  wire n647bar;
  wire n648bar;
  wire n649bar;
  wire n650bar;
  wire n651bar;
  wire n652bar;
  wire n653bar;
  wire n654bar;
  wire n655bar;
  wire n656bar;
  wire n657bar;
  wire n658bar;
  wire n659bar;
  wire n660bar;
  wire n661bar;
  wire n662bar;
  wire n663bar;
  wire n664bar;
  wire n665bar;
  wire n666bar;
  wire n667bar;
  wire n668bar;
  wire n669bar;
  wire n670bar;
  wire n671bar;
  wire n672bar;
  wire n673bar;
  wire n674bar;
  wire n675bar;
  wire n676bar;
  wire n677bar;
  wire n678bar;
  wire n679bar;
  wire n680bar;
  wire n681bar;
  wire n682bar;
  wire n683bar;
  wire n684bar;
  wire n685bar;
  wire n686bar;
  wire n687bar;
  wire n688bar;
  wire n689bar;
  wire n690bar;
  wire n691bar;
  wire n692bar;
  wire n693bar;
  wire n694bar;
  wire n695bar;
  wire n696bar;
  wire n697bar;
  wire n698bar;
  wire n699bar;
  wire n700bar;
  wire n701bar;
  wire n702bar;
  wire n703bar;
  wire n704bar;
  wire n705bar;
  wire n706bar;
  wire n707bar;
  wire n708bar;
  wire n709bar;
  wire n710bar;
  wire n711bar;
  wire n712bar;
  wire n713bar;
  wire n714bar;
  wire n715bar;
  wire n716bar;
  wire n717bar;
  wire n718bar;
  wire n719bar;
  wire n720bar;
  wire n721bar;
  wire n722bar;
  wire n723bar;
  wire n724bar;
  wire n725bar;
  wire n726bar;
  wire n727bar;
  wire n728bar;
  wire n729bar;
  wire n730bar;
  wire n731bar;
  wire n732bar;
  wire n733bar;
  wire n734bar;
  wire n735bar;
  wire n736bar;
  wire n737bar;
  wire n738bar;
  wire n739bar;
  wire n740bar;
  wire n741bar;
  wire n742bar;
  wire n743bar;
  wire n744bar;
  wire n745bar;
  wire n746bar;
  wire n747bar;
  wire n748bar;
  wire n749bar;
  wire n750bar;
  wire n751bar;
  wire n752bar;
  wire n753bar;
  wire n754bar;
  wire n755bar;
  wire n756bar;
  wire n757bar;
  wire n758bar;
  wire n759bar;
  wire n760bar;
  wire n761bar;
  wire n762bar;
  wire n763bar;
  wire n764bar;
  wire n765bar;
  wire n766bar;
  wire n767bar;
  wire n768bar;
  wire n769bar;
  wire n770bar;
  wire n771bar;
  wire n772bar;
  wire n773bar;
  wire n774bar;
  wire n775bar;
  wire n776bar;
  wire n777bar;
  wire n778bar;
  wire n779bar;
  wire n780bar;
  wire n781bar;
  wire n782bar;
  wire n783bar;
  wire n784bar;
  wire n785bar;
  wire n786bar;
  wire n787bar;
  wire n788bar;
  wire n789bar;
  wire n790bar;
  wire n791bar;
  wire n792bar;
  wire n793bar;
  wire n794bar;
  wire n795bar;
  wire n796bar;
  wire n797bar;
  wire n798bar;
  wire n799bar;
  wire n800bar;
  wire n801bar;
  wire n802bar;
  wire n803bar;
  wire n804bar;
  wire n805bar;
  wire n806bar;
  wire n807bar;
  wire n808bar;
  wire n809bar;
  wire n810bar;
  wire n811bar;
  wire n812bar;
  wire n813bar;
  wire n814bar;
  wire n815bar;
  wire n816bar;
  wire n817bar;
  wire n818bar;
  wire n819bar;
  wire n820bar;
  wire n821bar;
  wire n822bar;
  wire n823bar;
  wire n824bar;
  wire n825bar;
  wire n826bar;
  wire n827bar;
  wire n828bar;
  wire n829bar;
  wire n830bar;
  wire n831bar;
  wire n832bar;
  wire n833bar;
  wire n834bar;
  wire n835bar;
  wire n836bar;
  wire n837bar;
  wire n838bar;
  wire n839bar;
  wire n840bar;
  wire n841bar;
  wire n842bar;
  wire n843bar;
  wire n844bar;
  wire n845bar;
  wire n846bar;
  wire n847bar;
  wire n848bar;
  wire n849bar;
  wire n850bar;
  wire n851bar;
  wire n852bar;
  wire n853bar;
  wire n854bar;
  wire n855bar;
  wire n856bar;
  wire n857bar;
  wire n858bar;
  wire n859bar;
  wire n860bar;
  wire n861bar;
  wire n862bar;
  wire n863bar;
  wire n864bar;
  wire n865bar;
  wire n866bar;
  wire n867bar;
  wire n868bar;
  wire n869bar;
  wire n870bar;
  wire n871bar;
  wire n872bar;
  wire n873bar;
  wire n874bar;
  wire n875bar;
  wire n876bar;
  wire n877bar;
  wire n878bar;
  wire n879bar;
  wire n880bar;
  wire n881bar;
  wire n882bar;
  wire n883bar;
  wire n884bar;
  wire n885bar;
  wire n886bar;
  wire n887bar;
  wire n888bar;
  wire n889bar;
  wire n890bar;
  wire n891bar;
  wire n892bar;
  wire n893bar;
  wire n894bar;
  wire n895bar;
  wire n896bar;
  wire n897bar;
  wire n898bar;
  wire n899bar;
  wire n900bar;
  wire n901bar;
  wire n902bar;
  wire n903bar;
  wire n904bar;
  wire n905bar;
  wire n906bar;
  wire n907bar;
  wire n908bar;
  wire n909bar;
  wire n910bar;
  wire n911bar;
  wire n912bar;
  wire n913bar;
  wire n914bar;
  wire n915bar;
  wire n916bar;
  wire n917bar;
  wire n918bar;
  wire n919bar;
  wire n920bar;
  wire n921bar;
  wire n922bar;
  wire n923bar;
  wire n924bar;
  wire n925bar;
  wire n926bar;
  wire n927bar;
  wire n928bar;
  wire n929bar;
  wire n930bar;
  wire n931bar;
  wire n932bar;
  wire n933bar;
  wire n934bar;
  wire n935bar;
  wire n936bar;
  wire n937bar;
  wire n938bar;
  wire n939bar;
  wire n940bar;
  wire n941bar;
  wire n942bar;
  wire n943bar;
  wire n944bar;
  wire n945bar;
  wire n946bar;
  wire n947bar;
  wire n948bar;
  wire n949bar;
  wire n950bar;
  wire n951bar;
  wire n952bar;
  wire n953bar;
  wire n954bar;
  wire n955bar;
  wire n956bar;
  wire n957bar;
  wire n958bar;
  wire n959bar;
  wire n960bar;
  wire n961bar;
  wire n962bar;
  wire n963bar;
  wire n964bar;
  wire n965bar;
  wire n966bar;
  wire n967bar;
  wire n968bar;
  wire n969bar;
  wire n970bar;
  wire n971bar;
  wire n972bar;
//wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];
  //OR U1
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1 (
    .O(out[7]),
    .I0(n972),
    .I1(n971)
  );
  //AND U1bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1bar (
    .O(outbar[7]),
    .I0(n972bar),
    .I1(n971bar)
  );
  //OR U2
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2 (
    .O(n971),
    .I0(n970),
    .I1(n969)
  );
  //AND U2bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2bar (
    .O(n971bar),
    .I0(n970bar),
    .I1(n969bar)
  );
  //OR U3
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3 (
    .O(n969),
    .I0(n968),
    .I1(n967)
  );
  //AND U3bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3bar (
    .O(n969bar),
    .I0(n968bar),
    .I1(n967bar)
  );
  //OR U4
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4 (
    .O(n967),
    .I0(n966),
    .I1(n965)
  );
  //AND U4bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4bar (
    .O(n967bar),
    .I0(n966bar),
    .I1(n965bar)
  );
  //OR U5
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5 (
    .O(n968),
    .I0(n964),
    .I1(n963)
  );
  //AND U5bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5bar (
    .O(n968bar),
    .I0(n964bar),
    .I1(n963bar)
  );
  //OR U6
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6 (
    .O(n963),
    .I0(in[116]),
    .I1(n962)
  );
  //AND U6bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6bar (
    .O(n963bar),
    .I0(inbar[116]),
    .I1(n962bar)
  );
  //OR U7
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7 (
    .O(n970),
    .I0(n961),
    .I1(n960)
  );
  //AND U7bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7bar (
    .O(n970bar),
    .I0(n961bar),
    .I1(n960bar)
  );
  //OR U8
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8 (
    .O(n960),
    .I0(in[150]),
    .I1(in[127])
  );
  //AND U8bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8bar (
    .O(n960bar),
    .I0(inbar[150]),
    .I1(inbar[127])
  );
  //OR U9
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9 (
    .O(n961),
    .I0(in[160]),
    .I1(n959)
  );
  //AND U9bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9bar (
    .O(n961bar),
    .I0(inbar[160]),
    .I1(n959bar)
  );
  //OR U10
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10 (
    .O(n959),
    .I0(in[252]),
    .I1(in[168])
  );
  //AND U10bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10bar (
    .O(n959bar),
    .I0(inbar[252]),
    .I1(inbar[168])
  );
  //OR U11
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11 (
    .O(n972),
    .I0(n958),
    .I1(n957)
  );
  //AND U11bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11bar (
    .O(n972bar),
    .I0(n958bar),
    .I1(n957bar)
  );
  //OR U12
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12 (
    .O(n957),
    .I0(n956),
    .I1(n955)
  );
  //AND U12bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12bar (
    .O(n957bar),
    .I0(n956bar),
    .I1(n955bar)
  );
  //OR U13
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13 (
    .O(n955),
    .I0(in_17),
    .I1(in[96])
  );
  //AND U13bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13bar (
    .O(n955bar),
    .I0(in_17bar),
    .I1(inbar[96])
  );
  //OR U14
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14 (
    .O(n956),
    .I0(in_23),
    .I1(n954)
  );
  //AND U14bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14bar (
    .O(n956bar),
    .I0(in_23bar),
    .I1(n954bar)
  );
  //OR U15
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15 (
    .O(n954),
    .I0(in_31),
    .I1(in_26)
  );
  //AND U15bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15bar (
    .O(n954bar),
    .I0(in_31bar),
    .I1(in_26bar)
  );
  //OR U16
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16 (
    .O(n958),
    .I0(n953),
    .I1(n952)
  );
  //AND U16bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16bar (
    .O(n958bar),
    .I0(n953bar),
    .I1(n952bar)
  );
  //OR U17
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U17 (
    .O(n952),
    .I0(in_58),
    .I1(in_4)
  );
  //AND U17bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U17bar (
    .O(n952bar),
    .I0(in_58bar),
    .I1(in_4bar)
  );
  //OR U18
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U18 (
    .O(n953),
    .I0(in_59),
    .I1(n951)
  );
  //AND U18bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U18bar (
    .O(n953bar),
    .I0(in_59bar),
    .I1(n951bar)
  );
  //OR U19
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U19 (
    .O(n951),
    .I0(in_71),
    .I1(in_62)
  );
  //AND U19bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U19bar (
    .O(n951bar),
    .I0(in_71bar),
    .I1(in_62bar)
  );
  //OR U20
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U20 (
    .O(out[6]),
    .I0(n950),
    .I1(n949)
  );
  //AND U20bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U20bar (
    .O(outbar[6]),
    .I0(n950bar),
    .I1(n949bar)
  );
  //OR U21
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U21 (
    .O(n949),
    .I0(n948),
    .I1(n947)
  );
  //AND U21bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U21bar (
    .O(n949bar),
    .I0(n948bar),
    .I1(n947bar)
  );
  //OR U22
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U22 (
    .O(n947),
    .I0(n946),
    .I1(n945)
  );
  //AND U22bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U22bar (
    .O(n947bar),
    .I0(n946bar),
    .I1(n945bar)
  );
  //OR U23
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U23 (
    .O(n945),
    .I0(n944),
    .I1(n943)
  );
  //AND U23bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U23bar (
    .O(n945bar),
    .I0(n944bar),
    .I1(n943bar)
  );
  //OR U24
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U24 (
    .O(n946),
    .I0(n942),
    .I1(n941)
  );
  //AND U24bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U24bar (
    .O(n946bar),
    .I0(n942bar),
    .I1(n941bar)
  );
  //OR U25
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U25 (
    .O(n941),
    .I0(in[101]),
    .I1(n940)
  );
  //AND U25bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U25bar (
    .O(n941bar),
    .I0(inbar[101]),
    .I1(n940bar)
  );
  //OR U26
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U26 (
    .O(n948),
    .I0(n939),
    .I1(n938)
  );
  //AND U26bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U26bar (
    .O(n948bar),
    .I0(n939bar),
    .I1(n938bar)
  );
  //OR U27
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U27 (
    .O(n938),
    .I0(in[114]),
    .I1(in[104])
  );
  //AND U27bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U27bar (
    .O(n938bar),
    .I0(inbar[114]),
    .I1(inbar[104])
  );
  //OR U28
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U28 (
    .O(n939),
    .I0(in[128]),
    .I1(n937)
  );
  //AND U28bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U28bar (
    .O(n939bar),
    .I0(inbar[128]),
    .I1(n937bar)
  );
  //OR U29
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U29 (
    .O(n937),
    .I0(in[136]),
    .I1(in[134])
  );
  //AND U29bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U29bar (
    .O(n937bar),
    .I0(inbar[136]),
    .I1(inbar[134])
  );
  //OR U30
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U30 (
    .O(n950),
    .I0(n936),
    .I1(n935)
  );
  //AND U30bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U30bar (
    .O(n950bar),
    .I0(n936bar),
    .I1(n935bar)
  );
  //OR U31
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U31 (
    .O(n935),
    .I0(n934),
    .I1(n933)
  );
  //AND U31bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U31bar (
    .O(n935bar),
    .I0(n934bar),
    .I1(n933bar)
  );
  //OR U32
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U32 (
    .O(n933),
    .I0(in[177]),
    .I1(in[164])
  );
  //AND U32bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U32bar (
    .O(n933bar),
    .I0(inbar[177]),
    .I1(inbar[164])
  );
  //OR U33
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U33 (
    .O(n934),
    .I0(in[212]),
    .I1(n932)
  );
  //AND U33bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U33bar (
    .O(n934bar),
    .I0(inbar[212]),
    .I1(n932bar)
  );
  //OR U34
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U34 (
    .O(n932),
    .I0(in[248]),
    .I1(in[221])
  );
  //AND U34bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U34bar (
    .O(n932bar),
    .I0(inbar[248]),
    .I1(inbar[221])
  );
  //OR U35
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U35 (
    .O(n936),
    .I0(n931),
    .I1(n930)
  );
  //AND U35bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U35bar (
    .O(n936bar),
    .I0(n931bar),
    .I1(n930bar)
  );
  //OR U36
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U36 (
    .O(n930),
    .I0(in_18),
    .I1(in[93])
  );
  //AND U36bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U36bar (
    .O(n930bar),
    .I0(in_18bar),
    .I1(inbar[93])
  );
  //OR U37
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U37 (
    .O(n931),
    .I0(in_31),
    .I1(n929)
  );
  //AND U37bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U37bar (
    .O(n931bar),
    .I0(in_31bar),
    .I1(n929bar)
  );
  //OR U38
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U38 (
    .O(n929),
    .I0(in_7),
    .I1(in_39)
  );
  //AND U38bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U38bar (
    .O(n929bar),
    .I0(in_7bar),
    .I1(in_39bar)
  );
  //OR U39
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U39 (
    .O(out[5]),
    .I0(n928),
    .I1(n927)
  );
  //AND U39bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U39bar (
    .O(outbar[5]),
    .I0(n928bar),
    .I1(n927bar)
  );
  //OR U40
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U40 (
    .O(n927),
    .I0(n926),
    .I1(n925)
  );
  //AND U40bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U40bar (
    .O(n927bar),
    .I0(n926bar),
    .I1(n925bar)
  );
  //OR U41
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U41 (
    .O(n925),
    .I0(n924),
    .I1(n923)
  );
  //AND U41bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U41bar (
    .O(n925bar),
    .I0(n924bar),
    .I1(n923bar)
  );
  //OR U42
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U42 (
    .O(n923),
    .I0(n922),
    .I1(n921)
  );
  //AND U42bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U42bar (
    .O(n923bar),
    .I0(n922bar),
    .I1(n921bar)
  );
  //OR U43
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U43 (
    .O(n924),
    .I0(n940),
    .I1(n920)
  );
  //AND U43bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U43bar (
    .O(n924bar),
    .I0(n940bar),
    .I1(n920bar)
  );
  //OR U44
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U44 (
    .O(n920),
    .I0(in[111]),
    .I1(n919)
  );
  //AND U44bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U44bar (
    .O(n920bar),
    .I0(inbar[111]),
    .I1(n919bar)
  );
  //OR U45
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U45 (
    .O(n940),
    .I0(n918),
    .I1(n917)
  );
  //AND U45bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U45bar (
    .O(n940bar),
    .I0(n918bar),
    .I1(n917bar)
  );
  //OR U46
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U46 (
    .O(n917),
    .I0(n916),
    .I1(n915)
  );
  //AND U46bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U46bar (
    .O(n917bar),
    .I0(n916bar),
    .I1(n915bar)
  );
  //OR U47
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U47 (
    .O(n915),
    .I0(n914),
    .I1(n913)
  );
  //AND U47bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U47bar (
    .O(n915bar),
    .I0(n914bar),
    .I1(n913bar)
  );
  //OR U48
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U48 (
    .O(n913),
    .I0(in[140]),
    .I1(in[131])
  );
  //AND U48bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U48bar (
    .O(n913bar),
    .I0(inbar[140]),
    .I1(inbar[131])
  );
  //OR U49
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U49 (
    .O(n914),
    .I0(in[160]),
    .I1(in[144])
  );
  //AND U49bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U49bar (
    .O(n914bar),
    .I0(inbar[160]),
    .I1(inbar[144])
  );
  //OR U50
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U50 (
    .O(n916),
    .I0(n912),
    .I1(n911)
  );
  //AND U50bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U50bar (
    .O(n916bar),
    .I0(n912bar),
    .I1(n911bar)
  );
  //OR U51
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U51 (
    .O(n911),
    .I0(in[179]),
    .I1(in[174])
  );
  //AND U51bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U51bar (
    .O(n911bar),
    .I0(inbar[179]),
    .I1(inbar[174])
  );
  //OR U52
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U52 (
    .O(n912),
    .I0(in[188]),
    .I1(in[184])
  );
  //AND U52bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U52bar (
    .O(n912bar),
    .I0(inbar[188]),
    .I1(inbar[184])
  );
  //OR U53
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U53 (
    .O(n918),
    .I0(n910),
    .I1(n909)
  );
  //AND U53bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U53bar (
    .O(n918bar),
    .I0(n910bar),
    .I1(n909bar)
  );
  //OR U54
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U54 (
    .O(n909),
    .I0(n908),
    .I1(n907)
  );
  //AND U54bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U54bar (
    .O(n909bar),
    .I0(n908bar),
    .I1(n907bar)
  );
  //OR U55
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U55 (
    .O(n907),
    .I0(in[216]),
    .I1(in[200])
  );
  //AND U55bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U55bar (
    .O(n907bar),
    .I0(inbar[216]),
    .I1(inbar[200])
  );
  //OR U56
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U56 (
    .O(n908),
    .I0(in[228]),
    .I1(in[224])
  );
  //AND U56bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U56bar (
    .O(n908bar),
    .I0(inbar[228]),
    .I1(inbar[224])
  );
  //OR U57
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U57 (
    .O(n910),
    .I0(n906),
    .I1(n905)
  );
  //AND U57bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U57bar (
    .O(n910bar),
    .I0(n906bar),
    .I1(n905bar)
  );
  //OR U58
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U58 (
    .O(n905),
    .I0(in[247]),
    .I1(in[235])
  );
  //AND U58bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U58bar (
    .O(n905bar),
    .I0(inbar[247]),
    .I1(inbar[235])
  );
  //OR U59
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U59 (
    .O(n906),
    .I0(in_42),
    .I1(in[83])
  );
  //AND U59bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U59bar (
    .O(n906bar),
    .I0(in_42bar),
    .I1(inbar[83])
  );
  //OR U60
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U60 (
    .O(n926),
    .I0(n904),
    .I1(n903)
  );
  //AND U60bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U60bar (
    .O(n926bar),
    .I0(n904bar),
    .I1(n903bar)
  );
  //OR U61
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U61 (
    .O(n903),
    .I0(in[166]),
    .I1(in[123])
  );
  //AND U61bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U61bar (
    .O(n903bar),
    .I0(inbar[166]),
    .I1(inbar[123])
  );
  //OR U62
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U62 (
    .O(n904),
    .I0(in[170]),
    .I1(n902)
  );
  //AND U62bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U62bar (
    .O(n904bar),
    .I0(inbar[170]),
    .I1(n902bar)
  );
  //OR U63
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U63 (
    .O(n902),
    .I0(in[194]),
    .I1(in[183])
  );
  //AND U63bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U63bar (
    .O(n902bar),
    .I0(inbar[194]),
    .I1(inbar[183])
  );
  //OR U64
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U64 (
    .O(n928),
    .I0(n901),
    .I1(n900)
  );
  //AND U64bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U64bar (
    .O(n928bar),
    .I0(n901bar),
    .I1(n900bar)
  );
  //OR U65
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U65 (
    .O(n900),
    .I0(n899),
    .I1(n898)
  );
  //AND U65bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U65bar (
    .O(n900bar),
    .I0(n899bar),
    .I1(n898bar)
  );
  //OR U66
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U66 (
    .O(n898),
    .I0(in[241]),
    .I1(in[238])
  );
  //AND U66bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U66bar (
    .O(n898bar),
    .I0(inbar[241]),
    .I1(inbar[238])
  );
  //OR U67
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U67 (
    .O(n899),
    .I0(in[250]),
    .I1(n897)
  );
  //AND U67bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U67bar (
    .O(n899bar),
    .I0(inbar[250]),
    .I1(n897bar)
  );
  //OR U68
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U68 (
    .O(n897),
    .I0(in_24),
    .I1(in[84])
  );
  //AND U68bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U68bar (
    .O(n897bar),
    .I0(in_24bar),
    .I1(inbar[84])
  );
  //OR U69
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U69 (
    .O(n901),
    .I0(n896),
    .I1(n895)
  );
  //AND U69bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U69bar (
    .O(n901bar),
    .I0(n896bar),
    .I1(n895bar)
  );
  //OR U70
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U70 (
    .O(n895),
    .I0(in_41),
    .I1(in_29)
  );
  //AND U70bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U70bar (
    .O(n895bar),
    .I0(in_41bar),
    .I1(in_29bar)
  );
  //OR U71
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U71 (
    .O(n896),
    .I0(in_66),
    .I1(n894)
  );
  //AND U71bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U71bar (
    .O(n896bar),
    .I0(in_66bar),
    .I1(n894bar)
  );
  //OR U72
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U72 (
    .O(n894),
    .I0(in_76),
    .I1(in_71)
  );
  //AND U72bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U72bar (
    .O(n894bar),
    .I0(in_76bar),
    .I1(in_71bar)
  );
  //OR U73
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U73 (
    .O(out[4]),
    .I0(n893),
    .I1(n892)
  );
  //AND U73bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U73bar (
    .O(outbar[4]),
    .I0(n893bar),
    .I1(n892bar)
  );
  //OR U74
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U74 (
    .O(n892),
    .I0(n891),
    .I1(n890)
  );
  //AND U74bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U74bar (
    .O(n892bar),
    .I0(n891bar),
    .I1(n890bar)
  );
  //OR U75
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U75 (
    .O(n890),
    .I0(n889),
    .I1(n888)
  );
  //AND U75bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U75bar (
    .O(n890bar),
    .I0(n889bar),
    .I1(n888bar)
  );
  //OR U76
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U76 (
    .O(n888),
    .I0(n922),
    .I1(n887)
  );
  //AND U76bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U76bar (
    .O(n888bar),
    .I0(n922bar),
    .I1(n887bar)
  );
  //OR U77
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U77 (
    .O(n922),
    .I0(n886),
    .I1(n885)
  );
  //AND U77bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U77bar (
    .O(n922bar),
    .I0(n886bar),
    .I1(n885bar)
  );
  //OR U78
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U78 (
    .O(n885),
    .I0(n884),
    .I1(n883)
  );
  //AND U78bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U78bar (
    .O(n885bar),
    .I0(n884bar),
    .I1(n883bar)
  );
  //OR U79
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U79 (
    .O(n883),
    .I0(n882),
    .I1(n881)
  );
  //AND U79bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U79bar (
    .O(n883bar),
    .I0(n882bar),
    .I1(n881bar)
  );
  //OR U80
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U80 (
    .O(n881),
    .I0(in[118]),
    .I1(in[109])
  );
  //AND U80bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U80bar (
    .O(n881bar),
    .I0(inbar[118]),
    .I1(inbar[109])
  );
  //OR U81
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U81 (
    .O(n882),
    .I0(in[139]),
    .I1(in[120])
  );
  //AND U81bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U81bar (
    .O(n882bar),
    .I0(inbar[139]),
    .I1(inbar[120])
  );
  //OR U82
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U82 (
    .O(n884),
    .I0(n880),
    .I1(n879)
  );
  //AND U82bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U82bar (
    .O(n884bar),
    .I0(n880bar),
    .I1(n879bar)
  );
  //OR U83
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U83 (
    .O(n879),
    .I0(in[198]),
    .I1(in[154])
  );
  //AND U83bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U83bar (
    .O(n879bar),
    .I0(inbar[198]),
    .I1(inbar[154])
  );
  //OR U84
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U84 (
    .O(n880),
    .I0(in[210]),
    .I1(in[205])
  );
  //AND U84bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U84bar (
    .O(n880bar),
    .I0(inbar[210]),
    .I1(inbar[205])
  );
  //OR U85
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U85 (
    .O(n886),
    .I0(n878),
    .I1(n877)
  );
  //AND U85bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U85bar (
    .O(n886bar),
    .I0(n878bar),
    .I1(n877bar)
  );
  //OR U86
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U86 (
    .O(n877),
    .I0(n876),
    .I1(n875)
  );
  //AND U86bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U86bar (
    .O(n877bar),
    .I0(n876bar),
    .I1(n875bar)
  );
  //OR U87
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U87 (
    .O(n875),
    .I0(in[219]),
    .I1(in[217])
  );
  //AND U87bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U87bar (
    .O(n875bar),
    .I0(inbar[219]),
    .I1(inbar[217])
  );
  //OR U88
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U88 (
    .O(n876),
    .I0(in[86]),
    .I1(in[252])
  );
  //AND U88bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U88bar (
    .O(n876bar),
    .I0(inbar[86]),
    .I1(inbar[252])
  );
  //OR U89
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U89 (
    .O(n878),
    .I0(n874),
    .I1(n873)
  );
  //AND U89bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U89bar (
    .O(n878bar),
    .I0(n874bar),
    .I1(n873bar)
  );
  //OR U90
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U90 (
    .O(n873),
    .I0(in_40),
    .I1(in[91])
  );
  //AND U90bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U90bar (
    .O(n873bar),
    .I0(in_40bar),
    .I1(inbar[91])
  );
  //OR U91
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U91 (
    .O(n874),
    .I0(in_8),
    .I1(in_46)
  );
  //AND U91bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U91bar (
    .O(n874bar),
    .I0(in_8bar),
    .I1(in_46bar)
  );
  //OR U92
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U92 (
    .O(n889),
    .I0(n872),
    .I1(n871)
  );
  //AND U92bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U92bar (
    .O(n889bar),
    .I0(n872bar),
    .I1(n871bar)
  );
  //OR U93
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U93 (
    .O(n871),
    .I0(in[117]),
    .I1(n943)
  );
  //AND U93bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U93bar (
    .O(n871bar),
    .I0(inbar[117]),
    .I1(n943bar)
  );
  //OR U94
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U94 (
    .O(n943),
    .I0(n870),
    .I1(n869)
  );
  //AND U94bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U94bar (
    .O(n943bar),
    .I0(n870bar),
    .I1(n869bar)
  );
  //OR U95
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U95 (
    .O(n869),
    .I0(n868),
    .I1(n867)
  );
  //AND U95bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U95bar (
    .O(n869bar),
    .I0(n868bar),
    .I1(n867bar)
  );
  //OR U96
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U96 (
    .O(n867),
    .I0(n866),
    .I1(n865)
  );
  //AND U96bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U96bar (
    .O(n867bar),
    .I0(n866bar),
    .I1(n865bar)
  );
  //OR U97
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U97 (
    .O(n865),
    .I0(n864),
    .I1(n863)
  );
  //AND U97bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U97bar (
    .O(n865bar),
    .I0(n864bar),
    .I1(n863bar)
  );
  //OR U98
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U98 (
    .O(n866),
    .I0(in[108]),
    .I1(n919)
  );
  //AND U98bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U98bar (
    .O(n866bar),
    .I0(inbar[108]),
    .I1(n919bar)
  );
  //OR U99
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U99 (
    .O(n919),
    .I0(n862),
    .I1(n861)
  );
  //AND U99bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U99bar (
    .O(n919bar),
    .I0(n862bar),
    .I1(n861bar)
  );
  //OR U100
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U100 (
    .O(n861),
    .I0(n860),
    .I1(n859)
  );
  //AND U100bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U100bar (
    .O(n861bar),
    .I0(n860bar),
    .I1(n859bar)
  );
  //OR U101
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U101 (
    .O(n859),
    .I0(n858),
    .I1(n857)
  );
  //AND U101bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U101bar (
    .O(n859bar),
    .I0(n858bar),
    .I1(n857bar)
  );
  //OR U102
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U102 (
    .O(n857),
    .I0(in[119]),
    .I1(in[105])
  );
  //AND U102bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U102bar (
    .O(n857bar),
    .I0(inbar[119]),
    .I1(inbar[105])
  );
  //OR U103
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U103 (
    .O(n858),
    .I0(in[186]),
    .I1(in[175])
  );
  //AND U103bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U103bar (
    .O(n858bar),
    .I0(inbar[186]),
    .I1(inbar[175])
  );
  //OR U104
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U104 (
    .O(n860),
    .I0(n856),
    .I1(n855)
  );
  //AND U104bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U104bar (
    .O(n860bar),
    .I0(n856bar),
    .I1(n855bar)
  );
  //OR U105
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U105 (
    .O(n855),
    .I0(in[202]),
    .I1(in[193])
  );
  //AND U105bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U105bar (
    .O(n855bar),
    .I0(inbar[202]),
    .I1(inbar[193])
  );
  //OR U106
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U106 (
    .O(n856),
    .I0(in[225]),
    .I1(in[208])
  );
  //AND U106bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U106bar (
    .O(n856bar),
    .I0(inbar[225]),
    .I1(inbar[208])
  );
  //OR U107
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U107 (
    .O(n862),
    .I0(n854),
    .I1(n853)
  );
  //AND U107bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U107bar (
    .O(n862bar),
    .I0(n854bar),
    .I1(n853bar)
  );
  //OR U108
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U108 (
    .O(n853),
    .I0(n852),
    .I1(n851)
  );
  //AND U108bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U108bar (
    .O(n853bar),
    .I0(n852bar),
    .I1(n851bar)
  );
  //OR U109
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U109 (
    .O(n851),
    .I0(in_1),
    .I1(in[85])
  );
  //AND U109bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U109bar (
    .O(n851bar),
    .I0(in_1bar),
    .I1(inbar[85])
  );
  //OR U110
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U110 (
    .O(n852),
    .I0(in_23),
    .I1(in_19)
  );
  //AND U110bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U110bar (
    .O(n852bar),
    .I0(in_23bar),
    .I1(in_19bar)
  );
  //OR U111
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U111 (
    .O(n854),
    .I0(n850),
    .I1(n849)
  );
  //AND U111bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U111bar (
    .O(n854bar),
    .I0(n850bar),
    .I1(n849bar)
  );
  //OR U112
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U112 (
    .O(n849),
    .I0(in_43),
    .I1(in_33)
  );
  //AND U112bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U112bar (
    .O(n849bar),
    .I0(in_43bar),
    .I1(in_33bar)
  );
  //OR U113
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U113 (
    .O(n850),
    .I0(in_63),
    .I1(in_44)
  );
  //AND U113bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U113bar (
    .O(n850bar),
    .I0(in_63bar),
    .I1(in_44bar)
  );
  //OR U114
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U114 (
    .O(n868),
    .I0(n848),
    .I1(n847)
  );
  //AND U114bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U114bar (
    .O(n868bar),
    .I0(n848bar),
    .I1(n847bar)
  );
  //OR U115
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U115 (
    .O(n847),
    .I0(in[141]),
    .I1(in[112])
  );
  //AND U115bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U115bar (
    .O(n847bar),
    .I0(inbar[141]),
    .I1(inbar[112])
  );
  //OR U116
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U116 (
    .O(n848),
    .I0(in[147]),
    .I1(n846)
  );
  //AND U116bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U116bar (
    .O(n848bar),
    .I0(inbar[147]),
    .I1(n846bar)
  );
  //OR U117
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U117 (
    .O(n846),
    .I0(in[181]),
    .I1(in[167])
  );
  //AND U117bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U117bar (
    .O(n846bar),
    .I0(inbar[181]),
    .I1(inbar[167])
  );
  //OR U118
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U118 (
    .O(n870),
    .I0(n845),
    .I1(n844)
  );
  //AND U118bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U118bar (
    .O(n870bar),
    .I0(n845bar),
    .I1(n844bar)
  );
  //OR U119
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U119 (
    .O(n844),
    .I0(n843),
    .I1(n842)
  );
  //AND U119bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U119bar (
    .O(n844bar),
    .I0(n843bar),
    .I1(n842bar)
  );
  //OR U120
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U120 (
    .O(n842),
    .I0(in[229]),
    .I1(in[201])
  );
  //AND U120bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U120bar (
    .O(n842bar),
    .I0(inbar[229]),
    .I1(inbar[201])
  );
  //OR U121
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U121 (
    .O(n843),
    .I0(in[237]),
    .I1(n841)
  );
  //AND U121bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U121bar (
    .O(n843bar),
    .I0(inbar[237]),
    .I1(n841bar)
  );
  //OR U122
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U122 (
    .O(n841),
    .I0(in[94]),
    .I1(in[253])
  );
  //AND U122bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U122bar (
    .O(n841bar),
    .I0(inbar[94]),
    .I1(inbar[253])
  );
  //OR U123
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U123 (
    .O(n845),
    .I0(n840),
    .I1(n839)
  );
  //AND U123bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U123bar (
    .O(n845bar),
    .I0(n840bar),
    .I1(n839bar)
  );
  //OR U124
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U124 (
    .O(n839),
    .I0(in_21),
    .I1(in[96])
  );
  //AND U124bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U124bar (
    .O(n839bar),
    .I0(in_21bar),
    .I1(inbar[96])
  );
  //OR U125
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U125 (
    .O(n840),
    .I0(in_25),
    .I1(n838)
  );
  //AND U125bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U125bar (
    .O(n840bar),
    .I0(in_25bar),
    .I1(n838bar)
  );
  //OR U126
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U126 (
    .O(n838),
    .I0(in_81),
    .I1(in_45)
  );
  //AND U126bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U126bar (
    .O(n838bar),
    .I0(in_81bar),
    .I1(in_45bar)
  );
  //OR U127
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U127 (
    .O(n891),
    .I0(n837),
    .I1(n836)
  );
  //AND U127bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U127bar (
    .O(n891bar),
    .I0(n837bar),
    .I1(n836bar)
  );
  //OR U128
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U128 (
    .O(n836),
    .I0(in[142]),
    .I1(in[124])
  );
  //AND U128bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U128bar (
    .O(n836bar),
    .I0(inbar[142]),
    .I1(inbar[124])
  );
  //OR U129
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U129 (
    .O(n837),
    .I0(in[150]),
    .I1(n835)
  );
  //AND U129bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U129bar (
    .O(n837bar),
    .I0(inbar[150]),
    .I1(n835bar)
  );
  //OR U130
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U130 (
    .O(n835),
    .I0(in[172]),
    .I1(in[155])
  );
  //AND U130bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U130bar (
    .O(n835bar),
    .I0(inbar[172]),
    .I1(inbar[155])
  );
  //OR U131
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U131 (
    .O(n893),
    .I0(n834),
    .I1(n833)
  );
  //AND U131bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U131bar (
    .O(n893bar),
    .I0(n834bar),
    .I1(n833bar)
  );
  //OR U132
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U132 (
    .O(n833),
    .I0(n832),
    .I1(n831)
  );
  //AND U132bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U132bar (
    .O(n833bar),
    .I0(n832bar),
    .I1(n831bar)
  );
  //OR U133
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U133 (
    .O(n831),
    .I0(in[196]),
    .I1(in[173])
  );
  //AND U133bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U133bar (
    .O(n831bar),
    .I0(inbar[196]),
    .I1(inbar[173])
  );
  //OR U134
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U134 (
    .O(n832),
    .I0(in[222]),
    .I1(n830)
  );
  //AND U134bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U134bar (
    .O(n832bar),
    .I0(inbar[222]),
    .I1(n830bar)
  );
  //OR U135
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U135 (
    .O(n830),
    .I0(in[227]),
    .I1(in[226])
  );
  //AND U135bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U135bar (
    .O(n830bar),
    .I0(inbar[227]),
    .I1(inbar[226])
  );
  //OR U136
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U136 (
    .O(n834),
    .I0(n829),
    .I1(n828)
  );
  //AND U136bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U136bar (
    .O(n834bar),
    .I0(n829bar),
    .I1(n828bar)
  );
  //OR U137
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U137 (
    .O(n828),
    .I0(in[249]),
    .I1(in[231])
  );
  //AND U137bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U137bar (
    .O(n828bar),
    .I0(inbar[249]),
    .I1(inbar[231])
  );
  //OR U138
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U138 (
    .O(n829),
    .I0(in_28),
    .I1(n827)
  );
  //AND U138bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U138bar (
    .O(n829bar),
    .I0(in_28bar),
    .I1(n827bar)
  );
  //OR U139
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U139 (
    .O(n827),
    .I0(in_52),
    .I1(in_47)
  );
  //AND U139bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U139bar (
    .O(n827bar),
    .I0(in_52bar),
    .I1(in_47bar)
  );
  //OR U140
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U140 (
    .O(out[3]),
    .I0(n826),
    .I1(n825)
  );
  //AND U140bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U140bar (
    .O(outbar[3]),
    .I0(n826bar),
    .I1(n825bar)
  );
  //OR U141
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U141 (
    .O(n825),
    .I0(n824),
    .I1(n823)
  );
  //AND U141bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U141bar (
    .O(n825bar),
    .I0(n824bar),
    .I1(n823bar)
  );
  //OR U142
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U142 (
    .O(n823),
    .I0(n822),
    .I1(n821)
  );
  //AND U142bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U142bar (
    .O(n823bar),
    .I0(n822bar),
    .I1(n821bar)
  );
  //OR U143
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U143 (
    .O(n821),
    .I0(n820),
    .I1(n819)
  );
  //AND U143bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U143bar (
    .O(n821bar),
    .I0(n820bar),
    .I1(n819bar)
  );
  //OR U144
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U144 (
    .O(n822),
    .I0(n964),
    .I1(n818)
  );
  //AND U144bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U144bar (
    .O(n822bar),
    .I0(n964bar),
    .I1(n818bar)
  );
  //OR U145
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U145 (
    .O(n818),
    .I0(in[118]),
    .I1(n817)
  );
  //AND U145bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U145bar (
    .O(n818bar),
    .I0(inbar[118]),
    .I1(n817bar)
  );
  //OR U146
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U146 (
    .O(n964),
    .I0(n816),
    .I1(n815)
  );
  //AND U146bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U146bar (
    .O(n964bar),
    .I0(n816bar),
    .I1(n815bar)
  );
  //OR U147
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U147 (
    .O(n815),
    .I0(n814),
    .I1(n813)
  );
  //AND U147bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U147bar (
    .O(n815bar),
    .I0(n814bar),
    .I1(n813bar)
  );
  //OR U148
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U148 (
    .O(n813),
    .I0(n812),
    .I1(n811)
  );
  //AND U148bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U148bar (
    .O(n813bar),
    .I0(n812bar),
    .I1(n811bar)
  );
  //OR U149
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U149 (
    .O(n811),
    .I0(in[122]),
    .I1(in[111])
  );
  //AND U149bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U149bar (
    .O(n811bar),
    .I0(inbar[122]),
    .I1(inbar[111])
  );
  //OR U150
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U150 (
    .O(n812),
    .I0(in[154]),
    .I1(in[151])
  );
  //AND U150bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U150bar (
    .O(n812bar),
    .I0(inbar[154]),
    .I1(inbar[151])
  );
  //OR U151
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U151 (
    .O(n814),
    .I0(n810),
    .I1(n809)
  );
  //AND U151bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U151bar (
    .O(n814bar),
    .I0(n810bar),
    .I1(n809bar)
  );
  //OR U152
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U152 (
    .O(n809),
    .I0(in[187]),
    .I1(in[177])
  );
  //AND U152bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U152bar (
    .O(n809bar),
    .I0(inbar[187]),
    .I1(inbar[177])
  );
  //OR U153
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U153 (
    .O(n810),
    .I0(in[200]),
    .I1(in[192])
  );
  //AND U153bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U153bar (
    .O(n810bar),
    .I0(inbar[200]),
    .I1(inbar[192])
  );
  //OR U154
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U154 (
    .O(n816),
    .I0(n808),
    .I1(n807)
  );
  //AND U154bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U154bar (
    .O(n816bar),
    .I0(n808bar),
    .I1(n807bar)
  );
  //OR U155
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U155 (
    .O(n807),
    .I0(n806),
    .I1(n805)
  );
  //AND U155bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U155bar (
    .O(n807bar),
    .I0(n806bar),
    .I1(n805bar)
  );
  //OR U156
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U156 (
    .O(n805),
    .I0(in[225]),
    .I1(in[207])
  );
  //AND U156bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U156bar (
    .O(n805bar),
    .I0(inbar[225]),
    .I1(inbar[207])
  );
  //OR U157
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U157 (
    .O(n806),
    .I0(in[98]),
    .I1(in[226])
  );
  //AND U157bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U157bar (
    .O(n806bar),
    .I0(inbar[98]),
    .I1(inbar[226])
  );
  //OR U158
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U158 (
    .O(n808),
    .I0(n804),
    .I1(n803)
  );
  //AND U158bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U158bar (
    .O(n808bar),
    .I0(n804bar),
    .I1(n803bar)
  );
  //OR U159
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U159 (
    .O(n803),
    .I0(in_20),
    .I1(in_16)
  );
  //AND U159bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U159bar (
    .O(n803bar),
    .I0(in_20bar),
    .I1(in_16bar)
  );
  //OR U160
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U160 (
    .O(n804),
    .I0(in_55),
    .I1(in_45)
  );
  //AND U160bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U160bar (
    .O(n804bar),
    .I0(in_55bar),
    .I1(in_45bar)
  );
  //OR U161
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U161 (
    .O(n824),
    .I0(n802),
    .I1(n801)
  );
  //AND U161bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U161bar (
    .O(n824bar),
    .I0(n802bar),
    .I1(n801bar)
  );
  //OR U162
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U162 (
    .O(n801),
    .I0(in[162]),
    .I1(in[149])
  );
  //AND U162bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U162bar (
    .O(n801bar),
    .I0(inbar[162]),
    .I1(inbar[149])
  );
  //OR U163
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U163 (
    .O(n802),
    .I0(in[163]),
    .I1(n800)
  );
  //AND U163bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U163bar (
    .O(n802bar),
    .I0(inbar[163]),
    .I1(n800bar)
  );
  //OR U164
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U164 (
    .O(n800),
    .I0(in[191]),
    .I1(in[189])
  );
  //AND U164bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U164bar (
    .O(n800bar),
    .I0(inbar[191]),
    .I1(inbar[189])
  );
  //OR U165
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U165 (
    .O(n826),
    .I0(n799),
    .I1(n798)
  );
  //AND U165bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U165bar (
    .O(n826bar),
    .I0(n799bar),
    .I1(n798bar)
  );
  //OR U166
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U166 (
    .O(n798),
    .I0(n797),
    .I1(n796)
  );
  //AND U166bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U166bar (
    .O(n798bar),
    .I0(n797bar),
    .I1(n796bar)
  );
  //OR U167
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U167 (
    .O(n796),
    .I0(in[212]),
    .I1(in[193])
  );
  //AND U167bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U167bar (
    .O(n796bar),
    .I0(inbar[212]),
    .I1(inbar[193])
  );
  //OR U168
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U168 (
    .O(n797),
    .I0(in[238]),
    .I1(n795)
  );
  //AND U168bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U168bar (
    .O(n797bar),
    .I0(inbar[238]),
    .I1(n795bar)
  );
  //OR U169
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U169 (
    .O(n795),
    .I0(in[88]),
    .I1(in[247])
  );
  //AND U169bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U169bar (
    .O(n795bar),
    .I0(inbar[88]),
    .I1(inbar[247])
  );
  //OR U170
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U170 (
    .O(n799),
    .I0(n794),
    .I1(n793)
  );
  //AND U170bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U170bar (
    .O(n799bar),
    .I0(n794bar),
    .I1(n793bar)
  );
  //OR U171
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U171 (
    .O(n793),
    .I0(in[94]),
    .I1(in[92])
  );
  //AND U171bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U171bar (
    .O(n793bar),
    .I0(inbar[94]),
    .I1(inbar[92])
  );
  //OR U172
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U172 (
    .O(n794),
    .I0(in_52),
    .I1(n792)
  );
  //AND U172bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U172bar (
    .O(n794bar),
    .I0(in_52bar),
    .I1(n792bar)
  );
  //OR U173
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U173 (
    .O(n792),
    .I0(in_70),
    .I1(in_67)
  );
  //AND U173bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U173bar (
    .O(n792bar),
    .I0(in_70bar),
    .I1(in_67bar)
  );
  //OR U174
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U174 (
    .O(out[2]),
    .I0(n791),
    .I1(n790)
  );
  //AND U174bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U174bar (
    .O(outbar[2]),
    .I0(n791bar),
    .I1(n790bar)
  );
  //OR U175
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U175 (
    .O(n790),
    .I0(n789),
    .I1(n788)
  );
  //AND U175bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U175bar (
    .O(n790bar),
    .I0(n789bar),
    .I1(n788bar)
  );
  //OR U176
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U176 (
    .O(n788),
    .I0(n787),
    .I1(n786)
  );
  //AND U176bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U176bar (
    .O(n788bar),
    .I0(n787bar),
    .I1(n786bar)
  );
  //OR U177
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U177 (
    .O(n786),
    .I0(n819),
    .I1(n785)
  );
  //AND U177bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U177bar (
    .O(n786bar),
    .I0(n819bar),
    .I1(n785bar)
  );
  //OR U178
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U178 (
    .O(n819),
    .I0(n784),
    .I1(n783)
  );
  //AND U178bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U178bar (
    .O(n819bar),
    .I0(n784bar),
    .I1(n783bar)
  );
  //OR U179
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U179 (
    .O(n783),
    .I0(n782),
    .I1(n781)
  );
  //AND U179bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U179bar (
    .O(n783bar),
    .I0(n782bar),
    .I1(n781bar)
  );
  //OR U180
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U180 (
    .O(n781),
    .I0(n780),
    .I1(n779)
  );
  //AND U180bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U180bar (
    .O(n781bar),
    .I0(n780bar),
    .I1(n779bar)
  );
  //OR U181
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U181 (
    .O(n779),
    .I0(n962),
    .I1(n778)
  );
  //AND U181bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U181bar (
    .O(n779bar),
    .I0(n962bar),
    .I1(n778bar)
  );
  //OR U182
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U182 (
    .O(n962),
    .I0(n777),
    .I1(n776)
  );
  //AND U182bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U182bar (
    .O(n962bar),
    .I0(n777bar),
    .I1(n776bar)
  );
  //OR U183
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U183 (
    .O(n776),
    .I0(n775),
    .I1(n774)
  );
  //AND U183bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U183bar (
    .O(n776bar),
    .I0(n775bar),
    .I1(n774bar)
  );
  //OR U184
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U184 (
    .O(n774),
    .I0(n773),
    .I1(n772)
  );
  //AND U184bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U184bar (
    .O(n774bar),
    .I0(n773bar),
    .I1(n772bar)
  );
  //OR U185
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U185 (
    .O(n772),
    .I0(in[131]),
    .I1(in[120])
  );
  //AND U185bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U185bar (
    .O(n772bar),
    .I0(inbar[131]),
    .I1(inbar[120])
  );
  //OR U186
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U186 (
    .O(n773),
    .I0(in[153]),
    .I1(in[147])
  );
  //AND U186bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U186bar (
    .O(n773bar),
    .I0(inbar[153]),
    .I1(inbar[147])
  );
  //OR U187
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U187 (
    .O(n775),
    .I0(n771),
    .I1(n770)
  );
  //AND U187bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U187bar (
    .O(n775bar),
    .I0(n771bar),
    .I1(n770bar)
  );
  //OR U188
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U188 (
    .O(n770),
    .I0(in[170]),
    .I1(in[156])
  );
  //AND U188bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U188bar (
    .O(n770bar),
    .I0(inbar[170]),
    .I1(inbar[156])
  );
  //OR U189
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U189 (
    .O(n771),
    .I0(in[223]),
    .I1(in[190])
  );
  //AND U189bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U189bar (
    .O(n771bar),
    .I0(inbar[223]),
    .I1(inbar[190])
  );
  //OR U190
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U190 (
    .O(n777),
    .I0(n769),
    .I1(n768)
  );
  //AND U190bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U190bar (
    .O(n777bar),
    .I0(n769bar),
    .I1(n768bar)
  );
  //OR U191
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U191 (
    .O(n768),
    .I0(n767),
    .I1(n766)
  );
  //AND U191bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U191bar (
    .O(n768bar),
    .I0(n767bar),
    .I1(n766bar)
  );
  //OR U192
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U192 (
    .O(n766),
    .I0(in[236]),
    .I1(in[230])
  );
  //AND U192bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U192bar (
    .O(n766bar),
    .I0(inbar[236]),
    .I1(inbar[230])
  );
  //OR U193
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U193 (
    .O(n767),
    .I0(in[85]),
    .I1(in[240])
  );
  //AND U193bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U193bar (
    .O(n767bar),
    .I0(inbar[85]),
    .I1(inbar[240])
  );
  //OR U194
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U194 (
    .O(n769),
    .I0(n765),
    .I1(n764)
  );
  //AND U194bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U194bar (
    .O(n769bar),
    .I0(n765bar),
    .I1(n764bar)
  );
  //OR U195
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U195 (
    .O(n764),
    .I0(in_12),
    .I1(in[90])
  );
  //AND U195bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U195bar (
    .O(n764bar),
    .I0(in_12bar),
    .I1(inbar[90])
  );
  //OR U196
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U196 (
    .O(n765),
    .I0(in_39),
    .I1(in_28)
  );
  //AND U196bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U196bar (
    .O(n765bar),
    .I0(in_39bar),
    .I1(in_28bar)
  );
  //OR U197
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U197 (
    .O(n780),
    .I0(in[109]),
    .I1(n763)
  );
  //AND U197bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U197bar (
    .O(n780bar),
    .I0(inbar[109]),
    .I1(n763bar)
  );
  //OR U198
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U198 (
    .O(n782),
    .I0(n762),
    .I1(n761)
  );
  //AND U198bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U198bar (
    .O(n782bar),
    .I0(n762bar),
    .I1(n761bar)
  );
  //OR U199
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U199 (
    .O(n761),
    .I0(in[138]),
    .I1(in[129])
  );
  //AND U199bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U199bar (
    .O(n761bar),
    .I0(inbar[138]),
    .I1(inbar[129])
  );
  //OR U200
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U200 (
    .O(n762),
    .I0(in[157]),
    .I1(n760)
  );
  //AND U200bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U200bar (
    .O(n762bar),
    .I0(inbar[157]),
    .I1(n760bar)
  );
  //OR U201
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U201 (
    .O(n760),
    .I0(in[182]),
    .I1(in[167])
  );
  //AND U201bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U201bar (
    .O(n760bar),
    .I0(inbar[182]),
    .I1(inbar[167])
  );
  //OR U202
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U202 (
    .O(n784),
    .I0(n759),
    .I1(n758)
  );
  //AND U202bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U202bar (
    .O(n784bar),
    .I0(n759bar),
    .I1(n758bar)
  );
  //OR U203
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U203 (
    .O(n758),
    .I0(n757),
    .I1(n756)
  );
  //AND U203bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U203bar (
    .O(n758bar),
    .I0(n757bar),
    .I1(n756bar)
  );
  //OR U204
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U204 (
    .O(n756),
    .I0(in[195]),
    .I1(in[184])
  );
  //AND U204bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U204bar (
    .O(n756bar),
    .I0(inbar[195]),
    .I1(inbar[184])
  );
  //OR U205
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U205 (
    .O(n757),
    .I0(in[196]),
    .I1(n755)
  );
  //AND U205bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U205bar (
    .O(n757bar),
    .I0(inbar[196]),
    .I1(n755bar)
  );
  //OR U206
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U206 (
    .O(n755),
    .I0(in[215]),
    .I1(in[209])
  );
  //AND U206bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U206bar (
    .O(n755bar),
    .I0(inbar[215]),
    .I1(inbar[209])
  );
  //OR U207
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U207 (
    .O(n759),
    .I0(n754),
    .I1(n753)
  );
  //AND U207bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U207bar (
    .O(n759bar),
    .I0(n754bar),
    .I1(n753bar)
  );
  //OR U208
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U208 (
    .O(n753),
    .I0(in[93]),
    .I1(in[233])
  );
  //AND U208bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U208bar (
    .O(n753bar),
    .I0(inbar[93]),
    .I1(inbar[233])
  );
  //OR U209
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U209 (
    .O(n754),
    .I0(in_1),
    .I1(n752)
  );
  //AND U209bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U209bar (
    .O(n754bar),
    .I0(in_1bar),
    .I1(n752bar)
  );
  //OR U210
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U210 (
    .O(n752),
    .I0(in_69),
    .I1(in_66)
  );
  //AND U210bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U210bar (
    .O(n752bar),
    .I0(in_69bar),
    .I1(in_66bar)
  );
  //OR U211
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U211 (
    .O(n787),
    .I0(n966),
    .I1(n751)
  );
  //AND U211bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U211bar (
    .O(n787bar),
    .I0(n966bar),
    .I1(n751bar)
  );
  //OR U212
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U212 (
    .O(n751),
    .I0(in[134]),
    .I1(n750)
  );
  //AND U212bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U212bar (
    .O(n751bar),
    .I0(inbar[134]),
    .I1(n750bar)
  );
  //OR U213
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U213 (
    .O(n966),
    .I0(n749),
    .I1(n748)
  );
  //AND U213bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U213bar (
    .O(n966bar),
    .I0(n749bar),
    .I1(n748bar)
  );
  //OR U214
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U214 (
    .O(n748),
    .I0(n747),
    .I1(n746)
  );
  //AND U214bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U214bar (
    .O(n748bar),
    .I0(n747bar),
    .I1(n746bar)
  );
  //OR U215
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U215 (
    .O(n746),
    .I0(n745),
    .I1(n744)
  );
  //AND U215bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U215bar (
    .O(n746bar),
    .I0(n745bar),
    .I1(n744bar)
  );
  //OR U216
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U216 (
    .O(n744),
    .I0(in[136]),
    .I1(in[121])
  );
  //AND U216bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U216bar (
    .O(n744bar),
    .I0(inbar[136]),
    .I1(inbar[121])
  );
  //OR U217
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U217 (
    .O(n745),
    .I0(in[186]),
    .I1(in[174])
  );
  //AND U217bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U217bar (
    .O(n745bar),
    .I0(inbar[186]),
    .I1(inbar[174])
  );
  //OR U218
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U218 (
    .O(n747),
    .I0(n743),
    .I1(n742)
  );
  //AND U218bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U218bar (
    .O(n747bar),
    .I0(n743bar),
    .I1(n742bar)
  );
  //OR U219
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U219 (
    .O(n742),
    .I0(in[198]),
    .I1(in[197])
  );
  //AND U219bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U219bar (
    .O(n742bar),
    .I0(inbar[198]),
    .I1(inbar[197])
  );
  //OR U220
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U220 (
    .O(n743),
    .I0(in[214]),
    .I1(in[199])
  );
  //AND U220bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U220bar (
    .O(n743bar),
    .I0(inbar[214]),
    .I1(inbar[199])
  );
  //OR U221
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U221 (
    .O(n749),
    .I0(n741),
    .I1(n740)
  );
  //AND U221bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U221bar (
    .O(n749bar),
    .I0(n741bar),
    .I1(n740bar)
  );
  //OR U222
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U222 (
    .O(n740),
    .I0(n739),
    .I1(n738)
  );
  //AND U222bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U222bar (
    .O(n740bar),
    .I0(n739bar),
    .I1(n738bar)
  );
  //OR U223
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U223 (
    .O(n738),
    .I0(in[231]),
    .I1(in[220])
  );
  //AND U223bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U223bar (
    .O(n738bar),
    .I0(inbar[231]),
    .I1(inbar[220])
  );
  //OR U224
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U224 (
    .O(n739),
    .I0(in_25),
    .I1(in[245])
  );
  //AND U224bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U224bar (
    .O(n739bar),
    .I0(in_25bar),
    .I1(inbar[245])
  );
  //OR U225
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U225 (
    .O(n741),
    .I0(n737),
    .I1(n736)
  );
  //AND U225bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U225bar (
    .O(n741bar),
    .I0(n737bar),
    .I1(n736bar)
  );
  //OR U226
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U226 (
    .O(n736),
    .I0(in_53),
    .I1(in_29)
  );
  //AND U226bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U226bar (
    .O(n736bar),
    .I0(in_53bar),
    .I1(in_29bar)
  );
  //OR U227
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U227 (
    .O(n737),
    .I0(in_79),
    .I1(in_74)
  );
  //AND U227bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U227bar (
    .O(n737bar),
    .I0(in_79bar),
    .I1(in_74bar)
  );
  //OR U228
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U228 (
    .O(n789),
    .I0(n735),
    .I1(n734)
  );
  //AND U228bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U228bar (
    .O(n789bar),
    .I0(n735bar),
    .I1(n734bar)
  );
  //OR U229
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U229 (
    .O(n734),
    .I0(in[152]),
    .I1(in[140])
  );
  //AND U229bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U229bar (
    .O(n734bar),
    .I0(inbar[152]),
    .I1(inbar[140])
  );
  //OR U230
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U230 (
    .O(n735),
    .I0(in[155]),
    .I1(n733)
  );
  //AND U230bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U230bar (
    .O(n735bar),
    .I0(inbar[155]),
    .I1(n733bar)
  );
  //OR U231
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U231 (
    .O(n733),
    .I0(in[166]),
    .I1(in[165])
  );
  //AND U231bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U231bar (
    .O(n733bar),
    .I0(inbar[166]),
    .I1(inbar[165])
  );
  //OR U232
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U232 (
    .O(n791),
    .I0(n732),
    .I1(n731)
  );
  //AND U232bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U232bar (
    .O(n791bar),
    .I0(n732bar),
    .I1(n731bar)
  );
  //OR U233
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U233 (
    .O(n731),
    .I0(n730),
    .I1(n729)
  );
  //AND U233bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U233bar (
    .O(n731bar),
    .I0(n730bar),
    .I1(n729bar)
  );
  //OR U234
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U234 (
    .O(n729),
    .I0(in[202]),
    .I1(in[185])
  );
  //AND U234bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U234bar (
    .O(n729bar),
    .I0(inbar[202]),
    .I1(inbar[185])
  );
  //OR U235
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U235 (
    .O(n730),
    .I0(in[211]),
    .I1(n728)
  );
  //AND U235bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U235bar (
    .O(n730bar),
    .I0(inbar[211]),
    .I1(n728bar)
  );
  //OR U236
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U236 (
    .O(n728),
    .I0(in[255]),
    .I1(in[253])
  );
  //AND U236bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U236bar (
    .O(n728bar),
    .I0(inbar[255]),
    .I1(inbar[253])
  );
  //OR U237
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U237 (
    .O(n732),
    .I0(n727),
    .I1(n726)
  );
  //AND U237bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U237bar (
    .O(n732bar),
    .I0(n727bar),
    .I1(n726bar)
  );
  //OR U238
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U238 (
    .O(n726),
    .I0(in_35),
    .I1(in_15)
  );
  //AND U238bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U238bar (
    .O(n726bar),
    .I0(in_35bar),
    .I1(in_15bar)
  );
  //OR U239
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U239 (
    .O(n727),
    .I0(in_36),
    .I1(n725)
  );
  //AND U239bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U239bar (
    .O(n727bar),
    .I0(in_36bar),
    .I1(n725bar)
  );
  //OR U240
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U240 (
    .O(n725),
    .I0(in_48),
    .I1(in_40)
  );
  //AND U240bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U240bar (
    .O(n725bar),
    .I0(in_48bar),
    .I1(in_40bar)
  );
  //OR U241
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U241 (
    .O(out[1]),
    .I0(n724),
    .I1(n723)
  );
  //AND U241bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U241bar (
    .O(outbar[1]),
    .I0(n724bar),
    .I1(n723bar)
  );
  //OR U242
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U242 (
    .O(n723),
    .I0(n722),
    .I1(n721)
  );
  //AND U242bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U242bar (
    .O(n723bar),
    .I0(n722bar),
    .I1(n721bar)
  );
  //OR U243
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U243 (
    .O(n721),
    .I0(n720),
    .I1(n719)
  );
  //AND U243bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U243bar (
    .O(n721bar),
    .I0(n720bar),
    .I1(n719bar)
  );
  //OR U244
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U244 (
    .O(n719),
    .I0(n921),
    .I1(n887)
  );
  //AND U244bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U244bar (
    .O(n719bar),
    .I0(n921bar),
    .I1(n887bar)
  );
  //OR U245
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U245 (
    .O(n887),
    .I0(n718),
    .I1(n717)
  );
  //AND U245bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U245bar (
    .O(n887bar),
    .I0(n718bar),
    .I1(n717bar)
  );
  //OR U246
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U246 (
    .O(n717),
    .I0(n716),
    .I1(n715)
  );
  //AND U246bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U246bar (
    .O(n717bar),
    .I0(n716bar),
    .I1(n715bar)
  );
  //OR U247
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U247 (
    .O(n715),
    .I0(n714),
    .I1(n713)
  );
  //AND U247bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U247bar (
    .O(n715bar),
    .I0(n714bar),
    .I1(n713bar)
  );
  //OR U248
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U248 (
    .O(n713),
    .I0(in[116]),
    .I1(in[110])
  );
  //AND U248bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U248bar (
    .O(n713bar),
    .I0(inbar[116]),
    .I1(inbar[110])
  );
  //OR U249
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U249 (
    .O(n714),
    .I0(in[133]),
    .I1(in[130])
  );
  //AND U249bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U249bar (
    .O(n714bar),
    .I0(inbar[133]),
    .I1(inbar[130])
  );
  //OR U250
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U250 (
    .O(n716),
    .I0(n712),
    .I1(n711)
  );
  //AND U250bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U250bar (
    .O(n716bar),
    .I0(n712bar),
    .I1(n711bar)
  );
  //OR U251
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U251 (
    .O(n711),
    .I0(in[203]),
    .I1(in[135])
  );
  //AND U251bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U251bar (
    .O(n711bar),
    .I0(inbar[203]),
    .I1(inbar[135])
  );
  //OR U252
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U252 (
    .O(n712),
    .I0(in[232]),
    .I1(in[223])
  );
  //AND U252bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U252bar (
    .O(n712bar),
    .I0(inbar[232]),
    .I1(inbar[223])
  );
  //OR U253
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U253 (
    .O(n718),
    .I0(n710),
    .I1(n709)
  );
  //AND U253bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U253bar (
    .O(n718bar),
    .I0(n710bar),
    .I1(n709bar)
  );
  //OR U254
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U254 (
    .O(n709),
    .I0(n708),
    .I1(n707)
  );
  //AND U254bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U254bar (
    .O(n709bar),
    .I0(n708bar),
    .I1(n707bar)
  );
  //OR U255
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U255 (
    .O(n707),
    .I0(in[255]),
    .I1(in[233])
  );
  //AND U255bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U255bar (
    .O(n707bar),
    .I0(inbar[255]),
    .I1(inbar[233])
  );
  //OR U256
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U256 (
    .O(n708),
    .I0(in_53),
    .I1(in_34)
  );
  //AND U256bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U256bar (
    .O(n708bar),
    .I0(in_53bar),
    .I1(in_34bar)
  );
  //OR U257
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U257 (
    .O(n710),
    .I0(n706),
    .I1(n705)
  );
  //AND U257bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U257bar (
    .O(n710bar),
    .I0(n706bar),
    .I1(n705bar)
  );
  //OR U258
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U258 (
    .O(n705),
    .I0(in_57),
    .I1(in_55)
  );
  //AND U258bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U258bar (
    .O(n705bar),
    .I0(in_57bar),
    .I1(in_55bar)
  );
  //OR U259
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U259 (
    .O(n706),
    .I0(in_68),
    .I1(in_67)
  );
  //AND U259bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U259bar (
    .O(n706bar),
    .I0(in_68bar),
    .I1(in_67bar)
  );
  //OR U260
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U260 (
    .O(n921),
    .I0(n704),
    .I1(n703)
  );
  //AND U260bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U260bar (
    .O(n921bar),
    .I0(n704bar),
    .I1(n703bar)
  );
  //OR U261
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U261 (
    .O(n703),
    .I0(n702),
    .I1(n701)
  );
  //AND U261bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U261bar (
    .O(n703bar),
    .I0(n702bar),
    .I1(n701bar)
  );
  //OR U262
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U262 (
    .O(n701),
    .I0(n700),
    .I1(n699)
  );
  //AND U262bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U262bar (
    .O(n701bar),
    .I0(n700bar),
    .I1(n699bar)
  );
  //OR U263
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U263 (
    .O(n699),
    .I0(n944),
    .I1(n872)
  );
  //AND U263bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U263bar (
    .O(n699bar),
    .I0(n944bar),
    .I1(n872bar)
  );
  //OR U264
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U264 (
    .O(n872),
    .I0(n698),
    .I1(n697)
  );
  //AND U264bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U264bar (
    .O(n872bar),
    .I0(n698bar),
    .I1(n697bar)
  );
  //OR U265
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U265 (
    .O(n697),
    .I0(n696),
    .I1(n695)
  );
  //AND U265bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U265bar (
    .O(n697bar),
    .I0(n696bar),
    .I1(n695bar)
  );
  //OR U266
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U266 (
    .O(n695),
    .I0(n694),
    .I1(n693)
  );
  //AND U266bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U266bar (
    .O(n695bar),
    .I0(n694bar),
    .I1(n693bar)
  );
  //OR U267
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U267 (
    .O(n693),
    .I0(in[121]),
    .I1(in[102])
  );
  //AND U267bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U267bar (
    .O(n693bar),
    .I0(inbar[121]),
    .I1(inbar[102])
  );
  //OR U268
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U268 (
    .O(n694),
    .I0(in[162]),
    .I1(in[161])
  );
  //AND U268bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U268bar (
    .O(n694bar),
    .I0(inbar[162]),
    .I1(inbar[161])
  );
  //OR U269
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U269 (
    .O(n696),
    .I0(n692),
    .I1(n691)
  );
  //AND U269bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U269bar (
    .O(n696bar),
    .I0(n692bar),
    .I1(n691bar)
  );
  //OR U270
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U270 (
    .O(n691),
    .I0(in[192]),
    .I1(in[178])
  );
  //AND U270bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U270bar (
    .O(n691bar),
    .I0(inbar[192]),
    .I1(inbar[178])
  );
  //OR U271
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U271 (
    .O(n692),
    .I0(in[244]),
    .I1(in[209])
  );
  //AND U271bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U271bar (
    .O(n692bar),
    .I0(inbar[244]),
    .I1(inbar[209])
  );
  //OR U272
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U272 (
    .O(n698),
    .I0(n690),
    .I1(n689)
  );
  //AND U272bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U272bar (
    .O(n698bar),
    .I0(n690bar),
    .I1(n689bar)
  );
  //OR U273
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U273 (
    .O(n689),
    .I0(n688),
    .I1(n687)
  );
  //AND U273bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U273bar (
    .O(n689bar),
    .I0(n688bar),
    .I1(n687bar)
  );
  //OR U274
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U274 (
    .O(n687),
    .I0(in[90]),
    .I1(in[254])
  );
  //AND U274bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U274bar (
    .O(n687bar),
    .I0(inbar[90]),
    .I1(inbar[254])
  );
  //OR U275
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U275 (
    .O(n688),
    .I0(in_36),
    .I1(in_32)
  );
  //AND U275bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U275bar (
    .O(n688bar),
    .I0(in_36bar),
    .I1(in_32bar)
  );
  //OR U276
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U276 (
    .O(n690),
    .I0(n686),
    .I1(n685)
  );
  //AND U276bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U276bar (
    .O(n690bar),
    .I0(n686bar),
    .I1(n685bar)
  );
  //OR U277
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U277 (
    .O(n685),
    .I0(in_62),
    .I1(in_37)
  );
  //AND U277bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U277bar (
    .O(n685bar),
    .I0(in_62bar),
    .I1(in_37bar)
  );
  //OR U278
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U278 (
    .O(n686),
    .I0(in_75),
    .I1(in_73)
  );
  //AND U278bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U278bar (
    .O(n686bar),
    .I0(in_75bar),
    .I1(in_73bar)
  );
  //OR U279
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U279 (
    .O(n944),
    .I0(n684),
    .I1(n683)
  );
  //AND U279bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U279bar (
    .O(n944bar),
    .I0(n684bar),
    .I1(n683bar)
  );
  //OR U280
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U280 (
    .O(n683),
    .I0(n682),
    .I1(n681)
  );
  //AND U280bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U280bar (
    .O(n683bar),
    .I0(n682bar),
    .I1(n681bar)
  );
  //OR U281
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U281 (
    .O(n681),
    .I0(n680),
    .I1(n679)
  );
  //AND U281bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U281bar (
    .O(n681bar),
    .I0(n680bar),
    .I1(n679bar)
  );
  //OR U282
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U282 (
    .O(n679),
    .I0(in[171]),
    .I1(in[153])
  );
  //AND U282bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U282bar (
    .O(n679bar),
    .I0(inbar[171]),
    .I1(inbar[153])
  );
  //OR U283
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U283 (
    .O(n680),
    .I0(in[187]),
    .I1(in[176])
  );
  //AND U283bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U283bar (
    .O(n680bar),
    .I0(inbar[187]),
    .I1(inbar[176])
  );
  //OR U284
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U284 (
    .O(n682),
    .I0(n678),
    .I1(n677)
  );
  //AND U284bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U284bar (
    .O(n682bar),
    .I0(n678bar),
    .I1(n677bar)
  );
  //OR U285
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U285 (
    .O(n677),
    .I0(in[245]),
    .I1(in[211])
  );
  //AND U285bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U285bar (
    .O(n677bar),
    .I0(inbar[245]),
    .I1(inbar[211])
  );
  //OR U286
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U286 (
    .O(n678),
    .I0(in[97]),
    .I1(in[88])
  );
  //AND U286bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U286bar (
    .O(n678bar),
    .I0(inbar[97]),
    .I1(inbar[88])
  );
  //OR U287
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U287 (
    .O(n684),
    .I0(n676),
    .I1(n675)
  );
  //AND U287bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U287bar (
    .O(n684bar),
    .I0(n676bar),
    .I1(n675bar)
  );
  //OR U288
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U288 (
    .O(n675),
    .I0(n674),
    .I1(n673)
  );
  //AND U288bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U288bar (
    .O(n675bar),
    .I0(n674bar),
    .I1(n673bar)
  );
  //OR U289
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U289 (
    .O(n673),
    .I0(in_10),
    .I1(in_0)
  );
  //AND U289bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U289bar (
    .O(n673bar),
    .I0(in_10bar),
    .I1(in_0bar)
  );
  //OR U290
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U290 (
    .O(n674),
    .I0(in_59),
    .I1(in_5)
  );
  //AND U290bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U290bar (
    .O(n674bar),
    .I0(in_59bar),
    .I1(in_5bar)
  );
  //OR U291
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U291 (
    .O(n676),
    .I0(n672),
    .I1(n671)
  );
  //AND U291bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U291bar (
    .O(n676bar),
    .I0(n672bar),
    .I1(n671bar)
  );
  //OR U292
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U292 (
    .O(n671),
    .I0(in_60),
    .I1(in_6)
  );
  //AND U292bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U292bar (
    .O(n671bar),
    .I0(in_60bar),
    .I1(in_6bar)
  );
  //OR U293
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U293 (
    .O(n672),
    .I0(in_77),
    .I1(in_69)
  );
  //AND U293bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U293bar (
    .O(n672bar),
    .I0(in_77bar),
    .I1(in_69bar)
  );
  //OR U294
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U294 (
    .O(n700),
    .I0(in[113]),
    .I1(n864)
  );
  //AND U294bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U294bar (
    .O(n700bar),
    .I0(inbar[113]),
    .I1(n864bar)
  );
  //OR U295
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U295 (
    .O(n864),
    .I0(n670),
    .I1(n669)
  );
  //AND U295bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U295bar (
    .O(n864bar),
    .I0(n670bar),
    .I1(n669bar)
  );
  //OR U296
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U296 (
    .O(n669),
    .I0(n668),
    .I1(n667)
  );
  //AND U296bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U296bar (
    .O(n669bar),
    .I0(n668bar),
    .I1(n667bar)
  );
  //OR U297
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U297 (
    .O(n667),
    .I0(n666),
    .I1(n665)
  );
  //AND U297bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U297bar (
    .O(n667bar),
    .I0(n666bar),
    .I1(n665bar)
  );
  //OR U298
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U298 (
    .O(n665),
    .I0(in[125]),
    .I1(in[107])
  );
  //AND U298bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U298bar (
    .O(n665bar),
    .I0(inbar[125]),
    .I1(inbar[107])
  );
  //OR U299
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U299 (
    .O(n666),
    .I0(in[138]),
    .I1(in[126])
  );
  //AND U299bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U299bar (
    .O(n666bar),
    .I0(inbar[138]),
    .I1(inbar[126])
  );
  //OR U300
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U300 (
    .O(n668),
    .I0(n664),
    .I1(n663)
  );
  //AND U300bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U300bar (
    .O(n668bar),
    .I0(n664bar),
    .I1(n663bar)
  );
  //OR U301
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U301 (
    .O(n663),
    .I0(in[189]),
    .I1(in[143])
  );
  //AND U301bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U301bar (
    .O(n663bar),
    .I0(inbar[189]),
    .I1(inbar[143])
  );
  //OR U302
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U302 (
    .O(n664),
    .I0(in[99]),
    .I1(in[214])
  );
  //AND U302bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U302bar (
    .O(n664bar),
    .I0(inbar[99]),
    .I1(inbar[214])
  );
  //OR U303
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U303 (
    .O(n670),
    .I0(n662),
    .I1(n661)
  );
  //AND U303bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U303bar (
    .O(n670bar),
    .I0(n662bar),
    .I1(n661bar)
  );
  //OR U304
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U304 (
    .O(n661),
    .I0(n660),
    .I1(n659)
  );
  //AND U304bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U304bar (
    .O(n661bar),
    .I0(n660bar),
    .I1(n659bar)
  );
  //OR U305
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U305 (
    .O(n659),
    .I0(in_15),
    .I1(in_12)
  );
  //AND U305bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U305bar (
    .O(n659bar),
    .I0(in_15bar),
    .I1(in_12bar)
  );
  //OR U306
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U306 (
    .O(n660),
    .I0(in_20),
    .I1(in_2)
  );
  //AND U306bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U306bar (
    .O(n660bar),
    .I0(in_20bar),
    .I1(in_2bar)
  );
  //OR U307
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U307 (
    .O(n662),
    .I0(n658),
    .I1(n657)
  );
  //AND U307bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U307bar (
    .O(n662bar),
    .I0(n658bar),
    .I1(n657bar)
  );
  //OR U308
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U308 (
    .O(n657),
    .I0(in_30),
    .I1(in_3)
  );
  //AND U308bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U308bar (
    .O(n657bar),
    .I0(in_30bar),
    .I1(in_3bar)
  );
  //OR U309
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U309 (
    .O(n658),
    .I0(in_4),
    .I1(in_38)
  );
  //AND U309bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U309bar (
    .O(n658bar),
    .I0(in_4bar),
    .I1(in_38bar)
  );
  //OR U310
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U310 (
    .O(n702),
    .I0(n656),
    .I1(n655)
  );
  //AND U310bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U310bar (
    .O(n702bar),
    .I0(n656bar),
    .I1(n655bar)
  );
  //OR U311
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U311 (
    .O(n655),
    .I0(in[148]),
    .I1(in[137])
  );
  //AND U311bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U311bar (
    .O(n655bar),
    .I0(inbar[148]),
    .I1(inbar[137])
  );
  //OR U312
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U312 (
    .O(n656),
    .I0(in[149]),
    .I1(n654)
  );
  //AND U312bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U312bar (
    .O(n656bar),
    .I0(inbar[149]),
    .I1(n654bar)
  );
  //OR U313
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U313 (
    .O(n654),
    .I0(in[195]),
    .I1(in[190])
  );
  //AND U313bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U313bar (
    .O(n654bar),
    .I0(inbar[195]),
    .I1(inbar[190])
  );
  //OR U314
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U314 (
    .O(n704),
    .I0(n653),
    .I1(n652)
  );
  //AND U314bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U314bar (
    .O(n704bar),
    .I0(n653bar),
    .I1(n652bar)
  );
  //OR U315
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U315 (
    .O(n652),
    .I0(n651),
    .I1(n650)
  );
  //AND U315bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U315bar (
    .O(n652bar),
    .I0(n651bar),
    .I1(n650bar)
  );
  //OR U316
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U316 (
    .O(n650),
    .I0(in[98]),
    .I1(in[197])
  );
  //AND U316bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U316bar (
    .O(n650bar),
    .I0(inbar[98]),
    .I1(inbar[197])
  );
  //OR U317
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U317 (
    .O(n651),
    .I0(in_11),
    .I1(n649)
  );
  //AND U317bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U317bar (
    .O(n651bar),
    .I0(in_11bar),
    .I1(n649bar)
  );
  //OR U318
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U318 (
    .O(n649),
    .I0(in_26),
    .I1(in_14)
  );
  //AND U318bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U318bar (
    .O(n649bar),
    .I0(in_26bar),
    .I1(in_14bar)
  );
  //OR U319
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U319 (
    .O(n653),
    .I0(n648),
    .I1(n647)
  );
  //AND U319bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U319bar (
    .O(n653bar),
    .I0(n648bar),
    .I1(n647bar)
  );
  //OR U320
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U320 (
    .O(n647),
    .I0(in_35),
    .I1(in_27)
  );
  //AND U320bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U320bar (
    .O(n647bar),
    .I0(in_35bar),
    .I1(in_27bar)
  );
  //OR U321
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U321 (
    .O(n648),
    .I0(in_50),
    .I1(n646)
  );
  //AND U321bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U321bar (
    .O(n648bar),
    .I0(in_50bar),
    .I1(n646bar)
  );
  //OR U322
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U322 (
    .O(n646),
    .I0(in_78),
    .I1(in_61)
  );
  //AND U322bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U322bar (
    .O(n646bar),
    .I0(in_78bar),
    .I1(in_61bar)
  );
  //OR U323
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U323 (
    .O(n720),
    .I0(n942),
    .I1(n645)
  );
  //AND U323bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U323bar (
    .O(n720bar),
    .I0(n942bar),
    .I1(n645bar)
  );
  //OR U324
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U324 (
    .O(n645),
    .I0(in[106]),
    .I1(n863)
  );
  //AND U324bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U324bar (
    .O(n645bar),
    .I0(inbar[106]),
    .I1(n863bar)
  );
  //OR U325
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U325 (
    .O(n863),
    .I0(n644),
    .I1(n643)
  );
  //AND U325bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U325bar (
    .O(n863bar),
    .I0(n644bar),
    .I1(n643bar)
  );
  //OR U326
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U326 (
    .O(n643),
    .I0(n642),
    .I1(n641)
  );
  //AND U326bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U326bar (
    .O(n643bar),
    .I0(n642bar),
    .I1(n641bar)
  );
  //OR U327
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U327 (
    .O(n641),
    .I0(n640),
    .I1(n639)
  );
  //AND U327bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U327bar (
    .O(n641bar),
    .I0(n640bar),
    .I1(n639bar)
  );
  //OR U328
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U328 (
    .O(n639),
    .I0(in[127]),
    .I1(in[122])
  );
  //AND U328bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U328bar (
    .O(n639bar),
    .I0(inbar[127]),
    .I1(inbar[122])
  );
  //OR U329
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U329 (
    .O(n640),
    .I0(in[156]),
    .I1(in[132])
  );
  //AND U329bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U329bar (
    .O(n640bar),
    .I0(inbar[156]),
    .I1(inbar[132])
  );
  //OR U330
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U330 (
    .O(n642),
    .I0(n638),
    .I1(n637)
  );
  //AND U330bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U330bar (
    .O(n642bar),
    .I0(n638bar),
    .I1(n637bar)
  );
  //OR U331
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U331 (
    .O(n637),
    .I0(in[159]),
    .I1(in[157])
  );
  //AND U331bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U331bar (
    .O(n637bar),
    .I0(inbar[159]),
    .I1(inbar[157])
  );
  //OR U332
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U332 (
    .O(n638),
    .I0(in[185]),
    .I1(in[169])
  );
  //AND U332bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U332bar (
    .O(n638bar),
    .I0(inbar[185]),
    .I1(inbar[169])
  );
  //OR U333
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U333 (
    .O(n644),
    .I0(n636),
    .I1(n635)
  );
  //AND U333bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U333bar (
    .O(n644bar),
    .I0(n636bar),
    .I1(n635bar)
  );
  //OR U334
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U334 (
    .O(n635),
    .I0(n634),
    .I1(n633)
  );
  //AND U334bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U334bar (
    .O(n635bar),
    .I0(n634bar),
    .I1(n633bar)
  );
  //OR U335
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U335 (
    .O(n633),
    .I0(in[239]),
    .I1(in[218])
  );
  //AND U335bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U335bar (
    .O(n633bar),
    .I0(inbar[239]),
    .I1(inbar[218])
  );
  //OR U336
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U336 (
    .O(n634),
    .I0(in_13),
    .I1(in[87])
  );
  //AND U336bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U336bar (
    .O(n634bar),
    .I0(in_13bar),
    .I1(inbar[87])
  );
  //OR U337
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U337 (
    .O(n636),
    .I0(n632),
    .I1(n631)
  );
  //AND U337bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U337bar (
    .O(n636bar),
    .I0(n632bar),
    .I1(n631bar)
  );
  //OR U338
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U338 (
    .O(n631),
    .I0(in_72),
    .I1(in_70)
  );
  //AND U338bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U338bar (
    .O(n631bar),
    .I0(in_72bar),
    .I1(in_70bar)
  );
  //OR U339
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U339 (
    .O(n632),
    .I0(in_80),
    .I1(in_74)
  );
  //AND U339bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U339bar (
    .O(n632bar),
    .I0(in_80bar),
    .I1(in_74bar)
  );
  //OR U340
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U340 (
    .O(n942),
    .I0(n630),
    .I1(n629)
  );
  //AND U340bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U340bar (
    .O(n942bar),
    .I0(n630bar),
    .I1(n629bar)
  );
  //OR U341
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U341 (
    .O(n629),
    .I0(n628),
    .I1(n627)
  );
  //AND U341bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U341bar (
    .O(n629bar),
    .I0(n628bar),
    .I1(n627bar)
  );
  //OR U342
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U342 (
    .O(n627),
    .I0(n626),
    .I1(n625)
  );
  //AND U342bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U342bar (
    .O(n627bar),
    .I0(n626bar),
    .I1(n625bar)
  );
  //OR U343
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U343 (
    .O(n625),
    .I0(in[146]),
    .I1(in[100])
  );
  //AND U343bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U343bar (
    .O(n625bar),
    .I0(inbar[146]),
    .I1(inbar[100])
  );
  //OR U344
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U344 (
    .O(n626),
    .I0(in[168]),
    .I1(in[152])
  );
  //AND U344bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U344bar (
    .O(n626bar),
    .I0(inbar[168]),
    .I1(inbar[152])
  );
  //OR U345
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U345 (
    .O(n628),
    .I0(n624),
    .I1(n623)
  );
  //AND U345bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U345bar (
    .O(n628bar),
    .I0(n624bar),
    .I1(n623bar)
  );
  //OR U346
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U346 (
    .O(n623),
    .I0(in[199]),
    .I1(in[182])
  );
  //AND U346bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U346bar (
    .O(n623bar),
    .I0(inbar[199]),
    .I1(inbar[182])
  );
  //OR U347
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U347 (
    .O(n624),
    .I0(in[236]),
    .I1(in[204])
  );
  //AND U347bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U347bar (
    .O(n624bar),
    .I0(inbar[236]),
    .I1(inbar[204])
  );
  //OR U348
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U348 (
    .O(n630),
    .I0(n622),
    .I1(n621)
  );
  //AND U348bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U348bar (
    .O(n630bar),
    .I0(n622bar),
    .I1(n621bar)
  );
  //OR U349
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U349 (
    .O(n621),
    .I0(n620),
    .I1(n619)
  );
  //AND U349bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U349bar (
    .O(n621bar),
    .I0(n620bar),
    .I1(n619bar)
  );
  //OR U350
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U350 (
    .O(n619),
    .I0(in[89]),
    .I1(in[246])
  );
  //AND U350bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U350bar (
    .O(n619bar),
    .I0(inbar[89]),
    .I1(inbar[246])
  );
  //OR U351
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U351 (
    .O(n620),
    .I0(in[95]),
    .I1(in[92])
  );
  //AND U351bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U351bar (
    .O(n620bar),
    .I0(inbar[95]),
    .I1(inbar[92])
  );
  //OR U352
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U352 (
    .O(n622),
    .I0(n618),
    .I1(n617)
  );
  //AND U352bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U352bar (
    .O(n622bar),
    .I0(n618bar),
    .I1(n617bar)
  );
  //OR U353
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U353 (
    .O(n617),
    .I0(in_22),
    .I1(in_16)
  );
  //AND U353bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U353bar (
    .O(n617bar),
    .I0(in_22bar),
    .I1(in_16bar)
  );
  //OR U354
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U354 (
    .O(n618),
    .I0(in_51),
    .I1(in_49)
  );
  //AND U354bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U354bar (
    .O(n618bar),
    .I0(in_51bar),
    .I1(in_49bar)
  );
  //OR U355
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U355 (
    .O(n722),
    .I0(n616),
    .I1(n615)
  );
  //AND U355bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U355bar (
    .O(n722bar),
    .I0(n616bar),
    .I1(n615bar)
  );
  //OR U356
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U356 (
    .O(n615),
    .I0(in[158]),
    .I1(in[115])
  );
  //AND U356bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U356bar (
    .O(n615bar),
    .I0(inbar[158]),
    .I1(inbar[115])
  );
  //OR U357
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U357 (
    .O(n616),
    .I0(in[163]),
    .I1(n614)
  );
  //AND U357bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U357bar (
    .O(n616bar),
    .I0(inbar[163]),
    .I1(n614bar)
  );
  //OR U358
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U358 (
    .O(n614),
    .I0(in[206]),
    .I1(in[165])
  );
  //AND U358bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U358bar (
    .O(n614bar),
    .I0(inbar[206]),
    .I1(inbar[165])
  );
  //OR U359
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U359 (
    .O(n724),
    .I0(n613),
    .I1(n612)
  );
  //AND U359bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U359bar (
    .O(n724bar),
    .I0(n613bar),
    .I1(n612bar)
  );
  //OR U360
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U360 (
    .O(n612),
    .I0(n611),
    .I1(n610)
  );
  //AND U360bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U360bar (
    .O(n612bar),
    .I0(n611bar),
    .I1(n610bar)
  );
  //OR U361
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U361 (
    .O(n610),
    .I0(in[213]),
    .I1(in[207])
  );
  //AND U361bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U361bar (
    .O(n610bar),
    .I0(inbar[213]),
    .I1(inbar[207])
  );
  //OR U362
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U362 (
    .O(n611),
    .I0(in[215]),
    .I1(n609)
  );
  //AND U362bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U362bar (
    .O(n611bar),
    .I0(inbar[215]),
    .I1(n609bar)
  );
  //OR U363
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U363 (
    .O(n609),
    .I0(in[230]),
    .I1(in[220])
  );
  //AND U363bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U363bar (
    .O(n609bar),
    .I0(inbar[230]),
    .I1(inbar[220])
  );
  //OR U364
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U364 (
    .O(n613),
    .I0(n608),
    .I1(n607)
  );
  //AND U364bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U364bar (
    .O(n613bar),
    .I0(n608bar),
    .I1(n607bar)
  );
  //OR U365
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U365 (
    .O(n607),
    .I0(in[251]),
    .I1(in[234])
  );
  //AND U365bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U365bar (
    .O(n607bar),
    .I0(inbar[251]),
    .I1(inbar[234])
  );
  //OR U366
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U366 (
    .O(n608),
    .I0(in_17),
    .I1(n606)
  );
  //AND U366bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U366bar (
    .O(n608bar),
    .I0(in_17bar),
    .I1(n606bar)
  );
  //OR U367
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U367 (
    .O(n606),
    .I0(in_65),
    .I1(in_56)
  );
  //AND U367bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U367bar (
    .O(n606bar),
    .I0(in_65bar),
    .I1(in_56bar)
  );
  //OR U368
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U368 (
    .O(out[0]),
    .I0(n605),
    .I1(n604)
  );
  //AND U368bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U368bar (
    .O(outbar[0]),
    .I0(n605bar),
    .I1(n604bar)
  );
  //OR U369
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U369 (
    .O(n604),
    .I0(n603),
    .I1(n602)
  );
  //AND U369bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U369bar (
    .O(n604bar),
    .I0(n603bar),
    .I1(n602bar)
  );
  //OR U370
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U370 (
    .O(n602),
    .I0(n601),
    .I1(n600)
  );
  //AND U370bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U370bar (
    .O(n602bar),
    .I0(n601bar),
    .I1(n600bar)
  );
  //OR U371
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U371 (
    .O(n600),
    .I0(n820),
    .I1(n785)
  );
  //AND U371bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U371bar (
    .O(n600bar),
    .I0(n820bar),
    .I1(n785bar)
  );
  //OR U372
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U372 (
    .O(n785),
    .I0(n599),
    .I1(n598)
  );
  //AND U372bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U372bar (
    .O(n785bar),
    .I0(n599bar),
    .I1(n598bar)
  );
  //OR U373
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U373 (
    .O(n598),
    .I0(n597),
    .I1(n596)
  );
  //AND U373bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U373bar (
    .O(n598bar),
    .I0(n597bar),
    .I1(n596bar)
  );
  //OR U374
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U374 (
    .O(n596),
    .I0(n595),
    .I1(n594)
  );
  //AND U374bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U374bar (
    .O(n596bar),
    .I0(n595bar),
    .I1(n594bar)
  );
  //OR U375
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U375 (
    .O(n594),
    .I0(in[135]),
    .I1(in[104])
  );
  //AND U375bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U375bar (
    .O(n594bar),
    .I0(inbar[135]),
    .I1(inbar[104])
  );
  //OR U376
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U376 (
    .O(n595),
    .I0(in[188]),
    .I1(in[178])
  );
  //AND U376bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U376bar (
    .O(n595bar),
    .I0(inbar[188]),
    .I1(inbar[178])
  );
  //OR U377
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U377 (
    .O(n597),
    .I0(n593),
    .I1(n592)
  );
  //AND U377bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U377bar (
    .O(n597bar),
    .I0(n593bar),
    .I1(n592bar)
  );
  //OR U378
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U378 (
    .O(n592),
    .I0(in[217]),
    .I1(in[194])
  );
  //AND U378bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U378bar (
    .O(n592bar),
    .I0(inbar[217]),
    .I1(inbar[194])
  );
  //OR U379
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U379 (
    .O(n593),
    .I0(in[237]),
    .I1(in[218])
  );
  //AND U379bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U379bar (
    .O(n593bar),
    .I0(inbar[237]),
    .I1(inbar[218])
  );
  //OR U380
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U380 (
    .O(n599),
    .I0(n591),
    .I1(n590)
  );
  //AND U380bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U380bar (
    .O(n599bar),
    .I0(n591bar),
    .I1(n590bar)
  );
  //OR U381
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U381 (
    .O(n590),
    .I0(n589),
    .I1(n588)
  );
  //AND U381bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U381bar (
    .O(n590bar),
    .I0(n589bar),
    .I1(n588bar)
  );
  //OR U382
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U382 (
    .O(n588),
    .I0(in_2),
    .I1(in_10)
  );
  //AND U382bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U382bar (
    .O(n588bar),
    .I0(in_2bar),
    .I1(in_10bar)
  );
  //OR U383
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U383 (
    .O(n589),
    .I0(in_47),
    .I1(in_22)
  );
  //AND U383bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U383bar (
    .O(n589bar),
    .I0(in_47bar),
    .I1(in_22bar)
  );
  //OR U384
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U384 (
    .O(n591),
    .I0(n587),
    .I1(n586)
  );
  //AND U384bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U384bar (
    .O(n591bar),
    .I0(n587bar),
    .I1(n586bar)
  );
  //OR U385
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U385 (
    .O(n586),
    .I0(in_56),
    .I1(in_54)
  );
  //AND U385bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U385bar (
    .O(n586bar),
    .I0(in_56bar),
    .I1(in_54bar)
  );
  //OR U386
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U386 (
    .O(n587),
    .I0(in_63),
    .I1(in_61)
  );
  //AND U386bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U386bar (
    .O(n587bar),
    .I0(in_63bar),
    .I1(in_61bar)
  );
  //OR U387
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U387 (
    .O(n820),
    .I0(n585),
    .I1(n584)
  );
  //AND U387bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U387bar (
    .O(n820bar),
    .I0(n585bar),
    .I1(n584bar)
  );
  //OR U388
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U388 (
    .O(n584),
    .I0(n583),
    .I1(n582)
  );
  //AND U388bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U388bar (
    .O(n584bar),
    .I0(n583bar),
    .I1(n582bar)
  );
  //OR U389
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U389 (
    .O(n582),
    .I0(n581),
    .I1(n580)
  );
  //AND U389bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U389bar (
    .O(n582bar),
    .I0(n581bar),
    .I1(n580bar)
  );
  //OR U390
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U390 (
    .O(n580),
    .I0(in[158]),
    .I1(in[142])
  );
  //AND U390bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U390bar (
    .O(n580bar),
    .I0(inbar[158]),
    .I1(inbar[142])
  );
  //OR U391
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U391 (
    .O(n581),
    .I0(in[175]),
    .I1(in[164])
  );
  //AND U391bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U391bar (
    .O(n581bar),
    .I0(inbar[175]),
    .I1(inbar[164])
  );
  //OR U392
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U392 (
    .O(n583),
    .I0(n579),
    .I1(n578)
  );
  //AND U392bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U392bar (
    .O(n583bar),
    .I0(n579bar),
    .I1(n578bar)
  );
  //OR U393
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U393 (
    .O(n578),
    .I0(in[228]),
    .I1(in[204])
  );
  //AND U393bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U393bar (
    .O(n578bar),
    .I0(inbar[228]),
    .I1(inbar[204])
  );
  //OR U394
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U394 (
    .O(n579),
    .I0(in[91]),
    .I1(in[87])
  );
  //AND U394bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U394bar (
    .O(n579bar),
    .I0(inbar[91]),
    .I1(inbar[87])
  );
  //OR U395
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U395 (
    .O(n585),
    .I0(n577),
    .I1(n576)
  );
  //AND U395bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U395bar (
    .O(n585bar),
    .I0(n577bar),
    .I1(n576bar)
  );
  //OR U396
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U396 (
    .O(n576),
    .I0(n575),
    .I1(n574)
  );
  //AND U396bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U396bar (
    .O(n576bar),
    .I0(n575bar),
    .I1(n574bar)
  );
  //OR U397
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U397 (
    .O(n574),
    .I0(in_21),
    .I1(in_11)
  );
  //AND U397bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U397bar (
    .O(n574bar),
    .I0(in_21bar),
    .I1(in_11bar)
  );
  //OR U398
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U398 (
    .O(n575),
    .I0(in_5),
    .I1(in_3)
  );
  //AND U398bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U398bar (
    .O(n575bar),
    .I0(in_5bar),
    .I1(in_3bar)
  );
  //OR U399
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U399 (
    .O(n577),
    .I0(n573),
    .I1(n572)
  );
  //AND U399bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U399bar (
    .O(n577bar),
    .I0(n573bar),
    .I1(n572bar)
  );
  //OR U400
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U400 (
    .O(n572),
    .I0(in_68),
    .I1(in_64)
  );
  //AND U400bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U400bar (
    .O(n572bar),
    .I0(in_68bar),
    .I1(in_64bar)
  );
  //OR U401
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U401 (
    .O(n573),
    .I0(in_76),
    .I1(in_73)
  );
  //AND U401bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U401bar (
    .O(n573bar),
    .I0(in_76bar),
    .I1(in_73bar)
  );
  //OR U402
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U402 (
    .O(n601),
    .I0(n778),
    .I1(n571)
  );
  //AND U402bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U402bar (
    .O(n601bar),
    .I0(n778bar),
    .I1(n571bar)
  );
  //OR U403
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U403 (
    .O(n571),
    .I0(in[100]),
    .I1(n965)
  );
  //AND U403bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U403bar (
    .O(n571bar),
    .I0(inbar[100]),
    .I1(n965bar)
  );
  //OR U404
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U404 (
    .O(n965),
    .I0(n570),
    .I1(n569)
  );
  //AND U404bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U404bar (
    .O(n965bar),
    .I0(n570bar),
    .I1(n569bar)
  );
  //OR U405
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U405 (
    .O(n569),
    .I0(n568),
    .I1(n567)
  );
  //AND U405bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U405bar (
    .O(n569bar),
    .I0(n568bar),
    .I1(n567bar)
  );
  //OR U406
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U406 (
    .O(n567),
    .I0(n566),
    .I1(n565)
  );
  //AND U406bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U406bar (
    .O(n567bar),
    .I0(n566bar),
    .I1(n565bar)
  );
  //OR U407
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U407 (
    .O(n565),
    .I0(n817),
    .I1(n750)
  );
  //AND U407bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U407bar (
    .O(n565bar),
    .I0(n817bar),
    .I1(n750bar)
  );
  //OR U408
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U408 (
    .O(n750),
    .I0(n564),
    .I1(n563)
  );
  //AND U408bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U408bar (
    .O(n750bar),
    .I0(n564bar),
    .I1(n563bar)
  );
  //OR U409
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U409 (
    .O(n563),
    .I0(n562),
    .I1(n561)
  );
  //AND U409bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U409bar (
    .O(n563bar),
    .I0(n562bar),
    .I1(n561bar)
  );
  //OR U410
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U410 (
    .O(n561),
    .I0(n560),
    .I1(n559)
  );
  //AND U410bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U410bar (
    .O(n561bar),
    .I0(n560bar),
    .I1(n559bar)
  );
  //OR U411
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U411 (
    .O(n559),
    .I0(in[119]),
    .I1(in[103])
  );
  //AND U411bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U411bar (
    .O(n559bar),
    .I0(inbar[119]),
    .I1(inbar[103])
  );
  //OR U412
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U412 (
    .O(n560),
    .I0(in[137]),
    .I1(in[133])
  );
  //AND U412bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U412bar (
    .O(n560bar),
    .I0(inbar[137]),
    .I1(inbar[133])
  );
  //OR U413
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U413 (
    .O(n562),
    .I0(n558),
    .I1(n557)
  );
  //AND U413bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U413bar (
    .O(n562bar),
    .I0(n558bar),
    .I1(n557bar)
  );
  //OR U414
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U414 (
    .O(n557),
    .I0(in[176]),
    .I1(in[173])
  );
  //AND U414bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U414bar (
    .O(n557bar),
    .I0(inbar[176]),
    .I1(inbar[173])
  );
  //OR U415
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U415 (
    .O(n558),
    .I0(in[210]),
    .I1(in[181])
  );
  //AND U415bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U415bar (
    .O(n558bar),
    .I0(inbar[210]),
    .I1(inbar[181])
  );
  //OR U416
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U416 (
    .O(n564),
    .I0(n556),
    .I1(n555)
  );
  //AND U416bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U416bar (
    .O(n564bar),
    .I0(n556bar),
    .I1(n555bar)
  );
  //OR U417
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U417 (
    .O(n555),
    .I0(n554),
    .I1(n553)
  );
  //AND U417bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U417bar (
    .O(n555bar),
    .I0(n554bar),
    .I1(n553bar)
  );
  //OR U418
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U418 (
    .O(n553),
    .I0(in_13),
    .I1(in[234])
  );
  //AND U418bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U418bar (
    .O(n553bar),
    .I0(in_13bar),
    .I1(inbar[234])
  );
  //OR U419
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U419 (
    .O(n554),
    .I0(in_38),
    .I1(in_32)
  );
  //AND U419bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U419bar (
    .O(n554bar),
    .I0(in_38bar),
    .I1(in_32bar)
  );
  //OR U420
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U420 (
    .O(n556),
    .I0(n552),
    .I1(n551)
  );
  //AND U420bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U420bar (
    .O(n556bar),
    .I0(n552bar),
    .I1(n551bar)
  );
  //OR U421
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U421 (
    .O(n551),
    .I0(in_42),
    .I1(in_41)
  );
  //AND U421bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U421bar (
    .O(n551bar),
    .I0(in_42bar),
    .I1(in_41bar)
  );
  //OR U422
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U422 (
    .O(n552),
    .I0(in_7),
    .I1(in_49)
  );
  //AND U422bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U422bar (
    .O(n552bar),
    .I0(in_7bar),
    .I1(in_49bar)
  );
  //OR U423
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U423 (
    .O(n817),
    .I0(n550),
    .I1(n549)
  );
  //AND U423bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U423bar (
    .O(n817bar),
    .I0(n550bar),
    .I1(n549bar)
  );
  //OR U424
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U424 (
    .O(n549),
    .I0(n548),
    .I1(n547)
  );
  //AND U424bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U424bar (
    .O(n549bar),
    .I0(n548bar),
    .I1(n547bar)
  );
  //OR U425
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U425 (
    .O(n547),
    .I0(n546),
    .I1(n545)
  );
  //AND U425bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U425bar (
    .O(n547bar),
    .I0(n546bar),
    .I1(n545bar)
  );
  //OR U426
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U426 (
    .O(n545),
    .I0(in[159]),
    .I1(in[105])
  );
  //AND U426bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U426bar (
    .O(n545bar),
    .I0(inbar[159]),
    .I1(inbar[105])
  );
  //OR U427
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U427 (
    .O(n546),
    .I0(in[206]),
    .I1(in[183])
  );
  //AND U427bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U427bar (
    .O(n546bar),
    .I0(inbar[206]),
    .I1(inbar[183])
  );
  //OR U428
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U428 (
    .O(n548),
    .I0(n544),
    .I1(n543)
  );
  //AND U428bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U428bar (
    .O(n548bar),
    .I0(n544bar),
    .I1(n543bar)
  );
  //OR U429
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U429 (
    .O(n543),
    .I0(in[229]),
    .I1(in[219])
  );
  //AND U429bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U429bar (
    .O(n543bar),
    .I0(inbar[229]),
    .I1(inbar[219])
  );
  //OR U430
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U430 (
    .O(n544),
    .I0(in[235]),
    .I1(in[232])
  );
  //AND U430bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U430bar (
    .O(n544bar),
    .I0(inbar[235]),
    .I1(inbar[232])
  );
  //OR U431
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U431 (
    .O(n550),
    .I0(n542),
    .I1(n541)
  );
  //AND U431bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U431bar (
    .O(n550bar),
    .I0(n542bar),
    .I1(n541bar)
  );
  //OR U432
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U432 (
    .O(n541),
    .I0(n540),
    .I1(n539)
  );
  //AND U432bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U432bar (
    .O(n541bar),
    .I0(n540bar),
    .I1(n539bar)
  );
  //OR U433
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U433 (
    .O(n539),
    .I0(in[249]),
    .I1(in[242])
  );
  //AND U433bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U433bar (
    .O(n539bar),
    .I0(inbar[249]),
    .I1(inbar[242])
  );
  //OR U434
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U434 (
    .O(n540),
    .I0(in[89]),
    .I1(in[254])
  );
  //AND U434bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U434bar (
    .O(n540bar),
    .I0(inbar[89]),
    .I1(inbar[254])
  );
  //OR U435
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U435 (
    .O(n542),
    .I0(n538),
    .I1(n537)
  );
  //AND U435bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U435bar (
    .O(n542bar),
    .I0(n538bar),
    .I1(n537bar)
  );
  //OR U436
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U436 (
    .O(n537),
    .I0(in_14),
    .I1(in[99])
  );
  //AND U436bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U436bar (
    .O(n537bar),
    .I0(in_14bar),
    .I1(inbar[99])
  );
  //OR U437
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U437 (
    .O(n538),
    .I0(in_60),
    .I1(in_18)
  );
  //AND U437bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U437bar (
    .O(n538bar),
    .I0(in_60bar),
    .I1(in_18bar)
  );
  //OR U438
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U438 (
    .O(n566),
    .I0(in[113]),
    .I1(n763)
  );
  //AND U438bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U438bar (
    .O(n566bar),
    .I0(inbar[113]),
    .I1(n763bar)
  );
  //OR U439
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U439 (
    .O(n763),
    .I0(n536),
    .I1(n535)
  );
  //AND U439bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U439bar (
    .O(n763bar),
    .I0(n536bar),
    .I1(n535bar)
  );
  //OR U440
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U440 (
    .O(n535),
    .I0(n534),
    .I1(n533)
  );
  //AND U440bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U440bar (
    .O(n535bar),
    .I0(n534bar),
    .I1(n533bar)
  );
  //OR U441
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U441 (
    .O(n533),
    .I0(n532),
    .I1(n531)
  );
  //AND U441bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U441bar (
    .O(n533bar),
    .I0(n532bar),
    .I1(n531bar)
  );
  //OR U442
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U442 (
    .O(n531),
    .I0(in[115]),
    .I1(in[110])
  );
  //AND U442bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U442bar (
    .O(n531bar),
    .I0(inbar[115]),
    .I1(inbar[110])
  );
  //OR U443
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U443 (
    .O(n532),
    .I0(in[125]),
    .I1(in[117])
  );
  //AND U443bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U443bar (
    .O(n532bar),
    .I0(inbar[125]),
    .I1(inbar[117])
  );
  //OR U444
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U444 (
    .O(n534),
    .I0(n530),
    .I1(n529)
  );
  //AND U444bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U444bar (
    .O(n534bar),
    .I0(n530bar),
    .I1(n529bar)
  );
  //OR U445
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U445 (
    .O(n529),
    .I0(in[180]),
    .I1(in[128])
  );
  //AND U445bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U445bar (
    .O(n529bar),
    .I0(inbar[180]),
    .I1(inbar[128])
  );
  //OR U446
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U446 (
    .O(n530),
    .I0(in[205]),
    .I1(in[201])
  );
  //AND U446bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U446bar (
    .O(n530bar),
    .I0(inbar[205]),
    .I1(inbar[201])
  );
  //OR U447
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U447 (
    .O(n536),
    .I0(n528),
    .I1(n527)
  );
  //AND U447bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U447bar (
    .O(n536bar),
    .I0(n528bar),
    .I1(n527bar)
  );
  //OR U448
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U448 (
    .O(n527),
    .I0(n526),
    .I1(n525)
  );
  //AND U448bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U448bar (
    .O(n527bar),
    .I0(n526bar),
    .I1(n525bar)
  );
  //OR U449
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U449 (
    .O(n525),
    .I0(in[244]),
    .I1(in[239])
  );
  //AND U449bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U449bar (
    .O(n525bar),
    .I0(inbar[244]),
    .I1(inbar[239])
  );
  //OR U450
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U450 (
    .O(n526),
    .I0(in[95]),
    .I1(in[83])
  );
  //AND U450bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U450bar (
    .O(n526bar),
    .I0(inbar[95]),
    .I1(inbar[83])
  );
  //OR U451
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U451 (
    .O(n528),
    .I0(n524),
    .I1(n523)
  );
  //AND U451bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U451bar (
    .O(n528bar),
    .I0(n524bar),
    .I1(n523bar)
  );
  //OR U452
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U452 (
    .O(n523),
    .I0(in_24),
    .I1(in[97])
  );
  //AND U452bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U452bar (
    .O(n523bar),
    .I0(in_24bar),
    .I1(inbar[97])
  );
  //OR U453
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U453 (
    .O(n524),
    .I0(in_33),
    .I1(in_27)
  );
  //AND U453bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U453bar (
    .O(n524bar),
    .I0(in_33bar),
    .I1(in_27bar)
  );
  //OR U454
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U454 (
    .O(n568),
    .I0(n522),
    .I1(n521)
  );
  //AND U454bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U454bar (
    .O(n568bar),
    .I0(n522bar),
    .I1(n521bar)
  );
  //OR U455
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U455 (
    .O(n521),
    .I0(in[145]),
    .I1(in[126])
  );
  //AND U455bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U455bar (
    .O(n521bar),
    .I0(inbar[145]),
    .I1(inbar[126])
  );
  //OR U456
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U456 (
    .O(n522),
    .I0(in[169]),
    .I1(n520)
  );
  //AND U456bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U456bar (
    .O(n522bar),
    .I0(inbar[169]),
    .I1(n520bar)
  );
  //OR U457
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U457 (
    .O(n520),
    .I0(in[221]),
    .I1(in[172])
  );
  //AND U457bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U457bar (
    .O(n520bar),
    .I0(inbar[221]),
    .I1(inbar[172])
  );
  //OR U458
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U458 (
    .O(n570),
    .I0(n519),
    .I1(n518)
  );
  //AND U458bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U458bar (
    .O(n570bar),
    .I0(n519bar),
    .I1(n518bar)
  );
  //OR U459
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U459 (
    .O(n518),
    .I0(n517),
    .I1(n516)
  );
  //AND U459bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U459bar (
    .O(n518bar),
    .I0(n517bar),
    .I1(n516bar)
  );
  //OR U460
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U460 (
    .O(n516),
    .I0(in[241]),
    .I1(in[224])
  );
  //AND U460bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U460bar (
    .O(n516bar),
    .I0(inbar[241]),
    .I1(inbar[224])
  );
  //OR U461
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U461 (
    .O(n517),
    .I0(in[86]),
    .I1(n515)
  );
  //AND U461bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U461bar (
    .O(n517bar),
    .I0(inbar[86]),
    .I1(n515bar)
  );
  //OR U462
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U462 (
    .O(n515),
    .I0(in_43),
    .I1(in_34)
  );
  //AND U462bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U462bar (
    .O(n515bar),
    .I0(in_43bar),
    .I1(in_34bar)
  );
  //OR U463
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U463 (
    .O(n519),
    .I0(n514),
    .I1(n513)
  );
  //AND U463bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U463bar (
    .O(n519bar),
    .I0(n514bar),
    .I1(n513bar)
  );
  //OR U464
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U464 (
    .O(n513),
    .I0(in_65),
    .I1(in_51)
  );
  //AND U464bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U464bar (
    .O(n513bar),
    .I0(in_65bar),
    .I1(in_51bar)
  );
  //OR U465
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U465 (
    .O(n514),
    .I0(in_75),
    .I1(n512)
  );
  //AND U465bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U465bar (
    .O(n514bar),
    .I0(in_75bar),
    .I1(n512bar)
  );
  //OR U466
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U466 (
    .O(n512),
    .I0(in_81),
    .I1(in_77)
  );
  //AND U466bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U466bar (
    .O(n512bar),
    .I0(in_81bar),
    .I1(in_77bar)
  );
  //OR U467
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U467 (
    .O(n778),
    .I0(n511),
    .I1(n510)
  );
  //AND U467bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U467bar (
    .O(n778bar),
    .I0(n511bar),
    .I1(n510bar)
  );
  //OR U468
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U468 (
    .O(n510),
    .I0(n509),
    .I1(n508)
  );
  //AND U468bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U468bar (
    .O(n510bar),
    .I0(n509bar),
    .I1(n508bar)
  );
  //OR U469
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U469 (
    .O(n508),
    .I0(n507),
    .I1(n506)
  );
  //AND U469bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U469bar (
    .O(n508bar),
    .I0(n507bar),
    .I1(n506bar)
  );
  //OR U470
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U470 (
    .O(n506),
    .I0(in[107]),
    .I1(in[101])
  );
  //AND U470bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U470bar (
    .O(n506bar),
    .I0(inbar[107]),
    .I1(inbar[101])
  );
  //OR U471
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U471 (
    .O(n507),
    .I0(in[139]),
    .I1(in[132])
  );
  //AND U471bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U471bar (
    .O(n507bar),
    .I0(inbar[139]),
    .I1(inbar[132])
  );
  //OR U472
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U472 (
    .O(n509),
    .I0(n505),
    .I1(n504)
  );
  //AND U472bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U472bar (
    .O(n509bar),
    .I0(n505bar),
    .I1(n504bar)
  );
  //OR U473
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U473 (
    .O(n504),
    .I0(in[146]),
    .I1(in[141])
  );
  //AND U473bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U473bar (
    .O(n504bar),
    .I0(inbar[146]),
    .I1(inbar[141])
  );
  //OR U474
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U474 (
    .O(n505),
    .I0(in[203]),
    .I1(in[179])
  );
  //AND U474bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U474bar (
    .O(n505bar),
    .I0(inbar[203]),
    .I1(inbar[179])
  );
  //OR U475
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U475 (
    .O(n511),
    .I0(n503),
    .I1(n502)
  );
  //AND U475bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U475bar (
    .O(n511bar),
    .I0(n503bar),
    .I1(n502bar)
  );
  //OR U476
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U476 (
    .O(n502),
    .I0(n501),
    .I1(n500)
  );
  //AND U476bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U476bar (
    .O(n502bar),
    .I0(n501bar),
    .I1(n500bar)
  );
  //OR U477
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U477 (
    .O(n500),
    .I0(in[243]),
    .I1(in[222])
  );
  //AND U477bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U477bar (
    .O(n500bar),
    .I0(inbar[243]),
    .I1(inbar[222])
  );
  //OR U478
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U478 (
    .O(n501),
    .I0(in[251]),
    .I1(in[250])
  );
  //AND U478bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U478bar (
    .O(n501bar),
    .I0(inbar[251]),
    .I1(inbar[250])
  );
  //OR U479
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U479 (
    .O(n503),
    .I0(n499),
    .I1(n498)
  );
  //AND U479bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U479bar (
    .O(n503bar),
    .I0(n499bar),
    .I1(n498bar)
  );
  //OR U480
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U480 (
    .O(n498),
    .I0(in_37),
    .I1(in_19)
  );
  //AND U480bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U480bar (
    .O(n498bar),
    .I0(in_37bar),
    .I1(in_19bar)
  );
  //OR U481
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U481 (
    .O(n499),
    .I0(in_78),
    .I1(in_6)
  );
  //AND U481bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U481bar (
    .O(n499bar),
    .I0(in_78bar),
    .I1(in_6bar)
  );
  //OR U482
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U482 (
    .O(n603),
    .I0(n497),
    .I1(n496)
  );
  //AND U482bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U482bar (
    .O(n603bar),
    .I0(n497bar),
    .I1(n496bar)
  );
  //OR U483
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U483 (
    .O(n496),
    .I0(in[112]),
    .I1(in[102])
  );
  //AND U483bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U483bar (
    .O(n496bar),
    .I0(inbar[112]),
    .I1(inbar[102])
  );
  //OR U484
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U484 (
    .O(n497),
    .I0(in[123]),
    .I1(n495)
  );
  //AND U484bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U484bar (
    .O(n497bar),
    .I0(inbar[123]),
    .I1(n495bar)
  );
  //OR U485
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U485 (
    .O(n495),
    .I0(in[143]),
    .I1(in[130])
  );
  //AND U485bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U485bar (
    .O(n495bar),
    .I0(inbar[143]),
    .I1(inbar[130])
  );
  //OR U486
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U486 (
    .O(n605),
    .I0(n494),
    .I1(n493)
  );
  //AND U486bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U486bar (
    .O(n605bar),
    .I0(n494bar),
    .I1(n493bar)
  );
  //OR U487
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U487 (
    .O(n493),
    .I0(n492),
    .I1(n491)
  );
  //AND U487bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U487bar (
    .O(n493bar),
    .I0(n492bar),
    .I1(n491bar)
  );
  //OR U488
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U488 (
    .O(n491),
    .I0(in[216]),
    .I1(in[213])
  );
  //AND U488bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U488bar (
    .O(n491bar),
    .I0(inbar[216]),
    .I1(inbar[213])
  );
  //OR U489
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U489 (
    .O(n492),
    .I0(in[227]),
    .I1(n490)
  );
  //AND U489bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U489bar (
    .O(n492bar),
    .I0(inbar[227]),
    .I1(n490bar)
  );
  //OR U490
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U490 (
    .O(n490),
    .I0(in_0),
    .I1(in[248])
  );
  //AND U490bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U490bar (
    .O(n490bar),
    .I0(in_0bar),
    .I1(inbar[248])
  );
  //OR U491
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U491 (
    .O(n494),
    .I0(n489),
    .I1(n488)
  );
  //AND U491bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U491bar (
    .O(n494bar),
    .I0(n489bar),
    .I1(n488bar)
  );
  //OR U492
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U492 (
    .O(n488),
    .I0(in_46),
    .I1(in_44)
  );
  //AND U492bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U492bar (
    .O(n488bar),
    .I0(in_46bar),
    .I1(in_44bar)
  );
  //OR U493
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U493 (
    .O(n489),
    .I0(in_50),
    .I1(n487)
  );
  //AND U493bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U493bar (
    .O(n489bar),
    .I0(in_50bar),
    .I1(n487bar)
  );
  //OR U494
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U494 (
    .O(n487),
    .I0(in_9),
    .I1(in_80)
  );
  //AND U494bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U494bar (
    .O(n487bar),
    .I0(in_9bar),
    .I1(in_80bar)
  );
endmodule

module sBox_12 ( in, out );

  input wire [7:0] in;
//input_done

  output wire [7:0] out;
//output_done

  wire [255:0] decodeOut;
//wire_done

  decode_12 dec ( .in(in), .out(decodeOut) );
  encode_12 enc ( .in(decodeOut), .out(out) );
endmodule

module CD2_49 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD2_50 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD2_51 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD2_52 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD4_25 ( a, b, y );

  input wire [3:0] a;
  input wire [3:0] b;
  wire [3:0] abar;
  wire [3:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
//input_done

  output wire [15:0] y;
  wire [15:0] ybar;
//output_done

//wire_done

  //AND U1
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1 (
    .O(y[9]),
    .I0(b[1]),
    .I1(a[2])
  );
  //OR U1bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1bar (
    .O(ybar[9]),
    .I0(bbar[1]),
    .I1(abar[2])
  );
  //AND U2
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2 (
    .O(y[8]),
    .I0(b[0]),
    .I1(a[2])
  );
  //OR U2bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2bar (
    .O(ybar[8]),
    .I0(bbar[0]),
    .I1(abar[2])
  );
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[7]),
    .I0(b[3]),
    .I1(a[1])
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[7]),
    .I0(bbar[3]),
    .I1(abar[1])
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[6]),
    .I0(b[2]),
    .I1(a[1])
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[6]),
    .I0(bbar[2]),
    .I1(abar[1])
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[5]),
    .I0(a[1]),
    .I1(b[1])
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[5]),
    .I0(abar[1]),
    .I1(bbar[1])
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[4]),
    .I0(a[1]),
    .I1(b[0])
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[4]),
    .I0(abar[1]),
    .I1(bbar[0])
  );
  //AND U7
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7 (
    .O(y[3]),
    .I0(a[0]),
    .I1(b[3])
  );
  //OR U7bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7bar (
    .O(ybar[3]),
    .I0(abar[0]),
    .I1(bbar[3])
  );
  //AND U8
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8 (
    .O(y[2]),
    .I0(a[0]),
    .I1(b[2])
  );
  //OR U8bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8bar (
    .O(ybar[2]),
    .I0(abar[0]),
    .I1(bbar[2])
  );
  //AND U9
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9 (
    .O(y[1]),
    .I0(a[0]),
    .I1(b[1])
  );
  //OR U9bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9bar (
    .O(ybar[1]),
    .I0(abar[0]),
    .I1(bbar[1])
  );
  //AND U10
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10 (
    .O(y[15]),
    .I0(a[3]),
    .I1(b[3])
  );
  //OR U10bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10bar (
    .O(ybar[15]),
    .I0(abar[3]),
    .I1(bbar[3])
  );
  //AND U11
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11 (
    .O(y[14]),
    .I0(a[3]),
    .I1(b[2])
  );
  //OR U11bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11bar (
    .O(ybar[14]),
    .I0(abar[3]),
    .I1(bbar[2])
  );
  //AND U12
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12 (
    .O(y[13]),
    .I0(a[3]),
    .I1(b[1])
  );
  //OR U12bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12bar (
    .O(ybar[13]),
    .I0(abar[3]),
    .I1(bbar[1])
  );
  //AND U13
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13 (
    .O(y[12]),
    .I0(a[3]),
    .I1(b[0])
  );
  //OR U13bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13bar (
    .O(ybar[12]),
    .I0(abar[3]),
    .I1(bbar[0])
  );
  //AND U14
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14 (
    .O(y[11]),
    .I0(b[3]),
    .I1(a[2])
  );
  //OR U14bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14bar (
    .O(ybar[11]),
    .I0(bbar[3]),
    .I1(abar[2])
  );
  //AND U15
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15 (
    .O(y[10]),
    .I0(b[2]),
    .I1(a[2])
  );
  //OR U15bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15bar (
    .O(ybar[10]),
    .I0(bbar[2]),
    .I1(abar[2])
  );
  //AND U16
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16 (
    .O(y[0]),
    .I0(a[0]),
    .I1(b[0])
  );
  //OR U16bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16bar (
    .O(ybar[0]),
    .I0(abar[0]),
    .I1(bbar[0])
  );
endmodule

module CD4_26 ( a, b, y );

  input wire [3:0] a;
  input wire [3:0] b;
  wire [3:0] abar;
  wire [3:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
//input_done

  output wire [15:0] y;
  wire [15:0] ybar;
//output_done

//wire_done

  //AND U1
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1 (
    .O(y[9]),
    .I0(b[1]),
    .I1(a[2])
  );
  //OR U1bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1bar (
    .O(ybar[9]),
    .I0(bbar[1]),
    .I1(abar[2])
  );
  //AND U2
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2 (
    .O(y[8]),
    .I0(b[0]),
    .I1(a[2])
  );
  //OR U2bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2bar (
    .O(ybar[8]),
    .I0(bbar[0]),
    .I1(abar[2])
  );
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[7]),
    .I0(b[3]),
    .I1(a[1])
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[7]),
    .I0(bbar[3]),
    .I1(abar[1])
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[6]),
    .I0(b[2]),
    .I1(a[1])
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[6]),
    .I0(bbar[2]),
    .I1(abar[1])
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[5]),
    .I0(a[1]),
    .I1(b[1])
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[5]),
    .I0(abar[1]),
    .I1(bbar[1])
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[4]),
    .I0(a[1]),
    .I1(b[0])
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[4]),
    .I0(abar[1]),
    .I1(bbar[0])
  );
  //AND U7
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7 (
    .O(y[3]),
    .I0(a[0]),
    .I1(b[3])
  );
  //OR U7bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7bar (
    .O(ybar[3]),
    .I0(abar[0]),
    .I1(bbar[3])
  );
  //AND U8
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8 (
    .O(y[2]),
    .I0(a[0]),
    .I1(b[2])
  );
  //OR U8bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8bar (
    .O(ybar[2]),
    .I0(abar[0]),
    .I1(bbar[2])
  );
  //AND U9
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9 (
    .O(y[1]),
    .I0(a[0]),
    .I1(b[1])
  );
  //OR U9bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9bar (
    .O(ybar[1]),
    .I0(abar[0]),
    .I1(bbar[1])
  );
  //AND U10
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10 (
    .O(y[15]),
    .I0(a[3]),
    .I1(b[3])
  );
  //OR U10bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10bar (
    .O(ybar[15]),
    .I0(abar[3]),
    .I1(bbar[3])
  );
  //AND U11
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11 (
    .O(y[14]),
    .I0(a[3]),
    .I1(b[2])
  );
  //OR U11bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11bar (
    .O(ybar[14]),
    .I0(abar[3]),
    .I1(bbar[2])
  );
  //AND U12
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12 (
    .O(y[13]),
    .I0(a[3]),
    .I1(b[1])
  );
  //OR U12bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12bar (
    .O(ybar[13]),
    .I0(abar[3]),
    .I1(bbar[1])
  );
  //AND U13
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13 (
    .O(y[12]),
    .I0(a[3]),
    .I1(b[0])
  );
  //OR U13bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13bar (
    .O(ybar[12]),
    .I0(abar[3]),
    .I1(bbar[0])
  );
  //AND U14
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14 (
    .O(y[11]),
    .I0(b[3]),
    .I1(a[2])
  );
  //OR U14bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14bar (
    .O(ybar[11]),
    .I0(bbar[3]),
    .I1(abar[2])
  );
  //AND U15
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15 (
    .O(y[10]),
    .I0(b[2]),
    .I1(a[2])
  );
  //OR U15bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15bar (
    .O(ybar[10]),
    .I0(bbar[2]),
    .I1(abar[2])
  );
  //AND U16
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16 (
    .O(y[0]),
    .I0(a[0]),
    .I1(b[0])
  );
  //OR U16bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16bar (
    .O(ybar[0]),
    .I0(abar[0]),
    .I1(bbar[0])
  );
endmodule

module CD16_13 ( a, b, y );

  input wire [15:0] a;
  input wire [15:0] b;
  wire [15:0] abar;
  wire [15:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign abar[8] = ~a[8];
  assign abar[9] = ~a[9];
  assign abar[10] = ~a[10];
  assign abar[11] = ~a[11];
  assign abar[12] = ~a[12];
  assign abar[13] = ~a[13];
  assign abar[14] = ~a[14];
  assign abar[15] = ~a[15];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign bbar[8] = ~b[8];
  assign bbar[9] = ~b[9];
  assign bbar[10] = ~b[10];
  assign bbar[11] = ~b[11];
  assign bbar[12] = ~b[12];
  assign bbar[13] = ~b[13];
  assign bbar[14] = ~b[14];
  assign bbar[15] = ~b[15];
//input_done

  output wire [255:0] y;
  wire [255:0] ybar;
//output_done

//wire_done

  //AND U1
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1 (
    .O(y[9]),
    .I0(b[9]),
    .I1(a[0])
  );
  //OR U1bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1bar (
    .O(ybar[9]),
    .I0(bbar[9]),
    .I1(abar[0])
  );
  //AND U2
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2 (
    .O(y[99]),
    .I0(b[3]),
    .I1(a[6])
  );
  //OR U2bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2bar (
    .O(ybar[99]),
    .I0(bbar[3]),
    .I1(abar[6])
  );
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[98]),
    .I0(b[2]),
    .I1(a[6])
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[98]),
    .I0(bbar[2]),
    .I1(abar[6])
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[97]),
    .I0(b[1]),
    .I1(a[6])
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[97]),
    .I0(bbar[1]),
    .I1(abar[6])
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[96]),
    .I0(b[0]),
    .I1(a[6])
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[96]),
    .I0(bbar[0]),
    .I1(abar[6])
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[95]),
    .I0(b[15]),
    .I1(a[5])
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[95]),
    .I0(bbar[15]),
    .I1(abar[5])
  );
  //AND U7
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7 (
    .O(y[94]),
    .I0(b[14]),
    .I1(a[5])
  );
  //OR U7bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7bar (
    .O(ybar[94]),
    .I0(bbar[14]),
    .I1(abar[5])
  );
  //AND U8
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8 (
    .O(y[93]),
    .I0(b[13]),
    .I1(a[5])
  );
  //OR U8bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8bar (
    .O(ybar[93]),
    .I0(bbar[13]),
    .I1(abar[5])
  );
  //AND U9
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9 (
    .O(y[92]),
    .I0(b[12]),
    .I1(a[5])
  );
  //OR U9bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9bar (
    .O(ybar[92]),
    .I0(bbar[12]),
    .I1(abar[5])
  );
  //AND U10
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10 (
    .O(y[91]),
    .I0(b[11]),
    .I1(a[5])
  );
  //OR U10bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10bar (
    .O(ybar[91]),
    .I0(bbar[11]),
    .I1(abar[5])
  );
  //AND U11
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11 (
    .O(y[90]),
    .I0(b[10]),
    .I1(a[5])
  );
  //OR U11bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11bar (
    .O(ybar[90]),
    .I0(bbar[10]),
    .I1(abar[5])
  );
  //AND U12
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12 (
    .O(y[8]),
    .I0(b[8]),
    .I1(a[0])
  );
  //OR U12bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12bar (
    .O(ybar[8]),
    .I0(bbar[8]),
    .I1(abar[0])
  );
  //AND U13
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13 (
    .O(y[89]),
    .I0(a[5]),
    .I1(b[9])
  );
  //OR U13bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13bar (
    .O(ybar[89]),
    .I0(abar[5]),
    .I1(bbar[9])
  );
  //AND U14
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14 (
    .O(y[88]),
    .I0(b[8]),
    .I1(a[5])
  );
  //OR U14bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14bar (
    .O(ybar[88]),
    .I0(bbar[8]),
    .I1(abar[5])
  );
  //AND U15
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15 (
    .O(y[87]),
    .I0(b[7]),
    .I1(a[5])
  );
  //OR U15bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15bar (
    .O(ybar[87]),
    .I0(bbar[7]),
    .I1(abar[5])
  );
  //AND U16
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16 (
    .O(y[86]),
    .I0(b[6]),
    .I1(a[5])
  );
  //OR U16bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16bar (
    .O(ybar[86]),
    .I0(bbar[6]),
    .I1(abar[5])
  );
  //AND U17
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U17 (
    .O(y[85]),
    .I0(b[5]),
    .I1(a[5])
  );
  //OR U17bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U17bar (
    .O(ybar[85]),
    .I0(bbar[5]),
    .I1(abar[5])
  );
  //AND U18
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U18 (
    .O(y[84]),
    .I0(b[4]),
    .I1(a[5])
  );
  //OR U18bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U18bar (
    .O(ybar[84]),
    .I0(bbar[4]),
    .I1(abar[5])
  );
  //AND U19
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U19 (
    .O(y[83]),
    .I0(a[5]),
    .I1(b[3])
  );
  //OR U19bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U19bar (
    .O(ybar[83]),
    .I0(abar[5]),
    .I1(bbar[3])
  );
  //AND U20
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U20 (
    .O(y[82]),
    .I0(a[5]),
    .I1(b[2])
  );
  //OR U20bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U20bar (
    .O(ybar[82]),
    .I0(abar[5]),
    .I1(bbar[2])
  );
  //AND U21
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U21 (
    .O(y[81]),
    .I0(a[5]),
    .I1(b[1])
  );
  //OR U21bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U21bar (
    .O(ybar[81]),
    .I0(abar[5]),
    .I1(bbar[1])
  );
  //AND U22
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U22 (
    .O(y[80]),
    .I0(a[5]),
    .I1(b[0])
  );
  //OR U22bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U22bar (
    .O(ybar[80]),
    .I0(abar[5]),
    .I1(bbar[0])
  );
  //AND U23
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U23 (
    .O(y[7]),
    .I0(b[7]),
    .I1(a[0])
  );
  //OR U23bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U23bar (
    .O(ybar[7]),
    .I0(bbar[7]),
    .I1(abar[0])
  );
  //AND U24
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U24 (
    .O(y[79]),
    .I0(a[4]),
    .I1(b[15])
  );
  //OR U24bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U24bar (
    .O(ybar[79]),
    .I0(abar[4]),
    .I1(bbar[15])
  );
  //AND U25
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U25 (
    .O(y[78]),
    .I0(a[4]),
    .I1(b[14])
  );
  //OR U25bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U25bar (
    .O(ybar[78]),
    .I0(abar[4]),
    .I1(bbar[14])
  );
  //AND U26
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U26 (
    .O(y[77]),
    .I0(a[4]),
    .I1(b[13])
  );
  //OR U26bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U26bar (
    .O(ybar[77]),
    .I0(abar[4]),
    .I1(bbar[13])
  );
  //AND U27
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U27 (
    .O(y[76]),
    .I0(a[4]),
    .I1(b[12])
  );
  //OR U27bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U27bar (
    .O(ybar[76]),
    .I0(abar[4]),
    .I1(bbar[12])
  );
  //AND U28
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U28 (
    .O(y[75]),
    .I0(a[4]),
    .I1(b[11])
  );
  //OR U28bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U28bar (
    .O(ybar[75]),
    .I0(abar[4]),
    .I1(bbar[11])
  );
  //AND U29
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U29 (
    .O(y[74]),
    .I0(a[4]),
    .I1(b[10])
  );
  //OR U29bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U29bar (
    .O(ybar[74]),
    .I0(abar[4]),
    .I1(bbar[10])
  );
  //AND U30
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U30 (
    .O(y[73]),
    .I0(a[4]),
    .I1(b[9])
  );
  //OR U30bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U30bar (
    .O(ybar[73]),
    .I0(abar[4]),
    .I1(bbar[9])
  );
  //AND U31
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U31 (
    .O(y[72]),
    .I0(a[4]),
    .I1(b[8])
  );
  //OR U31bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U31bar (
    .O(ybar[72]),
    .I0(abar[4]),
    .I1(bbar[8])
  );
  //AND U32
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U32 (
    .O(y[71]),
    .I0(a[4]),
    .I1(b[7])
  );
  //OR U32bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U32bar (
    .O(ybar[71]),
    .I0(abar[4]),
    .I1(bbar[7])
  );
  //AND U33
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U33 (
    .O(y[70]),
    .I0(a[4]),
    .I1(b[6])
  );
  //OR U33bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U33bar (
    .O(ybar[70]),
    .I0(abar[4]),
    .I1(bbar[6])
  );
  //AND U34
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U34 (
    .O(y[6]),
    .I0(b[6]),
    .I1(a[0])
  );
  //OR U34bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U34bar (
    .O(ybar[6]),
    .I0(bbar[6]),
    .I1(abar[0])
  );
  //AND U35
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U35 (
    .O(y[69]),
    .I0(a[4]),
    .I1(b[5])
  );
  //OR U35bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U35bar (
    .O(ybar[69]),
    .I0(abar[4]),
    .I1(bbar[5])
  );
  //AND U36
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U36 (
    .O(y[68]),
    .I0(a[4]),
    .I1(b[4])
  );
  //OR U36bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U36bar (
    .O(ybar[68]),
    .I0(abar[4]),
    .I1(bbar[4])
  );
  //AND U37
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U37 (
    .O(y[67]),
    .I0(a[4]),
    .I1(b[3])
  );
  //OR U37bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U37bar (
    .O(ybar[67]),
    .I0(abar[4]),
    .I1(bbar[3])
  );
  //AND U38
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U38 (
    .O(y[66]),
    .I0(a[4]),
    .I1(b[2])
  );
  //OR U38bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U38bar (
    .O(ybar[66]),
    .I0(abar[4]),
    .I1(bbar[2])
  );
  //AND U39
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U39 (
    .O(y[65]),
    .I0(a[4]),
    .I1(b[1])
  );
  //OR U39bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U39bar (
    .O(ybar[65]),
    .I0(abar[4]),
    .I1(bbar[1])
  );
  //AND U40
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U40 (
    .O(y[64]),
    .I0(a[4]),
    .I1(b[0])
  );
  //OR U40bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U40bar (
    .O(ybar[64]),
    .I0(abar[4]),
    .I1(bbar[0])
  );
  //AND U41
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U41 (
    .O(y[63]),
    .I0(a[3]),
    .I1(b[15])
  );
  //OR U41bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U41bar (
    .O(ybar[63]),
    .I0(abar[3]),
    .I1(bbar[15])
  );
  //AND U42
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U42 (
    .O(y[62]),
    .I0(a[3]),
    .I1(b[14])
  );
  //OR U42bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U42bar (
    .O(ybar[62]),
    .I0(abar[3]),
    .I1(bbar[14])
  );
  //AND U43
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U43 (
    .O(y[61]),
    .I0(a[3]),
    .I1(b[13])
  );
  //OR U43bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U43bar (
    .O(ybar[61]),
    .I0(abar[3]),
    .I1(bbar[13])
  );
  //AND U44
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U44 (
    .O(y[60]),
    .I0(a[3]),
    .I1(b[12])
  );
  //OR U44bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U44bar (
    .O(ybar[60]),
    .I0(abar[3]),
    .I1(bbar[12])
  );
  //AND U45
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U45 (
    .O(y[5]),
    .I0(b[5]),
    .I1(a[0])
  );
  //OR U45bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U45bar (
    .O(ybar[5]),
    .I0(bbar[5]),
    .I1(abar[0])
  );
  //AND U46
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U46 (
    .O(y[59]),
    .I0(a[3]),
    .I1(b[11])
  );
  //OR U46bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U46bar (
    .O(ybar[59]),
    .I0(abar[3]),
    .I1(bbar[11])
  );
  //AND U47
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U47 (
    .O(y[58]),
    .I0(a[3]),
    .I1(b[10])
  );
  //OR U47bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U47bar (
    .O(ybar[58]),
    .I0(abar[3]),
    .I1(bbar[10])
  );
  //AND U48
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U48 (
    .O(y[57]),
    .I0(a[3]),
    .I1(b[9])
  );
  //OR U48bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U48bar (
    .O(ybar[57]),
    .I0(abar[3]),
    .I1(bbar[9])
  );
  //AND U49
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U49 (
    .O(y[56]),
    .I0(a[3]),
    .I1(b[8])
  );
  //OR U49bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U49bar (
    .O(ybar[56]),
    .I0(abar[3]),
    .I1(bbar[8])
  );
  //AND U50
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U50 (
    .O(y[55]),
    .I0(a[3]),
    .I1(b[7])
  );
  //OR U50bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U50bar (
    .O(ybar[55]),
    .I0(abar[3]),
    .I1(bbar[7])
  );
  //AND U51
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U51 (
    .O(y[54]),
    .I0(a[3]),
    .I1(b[6])
  );
  //OR U51bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U51bar (
    .O(ybar[54]),
    .I0(abar[3]),
    .I1(bbar[6])
  );
  //AND U52
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U52 (
    .O(y[53]),
    .I0(a[3]),
    .I1(b[5])
  );
  //OR U52bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U52bar (
    .O(ybar[53]),
    .I0(abar[3]),
    .I1(bbar[5])
  );
  //AND U53
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U53 (
    .O(y[52]),
    .I0(a[3]),
    .I1(b[4])
  );
  //OR U53bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U53bar (
    .O(ybar[52]),
    .I0(abar[3]),
    .I1(bbar[4])
  );
  //AND U54
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U54 (
    .O(y[51]),
    .I0(a[3]),
    .I1(b[3])
  );
  //OR U54bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U54bar (
    .O(ybar[51]),
    .I0(abar[3]),
    .I1(bbar[3])
  );
  //AND U55
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U55 (
    .O(y[50]),
    .I0(a[3]),
    .I1(b[2])
  );
  //OR U55bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U55bar (
    .O(ybar[50]),
    .I0(abar[3]),
    .I1(bbar[2])
  );
  //AND U56
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U56 (
    .O(y[4]),
    .I0(b[4]),
    .I1(a[0])
  );
  //OR U56bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U56bar (
    .O(ybar[4]),
    .I0(bbar[4]),
    .I1(abar[0])
  );
  //AND U57
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U57 (
    .O(y[49]),
    .I0(a[3]),
    .I1(b[1])
  );
  //OR U57bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U57bar (
    .O(ybar[49]),
    .I0(abar[3]),
    .I1(bbar[1])
  );
  //AND U58
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U58 (
    .O(y[48]),
    .I0(a[3]),
    .I1(b[0])
  );
  //OR U58bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U58bar (
    .O(ybar[48]),
    .I0(abar[3]),
    .I1(bbar[0])
  );
  //AND U59
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U59 (
    .O(y[47]),
    .I0(a[2]),
    .I1(b[15])
  );
  //OR U59bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U59bar (
    .O(ybar[47]),
    .I0(abar[2]),
    .I1(bbar[15])
  );
  //AND U60
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U60 (
    .O(y[46]),
    .I0(a[2]),
    .I1(b[14])
  );
  //OR U60bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U60bar (
    .O(ybar[46]),
    .I0(abar[2]),
    .I1(bbar[14])
  );
  //AND U61
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U61 (
    .O(y[45]),
    .I0(a[2]),
    .I1(b[13])
  );
  //OR U61bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U61bar (
    .O(ybar[45]),
    .I0(abar[2]),
    .I1(bbar[13])
  );
  //AND U62
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U62 (
    .O(y[44]),
    .I0(a[2]),
    .I1(b[12])
  );
  //OR U62bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U62bar (
    .O(ybar[44]),
    .I0(abar[2]),
    .I1(bbar[12])
  );
  //AND U63
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U63 (
    .O(y[43]),
    .I0(a[2]),
    .I1(b[11])
  );
  //OR U63bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U63bar (
    .O(ybar[43]),
    .I0(abar[2]),
    .I1(bbar[11])
  );
  //AND U64
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U64 (
    .O(y[42]),
    .I0(a[2]),
    .I1(b[10])
  );
  //OR U64bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U64bar (
    .O(ybar[42]),
    .I0(abar[2]),
    .I1(bbar[10])
  );
  //AND U65
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U65 (
    .O(y[41]),
    .I0(a[2]),
    .I1(b[9])
  );
  //OR U65bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U65bar (
    .O(ybar[41]),
    .I0(abar[2]),
    .I1(bbar[9])
  );
  //AND U66
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U66 (
    .O(y[40]),
    .I0(a[2]),
    .I1(b[8])
  );
  //OR U66bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U66bar (
    .O(ybar[40]),
    .I0(abar[2]),
    .I1(bbar[8])
  );
  //AND U67
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U67 (
    .O(y[3]),
    .I0(b[3]),
    .I1(a[0])
  );
  //OR U67bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U67bar (
    .O(ybar[3]),
    .I0(bbar[3]),
    .I1(abar[0])
  );
  //AND U68
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U68 (
    .O(y[39]),
    .I0(a[2]),
    .I1(b[7])
  );
  //OR U68bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U68bar (
    .O(ybar[39]),
    .I0(abar[2]),
    .I1(bbar[7])
  );
  //AND U69
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U69 (
    .O(y[38]),
    .I0(a[2]),
    .I1(b[6])
  );
  //OR U69bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U69bar (
    .O(ybar[38]),
    .I0(abar[2]),
    .I1(bbar[6])
  );
  //AND U70
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U70 (
    .O(y[37]),
    .I0(a[2]),
    .I1(b[5])
  );
  //OR U70bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U70bar (
    .O(ybar[37]),
    .I0(abar[2]),
    .I1(bbar[5])
  );
  //AND U71
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U71 (
    .O(y[36]),
    .I0(a[2]),
    .I1(b[4])
  );
  //OR U71bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U71bar (
    .O(ybar[36]),
    .I0(abar[2]),
    .I1(bbar[4])
  );
  //AND U72
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U72 (
    .O(y[35]),
    .I0(a[2]),
    .I1(b[3])
  );
  //OR U72bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U72bar (
    .O(ybar[35]),
    .I0(abar[2]),
    .I1(bbar[3])
  );
  //AND U73
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U73 (
    .O(y[34]),
    .I0(a[2]),
    .I1(b[2])
  );
  //OR U73bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U73bar (
    .O(ybar[34]),
    .I0(abar[2]),
    .I1(bbar[2])
  );
  //AND U74
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U74 (
    .O(y[33]),
    .I0(a[2]),
    .I1(b[1])
  );
  //OR U74bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U74bar (
    .O(ybar[33]),
    .I0(abar[2]),
    .I1(bbar[1])
  );
  //AND U75
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U75 (
    .O(y[32]),
    .I0(a[2]),
    .I1(b[0])
  );
  //OR U75bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U75bar (
    .O(ybar[32]),
    .I0(abar[2]),
    .I1(bbar[0])
  );
  //AND U76
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U76 (
    .O(y[31]),
    .I0(a[1]),
    .I1(b[15])
  );
  //OR U76bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U76bar (
    .O(ybar[31]),
    .I0(abar[1]),
    .I1(bbar[15])
  );
  //AND U77
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U77 (
    .O(y[30]),
    .I0(a[1]),
    .I1(b[14])
  );
  //OR U77bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U77bar (
    .O(ybar[30]),
    .I0(abar[1]),
    .I1(bbar[14])
  );
  //AND U78
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U78 (
    .O(y[2]),
    .I0(b[2]),
    .I1(a[0])
  );
  //OR U78bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U78bar (
    .O(ybar[2]),
    .I0(bbar[2]),
    .I1(abar[0])
  );
  //AND U79
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U79 (
    .O(y[29]),
    .I0(a[1]),
    .I1(b[13])
  );
  //OR U79bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U79bar (
    .O(ybar[29]),
    .I0(abar[1]),
    .I1(bbar[13])
  );
  //AND U80
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U80 (
    .O(y[28]),
    .I0(a[1]),
    .I1(b[12])
  );
  //OR U80bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U80bar (
    .O(ybar[28]),
    .I0(abar[1]),
    .I1(bbar[12])
  );
  //AND U81
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U81 (
    .O(y[27]),
    .I0(a[1]),
    .I1(b[11])
  );
  //OR U81bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U81bar (
    .O(ybar[27]),
    .I0(abar[1]),
    .I1(bbar[11])
  );
  //AND U82
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U82 (
    .O(y[26]),
    .I0(a[1]),
    .I1(b[10])
  );
  //OR U82bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U82bar (
    .O(ybar[26]),
    .I0(abar[1]),
    .I1(bbar[10])
  );
  //AND U83
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U83 (
    .O(y[25]),
    .I0(a[1]),
    .I1(b[9])
  );
  //OR U83bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U83bar (
    .O(ybar[25]),
    .I0(abar[1]),
    .I1(bbar[9])
  );
  //AND U84
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U84 (
    .O(y[255]),
    .I0(a[15]),
    .I1(b[15])
  );
  //OR U84bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U84bar (
    .O(ybar[255]),
    .I0(abar[15]),
    .I1(bbar[15])
  );
  //AND U85
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U85 (
    .O(y[254]),
    .I0(a[15]),
    .I1(b[14])
  );
  //OR U85bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U85bar (
    .O(ybar[254]),
    .I0(abar[15]),
    .I1(bbar[14])
  );
  //AND U86
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U86 (
    .O(y[253]),
    .I0(a[15]),
    .I1(b[13])
  );
  //OR U86bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U86bar (
    .O(ybar[253]),
    .I0(abar[15]),
    .I1(bbar[13])
  );
  //AND U87
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U87 (
    .O(y[252]),
    .I0(a[15]),
    .I1(b[12])
  );
  //OR U87bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U87bar (
    .O(ybar[252]),
    .I0(abar[15]),
    .I1(bbar[12])
  );
  //AND U88
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U88 (
    .O(y[251]),
    .I0(a[15]),
    .I1(b[11])
  );
  //OR U88bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U88bar (
    .O(ybar[251]),
    .I0(abar[15]),
    .I1(bbar[11])
  );
  //AND U89
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U89 (
    .O(y[250]),
    .I0(a[15]),
    .I1(b[10])
  );
  //OR U89bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U89bar (
    .O(ybar[250]),
    .I0(abar[15]),
    .I1(bbar[10])
  );
  //AND U90
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U90 (
    .O(y[24]),
    .I0(a[1]),
    .I1(b[8])
  );
  //OR U90bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U90bar (
    .O(ybar[24]),
    .I0(abar[1]),
    .I1(bbar[8])
  );
  //AND U91
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U91 (
    .O(y[249]),
    .I0(a[15]),
    .I1(b[9])
  );
  //OR U91bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U91bar (
    .O(ybar[249]),
    .I0(abar[15]),
    .I1(bbar[9])
  );
  //AND U92
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U92 (
    .O(y[248]),
    .I0(a[15]),
    .I1(b[8])
  );
  //OR U92bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U92bar (
    .O(ybar[248]),
    .I0(abar[15]),
    .I1(bbar[8])
  );
  //AND U93
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U93 (
    .O(y[247]),
    .I0(a[15]),
    .I1(b[7])
  );
  //OR U93bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U93bar (
    .O(ybar[247]),
    .I0(abar[15]),
    .I1(bbar[7])
  );
  //AND U94
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U94 (
    .O(y[246]),
    .I0(a[15]),
    .I1(b[6])
  );
  //OR U94bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U94bar (
    .O(ybar[246]),
    .I0(abar[15]),
    .I1(bbar[6])
  );
  //AND U95
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U95 (
    .O(y[245]),
    .I0(a[15]),
    .I1(b[5])
  );
  //OR U95bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U95bar (
    .O(ybar[245]),
    .I0(abar[15]),
    .I1(bbar[5])
  );
  //AND U96
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U96 (
    .O(y[244]),
    .I0(a[15]),
    .I1(b[4])
  );
  //OR U96bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U96bar (
    .O(ybar[244]),
    .I0(abar[15]),
    .I1(bbar[4])
  );
  //AND U97
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U97 (
    .O(y[243]),
    .I0(a[15]),
    .I1(b[3])
  );
  //OR U97bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U97bar (
    .O(ybar[243]),
    .I0(abar[15]),
    .I1(bbar[3])
  );
  //AND U98
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U98 (
    .O(y[242]),
    .I0(a[15]),
    .I1(b[2])
  );
  //OR U98bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U98bar (
    .O(ybar[242]),
    .I0(abar[15]),
    .I1(bbar[2])
  );
  //AND U99
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U99 (
    .O(y[241]),
    .I0(a[15]),
    .I1(b[1])
  );
  //OR U99bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U99bar (
    .O(ybar[241]),
    .I0(abar[15]),
    .I1(bbar[1])
  );
  //AND U100
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U100 (
    .O(y[240]),
    .I0(a[15]),
    .I1(b[0])
  );
  //OR U100bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U100bar (
    .O(ybar[240]),
    .I0(abar[15]),
    .I1(bbar[0])
  );
  //AND U101
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U101 (
    .O(y[23]),
    .I0(a[1]),
    .I1(b[7])
  );
  //OR U101bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U101bar (
    .O(ybar[23]),
    .I0(abar[1]),
    .I1(bbar[7])
  );
  //AND U102
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U102 (
    .O(y[239]),
    .I0(a[14]),
    .I1(b[15])
  );
  //OR U102bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U102bar (
    .O(ybar[239]),
    .I0(abar[14]),
    .I1(bbar[15])
  );
  //AND U103
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U103 (
    .O(y[238]),
    .I0(a[14]),
    .I1(b[14])
  );
  //OR U103bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U103bar (
    .O(ybar[238]),
    .I0(abar[14]),
    .I1(bbar[14])
  );
  //AND U104
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U104 (
    .O(y[237]),
    .I0(a[14]),
    .I1(b[13])
  );
  //OR U104bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U104bar (
    .O(ybar[237]),
    .I0(abar[14]),
    .I1(bbar[13])
  );
  //AND U105
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U105 (
    .O(y[236]),
    .I0(a[14]),
    .I1(b[12])
  );
  //OR U105bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U105bar (
    .O(ybar[236]),
    .I0(abar[14]),
    .I1(bbar[12])
  );
  //AND U106
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U106 (
    .O(y[235]),
    .I0(a[14]),
    .I1(b[11])
  );
  //OR U106bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U106bar (
    .O(ybar[235]),
    .I0(abar[14]),
    .I1(bbar[11])
  );
  //AND U107
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U107 (
    .O(y[234]),
    .I0(a[14]),
    .I1(b[10])
  );
  //OR U107bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U107bar (
    .O(ybar[234]),
    .I0(abar[14]),
    .I1(bbar[10])
  );
  //AND U108
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U108 (
    .O(y[233]),
    .I0(a[14]),
    .I1(b[9])
  );
  //OR U108bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U108bar (
    .O(ybar[233]),
    .I0(abar[14]),
    .I1(bbar[9])
  );
  //AND U109
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U109 (
    .O(y[232]),
    .I0(a[14]),
    .I1(b[8])
  );
  //OR U109bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U109bar (
    .O(ybar[232]),
    .I0(abar[14]),
    .I1(bbar[8])
  );
  //AND U110
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U110 (
    .O(y[231]),
    .I0(a[14]),
    .I1(b[7])
  );
  //OR U110bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U110bar (
    .O(ybar[231]),
    .I0(abar[14]),
    .I1(bbar[7])
  );
  //AND U111
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U111 (
    .O(y[230]),
    .I0(a[14]),
    .I1(b[6])
  );
  //OR U111bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U111bar (
    .O(ybar[230]),
    .I0(abar[14]),
    .I1(bbar[6])
  );
  //AND U112
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U112 (
    .O(y[22]),
    .I0(a[1]),
    .I1(b[6])
  );
  //OR U112bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U112bar (
    .O(ybar[22]),
    .I0(abar[1]),
    .I1(bbar[6])
  );
  //AND U113
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U113 (
    .O(y[229]),
    .I0(a[14]),
    .I1(b[5])
  );
  //OR U113bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U113bar (
    .O(ybar[229]),
    .I0(abar[14]),
    .I1(bbar[5])
  );
  //AND U114
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U114 (
    .O(y[228]),
    .I0(a[14]),
    .I1(b[4])
  );
  //OR U114bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U114bar (
    .O(ybar[228]),
    .I0(abar[14]),
    .I1(bbar[4])
  );
  //AND U115
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U115 (
    .O(y[227]),
    .I0(a[14]),
    .I1(b[3])
  );
  //OR U115bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U115bar (
    .O(ybar[227]),
    .I0(abar[14]),
    .I1(bbar[3])
  );
  //AND U116
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U116 (
    .O(y[226]),
    .I0(a[14]),
    .I1(b[2])
  );
  //OR U116bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U116bar (
    .O(ybar[226]),
    .I0(abar[14]),
    .I1(bbar[2])
  );
  //AND U117
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U117 (
    .O(y[225]),
    .I0(a[14]),
    .I1(b[1])
  );
  //OR U117bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U117bar (
    .O(ybar[225]),
    .I0(abar[14]),
    .I1(bbar[1])
  );
  //AND U118
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U118 (
    .O(y[224]),
    .I0(a[14]),
    .I1(b[0])
  );
  //OR U118bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U118bar (
    .O(ybar[224]),
    .I0(abar[14]),
    .I1(bbar[0])
  );
  //AND U119
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U119 (
    .O(y[223]),
    .I0(a[13]),
    .I1(b[15])
  );
  //OR U119bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U119bar (
    .O(ybar[223]),
    .I0(abar[13]),
    .I1(bbar[15])
  );
  //AND U120
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U120 (
    .O(y[222]),
    .I0(a[13]),
    .I1(b[14])
  );
  //OR U120bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U120bar (
    .O(ybar[222]),
    .I0(abar[13]),
    .I1(bbar[14])
  );
  //AND U121
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U121 (
    .O(y[221]),
    .I0(a[13]),
    .I1(b[13])
  );
  //OR U121bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U121bar (
    .O(ybar[221]),
    .I0(abar[13]),
    .I1(bbar[13])
  );
  //AND U122
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U122 (
    .O(y[220]),
    .I0(a[13]),
    .I1(b[12])
  );
  //OR U122bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U122bar (
    .O(ybar[220]),
    .I0(abar[13]),
    .I1(bbar[12])
  );
  //AND U123
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U123 (
    .O(y[21]),
    .I0(a[1]),
    .I1(b[5])
  );
  //OR U123bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U123bar (
    .O(ybar[21]),
    .I0(abar[1]),
    .I1(bbar[5])
  );
  //AND U124
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U124 (
    .O(y[219]),
    .I0(a[13]),
    .I1(b[11])
  );
  //OR U124bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U124bar (
    .O(ybar[219]),
    .I0(abar[13]),
    .I1(bbar[11])
  );
  //AND U125
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U125 (
    .O(y[218]),
    .I0(a[13]),
    .I1(b[10])
  );
  //OR U125bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U125bar (
    .O(ybar[218]),
    .I0(abar[13]),
    .I1(bbar[10])
  );
  //AND U126
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U126 (
    .O(y[217]),
    .I0(a[13]),
    .I1(b[9])
  );
  //OR U126bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U126bar (
    .O(ybar[217]),
    .I0(abar[13]),
    .I1(bbar[9])
  );
  //AND U127
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U127 (
    .O(y[216]),
    .I0(a[13]),
    .I1(b[8])
  );
  //OR U127bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U127bar (
    .O(ybar[216]),
    .I0(abar[13]),
    .I1(bbar[8])
  );
  //AND U128
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U128 (
    .O(y[215]),
    .I0(a[13]),
    .I1(b[7])
  );
  //OR U128bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U128bar (
    .O(ybar[215]),
    .I0(abar[13]),
    .I1(bbar[7])
  );
  //AND U129
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U129 (
    .O(y[214]),
    .I0(a[13]),
    .I1(b[6])
  );
  //OR U129bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U129bar (
    .O(ybar[214]),
    .I0(abar[13]),
    .I1(bbar[6])
  );
  //AND U130
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U130 (
    .O(y[213]),
    .I0(a[13]),
    .I1(b[5])
  );
  //OR U130bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U130bar (
    .O(ybar[213]),
    .I0(abar[13]),
    .I1(bbar[5])
  );
  //AND U131
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U131 (
    .O(y[212]),
    .I0(a[13]),
    .I1(b[4])
  );
  //OR U131bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U131bar (
    .O(ybar[212]),
    .I0(abar[13]),
    .I1(bbar[4])
  );
  //AND U132
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U132 (
    .O(y[211]),
    .I0(a[13]),
    .I1(b[3])
  );
  //OR U132bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U132bar (
    .O(ybar[211]),
    .I0(abar[13]),
    .I1(bbar[3])
  );
  //AND U133
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U133 (
    .O(y[210]),
    .I0(a[13]),
    .I1(b[2])
  );
  //OR U133bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U133bar (
    .O(ybar[210]),
    .I0(abar[13]),
    .I1(bbar[2])
  );
  //AND U134
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U134 (
    .O(y[20]),
    .I0(a[1]),
    .I1(b[4])
  );
  //OR U134bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U134bar (
    .O(ybar[20]),
    .I0(abar[1]),
    .I1(bbar[4])
  );
  //AND U135
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U135 (
    .O(y[209]),
    .I0(a[13]),
    .I1(b[1])
  );
  //OR U135bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U135bar (
    .O(ybar[209]),
    .I0(abar[13]),
    .I1(bbar[1])
  );
  //AND U136
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U136 (
    .O(y[208]),
    .I0(a[13]),
    .I1(b[0])
  );
  //OR U136bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U136bar (
    .O(ybar[208]),
    .I0(abar[13]),
    .I1(bbar[0])
  );
  //AND U137
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U137 (
    .O(y[207]),
    .I0(a[12]),
    .I1(b[15])
  );
  //OR U137bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U137bar (
    .O(ybar[207]),
    .I0(abar[12]),
    .I1(bbar[15])
  );
  //AND U138
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U138 (
    .O(y[206]),
    .I0(a[12]),
    .I1(b[14])
  );
  //OR U138bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U138bar (
    .O(ybar[206]),
    .I0(abar[12]),
    .I1(bbar[14])
  );
  //AND U139
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U139 (
    .O(y[205]),
    .I0(a[12]),
    .I1(b[13])
  );
  //OR U139bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U139bar (
    .O(ybar[205]),
    .I0(abar[12]),
    .I1(bbar[13])
  );
  //AND U140
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U140 (
    .O(y[204]),
    .I0(a[12]),
    .I1(b[12])
  );
  //OR U140bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U140bar (
    .O(ybar[204]),
    .I0(abar[12]),
    .I1(bbar[12])
  );
  //AND U141
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U141 (
    .O(y[203]),
    .I0(a[12]),
    .I1(b[11])
  );
  //OR U141bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U141bar (
    .O(ybar[203]),
    .I0(abar[12]),
    .I1(bbar[11])
  );
  //AND U142
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U142 (
    .O(y[202]),
    .I0(a[12]),
    .I1(b[10])
  );
  //OR U142bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U142bar (
    .O(ybar[202]),
    .I0(abar[12]),
    .I1(bbar[10])
  );
  //AND U143
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U143 (
    .O(y[201]),
    .I0(a[12]),
    .I1(b[9])
  );
  //OR U143bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U143bar (
    .O(ybar[201]),
    .I0(abar[12]),
    .I1(bbar[9])
  );
  //AND U144
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U144 (
    .O(y[200]),
    .I0(a[12]),
    .I1(b[8])
  );
  //OR U144bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U144bar (
    .O(ybar[200]),
    .I0(abar[12]),
    .I1(bbar[8])
  );
  //AND U145
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U145 (
    .O(y[1]),
    .I0(b[1]),
    .I1(a[0])
  );
  //OR U145bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U145bar (
    .O(ybar[1]),
    .I0(bbar[1]),
    .I1(abar[0])
  );
  //AND U146
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U146 (
    .O(y[19]),
    .I0(a[1]),
    .I1(b[3])
  );
  //OR U146bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U146bar (
    .O(ybar[19]),
    .I0(abar[1]),
    .I1(bbar[3])
  );
  //AND U147
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U147 (
    .O(y[199]),
    .I0(a[12]),
    .I1(b[7])
  );
  //OR U147bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U147bar (
    .O(ybar[199]),
    .I0(abar[12]),
    .I1(bbar[7])
  );
  //AND U148
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U148 (
    .O(y[198]),
    .I0(a[12]),
    .I1(b[6])
  );
  //OR U148bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U148bar (
    .O(ybar[198]),
    .I0(abar[12]),
    .I1(bbar[6])
  );
  //AND U149
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U149 (
    .O(y[197]),
    .I0(a[12]),
    .I1(b[5])
  );
  //OR U149bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U149bar (
    .O(ybar[197]),
    .I0(abar[12]),
    .I1(bbar[5])
  );
  //AND U150
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U150 (
    .O(y[196]),
    .I0(a[12]),
    .I1(b[4])
  );
  //OR U150bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U150bar (
    .O(ybar[196]),
    .I0(abar[12]),
    .I1(bbar[4])
  );
  //AND U151
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U151 (
    .O(y[195]),
    .I0(a[12]),
    .I1(b[3])
  );
  //OR U151bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U151bar (
    .O(ybar[195]),
    .I0(abar[12]),
    .I1(bbar[3])
  );
  //AND U152
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U152 (
    .O(y[194]),
    .I0(a[12]),
    .I1(b[2])
  );
  //OR U152bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U152bar (
    .O(ybar[194]),
    .I0(abar[12]),
    .I1(bbar[2])
  );
  //AND U153
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U153 (
    .O(y[193]),
    .I0(a[12]),
    .I1(b[1])
  );
  //OR U153bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U153bar (
    .O(ybar[193]),
    .I0(abar[12]),
    .I1(bbar[1])
  );
  //AND U154
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U154 (
    .O(y[192]),
    .I0(a[12]),
    .I1(b[0])
  );
  //OR U154bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U154bar (
    .O(ybar[192]),
    .I0(abar[12]),
    .I1(bbar[0])
  );
  //AND U155
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U155 (
    .O(y[191]),
    .I0(a[11]),
    .I1(b[15])
  );
  //OR U155bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U155bar (
    .O(ybar[191]),
    .I0(abar[11]),
    .I1(bbar[15])
  );
  //AND U156
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U156 (
    .O(y[190]),
    .I0(a[11]),
    .I1(b[14])
  );
  //OR U156bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U156bar (
    .O(ybar[190]),
    .I0(abar[11]),
    .I1(bbar[14])
  );
  //AND U157
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U157 (
    .O(y[18]),
    .I0(a[1]),
    .I1(b[2])
  );
  //OR U157bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U157bar (
    .O(ybar[18]),
    .I0(abar[1]),
    .I1(bbar[2])
  );
  //AND U158
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U158 (
    .O(y[189]),
    .I0(a[11]),
    .I1(b[13])
  );
  //OR U158bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U158bar (
    .O(ybar[189]),
    .I0(abar[11]),
    .I1(bbar[13])
  );
  //AND U159
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U159 (
    .O(y[188]),
    .I0(a[11]),
    .I1(b[12])
  );
  //OR U159bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U159bar (
    .O(ybar[188]),
    .I0(abar[11]),
    .I1(bbar[12])
  );
  //AND U160
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U160 (
    .O(y[187]),
    .I0(a[11]),
    .I1(b[11])
  );
  //OR U160bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U160bar (
    .O(ybar[187]),
    .I0(abar[11]),
    .I1(bbar[11])
  );
  //AND U161
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U161 (
    .O(y[186]),
    .I0(a[11]),
    .I1(b[10])
  );
  //OR U161bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U161bar (
    .O(ybar[186]),
    .I0(abar[11]),
    .I1(bbar[10])
  );
  //AND U162
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U162 (
    .O(y[185]),
    .I0(a[11]),
    .I1(b[9])
  );
  //OR U162bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U162bar (
    .O(ybar[185]),
    .I0(abar[11]),
    .I1(bbar[9])
  );
  //AND U163
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U163 (
    .O(y[184]),
    .I0(a[11]),
    .I1(b[8])
  );
  //OR U163bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U163bar (
    .O(ybar[184]),
    .I0(abar[11]),
    .I1(bbar[8])
  );
  //AND U164
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U164 (
    .O(y[183]),
    .I0(a[11]),
    .I1(b[7])
  );
  //OR U164bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U164bar (
    .O(ybar[183]),
    .I0(abar[11]),
    .I1(bbar[7])
  );
  //AND U165
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U165 (
    .O(y[182]),
    .I0(a[11]),
    .I1(b[6])
  );
  //OR U165bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U165bar (
    .O(ybar[182]),
    .I0(abar[11]),
    .I1(bbar[6])
  );
  //AND U166
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U166 (
    .O(y[181]),
    .I0(a[11]),
    .I1(b[5])
  );
  //OR U166bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U166bar (
    .O(ybar[181]),
    .I0(abar[11]),
    .I1(bbar[5])
  );
  //AND U167
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U167 (
    .O(y[180]),
    .I0(a[11]),
    .I1(b[4])
  );
  //OR U167bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U167bar (
    .O(ybar[180]),
    .I0(abar[11]),
    .I1(bbar[4])
  );
  //AND U168
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U168 (
    .O(y[17]),
    .I0(a[1]),
    .I1(b[1])
  );
  //OR U168bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U168bar (
    .O(ybar[17]),
    .I0(abar[1]),
    .I1(bbar[1])
  );
  //AND U169
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U169 (
    .O(y[179]),
    .I0(a[11]),
    .I1(b[3])
  );
  //OR U169bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U169bar (
    .O(ybar[179]),
    .I0(abar[11]),
    .I1(bbar[3])
  );
  //AND U170
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U170 (
    .O(y[178]),
    .I0(a[11]),
    .I1(b[2])
  );
  //OR U170bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U170bar (
    .O(ybar[178]),
    .I0(abar[11]),
    .I1(bbar[2])
  );
  //AND U171
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U171 (
    .O(y[177]),
    .I0(a[11]),
    .I1(b[1])
  );
  //OR U171bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U171bar (
    .O(ybar[177]),
    .I0(abar[11]),
    .I1(bbar[1])
  );
  //AND U172
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U172 (
    .O(y[176]),
    .I0(a[11]),
    .I1(b[0])
  );
  //OR U172bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U172bar (
    .O(ybar[176]),
    .I0(abar[11]),
    .I1(bbar[0])
  );
  //AND U173
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U173 (
    .O(y[175]),
    .I0(a[10]),
    .I1(b[15])
  );
  //OR U173bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U173bar (
    .O(ybar[175]),
    .I0(abar[10]),
    .I1(bbar[15])
  );
  //AND U174
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U174 (
    .O(y[174]),
    .I0(a[10]),
    .I1(b[14])
  );
  //OR U174bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U174bar (
    .O(ybar[174]),
    .I0(abar[10]),
    .I1(bbar[14])
  );
  //AND U175
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U175 (
    .O(y[173]),
    .I0(a[10]),
    .I1(b[13])
  );
  //OR U175bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U175bar (
    .O(ybar[173]),
    .I0(abar[10]),
    .I1(bbar[13])
  );
  //AND U176
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U176 (
    .O(y[172]),
    .I0(a[10]),
    .I1(b[12])
  );
  //OR U176bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U176bar (
    .O(ybar[172]),
    .I0(abar[10]),
    .I1(bbar[12])
  );
  //AND U177
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U177 (
    .O(y[171]),
    .I0(a[10]),
    .I1(b[11])
  );
  //OR U177bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U177bar (
    .O(ybar[171]),
    .I0(abar[10]),
    .I1(bbar[11])
  );
  //AND U178
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U178 (
    .O(y[170]),
    .I0(a[10]),
    .I1(b[10])
  );
  //OR U178bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U178bar (
    .O(ybar[170]),
    .I0(abar[10]),
    .I1(bbar[10])
  );
  //AND U179
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U179 (
    .O(y[16]),
    .I0(a[1]),
    .I1(b[0])
  );
  //OR U179bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U179bar (
    .O(ybar[16]),
    .I0(abar[1]),
    .I1(bbar[0])
  );
  //AND U180
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U180 (
    .O(y[169]),
    .I0(a[10]),
    .I1(b[9])
  );
  //OR U180bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U180bar (
    .O(ybar[169]),
    .I0(abar[10]),
    .I1(bbar[9])
  );
  //AND U181
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U181 (
    .O(y[168]),
    .I0(a[10]),
    .I1(b[8])
  );
  //OR U181bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U181bar (
    .O(ybar[168]),
    .I0(abar[10]),
    .I1(bbar[8])
  );
  //AND U182
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U182 (
    .O(y[167]),
    .I0(a[10]),
    .I1(b[7])
  );
  //OR U182bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U182bar (
    .O(ybar[167]),
    .I0(abar[10]),
    .I1(bbar[7])
  );
  //AND U183
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U183 (
    .O(y[166]),
    .I0(a[10]),
    .I1(b[6])
  );
  //OR U183bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U183bar (
    .O(ybar[166]),
    .I0(abar[10]),
    .I1(bbar[6])
  );
  //AND U184
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U184 (
    .O(y[165]),
    .I0(a[10]),
    .I1(b[5])
  );
  //OR U184bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U184bar (
    .O(ybar[165]),
    .I0(abar[10]),
    .I1(bbar[5])
  );
  //AND U185
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U185 (
    .O(y[164]),
    .I0(a[10]),
    .I1(b[4])
  );
  //OR U185bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U185bar (
    .O(ybar[164]),
    .I0(abar[10]),
    .I1(bbar[4])
  );
  //AND U186
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U186 (
    .O(y[163]),
    .I0(a[10]),
    .I1(b[3])
  );
  //OR U186bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U186bar (
    .O(ybar[163]),
    .I0(abar[10]),
    .I1(bbar[3])
  );
  //AND U187
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U187 (
    .O(y[162]),
    .I0(a[10]),
    .I1(b[2])
  );
  //OR U187bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U187bar (
    .O(ybar[162]),
    .I0(abar[10]),
    .I1(bbar[2])
  );
  //AND U188
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U188 (
    .O(y[161]),
    .I0(a[10]),
    .I1(b[1])
  );
  //OR U188bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U188bar (
    .O(ybar[161]),
    .I0(abar[10]),
    .I1(bbar[1])
  );
  //AND U189
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U189 (
    .O(y[160]),
    .I0(a[10]),
    .I1(b[0])
  );
  //OR U189bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U189bar (
    .O(ybar[160]),
    .I0(abar[10]),
    .I1(bbar[0])
  );
  //AND U190
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U190 (
    .O(y[15]),
    .I0(b[15]),
    .I1(a[0])
  );
  //OR U190bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U190bar (
    .O(ybar[15]),
    .I0(bbar[15]),
    .I1(abar[0])
  );
  //AND U191
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U191 (
    .O(y[159]),
    .I0(a[9]),
    .I1(b[15])
  );
  //OR U191bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U191bar (
    .O(ybar[159]),
    .I0(abar[9]),
    .I1(bbar[15])
  );
  //AND U192
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U192 (
    .O(y[158]),
    .I0(a[9]),
    .I1(b[14])
  );
  //OR U192bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U192bar (
    .O(ybar[158]),
    .I0(abar[9]),
    .I1(bbar[14])
  );
  //AND U193
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U193 (
    .O(y[157]),
    .I0(a[9]),
    .I1(b[13])
  );
  //OR U193bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U193bar (
    .O(ybar[157]),
    .I0(abar[9]),
    .I1(bbar[13])
  );
  //AND U194
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U194 (
    .O(y[156]),
    .I0(a[9]),
    .I1(b[12])
  );
  //OR U194bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U194bar (
    .O(ybar[156]),
    .I0(abar[9]),
    .I1(bbar[12])
  );
  //AND U195
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U195 (
    .O(y[155]),
    .I0(a[9]),
    .I1(b[11])
  );
  //OR U195bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U195bar (
    .O(ybar[155]),
    .I0(abar[9]),
    .I1(bbar[11])
  );
  //AND U196
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U196 (
    .O(y[154]),
    .I0(a[9]),
    .I1(b[10])
  );
  //OR U196bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U196bar (
    .O(ybar[154]),
    .I0(abar[9]),
    .I1(bbar[10])
  );
  //AND U197
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U197 (
    .O(y[153]),
    .I0(a[9]),
    .I1(b[9])
  );
  //OR U197bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U197bar (
    .O(ybar[153]),
    .I0(abar[9]),
    .I1(bbar[9])
  );
  //AND U198
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U198 (
    .O(y[152]),
    .I0(a[9]),
    .I1(b[8])
  );
  //OR U198bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U198bar (
    .O(ybar[152]),
    .I0(abar[9]),
    .I1(bbar[8])
  );
  //AND U199
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U199 (
    .O(y[151]),
    .I0(a[9]),
    .I1(b[7])
  );
  //OR U199bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U199bar (
    .O(ybar[151]),
    .I0(abar[9]),
    .I1(bbar[7])
  );
  //AND U200
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U200 (
    .O(y[150]),
    .I0(a[9]),
    .I1(b[6])
  );
  //OR U200bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U200bar (
    .O(ybar[150]),
    .I0(abar[9]),
    .I1(bbar[6])
  );
  //AND U201
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U201 (
    .O(y[14]),
    .I0(b[14]),
    .I1(a[0])
  );
  //OR U201bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U201bar (
    .O(ybar[14]),
    .I0(bbar[14]),
    .I1(abar[0])
  );
  //AND U202
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U202 (
    .O(y[149]),
    .I0(a[9]),
    .I1(b[5])
  );
  //OR U202bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U202bar (
    .O(ybar[149]),
    .I0(abar[9]),
    .I1(bbar[5])
  );
  //AND U203
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U203 (
    .O(y[148]),
    .I0(a[9]),
    .I1(b[4])
  );
  //OR U203bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U203bar (
    .O(ybar[148]),
    .I0(abar[9]),
    .I1(bbar[4])
  );
  //AND U204
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U204 (
    .O(y[147]),
    .I0(a[9]),
    .I1(b[3])
  );
  //OR U204bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U204bar (
    .O(ybar[147]),
    .I0(abar[9]),
    .I1(bbar[3])
  );
  //AND U205
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U205 (
    .O(y[146]),
    .I0(a[9]),
    .I1(b[2])
  );
  //OR U205bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U205bar (
    .O(ybar[146]),
    .I0(abar[9]),
    .I1(bbar[2])
  );
  //AND U206
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U206 (
    .O(y[145]),
    .I0(a[9]),
    .I1(b[1])
  );
  //OR U206bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U206bar (
    .O(ybar[145]),
    .I0(abar[9]),
    .I1(bbar[1])
  );
  //AND U207
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U207 (
    .O(y[144]),
    .I0(a[9]),
    .I1(b[0])
  );
  //OR U207bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U207bar (
    .O(ybar[144]),
    .I0(abar[9]),
    .I1(bbar[0])
  );
  //AND U208
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U208 (
    .O(y[143]),
    .I0(a[8]),
    .I1(b[15])
  );
  //OR U208bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U208bar (
    .O(ybar[143]),
    .I0(abar[8]),
    .I1(bbar[15])
  );
  //AND U209
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U209 (
    .O(y[142]),
    .I0(a[8]),
    .I1(b[14])
  );
  //OR U209bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U209bar (
    .O(ybar[142]),
    .I0(abar[8]),
    .I1(bbar[14])
  );
  //AND U210
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U210 (
    .O(y[141]),
    .I0(a[8]),
    .I1(b[13])
  );
  //OR U210bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U210bar (
    .O(ybar[141]),
    .I0(abar[8]),
    .I1(bbar[13])
  );
  //AND U211
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U211 (
    .O(y[140]),
    .I0(a[8]),
    .I1(b[12])
  );
  //OR U211bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U211bar (
    .O(ybar[140]),
    .I0(abar[8]),
    .I1(bbar[12])
  );
  //AND U212
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U212 (
    .O(y[13]),
    .I0(b[13]),
    .I1(a[0])
  );
  //OR U212bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U212bar (
    .O(ybar[13]),
    .I0(bbar[13]),
    .I1(abar[0])
  );
  //AND U213
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U213 (
    .O(y[139]),
    .I0(a[8]),
    .I1(b[11])
  );
  //OR U213bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U213bar (
    .O(ybar[139]),
    .I0(abar[8]),
    .I1(bbar[11])
  );
  //AND U214
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U214 (
    .O(y[138]),
    .I0(a[8]),
    .I1(b[10])
  );
  //OR U214bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U214bar (
    .O(ybar[138]),
    .I0(abar[8]),
    .I1(bbar[10])
  );
  //AND U215
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U215 (
    .O(y[137]),
    .I0(a[8]),
    .I1(b[9])
  );
  //OR U215bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U215bar (
    .O(ybar[137]),
    .I0(abar[8]),
    .I1(bbar[9])
  );
  //AND U216
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U216 (
    .O(y[136]),
    .I0(a[8]),
    .I1(b[8])
  );
  //OR U216bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U216bar (
    .O(ybar[136]),
    .I0(abar[8]),
    .I1(bbar[8])
  );
  //AND U217
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U217 (
    .O(y[135]),
    .I0(a[8]),
    .I1(b[7])
  );
  //OR U217bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U217bar (
    .O(ybar[135]),
    .I0(abar[8]),
    .I1(bbar[7])
  );
  //AND U218
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U218 (
    .O(y[134]),
    .I0(a[8]),
    .I1(b[6])
  );
  //OR U218bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U218bar (
    .O(ybar[134]),
    .I0(abar[8]),
    .I1(bbar[6])
  );
  //AND U219
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U219 (
    .O(y[133]),
    .I0(a[8]),
    .I1(b[5])
  );
  //OR U219bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U219bar (
    .O(ybar[133]),
    .I0(abar[8]),
    .I1(bbar[5])
  );
  //AND U220
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U220 (
    .O(y[132]),
    .I0(a[8]),
    .I1(b[4])
  );
  //OR U220bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U220bar (
    .O(ybar[132]),
    .I0(abar[8]),
    .I1(bbar[4])
  );
  //AND U221
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U221 (
    .O(y[131]),
    .I0(a[8]),
    .I1(b[3])
  );
  //OR U221bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U221bar (
    .O(ybar[131]),
    .I0(abar[8]),
    .I1(bbar[3])
  );
  //AND U222
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U222 (
    .O(y[130]),
    .I0(a[8]),
    .I1(b[2])
  );
  //OR U222bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U222bar (
    .O(ybar[130]),
    .I0(abar[8]),
    .I1(bbar[2])
  );
  //AND U223
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U223 (
    .O(y[12]),
    .I0(b[12]),
    .I1(a[0])
  );
  //OR U223bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U223bar (
    .O(ybar[12]),
    .I0(bbar[12]),
    .I1(abar[0])
  );
  //AND U224
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U224 (
    .O(y[129]),
    .I0(a[8]),
    .I1(b[1])
  );
  //OR U224bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U224bar (
    .O(ybar[129]),
    .I0(abar[8]),
    .I1(bbar[1])
  );
  //AND U225
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U225 (
    .O(y[128]),
    .I0(a[8]),
    .I1(b[0])
  );
  //OR U225bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U225bar (
    .O(ybar[128]),
    .I0(abar[8]),
    .I1(bbar[0])
  );
  //AND U226
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U226 (
    .O(y[127]),
    .I0(a[7]),
    .I1(b[15])
  );
  //OR U226bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U226bar (
    .O(ybar[127]),
    .I0(abar[7]),
    .I1(bbar[15])
  );
  //AND U227
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U227 (
    .O(y[126]),
    .I0(a[7]),
    .I1(b[14])
  );
  //OR U227bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U227bar (
    .O(ybar[126]),
    .I0(abar[7]),
    .I1(bbar[14])
  );
  //AND U228
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U228 (
    .O(y[125]),
    .I0(a[7]),
    .I1(b[13])
  );
  //OR U228bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U228bar (
    .O(ybar[125]),
    .I0(abar[7]),
    .I1(bbar[13])
  );
  //AND U229
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U229 (
    .O(y[124]),
    .I0(a[7]),
    .I1(b[12])
  );
  //OR U229bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U229bar (
    .O(ybar[124]),
    .I0(abar[7]),
    .I1(bbar[12])
  );
  //AND U230
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U230 (
    .O(y[123]),
    .I0(a[7]),
    .I1(b[11])
  );
  //OR U230bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U230bar (
    .O(ybar[123]),
    .I0(abar[7]),
    .I1(bbar[11])
  );
  //AND U231
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U231 (
    .O(y[122]),
    .I0(a[7]),
    .I1(b[10])
  );
  //OR U231bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U231bar (
    .O(ybar[122]),
    .I0(abar[7]),
    .I1(bbar[10])
  );
  //AND U232
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U232 (
    .O(y[121]),
    .I0(a[7]),
    .I1(b[9])
  );
  //OR U232bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U232bar (
    .O(ybar[121]),
    .I0(abar[7]),
    .I1(bbar[9])
  );
  //AND U233
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U233 (
    .O(y[120]),
    .I0(a[7]),
    .I1(b[8])
  );
  //OR U233bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U233bar (
    .O(ybar[120]),
    .I0(abar[7]),
    .I1(bbar[8])
  );
  //AND U234
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U234 (
    .O(y[11]),
    .I0(b[11]),
    .I1(a[0])
  );
  //OR U234bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U234bar (
    .O(ybar[11]),
    .I0(bbar[11]),
    .I1(abar[0])
  );
  //AND U235
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U235 (
    .O(y[119]),
    .I0(a[7]),
    .I1(b[7])
  );
  //OR U235bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U235bar (
    .O(ybar[119]),
    .I0(abar[7]),
    .I1(bbar[7])
  );
  //AND U236
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U236 (
    .O(y[118]),
    .I0(a[7]),
    .I1(b[6])
  );
  //OR U236bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U236bar (
    .O(ybar[118]),
    .I0(abar[7]),
    .I1(bbar[6])
  );
  //AND U237
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U237 (
    .O(y[117]),
    .I0(a[7]),
    .I1(b[5])
  );
  //OR U237bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U237bar (
    .O(ybar[117]),
    .I0(abar[7]),
    .I1(bbar[5])
  );
  //AND U238
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U238 (
    .O(y[116]),
    .I0(a[7]),
    .I1(b[4])
  );
  //OR U238bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U238bar (
    .O(ybar[116]),
    .I0(abar[7]),
    .I1(bbar[4])
  );
  //AND U239
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U239 (
    .O(y[115]),
    .I0(a[7]),
    .I1(b[3])
  );
  //OR U239bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U239bar (
    .O(ybar[115]),
    .I0(abar[7]),
    .I1(bbar[3])
  );
  //AND U240
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U240 (
    .O(y[114]),
    .I0(a[7]),
    .I1(b[2])
  );
  //OR U240bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U240bar (
    .O(ybar[114]),
    .I0(abar[7]),
    .I1(bbar[2])
  );
  //AND U241
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U241 (
    .O(y[113]),
    .I0(a[7]),
    .I1(b[1])
  );
  //OR U241bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U241bar (
    .O(ybar[113]),
    .I0(abar[7]),
    .I1(bbar[1])
  );
  //AND U242
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U242 (
    .O(y[112]),
    .I0(a[7]),
    .I1(b[0])
  );
  //OR U242bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U242bar (
    .O(ybar[112]),
    .I0(abar[7]),
    .I1(bbar[0])
  );
  //AND U243
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U243 (
    .O(y[111]),
    .I0(b[15]),
    .I1(a[6])
  );
  //OR U243bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U243bar (
    .O(ybar[111]),
    .I0(bbar[15]),
    .I1(abar[6])
  );
  //AND U244
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U244 (
    .O(y[110]),
    .I0(b[14]),
    .I1(a[6])
  );
  //OR U244bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U244bar (
    .O(ybar[110]),
    .I0(bbar[14]),
    .I1(abar[6])
  );
  //AND U245
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U245 (
    .O(y[10]),
    .I0(b[10]),
    .I1(a[0])
  );
  //OR U245bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U245bar (
    .O(ybar[10]),
    .I0(bbar[10]),
    .I1(abar[0])
  );
  //AND U246
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U246 (
    .O(y[109]),
    .I0(b[13]),
    .I1(a[6])
  );
  //OR U246bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U246bar (
    .O(ybar[109]),
    .I0(bbar[13]),
    .I1(abar[6])
  );
  //AND U247
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U247 (
    .O(y[108]),
    .I0(b[12]),
    .I1(a[6])
  );
  //OR U247bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U247bar (
    .O(ybar[108]),
    .I0(bbar[12]),
    .I1(abar[6])
  );
  //AND U248
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U248 (
    .O(y[107]),
    .I0(b[11]),
    .I1(a[6])
  );
  //OR U248bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U248bar (
    .O(ybar[107]),
    .I0(bbar[11]),
    .I1(abar[6])
  );
  //AND U249
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U249 (
    .O(y[106]),
    .I0(b[10]),
    .I1(a[6])
  );
  //OR U249bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U249bar (
    .O(ybar[106]),
    .I0(bbar[10]),
    .I1(abar[6])
  );
  //AND U250
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U250 (
    .O(y[105]),
    .I0(a[6]),
    .I1(b[9])
  );
  //OR U250bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U250bar (
    .O(ybar[105]),
    .I0(abar[6]),
    .I1(bbar[9])
  );
  //AND U251
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U251 (
    .O(y[104]),
    .I0(b[8]),
    .I1(a[6])
  );
  //OR U251bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U251bar (
    .O(ybar[104]),
    .I0(bbar[8]),
    .I1(abar[6])
  );
  //AND U252
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U252 (
    .O(y[103]),
    .I0(b[7]),
    .I1(a[6])
  );
  //OR U252bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U252bar (
    .O(ybar[103]),
    .I0(bbar[7]),
    .I1(abar[6])
  );
  //AND U253
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U253 (
    .O(y[102]),
    .I0(b[6]),
    .I1(a[6])
  );
  //OR U253bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U253bar (
    .O(ybar[102]),
    .I0(bbar[6]),
    .I1(abar[6])
  );
  //AND U254
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U254 (
    .O(y[101]),
    .I0(b[5]),
    .I1(a[6])
  );
  //OR U254bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U254bar (
    .O(ybar[101]),
    .I0(bbar[5]),
    .I1(abar[6])
  );
  //AND U255
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U255 (
    .O(y[100]),
    .I0(b[4]),
    .I1(a[6])
  );
  //OR U255bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U255bar (
    .O(ybar[100]),
    .I0(bbar[4]),
    .I1(abar[6])
  );
  //AND U256
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U256 (
    .O(y[0]),
    .I0(b[0]),
    .I1(a[0])
  );
  //OR U256bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U256bar (
    .O(ybar[0]),
    .I0(bbar[0]),
    .I1(abar[0])
  );
endmodule

module decode_13 ( in, out );

  input wire [7:0] in;
//input_done

  output wire [255:0] out;
//output_done

  wire [15:0] level1;
  wire [31:0] level2;
//wire_done

  CD2_52 cd_l1_1 ( .a(in[1]), .b(in[0]), .y(level1[3:0]) );
  CD2_51 cd_l1_2 ( .a(in[3]), .b(in[2]), .y(level1[7:4]) );
  CD2_50 cd_l1_3 ( .a(in[5]), .b(in[4]), .y(level1[11:8]) );
  CD2_49 cd_l1_4 ( .a(in[7]), .b(in[6]), .y(level1[15:12]) );
  CD4_26 cd_l2_1 ( .a(level1[7:4]), .b(level1[3:0]), .y(level2[15:0]) );
  CD4_25 cd_l2_2 ( .a(level1[15:12]), .b(level1[11:8]), .y(level2[31:16]) );
  CD16_13 cd_l3 ( .a(level2[31:16]), .b(level2[15:0]), .y(out) );
endmodule

module encode_13 ( in, out );

  input wire [255:0] in;
  wire [255:0] inbar;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
  assign inbar[8] = ~in[8];
  assign inbar[9] = ~in[9];
  assign inbar[10] = ~in[10];
  assign inbar[11] = ~in[11];
  assign inbar[12] = ~in[12];
  assign inbar[13] = ~in[13];
  assign inbar[14] = ~in[14];
  assign inbar[15] = ~in[15];
  assign inbar[16] = ~in[16];
  assign inbar[17] = ~in[17];
  assign inbar[18] = ~in[18];
  assign inbar[19] = ~in[19];
  assign inbar[20] = ~in[20];
  assign inbar[21] = ~in[21];
  assign inbar[22] = ~in[22];
  assign inbar[23] = ~in[23];
  assign inbar[24] = ~in[24];
  assign inbar[25] = ~in[25];
  assign inbar[26] = ~in[26];
  assign inbar[27] = ~in[27];
  assign inbar[28] = ~in[28];
  assign inbar[29] = ~in[29];
  assign inbar[30] = ~in[30];
  assign inbar[31] = ~in[31];
  assign inbar[32] = ~in[32];
  assign inbar[33] = ~in[33];
  assign inbar[34] = ~in[34];
  assign inbar[35] = ~in[35];
  assign inbar[36] = ~in[36];
  assign inbar[37] = ~in[37];
  assign inbar[38] = ~in[38];
  assign inbar[39] = ~in[39];
  assign inbar[40] = ~in[40];
  assign inbar[41] = ~in[41];
  assign inbar[42] = ~in[42];
  assign inbar[43] = ~in[43];
  assign inbar[44] = ~in[44];
  assign inbar[45] = ~in[45];
  assign inbar[46] = ~in[46];
  assign inbar[47] = ~in[47];
  assign inbar[48] = ~in[48];
  assign inbar[49] = ~in[49];
  assign inbar[50] = ~in[50];
  assign inbar[51] = ~in[51];
  assign inbar[52] = ~in[52];
  assign inbar[53] = ~in[53];
  assign inbar[54] = ~in[54];
  assign inbar[55] = ~in[55];
  assign inbar[56] = ~in[56];
  assign inbar[57] = ~in[57];
  assign inbar[58] = ~in[58];
  assign inbar[59] = ~in[59];
  assign inbar[60] = ~in[60];
  assign inbar[61] = ~in[61];
  assign inbar[62] = ~in[62];
  assign inbar[63] = ~in[63];
  assign inbar[64] = ~in[64];
  assign inbar[65] = ~in[65];
  assign inbar[66] = ~in[66];
  assign inbar[67] = ~in[67];
  assign inbar[68] = ~in[68];
  assign inbar[69] = ~in[69];
  assign inbar[70] = ~in[70];
  assign inbar[71] = ~in[71];
  assign inbar[72] = ~in[72];
  assign inbar[73] = ~in[73];
  assign inbar[74] = ~in[74];
  assign inbar[75] = ~in[75];
  assign inbar[76] = ~in[76];
  assign inbar[77] = ~in[77];
  assign inbar[78] = ~in[78];
  assign inbar[79] = ~in[79];
  assign inbar[80] = ~in[80];
  assign inbar[81] = ~in[81];
  assign inbar[82] = ~in[82];
  assign inbar[83] = ~in[83];
  assign inbar[84] = ~in[84];
  assign inbar[85] = ~in[85];
  assign inbar[86] = ~in[86];
  assign inbar[87] = ~in[87];
  assign inbar[88] = ~in[88];
  assign inbar[89] = ~in[89];
  assign inbar[90] = ~in[90];
  assign inbar[91] = ~in[91];
  assign inbar[92] = ~in[92];
  assign inbar[93] = ~in[93];
  assign inbar[94] = ~in[94];
  assign inbar[95] = ~in[95];
  assign inbar[96] = ~in[96];
  assign inbar[97] = ~in[97];
  assign inbar[98] = ~in[98];
  assign inbar[99] = ~in[99];
  assign inbar[100] = ~in[100];
  assign inbar[101] = ~in[101];
  assign inbar[102] = ~in[102];
  assign inbar[103] = ~in[103];
  assign inbar[104] = ~in[104];
  assign inbar[105] = ~in[105];
  assign inbar[106] = ~in[106];
  assign inbar[107] = ~in[107];
  assign inbar[108] = ~in[108];
  assign inbar[109] = ~in[109];
  assign inbar[110] = ~in[110];
  assign inbar[111] = ~in[111];
  assign inbar[112] = ~in[112];
  assign inbar[113] = ~in[113];
  assign inbar[114] = ~in[114];
  assign inbar[115] = ~in[115];
  assign inbar[116] = ~in[116];
  assign inbar[117] = ~in[117];
  assign inbar[118] = ~in[118];
  assign inbar[119] = ~in[119];
  assign inbar[120] = ~in[120];
  assign inbar[121] = ~in[121];
  assign inbar[122] = ~in[122];
  assign inbar[123] = ~in[123];
  assign inbar[124] = ~in[124];
  assign inbar[125] = ~in[125];
  assign inbar[126] = ~in[126];
  assign inbar[127] = ~in[127];
  assign inbar[128] = ~in[128];
  assign inbar[129] = ~in[129];
  assign inbar[130] = ~in[130];
  assign inbar[131] = ~in[131];
  assign inbar[132] = ~in[132];
  assign inbar[133] = ~in[133];
  assign inbar[134] = ~in[134];
  assign inbar[135] = ~in[135];
  assign inbar[136] = ~in[136];
  assign inbar[137] = ~in[137];
  assign inbar[138] = ~in[138];
  assign inbar[139] = ~in[139];
  assign inbar[140] = ~in[140];
  assign inbar[141] = ~in[141];
  assign inbar[142] = ~in[142];
  assign inbar[143] = ~in[143];
  assign inbar[144] = ~in[144];
  assign inbar[145] = ~in[145];
  assign inbar[146] = ~in[146];
  assign inbar[147] = ~in[147];
  assign inbar[148] = ~in[148];
  assign inbar[149] = ~in[149];
  assign inbar[150] = ~in[150];
  assign inbar[151] = ~in[151];
  assign inbar[152] = ~in[152];
  assign inbar[153] = ~in[153];
  assign inbar[154] = ~in[154];
  assign inbar[155] = ~in[155];
  assign inbar[156] = ~in[156];
  assign inbar[157] = ~in[157];
  assign inbar[158] = ~in[158];
  assign inbar[159] = ~in[159];
  assign inbar[160] = ~in[160];
  assign inbar[161] = ~in[161];
  assign inbar[162] = ~in[162];
  assign inbar[163] = ~in[163];
  assign inbar[164] = ~in[164];
  assign inbar[165] = ~in[165];
  assign inbar[166] = ~in[166];
  assign inbar[167] = ~in[167];
  assign inbar[168] = ~in[168];
  assign inbar[169] = ~in[169];
  assign inbar[170] = ~in[170];
  assign inbar[171] = ~in[171];
  assign inbar[172] = ~in[172];
  assign inbar[173] = ~in[173];
  assign inbar[174] = ~in[174];
  assign inbar[175] = ~in[175];
  assign inbar[176] = ~in[176];
  assign inbar[177] = ~in[177];
  assign inbar[178] = ~in[178];
  assign inbar[179] = ~in[179];
  assign inbar[180] = ~in[180];
  assign inbar[181] = ~in[181];
  assign inbar[182] = ~in[182];
  assign inbar[183] = ~in[183];
  assign inbar[184] = ~in[184];
  assign inbar[185] = ~in[185];
  assign inbar[186] = ~in[186];
  assign inbar[187] = ~in[187];
  assign inbar[188] = ~in[188];
  assign inbar[189] = ~in[189];
  assign inbar[190] = ~in[190];
  assign inbar[191] = ~in[191];
  assign inbar[192] = ~in[192];
  assign inbar[193] = ~in[193];
  assign inbar[194] = ~in[194];
  assign inbar[195] = ~in[195];
  assign inbar[196] = ~in[196];
  assign inbar[197] = ~in[197];
  assign inbar[198] = ~in[198];
  assign inbar[199] = ~in[199];
  assign inbar[200] = ~in[200];
  assign inbar[201] = ~in[201];
  assign inbar[202] = ~in[202];
  assign inbar[203] = ~in[203];
  assign inbar[204] = ~in[204];
  assign inbar[205] = ~in[205];
  assign inbar[206] = ~in[206];
  assign inbar[207] = ~in[207];
  assign inbar[208] = ~in[208];
  assign inbar[209] = ~in[209];
  assign inbar[210] = ~in[210];
  assign inbar[211] = ~in[211];
  assign inbar[212] = ~in[212];
  assign inbar[213] = ~in[213];
  assign inbar[214] = ~in[214];
  assign inbar[215] = ~in[215];
  assign inbar[216] = ~in[216];
  assign inbar[217] = ~in[217];
  assign inbar[218] = ~in[218];
  assign inbar[219] = ~in[219];
  assign inbar[220] = ~in[220];
  assign inbar[221] = ~in[221];
  assign inbar[222] = ~in[222];
  assign inbar[223] = ~in[223];
  assign inbar[224] = ~in[224];
  assign inbar[225] = ~in[225];
  assign inbar[226] = ~in[226];
  assign inbar[227] = ~in[227];
  assign inbar[228] = ~in[228];
  assign inbar[229] = ~in[229];
  assign inbar[230] = ~in[230];
  assign inbar[231] = ~in[231];
  assign inbar[232] = ~in[232];
  assign inbar[233] = ~in[233];
  assign inbar[234] = ~in[234];
  assign inbar[235] = ~in[235];
  assign inbar[236] = ~in[236];
  assign inbar[237] = ~in[237];
  assign inbar[238] = ~in[238];
  assign inbar[239] = ~in[239];
  assign inbar[240] = ~in[240];
  assign inbar[241] = ~in[241];
  assign inbar[242] = ~in[242];
  assign inbar[243] = ~in[243];
  assign inbar[244] = ~in[244];
  assign inbar[245] = ~in[245];
  assign inbar[246] = ~in[246];
  assign inbar[247] = ~in[247];
  assign inbar[248] = ~in[248];
  assign inbar[249] = ~in[249];
  assign inbar[250] = ~in[250];
  assign inbar[251] = ~in[251];
  assign inbar[252] = ~in[252];
  assign inbar[253] = ~in[253];
  assign inbar[254] = ~in[254];
  assign inbar[255] = ~in[255];
//input_done

  output wire [7:0] out;
  wire [7:0] outbar;
//output_done

  wire in_81;
  wire in_80;
  wire in_79;
  wire in_78;
  wire in_77;
  wire in_76;
  wire in_75;
  wire in_74;
  wire in_73;
  wire in_72;
  wire in_71;
  wire in_70;
  wire in_69;
  wire in_68;
  wire in_67;
  wire in_66;
  wire in_65;
  wire in_64;
  wire in_63;
  wire in_62;
  wire in_61;
  wire in_60;
  wire in_59;
  wire in_58;
  wire in_57;
  wire in_56;
  wire in_55;
  wire in_54;
  wire in_53;
  wire in_52;
  wire in_51;
  wire in_50;
  wire in_49;
  wire in_48;
  wire in_47;
  wire in_46;
  wire in_45;
  wire in_44;
  wire in_43;
  wire in_42;
  wire in_41;
  wire in_40;
  wire in_39;
  wire in_38;
  wire in_37;
  wire in_36;
  wire in_35;
  wire in_34;
  wire in_33;
  wire in_32;
  wire in_31;
  wire in_30;
  wire in_29;
  wire in_28;
  wire in_27;
  wire in_26;
  wire in_25;
  wire in_24;
  wire in_23;
  wire in_22;
  wire in_21;
  wire in_20;
  wire in_19;
  wire in_18;
  wire in_17;
  wire in_16;
  wire in_15;
  wire in_14;
  wire in_13;
  wire in_12;
  wire in_11;
  wire in_10;
  wire in_9;
  wire in_8;
  wire in_7;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_3;
  wire in_2;
  wire in_1;
  wire in_0;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire in_81bar;
  wire in_80bar;
  wire in_79bar;
  wire in_78bar;
  wire in_77bar;
  wire in_76bar;
  wire in_75bar;
  wire in_74bar;
  wire in_73bar;
  wire in_72bar;
  wire in_71bar;
  wire in_70bar;
  wire in_69bar;
  wire in_68bar;
  wire in_67bar;
  wire in_66bar;
  wire in_65bar;
  wire in_64bar;
  wire in_63bar;
  wire in_62bar;
  wire in_61bar;
  wire in_60bar;
  wire in_59bar;
  wire in_58bar;
  wire in_57bar;
  wire in_56bar;
  wire in_55bar;
  wire in_54bar;
  wire in_53bar;
  wire in_52bar;
  wire in_51bar;
  wire in_50bar;
  wire in_49bar;
  wire in_48bar;
  wire in_47bar;
  wire in_46bar;
  wire in_45bar;
  wire in_44bar;
  wire in_43bar;
  wire in_42bar;
  wire in_41bar;
  wire in_40bar;
  wire in_39bar;
  wire in_38bar;
  wire in_37bar;
  wire in_36bar;
  wire in_35bar;
  wire in_34bar;
  wire in_33bar;
  wire in_32bar;
  wire in_31bar;
  wire in_30bar;
  wire in_29bar;
  wire in_28bar;
  wire in_27bar;
  wire in_26bar;
  wire in_25bar;
  wire in_24bar;
  wire in_23bar;
  wire in_22bar;
  wire in_21bar;
  wire in_20bar;
  wire in_19bar;
  wire in_18bar;
  wire in_17bar;
  wire in_16bar;
  wire in_15bar;
  wire in_14bar;
  wire in_13bar;
  wire in_12bar;
  wire in_11bar;
  wire in_10bar;
  wire in_9bar;
  wire in_8bar;
  wire in_7bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_3bar;
  wire in_2bar;
  wire in_1bar;
  wire in_0bar;
  wire n487bar;
  wire n488bar;
  wire n489bar;
  wire n490bar;
  wire n491bar;
  wire n492bar;
  wire n493bar;
  wire n494bar;
  wire n495bar;
  wire n496bar;
  wire n497bar;
  wire n498bar;
  wire n499bar;
  wire n500bar;
  wire n501bar;
  wire n502bar;
  wire n503bar;
  wire n504bar;
  wire n505bar;
  wire n506bar;
  wire n507bar;
  wire n508bar;
  wire n509bar;
  wire n510bar;
  wire n511bar;
  wire n512bar;
  wire n513bar;
  wire n514bar;
  wire n515bar;
  wire n516bar;
  wire n517bar;
  wire n518bar;
  wire n519bar;
  wire n520bar;
  wire n521bar;
  wire n522bar;
  wire n523bar;
  wire n524bar;
  wire n525bar;
  wire n526bar;
  wire n527bar;
  wire n528bar;
  wire n529bar;
  wire n530bar;
  wire n531bar;
  wire n532bar;
  wire n533bar;
  wire n534bar;
  wire n535bar;
  wire n536bar;
  wire n537bar;
  wire n538bar;
  wire n539bar;
  wire n540bar;
  wire n541bar;
  wire n542bar;
  wire n543bar;
  wire n544bar;
  wire n545bar;
  wire n546bar;
  wire n547bar;
  wire n548bar;
  wire n549bar;
  wire n550bar;
  wire n551bar;
  wire n552bar;
  wire n553bar;
  wire n554bar;
  wire n555bar;
  wire n556bar;
  wire n557bar;
  wire n558bar;
  wire n559bar;
  wire n560bar;
  wire n561bar;
  wire n562bar;
  wire n563bar;
  wire n564bar;
  wire n565bar;
  wire n566bar;
  wire n567bar;
  wire n568bar;
  wire n569bar;
  wire n570bar;
  wire n571bar;
  wire n572bar;
  wire n573bar;
  wire n574bar;
  wire n575bar;
  wire n576bar;
  wire n577bar;
  wire n578bar;
  wire n579bar;
  wire n580bar;
  wire n581bar;
  wire n582bar;
  wire n583bar;
  wire n584bar;
  wire n585bar;
  wire n586bar;
  wire n587bar;
  wire n588bar;
  wire n589bar;
  wire n590bar;
  wire n591bar;
  wire n592bar;
  wire n593bar;
  wire n594bar;
  wire n595bar;
  wire n596bar;
  wire n597bar;
  wire n598bar;
  wire n599bar;
  wire n600bar;
  wire n601bar;
  wire n602bar;
  wire n603bar;
  wire n604bar;
  wire n605bar;
  wire n606bar;
  wire n607bar;
  wire n608bar;
  wire n609bar;
  wire n610bar;
  wire n611bar;
  wire n612bar;
  wire n613bar;
  wire n614bar;
  wire n615bar;
  wire n616bar;
  wire n617bar;
  wire n618bar;
  wire n619bar;
  wire n620bar;
  wire n621bar;
  wire n622bar;
  wire n623bar;
  wire n624bar;
  wire n625bar;
  wire n626bar;
  wire n627bar;
  wire n628bar;
  wire n629bar;
  wire n630bar;
  wire n631bar;
  wire n632bar;
  wire n633bar;
  wire n634bar;
  wire n635bar;
  wire n636bar;
  wire n637bar;
  wire n638bar;
  wire n639bar;
  wire n640bar;
  wire n641bar;
  wire n642bar;
  wire n643bar;
  wire n644bar;
  wire n645bar;
  wire n646bar;
  wire n647bar;
  wire n648bar;
  wire n649bar;
  wire n650bar;
  wire n651bar;
  wire n652bar;
  wire n653bar;
  wire n654bar;
  wire n655bar;
  wire n656bar;
  wire n657bar;
  wire n658bar;
  wire n659bar;
  wire n660bar;
  wire n661bar;
  wire n662bar;
  wire n663bar;
  wire n664bar;
  wire n665bar;
  wire n666bar;
  wire n667bar;
  wire n668bar;
  wire n669bar;
  wire n670bar;
  wire n671bar;
  wire n672bar;
  wire n673bar;
  wire n674bar;
  wire n675bar;
  wire n676bar;
  wire n677bar;
  wire n678bar;
  wire n679bar;
  wire n680bar;
  wire n681bar;
  wire n682bar;
  wire n683bar;
  wire n684bar;
  wire n685bar;
  wire n686bar;
  wire n687bar;
  wire n688bar;
  wire n689bar;
  wire n690bar;
  wire n691bar;
  wire n692bar;
  wire n693bar;
  wire n694bar;
  wire n695bar;
  wire n696bar;
  wire n697bar;
  wire n698bar;
  wire n699bar;
  wire n700bar;
  wire n701bar;
  wire n702bar;
  wire n703bar;
  wire n704bar;
  wire n705bar;
  wire n706bar;
  wire n707bar;
  wire n708bar;
  wire n709bar;
  wire n710bar;
  wire n711bar;
  wire n712bar;
  wire n713bar;
  wire n714bar;
  wire n715bar;
  wire n716bar;
  wire n717bar;
  wire n718bar;
  wire n719bar;
  wire n720bar;
  wire n721bar;
  wire n722bar;
  wire n723bar;
  wire n724bar;
  wire n725bar;
  wire n726bar;
  wire n727bar;
  wire n728bar;
  wire n729bar;
  wire n730bar;
  wire n731bar;
  wire n732bar;
  wire n733bar;
  wire n734bar;
  wire n735bar;
  wire n736bar;
  wire n737bar;
  wire n738bar;
  wire n739bar;
  wire n740bar;
  wire n741bar;
  wire n742bar;
  wire n743bar;
  wire n744bar;
  wire n745bar;
  wire n746bar;
  wire n747bar;
  wire n748bar;
  wire n749bar;
  wire n750bar;
  wire n751bar;
  wire n752bar;
  wire n753bar;
  wire n754bar;
  wire n755bar;
  wire n756bar;
  wire n757bar;
  wire n758bar;
  wire n759bar;
  wire n760bar;
  wire n761bar;
  wire n762bar;
  wire n763bar;
  wire n764bar;
  wire n765bar;
  wire n766bar;
  wire n767bar;
  wire n768bar;
  wire n769bar;
  wire n770bar;
  wire n771bar;
  wire n772bar;
  wire n773bar;
  wire n774bar;
  wire n775bar;
  wire n776bar;
  wire n777bar;
  wire n778bar;
  wire n779bar;
  wire n780bar;
  wire n781bar;
  wire n782bar;
  wire n783bar;
  wire n784bar;
  wire n785bar;
  wire n786bar;
  wire n787bar;
  wire n788bar;
  wire n789bar;
  wire n790bar;
  wire n791bar;
  wire n792bar;
  wire n793bar;
  wire n794bar;
  wire n795bar;
  wire n796bar;
  wire n797bar;
  wire n798bar;
  wire n799bar;
  wire n800bar;
  wire n801bar;
  wire n802bar;
  wire n803bar;
  wire n804bar;
  wire n805bar;
  wire n806bar;
  wire n807bar;
  wire n808bar;
  wire n809bar;
  wire n810bar;
  wire n811bar;
  wire n812bar;
  wire n813bar;
  wire n814bar;
  wire n815bar;
  wire n816bar;
  wire n817bar;
  wire n818bar;
  wire n819bar;
  wire n820bar;
  wire n821bar;
  wire n822bar;
  wire n823bar;
  wire n824bar;
  wire n825bar;
  wire n826bar;
  wire n827bar;
  wire n828bar;
  wire n829bar;
  wire n830bar;
  wire n831bar;
  wire n832bar;
  wire n833bar;
  wire n834bar;
  wire n835bar;
  wire n836bar;
  wire n837bar;
  wire n838bar;
  wire n839bar;
  wire n840bar;
  wire n841bar;
  wire n842bar;
  wire n843bar;
  wire n844bar;
  wire n845bar;
  wire n846bar;
  wire n847bar;
  wire n848bar;
  wire n849bar;
  wire n850bar;
  wire n851bar;
  wire n852bar;
  wire n853bar;
  wire n854bar;
  wire n855bar;
  wire n856bar;
  wire n857bar;
  wire n858bar;
  wire n859bar;
  wire n860bar;
  wire n861bar;
  wire n862bar;
  wire n863bar;
  wire n864bar;
  wire n865bar;
  wire n866bar;
  wire n867bar;
  wire n868bar;
  wire n869bar;
  wire n870bar;
  wire n871bar;
  wire n872bar;
  wire n873bar;
  wire n874bar;
  wire n875bar;
  wire n876bar;
  wire n877bar;
  wire n878bar;
  wire n879bar;
  wire n880bar;
  wire n881bar;
  wire n882bar;
  wire n883bar;
  wire n884bar;
  wire n885bar;
  wire n886bar;
  wire n887bar;
  wire n888bar;
  wire n889bar;
  wire n890bar;
  wire n891bar;
  wire n892bar;
  wire n893bar;
  wire n894bar;
  wire n895bar;
  wire n896bar;
  wire n897bar;
  wire n898bar;
  wire n899bar;
  wire n900bar;
  wire n901bar;
  wire n902bar;
  wire n903bar;
  wire n904bar;
  wire n905bar;
  wire n906bar;
  wire n907bar;
  wire n908bar;
  wire n909bar;
  wire n910bar;
  wire n911bar;
  wire n912bar;
  wire n913bar;
  wire n914bar;
  wire n915bar;
  wire n916bar;
  wire n917bar;
  wire n918bar;
  wire n919bar;
  wire n920bar;
  wire n921bar;
  wire n922bar;
  wire n923bar;
  wire n924bar;
  wire n925bar;
  wire n926bar;
  wire n927bar;
  wire n928bar;
  wire n929bar;
  wire n930bar;
  wire n931bar;
  wire n932bar;
  wire n933bar;
  wire n934bar;
  wire n935bar;
  wire n936bar;
  wire n937bar;
  wire n938bar;
  wire n939bar;
  wire n940bar;
  wire n941bar;
  wire n942bar;
  wire n943bar;
  wire n944bar;
  wire n945bar;
  wire n946bar;
  wire n947bar;
  wire n948bar;
  wire n949bar;
  wire n950bar;
  wire n951bar;
  wire n952bar;
  wire n953bar;
  wire n954bar;
  wire n955bar;
  wire n956bar;
  wire n957bar;
  wire n958bar;
  wire n959bar;
  wire n960bar;
  wire n961bar;
  wire n962bar;
  wire n963bar;
  wire n964bar;
  wire n965bar;
  wire n966bar;
  wire n967bar;
  wire n968bar;
  wire n969bar;
  wire n970bar;
  wire n971bar;
  wire n972bar;
//wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];
  //OR U1
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1 (
    .O(out[7]),
    .I0(n972),
    .I1(n971)
  );
  //AND U1bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1bar (
    .O(outbar[7]),
    .I0(n972bar),
    .I1(n971bar)
  );
  //OR U2
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2 (
    .O(n971),
    .I0(n970),
    .I1(n969)
  );
  //AND U2bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2bar (
    .O(n971bar),
    .I0(n970bar),
    .I1(n969bar)
  );
  //OR U3
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3 (
    .O(n969),
    .I0(n968),
    .I1(n967)
  );
  //AND U3bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3bar (
    .O(n969bar),
    .I0(n968bar),
    .I1(n967bar)
  );
  //OR U4
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4 (
    .O(n967),
    .I0(n966),
    .I1(n965)
  );
  //AND U4bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4bar (
    .O(n967bar),
    .I0(n966bar),
    .I1(n965bar)
  );
  //OR U5
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5 (
    .O(n968),
    .I0(n964),
    .I1(n963)
  );
  //AND U5bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5bar (
    .O(n968bar),
    .I0(n964bar),
    .I1(n963bar)
  );
  //OR U6
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6 (
    .O(n963),
    .I0(in[116]),
    .I1(n962)
  );
  //AND U6bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6bar (
    .O(n963bar),
    .I0(inbar[116]),
    .I1(n962bar)
  );
  //OR U7
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7 (
    .O(n970),
    .I0(n961),
    .I1(n960)
  );
  //AND U7bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7bar (
    .O(n970bar),
    .I0(n961bar),
    .I1(n960bar)
  );
  //OR U8
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8 (
    .O(n960),
    .I0(in[150]),
    .I1(in[127])
  );
  //AND U8bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8bar (
    .O(n960bar),
    .I0(inbar[150]),
    .I1(inbar[127])
  );
  //OR U9
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9 (
    .O(n961),
    .I0(in[160]),
    .I1(n959)
  );
  //AND U9bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9bar (
    .O(n961bar),
    .I0(inbar[160]),
    .I1(n959bar)
  );
  //OR U10
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10 (
    .O(n959),
    .I0(in[252]),
    .I1(in[168])
  );
  //AND U10bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10bar (
    .O(n959bar),
    .I0(inbar[252]),
    .I1(inbar[168])
  );
  //OR U11
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11 (
    .O(n972),
    .I0(n958),
    .I1(n957)
  );
  //AND U11bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11bar (
    .O(n972bar),
    .I0(n958bar),
    .I1(n957bar)
  );
  //OR U12
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12 (
    .O(n957),
    .I0(n956),
    .I1(n955)
  );
  //AND U12bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12bar (
    .O(n957bar),
    .I0(n956bar),
    .I1(n955bar)
  );
  //OR U13
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13 (
    .O(n955),
    .I0(in_17),
    .I1(in[96])
  );
  //AND U13bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13bar (
    .O(n955bar),
    .I0(in_17bar),
    .I1(inbar[96])
  );
  //OR U14
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14 (
    .O(n956),
    .I0(in_23),
    .I1(n954)
  );
  //AND U14bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14bar (
    .O(n956bar),
    .I0(in_23bar),
    .I1(n954bar)
  );
  //OR U15
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15 (
    .O(n954),
    .I0(in_31),
    .I1(in_26)
  );
  //AND U15bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15bar (
    .O(n954bar),
    .I0(in_31bar),
    .I1(in_26bar)
  );
  //OR U16
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16 (
    .O(n958),
    .I0(n953),
    .I1(n952)
  );
  //AND U16bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16bar (
    .O(n958bar),
    .I0(n953bar),
    .I1(n952bar)
  );
  //OR U17
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U17 (
    .O(n952),
    .I0(in_58),
    .I1(in_4)
  );
  //AND U17bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U17bar (
    .O(n952bar),
    .I0(in_58bar),
    .I1(in_4bar)
  );
  //OR U18
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U18 (
    .O(n953),
    .I0(in_59),
    .I1(n951)
  );
  //AND U18bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U18bar (
    .O(n953bar),
    .I0(in_59bar),
    .I1(n951bar)
  );
  //OR U19
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U19 (
    .O(n951),
    .I0(in_71),
    .I1(in_62)
  );
  //AND U19bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U19bar (
    .O(n951bar),
    .I0(in_71bar),
    .I1(in_62bar)
  );
  //OR U20
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U20 (
    .O(out[6]),
    .I0(n950),
    .I1(n949)
  );
  //AND U20bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U20bar (
    .O(outbar[6]),
    .I0(n950bar),
    .I1(n949bar)
  );
  //OR U21
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U21 (
    .O(n949),
    .I0(n948),
    .I1(n947)
  );
  //AND U21bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U21bar (
    .O(n949bar),
    .I0(n948bar),
    .I1(n947bar)
  );
  //OR U22
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U22 (
    .O(n947),
    .I0(n946),
    .I1(n945)
  );
  //AND U22bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U22bar (
    .O(n947bar),
    .I0(n946bar),
    .I1(n945bar)
  );
  //OR U23
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U23 (
    .O(n945),
    .I0(n944),
    .I1(n943)
  );
  //AND U23bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U23bar (
    .O(n945bar),
    .I0(n944bar),
    .I1(n943bar)
  );
  //OR U24
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U24 (
    .O(n946),
    .I0(n942),
    .I1(n941)
  );
  //AND U24bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U24bar (
    .O(n946bar),
    .I0(n942bar),
    .I1(n941bar)
  );
  //OR U25
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U25 (
    .O(n941),
    .I0(in[101]),
    .I1(n940)
  );
  //AND U25bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U25bar (
    .O(n941bar),
    .I0(inbar[101]),
    .I1(n940bar)
  );
  //OR U26
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U26 (
    .O(n948),
    .I0(n939),
    .I1(n938)
  );
  //AND U26bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U26bar (
    .O(n948bar),
    .I0(n939bar),
    .I1(n938bar)
  );
  //OR U27
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U27 (
    .O(n938),
    .I0(in[114]),
    .I1(in[104])
  );
  //AND U27bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U27bar (
    .O(n938bar),
    .I0(inbar[114]),
    .I1(inbar[104])
  );
  //OR U28
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U28 (
    .O(n939),
    .I0(in[128]),
    .I1(n937)
  );
  //AND U28bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U28bar (
    .O(n939bar),
    .I0(inbar[128]),
    .I1(n937bar)
  );
  //OR U29
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U29 (
    .O(n937),
    .I0(in[136]),
    .I1(in[134])
  );
  //AND U29bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U29bar (
    .O(n937bar),
    .I0(inbar[136]),
    .I1(inbar[134])
  );
  //OR U30
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U30 (
    .O(n950),
    .I0(n936),
    .I1(n935)
  );
  //AND U30bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U30bar (
    .O(n950bar),
    .I0(n936bar),
    .I1(n935bar)
  );
  //OR U31
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U31 (
    .O(n935),
    .I0(n934),
    .I1(n933)
  );
  //AND U31bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U31bar (
    .O(n935bar),
    .I0(n934bar),
    .I1(n933bar)
  );
  //OR U32
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U32 (
    .O(n933),
    .I0(in[177]),
    .I1(in[164])
  );
  //AND U32bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U32bar (
    .O(n933bar),
    .I0(inbar[177]),
    .I1(inbar[164])
  );
  //OR U33
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U33 (
    .O(n934),
    .I0(in[212]),
    .I1(n932)
  );
  //AND U33bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U33bar (
    .O(n934bar),
    .I0(inbar[212]),
    .I1(n932bar)
  );
  //OR U34
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U34 (
    .O(n932),
    .I0(in[248]),
    .I1(in[221])
  );
  //AND U34bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U34bar (
    .O(n932bar),
    .I0(inbar[248]),
    .I1(inbar[221])
  );
  //OR U35
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U35 (
    .O(n936),
    .I0(n931),
    .I1(n930)
  );
  //AND U35bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U35bar (
    .O(n936bar),
    .I0(n931bar),
    .I1(n930bar)
  );
  //OR U36
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U36 (
    .O(n930),
    .I0(in_18),
    .I1(in[93])
  );
  //AND U36bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U36bar (
    .O(n930bar),
    .I0(in_18bar),
    .I1(inbar[93])
  );
  //OR U37
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U37 (
    .O(n931),
    .I0(in_31),
    .I1(n929)
  );
  //AND U37bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U37bar (
    .O(n931bar),
    .I0(in_31bar),
    .I1(n929bar)
  );
  //OR U38
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U38 (
    .O(n929),
    .I0(in_7),
    .I1(in_39)
  );
  //AND U38bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U38bar (
    .O(n929bar),
    .I0(in_7bar),
    .I1(in_39bar)
  );
  //OR U39
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U39 (
    .O(out[5]),
    .I0(n928),
    .I1(n927)
  );
  //AND U39bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U39bar (
    .O(outbar[5]),
    .I0(n928bar),
    .I1(n927bar)
  );
  //OR U40
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U40 (
    .O(n927),
    .I0(n926),
    .I1(n925)
  );
  //AND U40bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U40bar (
    .O(n927bar),
    .I0(n926bar),
    .I1(n925bar)
  );
  //OR U41
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U41 (
    .O(n925),
    .I0(n924),
    .I1(n923)
  );
  //AND U41bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U41bar (
    .O(n925bar),
    .I0(n924bar),
    .I1(n923bar)
  );
  //OR U42
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U42 (
    .O(n923),
    .I0(n922),
    .I1(n921)
  );
  //AND U42bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U42bar (
    .O(n923bar),
    .I0(n922bar),
    .I1(n921bar)
  );
  //OR U43
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U43 (
    .O(n924),
    .I0(n940),
    .I1(n920)
  );
  //AND U43bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U43bar (
    .O(n924bar),
    .I0(n940bar),
    .I1(n920bar)
  );
  //OR U44
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U44 (
    .O(n920),
    .I0(in[111]),
    .I1(n919)
  );
  //AND U44bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U44bar (
    .O(n920bar),
    .I0(inbar[111]),
    .I1(n919bar)
  );
  //OR U45
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U45 (
    .O(n940),
    .I0(n918),
    .I1(n917)
  );
  //AND U45bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U45bar (
    .O(n940bar),
    .I0(n918bar),
    .I1(n917bar)
  );
  //OR U46
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U46 (
    .O(n917),
    .I0(n916),
    .I1(n915)
  );
  //AND U46bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U46bar (
    .O(n917bar),
    .I0(n916bar),
    .I1(n915bar)
  );
  //OR U47
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U47 (
    .O(n915),
    .I0(n914),
    .I1(n913)
  );
  //AND U47bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U47bar (
    .O(n915bar),
    .I0(n914bar),
    .I1(n913bar)
  );
  //OR U48
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U48 (
    .O(n913),
    .I0(in[140]),
    .I1(in[131])
  );
  //AND U48bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U48bar (
    .O(n913bar),
    .I0(inbar[140]),
    .I1(inbar[131])
  );
  //OR U49
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U49 (
    .O(n914),
    .I0(in[160]),
    .I1(in[144])
  );
  //AND U49bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U49bar (
    .O(n914bar),
    .I0(inbar[160]),
    .I1(inbar[144])
  );
  //OR U50
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U50 (
    .O(n916),
    .I0(n912),
    .I1(n911)
  );
  //AND U50bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U50bar (
    .O(n916bar),
    .I0(n912bar),
    .I1(n911bar)
  );
  //OR U51
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U51 (
    .O(n911),
    .I0(in[179]),
    .I1(in[174])
  );
  //AND U51bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U51bar (
    .O(n911bar),
    .I0(inbar[179]),
    .I1(inbar[174])
  );
  //OR U52
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U52 (
    .O(n912),
    .I0(in[188]),
    .I1(in[184])
  );
  //AND U52bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U52bar (
    .O(n912bar),
    .I0(inbar[188]),
    .I1(inbar[184])
  );
  //OR U53
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U53 (
    .O(n918),
    .I0(n910),
    .I1(n909)
  );
  //AND U53bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U53bar (
    .O(n918bar),
    .I0(n910bar),
    .I1(n909bar)
  );
  //OR U54
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U54 (
    .O(n909),
    .I0(n908),
    .I1(n907)
  );
  //AND U54bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U54bar (
    .O(n909bar),
    .I0(n908bar),
    .I1(n907bar)
  );
  //OR U55
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U55 (
    .O(n907),
    .I0(in[216]),
    .I1(in[200])
  );
  //AND U55bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U55bar (
    .O(n907bar),
    .I0(inbar[216]),
    .I1(inbar[200])
  );
  //OR U56
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U56 (
    .O(n908),
    .I0(in[228]),
    .I1(in[224])
  );
  //AND U56bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U56bar (
    .O(n908bar),
    .I0(inbar[228]),
    .I1(inbar[224])
  );
  //OR U57
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U57 (
    .O(n910),
    .I0(n906),
    .I1(n905)
  );
  //AND U57bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U57bar (
    .O(n910bar),
    .I0(n906bar),
    .I1(n905bar)
  );
  //OR U58
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U58 (
    .O(n905),
    .I0(in[247]),
    .I1(in[235])
  );
  //AND U58bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U58bar (
    .O(n905bar),
    .I0(inbar[247]),
    .I1(inbar[235])
  );
  //OR U59
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U59 (
    .O(n906),
    .I0(in_42),
    .I1(in[83])
  );
  //AND U59bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U59bar (
    .O(n906bar),
    .I0(in_42bar),
    .I1(inbar[83])
  );
  //OR U60
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U60 (
    .O(n926),
    .I0(n904),
    .I1(n903)
  );
  //AND U60bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U60bar (
    .O(n926bar),
    .I0(n904bar),
    .I1(n903bar)
  );
  //OR U61
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U61 (
    .O(n903),
    .I0(in[166]),
    .I1(in[123])
  );
  //AND U61bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U61bar (
    .O(n903bar),
    .I0(inbar[166]),
    .I1(inbar[123])
  );
  //OR U62
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U62 (
    .O(n904),
    .I0(in[170]),
    .I1(n902)
  );
  //AND U62bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U62bar (
    .O(n904bar),
    .I0(inbar[170]),
    .I1(n902bar)
  );
  //OR U63
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U63 (
    .O(n902),
    .I0(in[194]),
    .I1(in[183])
  );
  //AND U63bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U63bar (
    .O(n902bar),
    .I0(inbar[194]),
    .I1(inbar[183])
  );
  //OR U64
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U64 (
    .O(n928),
    .I0(n901),
    .I1(n900)
  );
  //AND U64bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U64bar (
    .O(n928bar),
    .I0(n901bar),
    .I1(n900bar)
  );
  //OR U65
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U65 (
    .O(n900),
    .I0(n899),
    .I1(n898)
  );
  //AND U65bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U65bar (
    .O(n900bar),
    .I0(n899bar),
    .I1(n898bar)
  );
  //OR U66
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U66 (
    .O(n898),
    .I0(in[241]),
    .I1(in[238])
  );
  //AND U66bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U66bar (
    .O(n898bar),
    .I0(inbar[241]),
    .I1(inbar[238])
  );
  //OR U67
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U67 (
    .O(n899),
    .I0(in[250]),
    .I1(n897)
  );
  //AND U67bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U67bar (
    .O(n899bar),
    .I0(inbar[250]),
    .I1(n897bar)
  );
  //OR U68
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U68 (
    .O(n897),
    .I0(in_24),
    .I1(in[84])
  );
  //AND U68bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U68bar (
    .O(n897bar),
    .I0(in_24bar),
    .I1(inbar[84])
  );
  //OR U69
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U69 (
    .O(n901),
    .I0(n896),
    .I1(n895)
  );
  //AND U69bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U69bar (
    .O(n901bar),
    .I0(n896bar),
    .I1(n895bar)
  );
  //OR U70
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U70 (
    .O(n895),
    .I0(in_41),
    .I1(in_29)
  );
  //AND U70bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U70bar (
    .O(n895bar),
    .I0(in_41bar),
    .I1(in_29bar)
  );
  //OR U71
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U71 (
    .O(n896),
    .I0(in_66),
    .I1(n894)
  );
  //AND U71bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U71bar (
    .O(n896bar),
    .I0(in_66bar),
    .I1(n894bar)
  );
  //OR U72
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U72 (
    .O(n894),
    .I0(in_76),
    .I1(in_71)
  );
  //AND U72bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U72bar (
    .O(n894bar),
    .I0(in_76bar),
    .I1(in_71bar)
  );
  //OR U73
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U73 (
    .O(out[4]),
    .I0(n893),
    .I1(n892)
  );
  //AND U73bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U73bar (
    .O(outbar[4]),
    .I0(n893bar),
    .I1(n892bar)
  );
  //OR U74
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U74 (
    .O(n892),
    .I0(n891),
    .I1(n890)
  );
  //AND U74bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U74bar (
    .O(n892bar),
    .I0(n891bar),
    .I1(n890bar)
  );
  //OR U75
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U75 (
    .O(n890),
    .I0(n889),
    .I1(n888)
  );
  //AND U75bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U75bar (
    .O(n890bar),
    .I0(n889bar),
    .I1(n888bar)
  );
  //OR U76
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U76 (
    .O(n888),
    .I0(n922),
    .I1(n887)
  );
  //AND U76bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U76bar (
    .O(n888bar),
    .I0(n922bar),
    .I1(n887bar)
  );
  //OR U77
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U77 (
    .O(n922),
    .I0(n886),
    .I1(n885)
  );
  //AND U77bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U77bar (
    .O(n922bar),
    .I0(n886bar),
    .I1(n885bar)
  );
  //OR U78
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U78 (
    .O(n885),
    .I0(n884),
    .I1(n883)
  );
  //AND U78bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U78bar (
    .O(n885bar),
    .I0(n884bar),
    .I1(n883bar)
  );
  //OR U79
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U79 (
    .O(n883),
    .I0(n882),
    .I1(n881)
  );
  //AND U79bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U79bar (
    .O(n883bar),
    .I0(n882bar),
    .I1(n881bar)
  );
  //OR U80
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U80 (
    .O(n881),
    .I0(in[118]),
    .I1(in[109])
  );
  //AND U80bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U80bar (
    .O(n881bar),
    .I0(inbar[118]),
    .I1(inbar[109])
  );
  //OR U81
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U81 (
    .O(n882),
    .I0(in[139]),
    .I1(in[120])
  );
  //AND U81bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U81bar (
    .O(n882bar),
    .I0(inbar[139]),
    .I1(inbar[120])
  );
  //OR U82
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U82 (
    .O(n884),
    .I0(n880),
    .I1(n879)
  );
  //AND U82bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U82bar (
    .O(n884bar),
    .I0(n880bar),
    .I1(n879bar)
  );
  //OR U83
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U83 (
    .O(n879),
    .I0(in[198]),
    .I1(in[154])
  );
  //AND U83bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U83bar (
    .O(n879bar),
    .I0(inbar[198]),
    .I1(inbar[154])
  );
  //OR U84
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U84 (
    .O(n880),
    .I0(in[210]),
    .I1(in[205])
  );
  //AND U84bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U84bar (
    .O(n880bar),
    .I0(inbar[210]),
    .I1(inbar[205])
  );
  //OR U85
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U85 (
    .O(n886),
    .I0(n878),
    .I1(n877)
  );
  //AND U85bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U85bar (
    .O(n886bar),
    .I0(n878bar),
    .I1(n877bar)
  );
  //OR U86
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U86 (
    .O(n877),
    .I0(n876),
    .I1(n875)
  );
  //AND U86bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U86bar (
    .O(n877bar),
    .I0(n876bar),
    .I1(n875bar)
  );
  //OR U87
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U87 (
    .O(n875),
    .I0(in[219]),
    .I1(in[217])
  );
  //AND U87bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U87bar (
    .O(n875bar),
    .I0(inbar[219]),
    .I1(inbar[217])
  );
  //OR U88
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U88 (
    .O(n876),
    .I0(in[86]),
    .I1(in[252])
  );
  //AND U88bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U88bar (
    .O(n876bar),
    .I0(inbar[86]),
    .I1(inbar[252])
  );
  //OR U89
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U89 (
    .O(n878),
    .I0(n874),
    .I1(n873)
  );
  //AND U89bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U89bar (
    .O(n878bar),
    .I0(n874bar),
    .I1(n873bar)
  );
  //OR U90
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U90 (
    .O(n873),
    .I0(in_40),
    .I1(in[91])
  );
  //AND U90bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U90bar (
    .O(n873bar),
    .I0(in_40bar),
    .I1(inbar[91])
  );
  //OR U91
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U91 (
    .O(n874),
    .I0(in_8),
    .I1(in_46)
  );
  //AND U91bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U91bar (
    .O(n874bar),
    .I0(in_8bar),
    .I1(in_46bar)
  );
  //OR U92
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U92 (
    .O(n889),
    .I0(n872),
    .I1(n871)
  );
  //AND U92bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U92bar (
    .O(n889bar),
    .I0(n872bar),
    .I1(n871bar)
  );
  //OR U93
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U93 (
    .O(n871),
    .I0(in[117]),
    .I1(n943)
  );
  //AND U93bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U93bar (
    .O(n871bar),
    .I0(inbar[117]),
    .I1(n943bar)
  );
  //OR U94
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U94 (
    .O(n943),
    .I0(n870),
    .I1(n869)
  );
  //AND U94bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U94bar (
    .O(n943bar),
    .I0(n870bar),
    .I1(n869bar)
  );
  //OR U95
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U95 (
    .O(n869),
    .I0(n868),
    .I1(n867)
  );
  //AND U95bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U95bar (
    .O(n869bar),
    .I0(n868bar),
    .I1(n867bar)
  );
  //OR U96
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U96 (
    .O(n867),
    .I0(n866),
    .I1(n865)
  );
  //AND U96bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U96bar (
    .O(n867bar),
    .I0(n866bar),
    .I1(n865bar)
  );
  //OR U97
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U97 (
    .O(n865),
    .I0(n864),
    .I1(n863)
  );
  //AND U97bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U97bar (
    .O(n865bar),
    .I0(n864bar),
    .I1(n863bar)
  );
  //OR U98
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U98 (
    .O(n866),
    .I0(in[108]),
    .I1(n919)
  );
  //AND U98bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U98bar (
    .O(n866bar),
    .I0(inbar[108]),
    .I1(n919bar)
  );
  //OR U99
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U99 (
    .O(n919),
    .I0(n862),
    .I1(n861)
  );
  //AND U99bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U99bar (
    .O(n919bar),
    .I0(n862bar),
    .I1(n861bar)
  );
  //OR U100
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U100 (
    .O(n861),
    .I0(n860),
    .I1(n859)
  );
  //AND U100bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U100bar (
    .O(n861bar),
    .I0(n860bar),
    .I1(n859bar)
  );
  //OR U101
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U101 (
    .O(n859),
    .I0(n858),
    .I1(n857)
  );
  //AND U101bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U101bar (
    .O(n859bar),
    .I0(n858bar),
    .I1(n857bar)
  );
  //OR U102
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U102 (
    .O(n857),
    .I0(in[119]),
    .I1(in[105])
  );
  //AND U102bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U102bar (
    .O(n857bar),
    .I0(inbar[119]),
    .I1(inbar[105])
  );
  //OR U103
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U103 (
    .O(n858),
    .I0(in[186]),
    .I1(in[175])
  );
  //AND U103bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U103bar (
    .O(n858bar),
    .I0(inbar[186]),
    .I1(inbar[175])
  );
  //OR U104
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U104 (
    .O(n860),
    .I0(n856),
    .I1(n855)
  );
  //AND U104bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U104bar (
    .O(n860bar),
    .I0(n856bar),
    .I1(n855bar)
  );
  //OR U105
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U105 (
    .O(n855),
    .I0(in[202]),
    .I1(in[193])
  );
  //AND U105bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U105bar (
    .O(n855bar),
    .I0(inbar[202]),
    .I1(inbar[193])
  );
  //OR U106
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U106 (
    .O(n856),
    .I0(in[225]),
    .I1(in[208])
  );
  //AND U106bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U106bar (
    .O(n856bar),
    .I0(inbar[225]),
    .I1(inbar[208])
  );
  //OR U107
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U107 (
    .O(n862),
    .I0(n854),
    .I1(n853)
  );
  //AND U107bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U107bar (
    .O(n862bar),
    .I0(n854bar),
    .I1(n853bar)
  );
  //OR U108
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U108 (
    .O(n853),
    .I0(n852),
    .I1(n851)
  );
  //AND U108bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U108bar (
    .O(n853bar),
    .I0(n852bar),
    .I1(n851bar)
  );
  //OR U109
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U109 (
    .O(n851),
    .I0(in_1),
    .I1(in[85])
  );
  //AND U109bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U109bar (
    .O(n851bar),
    .I0(in_1bar),
    .I1(inbar[85])
  );
  //OR U110
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U110 (
    .O(n852),
    .I0(in_23),
    .I1(in_19)
  );
  //AND U110bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U110bar (
    .O(n852bar),
    .I0(in_23bar),
    .I1(in_19bar)
  );
  //OR U111
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U111 (
    .O(n854),
    .I0(n850),
    .I1(n849)
  );
  //AND U111bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U111bar (
    .O(n854bar),
    .I0(n850bar),
    .I1(n849bar)
  );
  //OR U112
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U112 (
    .O(n849),
    .I0(in_43),
    .I1(in_33)
  );
  //AND U112bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U112bar (
    .O(n849bar),
    .I0(in_43bar),
    .I1(in_33bar)
  );
  //OR U113
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U113 (
    .O(n850),
    .I0(in_63),
    .I1(in_44)
  );
  //AND U113bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U113bar (
    .O(n850bar),
    .I0(in_63bar),
    .I1(in_44bar)
  );
  //OR U114
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U114 (
    .O(n868),
    .I0(n848),
    .I1(n847)
  );
  //AND U114bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U114bar (
    .O(n868bar),
    .I0(n848bar),
    .I1(n847bar)
  );
  //OR U115
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U115 (
    .O(n847),
    .I0(in[141]),
    .I1(in[112])
  );
  //AND U115bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U115bar (
    .O(n847bar),
    .I0(inbar[141]),
    .I1(inbar[112])
  );
  //OR U116
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U116 (
    .O(n848),
    .I0(in[147]),
    .I1(n846)
  );
  //AND U116bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U116bar (
    .O(n848bar),
    .I0(inbar[147]),
    .I1(n846bar)
  );
  //OR U117
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U117 (
    .O(n846),
    .I0(in[181]),
    .I1(in[167])
  );
  //AND U117bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U117bar (
    .O(n846bar),
    .I0(inbar[181]),
    .I1(inbar[167])
  );
  //OR U118
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U118 (
    .O(n870),
    .I0(n845),
    .I1(n844)
  );
  //AND U118bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U118bar (
    .O(n870bar),
    .I0(n845bar),
    .I1(n844bar)
  );
  //OR U119
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U119 (
    .O(n844),
    .I0(n843),
    .I1(n842)
  );
  //AND U119bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U119bar (
    .O(n844bar),
    .I0(n843bar),
    .I1(n842bar)
  );
  //OR U120
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U120 (
    .O(n842),
    .I0(in[229]),
    .I1(in[201])
  );
  //AND U120bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U120bar (
    .O(n842bar),
    .I0(inbar[229]),
    .I1(inbar[201])
  );
  //OR U121
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U121 (
    .O(n843),
    .I0(in[237]),
    .I1(n841)
  );
  //AND U121bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U121bar (
    .O(n843bar),
    .I0(inbar[237]),
    .I1(n841bar)
  );
  //OR U122
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U122 (
    .O(n841),
    .I0(in[94]),
    .I1(in[253])
  );
  //AND U122bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U122bar (
    .O(n841bar),
    .I0(inbar[94]),
    .I1(inbar[253])
  );
  //OR U123
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U123 (
    .O(n845),
    .I0(n840),
    .I1(n839)
  );
  //AND U123bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U123bar (
    .O(n845bar),
    .I0(n840bar),
    .I1(n839bar)
  );
  //OR U124
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U124 (
    .O(n839),
    .I0(in_21),
    .I1(in[96])
  );
  //AND U124bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U124bar (
    .O(n839bar),
    .I0(in_21bar),
    .I1(inbar[96])
  );
  //OR U125
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U125 (
    .O(n840),
    .I0(in_25),
    .I1(n838)
  );
  //AND U125bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U125bar (
    .O(n840bar),
    .I0(in_25bar),
    .I1(n838bar)
  );
  //OR U126
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U126 (
    .O(n838),
    .I0(in_81),
    .I1(in_45)
  );
  //AND U126bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U126bar (
    .O(n838bar),
    .I0(in_81bar),
    .I1(in_45bar)
  );
  //OR U127
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U127 (
    .O(n891),
    .I0(n837),
    .I1(n836)
  );
  //AND U127bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U127bar (
    .O(n891bar),
    .I0(n837bar),
    .I1(n836bar)
  );
  //OR U128
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U128 (
    .O(n836),
    .I0(in[142]),
    .I1(in[124])
  );
  //AND U128bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U128bar (
    .O(n836bar),
    .I0(inbar[142]),
    .I1(inbar[124])
  );
  //OR U129
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U129 (
    .O(n837),
    .I0(in[150]),
    .I1(n835)
  );
  //AND U129bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U129bar (
    .O(n837bar),
    .I0(inbar[150]),
    .I1(n835bar)
  );
  //OR U130
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U130 (
    .O(n835),
    .I0(in[172]),
    .I1(in[155])
  );
  //AND U130bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U130bar (
    .O(n835bar),
    .I0(inbar[172]),
    .I1(inbar[155])
  );
  //OR U131
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U131 (
    .O(n893),
    .I0(n834),
    .I1(n833)
  );
  //AND U131bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U131bar (
    .O(n893bar),
    .I0(n834bar),
    .I1(n833bar)
  );
  //OR U132
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U132 (
    .O(n833),
    .I0(n832),
    .I1(n831)
  );
  //AND U132bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U132bar (
    .O(n833bar),
    .I0(n832bar),
    .I1(n831bar)
  );
  //OR U133
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U133 (
    .O(n831),
    .I0(in[196]),
    .I1(in[173])
  );
  //AND U133bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U133bar (
    .O(n831bar),
    .I0(inbar[196]),
    .I1(inbar[173])
  );
  //OR U134
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U134 (
    .O(n832),
    .I0(in[222]),
    .I1(n830)
  );
  //AND U134bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U134bar (
    .O(n832bar),
    .I0(inbar[222]),
    .I1(n830bar)
  );
  //OR U135
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U135 (
    .O(n830),
    .I0(in[227]),
    .I1(in[226])
  );
  //AND U135bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U135bar (
    .O(n830bar),
    .I0(inbar[227]),
    .I1(inbar[226])
  );
  //OR U136
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U136 (
    .O(n834),
    .I0(n829),
    .I1(n828)
  );
  //AND U136bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U136bar (
    .O(n834bar),
    .I0(n829bar),
    .I1(n828bar)
  );
  //OR U137
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U137 (
    .O(n828),
    .I0(in[249]),
    .I1(in[231])
  );
  //AND U137bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U137bar (
    .O(n828bar),
    .I0(inbar[249]),
    .I1(inbar[231])
  );
  //OR U138
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U138 (
    .O(n829),
    .I0(in_28),
    .I1(n827)
  );
  //AND U138bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U138bar (
    .O(n829bar),
    .I0(in_28bar),
    .I1(n827bar)
  );
  //OR U139
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U139 (
    .O(n827),
    .I0(in_52),
    .I1(in_47)
  );
  //AND U139bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U139bar (
    .O(n827bar),
    .I0(in_52bar),
    .I1(in_47bar)
  );
  //OR U140
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U140 (
    .O(out[3]),
    .I0(n826),
    .I1(n825)
  );
  //AND U140bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U140bar (
    .O(outbar[3]),
    .I0(n826bar),
    .I1(n825bar)
  );
  //OR U141
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U141 (
    .O(n825),
    .I0(n824),
    .I1(n823)
  );
  //AND U141bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U141bar (
    .O(n825bar),
    .I0(n824bar),
    .I1(n823bar)
  );
  //OR U142
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U142 (
    .O(n823),
    .I0(n822),
    .I1(n821)
  );
  //AND U142bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U142bar (
    .O(n823bar),
    .I0(n822bar),
    .I1(n821bar)
  );
  //OR U143
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U143 (
    .O(n821),
    .I0(n820),
    .I1(n819)
  );
  //AND U143bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U143bar (
    .O(n821bar),
    .I0(n820bar),
    .I1(n819bar)
  );
  //OR U144
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U144 (
    .O(n822),
    .I0(n964),
    .I1(n818)
  );
  //AND U144bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U144bar (
    .O(n822bar),
    .I0(n964bar),
    .I1(n818bar)
  );
  //OR U145
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U145 (
    .O(n818),
    .I0(in[118]),
    .I1(n817)
  );
  //AND U145bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U145bar (
    .O(n818bar),
    .I0(inbar[118]),
    .I1(n817bar)
  );
  //OR U146
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U146 (
    .O(n964),
    .I0(n816),
    .I1(n815)
  );
  //AND U146bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U146bar (
    .O(n964bar),
    .I0(n816bar),
    .I1(n815bar)
  );
  //OR U147
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U147 (
    .O(n815),
    .I0(n814),
    .I1(n813)
  );
  //AND U147bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U147bar (
    .O(n815bar),
    .I0(n814bar),
    .I1(n813bar)
  );
  //OR U148
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U148 (
    .O(n813),
    .I0(n812),
    .I1(n811)
  );
  //AND U148bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U148bar (
    .O(n813bar),
    .I0(n812bar),
    .I1(n811bar)
  );
  //OR U149
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U149 (
    .O(n811),
    .I0(in[122]),
    .I1(in[111])
  );
  //AND U149bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U149bar (
    .O(n811bar),
    .I0(inbar[122]),
    .I1(inbar[111])
  );
  //OR U150
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U150 (
    .O(n812),
    .I0(in[154]),
    .I1(in[151])
  );
  //AND U150bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U150bar (
    .O(n812bar),
    .I0(inbar[154]),
    .I1(inbar[151])
  );
  //OR U151
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U151 (
    .O(n814),
    .I0(n810),
    .I1(n809)
  );
  //AND U151bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U151bar (
    .O(n814bar),
    .I0(n810bar),
    .I1(n809bar)
  );
  //OR U152
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U152 (
    .O(n809),
    .I0(in[187]),
    .I1(in[177])
  );
  //AND U152bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U152bar (
    .O(n809bar),
    .I0(inbar[187]),
    .I1(inbar[177])
  );
  //OR U153
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U153 (
    .O(n810),
    .I0(in[200]),
    .I1(in[192])
  );
  //AND U153bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U153bar (
    .O(n810bar),
    .I0(inbar[200]),
    .I1(inbar[192])
  );
  //OR U154
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U154 (
    .O(n816),
    .I0(n808),
    .I1(n807)
  );
  //AND U154bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U154bar (
    .O(n816bar),
    .I0(n808bar),
    .I1(n807bar)
  );
  //OR U155
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U155 (
    .O(n807),
    .I0(n806),
    .I1(n805)
  );
  //AND U155bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U155bar (
    .O(n807bar),
    .I0(n806bar),
    .I1(n805bar)
  );
  //OR U156
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U156 (
    .O(n805),
    .I0(in[225]),
    .I1(in[207])
  );
  //AND U156bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U156bar (
    .O(n805bar),
    .I0(inbar[225]),
    .I1(inbar[207])
  );
  //OR U157
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U157 (
    .O(n806),
    .I0(in[98]),
    .I1(in[226])
  );
  //AND U157bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U157bar (
    .O(n806bar),
    .I0(inbar[98]),
    .I1(inbar[226])
  );
  //OR U158
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U158 (
    .O(n808),
    .I0(n804),
    .I1(n803)
  );
  //AND U158bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U158bar (
    .O(n808bar),
    .I0(n804bar),
    .I1(n803bar)
  );
  //OR U159
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U159 (
    .O(n803),
    .I0(in_20),
    .I1(in_16)
  );
  //AND U159bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U159bar (
    .O(n803bar),
    .I0(in_20bar),
    .I1(in_16bar)
  );
  //OR U160
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U160 (
    .O(n804),
    .I0(in_55),
    .I1(in_45)
  );
  //AND U160bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U160bar (
    .O(n804bar),
    .I0(in_55bar),
    .I1(in_45bar)
  );
  //OR U161
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U161 (
    .O(n824),
    .I0(n802),
    .I1(n801)
  );
  //AND U161bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U161bar (
    .O(n824bar),
    .I0(n802bar),
    .I1(n801bar)
  );
  //OR U162
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U162 (
    .O(n801),
    .I0(in[162]),
    .I1(in[149])
  );
  //AND U162bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U162bar (
    .O(n801bar),
    .I0(inbar[162]),
    .I1(inbar[149])
  );
  //OR U163
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U163 (
    .O(n802),
    .I0(in[163]),
    .I1(n800)
  );
  //AND U163bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U163bar (
    .O(n802bar),
    .I0(inbar[163]),
    .I1(n800bar)
  );
  //OR U164
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U164 (
    .O(n800),
    .I0(in[191]),
    .I1(in[189])
  );
  //AND U164bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U164bar (
    .O(n800bar),
    .I0(inbar[191]),
    .I1(inbar[189])
  );
  //OR U165
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U165 (
    .O(n826),
    .I0(n799),
    .I1(n798)
  );
  //AND U165bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U165bar (
    .O(n826bar),
    .I0(n799bar),
    .I1(n798bar)
  );
  //OR U166
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U166 (
    .O(n798),
    .I0(n797),
    .I1(n796)
  );
  //AND U166bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U166bar (
    .O(n798bar),
    .I0(n797bar),
    .I1(n796bar)
  );
  //OR U167
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U167 (
    .O(n796),
    .I0(in[212]),
    .I1(in[193])
  );
  //AND U167bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U167bar (
    .O(n796bar),
    .I0(inbar[212]),
    .I1(inbar[193])
  );
  //OR U168
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U168 (
    .O(n797),
    .I0(in[238]),
    .I1(n795)
  );
  //AND U168bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U168bar (
    .O(n797bar),
    .I0(inbar[238]),
    .I1(n795bar)
  );
  //OR U169
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U169 (
    .O(n795),
    .I0(in[88]),
    .I1(in[247])
  );
  //AND U169bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U169bar (
    .O(n795bar),
    .I0(inbar[88]),
    .I1(inbar[247])
  );
  //OR U170
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U170 (
    .O(n799),
    .I0(n794),
    .I1(n793)
  );
  //AND U170bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U170bar (
    .O(n799bar),
    .I0(n794bar),
    .I1(n793bar)
  );
  //OR U171
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U171 (
    .O(n793),
    .I0(in[94]),
    .I1(in[92])
  );
  //AND U171bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U171bar (
    .O(n793bar),
    .I0(inbar[94]),
    .I1(inbar[92])
  );
  //OR U172
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U172 (
    .O(n794),
    .I0(in_52),
    .I1(n792)
  );
  //AND U172bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U172bar (
    .O(n794bar),
    .I0(in_52bar),
    .I1(n792bar)
  );
  //OR U173
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U173 (
    .O(n792),
    .I0(in_70),
    .I1(in_67)
  );
  //AND U173bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U173bar (
    .O(n792bar),
    .I0(in_70bar),
    .I1(in_67bar)
  );
  //OR U174
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U174 (
    .O(out[2]),
    .I0(n791),
    .I1(n790)
  );
  //AND U174bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U174bar (
    .O(outbar[2]),
    .I0(n791bar),
    .I1(n790bar)
  );
  //OR U175
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U175 (
    .O(n790),
    .I0(n789),
    .I1(n788)
  );
  //AND U175bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U175bar (
    .O(n790bar),
    .I0(n789bar),
    .I1(n788bar)
  );
  //OR U176
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U176 (
    .O(n788),
    .I0(n787),
    .I1(n786)
  );
  //AND U176bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U176bar (
    .O(n788bar),
    .I0(n787bar),
    .I1(n786bar)
  );
  //OR U177
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U177 (
    .O(n786),
    .I0(n819),
    .I1(n785)
  );
  //AND U177bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U177bar (
    .O(n786bar),
    .I0(n819bar),
    .I1(n785bar)
  );
  //OR U178
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U178 (
    .O(n819),
    .I0(n784),
    .I1(n783)
  );
  //AND U178bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U178bar (
    .O(n819bar),
    .I0(n784bar),
    .I1(n783bar)
  );
  //OR U179
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U179 (
    .O(n783),
    .I0(n782),
    .I1(n781)
  );
  //AND U179bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U179bar (
    .O(n783bar),
    .I0(n782bar),
    .I1(n781bar)
  );
  //OR U180
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U180 (
    .O(n781),
    .I0(n780),
    .I1(n779)
  );
  //AND U180bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U180bar (
    .O(n781bar),
    .I0(n780bar),
    .I1(n779bar)
  );
  //OR U181
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U181 (
    .O(n779),
    .I0(n962),
    .I1(n778)
  );
  //AND U181bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U181bar (
    .O(n779bar),
    .I0(n962bar),
    .I1(n778bar)
  );
  //OR U182
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U182 (
    .O(n962),
    .I0(n777),
    .I1(n776)
  );
  //AND U182bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U182bar (
    .O(n962bar),
    .I0(n777bar),
    .I1(n776bar)
  );
  //OR U183
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U183 (
    .O(n776),
    .I0(n775),
    .I1(n774)
  );
  //AND U183bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U183bar (
    .O(n776bar),
    .I0(n775bar),
    .I1(n774bar)
  );
  //OR U184
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U184 (
    .O(n774),
    .I0(n773),
    .I1(n772)
  );
  //AND U184bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U184bar (
    .O(n774bar),
    .I0(n773bar),
    .I1(n772bar)
  );
  //OR U185
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U185 (
    .O(n772),
    .I0(in[131]),
    .I1(in[120])
  );
  //AND U185bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U185bar (
    .O(n772bar),
    .I0(inbar[131]),
    .I1(inbar[120])
  );
  //OR U186
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U186 (
    .O(n773),
    .I0(in[153]),
    .I1(in[147])
  );
  //AND U186bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U186bar (
    .O(n773bar),
    .I0(inbar[153]),
    .I1(inbar[147])
  );
  //OR U187
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U187 (
    .O(n775),
    .I0(n771),
    .I1(n770)
  );
  //AND U187bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U187bar (
    .O(n775bar),
    .I0(n771bar),
    .I1(n770bar)
  );
  //OR U188
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U188 (
    .O(n770),
    .I0(in[170]),
    .I1(in[156])
  );
  //AND U188bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U188bar (
    .O(n770bar),
    .I0(inbar[170]),
    .I1(inbar[156])
  );
  //OR U189
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U189 (
    .O(n771),
    .I0(in[223]),
    .I1(in[190])
  );
  //AND U189bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U189bar (
    .O(n771bar),
    .I0(inbar[223]),
    .I1(inbar[190])
  );
  //OR U190
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U190 (
    .O(n777),
    .I0(n769),
    .I1(n768)
  );
  //AND U190bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U190bar (
    .O(n777bar),
    .I0(n769bar),
    .I1(n768bar)
  );
  //OR U191
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U191 (
    .O(n768),
    .I0(n767),
    .I1(n766)
  );
  //AND U191bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U191bar (
    .O(n768bar),
    .I0(n767bar),
    .I1(n766bar)
  );
  //OR U192
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U192 (
    .O(n766),
    .I0(in[236]),
    .I1(in[230])
  );
  //AND U192bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U192bar (
    .O(n766bar),
    .I0(inbar[236]),
    .I1(inbar[230])
  );
  //OR U193
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U193 (
    .O(n767),
    .I0(in[85]),
    .I1(in[240])
  );
  //AND U193bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U193bar (
    .O(n767bar),
    .I0(inbar[85]),
    .I1(inbar[240])
  );
  //OR U194
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U194 (
    .O(n769),
    .I0(n765),
    .I1(n764)
  );
  //AND U194bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U194bar (
    .O(n769bar),
    .I0(n765bar),
    .I1(n764bar)
  );
  //OR U195
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U195 (
    .O(n764),
    .I0(in_12),
    .I1(in[90])
  );
  //AND U195bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U195bar (
    .O(n764bar),
    .I0(in_12bar),
    .I1(inbar[90])
  );
  //OR U196
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U196 (
    .O(n765),
    .I0(in_39),
    .I1(in_28)
  );
  //AND U196bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U196bar (
    .O(n765bar),
    .I0(in_39bar),
    .I1(in_28bar)
  );
  //OR U197
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U197 (
    .O(n780),
    .I0(in[109]),
    .I1(n763)
  );
  //AND U197bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U197bar (
    .O(n780bar),
    .I0(inbar[109]),
    .I1(n763bar)
  );
  //OR U198
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U198 (
    .O(n782),
    .I0(n762),
    .I1(n761)
  );
  //AND U198bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U198bar (
    .O(n782bar),
    .I0(n762bar),
    .I1(n761bar)
  );
  //OR U199
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U199 (
    .O(n761),
    .I0(in[138]),
    .I1(in[129])
  );
  //AND U199bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U199bar (
    .O(n761bar),
    .I0(inbar[138]),
    .I1(inbar[129])
  );
  //OR U200
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U200 (
    .O(n762),
    .I0(in[157]),
    .I1(n760)
  );
  //AND U200bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U200bar (
    .O(n762bar),
    .I0(inbar[157]),
    .I1(n760bar)
  );
  //OR U201
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U201 (
    .O(n760),
    .I0(in[182]),
    .I1(in[167])
  );
  //AND U201bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U201bar (
    .O(n760bar),
    .I0(inbar[182]),
    .I1(inbar[167])
  );
  //OR U202
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U202 (
    .O(n784),
    .I0(n759),
    .I1(n758)
  );
  //AND U202bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U202bar (
    .O(n784bar),
    .I0(n759bar),
    .I1(n758bar)
  );
  //OR U203
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U203 (
    .O(n758),
    .I0(n757),
    .I1(n756)
  );
  //AND U203bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U203bar (
    .O(n758bar),
    .I0(n757bar),
    .I1(n756bar)
  );
  //OR U204
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U204 (
    .O(n756),
    .I0(in[195]),
    .I1(in[184])
  );
  //AND U204bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U204bar (
    .O(n756bar),
    .I0(inbar[195]),
    .I1(inbar[184])
  );
  //OR U205
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U205 (
    .O(n757),
    .I0(in[196]),
    .I1(n755)
  );
  //AND U205bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U205bar (
    .O(n757bar),
    .I0(inbar[196]),
    .I1(n755bar)
  );
  //OR U206
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U206 (
    .O(n755),
    .I0(in[215]),
    .I1(in[209])
  );
  //AND U206bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U206bar (
    .O(n755bar),
    .I0(inbar[215]),
    .I1(inbar[209])
  );
  //OR U207
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U207 (
    .O(n759),
    .I0(n754),
    .I1(n753)
  );
  //AND U207bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U207bar (
    .O(n759bar),
    .I0(n754bar),
    .I1(n753bar)
  );
  //OR U208
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U208 (
    .O(n753),
    .I0(in[93]),
    .I1(in[233])
  );
  //AND U208bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U208bar (
    .O(n753bar),
    .I0(inbar[93]),
    .I1(inbar[233])
  );
  //OR U209
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U209 (
    .O(n754),
    .I0(in_1),
    .I1(n752)
  );
  //AND U209bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U209bar (
    .O(n754bar),
    .I0(in_1bar),
    .I1(n752bar)
  );
  //OR U210
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U210 (
    .O(n752),
    .I0(in_69),
    .I1(in_66)
  );
  //AND U210bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U210bar (
    .O(n752bar),
    .I0(in_69bar),
    .I1(in_66bar)
  );
  //OR U211
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U211 (
    .O(n787),
    .I0(n966),
    .I1(n751)
  );
  //AND U211bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U211bar (
    .O(n787bar),
    .I0(n966bar),
    .I1(n751bar)
  );
  //OR U212
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U212 (
    .O(n751),
    .I0(in[134]),
    .I1(n750)
  );
  //AND U212bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U212bar (
    .O(n751bar),
    .I0(inbar[134]),
    .I1(n750bar)
  );
  //OR U213
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U213 (
    .O(n966),
    .I0(n749),
    .I1(n748)
  );
  //AND U213bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U213bar (
    .O(n966bar),
    .I0(n749bar),
    .I1(n748bar)
  );
  //OR U214
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U214 (
    .O(n748),
    .I0(n747),
    .I1(n746)
  );
  //AND U214bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U214bar (
    .O(n748bar),
    .I0(n747bar),
    .I1(n746bar)
  );
  //OR U215
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U215 (
    .O(n746),
    .I0(n745),
    .I1(n744)
  );
  //AND U215bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U215bar (
    .O(n746bar),
    .I0(n745bar),
    .I1(n744bar)
  );
  //OR U216
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U216 (
    .O(n744),
    .I0(in[136]),
    .I1(in[121])
  );
  //AND U216bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U216bar (
    .O(n744bar),
    .I0(inbar[136]),
    .I1(inbar[121])
  );
  //OR U217
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U217 (
    .O(n745),
    .I0(in[186]),
    .I1(in[174])
  );
  //AND U217bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U217bar (
    .O(n745bar),
    .I0(inbar[186]),
    .I1(inbar[174])
  );
  //OR U218
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U218 (
    .O(n747),
    .I0(n743),
    .I1(n742)
  );
  //AND U218bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U218bar (
    .O(n747bar),
    .I0(n743bar),
    .I1(n742bar)
  );
  //OR U219
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U219 (
    .O(n742),
    .I0(in[198]),
    .I1(in[197])
  );
  //AND U219bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U219bar (
    .O(n742bar),
    .I0(inbar[198]),
    .I1(inbar[197])
  );
  //OR U220
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U220 (
    .O(n743),
    .I0(in[214]),
    .I1(in[199])
  );
  //AND U220bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U220bar (
    .O(n743bar),
    .I0(inbar[214]),
    .I1(inbar[199])
  );
  //OR U221
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U221 (
    .O(n749),
    .I0(n741),
    .I1(n740)
  );
  //AND U221bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U221bar (
    .O(n749bar),
    .I0(n741bar),
    .I1(n740bar)
  );
  //OR U222
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U222 (
    .O(n740),
    .I0(n739),
    .I1(n738)
  );
  //AND U222bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U222bar (
    .O(n740bar),
    .I0(n739bar),
    .I1(n738bar)
  );
  //OR U223
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U223 (
    .O(n738),
    .I0(in[231]),
    .I1(in[220])
  );
  //AND U223bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U223bar (
    .O(n738bar),
    .I0(inbar[231]),
    .I1(inbar[220])
  );
  //OR U224
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U224 (
    .O(n739),
    .I0(in_25),
    .I1(in[245])
  );
  //AND U224bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U224bar (
    .O(n739bar),
    .I0(in_25bar),
    .I1(inbar[245])
  );
  //OR U225
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U225 (
    .O(n741),
    .I0(n737),
    .I1(n736)
  );
  //AND U225bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U225bar (
    .O(n741bar),
    .I0(n737bar),
    .I1(n736bar)
  );
  //OR U226
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U226 (
    .O(n736),
    .I0(in_53),
    .I1(in_29)
  );
  //AND U226bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U226bar (
    .O(n736bar),
    .I0(in_53bar),
    .I1(in_29bar)
  );
  //OR U227
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U227 (
    .O(n737),
    .I0(in_79),
    .I1(in_74)
  );
  //AND U227bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U227bar (
    .O(n737bar),
    .I0(in_79bar),
    .I1(in_74bar)
  );
  //OR U228
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U228 (
    .O(n789),
    .I0(n735),
    .I1(n734)
  );
  //AND U228bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U228bar (
    .O(n789bar),
    .I0(n735bar),
    .I1(n734bar)
  );
  //OR U229
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U229 (
    .O(n734),
    .I0(in[152]),
    .I1(in[140])
  );
  //AND U229bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U229bar (
    .O(n734bar),
    .I0(inbar[152]),
    .I1(inbar[140])
  );
  //OR U230
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U230 (
    .O(n735),
    .I0(in[155]),
    .I1(n733)
  );
  //AND U230bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U230bar (
    .O(n735bar),
    .I0(inbar[155]),
    .I1(n733bar)
  );
  //OR U231
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U231 (
    .O(n733),
    .I0(in[166]),
    .I1(in[165])
  );
  //AND U231bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U231bar (
    .O(n733bar),
    .I0(inbar[166]),
    .I1(inbar[165])
  );
  //OR U232
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U232 (
    .O(n791),
    .I0(n732),
    .I1(n731)
  );
  //AND U232bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U232bar (
    .O(n791bar),
    .I0(n732bar),
    .I1(n731bar)
  );
  //OR U233
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U233 (
    .O(n731),
    .I0(n730),
    .I1(n729)
  );
  //AND U233bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U233bar (
    .O(n731bar),
    .I0(n730bar),
    .I1(n729bar)
  );
  //OR U234
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U234 (
    .O(n729),
    .I0(in[202]),
    .I1(in[185])
  );
  //AND U234bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U234bar (
    .O(n729bar),
    .I0(inbar[202]),
    .I1(inbar[185])
  );
  //OR U235
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U235 (
    .O(n730),
    .I0(in[211]),
    .I1(n728)
  );
  //AND U235bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U235bar (
    .O(n730bar),
    .I0(inbar[211]),
    .I1(n728bar)
  );
  //OR U236
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U236 (
    .O(n728),
    .I0(in[255]),
    .I1(in[253])
  );
  //AND U236bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U236bar (
    .O(n728bar),
    .I0(inbar[255]),
    .I1(inbar[253])
  );
  //OR U237
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U237 (
    .O(n732),
    .I0(n727),
    .I1(n726)
  );
  //AND U237bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U237bar (
    .O(n732bar),
    .I0(n727bar),
    .I1(n726bar)
  );
  //OR U238
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U238 (
    .O(n726),
    .I0(in_35),
    .I1(in_15)
  );
  //AND U238bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U238bar (
    .O(n726bar),
    .I0(in_35bar),
    .I1(in_15bar)
  );
  //OR U239
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U239 (
    .O(n727),
    .I0(in_36),
    .I1(n725)
  );
  //AND U239bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U239bar (
    .O(n727bar),
    .I0(in_36bar),
    .I1(n725bar)
  );
  //OR U240
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U240 (
    .O(n725),
    .I0(in_48),
    .I1(in_40)
  );
  //AND U240bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U240bar (
    .O(n725bar),
    .I0(in_48bar),
    .I1(in_40bar)
  );
  //OR U241
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U241 (
    .O(out[1]),
    .I0(n724),
    .I1(n723)
  );
  //AND U241bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U241bar (
    .O(outbar[1]),
    .I0(n724bar),
    .I1(n723bar)
  );
  //OR U242
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U242 (
    .O(n723),
    .I0(n722),
    .I1(n721)
  );
  //AND U242bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U242bar (
    .O(n723bar),
    .I0(n722bar),
    .I1(n721bar)
  );
  //OR U243
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U243 (
    .O(n721),
    .I0(n720),
    .I1(n719)
  );
  //AND U243bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U243bar (
    .O(n721bar),
    .I0(n720bar),
    .I1(n719bar)
  );
  //OR U244
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U244 (
    .O(n719),
    .I0(n921),
    .I1(n887)
  );
  //AND U244bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U244bar (
    .O(n719bar),
    .I0(n921bar),
    .I1(n887bar)
  );
  //OR U245
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U245 (
    .O(n887),
    .I0(n718),
    .I1(n717)
  );
  //AND U245bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U245bar (
    .O(n887bar),
    .I0(n718bar),
    .I1(n717bar)
  );
  //OR U246
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U246 (
    .O(n717),
    .I0(n716),
    .I1(n715)
  );
  //AND U246bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U246bar (
    .O(n717bar),
    .I0(n716bar),
    .I1(n715bar)
  );
  //OR U247
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U247 (
    .O(n715),
    .I0(n714),
    .I1(n713)
  );
  //AND U247bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U247bar (
    .O(n715bar),
    .I0(n714bar),
    .I1(n713bar)
  );
  //OR U248
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U248 (
    .O(n713),
    .I0(in[116]),
    .I1(in[110])
  );
  //AND U248bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U248bar (
    .O(n713bar),
    .I0(inbar[116]),
    .I1(inbar[110])
  );
  //OR U249
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U249 (
    .O(n714),
    .I0(in[133]),
    .I1(in[130])
  );
  //AND U249bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U249bar (
    .O(n714bar),
    .I0(inbar[133]),
    .I1(inbar[130])
  );
  //OR U250
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U250 (
    .O(n716),
    .I0(n712),
    .I1(n711)
  );
  //AND U250bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U250bar (
    .O(n716bar),
    .I0(n712bar),
    .I1(n711bar)
  );
  //OR U251
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U251 (
    .O(n711),
    .I0(in[203]),
    .I1(in[135])
  );
  //AND U251bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U251bar (
    .O(n711bar),
    .I0(inbar[203]),
    .I1(inbar[135])
  );
  //OR U252
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U252 (
    .O(n712),
    .I0(in[232]),
    .I1(in[223])
  );
  //AND U252bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U252bar (
    .O(n712bar),
    .I0(inbar[232]),
    .I1(inbar[223])
  );
  //OR U253
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U253 (
    .O(n718),
    .I0(n710),
    .I1(n709)
  );
  //AND U253bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U253bar (
    .O(n718bar),
    .I0(n710bar),
    .I1(n709bar)
  );
  //OR U254
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U254 (
    .O(n709),
    .I0(n708),
    .I1(n707)
  );
  //AND U254bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U254bar (
    .O(n709bar),
    .I0(n708bar),
    .I1(n707bar)
  );
  //OR U255
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U255 (
    .O(n707),
    .I0(in[255]),
    .I1(in[233])
  );
  //AND U255bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U255bar (
    .O(n707bar),
    .I0(inbar[255]),
    .I1(inbar[233])
  );
  //OR U256
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U256 (
    .O(n708),
    .I0(in_53),
    .I1(in_34)
  );
  //AND U256bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U256bar (
    .O(n708bar),
    .I0(in_53bar),
    .I1(in_34bar)
  );
  //OR U257
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U257 (
    .O(n710),
    .I0(n706),
    .I1(n705)
  );
  //AND U257bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U257bar (
    .O(n710bar),
    .I0(n706bar),
    .I1(n705bar)
  );
  //OR U258
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U258 (
    .O(n705),
    .I0(in_57),
    .I1(in_55)
  );
  //AND U258bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U258bar (
    .O(n705bar),
    .I0(in_57bar),
    .I1(in_55bar)
  );
  //OR U259
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U259 (
    .O(n706),
    .I0(in_68),
    .I1(in_67)
  );
  //AND U259bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U259bar (
    .O(n706bar),
    .I0(in_68bar),
    .I1(in_67bar)
  );
  //OR U260
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U260 (
    .O(n921),
    .I0(n704),
    .I1(n703)
  );
  //AND U260bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U260bar (
    .O(n921bar),
    .I0(n704bar),
    .I1(n703bar)
  );
  //OR U261
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U261 (
    .O(n703),
    .I0(n702),
    .I1(n701)
  );
  //AND U261bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U261bar (
    .O(n703bar),
    .I0(n702bar),
    .I1(n701bar)
  );
  //OR U262
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U262 (
    .O(n701),
    .I0(n700),
    .I1(n699)
  );
  //AND U262bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U262bar (
    .O(n701bar),
    .I0(n700bar),
    .I1(n699bar)
  );
  //OR U263
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U263 (
    .O(n699),
    .I0(n944),
    .I1(n872)
  );
  //AND U263bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U263bar (
    .O(n699bar),
    .I0(n944bar),
    .I1(n872bar)
  );
  //OR U264
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U264 (
    .O(n872),
    .I0(n698),
    .I1(n697)
  );
  //AND U264bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U264bar (
    .O(n872bar),
    .I0(n698bar),
    .I1(n697bar)
  );
  //OR U265
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U265 (
    .O(n697),
    .I0(n696),
    .I1(n695)
  );
  //AND U265bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U265bar (
    .O(n697bar),
    .I0(n696bar),
    .I1(n695bar)
  );
  //OR U266
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U266 (
    .O(n695),
    .I0(n694),
    .I1(n693)
  );
  //AND U266bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U266bar (
    .O(n695bar),
    .I0(n694bar),
    .I1(n693bar)
  );
  //OR U267
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U267 (
    .O(n693),
    .I0(in[121]),
    .I1(in[102])
  );
  //AND U267bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U267bar (
    .O(n693bar),
    .I0(inbar[121]),
    .I1(inbar[102])
  );
  //OR U268
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U268 (
    .O(n694),
    .I0(in[162]),
    .I1(in[161])
  );
  //AND U268bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U268bar (
    .O(n694bar),
    .I0(inbar[162]),
    .I1(inbar[161])
  );
  //OR U269
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U269 (
    .O(n696),
    .I0(n692),
    .I1(n691)
  );
  //AND U269bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U269bar (
    .O(n696bar),
    .I0(n692bar),
    .I1(n691bar)
  );
  //OR U270
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U270 (
    .O(n691),
    .I0(in[192]),
    .I1(in[178])
  );
  //AND U270bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U270bar (
    .O(n691bar),
    .I0(inbar[192]),
    .I1(inbar[178])
  );
  //OR U271
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U271 (
    .O(n692),
    .I0(in[244]),
    .I1(in[209])
  );
  //AND U271bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U271bar (
    .O(n692bar),
    .I0(inbar[244]),
    .I1(inbar[209])
  );
  //OR U272
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U272 (
    .O(n698),
    .I0(n690),
    .I1(n689)
  );
  //AND U272bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U272bar (
    .O(n698bar),
    .I0(n690bar),
    .I1(n689bar)
  );
  //OR U273
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U273 (
    .O(n689),
    .I0(n688),
    .I1(n687)
  );
  //AND U273bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U273bar (
    .O(n689bar),
    .I0(n688bar),
    .I1(n687bar)
  );
  //OR U274
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U274 (
    .O(n687),
    .I0(in[90]),
    .I1(in[254])
  );
  //AND U274bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U274bar (
    .O(n687bar),
    .I0(inbar[90]),
    .I1(inbar[254])
  );
  //OR U275
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U275 (
    .O(n688),
    .I0(in_36),
    .I1(in_32)
  );
  //AND U275bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U275bar (
    .O(n688bar),
    .I0(in_36bar),
    .I1(in_32bar)
  );
  //OR U276
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U276 (
    .O(n690),
    .I0(n686),
    .I1(n685)
  );
  //AND U276bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U276bar (
    .O(n690bar),
    .I0(n686bar),
    .I1(n685bar)
  );
  //OR U277
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U277 (
    .O(n685),
    .I0(in_62),
    .I1(in_37)
  );
  //AND U277bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U277bar (
    .O(n685bar),
    .I0(in_62bar),
    .I1(in_37bar)
  );
  //OR U278
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U278 (
    .O(n686),
    .I0(in_75),
    .I1(in_73)
  );
  //AND U278bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U278bar (
    .O(n686bar),
    .I0(in_75bar),
    .I1(in_73bar)
  );
  //OR U279
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U279 (
    .O(n944),
    .I0(n684),
    .I1(n683)
  );
  //AND U279bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U279bar (
    .O(n944bar),
    .I0(n684bar),
    .I1(n683bar)
  );
  //OR U280
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U280 (
    .O(n683),
    .I0(n682),
    .I1(n681)
  );
  //AND U280bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U280bar (
    .O(n683bar),
    .I0(n682bar),
    .I1(n681bar)
  );
  //OR U281
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U281 (
    .O(n681),
    .I0(n680),
    .I1(n679)
  );
  //AND U281bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U281bar (
    .O(n681bar),
    .I0(n680bar),
    .I1(n679bar)
  );
  //OR U282
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U282 (
    .O(n679),
    .I0(in[171]),
    .I1(in[153])
  );
  //AND U282bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U282bar (
    .O(n679bar),
    .I0(inbar[171]),
    .I1(inbar[153])
  );
  //OR U283
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U283 (
    .O(n680),
    .I0(in[187]),
    .I1(in[176])
  );
  //AND U283bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U283bar (
    .O(n680bar),
    .I0(inbar[187]),
    .I1(inbar[176])
  );
  //OR U284
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U284 (
    .O(n682),
    .I0(n678),
    .I1(n677)
  );
  //AND U284bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U284bar (
    .O(n682bar),
    .I0(n678bar),
    .I1(n677bar)
  );
  //OR U285
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U285 (
    .O(n677),
    .I0(in[245]),
    .I1(in[211])
  );
  //AND U285bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U285bar (
    .O(n677bar),
    .I0(inbar[245]),
    .I1(inbar[211])
  );
  //OR U286
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U286 (
    .O(n678),
    .I0(in[97]),
    .I1(in[88])
  );
  //AND U286bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U286bar (
    .O(n678bar),
    .I0(inbar[97]),
    .I1(inbar[88])
  );
  //OR U287
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U287 (
    .O(n684),
    .I0(n676),
    .I1(n675)
  );
  //AND U287bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U287bar (
    .O(n684bar),
    .I0(n676bar),
    .I1(n675bar)
  );
  //OR U288
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U288 (
    .O(n675),
    .I0(n674),
    .I1(n673)
  );
  //AND U288bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U288bar (
    .O(n675bar),
    .I0(n674bar),
    .I1(n673bar)
  );
  //OR U289
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U289 (
    .O(n673),
    .I0(in_10),
    .I1(in_0)
  );
  //AND U289bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U289bar (
    .O(n673bar),
    .I0(in_10bar),
    .I1(in_0bar)
  );
  //OR U290
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U290 (
    .O(n674),
    .I0(in_59),
    .I1(in_5)
  );
  //AND U290bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U290bar (
    .O(n674bar),
    .I0(in_59bar),
    .I1(in_5bar)
  );
  //OR U291
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U291 (
    .O(n676),
    .I0(n672),
    .I1(n671)
  );
  //AND U291bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U291bar (
    .O(n676bar),
    .I0(n672bar),
    .I1(n671bar)
  );
  //OR U292
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U292 (
    .O(n671),
    .I0(in_60),
    .I1(in_6)
  );
  //AND U292bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U292bar (
    .O(n671bar),
    .I0(in_60bar),
    .I1(in_6bar)
  );
  //OR U293
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U293 (
    .O(n672),
    .I0(in_77),
    .I1(in_69)
  );
  //AND U293bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U293bar (
    .O(n672bar),
    .I0(in_77bar),
    .I1(in_69bar)
  );
  //OR U294
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U294 (
    .O(n700),
    .I0(in[113]),
    .I1(n864)
  );
  //AND U294bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U294bar (
    .O(n700bar),
    .I0(inbar[113]),
    .I1(n864bar)
  );
  //OR U295
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U295 (
    .O(n864),
    .I0(n670),
    .I1(n669)
  );
  //AND U295bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U295bar (
    .O(n864bar),
    .I0(n670bar),
    .I1(n669bar)
  );
  //OR U296
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U296 (
    .O(n669),
    .I0(n668),
    .I1(n667)
  );
  //AND U296bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U296bar (
    .O(n669bar),
    .I0(n668bar),
    .I1(n667bar)
  );
  //OR U297
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U297 (
    .O(n667),
    .I0(n666),
    .I1(n665)
  );
  //AND U297bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U297bar (
    .O(n667bar),
    .I0(n666bar),
    .I1(n665bar)
  );
  //OR U298
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U298 (
    .O(n665),
    .I0(in[125]),
    .I1(in[107])
  );
  //AND U298bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U298bar (
    .O(n665bar),
    .I0(inbar[125]),
    .I1(inbar[107])
  );
  //OR U299
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U299 (
    .O(n666),
    .I0(in[138]),
    .I1(in[126])
  );
  //AND U299bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U299bar (
    .O(n666bar),
    .I0(inbar[138]),
    .I1(inbar[126])
  );
  //OR U300
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U300 (
    .O(n668),
    .I0(n664),
    .I1(n663)
  );
  //AND U300bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U300bar (
    .O(n668bar),
    .I0(n664bar),
    .I1(n663bar)
  );
  //OR U301
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U301 (
    .O(n663),
    .I0(in[189]),
    .I1(in[143])
  );
  //AND U301bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U301bar (
    .O(n663bar),
    .I0(inbar[189]),
    .I1(inbar[143])
  );
  //OR U302
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U302 (
    .O(n664),
    .I0(in[99]),
    .I1(in[214])
  );
  //AND U302bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U302bar (
    .O(n664bar),
    .I0(inbar[99]),
    .I1(inbar[214])
  );
  //OR U303
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U303 (
    .O(n670),
    .I0(n662),
    .I1(n661)
  );
  //AND U303bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U303bar (
    .O(n670bar),
    .I0(n662bar),
    .I1(n661bar)
  );
  //OR U304
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U304 (
    .O(n661),
    .I0(n660),
    .I1(n659)
  );
  //AND U304bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U304bar (
    .O(n661bar),
    .I0(n660bar),
    .I1(n659bar)
  );
  //OR U305
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U305 (
    .O(n659),
    .I0(in_15),
    .I1(in_12)
  );
  //AND U305bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U305bar (
    .O(n659bar),
    .I0(in_15bar),
    .I1(in_12bar)
  );
  //OR U306
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U306 (
    .O(n660),
    .I0(in_20),
    .I1(in_2)
  );
  //AND U306bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U306bar (
    .O(n660bar),
    .I0(in_20bar),
    .I1(in_2bar)
  );
  //OR U307
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U307 (
    .O(n662),
    .I0(n658),
    .I1(n657)
  );
  //AND U307bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U307bar (
    .O(n662bar),
    .I0(n658bar),
    .I1(n657bar)
  );
  //OR U308
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U308 (
    .O(n657),
    .I0(in_30),
    .I1(in_3)
  );
  //AND U308bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U308bar (
    .O(n657bar),
    .I0(in_30bar),
    .I1(in_3bar)
  );
  //OR U309
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U309 (
    .O(n658),
    .I0(in_4),
    .I1(in_38)
  );
  //AND U309bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U309bar (
    .O(n658bar),
    .I0(in_4bar),
    .I1(in_38bar)
  );
  //OR U310
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U310 (
    .O(n702),
    .I0(n656),
    .I1(n655)
  );
  //AND U310bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U310bar (
    .O(n702bar),
    .I0(n656bar),
    .I1(n655bar)
  );
  //OR U311
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U311 (
    .O(n655),
    .I0(in[148]),
    .I1(in[137])
  );
  //AND U311bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U311bar (
    .O(n655bar),
    .I0(inbar[148]),
    .I1(inbar[137])
  );
  //OR U312
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U312 (
    .O(n656),
    .I0(in[149]),
    .I1(n654)
  );
  //AND U312bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U312bar (
    .O(n656bar),
    .I0(inbar[149]),
    .I1(n654bar)
  );
  //OR U313
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U313 (
    .O(n654),
    .I0(in[195]),
    .I1(in[190])
  );
  //AND U313bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U313bar (
    .O(n654bar),
    .I0(inbar[195]),
    .I1(inbar[190])
  );
  //OR U314
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U314 (
    .O(n704),
    .I0(n653),
    .I1(n652)
  );
  //AND U314bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U314bar (
    .O(n704bar),
    .I0(n653bar),
    .I1(n652bar)
  );
  //OR U315
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U315 (
    .O(n652),
    .I0(n651),
    .I1(n650)
  );
  //AND U315bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U315bar (
    .O(n652bar),
    .I0(n651bar),
    .I1(n650bar)
  );
  //OR U316
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U316 (
    .O(n650),
    .I0(in[98]),
    .I1(in[197])
  );
  //AND U316bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U316bar (
    .O(n650bar),
    .I0(inbar[98]),
    .I1(inbar[197])
  );
  //OR U317
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U317 (
    .O(n651),
    .I0(in_11),
    .I1(n649)
  );
  //AND U317bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U317bar (
    .O(n651bar),
    .I0(in_11bar),
    .I1(n649bar)
  );
  //OR U318
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U318 (
    .O(n649),
    .I0(in_26),
    .I1(in_14)
  );
  //AND U318bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U318bar (
    .O(n649bar),
    .I0(in_26bar),
    .I1(in_14bar)
  );
  //OR U319
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U319 (
    .O(n653),
    .I0(n648),
    .I1(n647)
  );
  //AND U319bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U319bar (
    .O(n653bar),
    .I0(n648bar),
    .I1(n647bar)
  );
  //OR U320
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U320 (
    .O(n647),
    .I0(in_35),
    .I1(in_27)
  );
  //AND U320bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U320bar (
    .O(n647bar),
    .I0(in_35bar),
    .I1(in_27bar)
  );
  //OR U321
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U321 (
    .O(n648),
    .I0(in_50),
    .I1(n646)
  );
  //AND U321bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U321bar (
    .O(n648bar),
    .I0(in_50bar),
    .I1(n646bar)
  );
  //OR U322
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U322 (
    .O(n646),
    .I0(in_78),
    .I1(in_61)
  );
  //AND U322bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U322bar (
    .O(n646bar),
    .I0(in_78bar),
    .I1(in_61bar)
  );
  //OR U323
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U323 (
    .O(n720),
    .I0(n942),
    .I1(n645)
  );
  //AND U323bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U323bar (
    .O(n720bar),
    .I0(n942bar),
    .I1(n645bar)
  );
  //OR U324
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U324 (
    .O(n645),
    .I0(in[106]),
    .I1(n863)
  );
  //AND U324bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U324bar (
    .O(n645bar),
    .I0(inbar[106]),
    .I1(n863bar)
  );
  //OR U325
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U325 (
    .O(n863),
    .I0(n644),
    .I1(n643)
  );
  //AND U325bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U325bar (
    .O(n863bar),
    .I0(n644bar),
    .I1(n643bar)
  );
  //OR U326
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U326 (
    .O(n643),
    .I0(n642),
    .I1(n641)
  );
  //AND U326bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U326bar (
    .O(n643bar),
    .I0(n642bar),
    .I1(n641bar)
  );
  //OR U327
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U327 (
    .O(n641),
    .I0(n640),
    .I1(n639)
  );
  //AND U327bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U327bar (
    .O(n641bar),
    .I0(n640bar),
    .I1(n639bar)
  );
  //OR U328
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U328 (
    .O(n639),
    .I0(in[127]),
    .I1(in[122])
  );
  //AND U328bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U328bar (
    .O(n639bar),
    .I0(inbar[127]),
    .I1(inbar[122])
  );
  //OR U329
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U329 (
    .O(n640),
    .I0(in[156]),
    .I1(in[132])
  );
  //AND U329bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U329bar (
    .O(n640bar),
    .I0(inbar[156]),
    .I1(inbar[132])
  );
  //OR U330
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U330 (
    .O(n642),
    .I0(n638),
    .I1(n637)
  );
  //AND U330bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U330bar (
    .O(n642bar),
    .I0(n638bar),
    .I1(n637bar)
  );
  //OR U331
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U331 (
    .O(n637),
    .I0(in[159]),
    .I1(in[157])
  );
  //AND U331bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U331bar (
    .O(n637bar),
    .I0(inbar[159]),
    .I1(inbar[157])
  );
  //OR U332
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U332 (
    .O(n638),
    .I0(in[185]),
    .I1(in[169])
  );
  //AND U332bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U332bar (
    .O(n638bar),
    .I0(inbar[185]),
    .I1(inbar[169])
  );
  //OR U333
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U333 (
    .O(n644),
    .I0(n636),
    .I1(n635)
  );
  //AND U333bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U333bar (
    .O(n644bar),
    .I0(n636bar),
    .I1(n635bar)
  );
  //OR U334
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U334 (
    .O(n635),
    .I0(n634),
    .I1(n633)
  );
  //AND U334bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U334bar (
    .O(n635bar),
    .I0(n634bar),
    .I1(n633bar)
  );
  //OR U335
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U335 (
    .O(n633),
    .I0(in[239]),
    .I1(in[218])
  );
  //AND U335bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U335bar (
    .O(n633bar),
    .I0(inbar[239]),
    .I1(inbar[218])
  );
  //OR U336
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U336 (
    .O(n634),
    .I0(in_13),
    .I1(in[87])
  );
  //AND U336bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U336bar (
    .O(n634bar),
    .I0(in_13bar),
    .I1(inbar[87])
  );
  //OR U337
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U337 (
    .O(n636),
    .I0(n632),
    .I1(n631)
  );
  //AND U337bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U337bar (
    .O(n636bar),
    .I0(n632bar),
    .I1(n631bar)
  );
  //OR U338
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U338 (
    .O(n631),
    .I0(in_72),
    .I1(in_70)
  );
  //AND U338bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U338bar (
    .O(n631bar),
    .I0(in_72bar),
    .I1(in_70bar)
  );
  //OR U339
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U339 (
    .O(n632),
    .I0(in_80),
    .I1(in_74)
  );
  //AND U339bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U339bar (
    .O(n632bar),
    .I0(in_80bar),
    .I1(in_74bar)
  );
  //OR U340
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U340 (
    .O(n942),
    .I0(n630),
    .I1(n629)
  );
  //AND U340bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U340bar (
    .O(n942bar),
    .I0(n630bar),
    .I1(n629bar)
  );
  //OR U341
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U341 (
    .O(n629),
    .I0(n628),
    .I1(n627)
  );
  //AND U341bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U341bar (
    .O(n629bar),
    .I0(n628bar),
    .I1(n627bar)
  );
  //OR U342
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U342 (
    .O(n627),
    .I0(n626),
    .I1(n625)
  );
  //AND U342bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U342bar (
    .O(n627bar),
    .I0(n626bar),
    .I1(n625bar)
  );
  //OR U343
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U343 (
    .O(n625),
    .I0(in[146]),
    .I1(in[100])
  );
  //AND U343bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U343bar (
    .O(n625bar),
    .I0(inbar[146]),
    .I1(inbar[100])
  );
  //OR U344
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U344 (
    .O(n626),
    .I0(in[168]),
    .I1(in[152])
  );
  //AND U344bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U344bar (
    .O(n626bar),
    .I0(inbar[168]),
    .I1(inbar[152])
  );
  //OR U345
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U345 (
    .O(n628),
    .I0(n624),
    .I1(n623)
  );
  //AND U345bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U345bar (
    .O(n628bar),
    .I0(n624bar),
    .I1(n623bar)
  );
  //OR U346
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U346 (
    .O(n623),
    .I0(in[199]),
    .I1(in[182])
  );
  //AND U346bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U346bar (
    .O(n623bar),
    .I0(inbar[199]),
    .I1(inbar[182])
  );
  //OR U347
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U347 (
    .O(n624),
    .I0(in[236]),
    .I1(in[204])
  );
  //AND U347bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U347bar (
    .O(n624bar),
    .I0(inbar[236]),
    .I1(inbar[204])
  );
  //OR U348
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U348 (
    .O(n630),
    .I0(n622),
    .I1(n621)
  );
  //AND U348bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U348bar (
    .O(n630bar),
    .I0(n622bar),
    .I1(n621bar)
  );
  //OR U349
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U349 (
    .O(n621),
    .I0(n620),
    .I1(n619)
  );
  //AND U349bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U349bar (
    .O(n621bar),
    .I0(n620bar),
    .I1(n619bar)
  );
  //OR U350
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U350 (
    .O(n619),
    .I0(in[89]),
    .I1(in[246])
  );
  //AND U350bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U350bar (
    .O(n619bar),
    .I0(inbar[89]),
    .I1(inbar[246])
  );
  //OR U351
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U351 (
    .O(n620),
    .I0(in[95]),
    .I1(in[92])
  );
  //AND U351bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U351bar (
    .O(n620bar),
    .I0(inbar[95]),
    .I1(inbar[92])
  );
  //OR U352
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U352 (
    .O(n622),
    .I0(n618),
    .I1(n617)
  );
  //AND U352bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U352bar (
    .O(n622bar),
    .I0(n618bar),
    .I1(n617bar)
  );
  //OR U353
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U353 (
    .O(n617),
    .I0(in_22),
    .I1(in_16)
  );
  //AND U353bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U353bar (
    .O(n617bar),
    .I0(in_22bar),
    .I1(in_16bar)
  );
  //OR U354
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U354 (
    .O(n618),
    .I0(in_51),
    .I1(in_49)
  );
  //AND U354bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U354bar (
    .O(n618bar),
    .I0(in_51bar),
    .I1(in_49bar)
  );
  //OR U355
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U355 (
    .O(n722),
    .I0(n616),
    .I1(n615)
  );
  //AND U355bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U355bar (
    .O(n722bar),
    .I0(n616bar),
    .I1(n615bar)
  );
  //OR U356
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U356 (
    .O(n615),
    .I0(in[158]),
    .I1(in[115])
  );
  //AND U356bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U356bar (
    .O(n615bar),
    .I0(inbar[158]),
    .I1(inbar[115])
  );
  //OR U357
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U357 (
    .O(n616),
    .I0(in[163]),
    .I1(n614)
  );
  //AND U357bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U357bar (
    .O(n616bar),
    .I0(inbar[163]),
    .I1(n614bar)
  );
  //OR U358
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U358 (
    .O(n614),
    .I0(in[206]),
    .I1(in[165])
  );
  //AND U358bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U358bar (
    .O(n614bar),
    .I0(inbar[206]),
    .I1(inbar[165])
  );
  //OR U359
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U359 (
    .O(n724),
    .I0(n613),
    .I1(n612)
  );
  //AND U359bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U359bar (
    .O(n724bar),
    .I0(n613bar),
    .I1(n612bar)
  );
  //OR U360
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U360 (
    .O(n612),
    .I0(n611),
    .I1(n610)
  );
  //AND U360bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U360bar (
    .O(n612bar),
    .I0(n611bar),
    .I1(n610bar)
  );
  //OR U361
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U361 (
    .O(n610),
    .I0(in[213]),
    .I1(in[207])
  );
  //AND U361bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U361bar (
    .O(n610bar),
    .I0(inbar[213]),
    .I1(inbar[207])
  );
  //OR U362
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U362 (
    .O(n611),
    .I0(in[215]),
    .I1(n609)
  );
  //AND U362bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U362bar (
    .O(n611bar),
    .I0(inbar[215]),
    .I1(n609bar)
  );
  //OR U363
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U363 (
    .O(n609),
    .I0(in[230]),
    .I1(in[220])
  );
  //AND U363bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U363bar (
    .O(n609bar),
    .I0(inbar[230]),
    .I1(inbar[220])
  );
  //OR U364
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U364 (
    .O(n613),
    .I0(n608),
    .I1(n607)
  );
  //AND U364bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U364bar (
    .O(n613bar),
    .I0(n608bar),
    .I1(n607bar)
  );
  //OR U365
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U365 (
    .O(n607),
    .I0(in[251]),
    .I1(in[234])
  );
  //AND U365bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U365bar (
    .O(n607bar),
    .I0(inbar[251]),
    .I1(inbar[234])
  );
  //OR U366
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U366 (
    .O(n608),
    .I0(in_17),
    .I1(n606)
  );
  //AND U366bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U366bar (
    .O(n608bar),
    .I0(in_17bar),
    .I1(n606bar)
  );
  //OR U367
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U367 (
    .O(n606),
    .I0(in_65),
    .I1(in_56)
  );
  //AND U367bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U367bar (
    .O(n606bar),
    .I0(in_65bar),
    .I1(in_56bar)
  );
  //OR U368
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U368 (
    .O(out[0]),
    .I0(n605),
    .I1(n604)
  );
  //AND U368bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U368bar (
    .O(outbar[0]),
    .I0(n605bar),
    .I1(n604bar)
  );
  //OR U369
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U369 (
    .O(n604),
    .I0(n603),
    .I1(n602)
  );
  //AND U369bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U369bar (
    .O(n604bar),
    .I0(n603bar),
    .I1(n602bar)
  );
  //OR U370
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U370 (
    .O(n602),
    .I0(n601),
    .I1(n600)
  );
  //AND U370bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U370bar (
    .O(n602bar),
    .I0(n601bar),
    .I1(n600bar)
  );
  //OR U371
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U371 (
    .O(n600),
    .I0(n820),
    .I1(n785)
  );
  //AND U371bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U371bar (
    .O(n600bar),
    .I0(n820bar),
    .I1(n785bar)
  );
  //OR U372
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U372 (
    .O(n785),
    .I0(n599),
    .I1(n598)
  );
  //AND U372bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U372bar (
    .O(n785bar),
    .I0(n599bar),
    .I1(n598bar)
  );
  //OR U373
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U373 (
    .O(n598),
    .I0(n597),
    .I1(n596)
  );
  //AND U373bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U373bar (
    .O(n598bar),
    .I0(n597bar),
    .I1(n596bar)
  );
  //OR U374
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U374 (
    .O(n596),
    .I0(n595),
    .I1(n594)
  );
  //AND U374bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U374bar (
    .O(n596bar),
    .I0(n595bar),
    .I1(n594bar)
  );
  //OR U375
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U375 (
    .O(n594),
    .I0(in[135]),
    .I1(in[104])
  );
  //AND U375bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U375bar (
    .O(n594bar),
    .I0(inbar[135]),
    .I1(inbar[104])
  );
  //OR U376
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U376 (
    .O(n595),
    .I0(in[188]),
    .I1(in[178])
  );
  //AND U376bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U376bar (
    .O(n595bar),
    .I0(inbar[188]),
    .I1(inbar[178])
  );
  //OR U377
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U377 (
    .O(n597),
    .I0(n593),
    .I1(n592)
  );
  //AND U377bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U377bar (
    .O(n597bar),
    .I0(n593bar),
    .I1(n592bar)
  );
  //OR U378
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U378 (
    .O(n592),
    .I0(in[217]),
    .I1(in[194])
  );
  //AND U378bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U378bar (
    .O(n592bar),
    .I0(inbar[217]),
    .I1(inbar[194])
  );
  //OR U379
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U379 (
    .O(n593),
    .I0(in[237]),
    .I1(in[218])
  );
  //AND U379bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U379bar (
    .O(n593bar),
    .I0(inbar[237]),
    .I1(inbar[218])
  );
  //OR U380
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U380 (
    .O(n599),
    .I0(n591),
    .I1(n590)
  );
  //AND U380bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U380bar (
    .O(n599bar),
    .I0(n591bar),
    .I1(n590bar)
  );
  //OR U381
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U381 (
    .O(n590),
    .I0(n589),
    .I1(n588)
  );
  //AND U381bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U381bar (
    .O(n590bar),
    .I0(n589bar),
    .I1(n588bar)
  );
  //OR U382
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U382 (
    .O(n588),
    .I0(in_2),
    .I1(in_10)
  );
  //AND U382bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U382bar (
    .O(n588bar),
    .I0(in_2bar),
    .I1(in_10bar)
  );
  //OR U383
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U383 (
    .O(n589),
    .I0(in_47),
    .I1(in_22)
  );
  //AND U383bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U383bar (
    .O(n589bar),
    .I0(in_47bar),
    .I1(in_22bar)
  );
  //OR U384
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U384 (
    .O(n591),
    .I0(n587),
    .I1(n586)
  );
  //AND U384bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U384bar (
    .O(n591bar),
    .I0(n587bar),
    .I1(n586bar)
  );
  //OR U385
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U385 (
    .O(n586),
    .I0(in_56),
    .I1(in_54)
  );
  //AND U385bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U385bar (
    .O(n586bar),
    .I0(in_56bar),
    .I1(in_54bar)
  );
  //OR U386
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U386 (
    .O(n587),
    .I0(in_63),
    .I1(in_61)
  );
  //AND U386bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U386bar (
    .O(n587bar),
    .I0(in_63bar),
    .I1(in_61bar)
  );
  //OR U387
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U387 (
    .O(n820),
    .I0(n585),
    .I1(n584)
  );
  //AND U387bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U387bar (
    .O(n820bar),
    .I0(n585bar),
    .I1(n584bar)
  );
  //OR U388
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U388 (
    .O(n584),
    .I0(n583),
    .I1(n582)
  );
  //AND U388bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U388bar (
    .O(n584bar),
    .I0(n583bar),
    .I1(n582bar)
  );
  //OR U389
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U389 (
    .O(n582),
    .I0(n581),
    .I1(n580)
  );
  //AND U389bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U389bar (
    .O(n582bar),
    .I0(n581bar),
    .I1(n580bar)
  );
  //OR U390
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U390 (
    .O(n580),
    .I0(in[158]),
    .I1(in[142])
  );
  //AND U390bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U390bar (
    .O(n580bar),
    .I0(inbar[158]),
    .I1(inbar[142])
  );
  //OR U391
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U391 (
    .O(n581),
    .I0(in[175]),
    .I1(in[164])
  );
  //AND U391bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U391bar (
    .O(n581bar),
    .I0(inbar[175]),
    .I1(inbar[164])
  );
  //OR U392
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U392 (
    .O(n583),
    .I0(n579),
    .I1(n578)
  );
  //AND U392bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U392bar (
    .O(n583bar),
    .I0(n579bar),
    .I1(n578bar)
  );
  //OR U393
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U393 (
    .O(n578),
    .I0(in[228]),
    .I1(in[204])
  );
  //AND U393bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U393bar (
    .O(n578bar),
    .I0(inbar[228]),
    .I1(inbar[204])
  );
  //OR U394
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U394 (
    .O(n579),
    .I0(in[91]),
    .I1(in[87])
  );
  //AND U394bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U394bar (
    .O(n579bar),
    .I0(inbar[91]),
    .I1(inbar[87])
  );
  //OR U395
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U395 (
    .O(n585),
    .I0(n577),
    .I1(n576)
  );
  //AND U395bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U395bar (
    .O(n585bar),
    .I0(n577bar),
    .I1(n576bar)
  );
  //OR U396
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U396 (
    .O(n576),
    .I0(n575),
    .I1(n574)
  );
  //AND U396bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U396bar (
    .O(n576bar),
    .I0(n575bar),
    .I1(n574bar)
  );
  //OR U397
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U397 (
    .O(n574),
    .I0(in_21),
    .I1(in_11)
  );
  //AND U397bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U397bar (
    .O(n574bar),
    .I0(in_21bar),
    .I1(in_11bar)
  );
  //OR U398
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U398 (
    .O(n575),
    .I0(in_5),
    .I1(in_3)
  );
  //AND U398bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U398bar (
    .O(n575bar),
    .I0(in_5bar),
    .I1(in_3bar)
  );
  //OR U399
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U399 (
    .O(n577),
    .I0(n573),
    .I1(n572)
  );
  //AND U399bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U399bar (
    .O(n577bar),
    .I0(n573bar),
    .I1(n572bar)
  );
  //OR U400
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U400 (
    .O(n572),
    .I0(in_68),
    .I1(in_64)
  );
  //AND U400bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U400bar (
    .O(n572bar),
    .I0(in_68bar),
    .I1(in_64bar)
  );
  //OR U401
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U401 (
    .O(n573),
    .I0(in_76),
    .I1(in_73)
  );
  //AND U401bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U401bar (
    .O(n573bar),
    .I0(in_76bar),
    .I1(in_73bar)
  );
  //OR U402
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U402 (
    .O(n601),
    .I0(n778),
    .I1(n571)
  );
  //AND U402bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U402bar (
    .O(n601bar),
    .I0(n778bar),
    .I1(n571bar)
  );
  //OR U403
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U403 (
    .O(n571),
    .I0(in[100]),
    .I1(n965)
  );
  //AND U403bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U403bar (
    .O(n571bar),
    .I0(inbar[100]),
    .I1(n965bar)
  );
  //OR U404
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U404 (
    .O(n965),
    .I0(n570),
    .I1(n569)
  );
  //AND U404bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U404bar (
    .O(n965bar),
    .I0(n570bar),
    .I1(n569bar)
  );
  //OR U405
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U405 (
    .O(n569),
    .I0(n568),
    .I1(n567)
  );
  //AND U405bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U405bar (
    .O(n569bar),
    .I0(n568bar),
    .I1(n567bar)
  );
  //OR U406
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U406 (
    .O(n567),
    .I0(n566),
    .I1(n565)
  );
  //AND U406bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U406bar (
    .O(n567bar),
    .I0(n566bar),
    .I1(n565bar)
  );
  //OR U407
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U407 (
    .O(n565),
    .I0(n817),
    .I1(n750)
  );
  //AND U407bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U407bar (
    .O(n565bar),
    .I0(n817bar),
    .I1(n750bar)
  );
  //OR U408
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U408 (
    .O(n750),
    .I0(n564),
    .I1(n563)
  );
  //AND U408bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U408bar (
    .O(n750bar),
    .I0(n564bar),
    .I1(n563bar)
  );
  //OR U409
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U409 (
    .O(n563),
    .I0(n562),
    .I1(n561)
  );
  //AND U409bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U409bar (
    .O(n563bar),
    .I0(n562bar),
    .I1(n561bar)
  );
  //OR U410
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U410 (
    .O(n561),
    .I0(n560),
    .I1(n559)
  );
  //AND U410bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U410bar (
    .O(n561bar),
    .I0(n560bar),
    .I1(n559bar)
  );
  //OR U411
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U411 (
    .O(n559),
    .I0(in[119]),
    .I1(in[103])
  );
  //AND U411bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U411bar (
    .O(n559bar),
    .I0(inbar[119]),
    .I1(inbar[103])
  );
  //OR U412
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U412 (
    .O(n560),
    .I0(in[137]),
    .I1(in[133])
  );
  //AND U412bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U412bar (
    .O(n560bar),
    .I0(inbar[137]),
    .I1(inbar[133])
  );
  //OR U413
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U413 (
    .O(n562),
    .I0(n558),
    .I1(n557)
  );
  //AND U413bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U413bar (
    .O(n562bar),
    .I0(n558bar),
    .I1(n557bar)
  );
  //OR U414
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U414 (
    .O(n557),
    .I0(in[176]),
    .I1(in[173])
  );
  //AND U414bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U414bar (
    .O(n557bar),
    .I0(inbar[176]),
    .I1(inbar[173])
  );
  //OR U415
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U415 (
    .O(n558),
    .I0(in[210]),
    .I1(in[181])
  );
  //AND U415bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U415bar (
    .O(n558bar),
    .I0(inbar[210]),
    .I1(inbar[181])
  );
  //OR U416
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U416 (
    .O(n564),
    .I0(n556),
    .I1(n555)
  );
  //AND U416bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U416bar (
    .O(n564bar),
    .I0(n556bar),
    .I1(n555bar)
  );
  //OR U417
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U417 (
    .O(n555),
    .I0(n554),
    .I1(n553)
  );
  //AND U417bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U417bar (
    .O(n555bar),
    .I0(n554bar),
    .I1(n553bar)
  );
  //OR U418
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U418 (
    .O(n553),
    .I0(in_13),
    .I1(in[234])
  );
  //AND U418bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U418bar (
    .O(n553bar),
    .I0(in_13bar),
    .I1(inbar[234])
  );
  //OR U419
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U419 (
    .O(n554),
    .I0(in_38),
    .I1(in_32)
  );
  //AND U419bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U419bar (
    .O(n554bar),
    .I0(in_38bar),
    .I1(in_32bar)
  );
  //OR U420
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U420 (
    .O(n556),
    .I0(n552),
    .I1(n551)
  );
  //AND U420bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U420bar (
    .O(n556bar),
    .I0(n552bar),
    .I1(n551bar)
  );
  //OR U421
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U421 (
    .O(n551),
    .I0(in_42),
    .I1(in_41)
  );
  //AND U421bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U421bar (
    .O(n551bar),
    .I0(in_42bar),
    .I1(in_41bar)
  );
  //OR U422
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U422 (
    .O(n552),
    .I0(in_7),
    .I1(in_49)
  );
  //AND U422bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U422bar (
    .O(n552bar),
    .I0(in_7bar),
    .I1(in_49bar)
  );
  //OR U423
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U423 (
    .O(n817),
    .I0(n550),
    .I1(n549)
  );
  //AND U423bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U423bar (
    .O(n817bar),
    .I0(n550bar),
    .I1(n549bar)
  );
  //OR U424
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U424 (
    .O(n549),
    .I0(n548),
    .I1(n547)
  );
  //AND U424bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U424bar (
    .O(n549bar),
    .I0(n548bar),
    .I1(n547bar)
  );
  //OR U425
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U425 (
    .O(n547),
    .I0(n546),
    .I1(n545)
  );
  //AND U425bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U425bar (
    .O(n547bar),
    .I0(n546bar),
    .I1(n545bar)
  );
  //OR U426
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U426 (
    .O(n545),
    .I0(in[159]),
    .I1(in[105])
  );
  //AND U426bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U426bar (
    .O(n545bar),
    .I0(inbar[159]),
    .I1(inbar[105])
  );
  //OR U427
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U427 (
    .O(n546),
    .I0(in[206]),
    .I1(in[183])
  );
  //AND U427bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U427bar (
    .O(n546bar),
    .I0(inbar[206]),
    .I1(inbar[183])
  );
  //OR U428
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U428 (
    .O(n548),
    .I0(n544),
    .I1(n543)
  );
  //AND U428bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U428bar (
    .O(n548bar),
    .I0(n544bar),
    .I1(n543bar)
  );
  //OR U429
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U429 (
    .O(n543),
    .I0(in[229]),
    .I1(in[219])
  );
  //AND U429bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U429bar (
    .O(n543bar),
    .I0(inbar[229]),
    .I1(inbar[219])
  );
  //OR U430
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U430 (
    .O(n544),
    .I0(in[235]),
    .I1(in[232])
  );
  //AND U430bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U430bar (
    .O(n544bar),
    .I0(inbar[235]),
    .I1(inbar[232])
  );
  //OR U431
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U431 (
    .O(n550),
    .I0(n542),
    .I1(n541)
  );
  //AND U431bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U431bar (
    .O(n550bar),
    .I0(n542bar),
    .I1(n541bar)
  );
  //OR U432
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U432 (
    .O(n541),
    .I0(n540),
    .I1(n539)
  );
  //AND U432bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U432bar (
    .O(n541bar),
    .I0(n540bar),
    .I1(n539bar)
  );
  //OR U433
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U433 (
    .O(n539),
    .I0(in[249]),
    .I1(in[242])
  );
  //AND U433bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U433bar (
    .O(n539bar),
    .I0(inbar[249]),
    .I1(inbar[242])
  );
  //OR U434
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U434 (
    .O(n540),
    .I0(in[89]),
    .I1(in[254])
  );
  //AND U434bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U434bar (
    .O(n540bar),
    .I0(inbar[89]),
    .I1(inbar[254])
  );
  //OR U435
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U435 (
    .O(n542),
    .I0(n538),
    .I1(n537)
  );
  //AND U435bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U435bar (
    .O(n542bar),
    .I0(n538bar),
    .I1(n537bar)
  );
  //OR U436
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U436 (
    .O(n537),
    .I0(in_14),
    .I1(in[99])
  );
  //AND U436bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U436bar (
    .O(n537bar),
    .I0(in_14bar),
    .I1(inbar[99])
  );
  //OR U437
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U437 (
    .O(n538),
    .I0(in_60),
    .I1(in_18)
  );
  //AND U437bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U437bar (
    .O(n538bar),
    .I0(in_60bar),
    .I1(in_18bar)
  );
  //OR U438
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U438 (
    .O(n566),
    .I0(in[113]),
    .I1(n763)
  );
  //AND U438bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U438bar (
    .O(n566bar),
    .I0(inbar[113]),
    .I1(n763bar)
  );
  //OR U439
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U439 (
    .O(n763),
    .I0(n536),
    .I1(n535)
  );
  //AND U439bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U439bar (
    .O(n763bar),
    .I0(n536bar),
    .I1(n535bar)
  );
  //OR U440
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U440 (
    .O(n535),
    .I0(n534),
    .I1(n533)
  );
  //AND U440bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U440bar (
    .O(n535bar),
    .I0(n534bar),
    .I1(n533bar)
  );
  //OR U441
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U441 (
    .O(n533),
    .I0(n532),
    .I1(n531)
  );
  //AND U441bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U441bar (
    .O(n533bar),
    .I0(n532bar),
    .I1(n531bar)
  );
  //OR U442
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U442 (
    .O(n531),
    .I0(in[115]),
    .I1(in[110])
  );
  //AND U442bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U442bar (
    .O(n531bar),
    .I0(inbar[115]),
    .I1(inbar[110])
  );
  //OR U443
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U443 (
    .O(n532),
    .I0(in[125]),
    .I1(in[117])
  );
  //AND U443bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U443bar (
    .O(n532bar),
    .I0(inbar[125]),
    .I1(inbar[117])
  );
  //OR U444
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U444 (
    .O(n534),
    .I0(n530),
    .I1(n529)
  );
  //AND U444bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U444bar (
    .O(n534bar),
    .I0(n530bar),
    .I1(n529bar)
  );
  //OR U445
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U445 (
    .O(n529),
    .I0(in[180]),
    .I1(in[128])
  );
  //AND U445bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U445bar (
    .O(n529bar),
    .I0(inbar[180]),
    .I1(inbar[128])
  );
  //OR U446
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U446 (
    .O(n530),
    .I0(in[205]),
    .I1(in[201])
  );
  //AND U446bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U446bar (
    .O(n530bar),
    .I0(inbar[205]),
    .I1(inbar[201])
  );
  //OR U447
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U447 (
    .O(n536),
    .I0(n528),
    .I1(n527)
  );
  //AND U447bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U447bar (
    .O(n536bar),
    .I0(n528bar),
    .I1(n527bar)
  );
  //OR U448
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U448 (
    .O(n527),
    .I0(n526),
    .I1(n525)
  );
  //AND U448bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U448bar (
    .O(n527bar),
    .I0(n526bar),
    .I1(n525bar)
  );
  //OR U449
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U449 (
    .O(n525),
    .I0(in[244]),
    .I1(in[239])
  );
  //AND U449bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U449bar (
    .O(n525bar),
    .I0(inbar[244]),
    .I1(inbar[239])
  );
  //OR U450
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U450 (
    .O(n526),
    .I0(in[95]),
    .I1(in[83])
  );
  //AND U450bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U450bar (
    .O(n526bar),
    .I0(inbar[95]),
    .I1(inbar[83])
  );
  //OR U451
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U451 (
    .O(n528),
    .I0(n524),
    .I1(n523)
  );
  //AND U451bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U451bar (
    .O(n528bar),
    .I0(n524bar),
    .I1(n523bar)
  );
  //OR U452
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U452 (
    .O(n523),
    .I0(in_24),
    .I1(in[97])
  );
  //AND U452bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U452bar (
    .O(n523bar),
    .I0(in_24bar),
    .I1(inbar[97])
  );
  //OR U453
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U453 (
    .O(n524),
    .I0(in_33),
    .I1(in_27)
  );
  //AND U453bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U453bar (
    .O(n524bar),
    .I0(in_33bar),
    .I1(in_27bar)
  );
  //OR U454
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U454 (
    .O(n568),
    .I0(n522),
    .I1(n521)
  );
  //AND U454bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U454bar (
    .O(n568bar),
    .I0(n522bar),
    .I1(n521bar)
  );
  //OR U455
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U455 (
    .O(n521),
    .I0(in[145]),
    .I1(in[126])
  );
  //AND U455bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U455bar (
    .O(n521bar),
    .I0(inbar[145]),
    .I1(inbar[126])
  );
  //OR U456
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U456 (
    .O(n522),
    .I0(in[169]),
    .I1(n520)
  );
  //AND U456bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U456bar (
    .O(n522bar),
    .I0(inbar[169]),
    .I1(n520bar)
  );
  //OR U457
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U457 (
    .O(n520),
    .I0(in[221]),
    .I1(in[172])
  );
  //AND U457bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U457bar (
    .O(n520bar),
    .I0(inbar[221]),
    .I1(inbar[172])
  );
  //OR U458
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U458 (
    .O(n570),
    .I0(n519),
    .I1(n518)
  );
  //AND U458bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U458bar (
    .O(n570bar),
    .I0(n519bar),
    .I1(n518bar)
  );
  //OR U459
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U459 (
    .O(n518),
    .I0(n517),
    .I1(n516)
  );
  //AND U459bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U459bar (
    .O(n518bar),
    .I0(n517bar),
    .I1(n516bar)
  );
  //OR U460
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U460 (
    .O(n516),
    .I0(in[241]),
    .I1(in[224])
  );
  //AND U460bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U460bar (
    .O(n516bar),
    .I0(inbar[241]),
    .I1(inbar[224])
  );
  //OR U461
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U461 (
    .O(n517),
    .I0(in[86]),
    .I1(n515)
  );
  //AND U461bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U461bar (
    .O(n517bar),
    .I0(inbar[86]),
    .I1(n515bar)
  );
  //OR U462
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U462 (
    .O(n515),
    .I0(in_43),
    .I1(in_34)
  );
  //AND U462bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U462bar (
    .O(n515bar),
    .I0(in_43bar),
    .I1(in_34bar)
  );
  //OR U463
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U463 (
    .O(n519),
    .I0(n514),
    .I1(n513)
  );
  //AND U463bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U463bar (
    .O(n519bar),
    .I0(n514bar),
    .I1(n513bar)
  );
  //OR U464
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U464 (
    .O(n513),
    .I0(in_65),
    .I1(in_51)
  );
  //AND U464bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U464bar (
    .O(n513bar),
    .I0(in_65bar),
    .I1(in_51bar)
  );
  //OR U465
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U465 (
    .O(n514),
    .I0(in_75),
    .I1(n512)
  );
  //AND U465bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U465bar (
    .O(n514bar),
    .I0(in_75bar),
    .I1(n512bar)
  );
  //OR U466
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U466 (
    .O(n512),
    .I0(in_81),
    .I1(in_77)
  );
  //AND U466bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U466bar (
    .O(n512bar),
    .I0(in_81bar),
    .I1(in_77bar)
  );
  //OR U467
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U467 (
    .O(n778),
    .I0(n511),
    .I1(n510)
  );
  //AND U467bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U467bar (
    .O(n778bar),
    .I0(n511bar),
    .I1(n510bar)
  );
  //OR U468
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U468 (
    .O(n510),
    .I0(n509),
    .I1(n508)
  );
  //AND U468bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U468bar (
    .O(n510bar),
    .I0(n509bar),
    .I1(n508bar)
  );
  //OR U469
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U469 (
    .O(n508),
    .I0(n507),
    .I1(n506)
  );
  //AND U469bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U469bar (
    .O(n508bar),
    .I0(n507bar),
    .I1(n506bar)
  );
  //OR U470
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U470 (
    .O(n506),
    .I0(in[107]),
    .I1(in[101])
  );
  //AND U470bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U470bar (
    .O(n506bar),
    .I0(inbar[107]),
    .I1(inbar[101])
  );
  //OR U471
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U471 (
    .O(n507),
    .I0(in[139]),
    .I1(in[132])
  );
  //AND U471bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U471bar (
    .O(n507bar),
    .I0(inbar[139]),
    .I1(inbar[132])
  );
  //OR U472
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U472 (
    .O(n509),
    .I0(n505),
    .I1(n504)
  );
  //AND U472bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U472bar (
    .O(n509bar),
    .I0(n505bar),
    .I1(n504bar)
  );
  //OR U473
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U473 (
    .O(n504),
    .I0(in[146]),
    .I1(in[141])
  );
  //AND U473bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U473bar (
    .O(n504bar),
    .I0(inbar[146]),
    .I1(inbar[141])
  );
  //OR U474
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U474 (
    .O(n505),
    .I0(in[203]),
    .I1(in[179])
  );
  //AND U474bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U474bar (
    .O(n505bar),
    .I0(inbar[203]),
    .I1(inbar[179])
  );
  //OR U475
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U475 (
    .O(n511),
    .I0(n503),
    .I1(n502)
  );
  //AND U475bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U475bar (
    .O(n511bar),
    .I0(n503bar),
    .I1(n502bar)
  );
  //OR U476
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U476 (
    .O(n502),
    .I0(n501),
    .I1(n500)
  );
  //AND U476bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U476bar (
    .O(n502bar),
    .I0(n501bar),
    .I1(n500bar)
  );
  //OR U477
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U477 (
    .O(n500),
    .I0(in[243]),
    .I1(in[222])
  );
  //AND U477bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U477bar (
    .O(n500bar),
    .I0(inbar[243]),
    .I1(inbar[222])
  );
  //OR U478
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U478 (
    .O(n501),
    .I0(in[251]),
    .I1(in[250])
  );
  //AND U478bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U478bar (
    .O(n501bar),
    .I0(inbar[251]),
    .I1(inbar[250])
  );
  //OR U479
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U479 (
    .O(n503),
    .I0(n499),
    .I1(n498)
  );
  //AND U479bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U479bar (
    .O(n503bar),
    .I0(n499bar),
    .I1(n498bar)
  );
  //OR U480
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U480 (
    .O(n498),
    .I0(in_37),
    .I1(in_19)
  );
  //AND U480bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U480bar (
    .O(n498bar),
    .I0(in_37bar),
    .I1(in_19bar)
  );
  //OR U481
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U481 (
    .O(n499),
    .I0(in_78),
    .I1(in_6)
  );
  //AND U481bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U481bar (
    .O(n499bar),
    .I0(in_78bar),
    .I1(in_6bar)
  );
  //OR U482
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U482 (
    .O(n603),
    .I0(n497),
    .I1(n496)
  );
  //AND U482bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U482bar (
    .O(n603bar),
    .I0(n497bar),
    .I1(n496bar)
  );
  //OR U483
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U483 (
    .O(n496),
    .I0(in[112]),
    .I1(in[102])
  );
  //AND U483bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U483bar (
    .O(n496bar),
    .I0(inbar[112]),
    .I1(inbar[102])
  );
  //OR U484
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U484 (
    .O(n497),
    .I0(in[123]),
    .I1(n495)
  );
  //AND U484bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U484bar (
    .O(n497bar),
    .I0(inbar[123]),
    .I1(n495bar)
  );
  //OR U485
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U485 (
    .O(n495),
    .I0(in[143]),
    .I1(in[130])
  );
  //AND U485bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U485bar (
    .O(n495bar),
    .I0(inbar[143]),
    .I1(inbar[130])
  );
  //OR U486
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U486 (
    .O(n605),
    .I0(n494),
    .I1(n493)
  );
  //AND U486bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U486bar (
    .O(n605bar),
    .I0(n494bar),
    .I1(n493bar)
  );
  //OR U487
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U487 (
    .O(n493),
    .I0(n492),
    .I1(n491)
  );
  //AND U487bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U487bar (
    .O(n493bar),
    .I0(n492bar),
    .I1(n491bar)
  );
  //OR U488
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U488 (
    .O(n491),
    .I0(in[216]),
    .I1(in[213])
  );
  //AND U488bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U488bar (
    .O(n491bar),
    .I0(inbar[216]),
    .I1(inbar[213])
  );
  //OR U489
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U489 (
    .O(n492),
    .I0(in[227]),
    .I1(n490)
  );
  //AND U489bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U489bar (
    .O(n492bar),
    .I0(inbar[227]),
    .I1(n490bar)
  );
  //OR U490
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U490 (
    .O(n490),
    .I0(in_0),
    .I1(in[248])
  );
  //AND U490bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U490bar (
    .O(n490bar),
    .I0(in_0bar),
    .I1(inbar[248])
  );
  //OR U491
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U491 (
    .O(n494),
    .I0(n489),
    .I1(n488)
  );
  //AND U491bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U491bar (
    .O(n494bar),
    .I0(n489bar),
    .I1(n488bar)
  );
  //OR U492
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U492 (
    .O(n488),
    .I0(in_46),
    .I1(in_44)
  );
  //AND U492bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U492bar (
    .O(n488bar),
    .I0(in_46bar),
    .I1(in_44bar)
  );
  //OR U493
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U493 (
    .O(n489),
    .I0(in_50),
    .I1(n487)
  );
  //AND U493bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U493bar (
    .O(n489bar),
    .I0(in_50bar),
    .I1(n487bar)
  );
  //OR U494
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U494 (
    .O(n487),
    .I0(in_9),
    .I1(in_80)
  );
  //AND U494bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U494bar (
    .O(n487bar),
    .I0(in_9bar),
    .I1(in_80bar)
  );
endmodule

module sBox_13 ( in, out );

  input wire [7:0] in;
//input_done

  output wire [7:0] out;
//output_done

  wire [255:0] decodeOut;
//wire_done

  decode_13 dec ( .in(in), .out(decodeOut) );
  encode_13 enc ( .in(decodeOut), .out(out) );
endmodule

module CD2_53 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD2_54 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD2_55 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD2_56 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD4_27 ( a, b, y );

  input wire [3:0] a;
  input wire [3:0] b;
  wire [3:0] abar;
  wire [3:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
//input_done

  output wire [15:0] y;
  wire [15:0] ybar;
//output_done

//wire_done

  //AND U1
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1 (
    .O(y[9]),
    .I0(b[1]),
    .I1(a[2])
  );
  //OR U1bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1bar (
    .O(ybar[9]),
    .I0(bbar[1]),
    .I1(abar[2])
  );
  //AND U2
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2 (
    .O(y[8]),
    .I0(b[0]),
    .I1(a[2])
  );
  //OR U2bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2bar (
    .O(ybar[8]),
    .I0(bbar[0]),
    .I1(abar[2])
  );
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[7]),
    .I0(b[3]),
    .I1(a[1])
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[7]),
    .I0(bbar[3]),
    .I1(abar[1])
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[6]),
    .I0(b[2]),
    .I1(a[1])
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[6]),
    .I0(bbar[2]),
    .I1(abar[1])
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[5]),
    .I0(a[1]),
    .I1(b[1])
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[5]),
    .I0(abar[1]),
    .I1(bbar[1])
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[4]),
    .I0(a[1]),
    .I1(b[0])
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[4]),
    .I0(abar[1]),
    .I1(bbar[0])
  );
  //AND U7
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7 (
    .O(y[3]),
    .I0(a[0]),
    .I1(b[3])
  );
  //OR U7bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7bar (
    .O(ybar[3]),
    .I0(abar[0]),
    .I1(bbar[3])
  );
  //AND U8
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8 (
    .O(y[2]),
    .I0(a[0]),
    .I1(b[2])
  );
  //OR U8bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8bar (
    .O(ybar[2]),
    .I0(abar[0]),
    .I1(bbar[2])
  );
  //AND U9
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9 (
    .O(y[1]),
    .I0(a[0]),
    .I1(b[1])
  );
  //OR U9bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9bar (
    .O(ybar[1]),
    .I0(abar[0]),
    .I1(bbar[1])
  );
  //AND U10
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10 (
    .O(y[15]),
    .I0(a[3]),
    .I1(b[3])
  );
  //OR U10bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10bar (
    .O(ybar[15]),
    .I0(abar[3]),
    .I1(bbar[3])
  );
  //AND U11
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11 (
    .O(y[14]),
    .I0(a[3]),
    .I1(b[2])
  );
  //OR U11bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11bar (
    .O(ybar[14]),
    .I0(abar[3]),
    .I1(bbar[2])
  );
  //AND U12
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12 (
    .O(y[13]),
    .I0(a[3]),
    .I1(b[1])
  );
  //OR U12bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12bar (
    .O(ybar[13]),
    .I0(abar[3]),
    .I1(bbar[1])
  );
  //AND U13
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13 (
    .O(y[12]),
    .I0(a[3]),
    .I1(b[0])
  );
  //OR U13bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13bar (
    .O(ybar[12]),
    .I0(abar[3]),
    .I1(bbar[0])
  );
  //AND U14
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14 (
    .O(y[11]),
    .I0(b[3]),
    .I1(a[2])
  );
  //OR U14bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14bar (
    .O(ybar[11]),
    .I0(bbar[3]),
    .I1(abar[2])
  );
  //AND U15
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15 (
    .O(y[10]),
    .I0(b[2]),
    .I1(a[2])
  );
  //OR U15bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15bar (
    .O(ybar[10]),
    .I0(bbar[2]),
    .I1(abar[2])
  );
  //AND U16
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16 (
    .O(y[0]),
    .I0(a[0]),
    .I1(b[0])
  );
  //OR U16bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16bar (
    .O(ybar[0]),
    .I0(abar[0]),
    .I1(bbar[0])
  );
endmodule

module CD4_28 ( a, b, y );

  input wire [3:0] a;
  input wire [3:0] b;
  wire [3:0] abar;
  wire [3:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
//input_done

  output wire [15:0] y;
  wire [15:0] ybar;
//output_done

//wire_done

  //AND U1
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1 (
    .O(y[9]),
    .I0(b[1]),
    .I1(a[2])
  );
  //OR U1bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1bar (
    .O(ybar[9]),
    .I0(bbar[1]),
    .I1(abar[2])
  );
  //AND U2
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2 (
    .O(y[8]),
    .I0(b[0]),
    .I1(a[2])
  );
  //OR U2bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2bar (
    .O(ybar[8]),
    .I0(bbar[0]),
    .I1(abar[2])
  );
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[7]),
    .I0(b[3]),
    .I1(a[1])
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[7]),
    .I0(bbar[3]),
    .I1(abar[1])
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[6]),
    .I0(b[2]),
    .I1(a[1])
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[6]),
    .I0(bbar[2]),
    .I1(abar[1])
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[5]),
    .I0(a[1]),
    .I1(b[1])
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[5]),
    .I0(abar[1]),
    .I1(bbar[1])
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[4]),
    .I0(a[1]),
    .I1(b[0])
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[4]),
    .I0(abar[1]),
    .I1(bbar[0])
  );
  //AND U7
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7 (
    .O(y[3]),
    .I0(a[0]),
    .I1(b[3])
  );
  //OR U7bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7bar (
    .O(ybar[3]),
    .I0(abar[0]),
    .I1(bbar[3])
  );
  //AND U8
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8 (
    .O(y[2]),
    .I0(a[0]),
    .I1(b[2])
  );
  //OR U8bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8bar (
    .O(ybar[2]),
    .I0(abar[0]),
    .I1(bbar[2])
  );
  //AND U9
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9 (
    .O(y[1]),
    .I0(a[0]),
    .I1(b[1])
  );
  //OR U9bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9bar (
    .O(ybar[1]),
    .I0(abar[0]),
    .I1(bbar[1])
  );
  //AND U10
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10 (
    .O(y[15]),
    .I0(a[3]),
    .I1(b[3])
  );
  //OR U10bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10bar (
    .O(ybar[15]),
    .I0(abar[3]),
    .I1(bbar[3])
  );
  //AND U11
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11 (
    .O(y[14]),
    .I0(a[3]),
    .I1(b[2])
  );
  //OR U11bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11bar (
    .O(ybar[14]),
    .I0(abar[3]),
    .I1(bbar[2])
  );
  //AND U12
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12 (
    .O(y[13]),
    .I0(a[3]),
    .I1(b[1])
  );
  //OR U12bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12bar (
    .O(ybar[13]),
    .I0(abar[3]),
    .I1(bbar[1])
  );
  //AND U13
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13 (
    .O(y[12]),
    .I0(a[3]),
    .I1(b[0])
  );
  //OR U13bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13bar (
    .O(ybar[12]),
    .I0(abar[3]),
    .I1(bbar[0])
  );
  //AND U14
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14 (
    .O(y[11]),
    .I0(b[3]),
    .I1(a[2])
  );
  //OR U14bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14bar (
    .O(ybar[11]),
    .I0(bbar[3]),
    .I1(abar[2])
  );
  //AND U15
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15 (
    .O(y[10]),
    .I0(b[2]),
    .I1(a[2])
  );
  //OR U15bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15bar (
    .O(ybar[10]),
    .I0(bbar[2]),
    .I1(abar[2])
  );
  //AND U16
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16 (
    .O(y[0]),
    .I0(a[0]),
    .I1(b[0])
  );
  //OR U16bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16bar (
    .O(ybar[0]),
    .I0(abar[0]),
    .I1(bbar[0])
  );
endmodule

module CD16_14 ( a, b, y );

  input wire [15:0] a;
  input wire [15:0] b;
  wire [15:0] abar;
  wire [15:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign abar[8] = ~a[8];
  assign abar[9] = ~a[9];
  assign abar[10] = ~a[10];
  assign abar[11] = ~a[11];
  assign abar[12] = ~a[12];
  assign abar[13] = ~a[13];
  assign abar[14] = ~a[14];
  assign abar[15] = ~a[15];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign bbar[8] = ~b[8];
  assign bbar[9] = ~b[9];
  assign bbar[10] = ~b[10];
  assign bbar[11] = ~b[11];
  assign bbar[12] = ~b[12];
  assign bbar[13] = ~b[13];
  assign bbar[14] = ~b[14];
  assign bbar[15] = ~b[15];
//input_done

  output wire [255:0] y;
  wire [255:0] ybar;
//output_done

//wire_done

  //AND U1
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1 (
    .O(y[9]),
    .I0(b[9]),
    .I1(a[0])
  );
  //OR U1bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1bar (
    .O(ybar[9]),
    .I0(bbar[9]),
    .I1(abar[0])
  );
  //AND U2
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2 (
    .O(y[99]),
    .I0(b[3]),
    .I1(a[6])
  );
  //OR U2bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2bar (
    .O(ybar[99]),
    .I0(bbar[3]),
    .I1(abar[6])
  );
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[98]),
    .I0(b[2]),
    .I1(a[6])
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[98]),
    .I0(bbar[2]),
    .I1(abar[6])
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[97]),
    .I0(b[1]),
    .I1(a[6])
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[97]),
    .I0(bbar[1]),
    .I1(abar[6])
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[96]),
    .I0(b[0]),
    .I1(a[6])
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[96]),
    .I0(bbar[0]),
    .I1(abar[6])
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[95]),
    .I0(b[15]),
    .I1(a[5])
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[95]),
    .I0(bbar[15]),
    .I1(abar[5])
  );
  //AND U7
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7 (
    .O(y[94]),
    .I0(b[14]),
    .I1(a[5])
  );
  //OR U7bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7bar (
    .O(ybar[94]),
    .I0(bbar[14]),
    .I1(abar[5])
  );
  //AND U8
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8 (
    .O(y[93]),
    .I0(b[13]),
    .I1(a[5])
  );
  //OR U8bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8bar (
    .O(ybar[93]),
    .I0(bbar[13]),
    .I1(abar[5])
  );
  //AND U9
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9 (
    .O(y[92]),
    .I0(b[12]),
    .I1(a[5])
  );
  //OR U9bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9bar (
    .O(ybar[92]),
    .I0(bbar[12]),
    .I1(abar[5])
  );
  //AND U10
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10 (
    .O(y[91]),
    .I0(b[11]),
    .I1(a[5])
  );
  //OR U10bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10bar (
    .O(ybar[91]),
    .I0(bbar[11]),
    .I1(abar[5])
  );
  //AND U11
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11 (
    .O(y[90]),
    .I0(b[10]),
    .I1(a[5])
  );
  //OR U11bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11bar (
    .O(ybar[90]),
    .I0(bbar[10]),
    .I1(abar[5])
  );
  //AND U12
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12 (
    .O(y[8]),
    .I0(b[8]),
    .I1(a[0])
  );
  //OR U12bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12bar (
    .O(ybar[8]),
    .I0(bbar[8]),
    .I1(abar[0])
  );
  //AND U13
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13 (
    .O(y[89]),
    .I0(a[5]),
    .I1(b[9])
  );
  //OR U13bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13bar (
    .O(ybar[89]),
    .I0(abar[5]),
    .I1(bbar[9])
  );
  //AND U14
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14 (
    .O(y[88]),
    .I0(b[8]),
    .I1(a[5])
  );
  //OR U14bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14bar (
    .O(ybar[88]),
    .I0(bbar[8]),
    .I1(abar[5])
  );
  //AND U15
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15 (
    .O(y[87]),
    .I0(b[7]),
    .I1(a[5])
  );
  //OR U15bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15bar (
    .O(ybar[87]),
    .I0(bbar[7]),
    .I1(abar[5])
  );
  //AND U16
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16 (
    .O(y[86]),
    .I0(b[6]),
    .I1(a[5])
  );
  //OR U16bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16bar (
    .O(ybar[86]),
    .I0(bbar[6]),
    .I1(abar[5])
  );
  //AND U17
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U17 (
    .O(y[85]),
    .I0(b[5]),
    .I1(a[5])
  );
  //OR U17bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U17bar (
    .O(ybar[85]),
    .I0(bbar[5]),
    .I1(abar[5])
  );
  //AND U18
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U18 (
    .O(y[84]),
    .I0(b[4]),
    .I1(a[5])
  );
  //OR U18bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U18bar (
    .O(ybar[84]),
    .I0(bbar[4]),
    .I1(abar[5])
  );
  //AND U19
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U19 (
    .O(y[83]),
    .I0(a[5]),
    .I1(b[3])
  );
  //OR U19bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U19bar (
    .O(ybar[83]),
    .I0(abar[5]),
    .I1(bbar[3])
  );
  //AND U20
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U20 (
    .O(y[82]),
    .I0(a[5]),
    .I1(b[2])
  );
  //OR U20bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U20bar (
    .O(ybar[82]),
    .I0(abar[5]),
    .I1(bbar[2])
  );
  //AND U21
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U21 (
    .O(y[81]),
    .I0(a[5]),
    .I1(b[1])
  );
  //OR U21bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U21bar (
    .O(ybar[81]),
    .I0(abar[5]),
    .I1(bbar[1])
  );
  //AND U22
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U22 (
    .O(y[80]),
    .I0(a[5]),
    .I1(b[0])
  );
  //OR U22bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U22bar (
    .O(ybar[80]),
    .I0(abar[5]),
    .I1(bbar[0])
  );
  //AND U23
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U23 (
    .O(y[7]),
    .I0(b[7]),
    .I1(a[0])
  );
  //OR U23bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U23bar (
    .O(ybar[7]),
    .I0(bbar[7]),
    .I1(abar[0])
  );
  //AND U24
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U24 (
    .O(y[79]),
    .I0(a[4]),
    .I1(b[15])
  );
  //OR U24bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U24bar (
    .O(ybar[79]),
    .I0(abar[4]),
    .I1(bbar[15])
  );
  //AND U25
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U25 (
    .O(y[78]),
    .I0(a[4]),
    .I1(b[14])
  );
  //OR U25bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U25bar (
    .O(ybar[78]),
    .I0(abar[4]),
    .I1(bbar[14])
  );
  //AND U26
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U26 (
    .O(y[77]),
    .I0(a[4]),
    .I1(b[13])
  );
  //OR U26bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U26bar (
    .O(ybar[77]),
    .I0(abar[4]),
    .I1(bbar[13])
  );
  //AND U27
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U27 (
    .O(y[76]),
    .I0(a[4]),
    .I1(b[12])
  );
  //OR U27bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U27bar (
    .O(ybar[76]),
    .I0(abar[4]),
    .I1(bbar[12])
  );
  //AND U28
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U28 (
    .O(y[75]),
    .I0(a[4]),
    .I1(b[11])
  );
  //OR U28bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U28bar (
    .O(ybar[75]),
    .I0(abar[4]),
    .I1(bbar[11])
  );
  //AND U29
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U29 (
    .O(y[74]),
    .I0(a[4]),
    .I1(b[10])
  );
  //OR U29bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U29bar (
    .O(ybar[74]),
    .I0(abar[4]),
    .I1(bbar[10])
  );
  //AND U30
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U30 (
    .O(y[73]),
    .I0(a[4]),
    .I1(b[9])
  );
  //OR U30bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U30bar (
    .O(ybar[73]),
    .I0(abar[4]),
    .I1(bbar[9])
  );
  //AND U31
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U31 (
    .O(y[72]),
    .I0(a[4]),
    .I1(b[8])
  );
  //OR U31bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U31bar (
    .O(ybar[72]),
    .I0(abar[4]),
    .I1(bbar[8])
  );
  //AND U32
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U32 (
    .O(y[71]),
    .I0(a[4]),
    .I1(b[7])
  );
  //OR U32bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U32bar (
    .O(ybar[71]),
    .I0(abar[4]),
    .I1(bbar[7])
  );
  //AND U33
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U33 (
    .O(y[70]),
    .I0(a[4]),
    .I1(b[6])
  );
  //OR U33bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U33bar (
    .O(ybar[70]),
    .I0(abar[4]),
    .I1(bbar[6])
  );
  //AND U34
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U34 (
    .O(y[6]),
    .I0(b[6]),
    .I1(a[0])
  );
  //OR U34bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U34bar (
    .O(ybar[6]),
    .I0(bbar[6]),
    .I1(abar[0])
  );
  //AND U35
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U35 (
    .O(y[69]),
    .I0(a[4]),
    .I1(b[5])
  );
  //OR U35bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U35bar (
    .O(ybar[69]),
    .I0(abar[4]),
    .I1(bbar[5])
  );
  //AND U36
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U36 (
    .O(y[68]),
    .I0(a[4]),
    .I1(b[4])
  );
  //OR U36bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U36bar (
    .O(ybar[68]),
    .I0(abar[4]),
    .I1(bbar[4])
  );
  //AND U37
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U37 (
    .O(y[67]),
    .I0(a[4]),
    .I1(b[3])
  );
  //OR U37bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U37bar (
    .O(ybar[67]),
    .I0(abar[4]),
    .I1(bbar[3])
  );
  //AND U38
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U38 (
    .O(y[66]),
    .I0(a[4]),
    .I1(b[2])
  );
  //OR U38bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U38bar (
    .O(ybar[66]),
    .I0(abar[4]),
    .I1(bbar[2])
  );
  //AND U39
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U39 (
    .O(y[65]),
    .I0(a[4]),
    .I1(b[1])
  );
  //OR U39bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U39bar (
    .O(ybar[65]),
    .I0(abar[4]),
    .I1(bbar[1])
  );
  //AND U40
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U40 (
    .O(y[64]),
    .I0(a[4]),
    .I1(b[0])
  );
  //OR U40bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U40bar (
    .O(ybar[64]),
    .I0(abar[4]),
    .I1(bbar[0])
  );
  //AND U41
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U41 (
    .O(y[63]),
    .I0(a[3]),
    .I1(b[15])
  );
  //OR U41bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U41bar (
    .O(ybar[63]),
    .I0(abar[3]),
    .I1(bbar[15])
  );
  //AND U42
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U42 (
    .O(y[62]),
    .I0(a[3]),
    .I1(b[14])
  );
  //OR U42bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U42bar (
    .O(ybar[62]),
    .I0(abar[3]),
    .I1(bbar[14])
  );
  //AND U43
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U43 (
    .O(y[61]),
    .I0(a[3]),
    .I1(b[13])
  );
  //OR U43bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U43bar (
    .O(ybar[61]),
    .I0(abar[3]),
    .I1(bbar[13])
  );
  //AND U44
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U44 (
    .O(y[60]),
    .I0(a[3]),
    .I1(b[12])
  );
  //OR U44bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U44bar (
    .O(ybar[60]),
    .I0(abar[3]),
    .I1(bbar[12])
  );
  //AND U45
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U45 (
    .O(y[5]),
    .I0(b[5]),
    .I1(a[0])
  );
  //OR U45bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U45bar (
    .O(ybar[5]),
    .I0(bbar[5]),
    .I1(abar[0])
  );
  //AND U46
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U46 (
    .O(y[59]),
    .I0(a[3]),
    .I1(b[11])
  );
  //OR U46bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U46bar (
    .O(ybar[59]),
    .I0(abar[3]),
    .I1(bbar[11])
  );
  //AND U47
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U47 (
    .O(y[58]),
    .I0(a[3]),
    .I1(b[10])
  );
  //OR U47bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U47bar (
    .O(ybar[58]),
    .I0(abar[3]),
    .I1(bbar[10])
  );
  //AND U48
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U48 (
    .O(y[57]),
    .I0(a[3]),
    .I1(b[9])
  );
  //OR U48bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U48bar (
    .O(ybar[57]),
    .I0(abar[3]),
    .I1(bbar[9])
  );
  //AND U49
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U49 (
    .O(y[56]),
    .I0(a[3]),
    .I1(b[8])
  );
  //OR U49bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U49bar (
    .O(ybar[56]),
    .I0(abar[3]),
    .I1(bbar[8])
  );
  //AND U50
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U50 (
    .O(y[55]),
    .I0(a[3]),
    .I1(b[7])
  );
  //OR U50bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U50bar (
    .O(ybar[55]),
    .I0(abar[3]),
    .I1(bbar[7])
  );
  //AND U51
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U51 (
    .O(y[54]),
    .I0(a[3]),
    .I1(b[6])
  );
  //OR U51bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U51bar (
    .O(ybar[54]),
    .I0(abar[3]),
    .I1(bbar[6])
  );
  //AND U52
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U52 (
    .O(y[53]),
    .I0(a[3]),
    .I1(b[5])
  );
  //OR U52bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U52bar (
    .O(ybar[53]),
    .I0(abar[3]),
    .I1(bbar[5])
  );
  //AND U53
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U53 (
    .O(y[52]),
    .I0(a[3]),
    .I1(b[4])
  );
  //OR U53bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U53bar (
    .O(ybar[52]),
    .I0(abar[3]),
    .I1(bbar[4])
  );
  //AND U54
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U54 (
    .O(y[51]),
    .I0(a[3]),
    .I1(b[3])
  );
  //OR U54bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U54bar (
    .O(ybar[51]),
    .I0(abar[3]),
    .I1(bbar[3])
  );
  //AND U55
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U55 (
    .O(y[50]),
    .I0(a[3]),
    .I1(b[2])
  );
  //OR U55bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U55bar (
    .O(ybar[50]),
    .I0(abar[3]),
    .I1(bbar[2])
  );
  //AND U56
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U56 (
    .O(y[4]),
    .I0(b[4]),
    .I1(a[0])
  );
  //OR U56bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U56bar (
    .O(ybar[4]),
    .I0(bbar[4]),
    .I1(abar[0])
  );
  //AND U57
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U57 (
    .O(y[49]),
    .I0(a[3]),
    .I1(b[1])
  );
  //OR U57bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U57bar (
    .O(ybar[49]),
    .I0(abar[3]),
    .I1(bbar[1])
  );
  //AND U58
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U58 (
    .O(y[48]),
    .I0(a[3]),
    .I1(b[0])
  );
  //OR U58bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U58bar (
    .O(ybar[48]),
    .I0(abar[3]),
    .I1(bbar[0])
  );
  //AND U59
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U59 (
    .O(y[47]),
    .I0(a[2]),
    .I1(b[15])
  );
  //OR U59bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U59bar (
    .O(ybar[47]),
    .I0(abar[2]),
    .I1(bbar[15])
  );
  //AND U60
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U60 (
    .O(y[46]),
    .I0(a[2]),
    .I1(b[14])
  );
  //OR U60bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U60bar (
    .O(ybar[46]),
    .I0(abar[2]),
    .I1(bbar[14])
  );
  //AND U61
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U61 (
    .O(y[45]),
    .I0(a[2]),
    .I1(b[13])
  );
  //OR U61bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U61bar (
    .O(ybar[45]),
    .I0(abar[2]),
    .I1(bbar[13])
  );
  //AND U62
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U62 (
    .O(y[44]),
    .I0(a[2]),
    .I1(b[12])
  );
  //OR U62bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U62bar (
    .O(ybar[44]),
    .I0(abar[2]),
    .I1(bbar[12])
  );
  //AND U63
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U63 (
    .O(y[43]),
    .I0(a[2]),
    .I1(b[11])
  );
  //OR U63bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U63bar (
    .O(ybar[43]),
    .I0(abar[2]),
    .I1(bbar[11])
  );
  //AND U64
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U64 (
    .O(y[42]),
    .I0(a[2]),
    .I1(b[10])
  );
  //OR U64bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U64bar (
    .O(ybar[42]),
    .I0(abar[2]),
    .I1(bbar[10])
  );
  //AND U65
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U65 (
    .O(y[41]),
    .I0(a[2]),
    .I1(b[9])
  );
  //OR U65bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U65bar (
    .O(ybar[41]),
    .I0(abar[2]),
    .I1(bbar[9])
  );
  //AND U66
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U66 (
    .O(y[40]),
    .I0(a[2]),
    .I1(b[8])
  );
  //OR U66bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U66bar (
    .O(ybar[40]),
    .I0(abar[2]),
    .I1(bbar[8])
  );
  //AND U67
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U67 (
    .O(y[3]),
    .I0(b[3]),
    .I1(a[0])
  );
  //OR U67bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U67bar (
    .O(ybar[3]),
    .I0(bbar[3]),
    .I1(abar[0])
  );
  //AND U68
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U68 (
    .O(y[39]),
    .I0(a[2]),
    .I1(b[7])
  );
  //OR U68bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U68bar (
    .O(ybar[39]),
    .I0(abar[2]),
    .I1(bbar[7])
  );
  //AND U69
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U69 (
    .O(y[38]),
    .I0(a[2]),
    .I1(b[6])
  );
  //OR U69bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U69bar (
    .O(ybar[38]),
    .I0(abar[2]),
    .I1(bbar[6])
  );
  //AND U70
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U70 (
    .O(y[37]),
    .I0(a[2]),
    .I1(b[5])
  );
  //OR U70bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U70bar (
    .O(ybar[37]),
    .I0(abar[2]),
    .I1(bbar[5])
  );
  //AND U71
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U71 (
    .O(y[36]),
    .I0(a[2]),
    .I1(b[4])
  );
  //OR U71bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U71bar (
    .O(ybar[36]),
    .I0(abar[2]),
    .I1(bbar[4])
  );
  //AND U72
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U72 (
    .O(y[35]),
    .I0(a[2]),
    .I1(b[3])
  );
  //OR U72bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U72bar (
    .O(ybar[35]),
    .I0(abar[2]),
    .I1(bbar[3])
  );
  //AND U73
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U73 (
    .O(y[34]),
    .I0(a[2]),
    .I1(b[2])
  );
  //OR U73bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U73bar (
    .O(ybar[34]),
    .I0(abar[2]),
    .I1(bbar[2])
  );
  //AND U74
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U74 (
    .O(y[33]),
    .I0(a[2]),
    .I1(b[1])
  );
  //OR U74bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U74bar (
    .O(ybar[33]),
    .I0(abar[2]),
    .I1(bbar[1])
  );
  //AND U75
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U75 (
    .O(y[32]),
    .I0(a[2]),
    .I1(b[0])
  );
  //OR U75bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U75bar (
    .O(ybar[32]),
    .I0(abar[2]),
    .I1(bbar[0])
  );
  //AND U76
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U76 (
    .O(y[31]),
    .I0(a[1]),
    .I1(b[15])
  );
  //OR U76bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U76bar (
    .O(ybar[31]),
    .I0(abar[1]),
    .I1(bbar[15])
  );
  //AND U77
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U77 (
    .O(y[30]),
    .I0(a[1]),
    .I1(b[14])
  );
  //OR U77bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U77bar (
    .O(ybar[30]),
    .I0(abar[1]),
    .I1(bbar[14])
  );
  //AND U78
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U78 (
    .O(y[2]),
    .I0(b[2]),
    .I1(a[0])
  );
  //OR U78bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U78bar (
    .O(ybar[2]),
    .I0(bbar[2]),
    .I1(abar[0])
  );
  //AND U79
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U79 (
    .O(y[29]),
    .I0(a[1]),
    .I1(b[13])
  );
  //OR U79bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U79bar (
    .O(ybar[29]),
    .I0(abar[1]),
    .I1(bbar[13])
  );
  //AND U80
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U80 (
    .O(y[28]),
    .I0(a[1]),
    .I1(b[12])
  );
  //OR U80bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U80bar (
    .O(ybar[28]),
    .I0(abar[1]),
    .I1(bbar[12])
  );
  //AND U81
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U81 (
    .O(y[27]),
    .I0(a[1]),
    .I1(b[11])
  );
  //OR U81bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U81bar (
    .O(ybar[27]),
    .I0(abar[1]),
    .I1(bbar[11])
  );
  //AND U82
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U82 (
    .O(y[26]),
    .I0(a[1]),
    .I1(b[10])
  );
  //OR U82bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U82bar (
    .O(ybar[26]),
    .I0(abar[1]),
    .I1(bbar[10])
  );
  //AND U83
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U83 (
    .O(y[25]),
    .I0(a[1]),
    .I1(b[9])
  );
  //OR U83bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U83bar (
    .O(ybar[25]),
    .I0(abar[1]),
    .I1(bbar[9])
  );
  //AND U84
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U84 (
    .O(y[255]),
    .I0(a[15]),
    .I1(b[15])
  );
  //OR U84bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U84bar (
    .O(ybar[255]),
    .I0(abar[15]),
    .I1(bbar[15])
  );
  //AND U85
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U85 (
    .O(y[254]),
    .I0(a[15]),
    .I1(b[14])
  );
  //OR U85bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U85bar (
    .O(ybar[254]),
    .I0(abar[15]),
    .I1(bbar[14])
  );
  //AND U86
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U86 (
    .O(y[253]),
    .I0(a[15]),
    .I1(b[13])
  );
  //OR U86bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U86bar (
    .O(ybar[253]),
    .I0(abar[15]),
    .I1(bbar[13])
  );
  //AND U87
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U87 (
    .O(y[252]),
    .I0(a[15]),
    .I1(b[12])
  );
  //OR U87bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U87bar (
    .O(ybar[252]),
    .I0(abar[15]),
    .I1(bbar[12])
  );
  //AND U88
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U88 (
    .O(y[251]),
    .I0(a[15]),
    .I1(b[11])
  );
  //OR U88bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U88bar (
    .O(ybar[251]),
    .I0(abar[15]),
    .I1(bbar[11])
  );
  //AND U89
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U89 (
    .O(y[250]),
    .I0(a[15]),
    .I1(b[10])
  );
  //OR U89bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U89bar (
    .O(ybar[250]),
    .I0(abar[15]),
    .I1(bbar[10])
  );
  //AND U90
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U90 (
    .O(y[24]),
    .I0(a[1]),
    .I1(b[8])
  );
  //OR U90bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U90bar (
    .O(ybar[24]),
    .I0(abar[1]),
    .I1(bbar[8])
  );
  //AND U91
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U91 (
    .O(y[249]),
    .I0(a[15]),
    .I1(b[9])
  );
  //OR U91bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U91bar (
    .O(ybar[249]),
    .I0(abar[15]),
    .I1(bbar[9])
  );
  //AND U92
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U92 (
    .O(y[248]),
    .I0(a[15]),
    .I1(b[8])
  );
  //OR U92bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U92bar (
    .O(ybar[248]),
    .I0(abar[15]),
    .I1(bbar[8])
  );
  //AND U93
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U93 (
    .O(y[247]),
    .I0(a[15]),
    .I1(b[7])
  );
  //OR U93bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U93bar (
    .O(ybar[247]),
    .I0(abar[15]),
    .I1(bbar[7])
  );
  //AND U94
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U94 (
    .O(y[246]),
    .I0(a[15]),
    .I1(b[6])
  );
  //OR U94bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U94bar (
    .O(ybar[246]),
    .I0(abar[15]),
    .I1(bbar[6])
  );
  //AND U95
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U95 (
    .O(y[245]),
    .I0(a[15]),
    .I1(b[5])
  );
  //OR U95bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U95bar (
    .O(ybar[245]),
    .I0(abar[15]),
    .I1(bbar[5])
  );
  //AND U96
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U96 (
    .O(y[244]),
    .I0(a[15]),
    .I1(b[4])
  );
  //OR U96bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U96bar (
    .O(ybar[244]),
    .I0(abar[15]),
    .I1(bbar[4])
  );
  //AND U97
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U97 (
    .O(y[243]),
    .I0(a[15]),
    .I1(b[3])
  );
  //OR U97bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U97bar (
    .O(ybar[243]),
    .I0(abar[15]),
    .I1(bbar[3])
  );
  //AND U98
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U98 (
    .O(y[242]),
    .I0(a[15]),
    .I1(b[2])
  );
  //OR U98bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U98bar (
    .O(ybar[242]),
    .I0(abar[15]),
    .I1(bbar[2])
  );
  //AND U99
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U99 (
    .O(y[241]),
    .I0(a[15]),
    .I1(b[1])
  );
  //OR U99bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U99bar (
    .O(ybar[241]),
    .I0(abar[15]),
    .I1(bbar[1])
  );
  //AND U100
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U100 (
    .O(y[240]),
    .I0(a[15]),
    .I1(b[0])
  );
  //OR U100bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U100bar (
    .O(ybar[240]),
    .I0(abar[15]),
    .I1(bbar[0])
  );
  //AND U101
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U101 (
    .O(y[23]),
    .I0(a[1]),
    .I1(b[7])
  );
  //OR U101bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U101bar (
    .O(ybar[23]),
    .I0(abar[1]),
    .I1(bbar[7])
  );
  //AND U102
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U102 (
    .O(y[239]),
    .I0(a[14]),
    .I1(b[15])
  );
  //OR U102bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U102bar (
    .O(ybar[239]),
    .I0(abar[14]),
    .I1(bbar[15])
  );
  //AND U103
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U103 (
    .O(y[238]),
    .I0(a[14]),
    .I1(b[14])
  );
  //OR U103bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U103bar (
    .O(ybar[238]),
    .I0(abar[14]),
    .I1(bbar[14])
  );
  //AND U104
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U104 (
    .O(y[237]),
    .I0(a[14]),
    .I1(b[13])
  );
  //OR U104bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U104bar (
    .O(ybar[237]),
    .I0(abar[14]),
    .I1(bbar[13])
  );
  //AND U105
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U105 (
    .O(y[236]),
    .I0(a[14]),
    .I1(b[12])
  );
  //OR U105bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U105bar (
    .O(ybar[236]),
    .I0(abar[14]),
    .I1(bbar[12])
  );
  //AND U106
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U106 (
    .O(y[235]),
    .I0(a[14]),
    .I1(b[11])
  );
  //OR U106bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U106bar (
    .O(ybar[235]),
    .I0(abar[14]),
    .I1(bbar[11])
  );
  //AND U107
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U107 (
    .O(y[234]),
    .I0(a[14]),
    .I1(b[10])
  );
  //OR U107bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U107bar (
    .O(ybar[234]),
    .I0(abar[14]),
    .I1(bbar[10])
  );
  //AND U108
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U108 (
    .O(y[233]),
    .I0(a[14]),
    .I1(b[9])
  );
  //OR U108bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U108bar (
    .O(ybar[233]),
    .I0(abar[14]),
    .I1(bbar[9])
  );
  //AND U109
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U109 (
    .O(y[232]),
    .I0(a[14]),
    .I1(b[8])
  );
  //OR U109bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U109bar (
    .O(ybar[232]),
    .I0(abar[14]),
    .I1(bbar[8])
  );
  //AND U110
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U110 (
    .O(y[231]),
    .I0(a[14]),
    .I1(b[7])
  );
  //OR U110bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U110bar (
    .O(ybar[231]),
    .I0(abar[14]),
    .I1(bbar[7])
  );
  //AND U111
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U111 (
    .O(y[230]),
    .I0(a[14]),
    .I1(b[6])
  );
  //OR U111bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U111bar (
    .O(ybar[230]),
    .I0(abar[14]),
    .I1(bbar[6])
  );
  //AND U112
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U112 (
    .O(y[22]),
    .I0(a[1]),
    .I1(b[6])
  );
  //OR U112bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U112bar (
    .O(ybar[22]),
    .I0(abar[1]),
    .I1(bbar[6])
  );
  //AND U113
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U113 (
    .O(y[229]),
    .I0(a[14]),
    .I1(b[5])
  );
  //OR U113bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U113bar (
    .O(ybar[229]),
    .I0(abar[14]),
    .I1(bbar[5])
  );
  //AND U114
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U114 (
    .O(y[228]),
    .I0(a[14]),
    .I1(b[4])
  );
  //OR U114bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U114bar (
    .O(ybar[228]),
    .I0(abar[14]),
    .I1(bbar[4])
  );
  //AND U115
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U115 (
    .O(y[227]),
    .I0(a[14]),
    .I1(b[3])
  );
  //OR U115bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U115bar (
    .O(ybar[227]),
    .I0(abar[14]),
    .I1(bbar[3])
  );
  //AND U116
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U116 (
    .O(y[226]),
    .I0(a[14]),
    .I1(b[2])
  );
  //OR U116bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U116bar (
    .O(ybar[226]),
    .I0(abar[14]),
    .I1(bbar[2])
  );
  //AND U117
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U117 (
    .O(y[225]),
    .I0(a[14]),
    .I1(b[1])
  );
  //OR U117bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U117bar (
    .O(ybar[225]),
    .I0(abar[14]),
    .I1(bbar[1])
  );
  //AND U118
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U118 (
    .O(y[224]),
    .I0(a[14]),
    .I1(b[0])
  );
  //OR U118bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U118bar (
    .O(ybar[224]),
    .I0(abar[14]),
    .I1(bbar[0])
  );
  //AND U119
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U119 (
    .O(y[223]),
    .I0(a[13]),
    .I1(b[15])
  );
  //OR U119bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U119bar (
    .O(ybar[223]),
    .I0(abar[13]),
    .I1(bbar[15])
  );
  //AND U120
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U120 (
    .O(y[222]),
    .I0(a[13]),
    .I1(b[14])
  );
  //OR U120bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U120bar (
    .O(ybar[222]),
    .I0(abar[13]),
    .I1(bbar[14])
  );
  //AND U121
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U121 (
    .O(y[221]),
    .I0(a[13]),
    .I1(b[13])
  );
  //OR U121bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U121bar (
    .O(ybar[221]),
    .I0(abar[13]),
    .I1(bbar[13])
  );
  //AND U122
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U122 (
    .O(y[220]),
    .I0(a[13]),
    .I1(b[12])
  );
  //OR U122bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U122bar (
    .O(ybar[220]),
    .I0(abar[13]),
    .I1(bbar[12])
  );
  //AND U123
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U123 (
    .O(y[21]),
    .I0(a[1]),
    .I1(b[5])
  );
  //OR U123bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U123bar (
    .O(ybar[21]),
    .I0(abar[1]),
    .I1(bbar[5])
  );
  //AND U124
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U124 (
    .O(y[219]),
    .I0(a[13]),
    .I1(b[11])
  );
  //OR U124bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U124bar (
    .O(ybar[219]),
    .I0(abar[13]),
    .I1(bbar[11])
  );
  //AND U125
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U125 (
    .O(y[218]),
    .I0(a[13]),
    .I1(b[10])
  );
  //OR U125bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U125bar (
    .O(ybar[218]),
    .I0(abar[13]),
    .I1(bbar[10])
  );
  //AND U126
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U126 (
    .O(y[217]),
    .I0(a[13]),
    .I1(b[9])
  );
  //OR U126bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U126bar (
    .O(ybar[217]),
    .I0(abar[13]),
    .I1(bbar[9])
  );
  //AND U127
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U127 (
    .O(y[216]),
    .I0(a[13]),
    .I1(b[8])
  );
  //OR U127bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U127bar (
    .O(ybar[216]),
    .I0(abar[13]),
    .I1(bbar[8])
  );
  //AND U128
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U128 (
    .O(y[215]),
    .I0(a[13]),
    .I1(b[7])
  );
  //OR U128bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U128bar (
    .O(ybar[215]),
    .I0(abar[13]),
    .I1(bbar[7])
  );
  //AND U129
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U129 (
    .O(y[214]),
    .I0(a[13]),
    .I1(b[6])
  );
  //OR U129bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U129bar (
    .O(ybar[214]),
    .I0(abar[13]),
    .I1(bbar[6])
  );
  //AND U130
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U130 (
    .O(y[213]),
    .I0(a[13]),
    .I1(b[5])
  );
  //OR U130bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U130bar (
    .O(ybar[213]),
    .I0(abar[13]),
    .I1(bbar[5])
  );
  //AND U131
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U131 (
    .O(y[212]),
    .I0(a[13]),
    .I1(b[4])
  );
  //OR U131bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U131bar (
    .O(ybar[212]),
    .I0(abar[13]),
    .I1(bbar[4])
  );
  //AND U132
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U132 (
    .O(y[211]),
    .I0(a[13]),
    .I1(b[3])
  );
  //OR U132bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U132bar (
    .O(ybar[211]),
    .I0(abar[13]),
    .I1(bbar[3])
  );
  //AND U133
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U133 (
    .O(y[210]),
    .I0(a[13]),
    .I1(b[2])
  );
  //OR U133bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U133bar (
    .O(ybar[210]),
    .I0(abar[13]),
    .I1(bbar[2])
  );
  //AND U134
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U134 (
    .O(y[20]),
    .I0(a[1]),
    .I1(b[4])
  );
  //OR U134bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U134bar (
    .O(ybar[20]),
    .I0(abar[1]),
    .I1(bbar[4])
  );
  //AND U135
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U135 (
    .O(y[209]),
    .I0(a[13]),
    .I1(b[1])
  );
  //OR U135bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U135bar (
    .O(ybar[209]),
    .I0(abar[13]),
    .I1(bbar[1])
  );
  //AND U136
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U136 (
    .O(y[208]),
    .I0(a[13]),
    .I1(b[0])
  );
  //OR U136bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U136bar (
    .O(ybar[208]),
    .I0(abar[13]),
    .I1(bbar[0])
  );
  //AND U137
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U137 (
    .O(y[207]),
    .I0(a[12]),
    .I1(b[15])
  );
  //OR U137bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U137bar (
    .O(ybar[207]),
    .I0(abar[12]),
    .I1(bbar[15])
  );
  //AND U138
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U138 (
    .O(y[206]),
    .I0(a[12]),
    .I1(b[14])
  );
  //OR U138bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U138bar (
    .O(ybar[206]),
    .I0(abar[12]),
    .I1(bbar[14])
  );
  //AND U139
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U139 (
    .O(y[205]),
    .I0(a[12]),
    .I1(b[13])
  );
  //OR U139bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U139bar (
    .O(ybar[205]),
    .I0(abar[12]),
    .I1(bbar[13])
  );
  //AND U140
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U140 (
    .O(y[204]),
    .I0(a[12]),
    .I1(b[12])
  );
  //OR U140bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U140bar (
    .O(ybar[204]),
    .I0(abar[12]),
    .I1(bbar[12])
  );
  //AND U141
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U141 (
    .O(y[203]),
    .I0(a[12]),
    .I1(b[11])
  );
  //OR U141bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U141bar (
    .O(ybar[203]),
    .I0(abar[12]),
    .I1(bbar[11])
  );
  //AND U142
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U142 (
    .O(y[202]),
    .I0(a[12]),
    .I1(b[10])
  );
  //OR U142bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U142bar (
    .O(ybar[202]),
    .I0(abar[12]),
    .I1(bbar[10])
  );
  //AND U143
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U143 (
    .O(y[201]),
    .I0(a[12]),
    .I1(b[9])
  );
  //OR U143bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U143bar (
    .O(ybar[201]),
    .I0(abar[12]),
    .I1(bbar[9])
  );
  //AND U144
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U144 (
    .O(y[200]),
    .I0(a[12]),
    .I1(b[8])
  );
  //OR U144bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U144bar (
    .O(ybar[200]),
    .I0(abar[12]),
    .I1(bbar[8])
  );
  //AND U145
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U145 (
    .O(y[1]),
    .I0(b[1]),
    .I1(a[0])
  );
  //OR U145bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U145bar (
    .O(ybar[1]),
    .I0(bbar[1]),
    .I1(abar[0])
  );
  //AND U146
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U146 (
    .O(y[19]),
    .I0(a[1]),
    .I1(b[3])
  );
  //OR U146bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U146bar (
    .O(ybar[19]),
    .I0(abar[1]),
    .I1(bbar[3])
  );
  //AND U147
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U147 (
    .O(y[199]),
    .I0(a[12]),
    .I1(b[7])
  );
  //OR U147bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U147bar (
    .O(ybar[199]),
    .I0(abar[12]),
    .I1(bbar[7])
  );
  //AND U148
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U148 (
    .O(y[198]),
    .I0(a[12]),
    .I1(b[6])
  );
  //OR U148bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U148bar (
    .O(ybar[198]),
    .I0(abar[12]),
    .I1(bbar[6])
  );
  //AND U149
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U149 (
    .O(y[197]),
    .I0(a[12]),
    .I1(b[5])
  );
  //OR U149bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U149bar (
    .O(ybar[197]),
    .I0(abar[12]),
    .I1(bbar[5])
  );
  //AND U150
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U150 (
    .O(y[196]),
    .I0(a[12]),
    .I1(b[4])
  );
  //OR U150bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U150bar (
    .O(ybar[196]),
    .I0(abar[12]),
    .I1(bbar[4])
  );
  //AND U151
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U151 (
    .O(y[195]),
    .I0(a[12]),
    .I1(b[3])
  );
  //OR U151bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U151bar (
    .O(ybar[195]),
    .I0(abar[12]),
    .I1(bbar[3])
  );
  //AND U152
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U152 (
    .O(y[194]),
    .I0(a[12]),
    .I1(b[2])
  );
  //OR U152bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U152bar (
    .O(ybar[194]),
    .I0(abar[12]),
    .I1(bbar[2])
  );
  //AND U153
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U153 (
    .O(y[193]),
    .I0(a[12]),
    .I1(b[1])
  );
  //OR U153bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U153bar (
    .O(ybar[193]),
    .I0(abar[12]),
    .I1(bbar[1])
  );
  //AND U154
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U154 (
    .O(y[192]),
    .I0(a[12]),
    .I1(b[0])
  );
  //OR U154bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U154bar (
    .O(ybar[192]),
    .I0(abar[12]),
    .I1(bbar[0])
  );
  //AND U155
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U155 (
    .O(y[191]),
    .I0(a[11]),
    .I1(b[15])
  );
  //OR U155bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U155bar (
    .O(ybar[191]),
    .I0(abar[11]),
    .I1(bbar[15])
  );
  //AND U156
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U156 (
    .O(y[190]),
    .I0(a[11]),
    .I1(b[14])
  );
  //OR U156bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U156bar (
    .O(ybar[190]),
    .I0(abar[11]),
    .I1(bbar[14])
  );
  //AND U157
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U157 (
    .O(y[18]),
    .I0(a[1]),
    .I1(b[2])
  );
  //OR U157bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U157bar (
    .O(ybar[18]),
    .I0(abar[1]),
    .I1(bbar[2])
  );
  //AND U158
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U158 (
    .O(y[189]),
    .I0(a[11]),
    .I1(b[13])
  );
  //OR U158bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U158bar (
    .O(ybar[189]),
    .I0(abar[11]),
    .I1(bbar[13])
  );
  //AND U159
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U159 (
    .O(y[188]),
    .I0(a[11]),
    .I1(b[12])
  );
  //OR U159bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U159bar (
    .O(ybar[188]),
    .I0(abar[11]),
    .I1(bbar[12])
  );
  //AND U160
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U160 (
    .O(y[187]),
    .I0(a[11]),
    .I1(b[11])
  );
  //OR U160bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U160bar (
    .O(ybar[187]),
    .I0(abar[11]),
    .I1(bbar[11])
  );
  //AND U161
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U161 (
    .O(y[186]),
    .I0(a[11]),
    .I1(b[10])
  );
  //OR U161bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U161bar (
    .O(ybar[186]),
    .I0(abar[11]),
    .I1(bbar[10])
  );
  //AND U162
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U162 (
    .O(y[185]),
    .I0(a[11]),
    .I1(b[9])
  );
  //OR U162bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U162bar (
    .O(ybar[185]),
    .I0(abar[11]),
    .I1(bbar[9])
  );
  //AND U163
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U163 (
    .O(y[184]),
    .I0(a[11]),
    .I1(b[8])
  );
  //OR U163bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U163bar (
    .O(ybar[184]),
    .I0(abar[11]),
    .I1(bbar[8])
  );
  //AND U164
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U164 (
    .O(y[183]),
    .I0(a[11]),
    .I1(b[7])
  );
  //OR U164bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U164bar (
    .O(ybar[183]),
    .I0(abar[11]),
    .I1(bbar[7])
  );
  //AND U165
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U165 (
    .O(y[182]),
    .I0(a[11]),
    .I1(b[6])
  );
  //OR U165bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U165bar (
    .O(ybar[182]),
    .I0(abar[11]),
    .I1(bbar[6])
  );
  //AND U166
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U166 (
    .O(y[181]),
    .I0(a[11]),
    .I1(b[5])
  );
  //OR U166bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U166bar (
    .O(ybar[181]),
    .I0(abar[11]),
    .I1(bbar[5])
  );
  //AND U167
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U167 (
    .O(y[180]),
    .I0(a[11]),
    .I1(b[4])
  );
  //OR U167bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U167bar (
    .O(ybar[180]),
    .I0(abar[11]),
    .I1(bbar[4])
  );
  //AND U168
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U168 (
    .O(y[17]),
    .I0(a[1]),
    .I1(b[1])
  );
  //OR U168bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U168bar (
    .O(ybar[17]),
    .I0(abar[1]),
    .I1(bbar[1])
  );
  //AND U169
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U169 (
    .O(y[179]),
    .I0(a[11]),
    .I1(b[3])
  );
  //OR U169bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U169bar (
    .O(ybar[179]),
    .I0(abar[11]),
    .I1(bbar[3])
  );
  //AND U170
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U170 (
    .O(y[178]),
    .I0(a[11]),
    .I1(b[2])
  );
  //OR U170bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U170bar (
    .O(ybar[178]),
    .I0(abar[11]),
    .I1(bbar[2])
  );
  //AND U171
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U171 (
    .O(y[177]),
    .I0(a[11]),
    .I1(b[1])
  );
  //OR U171bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U171bar (
    .O(ybar[177]),
    .I0(abar[11]),
    .I1(bbar[1])
  );
  //AND U172
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U172 (
    .O(y[176]),
    .I0(a[11]),
    .I1(b[0])
  );
  //OR U172bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U172bar (
    .O(ybar[176]),
    .I0(abar[11]),
    .I1(bbar[0])
  );
  //AND U173
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U173 (
    .O(y[175]),
    .I0(a[10]),
    .I1(b[15])
  );
  //OR U173bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U173bar (
    .O(ybar[175]),
    .I0(abar[10]),
    .I1(bbar[15])
  );
  //AND U174
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U174 (
    .O(y[174]),
    .I0(a[10]),
    .I1(b[14])
  );
  //OR U174bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U174bar (
    .O(ybar[174]),
    .I0(abar[10]),
    .I1(bbar[14])
  );
  //AND U175
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U175 (
    .O(y[173]),
    .I0(a[10]),
    .I1(b[13])
  );
  //OR U175bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U175bar (
    .O(ybar[173]),
    .I0(abar[10]),
    .I1(bbar[13])
  );
  //AND U176
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U176 (
    .O(y[172]),
    .I0(a[10]),
    .I1(b[12])
  );
  //OR U176bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U176bar (
    .O(ybar[172]),
    .I0(abar[10]),
    .I1(bbar[12])
  );
  //AND U177
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U177 (
    .O(y[171]),
    .I0(a[10]),
    .I1(b[11])
  );
  //OR U177bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U177bar (
    .O(ybar[171]),
    .I0(abar[10]),
    .I1(bbar[11])
  );
  //AND U178
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U178 (
    .O(y[170]),
    .I0(a[10]),
    .I1(b[10])
  );
  //OR U178bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U178bar (
    .O(ybar[170]),
    .I0(abar[10]),
    .I1(bbar[10])
  );
  //AND U179
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U179 (
    .O(y[16]),
    .I0(a[1]),
    .I1(b[0])
  );
  //OR U179bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U179bar (
    .O(ybar[16]),
    .I0(abar[1]),
    .I1(bbar[0])
  );
  //AND U180
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U180 (
    .O(y[169]),
    .I0(a[10]),
    .I1(b[9])
  );
  //OR U180bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U180bar (
    .O(ybar[169]),
    .I0(abar[10]),
    .I1(bbar[9])
  );
  //AND U181
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U181 (
    .O(y[168]),
    .I0(a[10]),
    .I1(b[8])
  );
  //OR U181bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U181bar (
    .O(ybar[168]),
    .I0(abar[10]),
    .I1(bbar[8])
  );
  //AND U182
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U182 (
    .O(y[167]),
    .I0(a[10]),
    .I1(b[7])
  );
  //OR U182bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U182bar (
    .O(ybar[167]),
    .I0(abar[10]),
    .I1(bbar[7])
  );
  //AND U183
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U183 (
    .O(y[166]),
    .I0(a[10]),
    .I1(b[6])
  );
  //OR U183bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U183bar (
    .O(ybar[166]),
    .I0(abar[10]),
    .I1(bbar[6])
  );
  //AND U184
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U184 (
    .O(y[165]),
    .I0(a[10]),
    .I1(b[5])
  );
  //OR U184bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U184bar (
    .O(ybar[165]),
    .I0(abar[10]),
    .I1(bbar[5])
  );
  //AND U185
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U185 (
    .O(y[164]),
    .I0(a[10]),
    .I1(b[4])
  );
  //OR U185bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U185bar (
    .O(ybar[164]),
    .I0(abar[10]),
    .I1(bbar[4])
  );
  //AND U186
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U186 (
    .O(y[163]),
    .I0(a[10]),
    .I1(b[3])
  );
  //OR U186bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U186bar (
    .O(ybar[163]),
    .I0(abar[10]),
    .I1(bbar[3])
  );
  //AND U187
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U187 (
    .O(y[162]),
    .I0(a[10]),
    .I1(b[2])
  );
  //OR U187bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U187bar (
    .O(ybar[162]),
    .I0(abar[10]),
    .I1(bbar[2])
  );
  //AND U188
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U188 (
    .O(y[161]),
    .I0(a[10]),
    .I1(b[1])
  );
  //OR U188bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U188bar (
    .O(ybar[161]),
    .I0(abar[10]),
    .I1(bbar[1])
  );
  //AND U189
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U189 (
    .O(y[160]),
    .I0(a[10]),
    .I1(b[0])
  );
  //OR U189bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U189bar (
    .O(ybar[160]),
    .I0(abar[10]),
    .I1(bbar[0])
  );
  //AND U190
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U190 (
    .O(y[15]),
    .I0(b[15]),
    .I1(a[0])
  );
  //OR U190bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U190bar (
    .O(ybar[15]),
    .I0(bbar[15]),
    .I1(abar[0])
  );
  //AND U191
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U191 (
    .O(y[159]),
    .I0(a[9]),
    .I1(b[15])
  );
  //OR U191bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U191bar (
    .O(ybar[159]),
    .I0(abar[9]),
    .I1(bbar[15])
  );
  //AND U192
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U192 (
    .O(y[158]),
    .I0(a[9]),
    .I1(b[14])
  );
  //OR U192bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U192bar (
    .O(ybar[158]),
    .I0(abar[9]),
    .I1(bbar[14])
  );
  //AND U193
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U193 (
    .O(y[157]),
    .I0(a[9]),
    .I1(b[13])
  );
  //OR U193bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U193bar (
    .O(ybar[157]),
    .I0(abar[9]),
    .I1(bbar[13])
  );
  //AND U194
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U194 (
    .O(y[156]),
    .I0(a[9]),
    .I1(b[12])
  );
  //OR U194bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U194bar (
    .O(ybar[156]),
    .I0(abar[9]),
    .I1(bbar[12])
  );
  //AND U195
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U195 (
    .O(y[155]),
    .I0(a[9]),
    .I1(b[11])
  );
  //OR U195bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U195bar (
    .O(ybar[155]),
    .I0(abar[9]),
    .I1(bbar[11])
  );
  //AND U196
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U196 (
    .O(y[154]),
    .I0(a[9]),
    .I1(b[10])
  );
  //OR U196bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U196bar (
    .O(ybar[154]),
    .I0(abar[9]),
    .I1(bbar[10])
  );
  //AND U197
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U197 (
    .O(y[153]),
    .I0(a[9]),
    .I1(b[9])
  );
  //OR U197bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U197bar (
    .O(ybar[153]),
    .I0(abar[9]),
    .I1(bbar[9])
  );
  //AND U198
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U198 (
    .O(y[152]),
    .I0(a[9]),
    .I1(b[8])
  );
  //OR U198bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U198bar (
    .O(ybar[152]),
    .I0(abar[9]),
    .I1(bbar[8])
  );
  //AND U199
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U199 (
    .O(y[151]),
    .I0(a[9]),
    .I1(b[7])
  );
  //OR U199bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U199bar (
    .O(ybar[151]),
    .I0(abar[9]),
    .I1(bbar[7])
  );
  //AND U200
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U200 (
    .O(y[150]),
    .I0(a[9]),
    .I1(b[6])
  );
  //OR U200bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U200bar (
    .O(ybar[150]),
    .I0(abar[9]),
    .I1(bbar[6])
  );
  //AND U201
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U201 (
    .O(y[14]),
    .I0(b[14]),
    .I1(a[0])
  );
  //OR U201bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U201bar (
    .O(ybar[14]),
    .I0(bbar[14]),
    .I1(abar[0])
  );
  //AND U202
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U202 (
    .O(y[149]),
    .I0(a[9]),
    .I1(b[5])
  );
  //OR U202bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U202bar (
    .O(ybar[149]),
    .I0(abar[9]),
    .I1(bbar[5])
  );
  //AND U203
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U203 (
    .O(y[148]),
    .I0(a[9]),
    .I1(b[4])
  );
  //OR U203bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U203bar (
    .O(ybar[148]),
    .I0(abar[9]),
    .I1(bbar[4])
  );
  //AND U204
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U204 (
    .O(y[147]),
    .I0(a[9]),
    .I1(b[3])
  );
  //OR U204bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U204bar (
    .O(ybar[147]),
    .I0(abar[9]),
    .I1(bbar[3])
  );
  //AND U205
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U205 (
    .O(y[146]),
    .I0(a[9]),
    .I1(b[2])
  );
  //OR U205bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U205bar (
    .O(ybar[146]),
    .I0(abar[9]),
    .I1(bbar[2])
  );
  //AND U206
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U206 (
    .O(y[145]),
    .I0(a[9]),
    .I1(b[1])
  );
  //OR U206bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U206bar (
    .O(ybar[145]),
    .I0(abar[9]),
    .I1(bbar[1])
  );
  //AND U207
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U207 (
    .O(y[144]),
    .I0(a[9]),
    .I1(b[0])
  );
  //OR U207bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U207bar (
    .O(ybar[144]),
    .I0(abar[9]),
    .I1(bbar[0])
  );
  //AND U208
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U208 (
    .O(y[143]),
    .I0(a[8]),
    .I1(b[15])
  );
  //OR U208bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U208bar (
    .O(ybar[143]),
    .I0(abar[8]),
    .I1(bbar[15])
  );
  //AND U209
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U209 (
    .O(y[142]),
    .I0(a[8]),
    .I1(b[14])
  );
  //OR U209bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U209bar (
    .O(ybar[142]),
    .I0(abar[8]),
    .I1(bbar[14])
  );
  //AND U210
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U210 (
    .O(y[141]),
    .I0(a[8]),
    .I1(b[13])
  );
  //OR U210bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U210bar (
    .O(ybar[141]),
    .I0(abar[8]),
    .I1(bbar[13])
  );
  //AND U211
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U211 (
    .O(y[140]),
    .I0(a[8]),
    .I1(b[12])
  );
  //OR U211bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U211bar (
    .O(ybar[140]),
    .I0(abar[8]),
    .I1(bbar[12])
  );
  //AND U212
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U212 (
    .O(y[13]),
    .I0(b[13]),
    .I1(a[0])
  );
  //OR U212bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U212bar (
    .O(ybar[13]),
    .I0(bbar[13]),
    .I1(abar[0])
  );
  //AND U213
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U213 (
    .O(y[139]),
    .I0(a[8]),
    .I1(b[11])
  );
  //OR U213bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U213bar (
    .O(ybar[139]),
    .I0(abar[8]),
    .I1(bbar[11])
  );
  //AND U214
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U214 (
    .O(y[138]),
    .I0(a[8]),
    .I1(b[10])
  );
  //OR U214bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U214bar (
    .O(ybar[138]),
    .I0(abar[8]),
    .I1(bbar[10])
  );
  //AND U215
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U215 (
    .O(y[137]),
    .I0(a[8]),
    .I1(b[9])
  );
  //OR U215bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U215bar (
    .O(ybar[137]),
    .I0(abar[8]),
    .I1(bbar[9])
  );
  //AND U216
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U216 (
    .O(y[136]),
    .I0(a[8]),
    .I1(b[8])
  );
  //OR U216bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U216bar (
    .O(ybar[136]),
    .I0(abar[8]),
    .I1(bbar[8])
  );
  //AND U217
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U217 (
    .O(y[135]),
    .I0(a[8]),
    .I1(b[7])
  );
  //OR U217bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U217bar (
    .O(ybar[135]),
    .I0(abar[8]),
    .I1(bbar[7])
  );
  //AND U218
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U218 (
    .O(y[134]),
    .I0(a[8]),
    .I1(b[6])
  );
  //OR U218bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U218bar (
    .O(ybar[134]),
    .I0(abar[8]),
    .I1(bbar[6])
  );
  //AND U219
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U219 (
    .O(y[133]),
    .I0(a[8]),
    .I1(b[5])
  );
  //OR U219bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U219bar (
    .O(ybar[133]),
    .I0(abar[8]),
    .I1(bbar[5])
  );
  //AND U220
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U220 (
    .O(y[132]),
    .I0(a[8]),
    .I1(b[4])
  );
  //OR U220bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U220bar (
    .O(ybar[132]),
    .I0(abar[8]),
    .I1(bbar[4])
  );
  //AND U221
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U221 (
    .O(y[131]),
    .I0(a[8]),
    .I1(b[3])
  );
  //OR U221bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U221bar (
    .O(ybar[131]),
    .I0(abar[8]),
    .I1(bbar[3])
  );
  //AND U222
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U222 (
    .O(y[130]),
    .I0(a[8]),
    .I1(b[2])
  );
  //OR U222bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U222bar (
    .O(ybar[130]),
    .I0(abar[8]),
    .I1(bbar[2])
  );
  //AND U223
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U223 (
    .O(y[12]),
    .I0(b[12]),
    .I1(a[0])
  );
  //OR U223bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U223bar (
    .O(ybar[12]),
    .I0(bbar[12]),
    .I1(abar[0])
  );
  //AND U224
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U224 (
    .O(y[129]),
    .I0(a[8]),
    .I1(b[1])
  );
  //OR U224bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U224bar (
    .O(ybar[129]),
    .I0(abar[8]),
    .I1(bbar[1])
  );
  //AND U225
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U225 (
    .O(y[128]),
    .I0(a[8]),
    .I1(b[0])
  );
  //OR U225bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U225bar (
    .O(ybar[128]),
    .I0(abar[8]),
    .I1(bbar[0])
  );
  //AND U226
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U226 (
    .O(y[127]),
    .I0(a[7]),
    .I1(b[15])
  );
  //OR U226bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U226bar (
    .O(ybar[127]),
    .I0(abar[7]),
    .I1(bbar[15])
  );
  //AND U227
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U227 (
    .O(y[126]),
    .I0(a[7]),
    .I1(b[14])
  );
  //OR U227bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U227bar (
    .O(ybar[126]),
    .I0(abar[7]),
    .I1(bbar[14])
  );
  //AND U228
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U228 (
    .O(y[125]),
    .I0(a[7]),
    .I1(b[13])
  );
  //OR U228bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U228bar (
    .O(ybar[125]),
    .I0(abar[7]),
    .I1(bbar[13])
  );
  //AND U229
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U229 (
    .O(y[124]),
    .I0(a[7]),
    .I1(b[12])
  );
  //OR U229bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U229bar (
    .O(ybar[124]),
    .I0(abar[7]),
    .I1(bbar[12])
  );
  //AND U230
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U230 (
    .O(y[123]),
    .I0(a[7]),
    .I1(b[11])
  );
  //OR U230bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U230bar (
    .O(ybar[123]),
    .I0(abar[7]),
    .I1(bbar[11])
  );
  //AND U231
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U231 (
    .O(y[122]),
    .I0(a[7]),
    .I1(b[10])
  );
  //OR U231bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U231bar (
    .O(ybar[122]),
    .I0(abar[7]),
    .I1(bbar[10])
  );
  //AND U232
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U232 (
    .O(y[121]),
    .I0(a[7]),
    .I1(b[9])
  );
  //OR U232bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U232bar (
    .O(ybar[121]),
    .I0(abar[7]),
    .I1(bbar[9])
  );
  //AND U233
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U233 (
    .O(y[120]),
    .I0(a[7]),
    .I1(b[8])
  );
  //OR U233bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U233bar (
    .O(ybar[120]),
    .I0(abar[7]),
    .I1(bbar[8])
  );
  //AND U234
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U234 (
    .O(y[11]),
    .I0(b[11]),
    .I1(a[0])
  );
  //OR U234bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U234bar (
    .O(ybar[11]),
    .I0(bbar[11]),
    .I1(abar[0])
  );
  //AND U235
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U235 (
    .O(y[119]),
    .I0(a[7]),
    .I1(b[7])
  );
  //OR U235bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U235bar (
    .O(ybar[119]),
    .I0(abar[7]),
    .I1(bbar[7])
  );
  //AND U236
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U236 (
    .O(y[118]),
    .I0(a[7]),
    .I1(b[6])
  );
  //OR U236bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U236bar (
    .O(ybar[118]),
    .I0(abar[7]),
    .I1(bbar[6])
  );
  //AND U237
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U237 (
    .O(y[117]),
    .I0(a[7]),
    .I1(b[5])
  );
  //OR U237bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U237bar (
    .O(ybar[117]),
    .I0(abar[7]),
    .I1(bbar[5])
  );
  //AND U238
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U238 (
    .O(y[116]),
    .I0(a[7]),
    .I1(b[4])
  );
  //OR U238bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U238bar (
    .O(ybar[116]),
    .I0(abar[7]),
    .I1(bbar[4])
  );
  //AND U239
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U239 (
    .O(y[115]),
    .I0(a[7]),
    .I1(b[3])
  );
  //OR U239bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U239bar (
    .O(ybar[115]),
    .I0(abar[7]),
    .I1(bbar[3])
  );
  //AND U240
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U240 (
    .O(y[114]),
    .I0(a[7]),
    .I1(b[2])
  );
  //OR U240bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U240bar (
    .O(ybar[114]),
    .I0(abar[7]),
    .I1(bbar[2])
  );
  //AND U241
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U241 (
    .O(y[113]),
    .I0(a[7]),
    .I1(b[1])
  );
  //OR U241bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U241bar (
    .O(ybar[113]),
    .I0(abar[7]),
    .I1(bbar[1])
  );
  //AND U242
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U242 (
    .O(y[112]),
    .I0(a[7]),
    .I1(b[0])
  );
  //OR U242bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U242bar (
    .O(ybar[112]),
    .I0(abar[7]),
    .I1(bbar[0])
  );
  //AND U243
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U243 (
    .O(y[111]),
    .I0(b[15]),
    .I1(a[6])
  );
  //OR U243bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U243bar (
    .O(ybar[111]),
    .I0(bbar[15]),
    .I1(abar[6])
  );
  //AND U244
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U244 (
    .O(y[110]),
    .I0(b[14]),
    .I1(a[6])
  );
  //OR U244bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U244bar (
    .O(ybar[110]),
    .I0(bbar[14]),
    .I1(abar[6])
  );
  //AND U245
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U245 (
    .O(y[10]),
    .I0(b[10]),
    .I1(a[0])
  );
  //OR U245bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U245bar (
    .O(ybar[10]),
    .I0(bbar[10]),
    .I1(abar[0])
  );
  //AND U246
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U246 (
    .O(y[109]),
    .I0(b[13]),
    .I1(a[6])
  );
  //OR U246bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U246bar (
    .O(ybar[109]),
    .I0(bbar[13]),
    .I1(abar[6])
  );
  //AND U247
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U247 (
    .O(y[108]),
    .I0(b[12]),
    .I1(a[6])
  );
  //OR U247bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U247bar (
    .O(ybar[108]),
    .I0(bbar[12]),
    .I1(abar[6])
  );
  //AND U248
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U248 (
    .O(y[107]),
    .I0(b[11]),
    .I1(a[6])
  );
  //OR U248bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U248bar (
    .O(ybar[107]),
    .I0(bbar[11]),
    .I1(abar[6])
  );
  //AND U249
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U249 (
    .O(y[106]),
    .I0(b[10]),
    .I1(a[6])
  );
  //OR U249bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U249bar (
    .O(ybar[106]),
    .I0(bbar[10]),
    .I1(abar[6])
  );
  //AND U250
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U250 (
    .O(y[105]),
    .I0(a[6]),
    .I1(b[9])
  );
  //OR U250bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U250bar (
    .O(ybar[105]),
    .I0(abar[6]),
    .I1(bbar[9])
  );
  //AND U251
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U251 (
    .O(y[104]),
    .I0(b[8]),
    .I1(a[6])
  );
  //OR U251bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U251bar (
    .O(ybar[104]),
    .I0(bbar[8]),
    .I1(abar[6])
  );
  //AND U252
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U252 (
    .O(y[103]),
    .I0(b[7]),
    .I1(a[6])
  );
  //OR U252bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U252bar (
    .O(ybar[103]),
    .I0(bbar[7]),
    .I1(abar[6])
  );
  //AND U253
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U253 (
    .O(y[102]),
    .I0(b[6]),
    .I1(a[6])
  );
  //OR U253bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U253bar (
    .O(ybar[102]),
    .I0(bbar[6]),
    .I1(abar[6])
  );
  //AND U254
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U254 (
    .O(y[101]),
    .I0(b[5]),
    .I1(a[6])
  );
  //OR U254bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U254bar (
    .O(ybar[101]),
    .I0(bbar[5]),
    .I1(abar[6])
  );
  //AND U255
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U255 (
    .O(y[100]),
    .I0(b[4]),
    .I1(a[6])
  );
  //OR U255bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U255bar (
    .O(ybar[100]),
    .I0(bbar[4]),
    .I1(abar[6])
  );
  //AND U256
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U256 (
    .O(y[0]),
    .I0(b[0]),
    .I1(a[0])
  );
  //OR U256bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U256bar (
    .O(ybar[0]),
    .I0(bbar[0]),
    .I1(abar[0])
  );
endmodule

module decode_14 ( in, out );

  input wire [7:0] in;
//input_done

  output wire [255:0] out;
//output_done

  wire [15:0] level1;
  wire [31:0] level2;
//wire_done

  CD2_56 cd_l1_1 ( .a(in[1]), .b(in[0]), .y(level1[3:0]) );
  CD2_55 cd_l1_2 ( .a(in[3]), .b(in[2]), .y(level1[7:4]) );
  CD2_54 cd_l1_3 ( .a(in[5]), .b(in[4]), .y(level1[11:8]) );
  CD2_53 cd_l1_4 ( .a(in[7]), .b(in[6]), .y(level1[15:12]) );
  CD4_28 cd_l2_1 ( .a(level1[7:4]), .b(level1[3:0]), .y(level2[15:0]) );
  CD4_27 cd_l2_2 ( .a(level1[15:12]), .b(level1[11:8]), .y(level2[31:16]) );
  CD16_14 cd_l3 ( .a(level2[31:16]), .b(level2[15:0]), .y(out) );
endmodule

module encode_14 ( in, out );

  input wire [255:0] in;
  wire [255:0] inbar;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
  assign inbar[8] = ~in[8];
  assign inbar[9] = ~in[9];
  assign inbar[10] = ~in[10];
  assign inbar[11] = ~in[11];
  assign inbar[12] = ~in[12];
  assign inbar[13] = ~in[13];
  assign inbar[14] = ~in[14];
  assign inbar[15] = ~in[15];
  assign inbar[16] = ~in[16];
  assign inbar[17] = ~in[17];
  assign inbar[18] = ~in[18];
  assign inbar[19] = ~in[19];
  assign inbar[20] = ~in[20];
  assign inbar[21] = ~in[21];
  assign inbar[22] = ~in[22];
  assign inbar[23] = ~in[23];
  assign inbar[24] = ~in[24];
  assign inbar[25] = ~in[25];
  assign inbar[26] = ~in[26];
  assign inbar[27] = ~in[27];
  assign inbar[28] = ~in[28];
  assign inbar[29] = ~in[29];
  assign inbar[30] = ~in[30];
  assign inbar[31] = ~in[31];
  assign inbar[32] = ~in[32];
  assign inbar[33] = ~in[33];
  assign inbar[34] = ~in[34];
  assign inbar[35] = ~in[35];
  assign inbar[36] = ~in[36];
  assign inbar[37] = ~in[37];
  assign inbar[38] = ~in[38];
  assign inbar[39] = ~in[39];
  assign inbar[40] = ~in[40];
  assign inbar[41] = ~in[41];
  assign inbar[42] = ~in[42];
  assign inbar[43] = ~in[43];
  assign inbar[44] = ~in[44];
  assign inbar[45] = ~in[45];
  assign inbar[46] = ~in[46];
  assign inbar[47] = ~in[47];
  assign inbar[48] = ~in[48];
  assign inbar[49] = ~in[49];
  assign inbar[50] = ~in[50];
  assign inbar[51] = ~in[51];
  assign inbar[52] = ~in[52];
  assign inbar[53] = ~in[53];
  assign inbar[54] = ~in[54];
  assign inbar[55] = ~in[55];
  assign inbar[56] = ~in[56];
  assign inbar[57] = ~in[57];
  assign inbar[58] = ~in[58];
  assign inbar[59] = ~in[59];
  assign inbar[60] = ~in[60];
  assign inbar[61] = ~in[61];
  assign inbar[62] = ~in[62];
  assign inbar[63] = ~in[63];
  assign inbar[64] = ~in[64];
  assign inbar[65] = ~in[65];
  assign inbar[66] = ~in[66];
  assign inbar[67] = ~in[67];
  assign inbar[68] = ~in[68];
  assign inbar[69] = ~in[69];
  assign inbar[70] = ~in[70];
  assign inbar[71] = ~in[71];
  assign inbar[72] = ~in[72];
  assign inbar[73] = ~in[73];
  assign inbar[74] = ~in[74];
  assign inbar[75] = ~in[75];
  assign inbar[76] = ~in[76];
  assign inbar[77] = ~in[77];
  assign inbar[78] = ~in[78];
  assign inbar[79] = ~in[79];
  assign inbar[80] = ~in[80];
  assign inbar[81] = ~in[81];
  assign inbar[82] = ~in[82];
  assign inbar[83] = ~in[83];
  assign inbar[84] = ~in[84];
  assign inbar[85] = ~in[85];
  assign inbar[86] = ~in[86];
  assign inbar[87] = ~in[87];
  assign inbar[88] = ~in[88];
  assign inbar[89] = ~in[89];
  assign inbar[90] = ~in[90];
  assign inbar[91] = ~in[91];
  assign inbar[92] = ~in[92];
  assign inbar[93] = ~in[93];
  assign inbar[94] = ~in[94];
  assign inbar[95] = ~in[95];
  assign inbar[96] = ~in[96];
  assign inbar[97] = ~in[97];
  assign inbar[98] = ~in[98];
  assign inbar[99] = ~in[99];
  assign inbar[100] = ~in[100];
  assign inbar[101] = ~in[101];
  assign inbar[102] = ~in[102];
  assign inbar[103] = ~in[103];
  assign inbar[104] = ~in[104];
  assign inbar[105] = ~in[105];
  assign inbar[106] = ~in[106];
  assign inbar[107] = ~in[107];
  assign inbar[108] = ~in[108];
  assign inbar[109] = ~in[109];
  assign inbar[110] = ~in[110];
  assign inbar[111] = ~in[111];
  assign inbar[112] = ~in[112];
  assign inbar[113] = ~in[113];
  assign inbar[114] = ~in[114];
  assign inbar[115] = ~in[115];
  assign inbar[116] = ~in[116];
  assign inbar[117] = ~in[117];
  assign inbar[118] = ~in[118];
  assign inbar[119] = ~in[119];
  assign inbar[120] = ~in[120];
  assign inbar[121] = ~in[121];
  assign inbar[122] = ~in[122];
  assign inbar[123] = ~in[123];
  assign inbar[124] = ~in[124];
  assign inbar[125] = ~in[125];
  assign inbar[126] = ~in[126];
  assign inbar[127] = ~in[127];
  assign inbar[128] = ~in[128];
  assign inbar[129] = ~in[129];
  assign inbar[130] = ~in[130];
  assign inbar[131] = ~in[131];
  assign inbar[132] = ~in[132];
  assign inbar[133] = ~in[133];
  assign inbar[134] = ~in[134];
  assign inbar[135] = ~in[135];
  assign inbar[136] = ~in[136];
  assign inbar[137] = ~in[137];
  assign inbar[138] = ~in[138];
  assign inbar[139] = ~in[139];
  assign inbar[140] = ~in[140];
  assign inbar[141] = ~in[141];
  assign inbar[142] = ~in[142];
  assign inbar[143] = ~in[143];
  assign inbar[144] = ~in[144];
  assign inbar[145] = ~in[145];
  assign inbar[146] = ~in[146];
  assign inbar[147] = ~in[147];
  assign inbar[148] = ~in[148];
  assign inbar[149] = ~in[149];
  assign inbar[150] = ~in[150];
  assign inbar[151] = ~in[151];
  assign inbar[152] = ~in[152];
  assign inbar[153] = ~in[153];
  assign inbar[154] = ~in[154];
  assign inbar[155] = ~in[155];
  assign inbar[156] = ~in[156];
  assign inbar[157] = ~in[157];
  assign inbar[158] = ~in[158];
  assign inbar[159] = ~in[159];
  assign inbar[160] = ~in[160];
  assign inbar[161] = ~in[161];
  assign inbar[162] = ~in[162];
  assign inbar[163] = ~in[163];
  assign inbar[164] = ~in[164];
  assign inbar[165] = ~in[165];
  assign inbar[166] = ~in[166];
  assign inbar[167] = ~in[167];
  assign inbar[168] = ~in[168];
  assign inbar[169] = ~in[169];
  assign inbar[170] = ~in[170];
  assign inbar[171] = ~in[171];
  assign inbar[172] = ~in[172];
  assign inbar[173] = ~in[173];
  assign inbar[174] = ~in[174];
  assign inbar[175] = ~in[175];
  assign inbar[176] = ~in[176];
  assign inbar[177] = ~in[177];
  assign inbar[178] = ~in[178];
  assign inbar[179] = ~in[179];
  assign inbar[180] = ~in[180];
  assign inbar[181] = ~in[181];
  assign inbar[182] = ~in[182];
  assign inbar[183] = ~in[183];
  assign inbar[184] = ~in[184];
  assign inbar[185] = ~in[185];
  assign inbar[186] = ~in[186];
  assign inbar[187] = ~in[187];
  assign inbar[188] = ~in[188];
  assign inbar[189] = ~in[189];
  assign inbar[190] = ~in[190];
  assign inbar[191] = ~in[191];
  assign inbar[192] = ~in[192];
  assign inbar[193] = ~in[193];
  assign inbar[194] = ~in[194];
  assign inbar[195] = ~in[195];
  assign inbar[196] = ~in[196];
  assign inbar[197] = ~in[197];
  assign inbar[198] = ~in[198];
  assign inbar[199] = ~in[199];
  assign inbar[200] = ~in[200];
  assign inbar[201] = ~in[201];
  assign inbar[202] = ~in[202];
  assign inbar[203] = ~in[203];
  assign inbar[204] = ~in[204];
  assign inbar[205] = ~in[205];
  assign inbar[206] = ~in[206];
  assign inbar[207] = ~in[207];
  assign inbar[208] = ~in[208];
  assign inbar[209] = ~in[209];
  assign inbar[210] = ~in[210];
  assign inbar[211] = ~in[211];
  assign inbar[212] = ~in[212];
  assign inbar[213] = ~in[213];
  assign inbar[214] = ~in[214];
  assign inbar[215] = ~in[215];
  assign inbar[216] = ~in[216];
  assign inbar[217] = ~in[217];
  assign inbar[218] = ~in[218];
  assign inbar[219] = ~in[219];
  assign inbar[220] = ~in[220];
  assign inbar[221] = ~in[221];
  assign inbar[222] = ~in[222];
  assign inbar[223] = ~in[223];
  assign inbar[224] = ~in[224];
  assign inbar[225] = ~in[225];
  assign inbar[226] = ~in[226];
  assign inbar[227] = ~in[227];
  assign inbar[228] = ~in[228];
  assign inbar[229] = ~in[229];
  assign inbar[230] = ~in[230];
  assign inbar[231] = ~in[231];
  assign inbar[232] = ~in[232];
  assign inbar[233] = ~in[233];
  assign inbar[234] = ~in[234];
  assign inbar[235] = ~in[235];
  assign inbar[236] = ~in[236];
  assign inbar[237] = ~in[237];
  assign inbar[238] = ~in[238];
  assign inbar[239] = ~in[239];
  assign inbar[240] = ~in[240];
  assign inbar[241] = ~in[241];
  assign inbar[242] = ~in[242];
  assign inbar[243] = ~in[243];
  assign inbar[244] = ~in[244];
  assign inbar[245] = ~in[245];
  assign inbar[246] = ~in[246];
  assign inbar[247] = ~in[247];
  assign inbar[248] = ~in[248];
  assign inbar[249] = ~in[249];
  assign inbar[250] = ~in[250];
  assign inbar[251] = ~in[251];
  assign inbar[252] = ~in[252];
  assign inbar[253] = ~in[253];
  assign inbar[254] = ~in[254];
  assign inbar[255] = ~in[255];
//input_done

  output wire [7:0] out;
  wire [7:0] outbar;
//output_done

  wire in_81;
  wire in_80;
  wire in_79;
  wire in_78;
  wire in_77;
  wire in_76;
  wire in_75;
  wire in_74;
  wire in_73;
  wire in_72;
  wire in_71;
  wire in_70;
  wire in_69;
  wire in_68;
  wire in_67;
  wire in_66;
  wire in_65;
  wire in_64;
  wire in_63;
  wire in_62;
  wire in_61;
  wire in_60;
  wire in_59;
  wire in_58;
  wire in_57;
  wire in_56;
  wire in_55;
  wire in_54;
  wire in_53;
  wire in_52;
  wire in_51;
  wire in_50;
  wire in_49;
  wire in_48;
  wire in_47;
  wire in_46;
  wire in_45;
  wire in_44;
  wire in_43;
  wire in_42;
  wire in_41;
  wire in_40;
  wire in_39;
  wire in_38;
  wire in_37;
  wire in_36;
  wire in_35;
  wire in_34;
  wire in_33;
  wire in_32;
  wire in_31;
  wire in_30;
  wire in_29;
  wire in_28;
  wire in_27;
  wire in_26;
  wire in_25;
  wire in_24;
  wire in_23;
  wire in_22;
  wire in_21;
  wire in_20;
  wire in_19;
  wire in_18;
  wire in_17;
  wire in_16;
  wire in_15;
  wire in_14;
  wire in_13;
  wire in_12;
  wire in_11;
  wire in_10;
  wire in_9;
  wire in_8;
  wire in_7;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_3;
  wire in_2;
  wire in_1;
  wire in_0;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire in_81bar;
  wire in_80bar;
  wire in_79bar;
  wire in_78bar;
  wire in_77bar;
  wire in_76bar;
  wire in_75bar;
  wire in_74bar;
  wire in_73bar;
  wire in_72bar;
  wire in_71bar;
  wire in_70bar;
  wire in_69bar;
  wire in_68bar;
  wire in_67bar;
  wire in_66bar;
  wire in_65bar;
  wire in_64bar;
  wire in_63bar;
  wire in_62bar;
  wire in_61bar;
  wire in_60bar;
  wire in_59bar;
  wire in_58bar;
  wire in_57bar;
  wire in_56bar;
  wire in_55bar;
  wire in_54bar;
  wire in_53bar;
  wire in_52bar;
  wire in_51bar;
  wire in_50bar;
  wire in_49bar;
  wire in_48bar;
  wire in_47bar;
  wire in_46bar;
  wire in_45bar;
  wire in_44bar;
  wire in_43bar;
  wire in_42bar;
  wire in_41bar;
  wire in_40bar;
  wire in_39bar;
  wire in_38bar;
  wire in_37bar;
  wire in_36bar;
  wire in_35bar;
  wire in_34bar;
  wire in_33bar;
  wire in_32bar;
  wire in_31bar;
  wire in_30bar;
  wire in_29bar;
  wire in_28bar;
  wire in_27bar;
  wire in_26bar;
  wire in_25bar;
  wire in_24bar;
  wire in_23bar;
  wire in_22bar;
  wire in_21bar;
  wire in_20bar;
  wire in_19bar;
  wire in_18bar;
  wire in_17bar;
  wire in_16bar;
  wire in_15bar;
  wire in_14bar;
  wire in_13bar;
  wire in_12bar;
  wire in_11bar;
  wire in_10bar;
  wire in_9bar;
  wire in_8bar;
  wire in_7bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_3bar;
  wire in_2bar;
  wire in_1bar;
  wire in_0bar;
  wire n487bar;
  wire n488bar;
  wire n489bar;
  wire n490bar;
  wire n491bar;
  wire n492bar;
  wire n493bar;
  wire n494bar;
  wire n495bar;
  wire n496bar;
  wire n497bar;
  wire n498bar;
  wire n499bar;
  wire n500bar;
  wire n501bar;
  wire n502bar;
  wire n503bar;
  wire n504bar;
  wire n505bar;
  wire n506bar;
  wire n507bar;
  wire n508bar;
  wire n509bar;
  wire n510bar;
  wire n511bar;
  wire n512bar;
  wire n513bar;
  wire n514bar;
  wire n515bar;
  wire n516bar;
  wire n517bar;
  wire n518bar;
  wire n519bar;
  wire n520bar;
  wire n521bar;
  wire n522bar;
  wire n523bar;
  wire n524bar;
  wire n525bar;
  wire n526bar;
  wire n527bar;
  wire n528bar;
  wire n529bar;
  wire n530bar;
  wire n531bar;
  wire n532bar;
  wire n533bar;
  wire n534bar;
  wire n535bar;
  wire n536bar;
  wire n537bar;
  wire n538bar;
  wire n539bar;
  wire n540bar;
  wire n541bar;
  wire n542bar;
  wire n543bar;
  wire n544bar;
  wire n545bar;
  wire n546bar;
  wire n547bar;
  wire n548bar;
  wire n549bar;
  wire n550bar;
  wire n551bar;
  wire n552bar;
  wire n553bar;
  wire n554bar;
  wire n555bar;
  wire n556bar;
  wire n557bar;
  wire n558bar;
  wire n559bar;
  wire n560bar;
  wire n561bar;
  wire n562bar;
  wire n563bar;
  wire n564bar;
  wire n565bar;
  wire n566bar;
  wire n567bar;
  wire n568bar;
  wire n569bar;
  wire n570bar;
  wire n571bar;
  wire n572bar;
  wire n573bar;
  wire n574bar;
  wire n575bar;
  wire n576bar;
  wire n577bar;
  wire n578bar;
  wire n579bar;
  wire n580bar;
  wire n581bar;
  wire n582bar;
  wire n583bar;
  wire n584bar;
  wire n585bar;
  wire n586bar;
  wire n587bar;
  wire n588bar;
  wire n589bar;
  wire n590bar;
  wire n591bar;
  wire n592bar;
  wire n593bar;
  wire n594bar;
  wire n595bar;
  wire n596bar;
  wire n597bar;
  wire n598bar;
  wire n599bar;
  wire n600bar;
  wire n601bar;
  wire n602bar;
  wire n603bar;
  wire n604bar;
  wire n605bar;
  wire n606bar;
  wire n607bar;
  wire n608bar;
  wire n609bar;
  wire n610bar;
  wire n611bar;
  wire n612bar;
  wire n613bar;
  wire n614bar;
  wire n615bar;
  wire n616bar;
  wire n617bar;
  wire n618bar;
  wire n619bar;
  wire n620bar;
  wire n621bar;
  wire n622bar;
  wire n623bar;
  wire n624bar;
  wire n625bar;
  wire n626bar;
  wire n627bar;
  wire n628bar;
  wire n629bar;
  wire n630bar;
  wire n631bar;
  wire n632bar;
  wire n633bar;
  wire n634bar;
  wire n635bar;
  wire n636bar;
  wire n637bar;
  wire n638bar;
  wire n639bar;
  wire n640bar;
  wire n641bar;
  wire n642bar;
  wire n643bar;
  wire n644bar;
  wire n645bar;
  wire n646bar;
  wire n647bar;
  wire n648bar;
  wire n649bar;
  wire n650bar;
  wire n651bar;
  wire n652bar;
  wire n653bar;
  wire n654bar;
  wire n655bar;
  wire n656bar;
  wire n657bar;
  wire n658bar;
  wire n659bar;
  wire n660bar;
  wire n661bar;
  wire n662bar;
  wire n663bar;
  wire n664bar;
  wire n665bar;
  wire n666bar;
  wire n667bar;
  wire n668bar;
  wire n669bar;
  wire n670bar;
  wire n671bar;
  wire n672bar;
  wire n673bar;
  wire n674bar;
  wire n675bar;
  wire n676bar;
  wire n677bar;
  wire n678bar;
  wire n679bar;
  wire n680bar;
  wire n681bar;
  wire n682bar;
  wire n683bar;
  wire n684bar;
  wire n685bar;
  wire n686bar;
  wire n687bar;
  wire n688bar;
  wire n689bar;
  wire n690bar;
  wire n691bar;
  wire n692bar;
  wire n693bar;
  wire n694bar;
  wire n695bar;
  wire n696bar;
  wire n697bar;
  wire n698bar;
  wire n699bar;
  wire n700bar;
  wire n701bar;
  wire n702bar;
  wire n703bar;
  wire n704bar;
  wire n705bar;
  wire n706bar;
  wire n707bar;
  wire n708bar;
  wire n709bar;
  wire n710bar;
  wire n711bar;
  wire n712bar;
  wire n713bar;
  wire n714bar;
  wire n715bar;
  wire n716bar;
  wire n717bar;
  wire n718bar;
  wire n719bar;
  wire n720bar;
  wire n721bar;
  wire n722bar;
  wire n723bar;
  wire n724bar;
  wire n725bar;
  wire n726bar;
  wire n727bar;
  wire n728bar;
  wire n729bar;
  wire n730bar;
  wire n731bar;
  wire n732bar;
  wire n733bar;
  wire n734bar;
  wire n735bar;
  wire n736bar;
  wire n737bar;
  wire n738bar;
  wire n739bar;
  wire n740bar;
  wire n741bar;
  wire n742bar;
  wire n743bar;
  wire n744bar;
  wire n745bar;
  wire n746bar;
  wire n747bar;
  wire n748bar;
  wire n749bar;
  wire n750bar;
  wire n751bar;
  wire n752bar;
  wire n753bar;
  wire n754bar;
  wire n755bar;
  wire n756bar;
  wire n757bar;
  wire n758bar;
  wire n759bar;
  wire n760bar;
  wire n761bar;
  wire n762bar;
  wire n763bar;
  wire n764bar;
  wire n765bar;
  wire n766bar;
  wire n767bar;
  wire n768bar;
  wire n769bar;
  wire n770bar;
  wire n771bar;
  wire n772bar;
  wire n773bar;
  wire n774bar;
  wire n775bar;
  wire n776bar;
  wire n777bar;
  wire n778bar;
  wire n779bar;
  wire n780bar;
  wire n781bar;
  wire n782bar;
  wire n783bar;
  wire n784bar;
  wire n785bar;
  wire n786bar;
  wire n787bar;
  wire n788bar;
  wire n789bar;
  wire n790bar;
  wire n791bar;
  wire n792bar;
  wire n793bar;
  wire n794bar;
  wire n795bar;
  wire n796bar;
  wire n797bar;
  wire n798bar;
  wire n799bar;
  wire n800bar;
  wire n801bar;
  wire n802bar;
  wire n803bar;
  wire n804bar;
  wire n805bar;
  wire n806bar;
  wire n807bar;
  wire n808bar;
  wire n809bar;
  wire n810bar;
  wire n811bar;
  wire n812bar;
  wire n813bar;
  wire n814bar;
  wire n815bar;
  wire n816bar;
  wire n817bar;
  wire n818bar;
  wire n819bar;
  wire n820bar;
  wire n821bar;
  wire n822bar;
  wire n823bar;
  wire n824bar;
  wire n825bar;
  wire n826bar;
  wire n827bar;
  wire n828bar;
  wire n829bar;
  wire n830bar;
  wire n831bar;
  wire n832bar;
  wire n833bar;
  wire n834bar;
  wire n835bar;
  wire n836bar;
  wire n837bar;
  wire n838bar;
  wire n839bar;
  wire n840bar;
  wire n841bar;
  wire n842bar;
  wire n843bar;
  wire n844bar;
  wire n845bar;
  wire n846bar;
  wire n847bar;
  wire n848bar;
  wire n849bar;
  wire n850bar;
  wire n851bar;
  wire n852bar;
  wire n853bar;
  wire n854bar;
  wire n855bar;
  wire n856bar;
  wire n857bar;
  wire n858bar;
  wire n859bar;
  wire n860bar;
  wire n861bar;
  wire n862bar;
  wire n863bar;
  wire n864bar;
  wire n865bar;
  wire n866bar;
  wire n867bar;
  wire n868bar;
  wire n869bar;
  wire n870bar;
  wire n871bar;
  wire n872bar;
  wire n873bar;
  wire n874bar;
  wire n875bar;
  wire n876bar;
  wire n877bar;
  wire n878bar;
  wire n879bar;
  wire n880bar;
  wire n881bar;
  wire n882bar;
  wire n883bar;
  wire n884bar;
  wire n885bar;
  wire n886bar;
  wire n887bar;
  wire n888bar;
  wire n889bar;
  wire n890bar;
  wire n891bar;
  wire n892bar;
  wire n893bar;
  wire n894bar;
  wire n895bar;
  wire n896bar;
  wire n897bar;
  wire n898bar;
  wire n899bar;
  wire n900bar;
  wire n901bar;
  wire n902bar;
  wire n903bar;
  wire n904bar;
  wire n905bar;
  wire n906bar;
  wire n907bar;
  wire n908bar;
  wire n909bar;
  wire n910bar;
  wire n911bar;
  wire n912bar;
  wire n913bar;
  wire n914bar;
  wire n915bar;
  wire n916bar;
  wire n917bar;
  wire n918bar;
  wire n919bar;
  wire n920bar;
  wire n921bar;
  wire n922bar;
  wire n923bar;
  wire n924bar;
  wire n925bar;
  wire n926bar;
  wire n927bar;
  wire n928bar;
  wire n929bar;
  wire n930bar;
  wire n931bar;
  wire n932bar;
  wire n933bar;
  wire n934bar;
  wire n935bar;
  wire n936bar;
  wire n937bar;
  wire n938bar;
  wire n939bar;
  wire n940bar;
  wire n941bar;
  wire n942bar;
  wire n943bar;
  wire n944bar;
  wire n945bar;
  wire n946bar;
  wire n947bar;
  wire n948bar;
  wire n949bar;
  wire n950bar;
  wire n951bar;
  wire n952bar;
  wire n953bar;
  wire n954bar;
  wire n955bar;
  wire n956bar;
  wire n957bar;
  wire n958bar;
  wire n959bar;
  wire n960bar;
  wire n961bar;
  wire n962bar;
  wire n963bar;
  wire n964bar;
  wire n965bar;
  wire n966bar;
  wire n967bar;
  wire n968bar;
  wire n969bar;
  wire n970bar;
  wire n971bar;
  wire n972bar;
//wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];
  //OR U1
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1 (
    .O(out[7]),
    .I0(n972),
    .I1(n971)
  );
  //AND U1bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1bar (
    .O(outbar[7]),
    .I0(n972bar),
    .I1(n971bar)
  );
  //OR U2
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2 (
    .O(n971),
    .I0(n970),
    .I1(n969)
  );
  //AND U2bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2bar (
    .O(n971bar),
    .I0(n970bar),
    .I1(n969bar)
  );
  //OR U3
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3 (
    .O(n969),
    .I0(n968),
    .I1(n967)
  );
  //AND U3bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3bar (
    .O(n969bar),
    .I0(n968bar),
    .I1(n967bar)
  );
  //OR U4
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4 (
    .O(n967),
    .I0(n966),
    .I1(n965)
  );
  //AND U4bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4bar (
    .O(n967bar),
    .I0(n966bar),
    .I1(n965bar)
  );
  //OR U5
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5 (
    .O(n968),
    .I0(n964),
    .I1(n963)
  );
  //AND U5bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5bar (
    .O(n968bar),
    .I0(n964bar),
    .I1(n963bar)
  );
  //OR U6
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6 (
    .O(n963),
    .I0(in[116]),
    .I1(n962)
  );
  //AND U6bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6bar (
    .O(n963bar),
    .I0(inbar[116]),
    .I1(n962bar)
  );
  //OR U7
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7 (
    .O(n970),
    .I0(n961),
    .I1(n960)
  );
  //AND U7bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7bar (
    .O(n970bar),
    .I0(n961bar),
    .I1(n960bar)
  );
  //OR U8
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8 (
    .O(n960),
    .I0(in[150]),
    .I1(in[127])
  );
  //AND U8bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8bar (
    .O(n960bar),
    .I0(inbar[150]),
    .I1(inbar[127])
  );
  //OR U9
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9 (
    .O(n961),
    .I0(in[160]),
    .I1(n959)
  );
  //AND U9bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9bar (
    .O(n961bar),
    .I0(inbar[160]),
    .I1(n959bar)
  );
  //OR U10
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10 (
    .O(n959),
    .I0(in[252]),
    .I1(in[168])
  );
  //AND U10bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10bar (
    .O(n959bar),
    .I0(inbar[252]),
    .I1(inbar[168])
  );
  //OR U11
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11 (
    .O(n972),
    .I0(n958),
    .I1(n957)
  );
  //AND U11bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11bar (
    .O(n972bar),
    .I0(n958bar),
    .I1(n957bar)
  );
  //OR U12
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12 (
    .O(n957),
    .I0(n956),
    .I1(n955)
  );
  //AND U12bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12bar (
    .O(n957bar),
    .I0(n956bar),
    .I1(n955bar)
  );
  //OR U13
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13 (
    .O(n955),
    .I0(in_17),
    .I1(in[96])
  );
  //AND U13bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13bar (
    .O(n955bar),
    .I0(in_17bar),
    .I1(inbar[96])
  );
  //OR U14
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14 (
    .O(n956),
    .I0(in_23),
    .I1(n954)
  );
  //AND U14bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14bar (
    .O(n956bar),
    .I0(in_23bar),
    .I1(n954bar)
  );
  //OR U15
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15 (
    .O(n954),
    .I0(in_31),
    .I1(in_26)
  );
  //AND U15bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15bar (
    .O(n954bar),
    .I0(in_31bar),
    .I1(in_26bar)
  );
  //OR U16
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16 (
    .O(n958),
    .I0(n953),
    .I1(n952)
  );
  //AND U16bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16bar (
    .O(n958bar),
    .I0(n953bar),
    .I1(n952bar)
  );
  //OR U17
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U17 (
    .O(n952),
    .I0(in_58),
    .I1(in_4)
  );
  //AND U17bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U17bar (
    .O(n952bar),
    .I0(in_58bar),
    .I1(in_4bar)
  );
  //OR U18
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U18 (
    .O(n953),
    .I0(in_59),
    .I1(n951)
  );
  //AND U18bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U18bar (
    .O(n953bar),
    .I0(in_59bar),
    .I1(n951bar)
  );
  //OR U19
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U19 (
    .O(n951),
    .I0(in_71),
    .I1(in_62)
  );
  //AND U19bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U19bar (
    .O(n951bar),
    .I0(in_71bar),
    .I1(in_62bar)
  );
  //OR U20
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U20 (
    .O(out[6]),
    .I0(n950),
    .I1(n949)
  );
  //AND U20bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U20bar (
    .O(outbar[6]),
    .I0(n950bar),
    .I1(n949bar)
  );
  //OR U21
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U21 (
    .O(n949),
    .I0(n948),
    .I1(n947)
  );
  //AND U21bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U21bar (
    .O(n949bar),
    .I0(n948bar),
    .I1(n947bar)
  );
  //OR U22
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U22 (
    .O(n947),
    .I0(n946),
    .I1(n945)
  );
  //AND U22bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U22bar (
    .O(n947bar),
    .I0(n946bar),
    .I1(n945bar)
  );
  //OR U23
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U23 (
    .O(n945),
    .I0(n944),
    .I1(n943)
  );
  //AND U23bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U23bar (
    .O(n945bar),
    .I0(n944bar),
    .I1(n943bar)
  );
  //OR U24
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U24 (
    .O(n946),
    .I0(n942),
    .I1(n941)
  );
  //AND U24bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U24bar (
    .O(n946bar),
    .I0(n942bar),
    .I1(n941bar)
  );
  //OR U25
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U25 (
    .O(n941),
    .I0(in[101]),
    .I1(n940)
  );
  //AND U25bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U25bar (
    .O(n941bar),
    .I0(inbar[101]),
    .I1(n940bar)
  );
  //OR U26
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U26 (
    .O(n948),
    .I0(n939),
    .I1(n938)
  );
  //AND U26bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U26bar (
    .O(n948bar),
    .I0(n939bar),
    .I1(n938bar)
  );
  //OR U27
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U27 (
    .O(n938),
    .I0(in[114]),
    .I1(in[104])
  );
  //AND U27bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U27bar (
    .O(n938bar),
    .I0(inbar[114]),
    .I1(inbar[104])
  );
  //OR U28
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U28 (
    .O(n939),
    .I0(in[128]),
    .I1(n937)
  );
  //AND U28bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U28bar (
    .O(n939bar),
    .I0(inbar[128]),
    .I1(n937bar)
  );
  //OR U29
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U29 (
    .O(n937),
    .I0(in[136]),
    .I1(in[134])
  );
  //AND U29bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U29bar (
    .O(n937bar),
    .I0(inbar[136]),
    .I1(inbar[134])
  );
  //OR U30
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U30 (
    .O(n950),
    .I0(n936),
    .I1(n935)
  );
  //AND U30bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U30bar (
    .O(n950bar),
    .I0(n936bar),
    .I1(n935bar)
  );
  //OR U31
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U31 (
    .O(n935),
    .I0(n934),
    .I1(n933)
  );
  //AND U31bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U31bar (
    .O(n935bar),
    .I0(n934bar),
    .I1(n933bar)
  );
  //OR U32
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U32 (
    .O(n933),
    .I0(in[177]),
    .I1(in[164])
  );
  //AND U32bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U32bar (
    .O(n933bar),
    .I0(inbar[177]),
    .I1(inbar[164])
  );
  //OR U33
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U33 (
    .O(n934),
    .I0(in[212]),
    .I1(n932)
  );
  //AND U33bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U33bar (
    .O(n934bar),
    .I0(inbar[212]),
    .I1(n932bar)
  );
  //OR U34
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U34 (
    .O(n932),
    .I0(in[248]),
    .I1(in[221])
  );
  //AND U34bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U34bar (
    .O(n932bar),
    .I0(inbar[248]),
    .I1(inbar[221])
  );
  //OR U35
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U35 (
    .O(n936),
    .I0(n931),
    .I1(n930)
  );
  //AND U35bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U35bar (
    .O(n936bar),
    .I0(n931bar),
    .I1(n930bar)
  );
  //OR U36
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U36 (
    .O(n930),
    .I0(in_18),
    .I1(in[93])
  );
  //AND U36bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U36bar (
    .O(n930bar),
    .I0(in_18bar),
    .I1(inbar[93])
  );
  //OR U37
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U37 (
    .O(n931),
    .I0(in_31),
    .I1(n929)
  );
  //AND U37bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U37bar (
    .O(n931bar),
    .I0(in_31bar),
    .I1(n929bar)
  );
  //OR U38
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U38 (
    .O(n929),
    .I0(in_7),
    .I1(in_39)
  );
  //AND U38bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U38bar (
    .O(n929bar),
    .I0(in_7bar),
    .I1(in_39bar)
  );
  //OR U39
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U39 (
    .O(out[5]),
    .I0(n928),
    .I1(n927)
  );
  //AND U39bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U39bar (
    .O(outbar[5]),
    .I0(n928bar),
    .I1(n927bar)
  );
  //OR U40
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U40 (
    .O(n927),
    .I0(n926),
    .I1(n925)
  );
  //AND U40bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U40bar (
    .O(n927bar),
    .I0(n926bar),
    .I1(n925bar)
  );
  //OR U41
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U41 (
    .O(n925),
    .I0(n924),
    .I1(n923)
  );
  //AND U41bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U41bar (
    .O(n925bar),
    .I0(n924bar),
    .I1(n923bar)
  );
  //OR U42
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U42 (
    .O(n923),
    .I0(n922),
    .I1(n921)
  );
  //AND U42bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U42bar (
    .O(n923bar),
    .I0(n922bar),
    .I1(n921bar)
  );
  //OR U43
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U43 (
    .O(n924),
    .I0(n940),
    .I1(n920)
  );
  //AND U43bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U43bar (
    .O(n924bar),
    .I0(n940bar),
    .I1(n920bar)
  );
  //OR U44
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U44 (
    .O(n920),
    .I0(in[111]),
    .I1(n919)
  );
  //AND U44bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U44bar (
    .O(n920bar),
    .I0(inbar[111]),
    .I1(n919bar)
  );
  //OR U45
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U45 (
    .O(n940),
    .I0(n918),
    .I1(n917)
  );
  //AND U45bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U45bar (
    .O(n940bar),
    .I0(n918bar),
    .I1(n917bar)
  );
  //OR U46
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U46 (
    .O(n917),
    .I0(n916),
    .I1(n915)
  );
  //AND U46bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U46bar (
    .O(n917bar),
    .I0(n916bar),
    .I1(n915bar)
  );
  //OR U47
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U47 (
    .O(n915),
    .I0(n914),
    .I1(n913)
  );
  //AND U47bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U47bar (
    .O(n915bar),
    .I0(n914bar),
    .I1(n913bar)
  );
  //OR U48
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U48 (
    .O(n913),
    .I0(in[140]),
    .I1(in[131])
  );
  //AND U48bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U48bar (
    .O(n913bar),
    .I0(inbar[140]),
    .I1(inbar[131])
  );
  //OR U49
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U49 (
    .O(n914),
    .I0(in[160]),
    .I1(in[144])
  );
  //AND U49bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U49bar (
    .O(n914bar),
    .I0(inbar[160]),
    .I1(inbar[144])
  );
  //OR U50
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U50 (
    .O(n916),
    .I0(n912),
    .I1(n911)
  );
  //AND U50bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U50bar (
    .O(n916bar),
    .I0(n912bar),
    .I1(n911bar)
  );
  //OR U51
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U51 (
    .O(n911),
    .I0(in[179]),
    .I1(in[174])
  );
  //AND U51bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U51bar (
    .O(n911bar),
    .I0(inbar[179]),
    .I1(inbar[174])
  );
  //OR U52
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U52 (
    .O(n912),
    .I0(in[188]),
    .I1(in[184])
  );
  //AND U52bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U52bar (
    .O(n912bar),
    .I0(inbar[188]),
    .I1(inbar[184])
  );
  //OR U53
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U53 (
    .O(n918),
    .I0(n910),
    .I1(n909)
  );
  //AND U53bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U53bar (
    .O(n918bar),
    .I0(n910bar),
    .I1(n909bar)
  );
  //OR U54
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U54 (
    .O(n909),
    .I0(n908),
    .I1(n907)
  );
  //AND U54bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U54bar (
    .O(n909bar),
    .I0(n908bar),
    .I1(n907bar)
  );
  //OR U55
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U55 (
    .O(n907),
    .I0(in[216]),
    .I1(in[200])
  );
  //AND U55bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U55bar (
    .O(n907bar),
    .I0(inbar[216]),
    .I1(inbar[200])
  );
  //OR U56
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U56 (
    .O(n908),
    .I0(in[228]),
    .I1(in[224])
  );
  //AND U56bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U56bar (
    .O(n908bar),
    .I0(inbar[228]),
    .I1(inbar[224])
  );
  //OR U57
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U57 (
    .O(n910),
    .I0(n906),
    .I1(n905)
  );
  //AND U57bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U57bar (
    .O(n910bar),
    .I0(n906bar),
    .I1(n905bar)
  );
  //OR U58
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U58 (
    .O(n905),
    .I0(in[247]),
    .I1(in[235])
  );
  //AND U58bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U58bar (
    .O(n905bar),
    .I0(inbar[247]),
    .I1(inbar[235])
  );
  //OR U59
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U59 (
    .O(n906),
    .I0(in_42),
    .I1(in[83])
  );
  //AND U59bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U59bar (
    .O(n906bar),
    .I0(in_42bar),
    .I1(inbar[83])
  );
  //OR U60
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U60 (
    .O(n926),
    .I0(n904),
    .I1(n903)
  );
  //AND U60bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U60bar (
    .O(n926bar),
    .I0(n904bar),
    .I1(n903bar)
  );
  //OR U61
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U61 (
    .O(n903),
    .I0(in[166]),
    .I1(in[123])
  );
  //AND U61bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U61bar (
    .O(n903bar),
    .I0(inbar[166]),
    .I1(inbar[123])
  );
  //OR U62
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U62 (
    .O(n904),
    .I0(in[170]),
    .I1(n902)
  );
  //AND U62bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U62bar (
    .O(n904bar),
    .I0(inbar[170]),
    .I1(n902bar)
  );
  //OR U63
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U63 (
    .O(n902),
    .I0(in[194]),
    .I1(in[183])
  );
  //AND U63bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U63bar (
    .O(n902bar),
    .I0(inbar[194]),
    .I1(inbar[183])
  );
  //OR U64
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U64 (
    .O(n928),
    .I0(n901),
    .I1(n900)
  );
  //AND U64bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U64bar (
    .O(n928bar),
    .I0(n901bar),
    .I1(n900bar)
  );
  //OR U65
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U65 (
    .O(n900),
    .I0(n899),
    .I1(n898)
  );
  //AND U65bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U65bar (
    .O(n900bar),
    .I0(n899bar),
    .I1(n898bar)
  );
  //OR U66
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U66 (
    .O(n898),
    .I0(in[241]),
    .I1(in[238])
  );
  //AND U66bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U66bar (
    .O(n898bar),
    .I0(inbar[241]),
    .I1(inbar[238])
  );
  //OR U67
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U67 (
    .O(n899),
    .I0(in[250]),
    .I1(n897)
  );
  //AND U67bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U67bar (
    .O(n899bar),
    .I0(inbar[250]),
    .I1(n897bar)
  );
  //OR U68
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U68 (
    .O(n897),
    .I0(in_24),
    .I1(in[84])
  );
  //AND U68bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U68bar (
    .O(n897bar),
    .I0(in_24bar),
    .I1(inbar[84])
  );
  //OR U69
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U69 (
    .O(n901),
    .I0(n896),
    .I1(n895)
  );
  //AND U69bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U69bar (
    .O(n901bar),
    .I0(n896bar),
    .I1(n895bar)
  );
  //OR U70
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U70 (
    .O(n895),
    .I0(in_41),
    .I1(in_29)
  );
  //AND U70bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U70bar (
    .O(n895bar),
    .I0(in_41bar),
    .I1(in_29bar)
  );
  //OR U71
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U71 (
    .O(n896),
    .I0(in_66),
    .I1(n894)
  );
  //AND U71bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U71bar (
    .O(n896bar),
    .I0(in_66bar),
    .I1(n894bar)
  );
  //OR U72
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U72 (
    .O(n894),
    .I0(in_76),
    .I1(in_71)
  );
  //AND U72bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U72bar (
    .O(n894bar),
    .I0(in_76bar),
    .I1(in_71bar)
  );
  //OR U73
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U73 (
    .O(out[4]),
    .I0(n893),
    .I1(n892)
  );
  //AND U73bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U73bar (
    .O(outbar[4]),
    .I0(n893bar),
    .I1(n892bar)
  );
  //OR U74
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U74 (
    .O(n892),
    .I0(n891),
    .I1(n890)
  );
  //AND U74bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U74bar (
    .O(n892bar),
    .I0(n891bar),
    .I1(n890bar)
  );
  //OR U75
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U75 (
    .O(n890),
    .I0(n889),
    .I1(n888)
  );
  //AND U75bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U75bar (
    .O(n890bar),
    .I0(n889bar),
    .I1(n888bar)
  );
  //OR U76
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U76 (
    .O(n888),
    .I0(n922),
    .I1(n887)
  );
  //AND U76bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U76bar (
    .O(n888bar),
    .I0(n922bar),
    .I1(n887bar)
  );
  //OR U77
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U77 (
    .O(n922),
    .I0(n886),
    .I1(n885)
  );
  //AND U77bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U77bar (
    .O(n922bar),
    .I0(n886bar),
    .I1(n885bar)
  );
  //OR U78
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U78 (
    .O(n885),
    .I0(n884),
    .I1(n883)
  );
  //AND U78bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U78bar (
    .O(n885bar),
    .I0(n884bar),
    .I1(n883bar)
  );
  //OR U79
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U79 (
    .O(n883),
    .I0(n882),
    .I1(n881)
  );
  //AND U79bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U79bar (
    .O(n883bar),
    .I0(n882bar),
    .I1(n881bar)
  );
  //OR U80
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U80 (
    .O(n881),
    .I0(in[118]),
    .I1(in[109])
  );
  //AND U80bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U80bar (
    .O(n881bar),
    .I0(inbar[118]),
    .I1(inbar[109])
  );
  //OR U81
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U81 (
    .O(n882),
    .I0(in[139]),
    .I1(in[120])
  );
  //AND U81bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U81bar (
    .O(n882bar),
    .I0(inbar[139]),
    .I1(inbar[120])
  );
  //OR U82
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U82 (
    .O(n884),
    .I0(n880),
    .I1(n879)
  );
  //AND U82bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U82bar (
    .O(n884bar),
    .I0(n880bar),
    .I1(n879bar)
  );
  //OR U83
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U83 (
    .O(n879),
    .I0(in[198]),
    .I1(in[154])
  );
  //AND U83bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U83bar (
    .O(n879bar),
    .I0(inbar[198]),
    .I1(inbar[154])
  );
  //OR U84
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U84 (
    .O(n880),
    .I0(in[210]),
    .I1(in[205])
  );
  //AND U84bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U84bar (
    .O(n880bar),
    .I0(inbar[210]),
    .I1(inbar[205])
  );
  //OR U85
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U85 (
    .O(n886),
    .I0(n878),
    .I1(n877)
  );
  //AND U85bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U85bar (
    .O(n886bar),
    .I0(n878bar),
    .I1(n877bar)
  );
  //OR U86
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U86 (
    .O(n877),
    .I0(n876),
    .I1(n875)
  );
  //AND U86bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U86bar (
    .O(n877bar),
    .I0(n876bar),
    .I1(n875bar)
  );
  //OR U87
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U87 (
    .O(n875),
    .I0(in[219]),
    .I1(in[217])
  );
  //AND U87bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U87bar (
    .O(n875bar),
    .I0(inbar[219]),
    .I1(inbar[217])
  );
  //OR U88
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U88 (
    .O(n876),
    .I0(in[86]),
    .I1(in[252])
  );
  //AND U88bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U88bar (
    .O(n876bar),
    .I0(inbar[86]),
    .I1(inbar[252])
  );
  //OR U89
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U89 (
    .O(n878),
    .I0(n874),
    .I1(n873)
  );
  //AND U89bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U89bar (
    .O(n878bar),
    .I0(n874bar),
    .I1(n873bar)
  );
  //OR U90
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U90 (
    .O(n873),
    .I0(in_40),
    .I1(in[91])
  );
  //AND U90bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U90bar (
    .O(n873bar),
    .I0(in_40bar),
    .I1(inbar[91])
  );
  //OR U91
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U91 (
    .O(n874),
    .I0(in_8),
    .I1(in_46)
  );
  //AND U91bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U91bar (
    .O(n874bar),
    .I0(in_8bar),
    .I1(in_46bar)
  );
  //OR U92
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U92 (
    .O(n889),
    .I0(n872),
    .I1(n871)
  );
  //AND U92bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U92bar (
    .O(n889bar),
    .I0(n872bar),
    .I1(n871bar)
  );
  //OR U93
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U93 (
    .O(n871),
    .I0(in[117]),
    .I1(n943)
  );
  //AND U93bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U93bar (
    .O(n871bar),
    .I0(inbar[117]),
    .I1(n943bar)
  );
  //OR U94
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U94 (
    .O(n943),
    .I0(n870),
    .I1(n869)
  );
  //AND U94bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U94bar (
    .O(n943bar),
    .I0(n870bar),
    .I1(n869bar)
  );
  //OR U95
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U95 (
    .O(n869),
    .I0(n868),
    .I1(n867)
  );
  //AND U95bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U95bar (
    .O(n869bar),
    .I0(n868bar),
    .I1(n867bar)
  );
  //OR U96
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U96 (
    .O(n867),
    .I0(n866),
    .I1(n865)
  );
  //AND U96bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U96bar (
    .O(n867bar),
    .I0(n866bar),
    .I1(n865bar)
  );
  //OR U97
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U97 (
    .O(n865),
    .I0(n864),
    .I1(n863)
  );
  //AND U97bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U97bar (
    .O(n865bar),
    .I0(n864bar),
    .I1(n863bar)
  );
  //OR U98
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U98 (
    .O(n866),
    .I0(in[108]),
    .I1(n919)
  );
  //AND U98bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U98bar (
    .O(n866bar),
    .I0(inbar[108]),
    .I1(n919bar)
  );
  //OR U99
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U99 (
    .O(n919),
    .I0(n862),
    .I1(n861)
  );
  //AND U99bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U99bar (
    .O(n919bar),
    .I0(n862bar),
    .I1(n861bar)
  );
  //OR U100
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U100 (
    .O(n861),
    .I0(n860),
    .I1(n859)
  );
  //AND U100bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U100bar (
    .O(n861bar),
    .I0(n860bar),
    .I1(n859bar)
  );
  //OR U101
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U101 (
    .O(n859),
    .I0(n858),
    .I1(n857)
  );
  //AND U101bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U101bar (
    .O(n859bar),
    .I0(n858bar),
    .I1(n857bar)
  );
  //OR U102
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U102 (
    .O(n857),
    .I0(in[119]),
    .I1(in[105])
  );
  //AND U102bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U102bar (
    .O(n857bar),
    .I0(inbar[119]),
    .I1(inbar[105])
  );
  //OR U103
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U103 (
    .O(n858),
    .I0(in[186]),
    .I1(in[175])
  );
  //AND U103bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U103bar (
    .O(n858bar),
    .I0(inbar[186]),
    .I1(inbar[175])
  );
  //OR U104
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U104 (
    .O(n860),
    .I0(n856),
    .I1(n855)
  );
  //AND U104bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U104bar (
    .O(n860bar),
    .I0(n856bar),
    .I1(n855bar)
  );
  //OR U105
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U105 (
    .O(n855),
    .I0(in[202]),
    .I1(in[193])
  );
  //AND U105bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U105bar (
    .O(n855bar),
    .I0(inbar[202]),
    .I1(inbar[193])
  );
  //OR U106
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U106 (
    .O(n856),
    .I0(in[225]),
    .I1(in[208])
  );
  //AND U106bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U106bar (
    .O(n856bar),
    .I0(inbar[225]),
    .I1(inbar[208])
  );
  //OR U107
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U107 (
    .O(n862),
    .I0(n854),
    .I1(n853)
  );
  //AND U107bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U107bar (
    .O(n862bar),
    .I0(n854bar),
    .I1(n853bar)
  );
  //OR U108
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U108 (
    .O(n853),
    .I0(n852),
    .I1(n851)
  );
  //AND U108bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U108bar (
    .O(n853bar),
    .I0(n852bar),
    .I1(n851bar)
  );
  //OR U109
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U109 (
    .O(n851),
    .I0(in_1),
    .I1(in[85])
  );
  //AND U109bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U109bar (
    .O(n851bar),
    .I0(in_1bar),
    .I1(inbar[85])
  );
  //OR U110
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U110 (
    .O(n852),
    .I0(in_23),
    .I1(in_19)
  );
  //AND U110bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U110bar (
    .O(n852bar),
    .I0(in_23bar),
    .I1(in_19bar)
  );
  //OR U111
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U111 (
    .O(n854),
    .I0(n850),
    .I1(n849)
  );
  //AND U111bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U111bar (
    .O(n854bar),
    .I0(n850bar),
    .I1(n849bar)
  );
  //OR U112
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U112 (
    .O(n849),
    .I0(in_43),
    .I1(in_33)
  );
  //AND U112bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U112bar (
    .O(n849bar),
    .I0(in_43bar),
    .I1(in_33bar)
  );
  //OR U113
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U113 (
    .O(n850),
    .I0(in_63),
    .I1(in_44)
  );
  //AND U113bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U113bar (
    .O(n850bar),
    .I0(in_63bar),
    .I1(in_44bar)
  );
  //OR U114
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U114 (
    .O(n868),
    .I0(n848),
    .I1(n847)
  );
  //AND U114bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U114bar (
    .O(n868bar),
    .I0(n848bar),
    .I1(n847bar)
  );
  //OR U115
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U115 (
    .O(n847),
    .I0(in[141]),
    .I1(in[112])
  );
  //AND U115bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U115bar (
    .O(n847bar),
    .I0(inbar[141]),
    .I1(inbar[112])
  );
  //OR U116
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U116 (
    .O(n848),
    .I0(in[147]),
    .I1(n846)
  );
  //AND U116bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U116bar (
    .O(n848bar),
    .I0(inbar[147]),
    .I1(n846bar)
  );
  //OR U117
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U117 (
    .O(n846),
    .I0(in[181]),
    .I1(in[167])
  );
  //AND U117bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U117bar (
    .O(n846bar),
    .I0(inbar[181]),
    .I1(inbar[167])
  );
  //OR U118
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U118 (
    .O(n870),
    .I0(n845),
    .I1(n844)
  );
  //AND U118bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U118bar (
    .O(n870bar),
    .I0(n845bar),
    .I1(n844bar)
  );
  //OR U119
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U119 (
    .O(n844),
    .I0(n843),
    .I1(n842)
  );
  //AND U119bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U119bar (
    .O(n844bar),
    .I0(n843bar),
    .I1(n842bar)
  );
  //OR U120
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U120 (
    .O(n842),
    .I0(in[229]),
    .I1(in[201])
  );
  //AND U120bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U120bar (
    .O(n842bar),
    .I0(inbar[229]),
    .I1(inbar[201])
  );
  //OR U121
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U121 (
    .O(n843),
    .I0(in[237]),
    .I1(n841)
  );
  //AND U121bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U121bar (
    .O(n843bar),
    .I0(inbar[237]),
    .I1(n841bar)
  );
  //OR U122
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U122 (
    .O(n841),
    .I0(in[94]),
    .I1(in[253])
  );
  //AND U122bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U122bar (
    .O(n841bar),
    .I0(inbar[94]),
    .I1(inbar[253])
  );
  //OR U123
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U123 (
    .O(n845),
    .I0(n840),
    .I1(n839)
  );
  //AND U123bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U123bar (
    .O(n845bar),
    .I0(n840bar),
    .I1(n839bar)
  );
  //OR U124
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U124 (
    .O(n839),
    .I0(in_21),
    .I1(in[96])
  );
  //AND U124bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U124bar (
    .O(n839bar),
    .I0(in_21bar),
    .I1(inbar[96])
  );
  //OR U125
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U125 (
    .O(n840),
    .I0(in_25),
    .I1(n838)
  );
  //AND U125bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U125bar (
    .O(n840bar),
    .I0(in_25bar),
    .I1(n838bar)
  );
  //OR U126
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U126 (
    .O(n838),
    .I0(in_81),
    .I1(in_45)
  );
  //AND U126bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U126bar (
    .O(n838bar),
    .I0(in_81bar),
    .I1(in_45bar)
  );
  //OR U127
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U127 (
    .O(n891),
    .I0(n837),
    .I1(n836)
  );
  //AND U127bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U127bar (
    .O(n891bar),
    .I0(n837bar),
    .I1(n836bar)
  );
  //OR U128
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U128 (
    .O(n836),
    .I0(in[142]),
    .I1(in[124])
  );
  //AND U128bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U128bar (
    .O(n836bar),
    .I0(inbar[142]),
    .I1(inbar[124])
  );
  //OR U129
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U129 (
    .O(n837),
    .I0(in[150]),
    .I1(n835)
  );
  //AND U129bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U129bar (
    .O(n837bar),
    .I0(inbar[150]),
    .I1(n835bar)
  );
  //OR U130
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U130 (
    .O(n835),
    .I0(in[172]),
    .I1(in[155])
  );
  //AND U130bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U130bar (
    .O(n835bar),
    .I0(inbar[172]),
    .I1(inbar[155])
  );
  //OR U131
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U131 (
    .O(n893),
    .I0(n834),
    .I1(n833)
  );
  //AND U131bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U131bar (
    .O(n893bar),
    .I0(n834bar),
    .I1(n833bar)
  );
  //OR U132
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U132 (
    .O(n833),
    .I0(n832),
    .I1(n831)
  );
  //AND U132bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U132bar (
    .O(n833bar),
    .I0(n832bar),
    .I1(n831bar)
  );
  //OR U133
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U133 (
    .O(n831),
    .I0(in[196]),
    .I1(in[173])
  );
  //AND U133bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U133bar (
    .O(n831bar),
    .I0(inbar[196]),
    .I1(inbar[173])
  );
  //OR U134
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U134 (
    .O(n832),
    .I0(in[222]),
    .I1(n830)
  );
  //AND U134bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U134bar (
    .O(n832bar),
    .I0(inbar[222]),
    .I1(n830bar)
  );
  //OR U135
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U135 (
    .O(n830),
    .I0(in[227]),
    .I1(in[226])
  );
  //AND U135bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U135bar (
    .O(n830bar),
    .I0(inbar[227]),
    .I1(inbar[226])
  );
  //OR U136
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U136 (
    .O(n834),
    .I0(n829),
    .I1(n828)
  );
  //AND U136bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U136bar (
    .O(n834bar),
    .I0(n829bar),
    .I1(n828bar)
  );
  //OR U137
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U137 (
    .O(n828),
    .I0(in[249]),
    .I1(in[231])
  );
  //AND U137bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U137bar (
    .O(n828bar),
    .I0(inbar[249]),
    .I1(inbar[231])
  );
  //OR U138
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U138 (
    .O(n829),
    .I0(in_28),
    .I1(n827)
  );
  //AND U138bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U138bar (
    .O(n829bar),
    .I0(in_28bar),
    .I1(n827bar)
  );
  //OR U139
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U139 (
    .O(n827),
    .I0(in_52),
    .I1(in_47)
  );
  //AND U139bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U139bar (
    .O(n827bar),
    .I0(in_52bar),
    .I1(in_47bar)
  );
  //OR U140
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U140 (
    .O(out[3]),
    .I0(n826),
    .I1(n825)
  );
  //AND U140bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U140bar (
    .O(outbar[3]),
    .I0(n826bar),
    .I1(n825bar)
  );
  //OR U141
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U141 (
    .O(n825),
    .I0(n824),
    .I1(n823)
  );
  //AND U141bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U141bar (
    .O(n825bar),
    .I0(n824bar),
    .I1(n823bar)
  );
  //OR U142
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U142 (
    .O(n823),
    .I0(n822),
    .I1(n821)
  );
  //AND U142bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U142bar (
    .O(n823bar),
    .I0(n822bar),
    .I1(n821bar)
  );
  //OR U143
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U143 (
    .O(n821),
    .I0(n820),
    .I1(n819)
  );
  //AND U143bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U143bar (
    .O(n821bar),
    .I0(n820bar),
    .I1(n819bar)
  );
  //OR U144
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U144 (
    .O(n822),
    .I0(n964),
    .I1(n818)
  );
  //AND U144bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U144bar (
    .O(n822bar),
    .I0(n964bar),
    .I1(n818bar)
  );
  //OR U145
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U145 (
    .O(n818),
    .I0(in[118]),
    .I1(n817)
  );
  //AND U145bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U145bar (
    .O(n818bar),
    .I0(inbar[118]),
    .I1(n817bar)
  );
  //OR U146
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U146 (
    .O(n964),
    .I0(n816),
    .I1(n815)
  );
  //AND U146bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U146bar (
    .O(n964bar),
    .I0(n816bar),
    .I1(n815bar)
  );
  //OR U147
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U147 (
    .O(n815),
    .I0(n814),
    .I1(n813)
  );
  //AND U147bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U147bar (
    .O(n815bar),
    .I0(n814bar),
    .I1(n813bar)
  );
  //OR U148
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U148 (
    .O(n813),
    .I0(n812),
    .I1(n811)
  );
  //AND U148bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U148bar (
    .O(n813bar),
    .I0(n812bar),
    .I1(n811bar)
  );
  //OR U149
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U149 (
    .O(n811),
    .I0(in[122]),
    .I1(in[111])
  );
  //AND U149bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U149bar (
    .O(n811bar),
    .I0(inbar[122]),
    .I1(inbar[111])
  );
  //OR U150
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U150 (
    .O(n812),
    .I0(in[154]),
    .I1(in[151])
  );
  //AND U150bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U150bar (
    .O(n812bar),
    .I0(inbar[154]),
    .I1(inbar[151])
  );
  //OR U151
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U151 (
    .O(n814),
    .I0(n810),
    .I1(n809)
  );
  //AND U151bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U151bar (
    .O(n814bar),
    .I0(n810bar),
    .I1(n809bar)
  );
  //OR U152
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U152 (
    .O(n809),
    .I0(in[187]),
    .I1(in[177])
  );
  //AND U152bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U152bar (
    .O(n809bar),
    .I0(inbar[187]),
    .I1(inbar[177])
  );
  //OR U153
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U153 (
    .O(n810),
    .I0(in[200]),
    .I1(in[192])
  );
  //AND U153bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U153bar (
    .O(n810bar),
    .I0(inbar[200]),
    .I1(inbar[192])
  );
  //OR U154
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U154 (
    .O(n816),
    .I0(n808),
    .I1(n807)
  );
  //AND U154bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U154bar (
    .O(n816bar),
    .I0(n808bar),
    .I1(n807bar)
  );
  //OR U155
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U155 (
    .O(n807),
    .I0(n806),
    .I1(n805)
  );
  //AND U155bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U155bar (
    .O(n807bar),
    .I0(n806bar),
    .I1(n805bar)
  );
  //OR U156
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U156 (
    .O(n805),
    .I0(in[225]),
    .I1(in[207])
  );
  //AND U156bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U156bar (
    .O(n805bar),
    .I0(inbar[225]),
    .I1(inbar[207])
  );
  //OR U157
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U157 (
    .O(n806),
    .I0(in[98]),
    .I1(in[226])
  );
  //AND U157bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U157bar (
    .O(n806bar),
    .I0(inbar[98]),
    .I1(inbar[226])
  );
  //OR U158
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U158 (
    .O(n808),
    .I0(n804),
    .I1(n803)
  );
  //AND U158bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U158bar (
    .O(n808bar),
    .I0(n804bar),
    .I1(n803bar)
  );
  //OR U159
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U159 (
    .O(n803),
    .I0(in_20),
    .I1(in_16)
  );
  //AND U159bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U159bar (
    .O(n803bar),
    .I0(in_20bar),
    .I1(in_16bar)
  );
  //OR U160
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U160 (
    .O(n804),
    .I0(in_55),
    .I1(in_45)
  );
  //AND U160bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U160bar (
    .O(n804bar),
    .I0(in_55bar),
    .I1(in_45bar)
  );
  //OR U161
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U161 (
    .O(n824),
    .I0(n802),
    .I1(n801)
  );
  //AND U161bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U161bar (
    .O(n824bar),
    .I0(n802bar),
    .I1(n801bar)
  );
  //OR U162
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U162 (
    .O(n801),
    .I0(in[162]),
    .I1(in[149])
  );
  //AND U162bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U162bar (
    .O(n801bar),
    .I0(inbar[162]),
    .I1(inbar[149])
  );
  //OR U163
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U163 (
    .O(n802),
    .I0(in[163]),
    .I1(n800)
  );
  //AND U163bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U163bar (
    .O(n802bar),
    .I0(inbar[163]),
    .I1(n800bar)
  );
  //OR U164
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U164 (
    .O(n800),
    .I0(in[191]),
    .I1(in[189])
  );
  //AND U164bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U164bar (
    .O(n800bar),
    .I0(inbar[191]),
    .I1(inbar[189])
  );
  //OR U165
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U165 (
    .O(n826),
    .I0(n799),
    .I1(n798)
  );
  //AND U165bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U165bar (
    .O(n826bar),
    .I0(n799bar),
    .I1(n798bar)
  );
  //OR U166
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U166 (
    .O(n798),
    .I0(n797),
    .I1(n796)
  );
  //AND U166bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U166bar (
    .O(n798bar),
    .I0(n797bar),
    .I1(n796bar)
  );
  //OR U167
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U167 (
    .O(n796),
    .I0(in[212]),
    .I1(in[193])
  );
  //AND U167bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U167bar (
    .O(n796bar),
    .I0(inbar[212]),
    .I1(inbar[193])
  );
  //OR U168
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U168 (
    .O(n797),
    .I0(in[238]),
    .I1(n795)
  );
  //AND U168bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U168bar (
    .O(n797bar),
    .I0(inbar[238]),
    .I1(n795bar)
  );
  //OR U169
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U169 (
    .O(n795),
    .I0(in[88]),
    .I1(in[247])
  );
  //AND U169bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U169bar (
    .O(n795bar),
    .I0(inbar[88]),
    .I1(inbar[247])
  );
  //OR U170
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U170 (
    .O(n799),
    .I0(n794),
    .I1(n793)
  );
  //AND U170bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U170bar (
    .O(n799bar),
    .I0(n794bar),
    .I1(n793bar)
  );
  //OR U171
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U171 (
    .O(n793),
    .I0(in[94]),
    .I1(in[92])
  );
  //AND U171bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U171bar (
    .O(n793bar),
    .I0(inbar[94]),
    .I1(inbar[92])
  );
  //OR U172
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U172 (
    .O(n794),
    .I0(in_52),
    .I1(n792)
  );
  //AND U172bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U172bar (
    .O(n794bar),
    .I0(in_52bar),
    .I1(n792bar)
  );
  //OR U173
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U173 (
    .O(n792),
    .I0(in_70),
    .I1(in_67)
  );
  //AND U173bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U173bar (
    .O(n792bar),
    .I0(in_70bar),
    .I1(in_67bar)
  );
  //OR U174
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U174 (
    .O(out[2]),
    .I0(n791),
    .I1(n790)
  );
  //AND U174bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U174bar (
    .O(outbar[2]),
    .I0(n791bar),
    .I1(n790bar)
  );
  //OR U175
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U175 (
    .O(n790),
    .I0(n789),
    .I1(n788)
  );
  //AND U175bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U175bar (
    .O(n790bar),
    .I0(n789bar),
    .I1(n788bar)
  );
  //OR U176
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U176 (
    .O(n788),
    .I0(n787),
    .I1(n786)
  );
  //AND U176bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U176bar (
    .O(n788bar),
    .I0(n787bar),
    .I1(n786bar)
  );
  //OR U177
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U177 (
    .O(n786),
    .I0(n819),
    .I1(n785)
  );
  //AND U177bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U177bar (
    .O(n786bar),
    .I0(n819bar),
    .I1(n785bar)
  );
  //OR U178
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U178 (
    .O(n819),
    .I0(n784),
    .I1(n783)
  );
  //AND U178bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U178bar (
    .O(n819bar),
    .I0(n784bar),
    .I1(n783bar)
  );
  //OR U179
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U179 (
    .O(n783),
    .I0(n782),
    .I1(n781)
  );
  //AND U179bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U179bar (
    .O(n783bar),
    .I0(n782bar),
    .I1(n781bar)
  );
  //OR U180
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U180 (
    .O(n781),
    .I0(n780),
    .I1(n779)
  );
  //AND U180bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U180bar (
    .O(n781bar),
    .I0(n780bar),
    .I1(n779bar)
  );
  //OR U181
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U181 (
    .O(n779),
    .I0(n962),
    .I1(n778)
  );
  //AND U181bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U181bar (
    .O(n779bar),
    .I0(n962bar),
    .I1(n778bar)
  );
  //OR U182
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U182 (
    .O(n962),
    .I0(n777),
    .I1(n776)
  );
  //AND U182bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U182bar (
    .O(n962bar),
    .I0(n777bar),
    .I1(n776bar)
  );
  //OR U183
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U183 (
    .O(n776),
    .I0(n775),
    .I1(n774)
  );
  //AND U183bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U183bar (
    .O(n776bar),
    .I0(n775bar),
    .I1(n774bar)
  );
  //OR U184
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U184 (
    .O(n774),
    .I0(n773),
    .I1(n772)
  );
  //AND U184bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U184bar (
    .O(n774bar),
    .I0(n773bar),
    .I1(n772bar)
  );
  //OR U185
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U185 (
    .O(n772),
    .I0(in[131]),
    .I1(in[120])
  );
  //AND U185bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U185bar (
    .O(n772bar),
    .I0(inbar[131]),
    .I1(inbar[120])
  );
  //OR U186
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U186 (
    .O(n773),
    .I0(in[153]),
    .I1(in[147])
  );
  //AND U186bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U186bar (
    .O(n773bar),
    .I0(inbar[153]),
    .I1(inbar[147])
  );
  //OR U187
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U187 (
    .O(n775),
    .I0(n771),
    .I1(n770)
  );
  //AND U187bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U187bar (
    .O(n775bar),
    .I0(n771bar),
    .I1(n770bar)
  );
  //OR U188
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U188 (
    .O(n770),
    .I0(in[170]),
    .I1(in[156])
  );
  //AND U188bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U188bar (
    .O(n770bar),
    .I0(inbar[170]),
    .I1(inbar[156])
  );
  //OR U189
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U189 (
    .O(n771),
    .I0(in[223]),
    .I1(in[190])
  );
  //AND U189bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U189bar (
    .O(n771bar),
    .I0(inbar[223]),
    .I1(inbar[190])
  );
  //OR U190
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U190 (
    .O(n777),
    .I0(n769),
    .I1(n768)
  );
  //AND U190bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U190bar (
    .O(n777bar),
    .I0(n769bar),
    .I1(n768bar)
  );
  //OR U191
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U191 (
    .O(n768),
    .I0(n767),
    .I1(n766)
  );
  //AND U191bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U191bar (
    .O(n768bar),
    .I0(n767bar),
    .I1(n766bar)
  );
  //OR U192
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U192 (
    .O(n766),
    .I0(in[236]),
    .I1(in[230])
  );
  //AND U192bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U192bar (
    .O(n766bar),
    .I0(inbar[236]),
    .I1(inbar[230])
  );
  //OR U193
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U193 (
    .O(n767),
    .I0(in[85]),
    .I1(in[240])
  );
  //AND U193bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U193bar (
    .O(n767bar),
    .I0(inbar[85]),
    .I1(inbar[240])
  );
  //OR U194
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U194 (
    .O(n769),
    .I0(n765),
    .I1(n764)
  );
  //AND U194bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U194bar (
    .O(n769bar),
    .I0(n765bar),
    .I1(n764bar)
  );
  //OR U195
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U195 (
    .O(n764),
    .I0(in_12),
    .I1(in[90])
  );
  //AND U195bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U195bar (
    .O(n764bar),
    .I0(in_12bar),
    .I1(inbar[90])
  );
  //OR U196
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U196 (
    .O(n765),
    .I0(in_39),
    .I1(in_28)
  );
  //AND U196bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U196bar (
    .O(n765bar),
    .I0(in_39bar),
    .I1(in_28bar)
  );
  //OR U197
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U197 (
    .O(n780),
    .I0(in[109]),
    .I1(n763)
  );
  //AND U197bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U197bar (
    .O(n780bar),
    .I0(inbar[109]),
    .I1(n763bar)
  );
  //OR U198
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U198 (
    .O(n782),
    .I0(n762),
    .I1(n761)
  );
  //AND U198bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U198bar (
    .O(n782bar),
    .I0(n762bar),
    .I1(n761bar)
  );
  //OR U199
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U199 (
    .O(n761),
    .I0(in[138]),
    .I1(in[129])
  );
  //AND U199bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U199bar (
    .O(n761bar),
    .I0(inbar[138]),
    .I1(inbar[129])
  );
  //OR U200
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U200 (
    .O(n762),
    .I0(in[157]),
    .I1(n760)
  );
  //AND U200bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U200bar (
    .O(n762bar),
    .I0(inbar[157]),
    .I1(n760bar)
  );
  //OR U201
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U201 (
    .O(n760),
    .I0(in[182]),
    .I1(in[167])
  );
  //AND U201bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U201bar (
    .O(n760bar),
    .I0(inbar[182]),
    .I1(inbar[167])
  );
  //OR U202
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U202 (
    .O(n784),
    .I0(n759),
    .I1(n758)
  );
  //AND U202bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U202bar (
    .O(n784bar),
    .I0(n759bar),
    .I1(n758bar)
  );
  //OR U203
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U203 (
    .O(n758),
    .I0(n757),
    .I1(n756)
  );
  //AND U203bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U203bar (
    .O(n758bar),
    .I0(n757bar),
    .I1(n756bar)
  );
  //OR U204
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U204 (
    .O(n756),
    .I0(in[195]),
    .I1(in[184])
  );
  //AND U204bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U204bar (
    .O(n756bar),
    .I0(inbar[195]),
    .I1(inbar[184])
  );
  //OR U205
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U205 (
    .O(n757),
    .I0(in[196]),
    .I1(n755)
  );
  //AND U205bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U205bar (
    .O(n757bar),
    .I0(inbar[196]),
    .I1(n755bar)
  );
  //OR U206
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U206 (
    .O(n755),
    .I0(in[215]),
    .I1(in[209])
  );
  //AND U206bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U206bar (
    .O(n755bar),
    .I0(inbar[215]),
    .I1(inbar[209])
  );
  //OR U207
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U207 (
    .O(n759),
    .I0(n754),
    .I1(n753)
  );
  //AND U207bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U207bar (
    .O(n759bar),
    .I0(n754bar),
    .I1(n753bar)
  );
  //OR U208
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U208 (
    .O(n753),
    .I0(in[93]),
    .I1(in[233])
  );
  //AND U208bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U208bar (
    .O(n753bar),
    .I0(inbar[93]),
    .I1(inbar[233])
  );
  //OR U209
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U209 (
    .O(n754),
    .I0(in_1),
    .I1(n752)
  );
  //AND U209bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U209bar (
    .O(n754bar),
    .I0(in_1bar),
    .I1(n752bar)
  );
  //OR U210
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U210 (
    .O(n752),
    .I0(in_69),
    .I1(in_66)
  );
  //AND U210bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U210bar (
    .O(n752bar),
    .I0(in_69bar),
    .I1(in_66bar)
  );
  //OR U211
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U211 (
    .O(n787),
    .I0(n966),
    .I1(n751)
  );
  //AND U211bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U211bar (
    .O(n787bar),
    .I0(n966bar),
    .I1(n751bar)
  );
  //OR U212
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U212 (
    .O(n751),
    .I0(in[134]),
    .I1(n750)
  );
  //AND U212bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U212bar (
    .O(n751bar),
    .I0(inbar[134]),
    .I1(n750bar)
  );
  //OR U213
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U213 (
    .O(n966),
    .I0(n749),
    .I1(n748)
  );
  //AND U213bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U213bar (
    .O(n966bar),
    .I0(n749bar),
    .I1(n748bar)
  );
  //OR U214
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U214 (
    .O(n748),
    .I0(n747),
    .I1(n746)
  );
  //AND U214bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U214bar (
    .O(n748bar),
    .I0(n747bar),
    .I1(n746bar)
  );
  //OR U215
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U215 (
    .O(n746),
    .I0(n745),
    .I1(n744)
  );
  //AND U215bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U215bar (
    .O(n746bar),
    .I0(n745bar),
    .I1(n744bar)
  );
  //OR U216
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U216 (
    .O(n744),
    .I0(in[136]),
    .I1(in[121])
  );
  //AND U216bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U216bar (
    .O(n744bar),
    .I0(inbar[136]),
    .I1(inbar[121])
  );
  //OR U217
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U217 (
    .O(n745),
    .I0(in[186]),
    .I1(in[174])
  );
  //AND U217bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U217bar (
    .O(n745bar),
    .I0(inbar[186]),
    .I1(inbar[174])
  );
  //OR U218
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U218 (
    .O(n747),
    .I0(n743),
    .I1(n742)
  );
  //AND U218bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U218bar (
    .O(n747bar),
    .I0(n743bar),
    .I1(n742bar)
  );
  //OR U219
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U219 (
    .O(n742),
    .I0(in[198]),
    .I1(in[197])
  );
  //AND U219bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U219bar (
    .O(n742bar),
    .I0(inbar[198]),
    .I1(inbar[197])
  );
  //OR U220
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U220 (
    .O(n743),
    .I0(in[214]),
    .I1(in[199])
  );
  //AND U220bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U220bar (
    .O(n743bar),
    .I0(inbar[214]),
    .I1(inbar[199])
  );
  //OR U221
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U221 (
    .O(n749),
    .I0(n741),
    .I1(n740)
  );
  //AND U221bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U221bar (
    .O(n749bar),
    .I0(n741bar),
    .I1(n740bar)
  );
  //OR U222
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U222 (
    .O(n740),
    .I0(n739),
    .I1(n738)
  );
  //AND U222bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U222bar (
    .O(n740bar),
    .I0(n739bar),
    .I1(n738bar)
  );
  //OR U223
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U223 (
    .O(n738),
    .I0(in[231]),
    .I1(in[220])
  );
  //AND U223bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U223bar (
    .O(n738bar),
    .I0(inbar[231]),
    .I1(inbar[220])
  );
  //OR U224
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U224 (
    .O(n739),
    .I0(in_25),
    .I1(in[245])
  );
  //AND U224bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U224bar (
    .O(n739bar),
    .I0(in_25bar),
    .I1(inbar[245])
  );
  //OR U225
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U225 (
    .O(n741),
    .I0(n737),
    .I1(n736)
  );
  //AND U225bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U225bar (
    .O(n741bar),
    .I0(n737bar),
    .I1(n736bar)
  );
  //OR U226
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U226 (
    .O(n736),
    .I0(in_53),
    .I1(in_29)
  );
  //AND U226bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U226bar (
    .O(n736bar),
    .I0(in_53bar),
    .I1(in_29bar)
  );
  //OR U227
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U227 (
    .O(n737),
    .I0(in_79),
    .I1(in_74)
  );
  //AND U227bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U227bar (
    .O(n737bar),
    .I0(in_79bar),
    .I1(in_74bar)
  );
  //OR U228
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U228 (
    .O(n789),
    .I0(n735),
    .I1(n734)
  );
  //AND U228bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U228bar (
    .O(n789bar),
    .I0(n735bar),
    .I1(n734bar)
  );
  //OR U229
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U229 (
    .O(n734),
    .I0(in[152]),
    .I1(in[140])
  );
  //AND U229bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U229bar (
    .O(n734bar),
    .I0(inbar[152]),
    .I1(inbar[140])
  );
  //OR U230
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U230 (
    .O(n735),
    .I0(in[155]),
    .I1(n733)
  );
  //AND U230bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U230bar (
    .O(n735bar),
    .I0(inbar[155]),
    .I1(n733bar)
  );
  //OR U231
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U231 (
    .O(n733),
    .I0(in[166]),
    .I1(in[165])
  );
  //AND U231bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U231bar (
    .O(n733bar),
    .I0(inbar[166]),
    .I1(inbar[165])
  );
  //OR U232
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U232 (
    .O(n791),
    .I0(n732),
    .I1(n731)
  );
  //AND U232bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U232bar (
    .O(n791bar),
    .I0(n732bar),
    .I1(n731bar)
  );
  //OR U233
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U233 (
    .O(n731),
    .I0(n730),
    .I1(n729)
  );
  //AND U233bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U233bar (
    .O(n731bar),
    .I0(n730bar),
    .I1(n729bar)
  );
  //OR U234
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U234 (
    .O(n729),
    .I0(in[202]),
    .I1(in[185])
  );
  //AND U234bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U234bar (
    .O(n729bar),
    .I0(inbar[202]),
    .I1(inbar[185])
  );
  //OR U235
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U235 (
    .O(n730),
    .I0(in[211]),
    .I1(n728)
  );
  //AND U235bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U235bar (
    .O(n730bar),
    .I0(inbar[211]),
    .I1(n728bar)
  );
  //OR U236
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U236 (
    .O(n728),
    .I0(in[255]),
    .I1(in[253])
  );
  //AND U236bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U236bar (
    .O(n728bar),
    .I0(inbar[255]),
    .I1(inbar[253])
  );
  //OR U237
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U237 (
    .O(n732),
    .I0(n727),
    .I1(n726)
  );
  //AND U237bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U237bar (
    .O(n732bar),
    .I0(n727bar),
    .I1(n726bar)
  );
  //OR U238
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U238 (
    .O(n726),
    .I0(in_35),
    .I1(in_15)
  );
  //AND U238bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U238bar (
    .O(n726bar),
    .I0(in_35bar),
    .I1(in_15bar)
  );
  //OR U239
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U239 (
    .O(n727),
    .I0(in_36),
    .I1(n725)
  );
  //AND U239bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U239bar (
    .O(n727bar),
    .I0(in_36bar),
    .I1(n725bar)
  );
  //OR U240
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U240 (
    .O(n725),
    .I0(in_48),
    .I1(in_40)
  );
  //AND U240bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U240bar (
    .O(n725bar),
    .I0(in_48bar),
    .I1(in_40bar)
  );
  //OR U241
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U241 (
    .O(out[1]),
    .I0(n724),
    .I1(n723)
  );
  //AND U241bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U241bar (
    .O(outbar[1]),
    .I0(n724bar),
    .I1(n723bar)
  );
  //OR U242
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U242 (
    .O(n723),
    .I0(n722),
    .I1(n721)
  );
  //AND U242bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U242bar (
    .O(n723bar),
    .I0(n722bar),
    .I1(n721bar)
  );
  //OR U243
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U243 (
    .O(n721),
    .I0(n720),
    .I1(n719)
  );
  //AND U243bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U243bar (
    .O(n721bar),
    .I0(n720bar),
    .I1(n719bar)
  );
  //OR U244
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U244 (
    .O(n719),
    .I0(n921),
    .I1(n887)
  );
  //AND U244bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U244bar (
    .O(n719bar),
    .I0(n921bar),
    .I1(n887bar)
  );
  //OR U245
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U245 (
    .O(n887),
    .I0(n718),
    .I1(n717)
  );
  //AND U245bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U245bar (
    .O(n887bar),
    .I0(n718bar),
    .I1(n717bar)
  );
  //OR U246
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U246 (
    .O(n717),
    .I0(n716),
    .I1(n715)
  );
  //AND U246bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U246bar (
    .O(n717bar),
    .I0(n716bar),
    .I1(n715bar)
  );
  //OR U247
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U247 (
    .O(n715),
    .I0(n714),
    .I1(n713)
  );
  //AND U247bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U247bar (
    .O(n715bar),
    .I0(n714bar),
    .I1(n713bar)
  );
  //OR U248
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U248 (
    .O(n713),
    .I0(in[116]),
    .I1(in[110])
  );
  //AND U248bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U248bar (
    .O(n713bar),
    .I0(inbar[116]),
    .I1(inbar[110])
  );
  //OR U249
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U249 (
    .O(n714),
    .I0(in[133]),
    .I1(in[130])
  );
  //AND U249bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U249bar (
    .O(n714bar),
    .I0(inbar[133]),
    .I1(inbar[130])
  );
  //OR U250
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U250 (
    .O(n716),
    .I0(n712),
    .I1(n711)
  );
  //AND U250bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U250bar (
    .O(n716bar),
    .I0(n712bar),
    .I1(n711bar)
  );
  //OR U251
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U251 (
    .O(n711),
    .I0(in[203]),
    .I1(in[135])
  );
  //AND U251bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U251bar (
    .O(n711bar),
    .I0(inbar[203]),
    .I1(inbar[135])
  );
  //OR U252
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U252 (
    .O(n712),
    .I0(in[232]),
    .I1(in[223])
  );
  //AND U252bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U252bar (
    .O(n712bar),
    .I0(inbar[232]),
    .I1(inbar[223])
  );
  //OR U253
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U253 (
    .O(n718),
    .I0(n710),
    .I1(n709)
  );
  //AND U253bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U253bar (
    .O(n718bar),
    .I0(n710bar),
    .I1(n709bar)
  );
  //OR U254
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U254 (
    .O(n709),
    .I0(n708),
    .I1(n707)
  );
  //AND U254bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U254bar (
    .O(n709bar),
    .I0(n708bar),
    .I1(n707bar)
  );
  //OR U255
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U255 (
    .O(n707),
    .I0(in[255]),
    .I1(in[233])
  );
  //AND U255bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U255bar (
    .O(n707bar),
    .I0(inbar[255]),
    .I1(inbar[233])
  );
  //OR U256
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U256 (
    .O(n708),
    .I0(in_53),
    .I1(in_34)
  );
  //AND U256bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U256bar (
    .O(n708bar),
    .I0(in_53bar),
    .I1(in_34bar)
  );
  //OR U257
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U257 (
    .O(n710),
    .I0(n706),
    .I1(n705)
  );
  //AND U257bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U257bar (
    .O(n710bar),
    .I0(n706bar),
    .I1(n705bar)
  );
  //OR U258
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U258 (
    .O(n705),
    .I0(in_57),
    .I1(in_55)
  );
  //AND U258bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U258bar (
    .O(n705bar),
    .I0(in_57bar),
    .I1(in_55bar)
  );
  //OR U259
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U259 (
    .O(n706),
    .I0(in_68),
    .I1(in_67)
  );
  //AND U259bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U259bar (
    .O(n706bar),
    .I0(in_68bar),
    .I1(in_67bar)
  );
  //OR U260
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U260 (
    .O(n921),
    .I0(n704),
    .I1(n703)
  );
  //AND U260bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U260bar (
    .O(n921bar),
    .I0(n704bar),
    .I1(n703bar)
  );
  //OR U261
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U261 (
    .O(n703),
    .I0(n702),
    .I1(n701)
  );
  //AND U261bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U261bar (
    .O(n703bar),
    .I0(n702bar),
    .I1(n701bar)
  );
  //OR U262
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U262 (
    .O(n701),
    .I0(n700),
    .I1(n699)
  );
  //AND U262bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U262bar (
    .O(n701bar),
    .I0(n700bar),
    .I1(n699bar)
  );
  //OR U263
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U263 (
    .O(n699),
    .I0(n944),
    .I1(n872)
  );
  //AND U263bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U263bar (
    .O(n699bar),
    .I0(n944bar),
    .I1(n872bar)
  );
  //OR U264
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U264 (
    .O(n872),
    .I0(n698),
    .I1(n697)
  );
  //AND U264bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U264bar (
    .O(n872bar),
    .I0(n698bar),
    .I1(n697bar)
  );
  //OR U265
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U265 (
    .O(n697),
    .I0(n696),
    .I1(n695)
  );
  //AND U265bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U265bar (
    .O(n697bar),
    .I0(n696bar),
    .I1(n695bar)
  );
  //OR U266
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U266 (
    .O(n695),
    .I0(n694),
    .I1(n693)
  );
  //AND U266bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U266bar (
    .O(n695bar),
    .I0(n694bar),
    .I1(n693bar)
  );
  //OR U267
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U267 (
    .O(n693),
    .I0(in[121]),
    .I1(in[102])
  );
  //AND U267bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U267bar (
    .O(n693bar),
    .I0(inbar[121]),
    .I1(inbar[102])
  );
  //OR U268
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U268 (
    .O(n694),
    .I0(in[162]),
    .I1(in[161])
  );
  //AND U268bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U268bar (
    .O(n694bar),
    .I0(inbar[162]),
    .I1(inbar[161])
  );
  //OR U269
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U269 (
    .O(n696),
    .I0(n692),
    .I1(n691)
  );
  //AND U269bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U269bar (
    .O(n696bar),
    .I0(n692bar),
    .I1(n691bar)
  );
  //OR U270
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U270 (
    .O(n691),
    .I0(in[192]),
    .I1(in[178])
  );
  //AND U270bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U270bar (
    .O(n691bar),
    .I0(inbar[192]),
    .I1(inbar[178])
  );
  //OR U271
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U271 (
    .O(n692),
    .I0(in[244]),
    .I1(in[209])
  );
  //AND U271bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U271bar (
    .O(n692bar),
    .I0(inbar[244]),
    .I1(inbar[209])
  );
  //OR U272
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U272 (
    .O(n698),
    .I0(n690),
    .I1(n689)
  );
  //AND U272bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U272bar (
    .O(n698bar),
    .I0(n690bar),
    .I1(n689bar)
  );
  //OR U273
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U273 (
    .O(n689),
    .I0(n688),
    .I1(n687)
  );
  //AND U273bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U273bar (
    .O(n689bar),
    .I0(n688bar),
    .I1(n687bar)
  );
  //OR U274
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U274 (
    .O(n687),
    .I0(in[90]),
    .I1(in[254])
  );
  //AND U274bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U274bar (
    .O(n687bar),
    .I0(inbar[90]),
    .I1(inbar[254])
  );
  //OR U275
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U275 (
    .O(n688),
    .I0(in_36),
    .I1(in_32)
  );
  //AND U275bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U275bar (
    .O(n688bar),
    .I0(in_36bar),
    .I1(in_32bar)
  );
  //OR U276
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U276 (
    .O(n690),
    .I0(n686),
    .I1(n685)
  );
  //AND U276bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U276bar (
    .O(n690bar),
    .I0(n686bar),
    .I1(n685bar)
  );
  //OR U277
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U277 (
    .O(n685),
    .I0(in_62),
    .I1(in_37)
  );
  //AND U277bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U277bar (
    .O(n685bar),
    .I0(in_62bar),
    .I1(in_37bar)
  );
  //OR U278
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U278 (
    .O(n686),
    .I0(in_75),
    .I1(in_73)
  );
  //AND U278bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U278bar (
    .O(n686bar),
    .I0(in_75bar),
    .I1(in_73bar)
  );
  //OR U279
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U279 (
    .O(n944),
    .I0(n684),
    .I1(n683)
  );
  //AND U279bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U279bar (
    .O(n944bar),
    .I0(n684bar),
    .I1(n683bar)
  );
  //OR U280
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U280 (
    .O(n683),
    .I0(n682),
    .I1(n681)
  );
  //AND U280bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U280bar (
    .O(n683bar),
    .I0(n682bar),
    .I1(n681bar)
  );
  //OR U281
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U281 (
    .O(n681),
    .I0(n680),
    .I1(n679)
  );
  //AND U281bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U281bar (
    .O(n681bar),
    .I0(n680bar),
    .I1(n679bar)
  );
  //OR U282
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U282 (
    .O(n679),
    .I0(in[171]),
    .I1(in[153])
  );
  //AND U282bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U282bar (
    .O(n679bar),
    .I0(inbar[171]),
    .I1(inbar[153])
  );
  //OR U283
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U283 (
    .O(n680),
    .I0(in[187]),
    .I1(in[176])
  );
  //AND U283bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U283bar (
    .O(n680bar),
    .I0(inbar[187]),
    .I1(inbar[176])
  );
  //OR U284
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U284 (
    .O(n682),
    .I0(n678),
    .I1(n677)
  );
  //AND U284bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U284bar (
    .O(n682bar),
    .I0(n678bar),
    .I1(n677bar)
  );
  //OR U285
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U285 (
    .O(n677),
    .I0(in[245]),
    .I1(in[211])
  );
  //AND U285bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U285bar (
    .O(n677bar),
    .I0(inbar[245]),
    .I1(inbar[211])
  );
  //OR U286
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U286 (
    .O(n678),
    .I0(in[97]),
    .I1(in[88])
  );
  //AND U286bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U286bar (
    .O(n678bar),
    .I0(inbar[97]),
    .I1(inbar[88])
  );
  //OR U287
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U287 (
    .O(n684),
    .I0(n676),
    .I1(n675)
  );
  //AND U287bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U287bar (
    .O(n684bar),
    .I0(n676bar),
    .I1(n675bar)
  );
  //OR U288
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U288 (
    .O(n675),
    .I0(n674),
    .I1(n673)
  );
  //AND U288bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U288bar (
    .O(n675bar),
    .I0(n674bar),
    .I1(n673bar)
  );
  //OR U289
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U289 (
    .O(n673),
    .I0(in_10),
    .I1(in_0)
  );
  //AND U289bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U289bar (
    .O(n673bar),
    .I0(in_10bar),
    .I1(in_0bar)
  );
  //OR U290
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U290 (
    .O(n674),
    .I0(in_59),
    .I1(in_5)
  );
  //AND U290bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U290bar (
    .O(n674bar),
    .I0(in_59bar),
    .I1(in_5bar)
  );
  //OR U291
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U291 (
    .O(n676),
    .I0(n672),
    .I1(n671)
  );
  //AND U291bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U291bar (
    .O(n676bar),
    .I0(n672bar),
    .I1(n671bar)
  );
  //OR U292
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U292 (
    .O(n671),
    .I0(in_60),
    .I1(in_6)
  );
  //AND U292bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U292bar (
    .O(n671bar),
    .I0(in_60bar),
    .I1(in_6bar)
  );
  //OR U293
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U293 (
    .O(n672),
    .I0(in_77),
    .I1(in_69)
  );
  //AND U293bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U293bar (
    .O(n672bar),
    .I0(in_77bar),
    .I1(in_69bar)
  );
  //OR U294
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U294 (
    .O(n700),
    .I0(in[113]),
    .I1(n864)
  );
  //AND U294bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U294bar (
    .O(n700bar),
    .I0(inbar[113]),
    .I1(n864bar)
  );
  //OR U295
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U295 (
    .O(n864),
    .I0(n670),
    .I1(n669)
  );
  //AND U295bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U295bar (
    .O(n864bar),
    .I0(n670bar),
    .I1(n669bar)
  );
  //OR U296
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U296 (
    .O(n669),
    .I0(n668),
    .I1(n667)
  );
  //AND U296bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U296bar (
    .O(n669bar),
    .I0(n668bar),
    .I1(n667bar)
  );
  //OR U297
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U297 (
    .O(n667),
    .I0(n666),
    .I1(n665)
  );
  //AND U297bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U297bar (
    .O(n667bar),
    .I0(n666bar),
    .I1(n665bar)
  );
  //OR U298
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U298 (
    .O(n665),
    .I0(in[125]),
    .I1(in[107])
  );
  //AND U298bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U298bar (
    .O(n665bar),
    .I0(inbar[125]),
    .I1(inbar[107])
  );
  //OR U299
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U299 (
    .O(n666),
    .I0(in[138]),
    .I1(in[126])
  );
  //AND U299bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U299bar (
    .O(n666bar),
    .I0(inbar[138]),
    .I1(inbar[126])
  );
  //OR U300
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U300 (
    .O(n668),
    .I0(n664),
    .I1(n663)
  );
  //AND U300bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U300bar (
    .O(n668bar),
    .I0(n664bar),
    .I1(n663bar)
  );
  //OR U301
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U301 (
    .O(n663),
    .I0(in[189]),
    .I1(in[143])
  );
  //AND U301bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U301bar (
    .O(n663bar),
    .I0(inbar[189]),
    .I1(inbar[143])
  );
  //OR U302
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U302 (
    .O(n664),
    .I0(in[99]),
    .I1(in[214])
  );
  //AND U302bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U302bar (
    .O(n664bar),
    .I0(inbar[99]),
    .I1(inbar[214])
  );
  //OR U303
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U303 (
    .O(n670),
    .I0(n662),
    .I1(n661)
  );
  //AND U303bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U303bar (
    .O(n670bar),
    .I0(n662bar),
    .I1(n661bar)
  );
  //OR U304
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U304 (
    .O(n661),
    .I0(n660),
    .I1(n659)
  );
  //AND U304bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U304bar (
    .O(n661bar),
    .I0(n660bar),
    .I1(n659bar)
  );
  //OR U305
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U305 (
    .O(n659),
    .I0(in_15),
    .I1(in_12)
  );
  //AND U305bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U305bar (
    .O(n659bar),
    .I0(in_15bar),
    .I1(in_12bar)
  );
  //OR U306
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U306 (
    .O(n660),
    .I0(in_20),
    .I1(in_2)
  );
  //AND U306bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U306bar (
    .O(n660bar),
    .I0(in_20bar),
    .I1(in_2bar)
  );
  //OR U307
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U307 (
    .O(n662),
    .I0(n658),
    .I1(n657)
  );
  //AND U307bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U307bar (
    .O(n662bar),
    .I0(n658bar),
    .I1(n657bar)
  );
  //OR U308
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U308 (
    .O(n657),
    .I0(in_30),
    .I1(in_3)
  );
  //AND U308bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U308bar (
    .O(n657bar),
    .I0(in_30bar),
    .I1(in_3bar)
  );
  //OR U309
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U309 (
    .O(n658),
    .I0(in_4),
    .I1(in_38)
  );
  //AND U309bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U309bar (
    .O(n658bar),
    .I0(in_4bar),
    .I1(in_38bar)
  );
  //OR U310
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U310 (
    .O(n702),
    .I0(n656),
    .I1(n655)
  );
  //AND U310bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U310bar (
    .O(n702bar),
    .I0(n656bar),
    .I1(n655bar)
  );
  //OR U311
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U311 (
    .O(n655),
    .I0(in[148]),
    .I1(in[137])
  );
  //AND U311bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U311bar (
    .O(n655bar),
    .I0(inbar[148]),
    .I1(inbar[137])
  );
  //OR U312
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U312 (
    .O(n656),
    .I0(in[149]),
    .I1(n654)
  );
  //AND U312bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U312bar (
    .O(n656bar),
    .I0(inbar[149]),
    .I1(n654bar)
  );
  //OR U313
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U313 (
    .O(n654),
    .I0(in[195]),
    .I1(in[190])
  );
  //AND U313bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U313bar (
    .O(n654bar),
    .I0(inbar[195]),
    .I1(inbar[190])
  );
  //OR U314
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U314 (
    .O(n704),
    .I0(n653),
    .I1(n652)
  );
  //AND U314bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U314bar (
    .O(n704bar),
    .I0(n653bar),
    .I1(n652bar)
  );
  //OR U315
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U315 (
    .O(n652),
    .I0(n651),
    .I1(n650)
  );
  //AND U315bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U315bar (
    .O(n652bar),
    .I0(n651bar),
    .I1(n650bar)
  );
  //OR U316
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U316 (
    .O(n650),
    .I0(in[98]),
    .I1(in[197])
  );
  //AND U316bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U316bar (
    .O(n650bar),
    .I0(inbar[98]),
    .I1(inbar[197])
  );
  //OR U317
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U317 (
    .O(n651),
    .I0(in_11),
    .I1(n649)
  );
  //AND U317bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U317bar (
    .O(n651bar),
    .I0(in_11bar),
    .I1(n649bar)
  );
  //OR U318
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U318 (
    .O(n649),
    .I0(in_26),
    .I1(in_14)
  );
  //AND U318bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U318bar (
    .O(n649bar),
    .I0(in_26bar),
    .I1(in_14bar)
  );
  //OR U319
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U319 (
    .O(n653),
    .I0(n648),
    .I1(n647)
  );
  //AND U319bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U319bar (
    .O(n653bar),
    .I0(n648bar),
    .I1(n647bar)
  );
  //OR U320
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U320 (
    .O(n647),
    .I0(in_35),
    .I1(in_27)
  );
  //AND U320bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U320bar (
    .O(n647bar),
    .I0(in_35bar),
    .I1(in_27bar)
  );
  //OR U321
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U321 (
    .O(n648),
    .I0(in_50),
    .I1(n646)
  );
  //AND U321bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U321bar (
    .O(n648bar),
    .I0(in_50bar),
    .I1(n646bar)
  );
  //OR U322
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U322 (
    .O(n646),
    .I0(in_78),
    .I1(in_61)
  );
  //AND U322bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U322bar (
    .O(n646bar),
    .I0(in_78bar),
    .I1(in_61bar)
  );
  //OR U323
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U323 (
    .O(n720),
    .I0(n942),
    .I1(n645)
  );
  //AND U323bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U323bar (
    .O(n720bar),
    .I0(n942bar),
    .I1(n645bar)
  );
  //OR U324
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U324 (
    .O(n645),
    .I0(in[106]),
    .I1(n863)
  );
  //AND U324bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U324bar (
    .O(n645bar),
    .I0(inbar[106]),
    .I1(n863bar)
  );
  //OR U325
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U325 (
    .O(n863),
    .I0(n644),
    .I1(n643)
  );
  //AND U325bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U325bar (
    .O(n863bar),
    .I0(n644bar),
    .I1(n643bar)
  );
  //OR U326
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U326 (
    .O(n643),
    .I0(n642),
    .I1(n641)
  );
  //AND U326bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U326bar (
    .O(n643bar),
    .I0(n642bar),
    .I1(n641bar)
  );
  //OR U327
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U327 (
    .O(n641),
    .I0(n640),
    .I1(n639)
  );
  //AND U327bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U327bar (
    .O(n641bar),
    .I0(n640bar),
    .I1(n639bar)
  );
  //OR U328
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U328 (
    .O(n639),
    .I0(in[127]),
    .I1(in[122])
  );
  //AND U328bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U328bar (
    .O(n639bar),
    .I0(inbar[127]),
    .I1(inbar[122])
  );
  //OR U329
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U329 (
    .O(n640),
    .I0(in[156]),
    .I1(in[132])
  );
  //AND U329bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U329bar (
    .O(n640bar),
    .I0(inbar[156]),
    .I1(inbar[132])
  );
  //OR U330
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U330 (
    .O(n642),
    .I0(n638),
    .I1(n637)
  );
  //AND U330bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U330bar (
    .O(n642bar),
    .I0(n638bar),
    .I1(n637bar)
  );
  //OR U331
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U331 (
    .O(n637),
    .I0(in[159]),
    .I1(in[157])
  );
  //AND U331bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U331bar (
    .O(n637bar),
    .I0(inbar[159]),
    .I1(inbar[157])
  );
  //OR U332
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U332 (
    .O(n638),
    .I0(in[185]),
    .I1(in[169])
  );
  //AND U332bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U332bar (
    .O(n638bar),
    .I0(inbar[185]),
    .I1(inbar[169])
  );
  //OR U333
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U333 (
    .O(n644),
    .I0(n636),
    .I1(n635)
  );
  //AND U333bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U333bar (
    .O(n644bar),
    .I0(n636bar),
    .I1(n635bar)
  );
  //OR U334
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U334 (
    .O(n635),
    .I0(n634),
    .I1(n633)
  );
  //AND U334bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U334bar (
    .O(n635bar),
    .I0(n634bar),
    .I1(n633bar)
  );
  //OR U335
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U335 (
    .O(n633),
    .I0(in[239]),
    .I1(in[218])
  );
  //AND U335bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U335bar (
    .O(n633bar),
    .I0(inbar[239]),
    .I1(inbar[218])
  );
  //OR U336
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U336 (
    .O(n634),
    .I0(in_13),
    .I1(in[87])
  );
  //AND U336bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U336bar (
    .O(n634bar),
    .I0(in_13bar),
    .I1(inbar[87])
  );
  //OR U337
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U337 (
    .O(n636),
    .I0(n632),
    .I1(n631)
  );
  //AND U337bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U337bar (
    .O(n636bar),
    .I0(n632bar),
    .I1(n631bar)
  );
  //OR U338
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U338 (
    .O(n631),
    .I0(in_72),
    .I1(in_70)
  );
  //AND U338bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U338bar (
    .O(n631bar),
    .I0(in_72bar),
    .I1(in_70bar)
  );
  //OR U339
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U339 (
    .O(n632),
    .I0(in_80),
    .I1(in_74)
  );
  //AND U339bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U339bar (
    .O(n632bar),
    .I0(in_80bar),
    .I1(in_74bar)
  );
  //OR U340
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U340 (
    .O(n942),
    .I0(n630),
    .I1(n629)
  );
  //AND U340bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U340bar (
    .O(n942bar),
    .I0(n630bar),
    .I1(n629bar)
  );
  //OR U341
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U341 (
    .O(n629),
    .I0(n628),
    .I1(n627)
  );
  //AND U341bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U341bar (
    .O(n629bar),
    .I0(n628bar),
    .I1(n627bar)
  );
  //OR U342
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U342 (
    .O(n627),
    .I0(n626),
    .I1(n625)
  );
  //AND U342bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U342bar (
    .O(n627bar),
    .I0(n626bar),
    .I1(n625bar)
  );
  //OR U343
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U343 (
    .O(n625),
    .I0(in[146]),
    .I1(in[100])
  );
  //AND U343bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U343bar (
    .O(n625bar),
    .I0(inbar[146]),
    .I1(inbar[100])
  );
  //OR U344
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U344 (
    .O(n626),
    .I0(in[168]),
    .I1(in[152])
  );
  //AND U344bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U344bar (
    .O(n626bar),
    .I0(inbar[168]),
    .I1(inbar[152])
  );
  //OR U345
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U345 (
    .O(n628),
    .I0(n624),
    .I1(n623)
  );
  //AND U345bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U345bar (
    .O(n628bar),
    .I0(n624bar),
    .I1(n623bar)
  );
  //OR U346
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U346 (
    .O(n623),
    .I0(in[199]),
    .I1(in[182])
  );
  //AND U346bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U346bar (
    .O(n623bar),
    .I0(inbar[199]),
    .I1(inbar[182])
  );
  //OR U347
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U347 (
    .O(n624),
    .I0(in[236]),
    .I1(in[204])
  );
  //AND U347bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U347bar (
    .O(n624bar),
    .I0(inbar[236]),
    .I1(inbar[204])
  );
  //OR U348
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U348 (
    .O(n630),
    .I0(n622),
    .I1(n621)
  );
  //AND U348bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U348bar (
    .O(n630bar),
    .I0(n622bar),
    .I1(n621bar)
  );
  //OR U349
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U349 (
    .O(n621),
    .I0(n620),
    .I1(n619)
  );
  //AND U349bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U349bar (
    .O(n621bar),
    .I0(n620bar),
    .I1(n619bar)
  );
  //OR U350
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U350 (
    .O(n619),
    .I0(in[89]),
    .I1(in[246])
  );
  //AND U350bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U350bar (
    .O(n619bar),
    .I0(inbar[89]),
    .I1(inbar[246])
  );
  //OR U351
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U351 (
    .O(n620),
    .I0(in[95]),
    .I1(in[92])
  );
  //AND U351bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U351bar (
    .O(n620bar),
    .I0(inbar[95]),
    .I1(inbar[92])
  );
  //OR U352
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U352 (
    .O(n622),
    .I0(n618),
    .I1(n617)
  );
  //AND U352bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U352bar (
    .O(n622bar),
    .I0(n618bar),
    .I1(n617bar)
  );
  //OR U353
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U353 (
    .O(n617),
    .I0(in_22),
    .I1(in_16)
  );
  //AND U353bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U353bar (
    .O(n617bar),
    .I0(in_22bar),
    .I1(in_16bar)
  );
  //OR U354
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U354 (
    .O(n618),
    .I0(in_51),
    .I1(in_49)
  );
  //AND U354bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U354bar (
    .O(n618bar),
    .I0(in_51bar),
    .I1(in_49bar)
  );
  //OR U355
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U355 (
    .O(n722),
    .I0(n616),
    .I1(n615)
  );
  //AND U355bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U355bar (
    .O(n722bar),
    .I0(n616bar),
    .I1(n615bar)
  );
  //OR U356
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U356 (
    .O(n615),
    .I0(in[158]),
    .I1(in[115])
  );
  //AND U356bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U356bar (
    .O(n615bar),
    .I0(inbar[158]),
    .I1(inbar[115])
  );
  //OR U357
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U357 (
    .O(n616),
    .I0(in[163]),
    .I1(n614)
  );
  //AND U357bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U357bar (
    .O(n616bar),
    .I0(inbar[163]),
    .I1(n614bar)
  );
  //OR U358
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U358 (
    .O(n614),
    .I0(in[206]),
    .I1(in[165])
  );
  //AND U358bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U358bar (
    .O(n614bar),
    .I0(inbar[206]),
    .I1(inbar[165])
  );
  //OR U359
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U359 (
    .O(n724),
    .I0(n613),
    .I1(n612)
  );
  //AND U359bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U359bar (
    .O(n724bar),
    .I0(n613bar),
    .I1(n612bar)
  );
  //OR U360
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U360 (
    .O(n612),
    .I0(n611),
    .I1(n610)
  );
  //AND U360bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U360bar (
    .O(n612bar),
    .I0(n611bar),
    .I1(n610bar)
  );
  //OR U361
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U361 (
    .O(n610),
    .I0(in[213]),
    .I1(in[207])
  );
  //AND U361bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U361bar (
    .O(n610bar),
    .I0(inbar[213]),
    .I1(inbar[207])
  );
  //OR U362
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U362 (
    .O(n611),
    .I0(in[215]),
    .I1(n609)
  );
  //AND U362bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U362bar (
    .O(n611bar),
    .I0(inbar[215]),
    .I1(n609bar)
  );
  //OR U363
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U363 (
    .O(n609),
    .I0(in[230]),
    .I1(in[220])
  );
  //AND U363bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U363bar (
    .O(n609bar),
    .I0(inbar[230]),
    .I1(inbar[220])
  );
  //OR U364
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U364 (
    .O(n613),
    .I0(n608),
    .I1(n607)
  );
  //AND U364bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U364bar (
    .O(n613bar),
    .I0(n608bar),
    .I1(n607bar)
  );
  //OR U365
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U365 (
    .O(n607),
    .I0(in[251]),
    .I1(in[234])
  );
  //AND U365bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U365bar (
    .O(n607bar),
    .I0(inbar[251]),
    .I1(inbar[234])
  );
  //OR U366
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U366 (
    .O(n608),
    .I0(in_17),
    .I1(n606)
  );
  //AND U366bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U366bar (
    .O(n608bar),
    .I0(in_17bar),
    .I1(n606bar)
  );
  //OR U367
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U367 (
    .O(n606),
    .I0(in_65),
    .I1(in_56)
  );
  //AND U367bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U367bar (
    .O(n606bar),
    .I0(in_65bar),
    .I1(in_56bar)
  );
  //OR U368
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U368 (
    .O(out[0]),
    .I0(n605),
    .I1(n604)
  );
  //AND U368bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U368bar (
    .O(outbar[0]),
    .I0(n605bar),
    .I1(n604bar)
  );
  //OR U369
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U369 (
    .O(n604),
    .I0(n603),
    .I1(n602)
  );
  //AND U369bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U369bar (
    .O(n604bar),
    .I0(n603bar),
    .I1(n602bar)
  );
  //OR U370
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U370 (
    .O(n602),
    .I0(n601),
    .I1(n600)
  );
  //AND U370bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U370bar (
    .O(n602bar),
    .I0(n601bar),
    .I1(n600bar)
  );
  //OR U371
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U371 (
    .O(n600),
    .I0(n820),
    .I1(n785)
  );
  //AND U371bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U371bar (
    .O(n600bar),
    .I0(n820bar),
    .I1(n785bar)
  );
  //OR U372
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U372 (
    .O(n785),
    .I0(n599),
    .I1(n598)
  );
  //AND U372bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U372bar (
    .O(n785bar),
    .I0(n599bar),
    .I1(n598bar)
  );
  //OR U373
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U373 (
    .O(n598),
    .I0(n597),
    .I1(n596)
  );
  //AND U373bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U373bar (
    .O(n598bar),
    .I0(n597bar),
    .I1(n596bar)
  );
  //OR U374
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U374 (
    .O(n596),
    .I0(n595),
    .I1(n594)
  );
  //AND U374bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U374bar (
    .O(n596bar),
    .I0(n595bar),
    .I1(n594bar)
  );
  //OR U375
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U375 (
    .O(n594),
    .I0(in[135]),
    .I1(in[104])
  );
  //AND U375bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U375bar (
    .O(n594bar),
    .I0(inbar[135]),
    .I1(inbar[104])
  );
  //OR U376
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U376 (
    .O(n595),
    .I0(in[188]),
    .I1(in[178])
  );
  //AND U376bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U376bar (
    .O(n595bar),
    .I0(inbar[188]),
    .I1(inbar[178])
  );
  //OR U377
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U377 (
    .O(n597),
    .I0(n593),
    .I1(n592)
  );
  //AND U377bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U377bar (
    .O(n597bar),
    .I0(n593bar),
    .I1(n592bar)
  );
  //OR U378
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U378 (
    .O(n592),
    .I0(in[217]),
    .I1(in[194])
  );
  //AND U378bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U378bar (
    .O(n592bar),
    .I0(inbar[217]),
    .I1(inbar[194])
  );
  //OR U379
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U379 (
    .O(n593),
    .I0(in[237]),
    .I1(in[218])
  );
  //AND U379bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U379bar (
    .O(n593bar),
    .I0(inbar[237]),
    .I1(inbar[218])
  );
  //OR U380
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U380 (
    .O(n599),
    .I0(n591),
    .I1(n590)
  );
  //AND U380bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U380bar (
    .O(n599bar),
    .I0(n591bar),
    .I1(n590bar)
  );
  //OR U381
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U381 (
    .O(n590),
    .I0(n589),
    .I1(n588)
  );
  //AND U381bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U381bar (
    .O(n590bar),
    .I0(n589bar),
    .I1(n588bar)
  );
  //OR U382
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U382 (
    .O(n588),
    .I0(in_2),
    .I1(in_10)
  );
  //AND U382bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U382bar (
    .O(n588bar),
    .I0(in_2bar),
    .I1(in_10bar)
  );
  //OR U383
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U383 (
    .O(n589),
    .I0(in_47),
    .I1(in_22)
  );
  //AND U383bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U383bar (
    .O(n589bar),
    .I0(in_47bar),
    .I1(in_22bar)
  );
  //OR U384
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U384 (
    .O(n591),
    .I0(n587),
    .I1(n586)
  );
  //AND U384bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U384bar (
    .O(n591bar),
    .I0(n587bar),
    .I1(n586bar)
  );
  //OR U385
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U385 (
    .O(n586),
    .I0(in_56),
    .I1(in_54)
  );
  //AND U385bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U385bar (
    .O(n586bar),
    .I0(in_56bar),
    .I1(in_54bar)
  );
  //OR U386
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U386 (
    .O(n587),
    .I0(in_63),
    .I1(in_61)
  );
  //AND U386bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U386bar (
    .O(n587bar),
    .I0(in_63bar),
    .I1(in_61bar)
  );
  //OR U387
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U387 (
    .O(n820),
    .I0(n585),
    .I1(n584)
  );
  //AND U387bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U387bar (
    .O(n820bar),
    .I0(n585bar),
    .I1(n584bar)
  );
  //OR U388
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U388 (
    .O(n584),
    .I0(n583),
    .I1(n582)
  );
  //AND U388bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U388bar (
    .O(n584bar),
    .I0(n583bar),
    .I1(n582bar)
  );
  //OR U389
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U389 (
    .O(n582),
    .I0(n581),
    .I1(n580)
  );
  //AND U389bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U389bar (
    .O(n582bar),
    .I0(n581bar),
    .I1(n580bar)
  );
  //OR U390
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U390 (
    .O(n580),
    .I0(in[158]),
    .I1(in[142])
  );
  //AND U390bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U390bar (
    .O(n580bar),
    .I0(inbar[158]),
    .I1(inbar[142])
  );
  //OR U391
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U391 (
    .O(n581),
    .I0(in[175]),
    .I1(in[164])
  );
  //AND U391bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U391bar (
    .O(n581bar),
    .I0(inbar[175]),
    .I1(inbar[164])
  );
  //OR U392
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U392 (
    .O(n583),
    .I0(n579),
    .I1(n578)
  );
  //AND U392bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U392bar (
    .O(n583bar),
    .I0(n579bar),
    .I1(n578bar)
  );
  //OR U393
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U393 (
    .O(n578),
    .I0(in[228]),
    .I1(in[204])
  );
  //AND U393bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U393bar (
    .O(n578bar),
    .I0(inbar[228]),
    .I1(inbar[204])
  );
  //OR U394
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U394 (
    .O(n579),
    .I0(in[91]),
    .I1(in[87])
  );
  //AND U394bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U394bar (
    .O(n579bar),
    .I0(inbar[91]),
    .I1(inbar[87])
  );
  //OR U395
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U395 (
    .O(n585),
    .I0(n577),
    .I1(n576)
  );
  //AND U395bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U395bar (
    .O(n585bar),
    .I0(n577bar),
    .I1(n576bar)
  );
  //OR U396
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U396 (
    .O(n576),
    .I0(n575),
    .I1(n574)
  );
  //AND U396bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U396bar (
    .O(n576bar),
    .I0(n575bar),
    .I1(n574bar)
  );
  //OR U397
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U397 (
    .O(n574),
    .I0(in_21),
    .I1(in_11)
  );
  //AND U397bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U397bar (
    .O(n574bar),
    .I0(in_21bar),
    .I1(in_11bar)
  );
  //OR U398
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U398 (
    .O(n575),
    .I0(in_5),
    .I1(in_3)
  );
  //AND U398bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U398bar (
    .O(n575bar),
    .I0(in_5bar),
    .I1(in_3bar)
  );
  //OR U399
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U399 (
    .O(n577),
    .I0(n573),
    .I1(n572)
  );
  //AND U399bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U399bar (
    .O(n577bar),
    .I0(n573bar),
    .I1(n572bar)
  );
  //OR U400
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U400 (
    .O(n572),
    .I0(in_68),
    .I1(in_64)
  );
  //AND U400bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U400bar (
    .O(n572bar),
    .I0(in_68bar),
    .I1(in_64bar)
  );
  //OR U401
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U401 (
    .O(n573),
    .I0(in_76),
    .I1(in_73)
  );
  //AND U401bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U401bar (
    .O(n573bar),
    .I0(in_76bar),
    .I1(in_73bar)
  );
  //OR U402
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U402 (
    .O(n601),
    .I0(n778),
    .I1(n571)
  );
  //AND U402bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U402bar (
    .O(n601bar),
    .I0(n778bar),
    .I1(n571bar)
  );
  //OR U403
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U403 (
    .O(n571),
    .I0(in[100]),
    .I1(n965)
  );
  //AND U403bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U403bar (
    .O(n571bar),
    .I0(inbar[100]),
    .I1(n965bar)
  );
  //OR U404
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U404 (
    .O(n965),
    .I0(n570),
    .I1(n569)
  );
  //AND U404bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U404bar (
    .O(n965bar),
    .I0(n570bar),
    .I1(n569bar)
  );
  //OR U405
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U405 (
    .O(n569),
    .I0(n568),
    .I1(n567)
  );
  //AND U405bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U405bar (
    .O(n569bar),
    .I0(n568bar),
    .I1(n567bar)
  );
  //OR U406
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U406 (
    .O(n567),
    .I0(n566),
    .I1(n565)
  );
  //AND U406bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U406bar (
    .O(n567bar),
    .I0(n566bar),
    .I1(n565bar)
  );
  //OR U407
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U407 (
    .O(n565),
    .I0(n817),
    .I1(n750)
  );
  //AND U407bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U407bar (
    .O(n565bar),
    .I0(n817bar),
    .I1(n750bar)
  );
  //OR U408
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U408 (
    .O(n750),
    .I0(n564),
    .I1(n563)
  );
  //AND U408bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U408bar (
    .O(n750bar),
    .I0(n564bar),
    .I1(n563bar)
  );
  //OR U409
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U409 (
    .O(n563),
    .I0(n562),
    .I1(n561)
  );
  //AND U409bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U409bar (
    .O(n563bar),
    .I0(n562bar),
    .I1(n561bar)
  );
  //OR U410
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U410 (
    .O(n561),
    .I0(n560),
    .I1(n559)
  );
  //AND U410bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U410bar (
    .O(n561bar),
    .I0(n560bar),
    .I1(n559bar)
  );
  //OR U411
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U411 (
    .O(n559),
    .I0(in[119]),
    .I1(in[103])
  );
  //AND U411bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U411bar (
    .O(n559bar),
    .I0(inbar[119]),
    .I1(inbar[103])
  );
  //OR U412
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U412 (
    .O(n560),
    .I0(in[137]),
    .I1(in[133])
  );
  //AND U412bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U412bar (
    .O(n560bar),
    .I0(inbar[137]),
    .I1(inbar[133])
  );
  //OR U413
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U413 (
    .O(n562),
    .I0(n558),
    .I1(n557)
  );
  //AND U413bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U413bar (
    .O(n562bar),
    .I0(n558bar),
    .I1(n557bar)
  );
  //OR U414
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U414 (
    .O(n557),
    .I0(in[176]),
    .I1(in[173])
  );
  //AND U414bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U414bar (
    .O(n557bar),
    .I0(inbar[176]),
    .I1(inbar[173])
  );
  //OR U415
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U415 (
    .O(n558),
    .I0(in[210]),
    .I1(in[181])
  );
  //AND U415bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U415bar (
    .O(n558bar),
    .I0(inbar[210]),
    .I1(inbar[181])
  );
  //OR U416
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U416 (
    .O(n564),
    .I0(n556),
    .I1(n555)
  );
  //AND U416bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U416bar (
    .O(n564bar),
    .I0(n556bar),
    .I1(n555bar)
  );
  //OR U417
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U417 (
    .O(n555),
    .I0(n554),
    .I1(n553)
  );
  //AND U417bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U417bar (
    .O(n555bar),
    .I0(n554bar),
    .I1(n553bar)
  );
  //OR U418
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U418 (
    .O(n553),
    .I0(in_13),
    .I1(in[234])
  );
  //AND U418bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U418bar (
    .O(n553bar),
    .I0(in_13bar),
    .I1(inbar[234])
  );
  //OR U419
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U419 (
    .O(n554),
    .I0(in_38),
    .I1(in_32)
  );
  //AND U419bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U419bar (
    .O(n554bar),
    .I0(in_38bar),
    .I1(in_32bar)
  );
  //OR U420
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U420 (
    .O(n556),
    .I0(n552),
    .I1(n551)
  );
  //AND U420bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U420bar (
    .O(n556bar),
    .I0(n552bar),
    .I1(n551bar)
  );
  //OR U421
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U421 (
    .O(n551),
    .I0(in_42),
    .I1(in_41)
  );
  //AND U421bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U421bar (
    .O(n551bar),
    .I0(in_42bar),
    .I1(in_41bar)
  );
  //OR U422
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U422 (
    .O(n552),
    .I0(in_7),
    .I1(in_49)
  );
  //AND U422bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U422bar (
    .O(n552bar),
    .I0(in_7bar),
    .I1(in_49bar)
  );
  //OR U423
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U423 (
    .O(n817),
    .I0(n550),
    .I1(n549)
  );
  //AND U423bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U423bar (
    .O(n817bar),
    .I0(n550bar),
    .I1(n549bar)
  );
  //OR U424
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U424 (
    .O(n549),
    .I0(n548),
    .I1(n547)
  );
  //AND U424bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U424bar (
    .O(n549bar),
    .I0(n548bar),
    .I1(n547bar)
  );
  //OR U425
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U425 (
    .O(n547),
    .I0(n546),
    .I1(n545)
  );
  //AND U425bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U425bar (
    .O(n547bar),
    .I0(n546bar),
    .I1(n545bar)
  );
  //OR U426
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U426 (
    .O(n545),
    .I0(in[159]),
    .I1(in[105])
  );
  //AND U426bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U426bar (
    .O(n545bar),
    .I0(inbar[159]),
    .I1(inbar[105])
  );
  //OR U427
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U427 (
    .O(n546),
    .I0(in[206]),
    .I1(in[183])
  );
  //AND U427bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U427bar (
    .O(n546bar),
    .I0(inbar[206]),
    .I1(inbar[183])
  );
  //OR U428
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U428 (
    .O(n548),
    .I0(n544),
    .I1(n543)
  );
  //AND U428bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U428bar (
    .O(n548bar),
    .I0(n544bar),
    .I1(n543bar)
  );
  //OR U429
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U429 (
    .O(n543),
    .I0(in[229]),
    .I1(in[219])
  );
  //AND U429bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U429bar (
    .O(n543bar),
    .I0(inbar[229]),
    .I1(inbar[219])
  );
  //OR U430
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U430 (
    .O(n544),
    .I0(in[235]),
    .I1(in[232])
  );
  //AND U430bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U430bar (
    .O(n544bar),
    .I0(inbar[235]),
    .I1(inbar[232])
  );
  //OR U431
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U431 (
    .O(n550),
    .I0(n542),
    .I1(n541)
  );
  //AND U431bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U431bar (
    .O(n550bar),
    .I0(n542bar),
    .I1(n541bar)
  );
  //OR U432
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U432 (
    .O(n541),
    .I0(n540),
    .I1(n539)
  );
  //AND U432bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U432bar (
    .O(n541bar),
    .I0(n540bar),
    .I1(n539bar)
  );
  //OR U433
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U433 (
    .O(n539),
    .I0(in[249]),
    .I1(in[242])
  );
  //AND U433bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U433bar (
    .O(n539bar),
    .I0(inbar[249]),
    .I1(inbar[242])
  );
  //OR U434
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U434 (
    .O(n540),
    .I0(in[89]),
    .I1(in[254])
  );
  //AND U434bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U434bar (
    .O(n540bar),
    .I0(inbar[89]),
    .I1(inbar[254])
  );
  //OR U435
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U435 (
    .O(n542),
    .I0(n538),
    .I1(n537)
  );
  //AND U435bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U435bar (
    .O(n542bar),
    .I0(n538bar),
    .I1(n537bar)
  );
  //OR U436
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U436 (
    .O(n537),
    .I0(in_14),
    .I1(in[99])
  );
  //AND U436bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U436bar (
    .O(n537bar),
    .I0(in_14bar),
    .I1(inbar[99])
  );
  //OR U437
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U437 (
    .O(n538),
    .I0(in_60),
    .I1(in_18)
  );
  //AND U437bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U437bar (
    .O(n538bar),
    .I0(in_60bar),
    .I1(in_18bar)
  );
  //OR U438
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U438 (
    .O(n566),
    .I0(in[113]),
    .I1(n763)
  );
  //AND U438bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U438bar (
    .O(n566bar),
    .I0(inbar[113]),
    .I1(n763bar)
  );
  //OR U439
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U439 (
    .O(n763),
    .I0(n536),
    .I1(n535)
  );
  //AND U439bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U439bar (
    .O(n763bar),
    .I0(n536bar),
    .I1(n535bar)
  );
  //OR U440
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U440 (
    .O(n535),
    .I0(n534),
    .I1(n533)
  );
  //AND U440bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U440bar (
    .O(n535bar),
    .I0(n534bar),
    .I1(n533bar)
  );
  //OR U441
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U441 (
    .O(n533),
    .I0(n532),
    .I1(n531)
  );
  //AND U441bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U441bar (
    .O(n533bar),
    .I0(n532bar),
    .I1(n531bar)
  );
  //OR U442
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U442 (
    .O(n531),
    .I0(in[115]),
    .I1(in[110])
  );
  //AND U442bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U442bar (
    .O(n531bar),
    .I0(inbar[115]),
    .I1(inbar[110])
  );
  //OR U443
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U443 (
    .O(n532),
    .I0(in[125]),
    .I1(in[117])
  );
  //AND U443bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U443bar (
    .O(n532bar),
    .I0(inbar[125]),
    .I1(inbar[117])
  );
  //OR U444
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U444 (
    .O(n534),
    .I0(n530),
    .I1(n529)
  );
  //AND U444bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U444bar (
    .O(n534bar),
    .I0(n530bar),
    .I1(n529bar)
  );
  //OR U445
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U445 (
    .O(n529),
    .I0(in[180]),
    .I1(in[128])
  );
  //AND U445bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U445bar (
    .O(n529bar),
    .I0(inbar[180]),
    .I1(inbar[128])
  );
  //OR U446
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U446 (
    .O(n530),
    .I0(in[205]),
    .I1(in[201])
  );
  //AND U446bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U446bar (
    .O(n530bar),
    .I0(inbar[205]),
    .I1(inbar[201])
  );
  //OR U447
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U447 (
    .O(n536),
    .I0(n528),
    .I1(n527)
  );
  //AND U447bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U447bar (
    .O(n536bar),
    .I0(n528bar),
    .I1(n527bar)
  );
  //OR U448
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U448 (
    .O(n527),
    .I0(n526),
    .I1(n525)
  );
  //AND U448bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U448bar (
    .O(n527bar),
    .I0(n526bar),
    .I1(n525bar)
  );
  //OR U449
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U449 (
    .O(n525),
    .I0(in[244]),
    .I1(in[239])
  );
  //AND U449bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U449bar (
    .O(n525bar),
    .I0(inbar[244]),
    .I1(inbar[239])
  );
  //OR U450
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U450 (
    .O(n526),
    .I0(in[95]),
    .I1(in[83])
  );
  //AND U450bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U450bar (
    .O(n526bar),
    .I0(inbar[95]),
    .I1(inbar[83])
  );
  //OR U451
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U451 (
    .O(n528),
    .I0(n524),
    .I1(n523)
  );
  //AND U451bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U451bar (
    .O(n528bar),
    .I0(n524bar),
    .I1(n523bar)
  );
  //OR U452
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U452 (
    .O(n523),
    .I0(in_24),
    .I1(in[97])
  );
  //AND U452bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U452bar (
    .O(n523bar),
    .I0(in_24bar),
    .I1(inbar[97])
  );
  //OR U453
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U453 (
    .O(n524),
    .I0(in_33),
    .I1(in_27)
  );
  //AND U453bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U453bar (
    .O(n524bar),
    .I0(in_33bar),
    .I1(in_27bar)
  );
  //OR U454
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U454 (
    .O(n568),
    .I0(n522),
    .I1(n521)
  );
  //AND U454bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U454bar (
    .O(n568bar),
    .I0(n522bar),
    .I1(n521bar)
  );
  //OR U455
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U455 (
    .O(n521),
    .I0(in[145]),
    .I1(in[126])
  );
  //AND U455bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U455bar (
    .O(n521bar),
    .I0(inbar[145]),
    .I1(inbar[126])
  );
  //OR U456
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U456 (
    .O(n522),
    .I0(in[169]),
    .I1(n520)
  );
  //AND U456bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U456bar (
    .O(n522bar),
    .I0(inbar[169]),
    .I1(n520bar)
  );
  //OR U457
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U457 (
    .O(n520),
    .I0(in[221]),
    .I1(in[172])
  );
  //AND U457bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U457bar (
    .O(n520bar),
    .I0(inbar[221]),
    .I1(inbar[172])
  );
  //OR U458
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U458 (
    .O(n570),
    .I0(n519),
    .I1(n518)
  );
  //AND U458bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U458bar (
    .O(n570bar),
    .I0(n519bar),
    .I1(n518bar)
  );
  //OR U459
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U459 (
    .O(n518),
    .I0(n517),
    .I1(n516)
  );
  //AND U459bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U459bar (
    .O(n518bar),
    .I0(n517bar),
    .I1(n516bar)
  );
  //OR U460
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U460 (
    .O(n516),
    .I0(in[241]),
    .I1(in[224])
  );
  //AND U460bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U460bar (
    .O(n516bar),
    .I0(inbar[241]),
    .I1(inbar[224])
  );
  //OR U461
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U461 (
    .O(n517),
    .I0(in[86]),
    .I1(n515)
  );
  //AND U461bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U461bar (
    .O(n517bar),
    .I0(inbar[86]),
    .I1(n515bar)
  );
  //OR U462
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U462 (
    .O(n515),
    .I0(in_43),
    .I1(in_34)
  );
  //AND U462bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U462bar (
    .O(n515bar),
    .I0(in_43bar),
    .I1(in_34bar)
  );
  //OR U463
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U463 (
    .O(n519),
    .I0(n514),
    .I1(n513)
  );
  //AND U463bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U463bar (
    .O(n519bar),
    .I0(n514bar),
    .I1(n513bar)
  );
  //OR U464
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U464 (
    .O(n513),
    .I0(in_65),
    .I1(in_51)
  );
  //AND U464bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U464bar (
    .O(n513bar),
    .I0(in_65bar),
    .I1(in_51bar)
  );
  //OR U465
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U465 (
    .O(n514),
    .I0(in_75),
    .I1(n512)
  );
  //AND U465bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U465bar (
    .O(n514bar),
    .I0(in_75bar),
    .I1(n512bar)
  );
  //OR U466
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U466 (
    .O(n512),
    .I0(in_81),
    .I1(in_77)
  );
  //AND U466bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U466bar (
    .O(n512bar),
    .I0(in_81bar),
    .I1(in_77bar)
  );
  //OR U467
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U467 (
    .O(n778),
    .I0(n511),
    .I1(n510)
  );
  //AND U467bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U467bar (
    .O(n778bar),
    .I0(n511bar),
    .I1(n510bar)
  );
  //OR U468
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U468 (
    .O(n510),
    .I0(n509),
    .I1(n508)
  );
  //AND U468bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U468bar (
    .O(n510bar),
    .I0(n509bar),
    .I1(n508bar)
  );
  //OR U469
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U469 (
    .O(n508),
    .I0(n507),
    .I1(n506)
  );
  //AND U469bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U469bar (
    .O(n508bar),
    .I0(n507bar),
    .I1(n506bar)
  );
  //OR U470
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U470 (
    .O(n506),
    .I0(in[107]),
    .I1(in[101])
  );
  //AND U470bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U470bar (
    .O(n506bar),
    .I0(inbar[107]),
    .I1(inbar[101])
  );
  //OR U471
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U471 (
    .O(n507),
    .I0(in[139]),
    .I1(in[132])
  );
  //AND U471bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U471bar (
    .O(n507bar),
    .I0(inbar[139]),
    .I1(inbar[132])
  );
  //OR U472
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U472 (
    .O(n509),
    .I0(n505),
    .I1(n504)
  );
  //AND U472bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U472bar (
    .O(n509bar),
    .I0(n505bar),
    .I1(n504bar)
  );
  //OR U473
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U473 (
    .O(n504),
    .I0(in[146]),
    .I1(in[141])
  );
  //AND U473bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U473bar (
    .O(n504bar),
    .I0(inbar[146]),
    .I1(inbar[141])
  );
  //OR U474
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U474 (
    .O(n505),
    .I0(in[203]),
    .I1(in[179])
  );
  //AND U474bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U474bar (
    .O(n505bar),
    .I0(inbar[203]),
    .I1(inbar[179])
  );
  //OR U475
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U475 (
    .O(n511),
    .I0(n503),
    .I1(n502)
  );
  //AND U475bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U475bar (
    .O(n511bar),
    .I0(n503bar),
    .I1(n502bar)
  );
  //OR U476
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U476 (
    .O(n502),
    .I0(n501),
    .I1(n500)
  );
  //AND U476bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U476bar (
    .O(n502bar),
    .I0(n501bar),
    .I1(n500bar)
  );
  //OR U477
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U477 (
    .O(n500),
    .I0(in[243]),
    .I1(in[222])
  );
  //AND U477bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U477bar (
    .O(n500bar),
    .I0(inbar[243]),
    .I1(inbar[222])
  );
  //OR U478
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U478 (
    .O(n501),
    .I0(in[251]),
    .I1(in[250])
  );
  //AND U478bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U478bar (
    .O(n501bar),
    .I0(inbar[251]),
    .I1(inbar[250])
  );
  //OR U479
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U479 (
    .O(n503),
    .I0(n499),
    .I1(n498)
  );
  //AND U479bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U479bar (
    .O(n503bar),
    .I0(n499bar),
    .I1(n498bar)
  );
  //OR U480
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U480 (
    .O(n498),
    .I0(in_37),
    .I1(in_19)
  );
  //AND U480bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U480bar (
    .O(n498bar),
    .I0(in_37bar),
    .I1(in_19bar)
  );
  //OR U481
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U481 (
    .O(n499),
    .I0(in_78),
    .I1(in_6)
  );
  //AND U481bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U481bar (
    .O(n499bar),
    .I0(in_78bar),
    .I1(in_6bar)
  );
  //OR U482
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U482 (
    .O(n603),
    .I0(n497),
    .I1(n496)
  );
  //AND U482bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U482bar (
    .O(n603bar),
    .I0(n497bar),
    .I1(n496bar)
  );
  //OR U483
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U483 (
    .O(n496),
    .I0(in[112]),
    .I1(in[102])
  );
  //AND U483bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U483bar (
    .O(n496bar),
    .I0(inbar[112]),
    .I1(inbar[102])
  );
  //OR U484
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U484 (
    .O(n497),
    .I0(in[123]),
    .I1(n495)
  );
  //AND U484bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U484bar (
    .O(n497bar),
    .I0(inbar[123]),
    .I1(n495bar)
  );
  //OR U485
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U485 (
    .O(n495),
    .I0(in[143]),
    .I1(in[130])
  );
  //AND U485bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U485bar (
    .O(n495bar),
    .I0(inbar[143]),
    .I1(inbar[130])
  );
  //OR U486
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U486 (
    .O(n605),
    .I0(n494),
    .I1(n493)
  );
  //AND U486bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U486bar (
    .O(n605bar),
    .I0(n494bar),
    .I1(n493bar)
  );
  //OR U487
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U487 (
    .O(n493),
    .I0(n492),
    .I1(n491)
  );
  //AND U487bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U487bar (
    .O(n493bar),
    .I0(n492bar),
    .I1(n491bar)
  );
  //OR U488
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U488 (
    .O(n491),
    .I0(in[216]),
    .I1(in[213])
  );
  //AND U488bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U488bar (
    .O(n491bar),
    .I0(inbar[216]),
    .I1(inbar[213])
  );
  //OR U489
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U489 (
    .O(n492),
    .I0(in[227]),
    .I1(n490)
  );
  //AND U489bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U489bar (
    .O(n492bar),
    .I0(inbar[227]),
    .I1(n490bar)
  );
  //OR U490
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U490 (
    .O(n490),
    .I0(in_0),
    .I1(in[248])
  );
  //AND U490bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U490bar (
    .O(n490bar),
    .I0(in_0bar),
    .I1(inbar[248])
  );
  //OR U491
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U491 (
    .O(n494),
    .I0(n489),
    .I1(n488)
  );
  //AND U491bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U491bar (
    .O(n494bar),
    .I0(n489bar),
    .I1(n488bar)
  );
  //OR U492
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U492 (
    .O(n488),
    .I0(in_46),
    .I1(in_44)
  );
  //AND U492bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U492bar (
    .O(n488bar),
    .I0(in_46bar),
    .I1(in_44bar)
  );
  //OR U493
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U493 (
    .O(n489),
    .I0(in_50),
    .I1(n487)
  );
  //AND U493bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U493bar (
    .O(n489bar),
    .I0(in_50bar),
    .I1(n487bar)
  );
  //OR U494
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U494 (
    .O(n487),
    .I0(in_9),
    .I1(in_80)
  );
  //AND U494bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U494bar (
    .O(n487bar),
    .I0(in_9bar),
    .I1(in_80bar)
  );
endmodule

module sBox_14 ( in, out );

  input wire [7:0] in;
//input_done

  output wire [7:0] out;
//output_done

  wire [255:0] decodeOut;
//wire_done

  decode_14 dec ( .in(in), .out(decodeOut) );
  encode_14 enc ( .in(decodeOut), .out(out) );
endmodule

module CD2_57 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD2_58 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD2_59 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD2_60 ( a, b, y );

  input wire a;
  input wire b;
  wire abar;
  wire bbar;
  assign abar = ~a;
  assign bbar = ~b;
//input_done

  output wire [3:0] y;
  wire [3:0] ybar;
//output_done

  wire n3;
  wire n4;
  wire n3bar;
  wire n4bar;
//wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[3]),
    .I0(b),
    .I1(a)
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[3]),
    .I0(bbar),
    .I1(abar)
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[2]),
    .I0(a),
    .I1(n3)
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[2]),
    .I0(abar),
    .I1(n3bar)
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[1]),
    .I0(b),
    .I1(n4)
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[1]),
    .I0(bbar),
    .I1(n4bar)
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[0]),
    .I0(n4),
    .I1(n3)
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[0]),
    .I0(n4bar),
    .I1(n3bar)
  );
endmodule

module CD4_29 ( a, b, y );

  input wire [3:0] a;
  input wire [3:0] b;
  wire [3:0] abar;
  wire [3:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
//input_done

  output wire [15:0] y;
  wire [15:0] ybar;
//output_done

//wire_done

  //AND U1
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1 (
    .O(y[9]),
    .I0(b[1]),
    .I1(a[2])
  );
  //OR U1bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1bar (
    .O(ybar[9]),
    .I0(bbar[1]),
    .I1(abar[2])
  );
  //AND U2
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2 (
    .O(y[8]),
    .I0(b[0]),
    .I1(a[2])
  );
  //OR U2bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2bar (
    .O(ybar[8]),
    .I0(bbar[0]),
    .I1(abar[2])
  );
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[7]),
    .I0(b[3]),
    .I1(a[1])
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[7]),
    .I0(bbar[3]),
    .I1(abar[1])
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[6]),
    .I0(b[2]),
    .I1(a[1])
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[6]),
    .I0(bbar[2]),
    .I1(abar[1])
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[5]),
    .I0(a[1]),
    .I1(b[1])
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[5]),
    .I0(abar[1]),
    .I1(bbar[1])
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[4]),
    .I0(a[1]),
    .I1(b[0])
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[4]),
    .I0(abar[1]),
    .I1(bbar[0])
  );
  //AND U7
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7 (
    .O(y[3]),
    .I0(a[0]),
    .I1(b[3])
  );
  //OR U7bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7bar (
    .O(ybar[3]),
    .I0(abar[0]),
    .I1(bbar[3])
  );
  //AND U8
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8 (
    .O(y[2]),
    .I0(a[0]),
    .I1(b[2])
  );
  //OR U8bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8bar (
    .O(ybar[2]),
    .I0(abar[0]),
    .I1(bbar[2])
  );
  //AND U9
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9 (
    .O(y[1]),
    .I0(a[0]),
    .I1(b[1])
  );
  //OR U9bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9bar (
    .O(ybar[1]),
    .I0(abar[0]),
    .I1(bbar[1])
  );
  //AND U10
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10 (
    .O(y[15]),
    .I0(a[3]),
    .I1(b[3])
  );
  //OR U10bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10bar (
    .O(ybar[15]),
    .I0(abar[3]),
    .I1(bbar[3])
  );
  //AND U11
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11 (
    .O(y[14]),
    .I0(a[3]),
    .I1(b[2])
  );
  //OR U11bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11bar (
    .O(ybar[14]),
    .I0(abar[3]),
    .I1(bbar[2])
  );
  //AND U12
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12 (
    .O(y[13]),
    .I0(a[3]),
    .I1(b[1])
  );
  //OR U12bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12bar (
    .O(ybar[13]),
    .I0(abar[3]),
    .I1(bbar[1])
  );
  //AND U13
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13 (
    .O(y[12]),
    .I0(a[3]),
    .I1(b[0])
  );
  //OR U13bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13bar (
    .O(ybar[12]),
    .I0(abar[3]),
    .I1(bbar[0])
  );
  //AND U14
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14 (
    .O(y[11]),
    .I0(b[3]),
    .I1(a[2])
  );
  //OR U14bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14bar (
    .O(ybar[11]),
    .I0(bbar[3]),
    .I1(abar[2])
  );
  //AND U15
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15 (
    .O(y[10]),
    .I0(b[2]),
    .I1(a[2])
  );
  //OR U15bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15bar (
    .O(ybar[10]),
    .I0(bbar[2]),
    .I1(abar[2])
  );
  //AND U16
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16 (
    .O(y[0]),
    .I0(a[0]),
    .I1(b[0])
  );
  //OR U16bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16bar (
    .O(ybar[0]),
    .I0(abar[0]),
    .I1(bbar[0])
  );
endmodule

module CD4_30 ( a, b, y );

  input wire [3:0] a;
  input wire [3:0] b;
  wire [3:0] abar;
  wire [3:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
//input_done

  output wire [15:0] y;
  wire [15:0] ybar;
//output_done

//wire_done

  //AND U1
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1 (
    .O(y[9]),
    .I0(b[1]),
    .I1(a[2])
  );
  //OR U1bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1bar (
    .O(ybar[9]),
    .I0(bbar[1]),
    .I1(abar[2])
  );
  //AND U2
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2 (
    .O(y[8]),
    .I0(b[0]),
    .I1(a[2])
  );
  //OR U2bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2bar (
    .O(ybar[8]),
    .I0(bbar[0]),
    .I1(abar[2])
  );
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[7]),
    .I0(b[3]),
    .I1(a[1])
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[7]),
    .I0(bbar[3]),
    .I1(abar[1])
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[6]),
    .I0(b[2]),
    .I1(a[1])
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[6]),
    .I0(bbar[2]),
    .I1(abar[1])
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[5]),
    .I0(a[1]),
    .I1(b[1])
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[5]),
    .I0(abar[1]),
    .I1(bbar[1])
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[4]),
    .I0(a[1]),
    .I1(b[0])
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[4]),
    .I0(abar[1]),
    .I1(bbar[0])
  );
  //AND U7
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7 (
    .O(y[3]),
    .I0(a[0]),
    .I1(b[3])
  );
  //OR U7bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7bar (
    .O(ybar[3]),
    .I0(abar[0]),
    .I1(bbar[3])
  );
  //AND U8
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8 (
    .O(y[2]),
    .I0(a[0]),
    .I1(b[2])
  );
  //OR U8bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8bar (
    .O(ybar[2]),
    .I0(abar[0]),
    .I1(bbar[2])
  );
  //AND U9
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9 (
    .O(y[1]),
    .I0(a[0]),
    .I1(b[1])
  );
  //OR U9bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9bar (
    .O(ybar[1]),
    .I0(abar[0]),
    .I1(bbar[1])
  );
  //AND U10
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10 (
    .O(y[15]),
    .I0(a[3]),
    .I1(b[3])
  );
  //OR U10bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10bar (
    .O(ybar[15]),
    .I0(abar[3]),
    .I1(bbar[3])
  );
  //AND U11
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11 (
    .O(y[14]),
    .I0(a[3]),
    .I1(b[2])
  );
  //OR U11bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11bar (
    .O(ybar[14]),
    .I0(abar[3]),
    .I1(bbar[2])
  );
  //AND U12
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12 (
    .O(y[13]),
    .I0(a[3]),
    .I1(b[1])
  );
  //OR U12bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12bar (
    .O(ybar[13]),
    .I0(abar[3]),
    .I1(bbar[1])
  );
  //AND U13
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13 (
    .O(y[12]),
    .I0(a[3]),
    .I1(b[0])
  );
  //OR U13bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13bar (
    .O(ybar[12]),
    .I0(abar[3]),
    .I1(bbar[0])
  );
  //AND U14
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14 (
    .O(y[11]),
    .I0(b[3]),
    .I1(a[2])
  );
  //OR U14bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14bar (
    .O(ybar[11]),
    .I0(bbar[3]),
    .I1(abar[2])
  );
  //AND U15
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15 (
    .O(y[10]),
    .I0(b[2]),
    .I1(a[2])
  );
  //OR U15bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15bar (
    .O(ybar[10]),
    .I0(bbar[2]),
    .I1(abar[2])
  );
  //AND U16
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16 (
    .O(y[0]),
    .I0(a[0]),
    .I1(b[0])
  );
  //OR U16bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16bar (
    .O(ybar[0]),
    .I0(abar[0]),
    .I1(bbar[0])
  );
endmodule

module CD16_15 ( a, b, y );

  input wire [15:0] a;
  input wire [15:0] b;
  wire [15:0] abar;
  wire [15:0] bbar;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign abar[8] = ~a[8];
  assign abar[9] = ~a[9];
  assign abar[10] = ~a[10];
  assign abar[11] = ~a[11];
  assign abar[12] = ~a[12];
  assign abar[13] = ~a[13];
  assign abar[14] = ~a[14];
  assign abar[15] = ~a[15];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign bbar[8] = ~b[8];
  assign bbar[9] = ~b[9];
  assign bbar[10] = ~b[10];
  assign bbar[11] = ~b[11];
  assign bbar[12] = ~b[12];
  assign bbar[13] = ~b[13];
  assign bbar[14] = ~b[14];
  assign bbar[15] = ~b[15];
//input_done

  output wire [255:0] y;
  wire [255:0] ybar;
//output_done

//wire_done

  //AND U1
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1 (
    .O(y[9]),
    .I0(b[9]),
    .I1(a[0])
  );
  //OR U1bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1bar (
    .O(ybar[9]),
    .I0(bbar[9]),
    .I1(abar[0])
  );
  //AND U2
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2 (
    .O(y[99]),
    .I0(b[3]),
    .I1(a[6])
  );
  //OR U2bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2bar (
    .O(ybar[99]),
    .I0(bbar[3]),
    .I1(abar[6])
  );
  //AND U3
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3 (
    .O(y[98]),
    .I0(b[2]),
    .I1(a[6])
  );
  //OR U3bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3bar (
    .O(ybar[98]),
    .I0(bbar[2]),
    .I1(abar[6])
  );
  //AND U4
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4 (
    .O(y[97]),
    .I0(b[1]),
    .I1(a[6])
  );
  //OR U4bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4bar (
    .O(ybar[97]),
    .I0(bbar[1]),
    .I1(abar[6])
  );
  //AND U5
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5 (
    .O(y[96]),
    .I0(b[0]),
    .I1(a[6])
  );
  //OR U5bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5bar (
    .O(ybar[96]),
    .I0(bbar[0]),
    .I1(abar[6])
  );
  //AND U6
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6 (
    .O(y[95]),
    .I0(b[15]),
    .I1(a[5])
  );
  //OR U6bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6bar (
    .O(ybar[95]),
    .I0(bbar[15]),
    .I1(abar[5])
  );
  //AND U7
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7 (
    .O(y[94]),
    .I0(b[14]),
    .I1(a[5])
  );
  //OR U7bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7bar (
    .O(ybar[94]),
    .I0(bbar[14]),
    .I1(abar[5])
  );
  //AND U8
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8 (
    .O(y[93]),
    .I0(b[13]),
    .I1(a[5])
  );
  //OR U8bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8bar (
    .O(ybar[93]),
    .I0(bbar[13]),
    .I1(abar[5])
  );
  //AND U9
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9 (
    .O(y[92]),
    .I0(b[12]),
    .I1(a[5])
  );
  //OR U9bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9bar (
    .O(ybar[92]),
    .I0(bbar[12]),
    .I1(abar[5])
  );
  //AND U10
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10 (
    .O(y[91]),
    .I0(b[11]),
    .I1(a[5])
  );
  //OR U10bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10bar (
    .O(ybar[91]),
    .I0(bbar[11]),
    .I1(abar[5])
  );
  //AND U11
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11 (
    .O(y[90]),
    .I0(b[10]),
    .I1(a[5])
  );
  //OR U11bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11bar (
    .O(ybar[90]),
    .I0(bbar[10]),
    .I1(abar[5])
  );
  //AND U12
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12 (
    .O(y[8]),
    .I0(b[8]),
    .I1(a[0])
  );
  //OR U12bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12bar (
    .O(ybar[8]),
    .I0(bbar[8]),
    .I1(abar[0])
  );
  //AND U13
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13 (
    .O(y[89]),
    .I0(a[5]),
    .I1(b[9])
  );
  //OR U13bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13bar (
    .O(ybar[89]),
    .I0(abar[5]),
    .I1(bbar[9])
  );
  //AND U14
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14 (
    .O(y[88]),
    .I0(b[8]),
    .I1(a[5])
  );
  //OR U14bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14bar (
    .O(ybar[88]),
    .I0(bbar[8]),
    .I1(abar[5])
  );
  //AND U15
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15 (
    .O(y[87]),
    .I0(b[7]),
    .I1(a[5])
  );
  //OR U15bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15bar (
    .O(ybar[87]),
    .I0(bbar[7]),
    .I1(abar[5])
  );
  //AND U16
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16 (
    .O(y[86]),
    .I0(b[6]),
    .I1(a[5])
  );
  //OR U16bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16bar (
    .O(ybar[86]),
    .I0(bbar[6]),
    .I1(abar[5])
  );
  //AND U17
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U17 (
    .O(y[85]),
    .I0(b[5]),
    .I1(a[5])
  );
  //OR U17bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U17bar (
    .O(ybar[85]),
    .I0(bbar[5]),
    .I1(abar[5])
  );
  //AND U18
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U18 (
    .O(y[84]),
    .I0(b[4]),
    .I1(a[5])
  );
  //OR U18bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U18bar (
    .O(ybar[84]),
    .I0(bbar[4]),
    .I1(abar[5])
  );
  //AND U19
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U19 (
    .O(y[83]),
    .I0(a[5]),
    .I1(b[3])
  );
  //OR U19bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U19bar (
    .O(ybar[83]),
    .I0(abar[5]),
    .I1(bbar[3])
  );
  //AND U20
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U20 (
    .O(y[82]),
    .I0(a[5]),
    .I1(b[2])
  );
  //OR U20bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U20bar (
    .O(ybar[82]),
    .I0(abar[5]),
    .I1(bbar[2])
  );
  //AND U21
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U21 (
    .O(y[81]),
    .I0(a[5]),
    .I1(b[1])
  );
  //OR U21bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U21bar (
    .O(ybar[81]),
    .I0(abar[5]),
    .I1(bbar[1])
  );
  //AND U22
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U22 (
    .O(y[80]),
    .I0(a[5]),
    .I1(b[0])
  );
  //OR U22bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U22bar (
    .O(ybar[80]),
    .I0(abar[5]),
    .I1(bbar[0])
  );
  //AND U23
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U23 (
    .O(y[7]),
    .I0(b[7]),
    .I1(a[0])
  );
  //OR U23bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U23bar (
    .O(ybar[7]),
    .I0(bbar[7]),
    .I1(abar[0])
  );
  //AND U24
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U24 (
    .O(y[79]),
    .I0(a[4]),
    .I1(b[15])
  );
  //OR U24bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U24bar (
    .O(ybar[79]),
    .I0(abar[4]),
    .I1(bbar[15])
  );
  //AND U25
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U25 (
    .O(y[78]),
    .I0(a[4]),
    .I1(b[14])
  );
  //OR U25bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U25bar (
    .O(ybar[78]),
    .I0(abar[4]),
    .I1(bbar[14])
  );
  //AND U26
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U26 (
    .O(y[77]),
    .I0(a[4]),
    .I1(b[13])
  );
  //OR U26bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U26bar (
    .O(ybar[77]),
    .I0(abar[4]),
    .I1(bbar[13])
  );
  //AND U27
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U27 (
    .O(y[76]),
    .I0(a[4]),
    .I1(b[12])
  );
  //OR U27bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U27bar (
    .O(ybar[76]),
    .I0(abar[4]),
    .I1(bbar[12])
  );
  //AND U28
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U28 (
    .O(y[75]),
    .I0(a[4]),
    .I1(b[11])
  );
  //OR U28bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U28bar (
    .O(ybar[75]),
    .I0(abar[4]),
    .I1(bbar[11])
  );
  //AND U29
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U29 (
    .O(y[74]),
    .I0(a[4]),
    .I1(b[10])
  );
  //OR U29bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U29bar (
    .O(ybar[74]),
    .I0(abar[4]),
    .I1(bbar[10])
  );
  //AND U30
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U30 (
    .O(y[73]),
    .I0(a[4]),
    .I1(b[9])
  );
  //OR U30bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U30bar (
    .O(ybar[73]),
    .I0(abar[4]),
    .I1(bbar[9])
  );
  //AND U31
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U31 (
    .O(y[72]),
    .I0(a[4]),
    .I1(b[8])
  );
  //OR U31bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U31bar (
    .O(ybar[72]),
    .I0(abar[4]),
    .I1(bbar[8])
  );
  //AND U32
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U32 (
    .O(y[71]),
    .I0(a[4]),
    .I1(b[7])
  );
  //OR U32bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U32bar (
    .O(ybar[71]),
    .I0(abar[4]),
    .I1(bbar[7])
  );
  //AND U33
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U33 (
    .O(y[70]),
    .I0(a[4]),
    .I1(b[6])
  );
  //OR U33bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U33bar (
    .O(ybar[70]),
    .I0(abar[4]),
    .I1(bbar[6])
  );
  //AND U34
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U34 (
    .O(y[6]),
    .I0(b[6]),
    .I1(a[0])
  );
  //OR U34bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U34bar (
    .O(ybar[6]),
    .I0(bbar[6]),
    .I1(abar[0])
  );
  //AND U35
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U35 (
    .O(y[69]),
    .I0(a[4]),
    .I1(b[5])
  );
  //OR U35bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U35bar (
    .O(ybar[69]),
    .I0(abar[4]),
    .I1(bbar[5])
  );
  //AND U36
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U36 (
    .O(y[68]),
    .I0(a[4]),
    .I1(b[4])
  );
  //OR U36bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U36bar (
    .O(ybar[68]),
    .I0(abar[4]),
    .I1(bbar[4])
  );
  //AND U37
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U37 (
    .O(y[67]),
    .I0(a[4]),
    .I1(b[3])
  );
  //OR U37bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U37bar (
    .O(ybar[67]),
    .I0(abar[4]),
    .I1(bbar[3])
  );
  //AND U38
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U38 (
    .O(y[66]),
    .I0(a[4]),
    .I1(b[2])
  );
  //OR U38bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U38bar (
    .O(ybar[66]),
    .I0(abar[4]),
    .I1(bbar[2])
  );
  //AND U39
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U39 (
    .O(y[65]),
    .I0(a[4]),
    .I1(b[1])
  );
  //OR U39bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U39bar (
    .O(ybar[65]),
    .I0(abar[4]),
    .I1(bbar[1])
  );
  //AND U40
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U40 (
    .O(y[64]),
    .I0(a[4]),
    .I1(b[0])
  );
  //OR U40bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U40bar (
    .O(ybar[64]),
    .I0(abar[4]),
    .I1(bbar[0])
  );
  //AND U41
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U41 (
    .O(y[63]),
    .I0(a[3]),
    .I1(b[15])
  );
  //OR U41bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U41bar (
    .O(ybar[63]),
    .I0(abar[3]),
    .I1(bbar[15])
  );
  //AND U42
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U42 (
    .O(y[62]),
    .I0(a[3]),
    .I1(b[14])
  );
  //OR U42bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U42bar (
    .O(ybar[62]),
    .I0(abar[3]),
    .I1(bbar[14])
  );
  //AND U43
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U43 (
    .O(y[61]),
    .I0(a[3]),
    .I1(b[13])
  );
  //OR U43bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U43bar (
    .O(ybar[61]),
    .I0(abar[3]),
    .I1(bbar[13])
  );
  //AND U44
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U44 (
    .O(y[60]),
    .I0(a[3]),
    .I1(b[12])
  );
  //OR U44bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U44bar (
    .O(ybar[60]),
    .I0(abar[3]),
    .I1(bbar[12])
  );
  //AND U45
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U45 (
    .O(y[5]),
    .I0(b[5]),
    .I1(a[0])
  );
  //OR U45bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U45bar (
    .O(ybar[5]),
    .I0(bbar[5]),
    .I1(abar[0])
  );
  //AND U46
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U46 (
    .O(y[59]),
    .I0(a[3]),
    .I1(b[11])
  );
  //OR U46bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U46bar (
    .O(ybar[59]),
    .I0(abar[3]),
    .I1(bbar[11])
  );
  //AND U47
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U47 (
    .O(y[58]),
    .I0(a[3]),
    .I1(b[10])
  );
  //OR U47bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U47bar (
    .O(ybar[58]),
    .I0(abar[3]),
    .I1(bbar[10])
  );
  //AND U48
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U48 (
    .O(y[57]),
    .I0(a[3]),
    .I1(b[9])
  );
  //OR U48bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U48bar (
    .O(ybar[57]),
    .I0(abar[3]),
    .I1(bbar[9])
  );
  //AND U49
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U49 (
    .O(y[56]),
    .I0(a[3]),
    .I1(b[8])
  );
  //OR U49bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U49bar (
    .O(ybar[56]),
    .I0(abar[3]),
    .I1(bbar[8])
  );
  //AND U50
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U50 (
    .O(y[55]),
    .I0(a[3]),
    .I1(b[7])
  );
  //OR U50bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U50bar (
    .O(ybar[55]),
    .I0(abar[3]),
    .I1(bbar[7])
  );
  //AND U51
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U51 (
    .O(y[54]),
    .I0(a[3]),
    .I1(b[6])
  );
  //OR U51bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U51bar (
    .O(ybar[54]),
    .I0(abar[3]),
    .I1(bbar[6])
  );
  //AND U52
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U52 (
    .O(y[53]),
    .I0(a[3]),
    .I1(b[5])
  );
  //OR U52bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U52bar (
    .O(ybar[53]),
    .I0(abar[3]),
    .I1(bbar[5])
  );
  //AND U53
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U53 (
    .O(y[52]),
    .I0(a[3]),
    .I1(b[4])
  );
  //OR U53bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U53bar (
    .O(ybar[52]),
    .I0(abar[3]),
    .I1(bbar[4])
  );
  //AND U54
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U54 (
    .O(y[51]),
    .I0(a[3]),
    .I1(b[3])
  );
  //OR U54bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U54bar (
    .O(ybar[51]),
    .I0(abar[3]),
    .I1(bbar[3])
  );
  //AND U55
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U55 (
    .O(y[50]),
    .I0(a[3]),
    .I1(b[2])
  );
  //OR U55bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U55bar (
    .O(ybar[50]),
    .I0(abar[3]),
    .I1(bbar[2])
  );
  //AND U56
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U56 (
    .O(y[4]),
    .I0(b[4]),
    .I1(a[0])
  );
  //OR U56bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U56bar (
    .O(ybar[4]),
    .I0(bbar[4]),
    .I1(abar[0])
  );
  //AND U57
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U57 (
    .O(y[49]),
    .I0(a[3]),
    .I1(b[1])
  );
  //OR U57bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U57bar (
    .O(ybar[49]),
    .I0(abar[3]),
    .I1(bbar[1])
  );
  //AND U58
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U58 (
    .O(y[48]),
    .I0(a[3]),
    .I1(b[0])
  );
  //OR U58bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U58bar (
    .O(ybar[48]),
    .I0(abar[3]),
    .I1(bbar[0])
  );
  //AND U59
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U59 (
    .O(y[47]),
    .I0(a[2]),
    .I1(b[15])
  );
  //OR U59bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U59bar (
    .O(ybar[47]),
    .I0(abar[2]),
    .I1(bbar[15])
  );
  //AND U60
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U60 (
    .O(y[46]),
    .I0(a[2]),
    .I1(b[14])
  );
  //OR U60bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U60bar (
    .O(ybar[46]),
    .I0(abar[2]),
    .I1(bbar[14])
  );
  //AND U61
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U61 (
    .O(y[45]),
    .I0(a[2]),
    .I1(b[13])
  );
  //OR U61bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U61bar (
    .O(ybar[45]),
    .I0(abar[2]),
    .I1(bbar[13])
  );
  //AND U62
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U62 (
    .O(y[44]),
    .I0(a[2]),
    .I1(b[12])
  );
  //OR U62bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U62bar (
    .O(ybar[44]),
    .I0(abar[2]),
    .I1(bbar[12])
  );
  //AND U63
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U63 (
    .O(y[43]),
    .I0(a[2]),
    .I1(b[11])
  );
  //OR U63bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U63bar (
    .O(ybar[43]),
    .I0(abar[2]),
    .I1(bbar[11])
  );
  //AND U64
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U64 (
    .O(y[42]),
    .I0(a[2]),
    .I1(b[10])
  );
  //OR U64bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U64bar (
    .O(ybar[42]),
    .I0(abar[2]),
    .I1(bbar[10])
  );
  //AND U65
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U65 (
    .O(y[41]),
    .I0(a[2]),
    .I1(b[9])
  );
  //OR U65bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U65bar (
    .O(ybar[41]),
    .I0(abar[2]),
    .I1(bbar[9])
  );
  //AND U66
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U66 (
    .O(y[40]),
    .I0(a[2]),
    .I1(b[8])
  );
  //OR U66bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U66bar (
    .O(ybar[40]),
    .I0(abar[2]),
    .I1(bbar[8])
  );
  //AND U67
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U67 (
    .O(y[3]),
    .I0(b[3]),
    .I1(a[0])
  );
  //OR U67bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U67bar (
    .O(ybar[3]),
    .I0(bbar[3]),
    .I1(abar[0])
  );
  //AND U68
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U68 (
    .O(y[39]),
    .I0(a[2]),
    .I1(b[7])
  );
  //OR U68bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U68bar (
    .O(ybar[39]),
    .I0(abar[2]),
    .I1(bbar[7])
  );
  //AND U69
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U69 (
    .O(y[38]),
    .I0(a[2]),
    .I1(b[6])
  );
  //OR U69bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U69bar (
    .O(ybar[38]),
    .I0(abar[2]),
    .I1(bbar[6])
  );
  //AND U70
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U70 (
    .O(y[37]),
    .I0(a[2]),
    .I1(b[5])
  );
  //OR U70bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U70bar (
    .O(ybar[37]),
    .I0(abar[2]),
    .I1(bbar[5])
  );
  //AND U71
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U71 (
    .O(y[36]),
    .I0(a[2]),
    .I1(b[4])
  );
  //OR U71bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U71bar (
    .O(ybar[36]),
    .I0(abar[2]),
    .I1(bbar[4])
  );
  //AND U72
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U72 (
    .O(y[35]),
    .I0(a[2]),
    .I1(b[3])
  );
  //OR U72bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U72bar (
    .O(ybar[35]),
    .I0(abar[2]),
    .I1(bbar[3])
  );
  //AND U73
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U73 (
    .O(y[34]),
    .I0(a[2]),
    .I1(b[2])
  );
  //OR U73bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U73bar (
    .O(ybar[34]),
    .I0(abar[2]),
    .I1(bbar[2])
  );
  //AND U74
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U74 (
    .O(y[33]),
    .I0(a[2]),
    .I1(b[1])
  );
  //OR U74bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U74bar (
    .O(ybar[33]),
    .I0(abar[2]),
    .I1(bbar[1])
  );
  //AND U75
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U75 (
    .O(y[32]),
    .I0(a[2]),
    .I1(b[0])
  );
  //OR U75bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U75bar (
    .O(ybar[32]),
    .I0(abar[2]),
    .I1(bbar[0])
  );
  //AND U76
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U76 (
    .O(y[31]),
    .I0(a[1]),
    .I1(b[15])
  );
  //OR U76bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U76bar (
    .O(ybar[31]),
    .I0(abar[1]),
    .I1(bbar[15])
  );
  //AND U77
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U77 (
    .O(y[30]),
    .I0(a[1]),
    .I1(b[14])
  );
  //OR U77bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U77bar (
    .O(ybar[30]),
    .I0(abar[1]),
    .I1(bbar[14])
  );
  //AND U78
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U78 (
    .O(y[2]),
    .I0(b[2]),
    .I1(a[0])
  );
  //OR U78bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U78bar (
    .O(ybar[2]),
    .I0(bbar[2]),
    .I1(abar[0])
  );
  //AND U79
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U79 (
    .O(y[29]),
    .I0(a[1]),
    .I1(b[13])
  );
  //OR U79bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U79bar (
    .O(ybar[29]),
    .I0(abar[1]),
    .I1(bbar[13])
  );
  //AND U80
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U80 (
    .O(y[28]),
    .I0(a[1]),
    .I1(b[12])
  );
  //OR U80bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U80bar (
    .O(ybar[28]),
    .I0(abar[1]),
    .I1(bbar[12])
  );
  //AND U81
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U81 (
    .O(y[27]),
    .I0(a[1]),
    .I1(b[11])
  );
  //OR U81bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U81bar (
    .O(ybar[27]),
    .I0(abar[1]),
    .I1(bbar[11])
  );
  //AND U82
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U82 (
    .O(y[26]),
    .I0(a[1]),
    .I1(b[10])
  );
  //OR U82bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U82bar (
    .O(ybar[26]),
    .I0(abar[1]),
    .I1(bbar[10])
  );
  //AND U83
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U83 (
    .O(y[25]),
    .I0(a[1]),
    .I1(b[9])
  );
  //OR U83bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U83bar (
    .O(ybar[25]),
    .I0(abar[1]),
    .I1(bbar[9])
  );
  //AND U84
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U84 (
    .O(y[255]),
    .I0(a[15]),
    .I1(b[15])
  );
  //OR U84bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U84bar (
    .O(ybar[255]),
    .I0(abar[15]),
    .I1(bbar[15])
  );
  //AND U85
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U85 (
    .O(y[254]),
    .I0(a[15]),
    .I1(b[14])
  );
  //OR U85bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U85bar (
    .O(ybar[254]),
    .I0(abar[15]),
    .I1(bbar[14])
  );
  //AND U86
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U86 (
    .O(y[253]),
    .I0(a[15]),
    .I1(b[13])
  );
  //OR U86bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U86bar (
    .O(ybar[253]),
    .I0(abar[15]),
    .I1(bbar[13])
  );
  //AND U87
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U87 (
    .O(y[252]),
    .I0(a[15]),
    .I1(b[12])
  );
  //OR U87bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U87bar (
    .O(ybar[252]),
    .I0(abar[15]),
    .I1(bbar[12])
  );
  //AND U88
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U88 (
    .O(y[251]),
    .I0(a[15]),
    .I1(b[11])
  );
  //OR U88bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U88bar (
    .O(ybar[251]),
    .I0(abar[15]),
    .I1(bbar[11])
  );
  //AND U89
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U89 (
    .O(y[250]),
    .I0(a[15]),
    .I1(b[10])
  );
  //OR U89bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U89bar (
    .O(ybar[250]),
    .I0(abar[15]),
    .I1(bbar[10])
  );
  //AND U90
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U90 (
    .O(y[24]),
    .I0(a[1]),
    .I1(b[8])
  );
  //OR U90bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U90bar (
    .O(ybar[24]),
    .I0(abar[1]),
    .I1(bbar[8])
  );
  //AND U91
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U91 (
    .O(y[249]),
    .I0(a[15]),
    .I1(b[9])
  );
  //OR U91bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U91bar (
    .O(ybar[249]),
    .I0(abar[15]),
    .I1(bbar[9])
  );
  //AND U92
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U92 (
    .O(y[248]),
    .I0(a[15]),
    .I1(b[8])
  );
  //OR U92bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U92bar (
    .O(ybar[248]),
    .I0(abar[15]),
    .I1(bbar[8])
  );
  //AND U93
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U93 (
    .O(y[247]),
    .I0(a[15]),
    .I1(b[7])
  );
  //OR U93bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U93bar (
    .O(ybar[247]),
    .I0(abar[15]),
    .I1(bbar[7])
  );
  //AND U94
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U94 (
    .O(y[246]),
    .I0(a[15]),
    .I1(b[6])
  );
  //OR U94bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U94bar (
    .O(ybar[246]),
    .I0(abar[15]),
    .I1(bbar[6])
  );
  //AND U95
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U95 (
    .O(y[245]),
    .I0(a[15]),
    .I1(b[5])
  );
  //OR U95bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U95bar (
    .O(ybar[245]),
    .I0(abar[15]),
    .I1(bbar[5])
  );
  //AND U96
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U96 (
    .O(y[244]),
    .I0(a[15]),
    .I1(b[4])
  );
  //OR U96bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U96bar (
    .O(ybar[244]),
    .I0(abar[15]),
    .I1(bbar[4])
  );
  //AND U97
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U97 (
    .O(y[243]),
    .I0(a[15]),
    .I1(b[3])
  );
  //OR U97bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U97bar (
    .O(ybar[243]),
    .I0(abar[15]),
    .I1(bbar[3])
  );
  //AND U98
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U98 (
    .O(y[242]),
    .I0(a[15]),
    .I1(b[2])
  );
  //OR U98bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U98bar (
    .O(ybar[242]),
    .I0(abar[15]),
    .I1(bbar[2])
  );
  //AND U99
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U99 (
    .O(y[241]),
    .I0(a[15]),
    .I1(b[1])
  );
  //OR U99bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U99bar (
    .O(ybar[241]),
    .I0(abar[15]),
    .I1(bbar[1])
  );
  //AND U100
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U100 (
    .O(y[240]),
    .I0(a[15]),
    .I1(b[0])
  );
  //OR U100bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U100bar (
    .O(ybar[240]),
    .I0(abar[15]),
    .I1(bbar[0])
  );
  //AND U101
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U101 (
    .O(y[23]),
    .I0(a[1]),
    .I1(b[7])
  );
  //OR U101bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U101bar (
    .O(ybar[23]),
    .I0(abar[1]),
    .I1(bbar[7])
  );
  //AND U102
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U102 (
    .O(y[239]),
    .I0(a[14]),
    .I1(b[15])
  );
  //OR U102bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U102bar (
    .O(ybar[239]),
    .I0(abar[14]),
    .I1(bbar[15])
  );
  //AND U103
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U103 (
    .O(y[238]),
    .I0(a[14]),
    .I1(b[14])
  );
  //OR U103bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U103bar (
    .O(ybar[238]),
    .I0(abar[14]),
    .I1(bbar[14])
  );
  //AND U104
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U104 (
    .O(y[237]),
    .I0(a[14]),
    .I1(b[13])
  );
  //OR U104bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U104bar (
    .O(ybar[237]),
    .I0(abar[14]),
    .I1(bbar[13])
  );
  //AND U105
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U105 (
    .O(y[236]),
    .I0(a[14]),
    .I1(b[12])
  );
  //OR U105bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U105bar (
    .O(ybar[236]),
    .I0(abar[14]),
    .I1(bbar[12])
  );
  //AND U106
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U106 (
    .O(y[235]),
    .I0(a[14]),
    .I1(b[11])
  );
  //OR U106bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U106bar (
    .O(ybar[235]),
    .I0(abar[14]),
    .I1(bbar[11])
  );
  //AND U107
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U107 (
    .O(y[234]),
    .I0(a[14]),
    .I1(b[10])
  );
  //OR U107bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U107bar (
    .O(ybar[234]),
    .I0(abar[14]),
    .I1(bbar[10])
  );
  //AND U108
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U108 (
    .O(y[233]),
    .I0(a[14]),
    .I1(b[9])
  );
  //OR U108bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U108bar (
    .O(ybar[233]),
    .I0(abar[14]),
    .I1(bbar[9])
  );
  //AND U109
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U109 (
    .O(y[232]),
    .I0(a[14]),
    .I1(b[8])
  );
  //OR U109bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U109bar (
    .O(ybar[232]),
    .I0(abar[14]),
    .I1(bbar[8])
  );
  //AND U110
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U110 (
    .O(y[231]),
    .I0(a[14]),
    .I1(b[7])
  );
  //OR U110bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U110bar (
    .O(ybar[231]),
    .I0(abar[14]),
    .I1(bbar[7])
  );
  //AND U111
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U111 (
    .O(y[230]),
    .I0(a[14]),
    .I1(b[6])
  );
  //OR U111bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U111bar (
    .O(ybar[230]),
    .I0(abar[14]),
    .I1(bbar[6])
  );
  //AND U112
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U112 (
    .O(y[22]),
    .I0(a[1]),
    .I1(b[6])
  );
  //OR U112bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U112bar (
    .O(ybar[22]),
    .I0(abar[1]),
    .I1(bbar[6])
  );
  //AND U113
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U113 (
    .O(y[229]),
    .I0(a[14]),
    .I1(b[5])
  );
  //OR U113bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U113bar (
    .O(ybar[229]),
    .I0(abar[14]),
    .I1(bbar[5])
  );
  //AND U114
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U114 (
    .O(y[228]),
    .I0(a[14]),
    .I1(b[4])
  );
  //OR U114bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U114bar (
    .O(ybar[228]),
    .I0(abar[14]),
    .I1(bbar[4])
  );
  //AND U115
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U115 (
    .O(y[227]),
    .I0(a[14]),
    .I1(b[3])
  );
  //OR U115bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U115bar (
    .O(ybar[227]),
    .I0(abar[14]),
    .I1(bbar[3])
  );
  //AND U116
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U116 (
    .O(y[226]),
    .I0(a[14]),
    .I1(b[2])
  );
  //OR U116bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U116bar (
    .O(ybar[226]),
    .I0(abar[14]),
    .I1(bbar[2])
  );
  //AND U117
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U117 (
    .O(y[225]),
    .I0(a[14]),
    .I1(b[1])
  );
  //OR U117bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U117bar (
    .O(ybar[225]),
    .I0(abar[14]),
    .I1(bbar[1])
  );
  //AND U118
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U118 (
    .O(y[224]),
    .I0(a[14]),
    .I1(b[0])
  );
  //OR U118bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U118bar (
    .O(ybar[224]),
    .I0(abar[14]),
    .I1(bbar[0])
  );
  //AND U119
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U119 (
    .O(y[223]),
    .I0(a[13]),
    .I1(b[15])
  );
  //OR U119bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U119bar (
    .O(ybar[223]),
    .I0(abar[13]),
    .I1(bbar[15])
  );
  //AND U120
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U120 (
    .O(y[222]),
    .I0(a[13]),
    .I1(b[14])
  );
  //OR U120bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U120bar (
    .O(ybar[222]),
    .I0(abar[13]),
    .I1(bbar[14])
  );
  //AND U121
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U121 (
    .O(y[221]),
    .I0(a[13]),
    .I1(b[13])
  );
  //OR U121bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U121bar (
    .O(ybar[221]),
    .I0(abar[13]),
    .I1(bbar[13])
  );
  //AND U122
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U122 (
    .O(y[220]),
    .I0(a[13]),
    .I1(b[12])
  );
  //OR U122bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U122bar (
    .O(ybar[220]),
    .I0(abar[13]),
    .I1(bbar[12])
  );
  //AND U123
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U123 (
    .O(y[21]),
    .I0(a[1]),
    .I1(b[5])
  );
  //OR U123bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U123bar (
    .O(ybar[21]),
    .I0(abar[1]),
    .I1(bbar[5])
  );
  //AND U124
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U124 (
    .O(y[219]),
    .I0(a[13]),
    .I1(b[11])
  );
  //OR U124bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U124bar (
    .O(ybar[219]),
    .I0(abar[13]),
    .I1(bbar[11])
  );
  //AND U125
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U125 (
    .O(y[218]),
    .I0(a[13]),
    .I1(b[10])
  );
  //OR U125bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U125bar (
    .O(ybar[218]),
    .I0(abar[13]),
    .I1(bbar[10])
  );
  //AND U126
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U126 (
    .O(y[217]),
    .I0(a[13]),
    .I1(b[9])
  );
  //OR U126bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U126bar (
    .O(ybar[217]),
    .I0(abar[13]),
    .I1(bbar[9])
  );
  //AND U127
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U127 (
    .O(y[216]),
    .I0(a[13]),
    .I1(b[8])
  );
  //OR U127bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U127bar (
    .O(ybar[216]),
    .I0(abar[13]),
    .I1(bbar[8])
  );
  //AND U128
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U128 (
    .O(y[215]),
    .I0(a[13]),
    .I1(b[7])
  );
  //OR U128bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U128bar (
    .O(ybar[215]),
    .I0(abar[13]),
    .I1(bbar[7])
  );
  //AND U129
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U129 (
    .O(y[214]),
    .I0(a[13]),
    .I1(b[6])
  );
  //OR U129bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U129bar (
    .O(ybar[214]),
    .I0(abar[13]),
    .I1(bbar[6])
  );
  //AND U130
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U130 (
    .O(y[213]),
    .I0(a[13]),
    .I1(b[5])
  );
  //OR U130bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U130bar (
    .O(ybar[213]),
    .I0(abar[13]),
    .I1(bbar[5])
  );
  //AND U131
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U131 (
    .O(y[212]),
    .I0(a[13]),
    .I1(b[4])
  );
  //OR U131bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U131bar (
    .O(ybar[212]),
    .I0(abar[13]),
    .I1(bbar[4])
  );
  //AND U132
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U132 (
    .O(y[211]),
    .I0(a[13]),
    .I1(b[3])
  );
  //OR U132bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U132bar (
    .O(ybar[211]),
    .I0(abar[13]),
    .I1(bbar[3])
  );
  //AND U133
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U133 (
    .O(y[210]),
    .I0(a[13]),
    .I1(b[2])
  );
  //OR U133bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U133bar (
    .O(ybar[210]),
    .I0(abar[13]),
    .I1(bbar[2])
  );
  //AND U134
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U134 (
    .O(y[20]),
    .I0(a[1]),
    .I1(b[4])
  );
  //OR U134bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U134bar (
    .O(ybar[20]),
    .I0(abar[1]),
    .I1(bbar[4])
  );
  //AND U135
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U135 (
    .O(y[209]),
    .I0(a[13]),
    .I1(b[1])
  );
  //OR U135bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U135bar (
    .O(ybar[209]),
    .I0(abar[13]),
    .I1(bbar[1])
  );
  //AND U136
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U136 (
    .O(y[208]),
    .I0(a[13]),
    .I1(b[0])
  );
  //OR U136bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U136bar (
    .O(ybar[208]),
    .I0(abar[13]),
    .I1(bbar[0])
  );
  //AND U137
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U137 (
    .O(y[207]),
    .I0(a[12]),
    .I1(b[15])
  );
  //OR U137bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U137bar (
    .O(ybar[207]),
    .I0(abar[12]),
    .I1(bbar[15])
  );
  //AND U138
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U138 (
    .O(y[206]),
    .I0(a[12]),
    .I1(b[14])
  );
  //OR U138bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U138bar (
    .O(ybar[206]),
    .I0(abar[12]),
    .I1(bbar[14])
  );
  //AND U139
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U139 (
    .O(y[205]),
    .I0(a[12]),
    .I1(b[13])
  );
  //OR U139bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U139bar (
    .O(ybar[205]),
    .I0(abar[12]),
    .I1(bbar[13])
  );
  //AND U140
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U140 (
    .O(y[204]),
    .I0(a[12]),
    .I1(b[12])
  );
  //OR U140bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U140bar (
    .O(ybar[204]),
    .I0(abar[12]),
    .I1(bbar[12])
  );
  //AND U141
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U141 (
    .O(y[203]),
    .I0(a[12]),
    .I1(b[11])
  );
  //OR U141bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U141bar (
    .O(ybar[203]),
    .I0(abar[12]),
    .I1(bbar[11])
  );
  //AND U142
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U142 (
    .O(y[202]),
    .I0(a[12]),
    .I1(b[10])
  );
  //OR U142bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U142bar (
    .O(ybar[202]),
    .I0(abar[12]),
    .I1(bbar[10])
  );
  //AND U143
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U143 (
    .O(y[201]),
    .I0(a[12]),
    .I1(b[9])
  );
  //OR U143bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U143bar (
    .O(ybar[201]),
    .I0(abar[12]),
    .I1(bbar[9])
  );
  //AND U144
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U144 (
    .O(y[200]),
    .I0(a[12]),
    .I1(b[8])
  );
  //OR U144bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U144bar (
    .O(ybar[200]),
    .I0(abar[12]),
    .I1(bbar[8])
  );
  //AND U145
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U145 (
    .O(y[1]),
    .I0(b[1]),
    .I1(a[0])
  );
  //OR U145bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U145bar (
    .O(ybar[1]),
    .I0(bbar[1]),
    .I1(abar[0])
  );
  //AND U146
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U146 (
    .O(y[19]),
    .I0(a[1]),
    .I1(b[3])
  );
  //OR U146bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U146bar (
    .O(ybar[19]),
    .I0(abar[1]),
    .I1(bbar[3])
  );
  //AND U147
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U147 (
    .O(y[199]),
    .I0(a[12]),
    .I1(b[7])
  );
  //OR U147bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U147bar (
    .O(ybar[199]),
    .I0(abar[12]),
    .I1(bbar[7])
  );
  //AND U148
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U148 (
    .O(y[198]),
    .I0(a[12]),
    .I1(b[6])
  );
  //OR U148bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U148bar (
    .O(ybar[198]),
    .I0(abar[12]),
    .I1(bbar[6])
  );
  //AND U149
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U149 (
    .O(y[197]),
    .I0(a[12]),
    .I1(b[5])
  );
  //OR U149bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U149bar (
    .O(ybar[197]),
    .I0(abar[12]),
    .I1(bbar[5])
  );
  //AND U150
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U150 (
    .O(y[196]),
    .I0(a[12]),
    .I1(b[4])
  );
  //OR U150bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U150bar (
    .O(ybar[196]),
    .I0(abar[12]),
    .I1(bbar[4])
  );
  //AND U151
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U151 (
    .O(y[195]),
    .I0(a[12]),
    .I1(b[3])
  );
  //OR U151bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U151bar (
    .O(ybar[195]),
    .I0(abar[12]),
    .I1(bbar[3])
  );
  //AND U152
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U152 (
    .O(y[194]),
    .I0(a[12]),
    .I1(b[2])
  );
  //OR U152bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U152bar (
    .O(ybar[194]),
    .I0(abar[12]),
    .I1(bbar[2])
  );
  //AND U153
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U153 (
    .O(y[193]),
    .I0(a[12]),
    .I1(b[1])
  );
  //OR U153bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U153bar (
    .O(ybar[193]),
    .I0(abar[12]),
    .I1(bbar[1])
  );
  //AND U154
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U154 (
    .O(y[192]),
    .I0(a[12]),
    .I1(b[0])
  );
  //OR U154bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U154bar (
    .O(ybar[192]),
    .I0(abar[12]),
    .I1(bbar[0])
  );
  //AND U155
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U155 (
    .O(y[191]),
    .I0(a[11]),
    .I1(b[15])
  );
  //OR U155bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U155bar (
    .O(ybar[191]),
    .I0(abar[11]),
    .I1(bbar[15])
  );
  //AND U156
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U156 (
    .O(y[190]),
    .I0(a[11]),
    .I1(b[14])
  );
  //OR U156bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U156bar (
    .O(ybar[190]),
    .I0(abar[11]),
    .I1(bbar[14])
  );
  //AND U157
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U157 (
    .O(y[18]),
    .I0(a[1]),
    .I1(b[2])
  );
  //OR U157bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U157bar (
    .O(ybar[18]),
    .I0(abar[1]),
    .I1(bbar[2])
  );
  //AND U158
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U158 (
    .O(y[189]),
    .I0(a[11]),
    .I1(b[13])
  );
  //OR U158bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U158bar (
    .O(ybar[189]),
    .I0(abar[11]),
    .I1(bbar[13])
  );
  //AND U159
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U159 (
    .O(y[188]),
    .I0(a[11]),
    .I1(b[12])
  );
  //OR U159bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U159bar (
    .O(ybar[188]),
    .I0(abar[11]),
    .I1(bbar[12])
  );
  //AND U160
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U160 (
    .O(y[187]),
    .I0(a[11]),
    .I1(b[11])
  );
  //OR U160bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U160bar (
    .O(ybar[187]),
    .I0(abar[11]),
    .I1(bbar[11])
  );
  //AND U161
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U161 (
    .O(y[186]),
    .I0(a[11]),
    .I1(b[10])
  );
  //OR U161bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U161bar (
    .O(ybar[186]),
    .I0(abar[11]),
    .I1(bbar[10])
  );
  //AND U162
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U162 (
    .O(y[185]),
    .I0(a[11]),
    .I1(b[9])
  );
  //OR U162bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U162bar (
    .O(ybar[185]),
    .I0(abar[11]),
    .I1(bbar[9])
  );
  //AND U163
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U163 (
    .O(y[184]),
    .I0(a[11]),
    .I1(b[8])
  );
  //OR U163bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U163bar (
    .O(ybar[184]),
    .I0(abar[11]),
    .I1(bbar[8])
  );
  //AND U164
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U164 (
    .O(y[183]),
    .I0(a[11]),
    .I1(b[7])
  );
  //OR U164bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U164bar (
    .O(ybar[183]),
    .I0(abar[11]),
    .I1(bbar[7])
  );
  //AND U165
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U165 (
    .O(y[182]),
    .I0(a[11]),
    .I1(b[6])
  );
  //OR U165bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U165bar (
    .O(ybar[182]),
    .I0(abar[11]),
    .I1(bbar[6])
  );
  //AND U166
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U166 (
    .O(y[181]),
    .I0(a[11]),
    .I1(b[5])
  );
  //OR U166bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U166bar (
    .O(ybar[181]),
    .I0(abar[11]),
    .I1(bbar[5])
  );
  //AND U167
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U167 (
    .O(y[180]),
    .I0(a[11]),
    .I1(b[4])
  );
  //OR U167bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U167bar (
    .O(ybar[180]),
    .I0(abar[11]),
    .I1(bbar[4])
  );
  //AND U168
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U168 (
    .O(y[17]),
    .I0(a[1]),
    .I1(b[1])
  );
  //OR U168bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U168bar (
    .O(ybar[17]),
    .I0(abar[1]),
    .I1(bbar[1])
  );
  //AND U169
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U169 (
    .O(y[179]),
    .I0(a[11]),
    .I1(b[3])
  );
  //OR U169bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U169bar (
    .O(ybar[179]),
    .I0(abar[11]),
    .I1(bbar[3])
  );
  //AND U170
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U170 (
    .O(y[178]),
    .I0(a[11]),
    .I1(b[2])
  );
  //OR U170bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U170bar (
    .O(ybar[178]),
    .I0(abar[11]),
    .I1(bbar[2])
  );
  //AND U171
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U171 (
    .O(y[177]),
    .I0(a[11]),
    .I1(b[1])
  );
  //OR U171bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U171bar (
    .O(ybar[177]),
    .I0(abar[11]),
    .I1(bbar[1])
  );
  //AND U172
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U172 (
    .O(y[176]),
    .I0(a[11]),
    .I1(b[0])
  );
  //OR U172bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U172bar (
    .O(ybar[176]),
    .I0(abar[11]),
    .I1(bbar[0])
  );
  //AND U173
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U173 (
    .O(y[175]),
    .I0(a[10]),
    .I1(b[15])
  );
  //OR U173bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U173bar (
    .O(ybar[175]),
    .I0(abar[10]),
    .I1(bbar[15])
  );
  //AND U174
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U174 (
    .O(y[174]),
    .I0(a[10]),
    .I1(b[14])
  );
  //OR U174bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U174bar (
    .O(ybar[174]),
    .I0(abar[10]),
    .I1(bbar[14])
  );
  //AND U175
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U175 (
    .O(y[173]),
    .I0(a[10]),
    .I1(b[13])
  );
  //OR U175bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U175bar (
    .O(ybar[173]),
    .I0(abar[10]),
    .I1(bbar[13])
  );
  //AND U176
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U176 (
    .O(y[172]),
    .I0(a[10]),
    .I1(b[12])
  );
  //OR U176bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U176bar (
    .O(ybar[172]),
    .I0(abar[10]),
    .I1(bbar[12])
  );
  //AND U177
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U177 (
    .O(y[171]),
    .I0(a[10]),
    .I1(b[11])
  );
  //OR U177bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U177bar (
    .O(ybar[171]),
    .I0(abar[10]),
    .I1(bbar[11])
  );
  //AND U178
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U178 (
    .O(y[170]),
    .I0(a[10]),
    .I1(b[10])
  );
  //OR U178bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U178bar (
    .O(ybar[170]),
    .I0(abar[10]),
    .I1(bbar[10])
  );
  //AND U179
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U179 (
    .O(y[16]),
    .I0(a[1]),
    .I1(b[0])
  );
  //OR U179bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U179bar (
    .O(ybar[16]),
    .I0(abar[1]),
    .I1(bbar[0])
  );
  //AND U180
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U180 (
    .O(y[169]),
    .I0(a[10]),
    .I1(b[9])
  );
  //OR U180bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U180bar (
    .O(ybar[169]),
    .I0(abar[10]),
    .I1(bbar[9])
  );
  //AND U181
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U181 (
    .O(y[168]),
    .I0(a[10]),
    .I1(b[8])
  );
  //OR U181bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U181bar (
    .O(ybar[168]),
    .I0(abar[10]),
    .I1(bbar[8])
  );
  //AND U182
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U182 (
    .O(y[167]),
    .I0(a[10]),
    .I1(b[7])
  );
  //OR U182bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U182bar (
    .O(ybar[167]),
    .I0(abar[10]),
    .I1(bbar[7])
  );
  //AND U183
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U183 (
    .O(y[166]),
    .I0(a[10]),
    .I1(b[6])
  );
  //OR U183bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U183bar (
    .O(ybar[166]),
    .I0(abar[10]),
    .I1(bbar[6])
  );
  //AND U184
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U184 (
    .O(y[165]),
    .I0(a[10]),
    .I1(b[5])
  );
  //OR U184bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U184bar (
    .O(ybar[165]),
    .I0(abar[10]),
    .I1(bbar[5])
  );
  //AND U185
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U185 (
    .O(y[164]),
    .I0(a[10]),
    .I1(b[4])
  );
  //OR U185bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U185bar (
    .O(ybar[164]),
    .I0(abar[10]),
    .I1(bbar[4])
  );
  //AND U186
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U186 (
    .O(y[163]),
    .I0(a[10]),
    .I1(b[3])
  );
  //OR U186bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U186bar (
    .O(ybar[163]),
    .I0(abar[10]),
    .I1(bbar[3])
  );
  //AND U187
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U187 (
    .O(y[162]),
    .I0(a[10]),
    .I1(b[2])
  );
  //OR U187bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U187bar (
    .O(ybar[162]),
    .I0(abar[10]),
    .I1(bbar[2])
  );
  //AND U188
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U188 (
    .O(y[161]),
    .I0(a[10]),
    .I1(b[1])
  );
  //OR U188bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U188bar (
    .O(ybar[161]),
    .I0(abar[10]),
    .I1(bbar[1])
  );
  //AND U189
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U189 (
    .O(y[160]),
    .I0(a[10]),
    .I1(b[0])
  );
  //OR U189bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U189bar (
    .O(ybar[160]),
    .I0(abar[10]),
    .I1(bbar[0])
  );
  //AND U190
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U190 (
    .O(y[15]),
    .I0(b[15]),
    .I1(a[0])
  );
  //OR U190bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U190bar (
    .O(ybar[15]),
    .I0(bbar[15]),
    .I1(abar[0])
  );
  //AND U191
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U191 (
    .O(y[159]),
    .I0(a[9]),
    .I1(b[15])
  );
  //OR U191bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U191bar (
    .O(ybar[159]),
    .I0(abar[9]),
    .I1(bbar[15])
  );
  //AND U192
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U192 (
    .O(y[158]),
    .I0(a[9]),
    .I1(b[14])
  );
  //OR U192bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U192bar (
    .O(ybar[158]),
    .I0(abar[9]),
    .I1(bbar[14])
  );
  //AND U193
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U193 (
    .O(y[157]),
    .I0(a[9]),
    .I1(b[13])
  );
  //OR U193bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U193bar (
    .O(ybar[157]),
    .I0(abar[9]),
    .I1(bbar[13])
  );
  //AND U194
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U194 (
    .O(y[156]),
    .I0(a[9]),
    .I1(b[12])
  );
  //OR U194bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U194bar (
    .O(ybar[156]),
    .I0(abar[9]),
    .I1(bbar[12])
  );
  //AND U195
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U195 (
    .O(y[155]),
    .I0(a[9]),
    .I1(b[11])
  );
  //OR U195bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U195bar (
    .O(ybar[155]),
    .I0(abar[9]),
    .I1(bbar[11])
  );
  //AND U196
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U196 (
    .O(y[154]),
    .I0(a[9]),
    .I1(b[10])
  );
  //OR U196bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U196bar (
    .O(ybar[154]),
    .I0(abar[9]),
    .I1(bbar[10])
  );
  //AND U197
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U197 (
    .O(y[153]),
    .I0(a[9]),
    .I1(b[9])
  );
  //OR U197bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U197bar (
    .O(ybar[153]),
    .I0(abar[9]),
    .I1(bbar[9])
  );
  //AND U198
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U198 (
    .O(y[152]),
    .I0(a[9]),
    .I1(b[8])
  );
  //OR U198bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U198bar (
    .O(ybar[152]),
    .I0(abar[9]),
    .I1(bbar[8])
  );
  //AND U199
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U199 (
    .O(y[151]),
    .I0(a[9]),
    .I1(b[7])
  );
  //OR U199bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U199bar (
    .O(ybar[151]),
    .I0(abar[9]),
    .I1(bbar[7])
  );
  //AND U200
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U200 (
    .O(y[150]),
    .I0(a[9]),
    .I1(b[6])
  );
  //OR U200bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U200bar (
    .O(ybar[150]),
    .I0(abar[9]),
    .I1(bbar[6])
  );
  //AND U201
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U201 (
    .O(y[14]),
    .I0(b[14]),
    .I1(a[0])
  );
  //OR U201bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U201bar (
    .O(ybar[14]),
    .I0(bbar[14]),
    .I1(abar[0])
  );
  //AND U202
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U202 (
    .O(y[149]),
    .I0(a[9]),
    .I1(b[5])
  );
  //OR U202bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U202bar (
    .O(ybar[149]),
    .I0(abar[9]),
    .I1(bbar[5])
  );
  //AND U203
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U203 (
    .O(y[148]),
    .I0(a[9]),
    .I1(b[4])
  );
  //OR U203bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U203bar (
    .O(ybar[148]),
    .I0(abar[9]),
    .I1(bbar[4])
  );
  //AND U204
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U204 (
    .O(y[147]),
    .I0(a[9]),
    .I1(b[3])
  );
  //OR U204bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U204bar (
    .O(ybar[147]),
    .I0(abar[9]),
    .I1(bbar[3])
  );
  //AND U205
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U205 (
    .O(y[146]),
    .I0(a[9]),
    .I1(b[2])
  );
  //OR U205bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U205bar (
    .O(ybar[146]),
    .I0(abar[9]),
    .I1(bbar[2])
  );
  //AND U206
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U206 (
    .O(y[145]),
    .I0(a[9]),
    .I1(b[1])
  );
  //OR U206bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U206bar (
    .O(ybar[145]),
    .I0(abar[9]),
    .I1(bbar[1])
  );
  //AND U207
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U207 (
    .O(y[144]),
    .I0(a[9]),
    .I1(b[0])
  );
  //OR U207bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U207bar (
    .O(ybar[144]),
    .I0(abar[9]),
    .I1(bbar[0])
  );
  //AND U208
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U208 (
    .O(y[143]),
    .I0(a[8]),
    .I1(b[15])
  );
  //OR U208bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U208bar (
    .O(ybar[143]),
    .I0(abar[8]),
    .I1(bbar[15])
  );
  //AND U209
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U209 (
    .O(y[142]),
    .I0(a[8]),
    .I1(b[14])
  );
  //OR U209bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U209bar (
    .O(ybar[142]),
    .I0(abar[8]),
    .I1(bbar[14])
  );
  //AND U210
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U210 (
    .O(y[141]),
    .I0(a[8]),
    .I1(b[13])
  );
  //OR U210bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U210bar (
    .O(ybar[141]),
    .I0(abar[8]),
    .I1(bbar[13])
  );
  //AND U211
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U211 (
    .O(y[140]),
    .I0(a[8]),
    .I1(b[12])
  );
  //OR U211bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U211bar (
    .O(ybar[140]),
    .I0(abar[8]),
    .I1(bbar[12])
  );
  //AND U212
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U212 (
    .O(y[13]),
    .I0(b[13]),
    .I1(a[0])
  );
  //OR U212bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U212bar (
    .O(ybar[13]),
    .I0(bbar[13]),
    .I1(abar[0])
  );
  //AND U213
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U213 (
    .O(y[139]),
    .I0(a[8]),
    .I1(b[11])
  );
  //OR U213bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U213bar (
    .O(ybar[139]),
    .I0(abar[8]),
    .I1(bbar[11])
  );
  //AND U214
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U214 (
    .O(y[138]),
    .I0(a[8]),
    .I1(b[10])
  );
  //OR U214bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U214bar (
    .O(ybar[138]),
    .I0(abar[8]),
    .I1(bbar[10])
  );
  //AND U215
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U215 (
    .O(y[137]),
    .I0(a[8]),
    .I1(b[9])
  );
  //OR U215bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U215bar (
    .O(ybar[137]),
    .I0(abar[8]),
    .I1(bbar[9])
  );
  //AND U216
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U216 (
    .O(y[136]),
    .I0(a[8]),
    .I1(b[8])
  );
  //OR U216bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U216bar (
    .O(ybar[136]),
    .I0(abar[8]),
    .I1(bbar[8])
  );
  //AND U217
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U217 (
    .O(y[135]),
    .I0(a[8]),
    .I1(b[7])
  );
  //OR U217bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U217bar (
    .O(ybar[135]),
    .I0(abar[8]),
    .I1(bbar[7])
  );
  //AND U218
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U218 (
    .O(y[134]),
    .I0(a[8]),
    .I1(b[6])
  );
  //OR U218bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U218bar (
    .O(ybar[134]),
    .I0(abar[8]),
    .I1(bbar[6])
  );
  //AND U219
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U219 (
    .O(y[133]),
    .I0(a[8]),
    .I1(b[5])
  );
  //OR U219bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U219bar (
    .O(ybar[133]),
    .I0(abar[8]),
    .I1(bbar[5])
  );
  //AND U220
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U220 (
    .O(y[132]),
    .I0(a[8]),
    .I1(b[4])
  );
  //OR U220bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U220bar (
    .O(ybar[132]),
    .I0(abar[8]),
    .I1(bbar[4])
  );
  //AND U221
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U221 (
    .O(y[131]),
    .I0(a[8]),
    .I1(b[3])
  );
  //OR U221bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U221bar (
    .O(ybar[131]),
    .I0(abar[8]),
    .I1(bbar[3])
  );
  //AND U222
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U222 (
    .O(y[130]),
    .I0(a[8]),
    .I1(b[2])
  );
  //OR U222bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U222bar (
    .O(ybar[130]),
    .I0(abar[8]),
    .I1(bbar[2])
  );
  //AND U223
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U223 (
    .O(y[12]),
    .I0(b[12]),
    .I1(a[0])
  );
  //OR U223bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U223bar (
    .O(ybar[12]),
    .I0(bbar[12]),
    .I1(abar[0])
  );
  //AND U224
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U224 (
    .O(y[129]),
    .I0(a[8]),
    .I1(b[1])
  );
  //OR U224bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U224bar (
    .O(ybar[129]),
    .I0(abar[8]),
    .I1(bbar[1])
  );
  //AND U225
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U225 (
    .O(y[128]),
    .I0(a[8]),
    .I1(b[0])
  );
  //OR U225bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U225bar (
    .O(ybar[128]),
    .I0(abar[8]),
    .I1(bbar[0])
  );
  //AND U226
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U226 (
    .O(y[127]),
    .I0(a[7]),
    .I1(b[15])
  );
  //OR U226bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U226bar (
    .O(ybar[127]),
    .I0(abar[7]),
    .I1(bbar[15])
  );
  //AND U227
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U227 (
    .O(y[126]),
    .I0(a[7]),
    .I1(b[14])
  );
  //OR U227bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U227bar (
    .O(ybar[126]),
    .I0(abar[7]),
    .I1(bbar[14])
  );
  //AND U228
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U228 (
    .O(y[125]),
    .I0(a[7]),
    .I1(b[13])
  );
  //OR U228bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U228bar (
    .O(ybar[125]),
    .I0(abar[7]),
    .I1(bbar[13])
  );
  //AND U229
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U229 (
    .O(y[124]),
    .I0(a[7]),
    .I1(b[12])
  );
  //OR U229bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U229bar (
    .O(ybar[124]),
    .I0(abar[7]),
    .I1(bbar[12])
  );
  //AND U230
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U230 (
    .O(y[123]),
    .I0(a[7]),
    .I1(b[11])
  );
  //OR U230bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U230bar (
    .O(ybar[123]),
    .I0(abar[7]),
    .I1(bbar[11])
  );
  //AND U231
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U231 (
    .O(y[122]),
    .I0(a[7]),
    .I1(b[10])
  );
  //OR U231bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U231bar (
    .O(ybar[122]),
    .I0(abar[7]),
    .I1(bbar[10])
  );
  //AND U232
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U232 (
    .O(y[121]),
    .I0(a[7]),
    .I1(b[9])
  );
  //OR U232bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U232bar (
    .O(ybar[121]),
    .I0(abar[7]),
    .I1(bbar[9])
  );
  //AND U233
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U233 (
    .O(y[120]),
    .I0(a[7]),
    .I1(b[8])
  );
  //OR U233bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U233bar (
    .O(ybar[120]),
    .I0(abar[7]),
    .I1(bbar[8])
  );
  //AND U234
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U234 (
    .O(y[11]),
    .I0(b[11]),
    .I1(a[0])
  );
  //OR U234bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U234bar (
    .O(ybar[11]),
    .I0(bbar[11]),
    .I1(abar[0])
  );
  //AND U235
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U235 (
    .O(y[119]),
    .I0(a[7]),
    .I1(b[7])
  );
  //OR U235bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U235bar (
    .O(ybar[119]),
    .I0(abar[7]),
    .I1(bbar[7])
  );
  //AND U236
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U236 (
    .O(y[118]),
    .I0(a[7]),
    .I1(b[6])
  );
  //OR U236bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U236bar (
    .O(ybar[118]),
    .I0(abar[7]),
    .I1(bbar[6])
  );
  //AND U237
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U237 (
    .O(y[117]),
    .I0(a[7]),
    .I1(b[5])
  );
  //OR U237bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U237bar (
    .O(ybar[117]),
    .I0(abar[7]),
    .I1(bbar[5])
  );
  //AND U238
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U238 (
    .O(y[116]),
    .I0(a[7]),
    .I1(b[4])
  );
  //OR U238bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U238bar (
    .O(ybar[116]),
    .I0(abar[7]),
    .I1(bbar[4])
  );
  //AND U239
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U239 (
    .O(y[115]),
    .I0(a[7]),
    .I1(b[3])
  );
  //OR U239bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U239bar (
    .O(ybar[115]),
    .I0(abar[7]),
    .I1(bbar[3])
  );
  //AND U240
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U240 (
    .O(y[114]),
    .I0(a[7]),
    .I1(b[2])
  );
  //OR U240bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U240bar (
    .O(ybar[114]),
    .I0(abar[7]),
    .I1(bbar[2])
  );
  //AND U241
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U241 (
    .O(y[113]),
    .I0(a[7]),
    .I1(b[1])
  );
  //OR U241bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U241bar (
    .O(ybar[113]),
    .I0(abar[7]),
    .I1(bbar[1])
  );
  //AND U242
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U242 (
    .O(y[112]),
    .I0(a[7]),
    .I1(b[0])
  );
  //OR U242bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U242bar (
    .O(ybar[112]),
    .I0(abar[7]),
    .I1(bbar[0])
  );
  //AND U243
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U243 (
    .O(y[111]),
    .I0(b[15]),
    .I1(a[6])
  );
  //OR U243bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U243bar (
    .O(ybar[111]),
    .I0(bbar[15]),
    .I1(abar[6])
  );
  //AND U244
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U244 (
    .O(y[110]),
    .I0(b[14]),
    .I1(a[6])
  );
  //OR U244bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U244bar (
    .O(ybar[110]),
    .I0(bbar[14]),
    .I1(abar[6])
  );
  //AND U245
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U245 (
    .O(y[10]),
    .I0(b[10]),
    .I1(a[0])
  );
  //OR U245bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U245bar (
    .O(ybar[10]),
    .I0(bbar[10]),
    .I1(abar[0])
  );
  //AND U246
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U246 (
    .O(y[109]),
    .I0(b[13]),
    .I1(a[6])
  );
  //OR U246bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U246bar (
    .O(ybar[109]),
    .I0(bbar[13]),
    .I1(abar[6])
  );
  //AND U247
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U247 (
    .O(y[108]),
    .I0(b[12]),
    .I1(a[6])
  );
  //OR U247bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U247bar (
    .O(ybar[108]),
    .I0(bbar[12]),
    .I1(abar[6])
  );
  //AND U248
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U248 (
    .O(y[107]),
    .I0(b[11]),
    .I1(a[6])
  );
  //OR U248bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U248bar (
    .O(ybar[107]),
    .I0(bbar[11]),
    .I1(abar[6])
  );
  //AND U249
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U249 (
    .O(y[106]),
    .I0(b[10]),
    .I1(a[6])
  );
  //OR U249bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U249bar (
    .O(ybar[106]),
    .I0(bbar[10]),
    .I1(abar[6])
  );
  //AND U250
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U250 (
    .O(y[105]),
    .I0(a[6]),
    .I1(b[9])
  );
  //OR U250bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U250bar (
    .O(ybar[105]),
    .I0(abar[6]),
    .I1(bbar[9])
  );
  //AND U251
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U251 (
    .O(y[104]),
    .I0(b[8]),
    .I1(a[6])
  );
  //OR U251bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U251bar (
    .O(ybar[104]),
    .I0(bbar[8]),
    .I1(abar[6])
  );
  //AND U252
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U252 (
    .O(y[103]),
    .I0(b[7]),
    .I1(a[6])
  );
  //OR U252bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U252bar (
    .O(ybar[103]),
    .I0(bbar[7]),
    .I1(abar[6])
  );
  //AND U253
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U253 (
    .O(y[102]),
    .I0(b[6]),
    .I1(a[6])
  );
  //OR U253bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U253bar (
    .O(ybar[102]),
    .I0(bbar[6]),
    .I1(abar[6])
  );
  //AND U254
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U254 (
    .O(y[101]),
    .I0(b[5]),
    .I1(a[6])
  );
  //OR U254bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U254bar (
    .O(ybar[101]),
    .I0(bbar[5]),
    .I1(abar[6])
  );
  //AND U255
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U255 (
    .O(y[100]),
    .I0(b[4]),
    .I1(a[6])
  );
  //OR U255bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U255bar (
    .O(ybar[100]),
    .I0(bbar[4]),
    .I1(abar[6])
  );
  //AND U256
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U256 (
    .O(y[0]),
    .I0(b[0]),
    .I1(a[0])
  );
  //OR U256bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U256bar (
    .O(ybar[0]),
    .I0(bbar[0]),
    .I1(abar[0])
  );
endmodule

module decode_15 ( in, out );

  input wire [7:0] in;
//input_done

  output wire [255:0] out;
//output_done

  wire [15:0] level1;
  wire [31:0] level2;
//wire_done

  CD2_60 cd_l1_1 ( .a(in[1]), .b(in[0]), .y(level1[3:0]) );
  CD2_59 cd_l1_2 ( .a(in[3]), .b(in[2]), .y(level1[7:4]) );
  CD2_58 cd_l1_3 ( .a(in[5]), .b(in[4]), .y(level1[11:8]) );
  CD2_57 cd_l1_4 ( .a(in[7]), .b(in[6]), .y(level1[15:12]) );
  CD4_30 cd_l2_1 ( .a(level1[7:4]), .b(level1[3:0]), .y(level2[15:0]) );
  CD4_29 cd_l2_2 ( .a(level1[15:12]), .b(level1[11:8]), .y(level2[31:16]) );
  CD16_15 cd_l3 ( .a(level2[31:16]), .b(level2[15:0]), .y(out) );
endmodule

module encode_15 ( in, out );

  input wire [255:0] in;
  wire [255:0] inbar;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
  assign inbar[8] = ~in[8];
  assign inbar[9] = ~in[9];
  assign inbar[10] = ~in[10];
  assign inbar[11] = ~in[11];
  assign inbar[12] = ~in[12];
  assign inbar[13] = ~in[13];
  assign inbar[14] = ~in[14];
  assign inbar[15] = ~in[15];
  assign inbar[16] = ~in[16];
  assign inbar[17] = ~in[17];
  assign inbar[18] = ~in[18];
  assign inbar[19] = ~in[19];
  assign inbar[20] = ~in[20];
  assign inbar[21] = ~in[21];
  assign inbar[22] = ~in[22];
  assign inbar[23] = ~in[23];
  assign inbar[24] = ~in[24];
  assign inbar[25] = ~in[25];
  assign inbar[26] = ~in[26];
  assign inbar[27] = ~in[27];
  assign inbar[28] = ~in[28];
  assign inbar[29] = ~in[29];
  assign inbar[30] = ~in[30];
  assign inbar[31] = ~in[31];
  assign inbar[32] = ~in[32];
  assign inbar[33] = ~in[33];
  assign inbar[34] = ~in[34];
  assign inbar[35] = ~in[35];
  assign inbar[36] = ~in[36];
  assign inbar[37] = ~in[37];
  assign inbar[38] = ~in[38];
  assign inbar[39] = ~in[39];
  assign inbar[40] = ~in[40];
  assign inbar[41] = ~in[41];
  assign inbar[42] = ~in[42];
  assign inbar[43] = ~in[43];
  assign inbar[44] = ~in[44];
  assign inbar[45] = ~in[45];
  assign inbar[46] = ~in[46];
  assign inbar[47] = ~in[47];
  assign inbar[48] = ~in[48];
  assign inbar[49] = ~in[49];
  assign inbar[50] = ~in[50];
  assign inbar[51] = ~in[51];
  assign inbar[52] = ~in[52];
  assign inbar[53] = ~in[53];
  assign inbar[54] = ~in[54];
  assign inbar[55] = ~in[55];
  assign inbar[56] = ~in[56];
  assign inbar[57] = ~in[57];
  assign inbar[58] = ~in[58];
  assign inbar[59] = ~in[59];
  assign inbar[60] = ~in[60];
  assign inbar[61] = ~in[61];
  assign inbar[62] = ~in[62];
  assign inbar[63] = ~in[63];
  assign inbar[64] = ~in[64];
  assign inbar[65] = ~in[65];
  assign inbar[66] = ~in[66];
  assign inbar[67] = ~in[67];
  assign inbar[68] = ~in[68];
  assign inbar[69] = ~in[69];
  assign inbar[70] = ~in[70];
  assign inbar[71] = ~in[71];
  assign inbar[72] = ~in[72];
  assign inbar[73] = ~in[73];
  assign inbar[74] = ~in[74];
  assign inbar[75] = ~in[75];
  assign inbar[76] = ~in[76];
  assign inbar[77] = ~in[77];
  assign inbar[78] = ~in[78];
  assign inbar[79] = ~in[79];
  assign inbar[80] = ~in[80];
  assign inbar[81] = ~in[81];
  assign inbar[82] = ~in[82];
  assign inbar[83] = ~in[83];
  assign inbar[84] = ~in[84];
  assign inbar[85] = ~in[85];
  assign inbar[86] = ~in[86];
  assign inbar[87] = ~in[87];
  assign inbar[88] = ~in[88];
  assign inbar[89] = ~in[89];
  assign inbar[90] = ~in[90];
  assign inbar[91] = ~in[91];
  assign inbar[92] = ~in[92];
  assign inbar[93] = ~in[93];
  assign inbar[94] = ~in[94];
  assign inbar[95] = ~in[95];
  assign inbar[96] = ~in[96];
  assign inbar[97] = ~in[97];
  assign inbar[98] = ~in[98];
  assign inbar[99] = ~in[99];
  assign inbar[100] = ~in[100];
  assign inbar[101] = ~in[101];
  assign inbar[102] = ~in[102];
  assign inbar[103] = ~in[103];
  assign inbar[104] = ~in[104];
  assign inbar[105] = ~in[105];
  assign inbar[106] = ~in[106];
  assign inbar[107] = ~in[107];
  assign inbar[108] = ~in[108];
  assign inbar[109] = ~in[109];
  assign inbar[110] = ~in[110];
  assign inbar[111] = ~in[111];
  assign inbar[112] = ~in[112];
  assign inbar[113] = ~in[113];
  assign inbar[114] = ~in[114];
  assign inbar[115] = ~in[115];
  assign inbar[116] = ~in[116];
  assign inbar[117] = ~in[117];
  assign inbar[118] = ~in[118];
  assign inbar[119] = ~in[119];
  assign inbar[120] = ~in[120];
  assign inbar[121] = ~in[121];
  assign inbar[122] = ~in[122];
  assign inbar[123] = ~in[123];
  assign inbar[124] = ~in[124];
  assign inbar[125] = ~in[125];
  assign inbar[126] = ~in[126];
  assign inbar[127] = ~in[127];
  assign inbar[128] = ~in[128];
  assign inbar[129] = ~in[129];
  assign inbar[130] = ~in[130];
  assign inbar[131] = ~in[131];
  assign inbar[132] = ~in[132];
  assign inbar[133] = ~in[133];
  assign inbar[134] = ~in[134];
  assign inbar[135] = ~in[135];
  assign inbar[136] = ~in[136];
  assign inbar[137] = ~in[137];
  assign inbar[138] = ~in[138];
  assign inbar[139] = ~in[139];
  assign inbar[140] = ~in[140];
  assign inbar[141] = ~in[141];
  assign inbar[142] = ~in[142];
  assign inbar[143] = ~in[143];
  assign inbar[144] = ~in[144];
  assign inbar[145] = ~in[145];
  assign inbar[146] = ~in[146];
  assign inbar[147] = ~in[147];
  assign inbar[148] = ~in[148];
  assign inbar[149] = ~in[149];
  assign inbar[150] = ~in[150];
  assign inbar[151] = ~in[151];
  assign inbar[152] = ~in[152];
  assign inbar[153] = ~in[153];
  assign inbar[154] = ~in[154];
  assign inbar[155] = ~in[155];
  assign inbar[156] = ~in[156];
  assign inbar[157] = ~in[157];
  assign inbar[158] = ~in[158];
  assign inbar[159] = ~in[159];
  assign inbar[160] = ~in[160];
  assign inbar[161] = ~in[161];
  assign inbar[162] = ~in[162];
  assign inbar[163] = ~in[163];
  assign inbar[164] = ~in[164];
  assign inbar[165] = ~in[165];
  assign inbar[166] = ~in[166];
  assign inbar[167] = ~in[167];
  assign inbar[168] = ~in[168];
  assign inbar[169] = ~in[169];
  assign inbar[170] = ~in[170];
  assign inbar[171] = ~in[171];
  assign inbar[172] = ~in[172];
  assign inbar[173] = ~in[173];
  assign inbar[174] = ~in[174];
  assign inbar[175] = ~in[175];
  assign inbar[176] = ~in[176];
  assign inbar[177] = ~in[177];
  assign inbar[178] = ~in[178];
  assign inbar[179] = ~in[179];
  assign inbar[180] = ~in[180];
  assign inbar[181] = ~in[181];
  assign inbar[182] = ~in[182];
  assign inbar[183] = ~in[183];
  assign inbar[184] = ~in[184];
  assign inbar[185] = ~in[185];
  assign inbar[186] = ~in[186];
  assign inbar[187] = ~in[187];
  assign inbar[188] = ~in[188];
  assign inbar[189] = ~in[189];
  assign inbar[190] = ~in[190];
  assign inbar[191] = ~in[191];
  assign inbar[192] = ~in[192];
  assign inbar[193] = ~in[193];
  assign inbar[194] = ~in[194];
  assign inbar[195] = ~in[195];
  assign inbar[196] = ~in[196];
  assign inbar[197] = ~in[197];
  assign inbar[198] = ~in[198];
  assign inbar[199] = ~in[199];
  assign inbar[200] = ~in[200];
  assign inbar[201] = ~in[201];
  assign inbar[202] = ~in[202];
  assign inbar[203] = ~in[203];
  assign inbar[204] = ~in[204];
  assign inbar[205] = ~in[205];
  assign inbar[206] = ~in[206];
  assign inbar[207] = ~in[207];
  assign inbar[208] = ~in[208];
  assign inbar[209] = ~in[209];
  assign inbar[210] = ~in[210];
  assign inbar[211] = ~in[211];
  assign inbar[212] = ~in[212];
  assign inbar[213] = ~in[213];
  assign inbar[214] = ~in[214];
  assign inbar[215] = ~in[215];
  assign inbar[216] = ~in[216];
  assign inbar[217] = ~in[217];
  assign inbar[218] = ~in[218];
  assign inbar[219] = ~in[219];
  assign inbar[220] = ~in[220];
  assign inbar[221] = ~in[221];
  assign inbar[222] = ~in[222];
  assign inbar[223] = ~in[223];
  assign inbar[224] = ~in[224];
  assign inbar[225] = ~in[225];
  assign inbar[226] = ~in[226];
  assign inbar[227] = ~in[227];
  assign inbar[228] = ~in[228];
  assign inbar[229] = ~in[229];
  assign inbar[230] = ~in[230];
  assign inbar[231] = ~in[231];
  assign inbar[232] = ~in[232];
  assign inbar[233] = ~in[233];
  assign inbar[234] = ~in[234];
  assign inbar[235] = ~in[235];
  assign inbar[236] = ~in[236];
  assign inbar[237] = ~in[237];
  assign inbar[238] = ~in[238];
  assign inbar[239] = ~in[239];
  assign inbar[240] = ~in[240];
  assign inbar[241] = ~in[241];
  assign inbar[242] = ~in[242];
  assign inbar[243] = ~in[243];
  assign inbar[244] = ~in[244];
  assign inbar[245] = ~in[245];
  assign inbar[246] = ~in[246];
  assign inbar[247] = ~in[247];
  assign inbar[248] = ~in[248];
  assign inbar[249] = ~in[249];
  assign inbar[250] = ~in[250];
  assign inbar[251] = ~in[251];
  assign inbar[252] = ~in[252];
  assign inbar[253] = ~in[253];
  assign inbar[254] = ~in[254];
  assign inbar[255] = ~in[255];
//input_done

  output wire [7:0] out;
  wire [7:0] outbar;
//output_done

  wire in_81;
  wire in_80;
  wire in_79;
  wire in_78;
  wire in_77;
  wire in_76;
  wire in_75;
  wire in_74;
  wire in_73;
  wire in_72;
  wire in_71;
  wire in_70;
  wire in_69;
  wire in_68;
  wire in_67;
  wire in_66;
  wire in_65;
  wire in_64;
  wire in_63;
  wire in_62;
  wire in_61;
  wire in_60;
  wire in_59;
  wire in_58;
  wire in_57;
  wire in_56;
  wire in_55;
  wire in_54;
  wire in_53;
  wire in_52;
  wire in_51;
  wire in_50;
  wire in_49;
  wire in_48;
  wire in_47;
  wire in_46;
  wire in_45;
  wire in_44;
  wire in_43;
  wire in_42;
  wire in_41;
  wire in_40;
  wire in_39;
  wire in_38;
  wire in_37;
  wire in_36;
  wire in_35;
  wire in_34;
  wire in_33;
  wire in_32;
  wire in_31;
  wire in_30;
  wire in_29;
  wire in_28;
  wire in_27;
  wire in_26;
  wire in_25;
  wire in_24;
  wire in_23;
  wire in_22;
  wire in_21;
  wire in_20;
  wire in_19;
  wire in_18;
  wire in_17;
  wire in_16;
  wire in_15;
  wire in_14;
  wire in_13;
  wire in_12;
  wire in_11;
  wire in_10;
  wire in_9;
  wire in_8;
  wire in_7;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_3;
  wire in_2;
  wire in_1;
  wire in_0;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire in_81bar;
  wire in_80bar;
  wire in_79bar;
  wire in_78bar;
  wire in_77bar;
  wire in_76bar;
  wire in_75bar;
  wire in_74bar;
  wire in_73bar;
  wire in_72bar;
  wire in_71bar;
  wire in_70bar;
  wire in_69bar;
  wire in_68bar;
  wire in_67bar;
  wire in_66bar;
  wire in_65bar;
  wire in_64bar;
  wire in_63bar;
  wire in_62bar;
  wire in_61bar;
  wire in_60bar;
  wire in_59bar;
  wire in_58bar;
  wire in_57bar;
  wire in_56bar;
  wire in_55bar;
  wire in_54bar;
  wire in_53bar;
  wire in_52bar;
  wire in_51bar;
  wire in_50bar;
  wire in_49bar;
  wire in_48bar;
  wire in_47bar;
  wire in_46bar;
  wire in_45bar;
  wire in_44bar;
  wire in_43bar;
  wire in_42bar;
  wire in_41bar;
  wire in_40bar;
  wire in_39bar;
  wire in_38bar;
  wire in_37bar;
  wire in_36bar;
  wire in_35bar;
  wire in_34bar;
  wire in_33bar;
  wire in_32bar;
  wire in_31bar;
  wire in_30bar;
  wire in_29bar;
  wire in_28bar;
  wire in_27bar;
  wire in_26bar;
  wire in_25bar;
  wire in_24bar;
  wire in_23bar;
  wire in_22bar;
  wire in_21bar;
  wire in_20bar;
  wire in_19bar;
  wire in_18bar;
  wire in_17bar;
  wire in_16bar;
  wire in_15bar;
  wire in_14bar;
  wire in_13bar;
  wire in_12bar;
  wire in_11bar;
  wire in_10bar;
  wire in_9bar;
  wire in_8bar;
  wire in_7bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_3bar;
  wire in_2bar;
  wire in_1bar;
  wire in_0bar;
  wire n487bar;
  wire n488bar;
  wire n489bar;
  wire n490bar;
  wire n491bar;
  wire n492bar;
  wire n493bar;
  wire n494bar;
  wire n495bar;
  wire n496bar;
  wire n497bar;
  wire n498bar;
  wire n499bar;
  wire n500bar;
  wire n501bar;
  wire n502bar;
  wire n503bar;
  wire n504bar;
  wire n505bar;
  wire n506bar;
  wire n507bar;
  wire n508bar;
  wire n509bar;
  wire n510bar;
  wire n511bar;
  wire n512bar;
  wire n513bar;
  wire n514bar;
  wire n515bar;
  wire n516bar;
  wire n517bar;
  wire n518bar;
  wire n519bar;
  wire n520bar;
  wire n521bar;
  wire n522bar;
  wire n523bar;
  wire n524bar;
  wire n525bar;
  wire n526bar;
  wire n527bar;
  wire n528bar;
  wire n529bar;
  wire n530bar;
  wire n531bar;
  wire n532bar;
  wire n533bar;
  wire n534bar;
  wire n535bar;
  wire n536bar;
  wire n537bar;
  wire n538bar;
  wire n539bar;
  wire n540bar;
  wire n541bar;
  wire n542bar;
  wire n543bar;
  wire n544bar;
  wire n545bar;
  wire n546bar;
  wire n547bar;
  wire n548bar;
  wire n549bar;
  wire n550bar;
  wire n551bar;
  wire n552bar;
  wire n553bar;
  wire n554bar;
  wire n555bar;
  wire n556bar;
  wire n557bar;
  wire n558bar;
  wire n559bar;
  wire n560bar;
  wire n561bar;
  wire n562bar;
  wire n563bar;
  wire n564bar;
  wire n565bar;
  wire n566bar;
  wire n567bar;
  wire n568bar;
  wire n569bar;
  wire n570bar;
  wire n571bar;
  wire n572bar;
  wire n573bar;
  wire n574bar;
  wire n575bar;
  wire n576bar;
  wire n577bar;
  wire n578bar;
  wire n579bar;
  wire n580bar;
  wire n581bar;
  wire n582bar;
  wire n583bar;
  wire n584bar;
  wire n585bar;
  wire n586bar;
  wire n587bar;
  wire n588bar;
  wire n589bar;
  wire n590bar;
  wire n591bar;
  wire n592bar;
  wire n593bar;
  wire n594bar;
  wire n595bar;
  wire n596bar;
  wire n597bar;
  wire n598bar;
  wire n599bar;
  wire n600bar;
  wire n601bar;
  wire n602bar;
  wire n603bar;
  wire n604bar;
  wire n605bar;
  wire n606bar;
  wire n607bar;
  wire n608bar;
  wire n609bar;
  wire n610bar;
  wire n611bar;
  wire n612bar;
  wire n613bar;
  wire n614bar;
  wire n615bar;
  wire n616bar;
  wire n617bar;
  wire n618bar;
  wire n619bar;
  wire n620bar;
  wire n621bar;
  wire n622bar;
  wire n623bar;
  wire n624bar;
  wire n625bar;
  wire n626bar;
  wire n627bar;
  wire n628bar;
  wire n629bar;
  wire n630bar;
  wire n631bar;
  wire n632bar;
  wire n633bar;
  wire n634bar;
  wire n635bar;
  wire n636bar;
  wire n637bar;
  wire n638bar;
  wire n639bar;
  wire n640bar;
  wire n641bar;
  wire n642bar;
  wire n643bar;
  wire n644bar;
  wire n645bar;
  wire n646bar;
  wire n647bar;
  wire n648bar;
  wire n649bar;
  wire n650bar;
  wire n651bar;
  wire n652bar;
  wire n653bar;
  wire n654bar;
  wire n655bar;
  wire n656bar;
  wire n657bar;
  wire n658bar;
  wire n659bar;
  wire n660bar;
  wire n661bar;
  wire n662bar;
  wire n663bar;
  wire n664bar;
  wire n665bar;
  wire n666bar;
  wire n667bar;
  wire n668bar;
  wire n669bar;
  wire n670bar;
  wire n671bar;
  wire n672bar;
  wire n673bar;
  wire n674bar;
  wire n675bar;
  wire n676bar;
  wire n677bar;
  wire n678bar;
  wire n679bar;
  wire n680bar;
  wire n681bar;
  wire n682bar;
  wire n683bar;
  wire n684bar;
  wire n685bar;
  wire n686bar;
  wire n687bar;
  wire n688bar;
  wire n689bar;
  wire n690bar;
  wire n691bar;
  wire n692bar;
  wire n693bar;
  wire n694bar;
  wire n695bar;
  wire n696bar;
  wire n697bar;
  wire n698bar;
  wire n699bar;
  wire n700bar;
  wire n701bar;
  wire n702bar;
  wire n703bar;
  wire n704bar;
  wire n705bar;
  wire n706bar;
  wire n707bar;
  wire n708bar;
  wire n709bar;
  wire n710bar;
  wire n711bar;
  wire n712bar;
  wire n713bar;
  wire n714bar;
  wire n715bar;
  wire n716bar;
  wire n717bar;
  wire n718bar;
  wire n719bar;
  wire n720bar;
  wire n721bar;
  wire n722bar;
  wire n723bar;
  wire n724bar;
  wire n725bar;
  wire n726bar;
  wire n727bar;
  wire n728bar;
  wire n729bar;
  wire n730bar;
  wire n731bar;
  wire n732bar;
  wire n733bar;
  wire n734bar;
  wire n735bar;
  wire n736bar;
  wire n737bar;
  wire n738bar;
  wire n739bar;
  wire n740bar;
  wire n741bar;
  wire n742bar;
  wire n743bar;
  wire n744bar;
  wire n745bar;
  wire n746bar;
  wire n747bar;
  wire n748bar;
  wire n749bar;
  wire n750bar;
  wire n751bar;
  wire n752bar;
  wire n753bar;
  wire n754bar;
  wire n755bar;
  wire n756bar;
  wire n757bar;
  wire n758bar;
  wire n759bar;
  wire n760bar;
  wire n761bar;
  wire n762bar;
  wire n763bar;
  wire n764bar;
  wire n765bar;
  wire n766bar;
  wire n767bar;
  wire n768bar;
  wire n769bar;
  wire n770bar;
  wire n771bar;
  wire n772bar;
  wire n773bar;
  wire n774bar;
  wire n775bar;
  wire n776bar;
  wire n777bar;
  wire n778bar;
  wire n779bar;
  wire n780bar;
  wire n781bar;
  wire n782bar;
  wire n783bar;
  wire n784bar;
  wire n785bar;
  wire n786bar;
  wire n787bar;
  wire n788bar;
  wire n789bar;
  wire n790bar;
  wire n791bar;
  wire n792bar;
  wire n793bar;
  wire n794bar;
  wire n795bar;
  wire n796bar;
  wire n797bar;
  wire n798bar;
  wire n799bar;
  wire n800bar;
  wire n801bar;
  wire n802bar;
  wire n803bar;
  wire n804bar;
  wire n805bar;
  wire n806bar;
  wire n807bar;
  wire n808bar;
  wire n809bar;
  wire n810bar;
  wire n811bar;
  wire n812bar;
  wire n813bar;
  wire n814bar;
  wire n815bar;
  wire n816bar;
  wire n817bar;
  wire n818bar;
  wire n819bar;
  wire n820bar;
  wire n821bar;
  wire n822bar;
  wire n823bar;
  wire n824bar;
  wire n825bar;
  wire n826bar;
  wire n827bar;
  wire n828bar;
  wire n829bar;
  wire n830bar;
  wire n831bar;
  wire n832bar;
  wire n833bar;
  wire n834bar;
  wire n835bar;
  wire n836bar;
  wire n837bar;
  wire n838bar;
  wire n839bar;
  wire n840bar;
  wire n841bar;
  wire n842bar;
  wire n843bar;
  wire n844bar;
  wire n845bar;
  wire n846bar;
  wire n847bar;
  wire n848bar;
  wire n849bar;
  wire n850bar;
  wire n851bar;
  wire n852bar;
  wire n853bar;
  wire n854bar;
  wire n855bar;
  wire n856bar;
  wire n857bar;
  wire n858bar;
  wire n859bar;
  wire n860bar;
  wire n861bar;
  wire n862bar;
  wire n863bar;
  wire n864bar;
  wire n865bar;
  wire n866bar;
  wire n867bar;
  wire n868bar;
  wire n869bar;
  wire n870bar;
  wire n871bar;
  wire n872bar;
  wire n873bar;
  wire n874bar;
  wire n875bar;
  wire n876bar;
  wire n877bar;
  wire n878bar;
  wire n879bar;
  wire n880bar;
  wire n881bar;
  wire n882bar;
  wire n883bar;
  wire n884bar;
  wire n885bar;
  wire n886bar;
  wire n887bar;
  wire n888bar;
  wire n889bar;
  wire n890bar;
  wire n891bar;
  wire n892bar;
  wire n893bar;
  wire n894bar;
  wire n895bar;
  wire n896bar;
  wire n897bar;
  wire n898bar;
  wire n899bar;
  wire n900bar;
  wire n901bar;
  wire n902bar;
  wire n903bar;
  wire n904bar;
  wire n905bar;
  wire n906bar;
  wire n907bar;
  wire n908bar;
  wire n909bar;
  wire n910bar;
  wire n911bar;
  wire n912bar;
  wire n913bar;
  wire n914bar;
  wire n915bar;
  wire n916bar;
  wire n917bar;
  wire n918bar;
  wire n919bar;
  wire n920bar;
  wire n921bar;
  wire n922bar;
  wire n923bar;
  wire n924bar;
  wire n925bar;
  wire n926bar;
  wire n927bar;
  wire n928bar;
  wire n929bar;
  wire n930bar;
  wire n931bar;
  wire n932bar;
  wire n933bar;
  wire n934bar;
  wire n935bar;
  wire n936bar;
  wire n937bar;
  wire n938bar;
  wire n939bar;
  wire n940bar;
  wire n941bar;
  wire n942bar;
  wire n943bar;
  wire n944bar;
  wire n945bar;
  wire n946bar;
  wire n947bar;
  wire n948bar;
  wire n949bar;
  wire n950bar;
  wire n951bar;
  wire n952bar;
  wire n953bar;
  wire n954bar;
  wire n955bar;
  wire n956bar;
  wire n957bar;
  wire n958bar;
  wire n959bar;
  wire n960bar;
  wire n961bar;
  wire n962bar;
  wire n963bar;
  wire n964bar;
  wire n965bar;
  wire n966bar;
  wire n967bar;
  wire n968bar;
  wire n969bar;
  wire n970bar;
  wire n971bar;
  wire n972bar;
//wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];
  //OR U1
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U1 (
    .O(out[7]),
    .I0(n972),
    .I1(n971)
  );
  //AND U1bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U1bar (
    .O(outbar[7]),
    .I0(n972bar),
    .I1(n971bar)
  );
  //OR U2
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U2 (
    .O(n971),
    .I0(n970),
    .I1(n969)
  );
  //AND U2bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U2bar (
    .O(n971bar),
    .I0(n970bar),
    .I1(n969bar)
  );
  //OR U3
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U3 (
    .O(n969),
    .I0(n968),
    .I1(n967)
  );
  //AND U3bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U3bar (
    .O(n969bar),
    .I0(n968bar),
    .I1(n967bar)
  );
  //OR U4
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U4 (
    .O(n967),
    .I0(n966),
    .I1(n965)
  );
  //AND U4bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U4bar (
    .O(n967bar),
    .I0(n966bar),
    .I1(n965bar)
  );
  //OR U5
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U5 (
    .O(n968),
    .I0(n964),
    .I1(n963)
  );
  //AND U5bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U5bar (
    .O(n968bar),
    .I0(n964bar),
    .I1(n963bar)
  );
  //OR U6
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U6 (
    .O(n963),
    .I0(in[116]),
    .I1(n962)
  );
  //AND U6bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U6bar (
    .O(n963bar),
    .I0(inbar[116]),
    .I1(n962bar)
  );
  //OR U7
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U7 (
    .O(n970),
    .I0(n961),
    .I1(n960)
  );
  //AND U7bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U7bar (
    .O(n970bar),
    .I0(n961bar),
    .I1(n960bar)
  );
  //OR U8
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U8 (
    .O(n960),
    .I0(in[150]),
    .I1(in[127])
  );
  //AND U8bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U8bar (
    .O(n960bar),
    .I0(inbar[150]),
    .I1(inbar[127])
  );
  //OR U9
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U9 (
    .O(n961),
    .I0(in[160]),
    .I1(n959)
  );
  //AND U9bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U9bar (
    .O(n961bar),
    .I0(inbar[160]),
    .I1(n959bar)
  );
  //OR U10
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U10 (
    .O(n959),
    .I0(in[252]),
    .I1(in[168])
  );
  //AND U10bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U10bar (
    .O(n959bar),
    .I0(inbar[252]),
    .I1(inbar[168])
  );
  //OR U11
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U11 (
    .O(n972),
    .I0(n958),
    .I1(n957)
  );
  //AND U11bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U11bar (
    .O(n972bar),
    .I0(n958bar),
    .I1(n957bar)
  );
  //OR U12
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U12 (
    .O(n957),
    .I0(n956),
    .I1(n955)
  );
  //AND U12bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U12bar (
    .O(n957bar),
    .I0(n956bar),
    .I1(n955bar)
  );
  //OR U13
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U13 (
    .O(n955),
    .I0(in_17),
    .I1(in[96])
  );
  //AND U13bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U13bar (
    .O(n955bar),
    .I0(in_17bar),
    .I1(inbar[96])
  );
  //OR U14
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U14 (
    .O(n956),
    .I0(in_23),
    .I1(n954)
  );
  //AND U14bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U14bar (
    .O(n956bar),
    .I0(in_23bar),
    .I1(n954bar)
  );
  //OR U15
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U15 (
    .O(n954),
    .I0(in_31),
    .I1(in_26)
  );
  //AND U15bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U15bar (
    .O(n954bar),
    .I0(in_31bar),
    .I1(in_26bar)
  );
  //OR U16
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U16 (
    .O(n958),
    .I0(n953),
    .I1(n952)
  );
  //AND U16bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U16bar (
    .O(n958bar),
    .I0(n953bar),
    .I1(n952bar)
  );
  //OR U17
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U17 (
    .O(n952),
    .I0(in_58),
    .I1(in_4)
  );
  //AND U17bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U17bar (
    .O(n952bar),
    .I0(in_58bar),
    .I1(in_4bar)
  );
  //OR U18
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U18 (
    .O(n953),
    .I0(in_59),
    .I1(n951)
  );
  //AND U18bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U18bar (
    .O(n953bar),
    .I0(in_59bar),
    .I1(n951bar)
  );
  //OR U19
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U19 (
    .O(n951),
    .I0(in_71),
    .I1(in_62)
  );
  //AND U19bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U19bar (
    .O(n951bar),
    .I0(in_71bar),
    .I1(in_62bar)
  );
  //OR U20
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U20 (
    .O(out[6]),
    .I0(n950),
    .I1(n949)
  );
  //AND U20bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U20bar (
    .O(outbar[6]),
    .I0(n950bar),
    .I1(n949bar)
  );
  //OR U21
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U21 (
    .O(n949),
    .I0(n948),
    .I1(n947)
  );
  //AND U21bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U21bar (
    .O(n949bar),
    .I0(n948bar),
    .I1(n947bar)
  );
  //OR U22
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U22 (
    .O(n947),
    .I0(n946),
    .I1(n945)
  );
  //AND U22bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U22bar (
    .O(n947bar),
    .I0(n946bar),
    .I1(n945bar)
  );
  //OR U23
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U23 (
    .O(n945),
    .I0(n944),
    .I1(n943)
  );
  //AND U23bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U23bar (
    .O(n945bar),
    .I0(n944bar),
    .I1(n943bar)
  );
  //OR U24
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U24 (
    .O(n946),
    .I0(n942),
    .I1(n941)
  );
  //AND U24bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U24bar (
    .O(n946bar),
    .I0(n942bar),
    .I1(n941bar)
  );
  //OR U25
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U25 (
    .O(n941),
    .I0(in[101]),
    .I1(n940)
  );
  //AND U25bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U25bar (
    .O(n941bar),
    .I0(inbar[101]),
    .I1(n940bar)
  );
  //OR U26
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U26 (
    .O(n948),
    .I0(n939),
    .I1(n938)
  );
  //AND U26bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U26bar (
    .O(n948bar),
    .I0(n939bar),
    .I1(n938bar)
  );
  //OR U27
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U27 (
    .O(n938),
    .I0(in[114]),
    .I1(in[104])
  );
  //AND U27bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U27bar (
    .O(n938bar),
    .I0(inbar[114]),
    .I1(inbar[104])
  );
  //OR U28
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U28 (
    .O(n939),
    .I0(in[128]),
    .I1(n937)
  );
  //AND U28bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U28bar (
    .O(n939bar),
    .I0(inbar[128]),
    .I1(n937bar)
  );
  //OR U29
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U29 (
    .O(n937),
    .I0(in[136]),
    .I1(in[134])
  );
  //AND U29bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U29bar (
    .O(n937bar),
    .I0(inbar[136]),
    .I1(inbar[134])
  );
  //OR U30
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U30 (
    .O(n950),
    .I0(n936),
    .I1(n935)
  );
  //AND U30bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U30bar (
    .O(n950bar),
    .I0(n936bar),
    .I1(n935bar)
  );
  //OR U31
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U31 (
    .O(n935),
    .I0(n934),
    .I1(n933)
  );
  //AND U31bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U31bar (
    .O(n935bar),
    .I0(n934bar),
    .I1(n933bar)
  );
  //OR U32
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U32 (
    .O(n933),
    .I0(in[177]),
    .I1(in[164])
  );
  //AND U32bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U32bar (
    .O(n933bar),
    .I0(inbar[177]),
    .I1(inbar[164])
  );
  //OR U33
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U33 (
    .O(n934),
    .I0(in[212]),
    .I1(n932)
  );
  //AND U33bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U33bar (
    .O(n934bar),
    .I0(inbar[212]),
    .I1(n932bar)
  );
  //OR U34
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U34 (
    .O(n932),
    .I0(in[248]),
    .I1(in[221])
  );
  //AND U34bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U34bar (
    .O(n932bar),
    .I0(inbar[248]),
    .I1(inbar[221])
  );
  //OR U35
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U35 (
    .O(n936),
    .I0(n931),
    .I1(n930)
  );
  //AND U35bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U35bar (
    .O(n936bar),
    .I0(n931bar),
    .I1(n930bar)
  );
  //OR U36
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U36 (
    .O(n930),
    .I0(in_18),
    .I1(in[93])
  );
  //AND U36bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U36bar (
    .O(n930bar),
    .I0(in_18bar),
    .I1(inbar[93])
  );
  //OR U37
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U37 (
    .O(n931),
    .I0(in_31),
    .I1(n929)
  );
  //AND U37bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U37bar (
    .O(n931bar),
    .I0(in_31bar),
    .I1(n929bar)
  );
  //OR U38
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U38 (
    .O(n929),
    .I0(in_7),
    .I1(in_39)
  );
  //AND U38bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U38bar (
    .O(n929bar),
    .I0(in_7bar),
    .I1(in_39bar)
  );
  //OR U39
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U39 (
    .O(out[5]),
    .I0(n928),
    .I1(n927)
  );
  //AND U39bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U39bar (
    .O(outbar[5]),
    .I0(n928bar),
    .I1(n927bar)
  );
  //OR U40
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U40 (
    .O(n927),
    .I0(n926),
    .I1(n925)
  );
  //AND U40bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U40bar (
    .O(n927bar),
    .I0(n926bar),
    .I1(n925bar)
  );
  //OR U41
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U41 (
    .O(n925),
    .I0(n924),
    .I1(n923)
  );
  //AND U41bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U41bar (
    .O(n925bar),
    .I0(n924bar),
    .I1(n923bar)
  );
  //OR U42
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U42 (
    .O(n923),
    .I0(n922),
    .I1(n921)
  );
  //AND U42bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U42bar (
    .O(n923bar),
    .I0(n922bar),
    .I1(n921bar)
  );
  //OR U43
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U43 (
    .O(n924),
    .I0(n940),
    .I1(n920)
  );
  //AND U43bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U43bar (
    .O(n924bar),
    .I0(n940bar),
    .I1(n920bar)
  );
  //OR U44
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U44 (
    .O(n920),
    .I0(in[111]),
    .I1(n919)
  );
  //AND U44bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U44bar (
    .O(n920bar),
    .I0(inbar[111]),
    .I1(n919bar)
  );
  //OR U45
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U45 (
    .O(n940),
    .I0(n918),
    .I1(n917)
  );
  //AND U45bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U45bar (
    .O(n940bar),
    .I0(n918bar),
    .I1(n917bar)
  );
  //OR U46
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U46 (
    .O(n917),
    .I0(n916),
    .I1(n915)
  );
  //AND U46bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U46bar (
    .O(n917bar),
    .I0(n916bar),
    .I1(n915bar)
  );
  //OR U47
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U47 (
    .O(n915),
    .I0(n914),
    .I1(n913)
  );
  //AND U47bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U47bar (
    .O(n915bar),
    .I0(n914bar),
    .I1(n913bar)
  );
  //OR U48
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U48 (
    .O(n913),
    .I0(in[140]),
    .I1(in[131])
  );
  //AND U48bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U48bar (
    .O(n913bar),
    .I0(inbar[140]),
    .I1(inbar[131])
  );
  //OR U49
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U49 (
    .O(n914),
    .I0(in[160]),
    .I1(in[144])
  );
  //AND U49bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U49bar (
    .O(n914bar),
    .I0(inbar[160]),
    .I1(inbar[144])
  );
  //OR U50
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U50 (
    .O(n916),
    .I0(n912),
    .I1(n911)
  );
  //AND U50bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U50bar (
    .O(n916bar),
    .I0(n912bar),
    .I1(n911bar)
  );
  //OR U51
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U51 (
    .O(n911),
    .I0(in[179]),
    .I1(in[174])
  );
  //AND U51bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U51bar (
    .O(n911bar),
    .I0(inbar[179]),
    .I1(inbar[174])
  );
  //OR U52
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U52 (
    .O(n912),
    .I0(in[188]),
    .I1(in[184])
  );
  //AND U52bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U52bar (
    .O(n912bar),
    .I0(inbar[188]),
    .I1(inbar[184])
  );
  //OR U53
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U53 (
    .O(n918),
    .I0(n910),
    .I1(n909)
  );
  //AND U53bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U53bar (
    .O(n918bar),
    .I0(n910bar),
    .I1(n909bar)
  );
  //OR U54
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U54 (
    .O(n909),
    .I0(n908),
    .I1(n907)
  );
  //AND U54bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U54bar (
    .O(n909bar),
    .I0(n908bar),
    .I1(n907bar)
  );
  //OR U55
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U55 (
    .O(n907),
    .I0(in[216]),
    .I1(in[200])
  );
  //AND U55bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U55bar (
    .O(n907bar),
    .I0(inbar[216]),
    .I1(inbar[200])
  );
  //OR U56
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U56 (
    .O(n908),
    .I0(in[228]),
    .I1(in[224])
  );
  //AND U56bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U56bar (
    .O(n908bar),
    .I0(inbar[228]),
    .I1(inbar[224])
  );
  //OR U57
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U57 (
    .O(n910),
    .I0(n906),
    .I1(n905)
  );
  //AND U57bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U57bar (
    .O(n910bar),
    .I0(n906bar),
    .I1(n905bar)
  );
  //OR U58
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U58 (
    .O(n905),
    .I0(in[247]),
    .I1(in[235])
  );
  //AND U58bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U58bar (
    .O(n905bar),
    .I0(inbar[247]),
    .I1(inbar[235])
  );
  //OR U59
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U59 (
    .O(n906),
    .I0(in_42),
    .I1(in[83])
  );
  //AND U59bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U59bar (
    .O(n906bar),
    .I0(in_42bar),
    .I1(inbar[83])
  );
  //OR U60
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U60 (
    .O(n926),
    .I0(n904),
    .I1(n903)
  );
  //AND U60bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U60bar (
    .O(n926bar),
    .I0(n904bar),
    .I1(n903bar)
  );
  //OR U61
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U61 (
    .O(n903),
    .I0(in[166]),
    .I1(in[123])
  );
  //AND U61bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U61bar (
    .O(n903bar),
    .I0(inbar[166]),
    .I1(inbar[123])
  );
  //OR U62
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U62 (
    .O(n904),
    .I0(in[170]),
    .I1(n902)
  );
  //AND U62bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U62bar (
    .O(n904bar),
    .I0(inbar[170]),
    .I1(n902bar)
  );
  //OR U63
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U63 (
    .O(n902),
    .I0(in[194]),
    .I1(in[183])
  );
  //AND U63bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U63bar (
    .O(n902bar),
    .I0(inbar[194]),
    .I1(inbar[183])
  );
  //OR U64
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U64 (
    .O(n928),
    .I0(n901),
    .I1(n900)
  );
  //AND U64bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U64bar (
    .O(n928bar),
    .I0(n901bar),
    .I1(n900bar)
  );
  //OR U65
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U65 (
    .O(n900),
    .I0(n899),
    .I1(n898)
  );
  //AND U65bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U65bar (
    .O(n900bar),
    .I0(n899bar),
    .I1(n898bar)
  );
  //OR U66
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U66 (
    .O(n898),
    .I0(in[241]),
    .I1(in[238])
  );
  //AND U66bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U66bar (
    .O(n898bar),
    .I0(inbar[241]),
    .I1(inbar[238])
  );
  //OR U67
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U67 (
    .O(n899),
    .I0(in[250]),
    .I1(n897)
  );
  //AND U67bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U67bar (
    .O(n899bar),
    .I0(inbar[250]),
    .I1(n897bar)
  );
  //OR U68
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U68 (
    .O(n897),
    .I0(in_24),
    .I1(in[84])
  );
  //AND U68bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U68bar (
    .O(n897bar),
    .I0(in_24bar),
    .I1(inbar[84])
  );
  //OR U69
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U69 (
    .O(n901),
    .I0(n896),
    .I1(n895)
  );
  //AND U69bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U69bar (
    .O(n901bar),
    .I0(n896bar),
    .I1(n895bar)
  );
  //OR U70
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U70 (
    .O(n895),
    .I0(in_41),
    .I1(in_29)
  );
  //AND U70bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U70bar (
    .O(n895bar),
    .I0(in_41bar),
    .I1(in_29bar)
  );
  //OR U71
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U71 (
    .O(n896),
    .I0(in_66),
    .I1(n894)
  );
  //AND U71bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U71bar (
    .O(n896bar),
    .I0(in_66bar),
    .I1(n894bar)
  );
  //OR U72
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U72 (
    .O(n894),
    .I0(in_76),
    .I1(in_71)
  );
  //AND U72bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U72bar (
    .O(n894bar),
    .I0(in_76bar),
    .I1(in_71bar)
  );
  //OR U73
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U73 (
    .O(out[4]),
    .I0(n893),
    .I1(n892)
  );
  //AND U73bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U73bar (
    .O(outbar[4]),
    .I0(n893bar),
    .I1(n892bar)
  );
  //OR U74
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U74 (
    .O(n892),
    .I0(n891),
    .I1(n890)
  );
  //AND U74bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U74bar (
    .O(n892bar),
    .I0(n891bar),
    .I1(n890bar)
  );
  //OR U75
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U75 (
    .O(n890),
    .I0(n889),
    .I1(n888)
  );
  //AND U75bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U75bar (
    .O(n890bar),
    .I0(n889bar),
    .I1(n888bar)
  );
  //OR U76
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U76 (
    .O(n888),
    .I0(n922),
    .I1(n887)
  );
  //AND U76bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U76bar (
    .O(n888bar),
    .I0(n922bar),
    .I1(n887bar)
  );
  //OR U77
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U77 (
    .O(n922),
    .I0(n886),
    .I1(n885)
  );
  //AND U77bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U77bar (
    .O(n922bar),
    .I0(n886bar),
    .I1(n885bar)
  );
  //OR U78
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U78 (
    .O(n885),
    .I0(n884),
    .I1(n883)
  );
  //AND U78bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U78bar (
    .O(n885bar),
    .I0(n884bar),
    .I1(n883bar)
  );
  //OR U79
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U79 (
    .O(n883),
    .I0(n882),
    .I1(n881)
  );
  //AND U79bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U79bar (
    .O(n883bar),
    .I0(n882bar),
    .I1(n881bar)
  );
  //OR U80
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U80 (
    .O(n881),
    .I0(in[118]),
    .I1(in[109])
  );
  //AND U80bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U80bar (
    .O(n881bar),
    .I0(inbar[118]),
    .I1(inbar[109])
  );
  //OR U81
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U81 (
    .O(n882),
    .I0(in[139]),
    .I1(in[120])
  );
  //AND U81bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U81bar (
    .O(n882bar),
    .I0(inbar[139]),
    .I1(inbar[120])
  );
  //OR U82
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U82 (
    .O(n884),
    .I0(n880),
    .I1(n879)
  );
  //AND U82bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U82bar (
    .O(n884bar),
    .I0(n880bar),
    .I1(n879bar)
  );
  //OR U83
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U83 (
    .O(n879),
    .I0(in[198]),
    .I1(in[154])
  );
  //AND U83bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U83bar (
    .O(n879bar),
    .I0(inbar[198]),
    .I1(inbar[154])
  );
  //OR U84
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U84 (
    .O(n880),
    .I0(in[210]),
    .I1(in[205])
  );
  //AND U84bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U84bar (
    .O(n880bar),
    .I0(inbar[210]),
    .I1(inbar[205])
  );
  //OR U85
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U85 (
    .O(n886),
    .I0(n878),
    .I1(n877)
  );
  //AND U85bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U85bar (
    .O(n886bar),
    .I0(n878bar),
    .I1(n877bar)
  );
  //OR U86
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U86 (
    .O(n877),
    .I0(n876),
    .I1(n875)
  );
  //AND U86bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U86bar (
    .O(n877bar),
    .I0(n876bar),
    .I1(n875bar)
  );
  //OR U87
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U87 (
    .O(n875),
    .I0(in[219]),
    .I1(in[217])
  );
  //AND U87bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U87bar (
    .O(n875bar),
    .I0(inbar[219]),
    .I1(inbar[217])
  );
  //OR U88
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U88 (
    .O(n876),
    .I0(in[86]),
    .I1(in[252])
  );
  //AND U88bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U88bar (
    .O(n876bar),
    .I0(inbar[86]),
    .I1(inbar[252])
  );
  //OR U89
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U89 (
    .O(n878),
    .I0(n874),
    .I1(n873)
  );
  //AND U89bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U89bar (
    .O(n878bar),
    .I0(n874bar),
    .I1(n873bar)
  );
  //OR U90
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U90 (
    .O(n873),
    .I0(in_40),
    .I1(in[91])
  );
  //AND U90bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U90bar (
    .O(n873bar),
    .I0(in_40bar),
    .I1(inbar[91])
  );
  //OR U91
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U91 (
    .O(n874),
    .I0(in_8),
    .I1(in_46)
  );
  //AND U91bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U91bar (
    .O(n874bar),
    .I0(in_8bar),
    .I1(in_46bar)
  );
  //OR U92
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U92 (
    .O(n889),
    .I0(n872),
    .I1(n871)
  );
  //AND U92bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U92bar (
    .O(n889bar),
    .I0(n872bar),
    .I1(n871bar)
  );
  //OR U93
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U93 (
    .O(n871),
    .I0(in[117]),
    .I1(n943)
  );
  //AND U93bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U93bar (
    .O(n871bar),
    .I0(inbar[117]),
    .I1(n943bar)
  );
  //OR U94
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U94 (
    .O(n943),
    .I0(n870),
    .I1(n869)
  );
  //AND U94bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U94bar (
    .O(n943bar),
    .I0(n870bar),
    .I1(n869bar)
  );
  //OR U95
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U95 (
    .O(n869),
    .I0(n868),
    .I1(n867)
  );
  //AND U95bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U95bar (
    .O(n869bar),
    .I0(n868bar),
    .I1(n867bar)
  );
  //OR U96
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U96 (
    .O(n867),
    .I0(n866),
    .I1(n865)
  );
  //AND U96bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U96bar (
    .O(n867bar),
    .I0(n866bar),
    .I1(n865bar)
  );
  //OR U97
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U97 (
    .O(n865),
    .I0(n864),
    .I1(n863)
  );
  //AND U97bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U97bar (
    .O(n865bar),
    .I0(n864bar),
    .I1(n863bar)
  );
  //OR U98
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U98 (
    .O(n866),
    .I0(in[108]),
    .I1(n919)
  );
  //AND U98bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U98bar (
    .O(n866bar),
    .I0(inbar[108]),
    .I1(n919bar)
  );
  //OR U99
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U99 (
    .O(n919),
    .I0(n862),
    .I1(n861)
  );
  //AND U99bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U99bar (
    .O(n919bar),
    .I0(n862bar),
    .I1(n861bar)
  );
  //OR U100
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U100 (
    .O(n861),
    .I0(n860),
    .I1(n859)
  );
  //AND U100bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U100bar (
    .O(n861bar),
    .I0(n860bar),
    .I1(n859bar)
  );
  //OR U101
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U101 (
    .O(n859),
    .I0(n858),
    .I1(n857)
  );
  //AND U101bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U101bar (
    .O(n859bar),
    .I0(n858bar),
    .I1(n857bar)
  );
  //OR U102
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U102 (
    .O(n857),
    .I0(in[119]),
    .I1(in[105])
  );
  //AND U102bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U102bar (
    .O(n857bar),
    .I0(inbar[119]),
    .I1(inbar[105])
  );
  //OR U103
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U103 (
    .O(n858),
    .I0(in[186]),
    .I1(in[175])
  );
  //AND U103bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U103bar (
    .O(n858bar),
    .I0(inbar[186]),
    .I1(inbar[175])
  );
  //OR U104
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U104 (
    .O(n860),
    .I0(n856),
    .I1(n855)
  );
  //AND U104bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U104bar (
    .O(n860bar),
    .I0(n856bar),
    .I1(n855bar)
  );
  //OR U105
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U105 (
    .O(n855),
    .I0(in[202]),
    .I1(in[193])
  );
  //AND U105bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U105bar (
    .O(n855bar),
    .I0(inbar[202]),
    .I1(inbar[193])
  );
  //OR U106
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U106 (
    .O(n856),
    .I0(in[225]),
    .I1(in[208])
  );
  //AND U106bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U106bar (
    .O(n856bar),
    .I0(inbar[225]),
    .I1(inbar[208])
  );
  //OR U107
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U107 (
    .O(n862),
    .I0(n854),
    .I1(n853)
  );
  //AND U107bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U107bar (
    .O(n862bar),
    .I0(n854bar),
    .I1(n853bar)
  );
  //OR U108
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U108 (
    .O(n853),
    .I0(n852),
    .I1(n851)
  );
  //AND U108bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U108bar (
    .O(n853bar),
    .I0(n852bar),
    .I1(n851bar)
  );
  //OR U109
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U109 (
    .O(n851),
    .I0(in_1),
    .I1(in[85])
  );
  //AND U109bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U109bar (
    .O(n851bar),
    .I0(in_1bar),
    .I1(inbar[85])
  );
  //OR U110
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U110 (
    .O(n852),
    .I0(in_23),
    .I1(in_19)
  );
  //AND U110bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U110bar (
    .O(n852bar),
    .I0(in_23bar),
    .I1(in_19bar)
  );
  //OR U111
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U111 (
    .O(n854),
    .I0(n850),
    .I1(n849)
  );
  //AND U111bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U111bar (
    .O(n854bar),
    .I0(n850bar),
    .I1(n849bar)
  );
  //OR U112
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U112 (
    .O(n849),
    .I0(in_43),
    .I1(in_33)
  );
  //AND U112bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U112bar (
    .O(n849bar),
    .I0(in_43bar),
    .I1(in_33bar)
  );
  //OR U113
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U113 (
    .O(n850),
    .I0(in_63),
    .I1(in_44)
  );
  //AND U113bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U113bar (
    .O(n850bar),
    .I0(in_63bar),
    .I1(in_44bar)
  );
  //OR U114
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U114 (
    .O(n868),
    .I0(n848),
    .I1(n847)
  );
  //AND U114bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U114bar (
    .O(n868bar),
    .I0(n848bar),
    .I1(n847bar)
  );
  //OR U115
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U115 (
    .O(n847),
    .I0(in[141]),
    .I1(in[112])
  );
  //AND U115bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U115bar (
    .O(n847bar),
    .I0(inbar[141]),
    .I1(inbar[112])
  );
  //OR U116
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U116 (
    .O(n848),
    .I0(in[147]),
    .I1(n846)
  );
  //AND U116bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U116bar (
    .O(n848bar),
    .I0(inbar[147]),
    .I1(n846bar)
  );
  //OR U117
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U117 (
    .O(n846),
    .I0(in[181]),
    .I1(in[167])
  );
  //AND U117bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U117bar (
    .O(n846bar),
    .I0(inbar[181]),
    .I1(inbar[167])
  );
  //OR U118
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U118 (
    .O(n870),
    .I0(n845),
    .I1(n844)
  );
  //AND U118bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U118bar (
    .O(n870bar),
    .I0(n845bar),
    .I1(n844bar)
  );
  //OR U119
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U119 (
    .O(n844),
    .I0(n843),
    .I1(n842)
  );
  //AND U119bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U119bar (
    .O(n844bar),
    .I0(n843bar),
    .I1(n842bar)
  );
  //OR U120
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U120 (
    .O(n842),
    .I0(in[229]),
    .I1(in[201])
  );
  //AND U120bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U120bar (
    .O(n842bar),
    .I0(inbar[229]),
    .I1(inbar[201])
  );
  //OR U121
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U121 (
    .O(n843),
    .I0(in[237]),
    .I1(n841)
  );
  //AND U121bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U121bar (
    .O(n843bar),
    .I0(inbar[237]),
    .I1(n841bar)
  );
  //OR U122
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U122 (
    .O(n841),
    .I0(in[94]),
    .I1(in[253])
  );
  //AND U122bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U122bar (
    .O(n841bar),
    .I0(inbar[94]),
    .I1(inbar[253])
  );
  //OR U123
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U123 (
    .O(n845),
    .I0(n840),
    .I1(n839)
  );
  //AND U123bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U123bar (
    .O(n845bar),
    .I0(n840bar),
    .I1(n839bar)
  );
  //OR U124
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U124 (
    .O(n839),
    .I0(in_21),
    .I1(in[96])
  );
  //AND U124bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U124bar (
    .O(n839bar),
    .I0(in_21bar),
    .I1(inbar[96])
  );
  //OR U125
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U125 (
    .O(n840),
    .I0(in_25),
    .I1(n838)
  );
  //AND U125bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U125bar (
    .O(n840bar),
    .I0(in_25bar),
    .I1(n838bar)
  );
  //OR U126
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U126 (
    .O(n838),
    .I0(in_81),
    .I1(in_45)
  );
  //AND U126bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U126bar (
    .O(n838bar),
    .I0(in_81bar),
    .I1(in_45bar)
  );
  //OR U127
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U127 (
    .O(n891),
    .I0(n837),
    .I1(n836)
  );
  //AND U127bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U127bar (
    .O(n891bar),
    .I0(n837bar),
    .I1(n836bar)
  );
  //OR U128
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U128 (
    .O(n836),
    .I0(in[142]),
    .I1(in[124])
  );
  //AND U128bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U128bar (
    .O(n836bar),
    .I0(inbar[142]),
    .I1(inbar[124])
  );
  //OR U129
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U129 (
    .O(n837),
    .I0(in[150]),
    .I1(n835)
  );
  //AND U129bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U129bar (
    .O(n837bar),
    .I0(inbar[150]),
    .I1(n835bar)
  );
  //OR U130
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U130 (
    .O(n835),
    .I0(in[172]),
    .I1(in[155])
  );
  //AND U130bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U130bar (
    .O(n835bar),
    .I0(inbar[172]),
    .I1(inbar[155])
  );
  //OR U131
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U131 (
    .O(n893),
    .I0(n834),
    .I1(n833)
  );
  //AND U131bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U131bar (
    .O(n893bar),
    .I0(n834bar),
    .I1(n833bar)
  );
  //OR U132
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U132 (
    .O(n833),
    .I0(n832),
    .I1(n831)
  );
  //AND U132bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U132bar (
    .O(n833bar),
    .I0(n832bar),
    .I1(n831bar)
  );
  //OR U133
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U133 (
    .O(n831),
    .I0(in[196]),
    .I1(in[173])
  );
  //AND U133bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U133bar (
    .O(n831bar),
    .I0(inbar[196]),
    .I1(inbar[173])
  );
  //OR U134
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U134 (
    .O(n832),
    .I0(in[222]),
    .I1(n830)
  );
  //AND U134bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U134bar (
    .O(n832bar),
    .I0(inbar[222]),
    .I1(n830bar)
  );
  //OR U135
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U135 (
    .O(n830),
    .I0(in[227]),
    .I1(in[226])
  );
  //AND U135bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U135bar (
    .O(n830bar),
    .I0(inbar[227]),
    .I1(inbar[226])
  );
  //OR U136
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U136 (
    .O(n834),
    .I0(n829),
    .I1(n828)
  );
  //AND U136bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U136bar (
    .O(n834bar),
    .I0(n829bar),
    .I1(n828bar)
  );
  //OR U137
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U137 (
    .O(n828),
    .I0(in[249]),
    .I1(in[231])
  );
  //AND U137bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U137bar (
    .O(n828bar),
    .I0(inbar[249]),
    .I1(inbar[231])
  );
  //OR U138
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U138 (
    .O(n829),
    .I0(in_28),
    .I1(n827)
  );
  //AND U138bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U138bar (
    .O(n829bar),
    .I0(in_28bar),
    .I1(n827bar)
  );
  //OR U139
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U139 (
    .O(n827),
    .I0(in_52),
    .I1(in_47)
  );
  //AND U139bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U139bar (
    .O(n827bar),
    .I0(in_52bar),
    .I1(in_47bar)
  );
  //OR U140
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U140 (
    .O(out[3]),
    .I0(n826),
    .I1(n825)
  );
  //AND U140bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U140bar (
    .O(outbar[3]),
    .I0(n826bar),
    .I1(n825bar)
  );
  //OR U141
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U141 (
    .O(n825),
    .I0(n824),
    .I1(n823)
  );
  //AND U141bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U141bar (
    .O(n825bar),
    .I0(n824bar),
    .I1(n823bar)
  );
  //OR U142
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U142 (
    .O(n823),
    .I0(n822),
    .I1(n821)
  );
  //AND U142bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U142bar (
    .O(n823bar),
    .I0(n822bar),
    .I1(n821bar)
  );
  //OR U143
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U143 (
    .O(n821),
    .I0(n820),
    .I1(n819)
  );
  //AND U143bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U143bar (
    .O(n821bar),
    .I0(n820bar),
    .I1(n819bar)
  );
  //OR U144
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U144 (
    .O(n822),
    .I0(n964),
    .I1(n818)
  );
  //AND U144bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U144bar (
    .O(n822bar),
    .I0(n964bar),
    .I1(n818bar)
  );
  //OR U145
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U145 (
    .O(n818),
    .I0(in[118]),
    .I1(n817)
  );
  //AND U145bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U145bar (
    .O(n818bar),
    .I0(inbar[118]),
    .I1(n817bar)
  );
  //OR U146
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U146 (
    .O(n964),
    .I0(n816),
    .I1(n815)
  );
  //AND U146bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U146bar (
    .O(n964bar),
    .I0(n816bar),
    .I1(n815bar)
  );
  //OR U147
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U147 (
    .O(n815),
    .I0(n814),
    .I1(n813)
  );
  //AND U147bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U147bar (
    .O(n815bar),
    .I0(n814bar),
    .I1(n813bar)
  );
  //OR U148
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U148 (
    .O(n813),
    .I0(n812),
    .I1(n811)
  );
  //AND U148bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U148bar (
    .O(n813bar),
    .I0(n812bar),
    .I1(n811bar)
  );
  //OR U149
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U149 (
    .O(n811),
    .I0(in[122]),
    .I1(in[111])
  );
  //AND U149bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U149bar (
    .O(n811bar),
    .I0(inbar[122]),
    .I1(inbar[111])
  );
  //OR U150
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U150 (
    .O(n812),
    .I0(in[154]),
    .I1(in[151])
  );
  //AND U150bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U150bar (
    .O(n812bar),
    .I0(inbar[154]),
    .I1(inbar[151])
  );
  //OR U151
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U151 (
    .O(n814),
    .I0(n810),
    .I1(n809)
  );
  //AND U151bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U151bar (
    .O(n814bar),
    .I0(n810bar),
    .I1(n809bar)
  );
  //OR U152
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U152 (
    .O(n809),
    .I0(in[187]),
    .I1(in[177])
  );
  //AND U152bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U152bar (
    .O(n809bar),
    .I0(inbar[187]),
    .I1(inbar[177])
  );
  //OR U153
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U153 (
    .O(n810),
    .I0(in[200]),
    .I1(in[192])
  );
  //AND U153bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U153bar (
    .O(n810bar),
    .I0(inbar[200]),
    .I1(inbar[192])
  );
  //OR U154
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U154 (
    .O(n816),
    .I0(n808),
    .I1(n807)
  );
  //AND U154bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U154bar (
    .O(n816bar),
    .I0(n808bar),
    .I1(n807bar)
  );
  //OR U155
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U155 (
    .O(n807),
    .I0(n806),
    .I1(n805)
  );
  //AND U155bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U155bar (
    .O(n807bar),
    .I0(n806bar),
    .I1(n805bar)
  );
  //OR U156
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U156 (
    .O(n805),
    .I0(in[225]),
    .I1(in[207])
  );
  //AND U156bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U156bar (
    .O(n805bar),
    .I0(inbar[225]),
    .I1(inbar[207])
  );
  //OR U157
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U157 (
    .O(n806),
    .I0(in[98]),
    .I1(in[226])
  );
  //AND U157bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U157bar (
    .O(n806bar),
    .I0(inbar[98]),
    .I1(inbar[226])
  );
  //OR U158
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U158 (
    .O(n808),
    .I0(n804),
    .I1(n803)
  );
  //AND U158bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U158bar (
    .O(n808bar),
    .I0(n804bar),
    .I1(n803bar)
  );
  //OR U159
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U159 (
    .O(n803),
    .I0(in_20),
    .I1(in_16)
  );
  //AND U159bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U159bar (
    .O(n803bar),
    .I0(in_20bar),
    .I1(in_16bar)
  );
  //OR U160
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U160 (
    .O(n804),
    .I0(in_55),
    .I1(in_45)
  );
  //AND U160bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U160bar (
    .O(n804bar),
    .I0(in_55bar),
    .I1(in_45bar)
  );
  //OR U161
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U161 (
    .O(n824),
    .I0(n802),
    .I1(n801)
  );
  //AND U161bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U161bar (
    .O(n824bar),
    .I0(n802bar),
    .I1(n801bar)
  );
  //OR U162
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U162 (
    .O(n801),
    .I0(in[162]),
    .I1(in[149])
  );
  //AND U162bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U162bar (
    .O(n801bar),
    .I0(inbar[162]),
    .I1(inbar[149])
  );
  //OR U163
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U163 (
    .O(n802),
    .I0(in[163]),
    .I1(n800)
  );
  //AND U163bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U163bar (
    .O(n802bar),
    .I0(inbar[163]),
    .I1(n800bar)
  );
  //OR U164
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U164 (
    .O(n800),
    .I0(in[191]),
    .I1(in[189])
  );
  //AND U164bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U164bar (
    .O(n800bar),
    .I0(inbar[191]),
    .I1(inbar[189])
  );
  //OR U165
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U165 (
    .O(n826),
    .I0(n799),
    .I1(n798)
  );
  //AND U165bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U165bar (
    .O(n826bar),
    .I0(n799bar),
    .I1(n798bar)
  );
  //OR U166
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U166 (
    .O(n798),
    .I0(n797),
    .I1(n796)
  );
  //AND U166bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U166bar (
    .O(n798bar),
    .I0(n797bar),
    .I1(n796bar)
  );
  //OR U167
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U167 (
    .O(n796),
    .I0(in[212]),
    .I1(in[193])
  );
  //AND U167bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U167bar (
    .O(n796bar),
    .I0(inbar[212]),
    .I1(inbar[193])
  );
  //OR U168
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U168 (
    .O(n797),
    .I0(in[238]),
    .I1(n795)
  );
  //AND U168bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U168bar (
    .O(n797bar),
    .I0(inbar[238]),
    .I1(n795bar)
  );
  //OR U169
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U169 (
    .O(n795),
    .I0(in[88]),
    .I1(in[247])
  );
  //AND U169bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U169bar (
    .O(n795bar),
    .I0(inbar[88]),
    .I1(inbar[247])
  );
  //OR U170
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U170 (
    .O(n799),
    .I0(n794),
    .I1(n793)
  );
  //AND U170bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U170bar (
    .O(n799bar),
    .I0(n794bar),
    .I1(n793bar)
  );
  //OR U171
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U171 (
    .O(n793),
    .I0(in[94]),
    .I1(in[92])
  );
  //AND U171bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U171bar (
    .O(n793bar),
    .I0(inbar[94]),
    .I1(inbar[92])
  );
  //OR U172
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U172 (
    .O(n794),
    .I0(in_52),
    .I1(n792)
  );
  //AND U172bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U172bar (
    .O(n794bar),
    .I0(in_52bar),
    .I1(n792bar)
  );
  //OR U173
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U173 (
    .O(n792),
    .I0(in_70),
    .I1(in_67)
  );
  //AND U173bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U173bar (
    .O(n792bar),
    .I0(in_70bar),
    .I1(in_67bar)
  );
  //OR U174
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U174 (
    .O(out[2]),
    .I0(n791),
    .I1(n790)
  );
  //AND U174bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U174bar (
    .O(outbar[2]),
    .I0(n791bar),
    .I1(n790bar)
  );
  //OR U175
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U175 (
    .O(n790),
    .I0(n789),
    .I1(n788)
  );
  //AND U175bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U175bar (
    .O(n790bar),
    .I0(n789bar),
    .I1(n788bar)
  );
  //OR U176
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U176 (
    .O(n788),
    .I0(n787),
    .I1(n786)
  );
  //AND U176bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U176bar (
    .O(n788bar),
    .I0(n787bar),
    .I1(n786bar)
  );
  //OR U177
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U177 (
    .O(n786),
    .I0(n819),
    .I1(n785)
  );
  //AND U177bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U177bar (
    .O(n786bar),
    .I0(n819bar),
    .I1(n785bar)
  );
  //OR U178
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U178 (
    .O(n819),
    .I0(n784),
    .I1(n783)
  );
  //AND U178bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U178bar (
    .O(n819bar),
    .I0(n784bar),
    .I1(n783bar)
  );
  //OR U179
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U179 (
    .O(n783),
    .I0(n782),
    .I1(n781)
  );
  //AND U179bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U179bar (
    .O(n783bar),
    .I0(n782bar),
    .I1(n781bar)
  );
  //OR U180
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U180 (
    .O(n781),
    .I0(n780),
    .I1(n779)
  );
  //AND U180bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U180bar (
    .O(n781bar),
    .I0(n780bar),
    .I1(n779bar)
  );
  //OR U181
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U181 (
    .O(n779),
    .I0(n962),
    .I1(n778)
  );
  //AND U181bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U181bar (
    .O(n779bar),
    .I0(n962bar),
    .I1(n778bar)
  );
  //OR U182
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U182 (
    .O(n962),
    .I0(n777),
    .I1(n776)
  );
  //AND U182bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U182bar (
    .O(n962bar),
    .I0(n777bar),
    .I1(n776bar)
  );
  //OR U183
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U183 (
    .O(n776),
    .I0(n775),
    .I1(n774)
  );
  //AND U183bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U183bar (
    .O(n776bar),
    .I0(n775bar),
    .I1(n774bar)
  );
  //OR U184
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U184 (
    .O(n774),
    .I0(n773),
    .I1(n772)
  );
  //AND U184bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U184bar (
    .O(n774bar),
    .I0(n773bar),
    .I1(n772bar)
  );
  //OR U185
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U185 (
    .O(n772),
    .I0(in[131]),
    .I1(in[120])
  );
  //AND U185bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U185bar (
    .O(n772bar),
    .I0(inbar[131]),
    .I1(inbar[120])
  );
  //OR U186
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U186 (
    .O(n773),
    .I0(in[153]),
    .I1(in[147])
  );
  //AND U186bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U186bar (
    .O(n773bar),
    .I0(inbar[153]),
    .I1(inbar[147])
  );
  //OR U187
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U187 (
    .O(n775),
    .I0(n771),
    .I1(n770)
  );
  //AND U187bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U187bar (
    .O(n775bar),
    .I0(n771bar),
    .I1(n770bar)
  );
  //OR U188
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U188 (
    .O(n770),
    .I0(in[170]),
    .I1(in[156])
  );
  //AND U188bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U188bar (
    .O(n770bar),
    .I0(inbar[170]),
    .I1(inbar[156])
  );
  //OR U189
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U189 (
    .O(n771),
    .I0(in[223]),
    .I1(in[190])
  );
  //AND U189bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U189bar (
    .O(n771bar),
    .I0(inbar[223]),
    .I1(inbar[190])
  );
  //OR U190
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U190 (
    .O(n777),
    .I0(n769),
    .I1(n768)
  );
  //AND U190bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U190bar (
    .O(n777bar),
    .I0(n769bar),
    .I1(n768bar)
  );
  //OR U191
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U191 (
    .O(n768),
    .I0(n767),
    .I1(n766)
  );
  //AND U191bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U191bar (
    .O(n768bar),
    .I0(n767bar),
    .I1(n766bar)
  );
  //OR U192
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U192 (
    .O(n766),
    .I0(in[236]),
    .I1(in[230])
  );
  //AND U192bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U192bar (
    .O(n766bar),
    .I0(inbar[236]),
    .I1(inbar[230])
  );
  //OR U193
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U193 (
    .O(n767),
    .I0(in[85]),
    .I1(in[240])
  );
  //AND U193bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U193bar (
    .O(n767bar),
    .I0(inbar[85]),
    .I1(inbar[240])
  );
  //OR U194
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U194 (
    .O(n769),
    .I0(n765),
    .I1(n764)
  );
  //AND U194bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U194bar (
    .O(n769bar),
    .I0(n765bar),
    .I1(n764bar)
  );
  //OR U195
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U195 (
    .O(n764),
    .I0(in_12),
    .I1(in[90])
  );
  //AND U195bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U195bar (
    .O(n764bar),
    .I0(in_12bar),
    .I1(inbar[90])
  );
  //OR U196
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U196 (
    .O(n765),
    .I0(in_39),
    .I1(in_28)
  );
  //AND U196bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U196bar (
    .O(n765bar),
    .I0(in_39bar),
    .I1(in_28bar)
  );
  //OR U197
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U197 (
    .O(n780),
    .I0(in[109]),
    .I1(n763)
  );
  //AND U197bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U197bar (
    .O(n780bar),
    .I0(inbar[109]),
    .I1(n763bar)
  );
  //OR U198
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U198 (
    .O(n782),
    .I0(n762),
    .I1(n761)
  );
  //AND U198bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U198bar (
    .O(n782bar),
    .I0(n762bar),
    .I1(n761bar)
  );
  //OR U199
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U199 (
    .O(n761),
    .I0(in[138]),
    .I1(in[129])
  );
  //AND U199bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U199bar (
    .O(n761bar),
    .I0(inbar[138]),
    .I1(inbar[129])
  );
  //OR U200
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U200 (
    .O(n762),
    .I0(in[157]),
    .I1(n760)
  );
  //AND U200bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U200bar (
    .O(n762bar),
    .I0(inbar[157]),
    .I1(n760bar)
  );
  //OR U201
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U201 (
    .O(n760),
    .I0(in[182]),
    .I1(in[167])
  );
  //AND U201bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U201bar (
    .O(n760bar),
    .I0(inbar[182]),
    .I1(inbar[167])
  );
  //OR U202
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U202 (
    .O(n784),
    .I0(n759),
    .I1(n758)
  );
  //AND U202bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U202bar (
    .O(n784bar),
    .I0(n759bar),
    .I1(n758bar)
  );
  //OR U203
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U203 (
    .O(n758),
    .I0(n757),
    .I1(n756)
  );
  //AND U203bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U203bar (
    .O(n758bar),
    .I0(n757bar),
    .I1(n756bar)
  );
  //OR U204
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U204 (
    .O(n756),
    .I0(in[195]),
    .I1(in[184])
  );
  //AND U204bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U204bar (
    .O(n756bar),
    .I0(inbar[195]),
    .I1(inbar[184])
  );
  //OR U205
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U205 (
    .O(n757),
    .I0(in[196]),
    .I1(n755)
  );
  //AND U205bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U205bar (
    .O(n757bar),
    .I0(inbar[196]),
    .I1(n755bar)
  );
  //OR U206
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U206 (
    .O(n755),
    .I0(in[215]),
    .I1(in[209])
  );
  //AND U206bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U206bar (
    .O(n755bar),
    .I0(inbar[215]),
    .I1(inbar[209])
  );
  //OR U207
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U207 (
    .O(n759),
    .I0(n754),
    .I1(n753)
  );
  //AND U207bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U207bar (
    .O(n759bar),
    .I0(n754bar),
    .I1(n753bar)
  );
  //OR U208
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U208 (
    .O(n753),
    .I0(in[93]),
    .I1(in[233])
  );
  //AND U208bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U208bar (
    .O(n753bar),
    .I0(inbar[93]),
    .I1(inbar[233])
  );
  //OR U209
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U209 (
    .O(n754),
    .I0(in_1),
    .I1(n752)
  );
  //AND U209bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U209bar (
    .O(n754bar),
    .I0(in_1bar),
    .I1(n752bar)
  );
  //OR U210
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U210 (
    .O(n752),
    .I0(in_69),
    .I1(in_66)
  );
  //AND U210bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U210bar (
    .O(n752bar),
    .I0(in_69bar),
    .I1(in_66bar)
  );
  //OR U211
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U211 (
    .O(n787),
    .I0(n966),
    .I1(n751)
  );
  //AND U211bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U211bar (
    .O(n787bar),
    .I0(n966bar),
    .I1(n751bar)
  );
  //OR U212
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U212 (
    .O(n751),
    .I0(in[134]),
    .I1(n750)
  );
  //AND U212bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U212bar (
    .O(n751bar),
    .I0(inbar[134]),
    .I1(n750bar)
  );
  //OR U213
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U213 (
    .O(n966),
    .I0(n749),
    .I1(n748)
  );
  //AND U213bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U213bar (
    .O(n966bar),
    .I0(n749bar),
    .I1(n748bar)
  );
  //OR U214
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U214 (
    .O(n748),
    .I0(n747),
    .I1(n746)
  );
  //AND U214bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U214bar (
    .O(n748bar),
    .I0(n747bar),
    .I1(n746bar)
  );
  //OR U215
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U215 (
    .O(n746),
    .I0(n745),
    .I1(n744)
  );
  //AND U215bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U215bar (
    .O(n746bar),
    .I0(n745bar),
    .I1(n744bar)
  );
  //OR U216
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U216 (
    .O(n744),
    .I0(in[136]),
    .I1(in[121])
  );
  //AND U216bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U216bar (
    .O(n744bar),
    .I0(inbar[136]),
    .I1(inbar[121])
  );
  //OR U217
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U217 (
    .O(n745),
    .I0(in[186]),
    .I1(in[174])
  );
  //AND U217bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U217bar (
    .O(n745bar),
    .I0(inbar[186]),
    .I1(inbar[174])
  );
  //OR U218
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U218 (
    .O(n747),
    .I0(n743),
    .I1(n742)
  );
  //AND U218bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U218bar (
    .O(n747bar),
    .I0(n743bar),
    .I1(n742bar)
  );
  //OR U219
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U219 (
    .O(n742),
    .I0(in[198]),
    .I1(in[197])
  );
  //AND U219bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U219bar (
    .O(n742bar),
    .I0(inbar[198]),
    .I1(inbar[197])
  );
  //OR U220
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U220 (
    .O(n743),
    .I0(in[214]),
    .I1(in[199])
  );
  //AND U220bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U220bar (
    .O(n743bar),
    .I0(inbar[214]),
    .I1(inbar[199])
  );
  //OR U221
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U221 (
    .O(n749),
    .I0(n741),
    .I1(n740)
  );
  //AND U221bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U221bar (
    .O(n749bar),
    .I0(n741bar),
    .I1(n740bar)
  );
  //OR U222
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U222 (
    .O(n740),
    .I0(n739),
    .I1(n738)
  );
  //AND U222bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U222bar (
    .O(n740bar),
    .I0(n739bar),
    .I1(n738bar)
  );
  //OR U223
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U223 (
    .O(n738),
    .I0(in[231]),
    .I1(in[220])
  );
  //AND U223bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U223bar (
    .O(n738bar),
    .I0(inbar[231]),
    .I1(inbar[220])
  );
  //OR U224
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U224 (
    .O(n739),
    .I0(in_25),
    .I1(in[245])
  );
  //AND U224bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U224bar (
    .O(n739bar),
    .I0(in_25bar),
    .I1(inbar[245])
  );
  //OR U225
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U225 (
    .O(n741),
    .I0(n737),
    .I1(n736)
  );
  //AND U225bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U225bar (
    .O(n741bar),
    .I0(n737bar),
    .I1(n736bar)
  );
  //OR U226
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U226 (
    .O(n736),
    .I0(in_53),
    .I1(in_29)
  );
  //AND U226bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U226bar (
    .O(n736bar),
    .I0(in_53bar),
    .I1(in_29bar)
  );
  //OR U227
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U227 (
    .O(n737),
    .I0(in_79),
    .I1(in_74)
  );
  //AND U227bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U227bar (
    .O(n737bar),
    .I0(in_79bar),
    .I1(in_74bar)
  );
  //OR U228
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U228 (
    .O(n789),
    .I0(n735),
    .I1(n734)
  );
  //AND U228bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U228bar (
    .O(n789bar),
    .I0(n735bar),
    .I1(n734bar)
  );
  //OR U229
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U229 (
    .O(n734),
    .I0(in[152]),
    .I1(in[140])
  );
  //AND U229bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U229bar (
    .O(n734bar),
    .I0(inbar[152]),
    .I1(inbar[140])
  );
  //OR U230
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U230 (
    .O(n735),
    .I0(in[155]),
    .I1(n733)
  );
  //AND U230bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U230bar (
    .O(n735bar),
    .I0(inbar[155]),
    .I1(n733bar)
  );
  //OR U231
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U231 (
    .O(n733),
    .I0(in[166]),
    .I1(in[165])
  );
  //AND U231bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U231bar (
    .O(n733bar),
    .I0(inbar[166]),
    .I1(inbar[165])
  );
  //OR U232
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U232 (
    .O(n791),
    .I0(n732),
    .I1(n731)
  );
  //AND U232bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U232bar (
    .O(n791bar),
    .I0(n732bar),
    .I1(n731bar)
  );
  //OR U233
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U233 (
    .O(n731),
    .I0(n730),
    .I1(n729)
  );
  //AND U233bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U233bar (
    .O(n731bar),
    .I0(n730bar),
    .I1(n729bar)
  );
  //OR U234
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U234 (
    .O(n729),
    .I0(in[202]),
    .I1(in[185])
  );
  //AND U234bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U234bar (
    .O(n729bar),
    .I0(inbar[202]),
    .I1(inbar[185])
  );
  //OR U235
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U235 (
    .O(n730),
    .I0(in[211]),
    .I1(n728)
  );
  //AND U235bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U235bar (
    .O(n730bar),
    .I0(inbar[211]),
    .I1(n728bar)
  );
  //OR U236
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U236 (
    .O(n728),
    .I0(in[255]),
    .I1(in[253])
  );
  //AND U236bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U236bar (
    .O(n728bar),
    .I0(inbar[255]),
    .I1(inbar[253])
  );
  //OR U237
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U237 (
    .O(n732),
    .I0(n727),
    .I1(n726)
  );
  //AND U237bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U237bar (
    .O(n732bar),
    .I0(n727bar),
    .I1(n726bar)
  );
  //OR U238
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U238 (
    .O(n726),
    .I0(in_35),
    .I1(in_15)
  );
  //AND U238bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U238bar (
    .O(n726bar),
    .I0(in_35bar),
    .I1(in_15bar)
  );
  //OR U239
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U239 (
    .O(n727),
    .I0(in_36),
    .I1(n725)
  );
  //AND U239bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U239bar (
    .O(n727bar),
    .I0(in_36bar),
    .I1(n725bar)
  );
  //OR U240
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U240 (
    .O(n725),
    .I0(in_48),
    .I1(in_40)
  );
  //AND U240bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U240bar (
    .O(n725bar),
    .I0(in_48bar),
    .I1(in_40bar)
  );
  //OR U241
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U241 (
    .O(out[1]),
    .I0(n724),
    .I1(n723)
  );
  //AND U241bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U241bar (
    .O(outbar[1]),
    .I0(n724bar),
    .I1(n723bar)
  );
  //OR U242
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U242 (
    .O(n723),
    .I0(n722),
    .I1(n721)
  );
  //AND U242bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U242bar (
    .O(n723bar),
    .I0(n722bar),
    .I1(n721bar)
  );
  //OR U243
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U243 (
    .O(n721),
    .I0(n720),
    .I1(n719)
  );
  //AND U243bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U243bar (
    .O(n721bar),
    .I0(n720bar),
    .I1(n719bar)
  );
  //OR U244
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U244 (
    .O(n719),
    .I0(n921),
    .I1(n887)
  );
  //AND U244bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U244bar (
    .O(n719bar),
    .I0(n921bar),
    .I1(n887bar)
  );
  //OR U245
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U245 (
    .O(n887),
    .I0(n718),
    .I1(n717)
  );
  //AND U245bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U245bar (
    .O(n887bar),
    .I0(n718bar),
    .I1(n717bar)
  );
  //OR U246
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U246 (
    .O(n717),
    .I0(n716),
    .I1(n715)
  );
  //AND U246bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U246bar (
    .O(n717bar),
    .I0(n716bar),
    .I1(n715bar)
  );
  //OR U247
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U247 (
    .O(n715),
    .I0(n714),
    .I1(n713)
  );
  //AND U247bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U247bar (
    .O(n715bar),
    .I0(n714bar),
    .I1(n713bar)
  );
  //OR U248
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U248 (
    .O(n713),
    .I0(in[116]),
    .I1(in[110])
  );
  //AND U248bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U248bar (
    .O(n713bar),
    .I0(inbar[116]),
    .I1(inbar[110])
  );
  //OR U249
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U249 (
    .O(n714),
    .I0(in[133]),
    .I1(in[130])
  );
  //AND U249bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U249bar (
    .O(n714bar),
    .I0(inbar[133]),
    .I1(inbar[130])
  );
  //OR U250
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U250 (
    .O(n716),
    .I0(n712),
    .I1(n711)
  );
  //AND U250bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U250bar (
    .O(n716bar),
    .I0(n712bar),
    .I1(n711bar)
  );
  //OR U251
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U251 (
    .O(n711),
    .I0(in[203]),
    .I1(in[135])
  );
  //AND U251bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U251bar (
    .O(n711bar),
    .I0(inbar[203]),
    .I1(inbar[135])
  );
  //OR U252
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U252 (
    .O(n712),
    .I0(in[232]),
    .I1(in[223])
  );
  //AND U252bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U252bar (
    .O(n712bar),
    .I0(inbar[232]),
    .I1(inbar[223])
  );
  //OR U253
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U253 (
    .O(n718),
    .I0(n710),
    .I1(n709)
  );
  //AND U253bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U253bar (
    .O(n718bar),
    .I0(n710bar),
    .I1(n709bar)
  );
  //OR U254
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U254 (
    .O(n709),
    .I0(n708),
    .I1(n707)
  );
  //AND U254bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U254bar (
    .O(n709bar),
    .I0(n708bar),
    .I1(n707bar)
  );
  //OR U255
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U255 (
    .O(n707),
    .I0(in[255]),
    .I1(in[233])
  );
  //AND U255bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U255bar (
    .O(n707bar),
    .I0(inbar[255]),
    .I1(inbar[233])
  );
  //OR U256
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U256 (
    .O(n708),
    .I0(in_53),
    .I1(in_34)
  );
  //AND U256bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U256bar (
    .O(n708bar),
    .I0(in_53bar),
    .I1(in_34bar)
  );
  //OR U257
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U257 (
    .O(n710),
    .I0(n706),
    .I1(n705)
  );
  //AND U257bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U257bar (
    .O(n710bar),
    .I0(n706bar),
    .I1(n705bar)
  );
  //OR U258
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U258 (
    .O(n705),
    .I0(in_57),
    .I1(in_55)
  );
  //AND U258bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U258bar (
    .O(n705bar),
    .I0(in_57bar),
    .I1(in_55bar)
  );
  //OR U259
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U259 (
    .O(n706),
    .I0(in_68),
    .I1(in_67)
  );
  //AND U259bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U259bar (
    .O(n706bar),
    .I0(in_68bar),
    .I1(in_67bar)
  );
  //OR U260
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U260 (
    .O(n921),
    .I0(n704),
    .I1(n703)
  );
  //AND U260bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U260bar (
    .O(n921bar),
    .I0(n704bar),
    .I1(n703bar)
  );
  //OR U261
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U261 (
    .O(n703),
    .I0(n702),
    .I1(n701)
  );
  //AND U261bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U261bar (
    .O(n703bar),
    .I0(n702bar),
    .I1(n701bar)
  );
  //OR U262
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U262 (
    .O(n701),
    .I0(n700),
    .I1(n699)
  );
  //AND U262bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U262bar (
    .O(n701bar),
    .I0(n700bar),
    .I1(n699bar)
  );
  //OR U263
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U263 (
    .O(n699),
    .I0(n944),
    .I1(n872)
  );
  //AND U263bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U263bar (
    .O(n699bar),
    .I0(n944bar),
    .I1(n872bar)
  );
  //OR U264
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U264 (
    .O(n872),
    .I0(n698),
    .I1(n697)
  );
  //AND U264bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U264bar (
    .O(n872bar),
    .I0(n698bar),
    .I1(n697bar)
  );
  //OR U265
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U265 (
    .O(n697),
    .I0(n696),
    .I1(n695)
  );
  //AND U265bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U265bar (
    .O(n697bar),
    .I0(n696bar),
    .I1(n695bar)
  );
  //OR U266
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U266 (
    .O(n695),
    .I0(n694),
    .I1(n693)
  );
  //AND U266bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U266bar (
    .O(n695bar),
    .I0(n694bar),
    .I1(n693bar)
  );
  //OR U267
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U267 (
    .O(n693),
    .I0(in[121]),
    .I1(in[102])
  );
  //AND U267bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U267bar (
    .O(n693bar),
    .I0(inbar[121]),
    .I1(inbar[102])
  );
  //OR U268
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U268 (
    .O(n694),
    .I0(in[162]),
    .I1(in[161])
  );
  //AND U268bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U268bar (
    .O(n694bar),
    .I0(inbar[162]),
    .I1(inbar[161])
  );
  //OR U269
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U269 (
    .O(n696),
    .I0(n692),
    .I1(n691)
  );
  //AND U269bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U269bar (
    .O(n696bar),
    .I0(n692bar),
    .I1(n691bar)
  );
  //OR U270
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U270 (
    .O(n691),
    .I0(in[192]),
    .I1(in[178])
  );
  //AND U270bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U270bar (
    .O(n691bar),
    .I0(inbar[192]),
    .I1(inbar[178])
  );
  //OR U271
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U271 (
    .O(n692),
    .I0(in[244]),
    .I1(in[209])
  );
  //AND U271bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U271bar (
    .O(n692bar),
    .I0(inbar[244]),
    .I1(inbar[209])
  );
  //OR U272
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U272 (
    .O(n698),
    .I0(n690),
    .I1(n689)
  );
  //AND U272bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U272bar (
    .O(n698bar),
    .I0(n690bar),
    .I1(n689bar)
  );
  //OR U273
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U273 (
    .O(n689),
    .I0(n688),
    .I1(n687)
  );
  //AND U273bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U273bar (
    .O(n689bar),
    .I0(n688bar),
    .I1(n687bar)
  );
  //OR U274
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U274 (
    .O(n687),
    .I0(in[90]),
    .I1(in[254])
  );
  //AND U274bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U274bar (
    .O(n687bar),
    .I0(inbar[90]),
    .I1(inbar[254])
  );
  //OR U275
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U275 (
    .O(n688),
    .I0(in_36),
    .I1(in_32)
  );
  //AND U275bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U275bar (
    .O(n688bar),
    .I0(in_36bar),
    .I1(in_32bar)
  );
  //OR U276
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U276 (
    .O(n690),
    .I0(n686),
    .I1(n685)
  );
  //AND U276bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U276bar (
    .O(n690bar),
    .I0(n686bar),
    .I1(n685bar)
  );
  //OR U277
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U277 (
    .O(n685),
    .I0(in_62),
    .I1(in_37)
  );
  //AND U277bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U277bar (
    .O(n685bar),
    .I0(in_62bar),
    .I1(in_37bar)
  );
  //OR U278
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U278 (
    .O(n686),
    .I0(in_75),
    .I1(in_73)
  );
  //AND U278bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U278bar (
    .O(n686bar),
    .I0(in_75bar),
    .I1(in_73bar)
  );
  //OR U279
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U279 (
    .O(n944),
    .I0(n684),
    .I1(n683)
  );
  //AND U279bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U279bar (
    .O(n944bar),
    .I0(n684bar),
    .I1(n683bar)
  );
  //OR U280
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U280 (
    .O(n683),
    .I0(n682),
    .I1(n681)
  );
  //AND U280bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U280bar (
    .O(n683bar),
    .I0(n682bar),
    .I1(n681bar)
  );
  //OR U281
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U281 (
    .O(n681),
    .I0(n680),
    .I1(n679)
  );
  //AND U281bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U281bar (
    .O(n681bar),
    .I0(n680bar),
    .I1(n679bar)
  );
  //OR U282
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U282 (
    .O(n679),
    .I0(in[171]),
    .I1(in[153])
  );
  //AND U282bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U282bar (
    .O(n679bar),
    .I0(inbar[171]),
    .I1(inbar[153])
  );
  //OR U283
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U283 (
    .O(n680),
    .I0(in[187]),
    .I1(in[176])
  );
  //AND U283bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U283bar (
    .O(n680bar),
    .I0(inbar[187]),
    .I1(inbar[176])
  );
  //OR U284
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U284 (
    .O(n682),
    .I0(n678),
    .I1(n677)
  );
  //AND U284bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U284bar (
    .O(n682bar),
    .I0(n678bar),
    .I1(n677bar)
  );
  //OR U285
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U285 (
    .O(n677),
    .I0(in[245]),
    .I1(in[211])
  );
  //AND U285bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U285bar (
    .O(n677bar),
    .I0(inbar[245]),
    .I1(inbar[211])
  );
  //OR U286
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U286 (
    .O(n678),
    .I0(in[97]),
    .I1(in[88])
  );
  //AND U286bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U286bar (
    .O(n678bar),
    .I0(inbar[97]),
    .I1(inbar[88])
  );
  //OR U287
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U287 (
    .O(n684),
    .I0(n676),
    .I1(n675)
  );
  //AND U287bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U287bar (
    .O(n684bar),
    .I0(n676bar),
    .I1(n675bar)
  );
  //OR U288
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U288 (
    .O(n675),
    .I0(n674),
    .I1(n673)
  );
  //AND U288bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U288bar (
    .O(n675bar),
    .I0(n674bar),
    .I1(n673bar)
  );
  //OR U289
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U289 (
    .O(n673),
    .I0(in_10),
    .I1(in_0)
  );
  //AND U289bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U289bar (
    .O(n673bar),
    .I0(in_10bar),
    .I1(in_0bar)
  );
  //OR U290
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U290 (
    .O(n674),
    .I0(in_59),
    .I1(in_5)
  );
  //AND U290bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U290bar (
    .O(n674bar),
    .I0(in_59bar),
    .I1(in_5bar)
  );
  //OR U291
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U291 (
    .O(n676),
    .I0(n672),
    .I1(n671)
  );
  //AND U291bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U291bar (
    .O(n676bar),
    .I0(n672bar),
    .I1(n671bar)
  );
  //OR U292
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U292 (
    .O(n671),
    .I0(in_60),
    .I1(in_6)
  );
  //AND U292bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U292bar (
    .O(n671bar),
    .I0(in_60bar),
    .I1(in_6bar)
  );
  //OR U293
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U293 (
    .O(n672),
    .I0(in_77),
    .I1(in_69)
  );
  //AND U293bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U293bar (
    .O(n672bar),
    .I0(in_77bar),
    .I1(in_69bar)
  );
  //OR U294
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U294 (
    .O(n700),
    .I0(in[113]),
    .I1(n864)
  );
  //AND U294bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U294bar (
    .O(n700bar),
    .I0(inbar[113]),
    .I1(n864bar)
  );
  //OR U295
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U295 (
    .O(n864),
    .I0(n670),
    .I1(n669)
  );
  //AND U295bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U295bar (
    .O(n864bar),
    .I0(n670bar),
    .I1(n669bar)
  );
  //OR U296
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U296 (
    .O(n669),
    .I0(n668),
    .I1(n667)
  );
  //AND U296bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U296bar (
    .O(n669bar),
    .I0(n668bar),
    .I1(n667bar)
  );
  //OR U297
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U297 (
    .O(n667),
    .I0(n666),
    .I1(n665)
  );
  //AND U297bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U297bar (
    .O(n667bar),
    .I0(n666bar),
    .I1(n665bar)
  );
  //OR U298
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U298 (
    .O(n665),
    .I0(in[125]),
    .I1(in[107])
  );
  //AND U298bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U298bar (
    .O(n665bar),
    .I0(inbar[125]),
    .I1(inbar[107])
  );
  //OR U299
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U299 (
    .O(n666),
    .I0(in[138]),
    .I1(in[126])
  );
  //AND U299bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U299bar (
    .O(n666bar),
    .I0(inbar[138]),
    .I1(inbar[126])
  );
  //OR U300
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U300 (
    .O(n668),
    .I0(n664),
    .I1(n663)
  );
  //AND U300bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U300bar (
    .O(n668bar),
    .I0(n664bar),
    .I1(n663bar)
  );
  //OR U301
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U301 (
    .O(n663),
    .I0(in[189]),
    .I1(in[143])
  );
  //AND U301bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U301bar (
    .O(n663bar),
    .I0(inbar[189]),
    .I1(inbar[143])
  );
  //OR U302
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U302 (
    .O(n664),
    .I0(in[99]),
    .I1(in[214])
  );
  //AND U302bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U302bar (
    .O(n664bar),
    .I0(inbar[99]),
    .I1(inbar[214])
  );
  //OR U303
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U303 (
    .O(n670),
    .I0(n662),
    .I1(n661)
  );
  //AND U303bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U303bar (
    .O(n670bar),
    .I0(n662bar),
    .I1(n661bar)
  );
  //OR U304
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U304 (
    .O(n661),
    .I0(n660),
    .I1(n659)
  );
  //AND U304bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U304bar (
    .O(n661bar),
    .I0(n660bar),
    .I1(n659bar)
  );
  //OR U305
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U305 (
    .O(n659),
    .I0(in_15),
    .I1(in_12)
  );
  //AND U305bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U305bar (
    .O(n659bar),
    .I0(in_15bar),
    .I1(in_12bar)
  );
  //OR U306
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U306 (
    .O(n660),
    .I0(in_20),
    .I1(in_2)
  );
  //AND U306bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U306bar (
    .O(n660bar),
    .I0(in_20bar),
    .I1(in_2bar)
  );
  //OR U307
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U307 (
    .O(n662),
    .I0(n658),
    .I1(n657)
  );
  //AND U307bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U307bar (
    .O(n662bar),
    .I0(n658bar),
    .I1(n657bar)
  );
  //OR U308
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U308 (
    .O(n657),
    .I0(in_30),
    .I1(in_3)
  );
  //AND U308bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U308bar (
    .O(n657bar),
    .I0(in_30bar),
    .I1(in_3bar)
  );
  //OR U309
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U309 (
    .O(n658),
    .I0(in_4),
    .I1(in_38)
  );
  //AND U309bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U309bar (
    .O(n658bar),
    .I0(in_4bar),
    .I1(in_38bar)
  );
  //OR U310
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U310 (
    .O(n702),
    .I0(n656),
    .I1(n655)
  );
  //AND U310bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U310bar (
    .O(n702bar),
    .I0(n656bar),
    .I1(n655bar)
  );
  //OR U311
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U311 (
    .O(n655),
    .I0(in[148]),
    .I1(in[137])
  );
  //AND U311bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U311bar (
    .O(n655bar),
    .I0(inbar[148]),
    .I1(inbar[137])
  );
  //OR U312
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U312 (
    .O(n656),
    .I0(in[149]),
    .I1(n654)
  );
  //AND U312bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U312bar (
    .O(n656bar),
    .I0(inbar[149]),
    .I1(n654bar)
  );
  //OR U313
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U313 (
    .O(n654),
    .I0(in[195]),
    .I1(in[190])
  );
  //AND U313bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U313bar (
    .O(n654bar),
    .I0(inbar[195]),
    .I1(inbar[190])
  );
  //OR U314
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U314 (
    .O(n704),
    .I0(n653),
    .I1(n652)
  );
  //AND U314bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U314bar (
    .O(n704bar),
    .I0(n653bar),
    .I1(n652bar)
  );
  //OR U315
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U315 (
    .O(n652),
    .I0(n651),
    .I1(n650)
  );
  //AND U315bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U315bar (
    .O(n652bar),
    .I0(n651bar),
    .I1(n650bar)
  );
  //OR U316
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U316 (
    .O(n650),
    .I0(in[98]),
    .I1(in[197])
  );
  //AND U316bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U316bar (
    .O(n650bar),
    .I0(inbar[98]),
    .I1(inbar[197])
  );
  //OR U317
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U317 (
    .O(n651),
    .I0(in_11),
    .I1(n649)
  );
  //AND U317bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U317bar (
    .O(n651bar),
    .I0(in_11bar),
    .I1(n649bar)
  );
  //OR U318
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U318 (
    .O(n649),
    .I0(in_26),
    .I1(in_14)
  );
  //AND U318bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U318bar (
    .O(n649bar),
    .I0(in_26bar),
    .I1(in_14bar)
  );
  //OR U319
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U319 (
    .O(n653),
    .I0(n648),
    .I1(n647)
  );
  //AND U319bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U319bar (
    .O(n653bar),
    .I0(n648bar),
    .I1(n647bar)
  );
  //OR U320
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U320 (
    .O(n647),
    .I0(in_35),
    .I1(in_27)
  );
  //AND U320bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U320bar (
    .O(n647bar),
    .I0(in_35bar),
    .I1(in_27bar)
  );
  //OR U321
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U321 (
    .O(n648),
    .I0(in_50),
    .I1(n646)
  );
  //AND U321bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U321bar (
    .O(n648bar),
    .I0(in_50bar),
    .I1(n646bar)
  );
  //OR U322
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U322 (
    .O(n646),
    .I0(in_78),
    .I1(in_61)
  );
  //AND U322bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U322bar (
    .O(n646bar),
    .I0(in_78bar),
    .I1(in_61bar)
  );
  //OR U323
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U323 (
    .O(n720),
    .I0(n942),
    .I1(n645)
  );
  //AND U323bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U323bar (
    .O(n720bar),
    .I0(n942bar),
    .I1(n645bar)
  );
  //OR U324
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U324 (
    .O(n645),
    .I0(in[106]),
    .I1(n863)
  );
  //AND U324bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U324bar (
    .O(n645bar),
    .I0(inbar[106]),
    .I1(n863bar)
  );
  //OR U325
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U325 (
    .O(n863),
    .I0(n644),
    .I1(n643)
  );
  //AND U325bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U325bar (
    .O(n863bar),
    .I0(n644bar),
    .I1(n643bar)
  );
  //OR U326
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U326 (
    .O(n643),
    .I0(n642),
    .I1(n641)
  );
  //AND U326bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U326bar (
    .O(n643bar),
    .I0(n642bar),
    .I1(n641bar)
  );
  //OR U327
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U327 (
    .O(n641),
    .I0(n640),
    .I1(n639)
  );
  //AND U327bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U327bar (
    .O(n641bar),
    .I0(n640bar),
    .I1(n639bar)
  );
  //OR U328
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U328 (
    .O(n639),
    .I0(in[127]),
    .I1(in[122])
  );
  //AND U328bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U328bar (
    .O(n639bar),
    .I0(inbar[127]),
    .I1(inbar[122])
  );
  //OR U329
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U329 (
    .O(n640),
    .I0(in[156]),
    .I1(in[132])
  );
  //AND U329bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U329bar (
    .O(n640bar),
    .I0(inbar[156]),
    .I1(inbar[132])
  );
  //OR U330
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U330 (
    .O(n642),
    .I0(n638),
    .I1(n637)
  );
  //AND U330bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U330bar (
    .O(n642bar),
    .I0(n638bar),
    .I1(n637bar)
  );
  //OR U331
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U331 (
    .O(n637),
    .I0(in[159]),
    .I1(in[157])
  );
  //AND U331bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U331bar (
    .O(n637bar),
    .I0(inbar[159]),
    .I1(inbar[157])
  );
  //OR U332
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U332 (
    .O(n638),
    .I0(in[185]),
    .I1(in[169])
  );
  //AND U332bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U332bar (
    .O(n638bar),
    .I0(inbar[185]),
    .I1(inbar[169])
  );
  //OR U333
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U333 (
    .O(n644),
    .I0(n636),
    .I1(n635)
  );
  //AND U333bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U333bar (
    .O(n644bar),
    .I0(n636bar),
    .I1(n635bar)
  );
  //OR U334
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U334 (
    .O(n635),
    .I0(n634),
    .I1(n633)
  );
  //AND U334bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U334bar (
    .O(n635bar),
    .I0(n634bar),
    .I1(n633bar)
  );
  //OR U335
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U335 (
    .O(n633),
    .I0(in[239]),
    .I1(in[218])
  );
  //AND U335bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U335bar (
    .O(n633bar),
    .I0(inbar[239]),
    .I1(inbar[218])
  );
  //OR U336
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U336 (
    .O(n634),
    .I0(in_13),
    .I1(in[87])
  );
  //AND U336bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U336bar (
    .O(n634bar),
    .I0(in_13bar),
    .I1(inbar[87])
  );
  //OR U337
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U337 (
    .O(n636),
    .I0(n632),
    .I1(n631)
  );
  //AND U337bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U337bar (
    .O(n636bar),
    .I0(n632bar),
    .I1(n631bar)
  );
  //OR U338
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U338 (
    .O(n631),
    .I0(in_72),
    .I1(in_70)
  );
  //AND U338bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U338bar (
    .O(n631bar),
    .I0(in_72bar),
    .I1(in_70bar)
  );
  //OR U339
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U339 (
    .O(n632),
    .I0(in_80),
    .I1(in_74)
  );
  //AND U339bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U339bar (
    .O(n632bar),
    .I0(in_80bar),
    .I1(in_74bar)
  );
  //OR U340
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U340 (
    .O(n942),
    .I0(n630),
    .I1(n629)
  );
  //AND U340bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U340bar (
    .O(n942bar),
    .I0(n630bar),
    .I1(n629bar)
  );
  //OR U341
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U341 (
    .O(n629),
    .I0(n628),
    .I1(n627)
  );
  //AND U341bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U341bar (
    .O(n629bar),
    .I0(n628bar),
    .I1(n627bar)
  );
  //OR U342
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U342 (
    .O(n627),
    .I0(n626),
    .I1(n625)
  );
  //AND U342bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U342bar (
    .O(n627bar),
    .I0(n626bar),
    .I1(n625bar)
  );
  //OR U343
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U343 (
    .O(n625),
    .I0(in[146]),
    .I1(in[100])
  );
  //AND U343bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U343bar (
    .O(n625bar),
    .I0(inbar[146]),
    .I1(inbar[100])
  );
  //OR U344
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U344 (
    .O(n626),
    .I0(in[168]),
    .I1(in[152])
  );
  //AND U344bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U344bar (
    .O(n626bar),
    .I0(inbar[168]),
    .I1(inbar[152])
  );
  //OR U345
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U345 (
    .O(n628),
    .I0(n624),
    .I1(n623)
  );
  //AND U345bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U345bar (
    .O(n628bar),
    .I0(n624bar),
    .I1(n623bar)
  );
  //OR U346
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U346 (
    .O(n623),
    .I0(in[199]),
    .I1(in[182])
  );
  //AND U346bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U346bar (
    .O(n623bar),
    .I0(inbar[199]),
    .I1(inbar[182])
  );
  //OR U347
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U347 (
    .O(n624),
    .I0(in[236]),
    .I1(in[204])
  );
  //AND U347bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U347bar (
    .O(n624bar),
    .I0(inbar[236]),
    .I1(inbar[204])
  );
  //OR U348
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U348 (
    .O(n630),
    .I0(n622),
    .I1(n621)
  );
  //AND U348bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U348bar (
    .O(n630bar),
    .I0(n622bar),
    .I1(n621bar)
  );
  //OR U349
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U349 (
    .O(n621),
    .I0(n620),
    .I1(n619)
  );
  //AND U349bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U349bar (
    .O(n621bar),
    .I0(n620bar),
    .I1(n619bar)
  );
  //OR U350
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U350 (
    .O(n619),
    .I0(in[89]),
    .I1(in[246])
  );
  //AND U350bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U350bar (
    .O(n619bar),
    .I0(inbar[89]),
    .I1(inbar[246])
  );
  //OR U351
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U351 (
    .O(n620),
    .I0(in[95]),
    .I1(in[92])
  );
  //AND U351bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U351bar (
    .O(n620bar),
    .I0(inbar[95]),
    .I1(inbar[92])
  );
  //OR U352
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U352 (
    .O(n622),
    .I0(n618),
    .I1(n617)
  );
  //AND U352bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U352bar (
    .O(n622bar),
    .I0(n618bar),
    .I1(n617bar)
  );
  //OR U353
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U353 (
    .O(n617),
    .I0(in_22),
    .I1(in_16)
  );
  //AND U353bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U353bar (
    .O(n617bar),
    .I0(in_22bar),
    .I1(in_16bar)
  );
  //OR U354
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U354 (
    .O(n618),
    .I0(in_51),
    .I1(in_49)
  );
  //AND U354bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U354bar (
    .O(n618bar),
    .I0(in_51bar),
    .I1(in_49bar)
  );
  //OR U355
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U355 (
    .O(n722),
    .I0(n616),
    .I1(n615)
  );
  //AND U355bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U355bar (
    .O(n722bar),
    .I0(n616bar),
    .I1(n615bar)
  );
  //OR U356
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U356 (
    .O(n615),
    .I0(in[158]),
    .I1(in[115])
  );
  //AND U356bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U356bar (
    .O(n615bar),
    .I0(inbar[158]),
    .I1(inbar[115])
  );
  //OR U357
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U357 (
    .O(n616),
    .I0(in[163]),
    .I1(n614)
  );
  //AND U357bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U357bar (
    .O(n616bar),
    .I0(inbar[163]),
    .I1(n614bar)
  );
  //OR U358
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U358 (
    .O(n614),
    .I0(in[206]),
    .I1(in[165])
  );
  //AND U358bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U358bar (
    .O(n614bar),
    .I0(inbar[206]),
    .I1(inbar[165])
  );
  //OR U359
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U359 (
    .O(n724),
    .I0(n613),
    .I1(n612)
  );
  //AND U359bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U359bar (
    .O(n724bar),
    .I0(n613bar),
    .I1(n612bar)
  );
  //OR U360
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U360 (
    .O(n612),
    .I0(n611),
    .I1(n610)
  );
  //AND U360bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U360bar (
    .O(n612bar),
    .I0(n611bar),
    .I1(n610bar)
  );
  //OR U361
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U361 (
    .O(n610),
    .I0(in[213]),
    .I1(in[207])
  );
  //AND U361bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U361bar (
    .O(n610bar),
    .I0(inbar[213]),
    .I1(inbar[207])
  );
  //OR U362
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U362 (
    .O(n611),
    .I0(in[215]),
    .I1(n609)
  );
  //AND U362bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U362bar (
    .O(n611bar),
    .I0(inbar[215]),
    .I1(n609bar)
  );
  //OR U363
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U363 (
    .O(n609),
    .I0(in[230]),
    .I1(in[220])
  );
  //AND U363bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U363bar (
    .O(n609bar),
    .I0(inbar[230]),
    .I1(inbar[220])
  );
  //OR U364
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U364 (
    .O(n613),
    .I0(n608),
    .I1(n607)
  );
  //AND U364bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U364bar (
    .O(n613bar),
    .I0(n608bar),
    .I1(n607bar)
  );
  //OR U365
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U365 (
    .O(n607),
    .I0(in[251]),
    .I1(in[234])
  );
  //AND U365bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U365bar (
    .O(n607bar),
    .I0(inbar[251]),
    .I1(inbar[234])
  );
  //OR U366
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U366 (
    .O(n608),
    .I0(in_17),
    .I1(n606)
  );
  //AND U366bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U366bar (
    .O(n608bar),
    .I0(in_17bar),
    .I1(n606bar)
  );
  //OR U367
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U367 (
    .O(n606),
    .I0(in_65),
    .I1(in_56)
  );
  //AND U367bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U367bar (
    .O(n606bar),
    .I0(in_65bar),
    .I1(in_56bar)
  );
  //OR U368
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U368 (
    .O(out[0]),
    .I0(n605),
    .I1(n604)
  );
  //AND U368bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U368bar (
    .O(outbar[0]),
    .I0(n605bar),
    .I1(n604bar)
  );
  //OR U369
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U369 (
    .O(n604),
    .I0(n603),
    .I1(n602)
  );
  //AND U369bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U369bar (
    .O(n604bar),
    .I0(n603bar),
    .I1(n602bar)
  );
  //OR U370
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U370 (
    .O(n602),
    .I0(n601),
    .I1(n600)
  );
  //AND U370bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U370bar (
    .O(n602bar),
    .I0(n601bar),
    .I1(n600bar)
  );
  //OR U371
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U371 (
    .O(n600),
    .I0(n820),
    .I1(n785)
  );
  //AND U371bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U371bar (
    .O(n600bar),
    .I0(n820bar),
    .I1(n785bar)
  );
  //OR U372
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U372 (
    .O(n785),
    .I0(n599),
    .I1(n598)
  );
  //AND U372bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U372bar (
    .O(n785bar),
    .I0(n599bar),
    .I1(n598bar)
  );
  //OR U373
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U373 (
    .O(n598),
    .I0(n597),
    .I1(n596)
  );
  //AND U373bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U373bar (
    .O(n598bar),
    .I0(n597bar),
    .I1(n596bar)
  );
  //OR U374
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U374 (
    .O(n596),
    .I0(n595),
    .I1(n594)
  );
  //AND U374bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U374bar (
    .O(n596bar),
    .I0(n595bar),
    .I1(n594bar)
  );
  //OR U375
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U375 (
    .O(n594),
    .I0(in[135]),
    .I1(in[104])
  );
  //AND U375bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U375bar (
    .O(n594bar),
    .I0(inbar[135]),
    .I1(inbar[104])
  );
  //OR U376
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U376 (
    .O(n595),
    .I0(in[188]),
    .I1(in[178])
  );
  //AND U376bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U376bar (
    .O(n595bar),
    .I0(inbar[188]),
    .I1(inbar[178])
  );
  //OR U377
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U377 (
    .O(n597),
    .I0(n593),
    .I1(n592)
  );
  //AND U377bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U377bar (
    .O(n597bar),
    .I0(n593bar),
    .I1(n592bar)
  );
  //OR U378
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U378 (
    .O(n592),
    .I0(in[217]),
    .I1(in[194])
  );
  //AND U378bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U378bar (
    .O(n592bar),
    .I0(inbar[217]),
    .I1(inbar[194])
  );
  //OR U379
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U379 (
    .O(n593),
    .I0(in[237]),
    .I1(in[218])
  );
  //AND U379bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U379bar (
    .O(n593bar),
    .I0(inbar[237]),
    .I1(inbar[218])
  );
  //OR U380
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U380 (
    .O(n599),
    .I0(n591),
    .I1(n590)
  );
  //AND U380bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U380bar (
    .O(n599bar),
    .I0(n591bar),
    .I1(n590bar)
  );
  //OR U381
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U381 (
    .O(n590),
    .I0(n589),
    .I1(n588)
  );
  //AND U381bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U381bar (
    .O(n590bar),
    .I0(n589bar),
    .I1(n588bar)
  );
  //OR U382
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U382 (
    .O(n588),
    .I0(in_2),
    .I1(in_10)
  );
  //AND U382bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U382bar (
    .O(n588bar),
    .I0(in_2bar),
    .I1(in_10bar)
  );
  //OR U383
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U383 (
    .O(n589),
    .I0(in_47),
    .I1(in_22)
  );
  //AND U383bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U383bar (
    .O(n589bar),
    .I0(in_47bar),
    .I1(in_22bar)
  );
  //OR U384
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U384 (
    .O(n591),
    .I0(n587),
    .I1(n586)
  );
  //AND U384bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U384bar (
    .O(n591bar),
    .I0(n587bar),
    .I1(n586bar)
  );
  //OR U385
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U385 (
    .O(n586),
    .I0(in_56),
    .I1(in_54)
  );
  //AND U385bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U385bar (
    .O(n586bar),
    .I0(in_56bar),
    .I1(in_54bar)
  );
  //OR U386
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U386 (
    .O(n587),
    .I0(in_63),
    .I1(in_61)
  );
  //AND U386bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U386bar (
    .O(n587bar),
    .I0(in_63bar),
    .I1(in_61bar)
  );
  //OR U387
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U387 (
    .O(n820),
    .I0(n585),
    .I1(n584)
  );
  //AND U387bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U387bar (
    .O(n820bar),
    .I0(n585bar),
    .I1(n584bar)
  );
  //OR U388
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U388 (
    .O(n584),
    .I0(n583),
    .I1(n582)
  );
  //AND U388bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U388bar (
    .O(n584bar),
    .I0(n583bar),
    .I1(n582bar)
  );
  //OR U389
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U389 (
    .O(n582),
    .I0(n581),
    .I1(n580)
  );
  //AND U389bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U389bar (
    .O(n582bar),
    .I0(n581bar),
    .I1(n580bar)
  );
  //OR U390
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U390 (
    .O(n580),
    .I0(in[158]),
    .I1(in[142])
  );
  //AND U390bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U390bar (
    .O(n580bar),
    .I0(inbar[158]),
    .I1(inbar[142])
  );
  //OR U391
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U391 (
    .O(n581),
    .I0(in[175]),
    .I1(in[164])
  );
  //AND U391bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U391bar (
    .O(n581bar),
    .I0(inbar[175]),
    .I1(inbar[164])
  );
  //OR U392
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U392 (
    .O(n583),
    .I0(n579),
    .I1(n578)
  );
  //AND U392bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U392bar (
    .O(n583bar),
    .I0(n579bar),
    .I1(n578bar)
  );
  //OR U393
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U393 (
    .O(n578),
    .I0(in[228]),
    .I1(in[204])
  );
  //AND U393bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U393bar (
    .O(n578bar),
    .I0(inbar[228]),
    .I1(inbar[204])
  );
  //OR U394
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U394 (
    .O(n579),
    .I0(in[91]),
    .I1(in[87])
  );
  //AND U394bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U394bar (
    .O(n579bar),
    .I0(inbar[91]),
    .I1(inbar[87])
  );
  //OR U395
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U395 (
    .O(n585),
    .I0(n577),
    .I1(n576)
  );
  //AND U395bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U395bar (
    .O(n585bar),
    .I0(n577bar),
    .I1(n576bar)
  );
  //OR U396
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U396 (
    .O(n576),
    .I0(n575),
    .I1(n574)
  );
  //AND U396bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U396bar (
    .O(n576bar),
    .I0(n575bar),
    .I1(n574bar)
  );
  //OR U397
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U397 (
    .O(n574),
    .I0(in_21),
    .I1(in_11)
  );
  //AND U397bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U397bar (
    .O(n574bar),
    .I0(in_21bar),
    .I1(in_11bar)
  );
  //OR U398
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U398 (
    .O(n575),
    .I0(in_5),
    .I1(in_3)
  );
  //AND U398bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U398bar (
    .O(n575bar),
    .I0(in_5bar),
    .I1(in_3bar)
  );
  //OR U399
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U399 (
    .O(n577),
    .I0(n573),
    .I1(n572)
  );
  //AND U399bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U399bar (
    .O(n577bar),
    .I0(n573bar),
    .I1(n572bar)
  );
  //OR U400
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U400 (
    .O(n572),
    .I0(in_68),
    .I1(in_64)
  );
  //AND U400bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U400bar (
    .O(n572bar),
    .I0(in_68bar),
    .I1(in_64bar)
  );
  //OR U401
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U401 (
    .O(n573),
    .I0(in_76),
    .I1(in_73)
  );
  //AND U401bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U401bar (
    .O(n573bar),
    .I0(in_76bar),
    .I1(in_73bar)
  );
  //OR U402
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U402 (
    .O(n601),
    .I0(n778),
    .I1(n571)
  );
  //AND U402bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U402bar (
    .O(n601bar),
    .I0(n778bar),
    .I1(n571bar)
  );
  //OR U403
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U403 (
    .O(n571),
    .I0(in[100]),
    .I1(n965)
  );
  //AND U403bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U403bar (
    .O(n571bar),
    .I0(inbar[100]),
    .I1(n965bar)
  );
  //OR U404
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U404 (
    .O(n965),
    .I0(n570),
    .I1(n569)
  );
  //AND U404bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U404bar (
    .O(n965bar),
    .I0(n570bar),
    .I1(n569bar)
  );
  //OR U405
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U405 (
    .O(n569),
    .I0(n568),
    .I1(n567)
  );
  //AND U405bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U405bar (
    .O(n569bar),
    .I0(n568bar),
    .I1(n567bar)
  );
  //OR U406
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U406 (
    .O(n567),
    .I0(n566),
    .I1(n565)
  );
  //AND U406bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U406bar (
    .O(n567bar),
    .I0(n566bar),
    .I1(n565bar)
  );
  //OR U407
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U407 (
    .O(n565),
    .I0(n817),
    .I1(n750)
  );
  //AND U407bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U407bar (
    .O(n565bar),
    .I0(n817bar),
    .I1(n750bar)
  );
  //OR U408
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U408 (
    .O(n750),
    .I0(n564),
    .I1(n563)
  );
  //AND U408bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U408bar (
    .O(n750bar),
    .I0(n564bar),
    .I1(n563bar)
  );
  //OR U409
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U409 (
    .O(n563),
    .I0(n562),
    .I1(n561)
  );
  //AND U409bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U409bar (
    .O(n563bar),
    .I0(n562bar),
    .I1(n561bar)
  );
  //OR U410
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U410 (
    .O(n561),
    .I0(n560),
    .I1(n559)
  );
  //AND U410bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U410bar (
    .O(n561bar),
    .I0(n560bar),
    .I1(n559bar)
  );
  //OR U411
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U411 (
    .O(n559),
    .I0(in[119]),
    .I1(in[103])
  );
  //AND U411bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U411bar (
    .O(n559bar),
    .I0(inbar[119]),
    .I1(inbar[103])
  );
  //OR U412
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U412 (
    .O(n560),
    .I0(in[137]),
    .I1(in[133])
  );
  //AND U412bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U412bar (
    .O(n560bar),
    .I0(inbar[137]),
    .I1(inbar[133])
  );
  //OR U413
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U413 (
    .O(n562),
    .I0(n558),
    .I1(n557)
  );
  //AND U413bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U413bar (
    .O(n562bar),
    .I0(n558bar),
    .I1(n557bar)
  );
  //OR U414
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U414 (
    .O(n557),
    .I0(in[176]),
    .I1(in[173])
  );
  //AND U414bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U414bar (
    .O(n557bar),
    .I0(inbar[176]),
    .I1(inbar[173])
  );
  //OR U415
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U415 (
    .O(n558),
    .I0(in[210]),
    .I1(in[181])
  );
  //AND U415bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U415bar (
    .O(n558bar),
    .I0(inbar[210]),
    .I1(inbar[181])
  );
  //OR U416
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U416 (
    .O(n564),
    .I0(n556),
    .I1(n555)
  );
  //AND U416bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U416bar (
    .O(n564bar),
    .I0(n556bar),
    .I1(n555bar)
  );
  //OR U417
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U417 (
    .O(n555),
    .I0(n554),
    .I1(n553)
  );
  //AND U417bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U417bar (
    .O(n555bar),
    .I0(n554bar),
    .I1(n553bar)
  );
  //OR U418
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U418 (
    .O(n553),
    .I0(in_13),
    .I1(in[234])
  );
  //AND U418bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U418bar (
    .O(n553bar),
    .I0(in_13bar),
    .I1(inbar[234])
  );
  //OR U419
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U419 (
    .O(n554),
    .I0(in_38),
    .I1(in_32)
  );
  //AND U419bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U419bar (
    .O(n554bar),
    .I0(in_38bar),
    .I1(in_32bar)
  );
  //OR U420
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U420 (
    .O(n556),
    .I0(n552),
    .I1(n551)
  );
  //AND U420bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U420bar (
    .O(n556bar),
    .I0(n552bar),
    .I1(n551bar)
  );
  //OR U421
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U421 (
    .O(n551),
    .I0(in_42),
    .I1(in_41)
  );
  //AND U421bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U421bar (
    .O(n551bar),
    .I0(in_42bar),
    .I1(in_41bar)
  );
  //OR U422
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U422 (
    .O(n552),
    .I0(in_7),
    .I1(in_49)
  );
  //AND U422bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U422bar (
    .O(n552bar),
    .I0(in_7bar),
    .I1(in_49bar)
  );
  //OR U423
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U423 (
    .O(n817),
    .I0(n550),
    .I1(n549)
  );
  //AND U423bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U423bar (
    .O(n817bar),
    .I0(n550bar),
    .I1(n549bar)
  );
  //OR U424
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U424 (
    .O(n549),
    .I0(n548),
    .I1(n547)
  );
  //AND U424bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U424bar (
    .O(n549bar),
    .I0(n548bar),
    .I1(n547bar)
  );
  //OR U425
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U425 (
    .O(n547),
    .I0(n546),
    .I1(n545)
  );
  //AND U425bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U425bar (
    .O(n547bar),
    .I0(n546bar),
    .I1(n545bar)
  );
  //OR U426
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U426 (
    .O(n545),
    .I0(in[159]),
    .I1(in[105])
  );
  //AND U426bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U426bar (
    .O(n545bar),
    .I0(inbar[159]),
    .I1(inbar[105])
  );
  //OR U427
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U427 (
    .O(n546),
    .I0(in[206]),
    .I1(in[183])
  );
  //AND U427bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U427bar (
    .O(n546bar),
    .I0(inbar[206]),
    .I1(inbar[183])
  );
  //OR U428
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U428 (
    .O(n548),
    .I0(n544),
    .I1(n543)
  );
  //AND U428bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U428bar (
    .O(n548bar),
    .I0(n544bar),
    .I1(n543bar)
  );
  //OR U429
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U429 (
    .O(n543),
    .I0(in[229]),
    .I1(in[219])
  );
  //AND U429bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U429bar (
    .O(n543bar),
    .I0(inbar[229]),
    .I1(inbar[219])
  );
  //OR U430
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U430 (
    .O(n544),
    .I0(in[235]),
    .I1(in[232])
  );
  //AND U430bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U430bar (
    .O(n544bar),
    .I0(inbar[235]),
    .I1(inbar[232])
  );
  //OR U431
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U431 (
    .O(n550),
    .I0(n542),
    .I1(n541)
  );
  //AND U431bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U431bar (
    .O(n550bar),
    .I0(n542bar),
    .I1(n541bar)
  );
  //OR U432
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U432 (
    .O(n541),
    .I0(n540),
    .I1(n539)
  );
  //AND U432bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U432bar (
    .O(n541bar),
    .I0(n540bar),
    .I1(n539bar)
  );
  //OR U433
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U433 (
    .O(n539),
    .I0(in[249]),
    .I1(in[242])
  );
  //AND U433bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U433bar (
    .O(n539bar),
    .I0(inbar[249]),
    .I1(inbar[242])
  );
  //OR U434
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U434 (
    .O(n540),
    .I0(in[89]),
    .I1(in[254])
  );
  //AND U434bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U434bar (
    .O(n540bar),
    .I0(inbar[89]),
    .I1(inbar[254])
  );
  //OR U435
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U435 (
    .O(n542),
    .I0(n538),
    .I1(n537)
  );
  //AND U435bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U435bar (
    .O(n542bar),
    .I0(n538bar),
    .I1(n537bar)
  );
  //OR U436
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U436 (
    .O(n537),
    .I0(in_14),
    .I1(in[99])
  );
  //AND U436bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U436bar (
    .O(n537bar),
    .I0(in_14bar),
    .I1(inbar[99])
  );
  //OR U437
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U437 (
    .O(n538),
    .I0(in_60),
    .I1(in_18)
  );
  //AND U437bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U437bar (
    .O(n538bar),
    .I0(in_60bar),
    .I1(in_18bar)
  );
  //OR U438
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U438 (
    .O(n566),
    .I0(in[113]),
    .I1(n763)
  );
  //AND U438bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U438bar (
    .O(n566bar),
    .I0(inbar[113]),
    .I1(n763bar)
  );
  //OR U439
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U439 (
    .O(n763),
    .I0(n536),
    .I1(n535)
  );
  //AND U439bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U439bar (
    .O(n763bar),
    .I0(n536bar),
    .I1(n535bar)
  );
  //OR U440
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U440 (
    .O(n535),
    .I0(n534),
    .I1(n533)
  );
  //AND U440bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U440bar (
    .O(n535bar),
    .I0(n534bar),
    .I1(n533bar)
  );
  //OR U441
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U441 (
    .O(n533),
    .I0(n532),
    .I1(n531)
  );
  //AND U441bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U441bar (
    .O(n533bar),
    .I0(n532bar),
    .I1(n531bar)
  );
  //OR U442
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U442 (
    .O(n531),
    .I0(in[115]),
    .I1(in[110])
  );
  //AND U442bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U442bar (
    .O(n531bar),
    .I0(inbar[115]),
    .I1(inbar[110])
  );
  //OR U443
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U443 (
    .O(n532),
    .I0(in[125]),
    .I1(in[117])
  );
  //AND U443bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U443bar (
    .O(n532bar),
    .I0(inbar[125]),
    .I1(inbar[117])
  );
  //OR U444
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U444 (
    .O(n534),
    .I0(n530),
    .I1(n529)
  );
  //AND U444bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U444bar (
    .O(n534bar),
    .I0(n530bar),
    .I1(n529bar)
  );
  //OR U445
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U445 (
    .O(n529),
    .I0(in[180]),
    .I1(in[128])
  );
  //AND U445bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U445bar (
    .O(n529bar),
    .I0(inbar[180]),
    .I1(inbar[128])
  );
  //OR U446
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U446 (
    .O(n530),
    .I0(in[205]),
    .I1(in[201])
  );
  //AND U446bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U446bar (
    .O(n530bar),
    .I0(inbar[205]),
    .I1(inbar[201])
  );
  //OR U447
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U447 (
    .O(n536),
    .I0(n528),
    .I1(n527)
  );
  //AND U447bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U447bar (
    .O(n536bar),
    .I0(n528bar),
    .I1(n527bar)
  );
  //OR U448
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U448 (
    .O(n527),
    .I0(n526),
    .I1(n525)
  );
  //AND U448bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U448bar (
    .O(n527bar),
    .I0(n526bar),
    .I1(n525bar)
  );
  //OR U449
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U449 (
    .O(n525),
    .I0(in[244]),
    .I1(in[239])
  );
  //AND U449bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U449bar (
    .O(n525bar),
    .I0(inbar[244]),
    .I1(inbar[239])
  );
  //OR U450
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U450 (
    .O(n526),
    .I0(in[95]),
    .I1(in[83])
  );
  //AND U450bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U450bar (
    .O(n526bar),
    .I0(inbar[95]),
    .I1(inbar[83])
  );
  //OR U451
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U451 (
    .O(n528),
    .I0(n524),
    .I1(n523)
  );
  //AND U451bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U451bar (
    .O(n528bar),
    .I0(n524bar),
    .I1(n523bar)
  );
  //OR U452
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U452 (
    .O(n523),
    .I0(in_24),
    .I1(in[97])
  );
  //AND U452bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U452bar (
    .O(n523bar),
    .I0(in_24bar),
    .I1(inbar[97])
  );
  //OR U453
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U453 (
    .O(n524),
    .I0(in_33),
    .I1(in_27)
  );
  //AND U453bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U453bar (
    .O(n524bar),
    .I0(in_33bar),
    .I1(in_27bar)
  );
  //OR U454
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U454 (
    .O(n568),
    .I0(n522),
    .I1(n521)
  );
  //AND U454bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U454bar (
    .O(n568bar),
    .I0(n522bar),
    .I1(n521bar)
  );
  //OR U455
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U455 (
    .O(n521),
    .I0(in[145]),
    .I1(in[126])
  );
  //AND U455bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U455bar (
    .O(n521bar),
    .I0(inbar[145]),
    .I1(inbar[126])
  );
  //OR U456
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U456 (
    .O(n522),
    .I0(in[169]),
    .I1(n520)
  );
  //AND U456bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U456bar (
    .O(n522bar),
    .I0(inbar[169]),
    .I1(n520bar)
  );
  //OR U457
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U457 (
    .O(n520),
    .I0(in[221]),
    .I1(in[172])
  );
  //AND U457bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U457bar (
    .O(n520bar),
    .I0(inbar[221]),
    .I1(inbar[172])
  );
  //OR U458
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U458 (
    .O(n570),
    .I0(n519),
    .I1(n518)
  );
  //AND U458bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U458bar (
    .O(n570bar),
    .I0(n519bar),
    .I1(n518bar)
  );
  //OR U459
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U459 (
    .O(n518),
    .I0(n517),
    .I1(n516)
  );
  //AND U459bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U459bar (
    .O(n518bar),
    .I0(n517bar),
    .I1(n516bar)
  );
  //OR U460
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U460 (
    .O(n516),
    .I0(in[241]),
    .I1(in[224])
  );
  //AND U460bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U460bar (
    .O(n516bar),
    .I0(inbar[241]),
    .I1(inbar[224])
  );
  //OR U461
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U461 (
    .O(n517),
    .I0(in[86]),
    .I1(n515)
  );
  //AND U461bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U461bar (
    .O(n517bar),
    .I0(inbar[86]),
    .I1(n515bar)
  );
  //OR U462
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U462 (
    .O(n515),
    .I0(in_43),
    .I1(in_34)
  );
  //AND U462bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U462bar (
    .O(n515bar),
    .I0(in_43bar),
    .I1(in_34bar)
  );
  //OR U463
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U463 (
    .O(n519),
    .I0(n514),
    .I1(n513)
  );
  //AND U463bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U463bar (
    .O(n519bar),
    .I0(n514bar),
    .I1(n513bar)
  );
  //OR U464
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U464 (
    .O(n513),
    .I0(in_65),
    .I1(in_51)
  );
  //AND U464bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U464bar (
    .O(n513bar),
    .I0(in_65bar),
    .I1(in_51bar)
  );
  //OR U465
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U465 (
    .O(n514),
    .I0(in_75),
    .I1(n512)
  );
  //AND U465bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U465bar (
    .O(n514bar),
    .I0(in_75bar),
    .I1(n512bar)
  );
  //OR U466
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U466 (
    .O(n512),
    .I0(in_81),
    .I1(in_77)
  );
  //AND U466bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U466bar (
    .O(n512bar),
    .I0(in_81bar),
    .I1(in_77bar)
  );
  //OR U467
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U467 (
    .O(n778),
    .I0(n511),
    .I1(n510)
  );
  //AND U467bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U467bar (
    .O(n778bar),
    .I0(n511bar),
    .I1(n510bar)
  );
  //OR U468
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U468 (
    .O(n510),
    .I0(n509),
    .I1(n508)
  );
  //AND U468bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U468bar (
    .O(n510bar),
    .I0(n509bar),
    .I1(n508bar)
  );
  //OR U469
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U469 (
    .O(n508),
    .I0(n507),
    .I1(n506)
  );
  //AND U469bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U469bar (
    .O(n508bar),
    .I0(n507bar),
    .I1(n506bar)
  );
  //OR U470
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U470 (
    .O(n506),
    .I0(in[107]),
    .I1(in[101])
  );
  //AND U470bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U470bar (
    .O(n506bar),
    .I0(inbar[107]),
    .I1(inbar[101])
  );
  //OR U471
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U471 (
    .O(n507),
    .I0(in[139]),
    .I1(in[132])
  );
  //AND U471bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U471bar (
    .O(n507bar),
    .I0(inbar[139]),
    .I1(inbar[132])
  );
  //OR U472
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U472 (
    .O(n509),
    .I0(n505),
    .I1(n504)
  );
  //AND U472bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U472bar (
    .O(n509bar),
    .I0(n505bar),
    .I1(n504bar)
  );
  //OR U473
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U473 (
    .O(n504),
    .I0(in[146]),
    .I1(in[141])
  );
  //AND U473bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U473bar (
    .O(n504bar),
    .I0(inbar[146]),
    .I1(inbar[141])
  );
  //OR U474
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U474 (
    .O(n505),
    .I0(in[203]),
    .I1(in[179])
  );
  //AND U474bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U474bar (
    .O(n505bar),
    .I0(inbar[203]),
    .I1(inbar[179])
  );
  //OR U475
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U475 (
    .O(n511),
    .I0(n503),
    .I1(n502)
  );
  //AND U475bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U475bar (
    .O(n511bar),
    .I0(n503bar),
    .I1(n502bar)
  );
  //OR U476
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U476 (
    .O(n502),
    .I0(n501),
    .I1(n500)
  );
  //AND U476bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U476bar (
    .O(n502bar),
    .I0(n501bar),
    .I1(n500bar)
  );
  //OR U477
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U477 (
    .O(n500),
    .I0(in[243]),
    .I1(in[222])
  );
  //AND U477bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U477bar (
    .O(n500bar),
    .I0(inbar[243]),
    .I1(inbar[222])
  );
  //OR U478
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U478 (
    .O(n501),
    .I0(in[251]),
    .I1(in[250])
  );
  //AND U478bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U478bar (
    .O(n501bar),
    .I0(inbar[251]),
    .I1(inbar[250])
  );
  //OR U479
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U479 (
    .O(n503),
    .I0(n499),
    .I1(n498)
  );
  //AND U479bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U479bar (
    .O(n503bar),
    .I0(n499bar),
    .I1(n498bar)
  );
  //OR U480
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U480 (
    .O(n498),
    .I0(in_37),
    .I1(in_19)
  );
  //AND U480bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U480bar (
    .O(n498bar),
    .I0(in_37bar),
    .I1(in_19bar)
  );
  //OR U481
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U481 (
    .O(n499),
    .I0(in_78),
    .I1(in_6)
  );
  //AND U481bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U481bar (
    .O(n499bar),
    .I0(in_78bar),
    .I1(in_6bar)
  );
  //OR U482
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U482 (
    .O(n603),
    .I0(n497),
    .I1(n496)
  );
  //AND U482bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U482bar (
    .O(n603bar),
    .I0(n497bar),
    .I1(n496bar)
  );
  //OR U483
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U483 (
    .O(n496),
    .I0(in[112]),
    .I1(in[102])
  );
  //AND U483bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U483bar (
    .O(n496bar),
    .I0(inbar[112]),
    .I1(inbar[102])
  );
  //OR U484
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U484 (
    .O(n497),
    .I0(in[123]),
    .I1(n495)
  );
  //AND U484bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U484bar (
    .O(n497bar),
    .I0(inbar[123]),
    .I1(n495bar)
  );
  //OR U485
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U485 (
    .O(n495),
    .I0(in[143]),
    .I1(in[130])
  );
  //AND U485bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U485bar (
    .O(n495bar),
    .I0(inbar[143]),
    .I1(inbar[130])
  );
  //OR U486
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U486 (
    .O(n605),
    .I0(n494),
    .I1(n493)
  );
  //AND U486bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U486bar (
    .O(n605bar),
    .I0(n494bar),
    .I1(n493bar)
  );
  //OR U487
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U487 (
    .O(n493),
    .I0(n492),
    .I1(n491)
  );
  //AND U487bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U487bar (
    .O(n493bar),
    .I0(n492bar),
    .I1(n491bar)
  );
  //OR U488
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U488 (
    .O(n491),
    .I0(in[216]),
    .I1(in[213])
  );
  //AND U488bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U488bar (
    .O(n491bar),
    .I0(inbar[216]),
    .I1(inbar[213])
  );
  //OR U489
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U489 (
    .O(n492),
    .I0(in[227]),
    .I1(n490)
  );
  //AND U489bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U489bar (
    .O(n492bar),
    .I0(inbar[227]),
    .I1(n490bar)
  );
  //OR U490
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U490 (
    .O(n490),
    .I0(in_0),
    .I1(in[248])
  );
  //AND U490bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U490bar (
    .O(n490bar),
    .I0(in_0bar),
    .I1(inbar[248])
  );
  //OR U491
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U491 (
    .O(n494),
    .I0(n489),
    .I1(n488)
  );
  //AND U491bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U491bar (
    .O(n494bar),
    .I0(n489bar),
    .I1(n488bar)
  );
  //OR U492
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U492 (
    .O(n488),
    .I0(in_46),
    .I1(in_44)
  );
  //AND U492bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U492bar (
    .O(n488bar),
    .I0(in_46bar),
    .I1(in_44bar)
  );
  //OR U493
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U493 (
    .O(n489),
    .I0(in_50),
    .I1(n487)
  );
  //AND U493bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U493bar (
    .O(n489bar),
    .I0(in_50bar),
    .I1(n487bar)
  );
  //OR U494
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U494 (
    .O(n487),
    .I0(in_9),
    .I1(in_80)
  );
  //AND U494bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U494bar (
    .O(n487bar),
    .I0(in_9bar),
    .I1(in_80bar)
  );
endmodule

module sBox_15 ( in, out );

  input wire [7:0] in;
//input_done

  output wire [7:0] out;
//output_done

  wire [255:0] decodeOut;
//wire_done

  decode_15 dec ( .in(in), .out(decodeOut) );
  encode_15 enc ( .in(decodeOut), .out(out) );
endmodule

module s_box_LUT ( in, out );

  input wire [127:0] in;
//input_done

  output [127:0] out;
//output_done

//wire_done

  sBox_15 s0 ( .in(in[127:120]), .out(out[127:120]) );
  sBox_14 s1 ( .in(in[119:112]), .out(out[119:112]) );
  sBox_13 s2 ( .in(in[111:104]), .out(out[111:104]) );
  sBox_12 s3 ( .in(in[103:96]), .out(out[103:96]) );
  sBox_11 s4 ( .in(in[95:88]), .out(out[95:88]) );
  sBox_10 s5 ( .in(in[87:80]), .out(out[87:80]) );
  sBox_9 s6 ( .in(in[79:72]), .out(out[79:72]) );
  sBox_8 s7 ( .in(in[71:64]), .out(out[71:64]) );
  sBox_7 s8 ( .in(in[63:56]), .out(out[63:56]) );
  sBox_6 s9 ( .in(in[55:48]), .out(out[55:48]) );
  sBox_5 s10 ( .in(in[47:40]), .out(out[47:40]) );
  sBox_4 s11 ( .in(in[39:32]), .out(out[39:32]) );
  sBox_3 s12 ( .in(in[31:24]), .out(out[31:24]) );
  sBox_2 s13 ( .in(in[23:16]), .out(out[23:16]) );
  sBox_1 s14 ( .in(in[15:8]), .out(out[15:8]) );
  sBox_0 s15 ( .in(in[7:0]), .out(out[7:0]) );
endmodule

//done
