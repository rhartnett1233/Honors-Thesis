`timescale 1ns / 1ps


module addRoundKey_Precharge_LUT ( data, databar, key, out, outbar );

  input wire [127:0] data;
  input wire [127:0] key;
  input wire [127:0] databar;
  wire [127:0] keybar;
  assign keybar[0] = ~key[0];
  assign keybar[1] = ~key[1];
  assign keybar[2] = ~key[2];
  assign keybar[3] = ~key[3];
  assign keybar[4] = ~key[4];
  assign keybar[5] = ~key[5];
  assign keybar[6] = ~key[6];
  assign keybar[7] = ~key[7];
  assign keybar[8] = ~key[8];
  assign keybar[9] = ~key[9];
  assign keybar[10] = ~key[10];
  assign keybar[11] = ~key[11];
  assign keybar[12] = ~key[12];
  assign keybar[13] = ~key[13];
  assign keybar[14] = ~key[14];
  assign keybar[15] = ~key[15];
  assign keybar[16] = ~key[16];
  assign keybar[17] = ~key[17];
  assign keybar[18] = ~key[18];
  assign keybar[19] = ~key[19];
  assign keybar[20] = ~key[20];
  assign keybar[21] = ~key[21];
  assign keybar[22] = ~key[22];
  assign keybar[23] = ~key[23];
  assign keybar[24] = ~key[24];
  assign keybar[25] = ~key[25];
  assign keybar[26] = ~key[26];
  assign keybar[27] = ~key[27];
  assign keybar[28] = ~key[28];
  assign keybar[29] = ~key[29];
  assign keybar[30] = ~key[30];
  assign keybar[31] = ~key[31];
  assign keybar[32] = ~key[32];
  assign keybar[33] = ~key[33];
  assign keybar[34] = ~key[34];
  assign keybar[35] = ~key[35];
  assign keybar[36] = ~key[36];
  assign keybar[37] = ~key[37];
  assign keybar[38] = ~key[38];
  assign keybar[39] = ~key[39];
  assign keybar[40] = ~key[40];
  assign keybar[41] = ~key[41];
  assign keybar[42] = ~key[42];
  assign keybar[43] = ~key[43];
  assign keybar[44] = ~key[44];
  assign keybar[45] = ~key[45];
  assign keybar[46] = ~key[46];
  assign keybar[47] = ~key[47];
  assign keybar[48] = ~key[48];
  assign keybar[49] = ~key[49];
  assign keybar[50] = ~key[50];
  assign keybar[51] = ~key[51];
  assign keybar[52] = ~key[52];
  assign keybar[53] = ~key[53];
  assign keybar[54] = ~key[54];
  assign keybar[55] = ~key[55];
  assign keybar[56] = ~key[56];
  assign keybar[57] = ~key[57];
  assign keybar[58] = ~key[58];
  assign keybar[59] = ~key[59];
  assign keybar[60] = ~key[60];
  assign keybar[61] = ~key[61];
  assign keybar[62] = ~key[62];
  assign keybar[63] = ~key[63];
  assign keybar[64] = ~key[64];
  assign keybar[65] = ~key[65];
  assign keybar[66] = ~key[66];
  assign keybar[67] = ~key[67];
  assign keybar[68] = ~key[68];
  assign keybar[69] = ~key[69];
  assign keybar[70] = ~key[70];
  assign keybar[71] = ~key[71];
  assign keybar[72] = ~key[72];
  assign keybar[73] = ~key[73];
  assign keybar[74] = ~key[74];
  assign keybar[75] = ~key[75];
  assign keybar[76] = ~key[76];
  assign keybar[77] = ~key[77];
  assign keybar[78] = ~key[78];
  assign keybar[79] = ~key[79];
  assign keybar[80] = ~key[80];
  assign keybar[81] = ~key[81];
  assign keybar[82] = ~key[82];
  assign keybar[83] = ~key[83];
  assign keybar[84] = ~key[84];
  assign keybar[85] = ~key[85];
  assign keybar[86] = ~key[86];
  assign keybar[87] = ~key[87];
  assign keybar[88] = ~key[88];
  assign keybar[89] = ~key[89];
  assign keybar[90] = ~key[90];
  assign keybar[91] = ~key[91];
  assign keybar[92] = ~key[92];
  assign keybar[93] = ~key[93];
  assign keybar[94] = ~key[94];
  assign keybar[95] = ~key[95];
  assign keybar[96] = ~key[96];
  assign keybar[97] = ~key[97];
  assign keybar[98] = ~key[98];
  assign keybar[99] = ~key[99];
  assign keybar[100] = ~key[100];
  assign keybar[101] = ~key[101];
  assign keybar[102] = ~key[102];
  assign keybar[103] = ~key[103];
  assign keybar[104] = ~key[104];
  assign keybar[105] = ~key[105];
  assign keybar[106] = ~key[106];
  assign keybar[107] = ~key[107];
  assign keybar[108] = ~key[108];
  assign keybar[109] = ~key[109];
  assign keybar[110] = ~key[110];
  assign keybar[111] = ~key[111];
  assign keybar[112] = ~key[112];
  assign keybar[113] = ~key[113];
  assign keybar[114] = ~key[114];
  assign keybar[115] = ~key[115];
  assign keybar[116] = ~key[116];
  assign keybar[117] = ~key[117];
  assign keybar[118] = ~key[118];
  assign keybar[119] = ~key[119];
  assign keybar[120] = ~key[120];
  assign keybar[121] = ~key[121];
  assign keybar[122] = ~key[122];
  assign keybar[123] = ~key[123];
  assign keybar[124] = ~key[124];
  assign keybar[125] = ~key[125];
  assign keybar[126] = ~key[126];
  assign keybar[127] = ~key[127];
//input_done

  output wire [127:0] out;
  output wire [127:0] outbar;
//output_done

  wire n1;
  wire n2;
  wire n3;
  wire n4;
  wire n5;
  wire n6;
  wire n7;
  wire n8;
  wire n9;
  wire n10;
  wire n11;
  wire n12;
  wire n13;
  wire n14;
  wire n15;
  wire n16;
  wire n17;
  wire n18;
  wire n19;
  wire n20;
  wire n21;
  wire n22;
  wire n23;
  wire n24;
  wire n25;
  wire n26;
  wire n27;
  wire n28;
  wire n29;
  wire n30;
  wire n31;
  wire n32;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n1bar;
  wire n2bar;
  wire n3bar;
  wire n4bar;
  wire n5bar;
  wire n6bar;
  wire n7bar;
  wire n8bar;
  wire n9bar;
  wire n10bar;
  wire n11bar;
  wire n12bar;
  wire n13bar;
  wire n14bar;
  wire n15bar;
  wire n16bar;
  wire n17bar;
  wire n18bar;
  wire n19bar;
  wire n20bar;
  wire n21bar;
  wire n22bar;
  wire n23bar;
  wire n24bar;
  wire n25bar;
  wire n26bar;
  wire n27bar;
  wire n28bar;
  wire n29bar;
  wire n30bar;
  wire n31bar;
  wire n32bar;
  wire n33bar;
  wire n34bar;
  wire n35bar;
  wire n36bar;
  wire n37bar;
  wire n38bar;
  wire n39bar;
  wire n40bar;
  wire n41bar;
  wire n42bar;
  wire n43bar;
  wire n44bar;
  wire n45bar;
  wire n46bar;
  wire n47bar;
  wire n48bar;
  wire n49bar;
  wire n50bar;
  wire n51bar;
  wire n52bar;
  wire n53bar;
  wire n54bar;
  wire n55bar;
  wire n56bar;
  wire n57bar;
  wire n58bar;
  wire n59bar;
  wire n60bar;
  wire n61bar;
  wire n62bar;
  wire n63bar;
  wire n64bar;
  wire n65bar;
  wire n66bar;
  wire n67bar;
  wire n68bar;
  wire n69bar;
  wire n70bar;
  wire n71bar;
  wire n72bar;
  wire n73bar;
  wire n74bar;
  wire n75bar;
  wire n76bar;
  wire n77bar;
  wire n78bar;
  wire n79bar;
  wire n80bar;
  wire n81bar;
  wire n82bar;
  wire n83bar;
  wire n84bar;
  wire n85bar;
  wire n86bar;
  wire n87bar;
  wire n88bar;
  wire n89bar;
  wire n90bar;
  wire n91bar;
  wire n92bar;
  wire n93bar;
  wire n94bar;
  wire n95bar;
  wire n96bar;
  wire n97bar;
  wire n98bar;
  wire n99bar;
  wire n100bar;
  wire n101bar;
  wire n102bar;
  wire n103bar;
  wire n104bar;
  wire n105bar;
  wire n106bar;
  wire n107bar;
  wire n108bar;
  wire n109bar;
  wire n110bar;
  wire n111bar;
  wire n112bar;
  wire n113bar;
  wire n114bar;
  wire n115bar;
  wire n116bar;
  wire n117bar;
  wire n118bar;
  wire n119bar;
  wire n120bar;
  wire n121bar;
  wire n122bar;
  wire n123bar;
  wire n124bar;
  wire n125bar;
  wire n126bar;
  wire n127bar;
  wire n128bar;
  wire n129bar;
  wire n130bar;
  wire n131bar;
  wire n132bar;
  wire n133bar;
  wire n134bar;
  wire n135bar;
  wire n136bar;
  wire n137bar;
  wire n138bar;
  wire n139bar;
  wire n140bar;
  wire n141bar;
  wire n142bar;
  wire n143bar;
  wire n144bar;
  wire n145bar;
  wire n146bar;
  wire n147bar;
  wire n148bar;
  wire n149bar;
  wire n150bar;
  wire n151bar;
  wire n152bar;
  wire n153bar;
  wire n154bar;
  wire n155bar;
  wire n156bar;
  wire n157bar;
  wire n158bar;
  wire n159bar;
  wire n160bar;
  wire n161bar;
  wire n162bar;
  wire n163bar;
  wire n164bar;
  wire n165bar;
  wire n166bar;
  wire n167bar;
  wire n168bar;
  wire n169bar;
  wire n170bar;
  wire n171bar;
  wire n172bar;
  wire n173bar;
  wire n174bar;
  wire n175bar;
  wire n176bar;
  wire n177bar;
  wire n178bar;
  wire n179bar;
  wire n180bar;
  wire n181bar;
  wire n182bar;
  wire n183bar;
  wire n184bar;
  wire n185bar;
  wire n186bar;
  wire n187bar;
  wire n188bar;
  wire n189bar;
  wire n190bar;
  wire n191bar;
  wire n192bar;
  wire n193bar;
  wire n194bar;
  wire n195bar;
  wire n196bar;
  wire n197bar;
  wire n198bar;
  wire n199bar;
  wire n200bar;
  wire n201bar;
  wire n202bar;
  wire n203bar;
  wire n204bar;
  wire n205bar;
  wire n206bar;
  wire n207bar;
  wire n208bar;
  wire n209bar;
  wire n210bar;
  wire n211bar;
  wire n212bar;
  wire n213bar;
  wire n214bar;
  wire n215bar;
  wire n216bar;
  wire n217bar;
  wire n218bar;
  wire n219bar;
  wire n220bar;
  wire n221bar;
  wire n222bar;
  wire n223bar;
  wire n224bar;
  wire n225bar;
  wire n226bar;
  wire n227bar;
  wire n228bar;
  wire n229bar;
  wire n230bar;
  wire n231bar;
  wire n232bar;
  wire n233bar;
  wire n234bar;
  wire n235bar;
  wire n236bar;
  wire n237bar;
  wire n238bar;
  wire n239bar;
  wire n240bar;
  wire n241bar;
  wire n242bar;
  wire n243bar;
  wire n244bar;
  wire n245bar;
  wire n246bar;
  wire n247bar;
  wire n248bar;
  wire n249bar;
  wire n250bar;
  wire n251bar;
  wire n252bar;
  wire n253bar;
  wire n254bar;
  wire n255bar;
  wire n256bar;
  wire n257bar;
  wire n258bar;
  wire n259bar;
  wire n260bar;
  wire n261bar;
  wire n262bar;
  wire n263bar;
  wire n264bar;
  wire n265bar;
  wire n266bar;
  wire n267bar;
  wire n268bar;
  wire n269bar;
  wire n270bar;
  wire n271bar;
  wire n272bar;
  wire n273bar;
  wire n274bar;
  wire n275bar;
  wire n276bar;
  wire n277bar;
  wire n278bar;
  wire n279bar;
  wire n280bar;
  wire n281bar;
  wire n282bar;
  wire n283bar;
  wire n284bar;
  wire n285bar;
  wire n286bar;
  wire n287bar;
  wire n288bar;
  wire n289bar;
  wire n290bar;
  wire n291bar;
  wire n292bar;
  wire n293bar;
  wire n294bar;
  wire n295bar;
  wire n296bar;
  wire n297bar;
  wire n298bar;
  wire n299bar;
  wire n300bar;
  wire n301bar;
  wire n302bar;
  wire n303bar;
  wire n304bar;
  wire n305bar;
  wire n306bar;
  wire n307bar;
  wire n308bar;
  wire n309bar;
  wire n310bar;
  wire n311bar;
  wire n312bar;
  wire n313bar;
  wire n314bar;
  wire n315bar;
  wire n316bar;
  wire n317bar;
  wire n318bar;
  wire n319bar;
  wire n320bar;
  wire n321bar;
  wire n322bar;
  wire n323bar;
  wire n324bar;
  wire n325bar;
  wire n326bar;
  wire n327bar;
  wire n328bar;
  wire n329bar;
  wire n330bar;
  wire n331bar;
  wire n332bar;
  wire n333bar;
  wire n334bar;
  wire n335bar;
  wire n336bar;
  wire n337bar;
  wire n338bar;
  wire n339bar;
  wire n340bar;
  wire n341bar;
  wire n342bar;
  wire n343bar;
  wire n344bar;
  wire n345bar;
  wire n346bar;
  wire n347bar;
  wire n348bar;
  wire n349bar;
  wire n350bar;
  wire n351bar;
  wire n352bar;
  wire n353bar;
  wire n354bar;
  wire n355bar;
  wire n356bar;
  wire n357bar;
  wire n358bar;
  wire n359bar;
  wire n360bar;
  wire n361bar;
  wire n362bar;
  wire n363bar;
  wire n364bar;
  wire n365bar;
  wire n366bar;
  wire n367bar;
  wire n368bar;
  wire n369bar;
  wire n370bar;
  wire n371bar;
  wire n372bar;
  wire n373bar;
  wire n374bar;
  wire n375bar;
  wire n376bar;
  wire n377bar;
  wire n378bar;
  wire n379bar;
  wire n380bar;
  wire n381bar;
  wire n382bar;
  wire n383bar;
  wire n384bar;
  wire n385bar;
  wire n386bar;
  wire n387bar;
  wire n388bar;
  wire n389bar;
  wire n390bar;
  wire n391bar;
  wire n392bar;
  wire n393bar;
  wire n394bar;
  wire n395bar;
  wire n396bar;
  wire n397bar;
  wire n398bar;
  wire n399bar;
  wire n400bar;
  wire n401bar;
  wire n402bar;
  wire n403bar;
  wire n404bar;
  wire n405bar;
  wire n406bar;
  wire n407bar;
  wire n408bar;
  wire n409bar;
  wire n410bar;
  wire n411bar;
  wire n412bar;
  wire n413bar;
  wire n414bar;
  wire n415bar;
  wire n416bar;
  wire n417bar;
  wire n418bar;
  wire n419bar;
  wire n420bar;
  wire n421bar;
  wire n422bar;
  wire n423bar;
  wire n424bar;
  wire n425bar;
  wire n426bar;
  wire n427bar;
  wire n428bar;
  wire n429bar;
  wire n430bar;
  wire n431bar;
  wire n432bar;
  wire n433bar;
  wire n434bar;
  wire n435bar;
  wire n436bar;
  wire n437bar;
  wire n438bar;
  wire n439bar;
  wire n440bar;
  wire n441bar;
  wire n442bar;
  wire n443bar;
  wire n444bar;
  wire n445bar;
  wire n446bar;
  wire n447bar;
  wire n448bar;
  wire n449bar;
  wire n450bar;
  wire n451bar;
  wire n452bar;
  wire n453bar;
  wire n454bar;
  wire n455bar;
  wire n456bar;
  wire n457bar;
  wire n458bar;
  wire n459bar;
  wire n460bar;
  wire n461bar;
  wire n462bar;
  wire n463bar;
  wire n464bar;
  wire n465bar;
  wire n466bar;
  wire n467bar;
  wire n468bar;
  wire n469bar;
  wire n470bar;
  wire n471bar;
  wire n472bar;
  wire n473bar;
  wire n474bar;
  wire n475bar;
  wire n476bar;
  wire n477bar;
  wire n478bar;
  wire n479bar;
  wire n480bar;
  wire n481bar;
  wire n482bar;
  wire n483bar;
  wire n484bar;
  wire n485bar;
  wire n486bar;
  wire n487bar;
  wire n488bar;
  wire n489bar;
  wire n490bar;
  wire n491bar;
  wire n492bar;
  wire n493bar;
  wire n494bar;
  wire n495bar;
  wire n496bar;
  wire n497bar;
  wire n498bar;
  wire n499bar;
  wire n500bar;
  wire n501bar;
  wire n502bar;
  wire n503bar;
  wire n504bar;
  wire n505bar;
  wire n506bar;
  wire n507bar;
  wire n508bar;
  wire n509bar;
  wire n510bar;
  wire n511bar;
  wire n512bar;
//wire_done

 //assign_done

  assign n1bar = n452;
  assign n1 = n452bar;
  assign n2bar = data[127];
  assign n2 = databar[127];
  assign n3bar = n454;
  assign n3 = n454bar;
  assign n4bar = data[126];
  assign n4 = databar[126];
  assign n5bar = n456;
  assign n5 = n456bar;
  assign n6bar = data[125];
  assign n6 = databar[125];
  assign n7bar = n458;
  assign n7 = n458bar;
  assign n8bar = data[124];
  assign n8 = databar[124];
  assign n9bar = n460;
  assign n9 = n460bar;
  assign n10bar = data[123];
  assign n10 = databar[123];
  assign n11bar = n462;
  assign n11 = n462bar;
  assign n12bar = data[122];
  assign n12 = databar[122];
  assign n13bar = n464;
  assign n13 = n464bar;
  assign n14bar = data[121];
  assign n14 = databar[121];
  assign n15bar = n466;
  assign n15 = n466bar;
  assign n16bar = data[120];
  assign n16 = databar[120];
  assign n17bar = n470;
  assign n17 = n470bar;
  assign n18bar = data[119];
  assign n18 = databar[119];
  assign n19bar = n472;
  assign n19 = n472bar;
  assign n20bar = data[118];
  assign n20 = databar[118];
  assign n21bar = n474;
  assign n21 = n474bar;
  assign n22bar = data[117];
  assign n22 = databar[117];
  assign n23bar = n476;
  assign n23 = n476bar;
  assign n24bar = data[116];
  assign n24 = databar[116];
  assign n25bar = n478;
  assign n25 = n478bar;
  assign n26bar = data[115];
  assign n26 = databar[115];
  assign n27bar = n480;
  assign n27 = n480bar;
  assign n28bar = data[114];
  assign n28 = databar[114];
  assign n29bar = n482;
  assign n29 = n482bar;
  assign n30bar = data[113];
  assign n30 = databar[113];
  assign n31bar = n484;
  assign n31 = n484bar;
  assign n32bar = data[112];
  assign n32 = databar[112];
  assign n33bar = n486;
  assign n33 = n486bar;
  assign n34bar = data[111];
  assign n34 = databar[111];
  assign n35bar = n488;
  assign n35 = n488bar;
  assign n36bar = data[110];
  assign n36 = databar[110];
  assign n37bar = n492;
  assign n37 = n492bar;
  assign n38bar = data[109];
  assign n38 = databar[109];
  assign n39bar = n494;
  assign n39 = n494bar;
  assign n40bar = data[108];
  assign n40 = databar[108];
  assign n41bar = n496;
  assign n41 = n496bar;
  assign n42bar = data[107];
  assign n42 = databar[107];
  assign n43bar = n498;
  assign n43 = n498bar;
  assign n44bar = data[106];
  assign n44 = databar[106];
  assign n45bar = n500;
  assign n45 = n500bar;
  assign n46bar = data[105];
  assign n46 = databar[105];
  assign n47bar = n502;
  assign n47 = n502bar;
  assign n48bar = data[104];
  assign n48 = databar[104];
  assign n49bar = n504;
  assign n49 = n504bar;
  assign n50bar = data[103];
  assign n50 = databar[103];
  assign n51bar = n506;
  assign n51 = n506bar;
  assign n52bar = data[102];
  assign n52 = databar[102];
  assign n53bar = n508;
  assign n53 = n508bar;
  assign n54bar = data[101];
  assign n54 = databar[101];
  assign n55bar = n510;
  assign n55 = n510bar;
  assign n56bar = data[100];
  assign n56 = databar[100];
  assign n57bar = n260;
  assign n57 = n260bar;
  assign n58bar = data[99];
  assign n58 = databar[99];
  assign n59bar = n262;
  assign n59 = n262bar;
  assign n60bar = data[98];
  assign n60 = databar[98];
  assign n61bar = n264;
  assign n61 = n264bar;
  assign n62bar = data[97];
  assign n62 = databar[97];
  assign n63bar = n266;
  assign n63 = n266bar;
  assign n64bar = data[96];
  assign n64 = databar[96];
  assign n65bar = n268;
  assign n65 = n268bar;
  assign n66bar = data[95];
  assign n66 = databar[95];
  assign n67bar = n270;
  assign n67 = n270bar;
  assign n68bar = data[94];
  assign n68 = databar[94];
  assign n69bar = n272;
  assign n69 = n272bar;
  assign n70bar = data[93];
  assign n70 = databar[93];
  assign n71bar = n274;
  assign n71 = n274bar;
  assign n72bar = data[92];
  assign n72 = databar[92];
  assign n73bar = n276;
  assign n73 = n276bar;
  assign n74bar = data[91];
  assign n74 = databar[91];
  assign n75bar = n278;
  assign n75 = n278bar;
  assign n76bar = data[90];
  assign n76 = databar[90];
  assign n77bar = n282;
  assign n77 = n282bar;
  assign n78bar = data[89];
  assign n78 = databar[89];
  assign n79bar = n284;
  assign n79 = n284bar;
  assign n80bar = data[88];
  assign n80 = databar[88];
  assign n81bar = n286;
  assign n81 = n286bar;
  assign n82bar = data[87];
  assign n82 = databar[87];
  assign n83bar = n288;
  assign n83 = n288bar;
  assign n84bar = data[86];
  assign n84 = databar[86];
  assign n85bar = n290;
  assign n85 = n290bar;
  assign n86bar = data[85];
  assign n86 = databar[85];
  assign n87bar = n292;
  assign n87 = n292bar;
  assign n88bar = data[84];
  assign n88 = databar[84];
  assign n89bar = n294;
  assign n89 = n294bar;
  assign n90bar = data[83];
  assign n90 = databar[83];
  assign n91bar = n296;
  assign n91 = n296bar;
  assign n92bar = data[82];
  assign n92 = databar[82];
  assign n93bar = n298;
  assign n93 = n298bar;
  assign n94bar = data[81];
  assign n94 = databar[81];
  assign n95bar = n300;
  assign n95 = n300bar;
  assign n96bar = data[80];
  assign n96 = databar[80];
  assign n97bar = n304;
  assign n97 = n304bar;
  assign n98bar = data[79];
  assign n98 = databar[79];
  assign n99bar = n306;
  assign n99 = n306bar;
  assign n100bar = data[78];
  assign n100 = databar[78];
  assign n101bar = n308;
  assign n101 = n308bar;
  assign n102bar = data[77];
  assign n102 = databar[77];
  assign n103bar = n310;
  assign n103 = n310bar;
  assign n104bar = data[76];
  assign n104 = databar[76];
  assign n105bar = n312;
  assign n105 = n312bar;
  assign n106bar = data[75];
  assign n106 = databar[75];
  assign n107bar = n314;
  assign n107 = n314bar;
  assign n108bar = data[74];
  assign n108 = databar[74];
  assign n109bar = n316;
  assign n109 = n316bar;
  assign n110bar = data[73];
  assign n110 = databar[73];
  assign n111bar = n318;
  assign n111 = n318bar;
  assign n112bar = data[72];
  assign n112 = databar[72];
  assign n113bar = n320;
  assign n113 = n320bar;
  assign n114bar = data[71];
  assign n114 = databar[71];
  assign n115bar = n322;
  assign n115 = n322bar;
  assign n116bar = data[70];
  assign n116 = databar[70];
  assign n117bar = n326;
  assign n117 = n326bar;
  assign n118bar = data[69];
  assign n118 = databar[69];
  assign n119bar = n328;
  assign n119 = n328bar;
  assign n120bar = data[68];
  assign n120 = databar[68];
  assign n121bar = n330;
  assign n121 = n330bar;
  assign n122bar = data[67];
  assign n122 = databar[67];
  assign n123bar = n332;
  assign n123 = n332bar;
  assign n124bar = data[66];
  assign n124 = databar[66];
  assign n125bar = n334;
  assign n125 = n334bar;
  assign n126bar = data[65];
  assign n126 = databar[65];
  assign n127bar = n336;
  assign n127 = n336bar;
  assign n128bar = data[64];
  assign n128 = databar[64];
  assign n129bar = n338;
  assign n129 = n338bar;
  assign n130bar = data[63];
  assign n130 = databar[63];
  assign n131bar = n340;
  assign n131 = n340bar;
  assign n132bar = data[62];
  assign n132 = databar[62];
  assign n133bar = n342;
  assign n133 = n342bar;
  assign n134bar = data[61];
  assign n134 = databar[61];
  assign n135bar = n344;
  assign n135 = n344bar;
  assign n136bar = data[60];
  assign n136 = databar[60];
  assign n137bar = n348;
  assign n137 = n348bar;
  assign n138bar = data[59];
  assign n138 = databar[59];
  assign n139bar = n350;
  assign n139 = n350bar;
  assign n140bar = data[58];
  assign n140 = databar[58];
  assign n141bar = n352;
  assign n141 = n352bar;
  assign n142bar = data[57];
  assign n142 = databar[57];
  assign n143bar = n354;
  assign n143 = n354bar;
  assign n144bar = data[56];
  assign n144 = databar[56];
  assign n145bar = n356;
  assign n145 = n356bar;
  assign n146bar = data[55];
  assign n146 = databar[55];
  assign n147bar = n358;
  assign n147 = n358bar;
  assign n148bar = data[54];
  assign n148 = databar[54];
  assign n149bar = n360;
  assign n149 = n360bar;
  assign n150bar = data[53];
  assign n150 = databar[53];
  assign n151bar = n362;
  assign n151 = n362bar;
  assign n152bar = data[52];
  assign n152 = databar[52];
  assign n153bar = n364;
  assign n153 = n364bar;
  assign n154bar = data[51];
  assign n154 = databar[51];
  assign n155bar = n366;
  assign n155 = n366bar;
  assign n156bar = data[50];
  assign n156 = databar[50];
  assign n157bar = n370;
  assign n157 = n370bar;
  assign n158bar = data[49];
  assign n158 = databar[49];
  assign n159bar = n372;
  assign n159 = n372bar;
  assign n160bar = data[48];
  assign n160 = databar[48];
  assign n161bar = n374;
  assign n161 = n374bar;
  assign n162bar = data[47];
  assign n162 = databar[47];
  assign n163bar = n376;
  assign n163 = n376bar;
  assign n164bar = data[46];
  assign n164 = databar[46];
  assign n165bar = n378;
  assign n165 = n378bar;
  assign n166bar = data[45];
  assign n166 = databar[45];
  assign n167bar = n380;
  assign n167 = n380bar;
  assign n168bar = data[44];
  assign n168 = databar[44];
  assign n169bar = n382;
  assign n169 = n382bar;
  assign n170bar = data[43];
  assign n170 = databar[43];
  assign n171bar = n384;
  assign n171 = n384bar;
  assign n172bar = data[42];
  assign n172 = databar[42];
  assign n173bar = n386;
  assign n173 = n386bar;
  assign n174bar = data[41];
  assign n174 = databar[41];
  assign n175bar = n388;
  assign n175 = n388bar;
  assign n176bar = data[40];
  assign n176 = databar[40];
  assign n177bar = n392;
  assign n177 = n392bar;
  assign n178bar = data[39];
  assign n178 = databar[39];
  assign n179bar = n394;
  assign n179 = n394bar;
  assign n180bar = data[38];
  assign n180 = databar[38];
  assign n181bar = n396;
  assign n181 = n396bar;
  assign n182bar = data[37];
  assign n182 = databar[37];
  assign n183bar = n398;
  assign n183 = n398bar;
  assign n184bar = data[36];
  assign n184 = databar[36];
  assign n185bar = n400;
  assign n185 = n400bar;
  assign n186bar = data[35];
  assign n186 = databar[35];
  assign n187bar = n402;
  assign n187 = n402bar;
  assign n188bar = data[34];
  assign n188 = databar[34];
  assign n189bar = n404;
  assign n189 = n404bar;
  assign n190bar = data[33];
  assign n190 = databar[33];
  assign n191bar = n406;
  assign n191 = n406bar;
  assign n192bar = data[32];
  assign n192 = databar[32];
  assign n193bar = n408;
  assign n193 = n408bar;
  assign n194bar = data[31];
  assign n194 = databar[31];
  assign n195bar = n410;
  assign n195 = n410bar;
  assign n196bar = data[30];
  assign n196 = databar[30];
  assign n197bar = n414;
  assign n197 = n414bar;
  assign n198bar = data[29];
  assign n198 = databar[29];
  assign n199bar = n416;
  assign n199 = n416bar;
  assign n200bar = data[28];
  assign n200 = databar[28];
  assign n201bar = n418;
  assign n201 = n418bar;
  assign n202bar = data[27];
  assign n202 = databar[27];
  assign n203bar = n420;
  assign n203 = n420bar;
  assign n204bar = data[26];
  assign n204 = databar[26];
  assign n205bar = n422;
  assign n205 = n422bar;
  assign n206bar = data[25];
  assign n206 = databar[25];
  assign n207bar = n424;
  assign n207 = n424bar;
  assign n208bar = data[24];
  assign n208 = databar[24];
  assign n209bar = n426;
  assign n209 = n426bar;
  assign n210bar = data[23];
  assign n210 = databar[23];
  assign n211bar = n428;
  assign n211 = n428bar;
  assign n212bar = data[22];
  assign n212 = databar[22];
  assign n213bar = n430;
  assign n213 = n430bar;
  assign n214bar = data[21];
  assign n214 = databar[21];
  assign n215bar = n432;
  assign n215 = n432bar;
  assign n216bar = data[20];
  assign n216 = databar[20];
  assign n217bar = n436;
  assign n217 = n436bar;
  assign n218bar = data[19];
  assign n218 = databar[19];
  assign n219bar = n438;
  assign n219 = n438bar;
  assign n220bar = data[18];
  assign n220 = databar[18];
  assign n221bar = n440;
  assign n221 = n440bar;
  assign n222bar = data[17];
  assign n222 = databar[17];
  assign n223bar = n442;
  assign n223 = n442bar;
  assign n224bar = data[16];
  assign n224 = databar[16];
  assign n225bar = n444;
  assign n225 = n444bar;
  assign n226bar = data[15];
  assign n226 = databar[15];
  assign n227bar = n446;
  assign n227 = n446bar;
  assign n228bar = data[14];
  assign n228 = databar[14];
  assign n229bar = n448;
  assign n229 = n448bar;
  assign n230bar = data[13];
  assign n230 = databar[13];
  assign n231bar = n450;
  assign n231 = n450bar;
  assign n232bar = data[12];
  assign n232 = databar[12];
  assign n233bar = n468;
  assign n233 = n468bar;
  assign n234bar = data[11];
  assign n234 = databar[11];
  assign n235bar = n490;
  assign n235 = n490bar;
  assign n236bar = data[10];
  assign n236 = databar[10];
  assign n237bar = n258;
  assign n237 = n258bar;
  assign n238bar = data[9];
  assign n238 = databar[9];
  assign n239bar = n280;
  assign n239 = n280bar;
  assign n240bar = data[8];
  assign n240 = databar[8];
  assign n241bar = n302;
  assign n241 = n302bar;
  assign n242bar = data[7];
  assign n242 = databar[7];
  assign n243bar = n324;
  assign n243 = n324bar;
  assign n244bar = data[6];
  assign n244 = databar[6];
  assign n245bar = n346;
  assign n245 = n346bar;
  assign n246bar = data[5];
  assign n246 = databar[5];
  assign n247bar = n368;
  assign n247 = n368bar;
  assign n248bar = data[4];
  assign n248 = databar[4];
  assign n249bar = n390;
  assign n249 = n390bar;
  assign n250bar = data[3];
  assign n250 = databar[3];
  assign n251bar = n412;
  assign n251 = n412bar;
  assign n252bar = data[2];
  assign n252 = databar[2];
  assign n253bar = n434;
  assign n253 = n434bar;
  assign n254bar = data[1];
  assign n254 = databar[1];
  assign n255bar = n512;
  assign n255 = n512bar;
  assign n256bar = data[0];
  assign n256 = databar[0];
  //OR U257
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U257 (
    .O(out[9]),
    .I0(n257),
    .I1(n237)
  );
  //AND U257bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U257bar (
    .O(outbar[9]),
    .I0(n257bar),
    .I1(n237bar)
  );
  //OR U258
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U258 (
    .O(n258),
    .I0(n238),
    .I1(key[9])
  );
  //AND U258bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U258bar (
    .O(n258bar),
    .I0(n238bar),
    .I1(keybar[9])
  );
  //AND U259
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U259 (
    .O(n257),
    .I0(key[9]),
    .I1(n238)
  );
  //OR U259bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U259bar (
    .O(n257bar),
    .I0(keybar[9]),
    .I1(n238bar)
  );
  //OR U260
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U260 (
    .O(out[99]),
    .I0(n259),
    .I1(n57)
  );
  //AND U260bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U260bar (
    .O(outbar[99]),
    .I0(n259bar),
    .I1(n57bar)
  );
  //OR U261
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U261 (
    .O(n260),
    .I0(n58),
    .I1(key[99])
  );
  //AND U261bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U261bar (
    .O(n260bar),
    .I0(n58bar),
    .I1(keybar[99])
  );
  //AND U262
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U262 (
    .O(n259),
    .I0(key[99]),
    .I1(n58)
  );
  //OR U262bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U262bar (
    .O(n259bar),
    .I0(keybar[99]),
    .I1(n58bar)
  );
  //OR U263
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U263 (
    .O(out[98]),
    .I0(n261),
    .I1(n59)
  );
  //AND U263bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U263bar (
    .O(outbar[98]),
    .I0(n261bar),
    .I1(n59bar)
  );
  //OR U264
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U264 (
    .O(n262),
    .I0(n60),
    .I1(key[98])
  );
  //AND U264bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U264bar (
    .O(n262bar),
    .I0(n60bar),
    .I1(keybar[98])
  );
  //AND U265
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U265 (
    .O(n261),
    .I0(key[98]),
    .I1(n60)
  );
  //OR U265bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U265bar (
    .O(n261bar),
    .I0(keybar[98]),
    .I1(n60bar)
  );
  //OR U266
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U266 (
    .O(out[97]),
    .I0(n263),
    .I1(n61)
  );
  //AND U266bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U266bar (
    .O(outbar[97]),
    .I0(n263bar),
    .I1(n61bar)
  );
  //OR U267
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U267 (
    .O(n264),
    .I0(n62),
    .I1(key[97])
  );
  //AND U267bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U267bar (
    .O(n264bar),
    .I0(n62bar),
    .I1(keybar[97])
  );
  //AND U268
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U268 (
    .O(n263),
    .I0(key[97]),
    .I1(n62)
  );
  //OR U268bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U268bar (
    .O(n263bar),
    .I0(keybar[97]),
    .I1(n62bar)
  );
  //OR U269
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U269 (
    .O(out[96]),
    .I0(n265),
    .I1(n63)
  );
  //AND U269bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U269bar (
    .O(outbar[96]),
    .I0(n265bar),
    .I1(n63bar)
  );
  //OR U270
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U270 (
    .O(n266),
    .I0(n64),
    .I1(key[96])
  );
  //AND U270bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U270bar (
    .O(n266bar),
    .I0(n64bar),
    .I1(keybar[96])
  );
  //AND U271
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U271 (
    .O(n265),
    .I0(key[96]),
    .I1(n64)
  );
  //OR U271bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U271bar (
    .O(n265bar),
    .I0(keybar[96]),
    .I1(n64bar)
  );
  //OR U272
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U272 (
    .O(out[95]),
    .I0(n267),
    .I1(n65)
  );
  //AND U272bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U272bar (
    .O(outbar[95]),
    .I0(n267bar),
    .I1(n65bar)
  );
  //OR U273
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U273 (
    .O(n268),
    .I0(n66),
    .I1(key[95])
  );
  //AND U273bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U273bar (
    .O(n268bar),
    .I0(n66bar),
    .I1(keybar[95])
  );
  //AND U274
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U274 (
    .O(n267),
    .I0(key[95]),
    .I1(n66)
  );
  //OR U274bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U274bar (
    .O(n267bar),
    .I0(keybar[95]),
    .I1(n66bar)
  );
  //OR U275
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U275 (
    .O(out[94]),
    .I0(n269),
    .I1(n67)
  );
  //AND U275bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U275bar (
    .O(outbar[94]),
    .I0(n269bar),
    .I1(n67bar)
  );
  //OR U276
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U276 (
    .O(n270),
    .I0(n68),
    .I1(key[94])
  );
  //AND U276bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U276bar (
    .O(n270bar),
    .I0(n68bar),
    .I1(keybar[94])
  );
  //AND U277
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U277 (
    .O(n269),
    .I0(key[94]),
    .I1(n68)
  );
  //OR U277bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U277bar (
    .O(n269bar),
    .I0(keybar[94]),
    .I1(n68bar)
  );
  //OR U278
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U278 (
    .O(out[93]),
    .I0(n271),
    .I1(n69)
  );
  //AND U278bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U278bar (
    .O(outbar[93]),
    .I0(n271bar),
    .I1(n69bar)
  );
  //OR U279
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U279 (
    .O(n272),
    .I0(n70),
    .I1(key[93])
  );
  //AND U279bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U279bar (
    .O(n272bar),
    .I0(n70bar),
    .I1(keybar[93])
  );
  //AND U280
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U280 (
    .O(n271),
    .I0(key[93]),
    .I1(n70)
  );
  //OR U280bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U280bar (
    .O(n271bar),
    .I0(keybar[93]),
    .I1(n70bar)
  );
  //OR U281
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U281 (
    .O(out[92]),
    .I0(n273),
    .I1(n71)
  );
  //AND U281bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U281bar (
    .O(outbar[92]),
    .I0(n273bar),
    .I1(n71bar)
  );
  //OR U282
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U282 (
    .O(n274),
    .I0(n72),
    .I1(key[92])
  );
  //AND U282bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U282bar (
    .O(n274bar),
    .I0(n72bar),
    .I1(keybar[92])
  );
  //AND U283
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U283 (
    .O(n273),
    .I0(key[92]),
    .I1(n72)
  );
  //OR U283bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U283bar (
    .O(n273bar),
    .I0(keybar[92]),
    .I1(n72bar)
  );
  //OR U284
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U284 (
    .O(out[91]),
    .I0(n275),
    .I1(n73)
  );
  //AND U284bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U284bar (
    .O(outbar[91]),
    .I0(n275bar),
    .I1(n73bar)
  );
  //OR U285
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U285 (
    .O(n276),
    .I0(n74),
    .I1(key[91])
  );
  //AND U285bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U285bar (
    .O(n276bar),
    .I0(n74bar),
    .I1(keybar[91])
  );
  //AND U286
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U286 (
    .O(n275),
    .I0(key[91]),
    .I1(n74)
  );
  //OR U286bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U286bar (
    .O(n275bar),
    .I0(keybar[91]),
    .I1(n74bar)
  );
  //OR U287
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U287 (
    .O(out[90]),
    .I0(n277),
    .I1(n75)
  );
  //AND U287bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U287bar (
    .O(outbar[90]),
    .I0(n277bar),
    .I1(n75bar)
  );
  //OR U288
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U288 (
    .O(n278),
    .I0(n76),
    .I1(key[90])
  );
  //AND U288bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U288bar (
    .O(n278bar),
    .I0(n76bar),
    .I1(keybar[90])
  );
  //AND U289
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U289 (
    .O(n277),
    .I0(key[90]),
    .I1(n76)
  );
  //OR U289bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U289bar (
    .O(n277bar),
    .I0(keybar[90]),
    .I1(n76bar)
  );
  //OR U290
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U290 (
    .O(out[8]),
    .I0(n279),
    .I1(n239)
  );
  //AND U290bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U290bar (
    .O(outbar[8]),
    .I0(n279bar),
    .I1(n239bar)
  );
  //OR U291
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U291 (
    .O(n280),
    .I0(n240),
    .I1(key[8])
  );
  //AND U291bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U291bar (
    .O(n280bar),
    .I0(n240bar),
    .I1(keybar[8])
  );
  //AND U292
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U292 (
    .O(n279),
    .I0(key[8]),
    .I1(n240)
  );
  //OR U292bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U292bar (
    .O(n279bar),
    .I0(keybar[8]),
    .I1(n240bar)
  );
  //OR U293
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U293 (
    .O(out[89]),
    .I0(n281),
    .I1(n77)
  );
  //AND U293bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U293bar (
    .O(outbar[89]),
    .I0(n281bar),
    .I1(n77bar)
  );
  //OR U294
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U294 (
    .O(n282),
    .I0(n78),
    .I1(key[89])
  );
  //AND U294bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U294bar (
    .O(n282bar),
    .I0(n78bar),
    .I1(keybar[89])
  );
  //AND U295
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U295 (
    .O(n281),
    .I0(key[89]),
    .I1(n78)
  );
  //OR U295bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U295bar (
    .O(n281bar),
    .I0(keybar[89]),
    .I1(n78bar)
  );
  //OR U296
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U296 (
    .O(out[88]),
    .I0(n283),
    .I1(n79)
  );
  //AND U296bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U296bar (
    .O(outbar[88]),
    .I0(n283bar),
    .I1(n79bar)
  );
  //OR U297
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U297 (
    .O(n284),
    .I0(n80),
    .I1(key[88])
  );
  //AND U297bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U297bar (
    .O(n284bar),
    .I0(n80bar),
    .I1(keybar[88])
  );
  //AND U298
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U298 (
    .O(n283),
    .I0(key[88]),
    .I1(n80)
  );
  //OR U298bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U298bar (
    .O(n283bar),
    .I0(keybar[88]),
    .I1(n80bar)
  );
  //OR U299
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U299 (
    .O(out[87]),
    .I0(n285),
    .I1(n81)
  );
  //AND U299bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U299bar (
    .O(outbar[87]),
    .I0(n285bar),
    .I1(n81bar)
  );
  //OR U300
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U300 (
    .O(n286),
    .I0(n82),
    .I1(key[87])
  );
  //AND U300bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U300bar (
    .O(n286bar),
    .I0(n82bar),
    .I1(keybar[87])
  );
  //AND U301
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U301 (
    .O(n285),
    .I0(key[87]),
    .I1(n82)
  );
  //OR U301bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U301bar (
    .O(n285bar),
    .I0(keybar[87]),
    .I1(n82bar)
  );
  //OR U302
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U302 (
    .O(out[86]),
    .I0(n287),
    .I1(n83)
  );
  //AND U302bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U302bar (
    .O(outbar[86]),
    .I0(n287bar),
    .I1(n83bar)
  );
  //OR U303
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U303 (
    .O(n288),
    .I0(n84),
    .I1(key[86])
  );
  //AND U303bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U303bar (
    .O(n288bar),
    .I0(n84bar),
    .I1(keybar[86])
  );
  //AND U304
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U304 (
    .O(n287),
    .I0(key[86]),
    .I1(n84)
  );
  //OR U304bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U304bar (
    .O(n287bar),
    .I0(keybar[86]),
    .I1(n84bar)
  );
  //OR U305
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U305 (
    .O(out[85]),
    .I0(n289),
    .I1(n85)
  );
  //AND U305bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U305bar (
    .O(outbar[85]),
    .I0(n289bar),
    .I1(n85bar)
  );
  //OR U306
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U306 (
    .O(n290),
    .I0(n86),
    .I1(key[85])
  );
  //AND U306bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U306bar (
    .O(n290bar),
    .I0(n86bar),
    .I1(keybar[85])
  );
  //AND U307
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U307 (
    .O(n289),
    .I0(key[85]),
    .I1(n86)
  );
  //OR U307bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U307bar (
    .O(n289bar),
    .I0(keybar[85]),
    .I1(n86bar)
  );
  //OR U308
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U308 (
    .O(out[84]),
    .I0(n291),
    .I1(n87)
  );
  //AND U308bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U308bar (
    .O(outbar[84]),
    .I0(n291bar),
    .I1(n87bar)
  );
  //OR U309
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U309 (
    .O(n292),
    .I0(n88),
    .I1(key[84])
  );
  //AND U309bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U309bar (
    .O(n292bar),
    .I0(n88bar),
    .I1(keybar[84])
  );
  //AND U310
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U310 (
    .O(n291),
    .I0(key[84]),
    .I1(n88)
  );
  //OR U310bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U310bar (
    .O(n291bar),
    .I0(keybar[84]),
    .I1(n88bar)
  );
  //OR U311
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U311 (
    .O(out[83]),
    .I0(n293),
    .I1(n89)
  );
  //AND U311bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U311bar (
    .O(outbar[83]),
    .I0(n293bar),
    .I1(n89bar)
  );
  //OR U312
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U312 (
    .O(n294),
    .I0(n90),
    .I1(key[83])
  );
  //AND U312bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U312bar (
    .O(n294bar),
    .I0(n90bar),
    .I1(keybar[83])
  );
  //AND U313
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U313 (
    .O(n293),
    .I0(key[83]),
    .I1(n90)
  );
  //OR U313bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U313bar (
    .O(n293bar),
    .I0(keybar[83]),
    .I1(n90bar)
  );
  //OR U314
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U314 (
    .O(out[82]),
    .I0(n295),
    .I1(n91)
  );
  //AND U314bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U314bar (
    .O(outbar[82]),
    .I0(n295bar),
    .I1(n91bar)
  );
  //OR U315
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U315 (
    .O(n296),
    .I0(n92),
    .I1(key[82])
  );
  //AND U315bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U315bar (
    .O(n296bar),
    .I0(n92bar),
    .I1(keybar[82])
  );
  //AND U316
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U316 (
    .O(n295),
    .I0(key[82]),
    .I1(n92)
  );
  //OR U316bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U316bar (
    .O(n295bar),
    .I0(keybar[82]),
    .I1(n92bar)
  );
  //OR U317
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U317 (
    .O(out[81]),
    .I0(n297),
    .I1(n93)
  );
  //AND U317bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U317bar (
    .O(outbar[81]),
    .I0(n297bar),
    .I1(n93bar)
  );
  //OR U318
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U318 (
    .O(n298),
    .I0(n94),
    .I1(key[81])
  );
  //AND U318bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U318bar (
    .O(n298bar),
    .I0(n94bar),
    .I1(keybar[81])
  );
  //AND U319
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U319 (
    .O(n297),
    .I0(key[81]),
    .I1(n94)
  );
  //OR U319bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U319bar (
    .O(n297bar),
    .I0(keybar[81]),
    .I1(n94bar)
  );
  //OR U320
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U320 (
    .O(out[80]),
    .I0(n299),
    .I1(n95)
  );
  //AND U320bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U320bar (
    .O(outbar[80]),
    .I0(n299bar),
    .I1(n95bar)
  );
  //OR U321
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U321 (
    .O(n300),
    .I0(n96),
    .I1(key[80])
  );
  //AND U321bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U321bar (
    .O(n300bar),
    .I0(n96bar),
    .I1(keybar[80])
  );
  //AND U322
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U322 (
    .O(n299),
    .I0(key[80]),
    .I1(n96)
  );
  //OR U322bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U322bar (
    .O(n299bar),
    .I0(keybar[80]),
    .I1(n96bar)
  );
  //OR U323
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U323 (
    .O(out[7]),
    .I0(n301),
    .I1(n241)
  );
  //AND U323bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U323bar (
    .O(outbar[7]),
    .I0(n301bar),
    .I1(n241bar)
  );
  //OR U324
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U324 (
    .O(n302),
    .I0(n242),
    .I1(key[7])
  );
  //AND U324bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U324bar (
    .O(n302bar),
    .I0(n242bar),
    .I1(keybar[7])
  );
  //AND U325
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U325 (
    .O(n301),
    .I0(key[7]),
    .I1(n242)
  );
  //OR U325bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U325bar (
    .O(n301bar),
    .I0(keybar[7]),
    .I1(n242bar)
  );
  //OR U326
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U326 (
    .O(out[79]),
    .I0(n303),
    .I1(n97)
  );
  //AND U326bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U326bar (
    .O(outbar[79]),
    .I0(n303bar),
    .I1(n97bar)
  );
  //OR U327
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U327 (
    .O(n304),
    .I0(n98),
    .I1(key[79])
  );
  //AND U327bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U327bar (
    .O(n304bar),
    .I0(n98bar),
    .I1(keybar[79])
  );
  //AND U328
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U328 (
    .O(n303),
    .I0(key[79]),
    .I1(n98)
  );
  //OR U328bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U328bar (
    .O(n303bar),
    .I0(keybar[79]),
    .I1(n98bar)
  );
  //OR U329
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U329 (
    .O(out[78]),
    .I0(n305),
    .I1(n99)
  );
  //AND U329bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U329bar (
    .O(outbar[78]),
    .I0(n305bar),
    .I1(n99bar)
  );
  //OR U330
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U330 (
    .O(n306),
    .I0(n100),
    .I1(key[78])
  );
  //AND U330bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U330bar (
    .O(n306bar),
    .I0(n100bar),
    .I1(keybar[78])
  );
  //AND U331
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U331 (
    .O(n305),
    .I0(key[78]),
    .I1(n100)
  );
  //OR U331bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U331bar (
    .O(n305bar),
    .I0(keybar[78]),
    .I1(n100bar)
  );
  //OR U332
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U332 (
    .O(out[77]),
    .I0(n307),
    .I1(n101)
  );
  //AND U332bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U332bar (
    .O(outbar[77]),
    .I0(n307bar),
    .I1(n101bar)
  );
  //OR U333
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U333 (
    .O(n308),
    .I0(n102),
    .I1(key[77])
  );
  //AND U333bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U333bar (
    .O(n308bar),
    .I0(n102bar),
    .I1(keybar[77])
  );
  //AND U334
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U334 (
    .O(n307),
    .I0(key[77]),
    .I1(n102)
  );
  //OR U334bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U334bar (
    .O(n307bar),
    .I0(keybar[77]),
    .I1(n102bar)
  );
  //OR U335
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U335 (
    .O(out[76]),
    .I0(n309),
    .I1(n103)
  );
  //AND U335bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U335bar (
    .O(outbar[76]),
    .I0(n309bar),
    .I1(n103bar)
  );
  //OR U336
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U336 (
    .O(n310),
    .I0(n104),
    .I1(key[76])
  );
  //AND U336bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U336bar (
    .O(n310bar),
    .I0(n104bar),
    .I1(keybar[76])
  );
  //AND U337
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U337 (
    .O(n309),
    .I0(key[76]),
    .I1(n104)
  );
  //OR U337bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U337bar (
    .O(n309bar),
    .I0(keybar[76]),
    .I1(n104bar)
  );
  //OR U338
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U338 (
    .O(out[75]),
    .I0(n311),
    .I1(n105)
  );
  //AND U338bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U338bar (
    .O(outbar[75]),
    .I0(n311bar),
    .I1(n105bar)
  );
  //OR U339
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U339 (
    .O(n312),
    .I0(n106),
    .I1(key[75])
  );
  //AND U339bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U339bar (
    .O(n312bar),
    .I0(n106bar),
    .I1(keybar[75])
  );
  //AND U340
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U340 (
    .O(n311),
    .I0(key[75]),
    .I1(n106)
  );
  //OR U340bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U340bar (
    .O(n311bar),
    .I0(keybar[75]),
    .I1(n106bar)
  );
  //OR U341
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U341 (
    .O(out[74]),
    .I0(n313),
    .I1(n107)
  );
  //AND U341bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U341bar (
    .O(outbar[74]),
    .I0(n313bar),
    .I1(n107bar)
  );
  //OR U342
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U342 (
    .O(n314),
    .I0(n108),
    .I1(key[74])
  );
  //AND U342bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U342bar (
    .O(n314bar),
    .I0(n108bar),
    .I1(keybar[74])
  );
  //AND U343
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U343 (
    .O(n313),
    .I0(key[74]),
    .I1(n108)
  );
  //OR U343bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U343bar (
    .O(n313bar),
    .I0(keybar[74]),
    .I1(n108bar)
  );
  //OR U344
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U344 (
    .O(out[73]),
    .I0(n315),
    .I1(n109)
  );
  //AND U344bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U344bar (
    .O(outbar[73]),
    .I0(n315bar),
    .I1(n109bar)
  );
  //OR U345
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U345 (
    .O(n316),
    .I0(n110),
    .I1(key[73])
  );
  //AND U345bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U345bar (
    .O(n316bar),
    .I0(n110bar),
    .I1(keybar[73])
  );
  //AND U346
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U346 (
    .O(n315),
    .I0(key[73]),
    .I1(n110)
  );
  //OR U346bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U346bar (
    .O(n315bar),
    .I0(keybar[73]),
    .I1(n110bar)
  );
  //OR U347
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U347 (
    .O(out[72]),
    .I0(n317),
    .I1(n111)
  );
  //AND U347bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U347bar (
    .O(outbar[72]),
    .I0(n317bar),
    .I1(n111bar)
  );
  //OR U348
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U348 (
    .O(n318),
    .I0(n112),
    .I1(key[72])
  );
  //AND U348bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U348bar (
    .O(n318bar),
    .I0(n112bar),
    .I1(keybar[72])
  );
  //AND U349
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U349 (
    .O(n317),
    .I0(key[72]),
    .I1(n112)
  );
  //OR U349bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U349bar (
    .O(n317bar),
    .I0(keybar[72]),
    .I1(n112bar)
  );
  //OR U350
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U350 (
    .O(out[71]),
    .I0(n319),
    .I1(n113)
  );
  //AND U350bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U350bar (
    .O(outbar[71]),
    .I0(n319bar),
    .I1(n113bar)
  );
  //OR U351
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U351 (
    .O(n320),
    .I0(n114),
    .I1(key[71])
  );
  //AND U351bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U351bar (
    .O(n320bar),
    .I0(n114bar),
    .I1(keybar[71])
  );
  //AND U352
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U352 (
    .O(n319),
    .I0(key[71]),
    .I1(n114)
  );
  //OR U352bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U352bar (
    .O(n319bar),
    .I0(keybar[71]),
    .I1(n114bar)
  );
  //OR U353
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U353 (
    .O(out[70]),
    .I0(n321),
    .I1(n115)
  );
  //AND U353bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U353bar (
    .O(outbar[70]),
    .I0(n321bar),
    .I1(n115bar)
  );
  //OR U354
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U354 (
    .O(n322),
    .I0(n116),
    .I1(key[70])
  );
  //AND U354bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U354bar (
    .O(n322bar),
    .I0(n116bar),
    .I1(keybar[70])
  );
  //AND U355
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U355 (
    .O(n321),
    .I0(key[70]),
    .I1(n116)
  );
  //OR U355bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U355bar (
    .O(n321bar),
    .I0(keybar[70]),
    .I1(n116bar)
  );
  //OR U356
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U356 (
    .O(out[6]),
    .I0(n323),
    .I1(n243)
  );
  //AND U356bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U356bar (
    .O(outbar[6]),
    .I0(n323bar),
    .I1(n243bar)
  );
  //OR U357
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U357 (
    .O(n324),
    .I0(n244),
    .I1(key[6])
  );
  //AND U357bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U357bar (
    .O(n324bar),
    .I0(n244bar),
    .I1(keybar[6])
  );
  //AND U358
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U358 (
    .O(n323),
    .I0(key[6]),
    .I1(n244)
  );
  //OR U358bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U358bar (
    .O(n323bar),
    .I0(keybar[6]),
    .I1(n244bar)
  );
  //OR U359
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U359 (
    .O(out[69]),
    .I0(n325),
    .I1(n117)
  );
  //AND U359bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U359bar (
    .O(outbar[69]),
    .I0(n325bar),
    .I1(n117bar)
  );
  //OR U360
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U360 (
    .O(n326),
    .I0(n118),
    .I1(key[69])
  );
  //AND U360bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U360bar (
    .O(n326bar),
    .I0(n118bar),
    .I1(keybar[69])
  );
  //AND U361
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U361 (
    .O(n325),
    .I0(key[69]),
    .I1(n118)
  );
  //OR U361bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U361bar (
    .O(n325bar),
    .I0(keybar[69]),
    .I1(n118bar)
  );
  //OR U362
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U362 (
    .O(out[68]),
    .I0(n327),
    .I1(n119)
  );
  //AND U362bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U362bar (
    .O(outbar[68]),
    .I0(n327bar),
    .I1(n119bar)
  );
  //OR U363
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U363 (
    .O(n328),
    .I0(n120),
    .I1(key[68])
  );
  //AND U363bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U363bar (
    .O(n328bar),
    .I0(n120bar),
    .I1(keybar[68])
  );
  //AND U364
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U364 (
    .O(n327),
    .I0(key[68]),
    .I1(n120)
  );
  //OR U364bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U364bar (
    .O(n327bar),
    .I0(keybar[68]),
    .I1(n120bar)
  );
  //OR U365
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U365 (
    .O(out[67]),
    .I0(n329),
    .I1(n121)
  );
  //AND U365bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U365bar (
    .O(outbar[67]),
    .I0(n329bar),
    .I1(n121bar)
  );
  //OR U366
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U366 (
    .O(n330),
    .I0(n122),
    .I1(key[67])
  );
  //AND U366bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U366bar (
    .O(n330bar),
    .I0(n122bar),
    .I1(keybar[67])
  );
  //AND U367
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U367 (
    .O(n329),
    .I0(key[67]),
    .I1(n122)
  );
  //OR U367bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U367bar (
    .O(n329bar),
    .I0(keybar[67]),
    .I1(n122bar)
  );
  //OR U368
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U368 (
    .O(out[66]),
    .I0(n331),
    .I1(n123)
  );
  //AND U368bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U368bar (
    .O(outbar[66]),
    .I0(n331bar),
    .I1(n123bar)
  );
  //OR U369
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U369 (
    .O(n332),
    .I0(n124),
    .I1(key[66])
  );
  //AND U369bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U369bar (
    .O(n332bar),
    .I0(n124bar),
    .I1(keybar[66])
  );
  //AND U370
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U370 (
    .O(n331),
    .I0(key[66]),
    .I1(n124)
  );
  //OR U370bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U370bar (
    .O(n331bar),
    .I0(keybar[66]),
    .I1(n124bar)
  );
  //OR U371
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U371 (
    .O(out[65]),
    .I0(n333),
    .I1(n125)
  );
  //AND U371bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U371bar (
    .O(outbar[65]),
    .I0(n333bar),
    .I1(n125bar)
  );
  //OR U372
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U372 (
    .O(n334),
    .I0(n126),
    .I1(key[65])
  );
  //AND U372bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U372bar (
    .O(n334bar),
    .I0(n126bar),
    .I1(keybar[65])
  );
  //AND U373
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U373 (
    .O(n333),
    .I0(key[65]),
    .I1(n126)
  );
  //OR U373bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U373bar (
    .O(n333bar),
    .I0(keybar[65]),
    .I1(n126bar)
  );
  //OR U374
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U374 (
    .O(out[64]),
    .I0(n335),
    .I1(n127)
  );
  //AND U374bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U374bar (
    .O(outbar[64]),
    .I0(n335bar),
    .I1(n127bar)
  );
  //OR U375
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U375 (
    .O(n336),
    .I0(n128),
    .I1(key[64])
  );
  //AND U375bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U375bar (
    .O(n336bar),
    .I0(n128bar),
    .I1(keybar[64])
  );
  //AND U376
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U376 (
    .O(n335),
    .I0(key[64]),
    .I1(n128)
  );
  //OR U376bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U376bar (
    .O(n335bar),
    .I0(keybar[64]),
    .I1(n128bar)
  );
  //OR U377
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U377 (
    .O(out[63]),
    .I0(n337),
    .I1(n129)
  );
  //AND U377bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U377bar (
    .O(outbar[63]),
    .I0(n337bar),
    .I1(n129bar)
  );
  //OR U378
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U378 (
    .O(n338),
    .I0(n130),
    .I1(key[63])
  );
  //AND U378bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U378bar (
    .O(n338bar),
    .I0(n130bar),
    .I1(keybar[63])
  );
  //AND U379
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U379 (
    .O(n337),
    .I0(key[63]),
    .I1(n130)
  );
  //OR U379bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U379bar (
    .O(n337bar),
    .I0(keybar[63]),
    .I1(n130bar)
  );
  //OR U380
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U380 (
    .O(out[62]),
    .I0(n339),
    .I1(n131)
  );
  //AND U380bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U380bar (
    .O(outbar[62]),
    .I0(n339bar),
    .I1(n131bar)
  );
  //OR U381
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U381 (
    .O(n340),
    .I0(n132),
    .I1(key[62])
  );
  //AND U381bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U381bar (
    .O(n340bar),
    .I0(n132bar),
    .I1(keybar[62])
  );
  //AND U382
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U382 (
    .O(n339),
    .I0(key[62]),
    .I1(n132)
  );
  //OR U382bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U382bar (
    .O(n339bar),
    .I0(keybar[62]),
    .I1(n132bar)
  );
  //OR U383
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U383 (
    .O(out[61]),
    .I0(n341),
    .I1(n133)
  );
  //AND U383bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U383bar (
    .O(outbar[61]),
    .I0(n341bar),
    .I1(n133bar)
  );
  //OR U384
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U384 (
    .O(n342),
    .I0(n134),
    .I1(key[61])
  );
  //AND U384bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U384bar (
    .O(n342bar),
    .I0(n134bar),
    .I1(keybar[61])
  );
  //AND U385
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U385 (
    .O(n341),
    .I0(key[61]),
    .I1(n134)
  );
  //OR U385bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U385bar (
    .O(n341bar),
    .I0(keybar[61]),
    .I1(n134bar)
  );
  //OR U386
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U386 (
    .O(out[60]),
    .I0(n343),
    .I1(n135)
  );
  //AND U386bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U386bar (
    .O(outbar[60]),
    .I0(n343bar),
    .I1(n135bar)
  );
  //OR U387
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U387 (
    .O(n344),
    .I0(n136),
    .I1(key[60])
  );
  //AND U387bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U387bar (
    .O(n344bar),
    .I0(n136bar),
    .I1(keybar[60])
  );
  //AND U388
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U388 (
    .O(n343),
    .I0(key[60]),
    .I1(n136)
  );
  //OR U388bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U388bar (
    .O(n343bar),
    .I0(keybar[60]),
    .I1(n136bar)
  );
  //OR U389
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U389 (
    .O(out[5]),
    .I0(n345),
    .I1(n245)
  );
  //AND U389bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U389bar (
    .O(outbar[5]),
    .I0(n345bar),
    .I1(n245bar)
  );
  //OR U390
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U390 (
    .O(n346),
    .I0(n246),
    .I1(key[5])
  );
  //AND U390bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U390bar (
    .O(n346bar),
    .I0(n246bar),
    .I1(keybar[5])
  );
  //AND U391
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U391 (
    .O(n345),
    .I0(key[5]),
    .I1(n246)
  );
  //OR U391bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U391bar (
    .O(n345bar),
    .I0(keybar[5]),
    .I1(n246bar)
  );
  //OR U392
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U392 (
    .O(out[59]),
    .I0(n347),
    .I1(n137)
  );
  //AND U392bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U392bar (
    .O(outbar[59]),
    .I0(n347bar),
    .I1(n137bar)
  );
  //OR U393
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U393 (
    .O(n348),
    .I0(n138),
    .I1(key[59])
  );
  //AND U393bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U393bar (
    .O(n348bar),
    .I0(n138bar),
    .I1(keybar[59])
  );
  //AND U394
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U394 (
    .O(n347),
    .I0(key[59]),
    .I1(n138)
  );
  //OR U394bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U394bar (
    .O(n347bar),
    .I0(keybar[59]),
    .I1(n138bar)
  );
  //OR U395
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U395 (
    .O(out[58]),
    .I0(n349),
    .I1(n139)
  );
  //AND U395bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U395bar (
    .O(outbar[58]),
    .I0(n349bar),
    .I1(n139bar)
  );
  //OR U396
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U396 (
    .O(n350),
    .I0(n140),
    .I1(key[58])
  );
  //AND U396bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U396bar (
    .O(n350bar),
    .I0(n140bar),
    .I1(keybar[58])
  );
  //AND U397
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U397 (
    .O(n349),
    .I0(key[58]),
    .I1(n140)
  );
  //OR U397bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U397bar (
    .O(n349bar),
    .I0(keybar[58]),
    .I1(n140bar)
  );
  //OR U398
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U398 (
    .O(out[57]),
    .I0(n351),
    .I1(n141)
  );
  //AND U398bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U398bar (
    .O(outbar[57]),
    .I0(n351bar),
    .I1(n141bar)
  );
  //OR U399
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U399 (
    .O(n352),
    .I0(n142),
    .I1(key[57])
  );
  //AND U399bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U399bar (
    .O(n352bar),
    .I0(n142bar),
    .I1(keybar[57])
  );
  //AND U400
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U400 (
    .O(n351),
    .I0(key[57]),
    .I1(n142)
  );
  //OR U400bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U400bar (
    .O(n351bar),
    .I0(keybar[57]),
    .I1(n142bar)
  );
  //OR U401
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U401 (
    .O(out[56]),
    .I0(n353),
    .I1(n143)
  );
  //AND U401bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U401bar (
    .O(outbar[56]),
    .I0(n353bar),
    .I1(n143bar)
  );
  //OR U402
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U402 (
    .O(n354),
    .I0(n144),
    .I1(key[56])
  );
  //AND U402bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U402bar (
    .O(n354bar),
    .I0(n144bar),
    .I1(keybar[56])
  );
  //AND U403
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U403 (
    .O(n353),
    .I0(key[56]),
    .I1(n144)
  );
  //OR U403bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U403bar (
    .O(n353bar),
    .I0(keybar[56]),
    .I1(n144bar)
  );
  //OR U404
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U404 (
    .O(out[55]),
    .I0(n355),
    .I1(n145)
  );
  //AND U404bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U404bar (
    .O(outbar[55]),
    .I0(n355bar),
    .I1(n145bar)
  );
  //OR U405
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U405 (
    .O(n356),
    .I0(n146),
    .I1(key[55])
  );
  //AND U405bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U405bar (
    .O(n356bar),
    .I0(n146bar),
    .I1(keybar[55])
  );
  //AND U406
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U406 (
    .O(n355),
    .I0(key[55]),
    .I1(n146)
  );
  //OR U406bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U406bar (
    .O(n355bar),
    .I0(keybar[55]),
    .I1(n146bar)
  );
  //OR U407
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U407 (
    .O(out[54]),
    .I0(n357),
    .I1(n147)
  );
  //AND U407bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U407bar (
    .O(outbar[54]),
    .I0(n357bar),
    .I1(n147bar)
  );
  //OR U408
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U408 (
    .O(n358),
    .I0(n148),
    .I1(key[54])
  );
  //AND U408bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U408bar (
    .O(n358bar),
    .I0(n148bar),
    .I1(keybar[54])
  );
  //AND U409
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U409 (
    .O(n357),
    .I0(key[54]),
    .I1(n148)
  );
  //OR U409bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U409bar (
    .O(n357bar),
    .I0(keybar[54]),
    .I1(n148bar)
  );
  //OR U410
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U410 (
    .O(out[53]),
    .I0(n359),
    .I1(n149)
  );
  //AND U410bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U410bar (
    .O(outbar[53]),
    .I0(n359bar),
    .I1(n149bar)
  );
  //OR U411
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U411 (
    .O(n360),
    .I0(n150),
    .I1(key[53])
  );
  //AND U411bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U411bar (
    .O(n360bar),
    .I0(n150bar),
    .I1(keybar[53])
  );
  //AND U412
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U412 (
    .O(n359),
    .I0(key[53]),
    .I1(n150)
  );
  //OR U412bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U412bar (
    .O(n359bar),
    .I0(keybar[53]),
    .I1(n150bar)
  );
  //OR U413
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U413 (
    .O(out[52]),
    .I0(n361),
    .I1(n151)
  );
  //AND U413bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U413bar (
    .O(outbar[52]),
    .I0(n361bar),
    .I1(n151bar)
  );
  //OR U414
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U414 (
    .O(n362),
    .I0(n152),
    .I1(key[52])
  );
  //AND U414bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U414bar (
    .O(n362bar),
    .I0(n152bar),
    .I1(keybar[52])
  );
  //AND U415
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U415 (
    .O(n361),
    .I0(key[52]),
    .I1(n152)
  );
  //OR U415bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U415bar (
    .O(n361bar),
    .I0(keybar[52]),
    .I1(n152bar)
  );
  //OR U416
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U416 (
    .O(out[51]),
    .I0(n363),
    .I1(n153)
  );
  //AND U416bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U416bar (
    .O(outbar[51]),
    .I0(n363bar),
    .I1(n153bar)
  );
  //OR U417
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U417 (
    .O(n364),
    .I0(n154),
    .I1(key[51])
  );
  //AND U417bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U417bar (
    .O(n364bar),
    .I0(n154bar),
    .I1(keybar[51])
  );
  //AND U418
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U418 (
    .O(n363),
    .I0(key[51]),
    .I1(n154)
  );
  //OR U418bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U418bar (
    .O(n363bar),
    .I0(keybar[51]),
    .I1(n154bar)
  );
  //OR U419
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U419 (
    .O(out[50]),
    .I0(n365),
    .I1(n155)
  );
  //AND U419bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U419bar (
    .O(outbar[50]),
    .I0(n365bar),
    .I1(n155bar)
  );
  //OR U420
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U420 (
    .O(n366),
    .I0(n156),
    .I1(key[50])
  );
  //AND U420bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U420bar (
    .O(n366bar),
    .I0(n156bar),
    .I1(keybar[50])
  );
  //AND U421
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U421 (
    .O(n365),
    .I0(key[50]),
    .I1(n156)
  );
  //OR U421bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U421bar (
    .O(n365bar),
    .I0(keybar[50]),
    .I1(n156bar)
  );
  //OR U422
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U422 (
    .O(out[4]),
    .I0(n367),
    .I1(n247)
  );
  //AND U422bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U422bar (
    .O(outbar[4]),
    .I0(n367bar),
    .I1(n247bar)
  );
  //OR U423
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U423 (
    .O(n368),
    .I0(n248),
    .I1(key[4])
  );
  //AND U423bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U423bar (
    .O(n368bar),
    .I0(n248bar),
    .I1(keybar[4])
  );
  //AND U424
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U424 (
    .O(n367),
    .I0(key[4]),
    .I1(n248)
  );
  //OR U424bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U424bar (
    .O(n367bar),
    .I0(keybar[4]),
    .I1(n248bar)
  );
  //OR U425
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U425 (
    .O(out[49]),
    .I0(n369),
    .I1(n157)
  );
  //AND U425bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U425bar (
    .O(outbar[49]),
    .I0(n369bar),
    .I1(n157bar)
  );
  //OR U426
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U426 (
    .O(n370),
    .I0(n158),
    .I1(key[49])
  );
  //AND U426bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U426bar (
    .O(n370bar),
    .I0(n158bar),
    .I1(keybar[49])
  );
  //AND U427
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U427 (
    .O(n369),
    .I0(key[49]),
    .I1(n158)
  );
  //OR U427bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U427bar (
    .O(n369bar),
    .I0(keybar[49]),
    .I1(n158bar)
  );
  //OR U428
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U428 (
    .O(out[48]),
    .I0(n371),
    .I1(n159)
  );
  //AND U428bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U428bar (
    .O(outbar[48]),
    .I0(n371bar),
    .I1(n159bar)
  );
  //OR U429
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U429 (
    .O(n372),
    .I0(n160),
    .I1(key[48])
  );
  //AND U429bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U429bar (
    .O(n372bar),
    .I0(n160bar),
    .I1(keybar[48])
  );
  //AND U430
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U430 (
    .O(n371),
    .I0(key[48]),
    .I1(n160)
  );
  //OR U430bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U430bar (
    .O(n371bar),
    .I0(keybar[48]),
    .I1(n160bar)
  );
  //OR U431
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U431 (
    .O(out[47]),
    .I0(n373),
    .I1(n161)
  );
  //AND U431bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U431bar (
    .O(outbar[47]),
    .I0(n373bar),
    .I1(n161bar)
  );
  //OR U432
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U432 (
    .O(n374),
    .I0(n162),
    .I1(key[47])
  );
  //AND U432bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U432bar (
    .O(n374bar),
    .I0(n162bar),
    .I1(keybar[47])
  );
  //AND U433
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U433 (
    .O(n373),
    .I0(key[47]),
    .I1(n162)
  );
  //OR U433bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U433bar (
    .O(n373bar),
    .I0(keybar[47]),
    .I1(n162bar)
  );
  //OR U434
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U434 (
    .O(out[46]),
    .I0(n375),
    .I1(n163)
  );
  //AND U434bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U434bar (
    .O(outbar[46]),
    .I0(n375bar),
    .I1(n163bar)
  );
  //OR U435
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U435 (
    .O(n376),
    .I0(n164),
    .I1(key[46])
  );
  //AND U435bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U435bar (
    .O(n376bar),
    .I0(n164bar),
    .I1(keybar[46])
  );
  //AND U436
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U436 (
    .O(n375),
    .I0(key[46]),
    .I1(n164)
  );
  //OR U436bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U436bar (
    .O(n375bar),
    .I0(keybar[46]),
    .I1(n164bar)
  );
  //OR U437
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U437 (
    .O(out[45]),
    .I0(n377),
    .I1(n165)
  );
  //AND U437bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U437bar (
    .O(outbar[45]),
    .I0(n377bar),
    .I1(n165bar)
  );
  //OR U438
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U438 (
    .O(n378),
    .I0(n166),
    .I1(key[45])
  );
  //AND U438bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U438bar (
    .O(n378bar),
    .I0(n166bar),
    .I1(keybar[45])
  );
  //AND U439
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U439 (
    .O(n377),
    .I0(key[45]),
    .I1(n166)
  );
  //OR U439bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U439bar (
    .O(n377bar),
    .I0(keybar[45]),
    .I1(n166bar)
  );
  //OR U440
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U440 (
    .O(out[44]),
    .I0(n379),
    .I1(n167)
  );
  //AND U440bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U440bar (
    .O(outbar[44]),
    .I0(n379bar),
    .I1(n167bar)
  );
  //OR U441
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U441 (
    .O(n380),
    .I0(n168),
    .I1(key[44])
  );
  //AND U441bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U441bar (
    .O(n380bar),
    .I0(n168bar),
    .I1(keybar[44])
  );
  //AND U442
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U442 (
    .O(n379),
    .I0(key[44]),
    .I1(n168)
  );
  //OR U442bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U442bar (
    .O(n379bar),
    .I0(keybar[44]),
    .I1(n168bar)
  );
  //OR U443
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U443 (
    .O(out[43]),
    .I0(n381),
    .I1(n169)
  );
  //AND U443bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U443bar (
    .O(outbar[43]),
    .I0(n381bar),
    .I1(n169bar)
  );
  //OR U444
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U444 (
    .O(n382),
    .I0(n170),
    .I1(key[43])
  );
  //AND U444bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U444bar (
    .O(n382bar),
    .I0(n170bar),
    .I1(keybar[43])
  );
  //AND U445
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U445 (
    .O(n381),
    .I0(key[43]),
    .I1(n170)
  );
  //OR U445bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U445bar (
    .O(n381bar),
    .I0(keybar[43]),
    .I1(n170bar)
  );
  //OR U446
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U446 (
    .O(out[42]),
    .I0(n383),
    .I1(n171)
  );
  //AND U446bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U446bar (
    .O(outbar[42]),
    .I0(n383bar),
    .I1(n171bar)
  );
  //OR U447
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U447 (
    .O(n384),
    .I0(n172),
    .I1(key[42])
  );
  //AND U447bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U447bar (
    .O(n384bar),
    .I0(n172bar),
    .I1(keybar[42])
  );
  //AND U448
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U448 (
    .O(n383),
    .I0(key[42]),
    .I1(n172)
  );
  //OR U448bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U448bar (
    .O(n383bar),
    .I0(keybar[42]),
    .I1(n172bar)
  );
  //OR U449
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U449 (
    .O(out[41]),
    .I0(n385),
    .I1(n173)
  );
  //AND U449bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U449bar (
    .O(outbar[41]),
    .I0(n385bar),
    .I1(n173bar)
  );
  //OR U450
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U450 (
    .O(n386),
    .I0(n174),
    .I1(key[41])
  );
  //AND U450bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U450bar (
    .O(n386bar),
    .I0(n174bar),
    .I1(keybar[41])
  );
  //AND U451
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U451 (
    .O(n385),
    .I0(key[41]),
    .I1(n174)
  );
  //OR U451bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U451bar (
    .O(n385bar),
    .I0(keybar[41]),
    .I1(n174bar)
  );
  //OR U452
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U452 (
    .O(out[40]),
    .I0(n387),
    .I1(n175)
  );
  //AND U452bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U452bar (
    .O(outbar[40]),
    .I0(n387bar),
    .I1(n175bar)
  );
  //OR U453
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U453 (
    .O(n388),
    .I0(n176),
    .I1(key[40])
  );
  //AND U453bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U453bar (
    .O(n388bar),
    .I0(n176bar),
    .I1(keybar[40])
  );
  //AND U454
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U454 (
    .O(n387),
    .I0(key[40]),
    .I1(n176)
  );
  //OR U454bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U454bar (
    .O(n387bar),
    .I0(keybar[40]),
    .I1(n176bar)
  );
  //OR U455
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U455 (
    .O(out[3]),
    .I0(n389),
    .I1(n249)
  );
  //AND U455bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U455bar (
    .O(outbar[3]),
    .I0(n389bar),
    .I1(n249bar)
  );
  //OR U456
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U456 (
    .O(n390),
    .I0(n250),
    .I1(key[3])
  );
  //AND U456bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U456bar (
    .O(n390bar),
    .I0(n250bar),
    .I1(keybar[3])
  );
  //AND U457
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U457 (
    .O(n389),
    .I0(key[3]),
    .I1(n250)
  );
  //OR U457bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U457bar (
    .O(n389bar),
    .I0(keybar[3]),
    .I1(n250bar)
  );
  //OR U458
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U458 (
    .O(out[39]),
    .I0(n391),
    .I1(n177)
  );
  //AND U458bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U458bar (
    .O(outbar[39]),
    .I0(n391bar),
    .I1(n177bar)
  );
  //OR U459
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U459 (
    .O(n392),
    .I0(n178),
    .I1(key[39])
  );
  //AND U459bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U459bar (
    .O(n392bar),
    .I0(n178bar),
    .I1(keybar[39])
  );
  //AND U460
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U460 (
    .O(n391),
    .I0(key[39]),
    .I1(n178)
  );
  //OR U460bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U460bar (
    .O(n391bar),
    .I0(keybar[39]),
    .I1(n178bar)
  );
  //OR U461
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U461 (
    .O(out[38]),
    .I0(n393),
    .I1(n179)
  );
  //AND U461bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U461bar (
    .O(outbar[38]),
    .I0(n393bar),
    .I1(n179bar)
  );
  //OR U462
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U462 (
    .O(n394),
    .I0(n180),
    .I1(key[38])
  );
  //AND U462bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U462bar (
    .O(n394bar),
    .I0(n180bar),
    .I1(keybar[38])
  );
  //AND U463
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U463 (
    .O(n393),
    .I0(key[38]),
    .I1(n180)
  );
  //OR U463bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U463bar (
    .O(n393bar),
    .I0(keybar[38]),
    .I1(n180bar)
  );
  //OR U464
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U464 (
    .O(out[37]),
    .I0(n395),
    .I1(n181)
  );
  //AND U464bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U464bar (
    .O(outbar[37]),
    .I0(n395bar),
    .I1(n181bar)
  );
  //OR U465
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U465 (
    .O(n396),
    .I0(n182),
    .I1(key[37])
  );
  //AND U465bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U465bar (
    .O(n396bar),
    .I0(n182bar),
    .I1(keybar[37])
  );
  //AND U466
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U466 (
    .O(n395),
    .I0(key[37]),
    .I1(n182)
  );
  //OR U466bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U466bar (
    .O(n395bar),
    .I0(keybar[37]),
    .I1(n182bar)
  );
  //OR U467
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U467 (
    .O(out[36]),
    .I0(n397),
    .I1(n183)
  );
  //AND U467bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U467bar (
    .O(outbar[36]),
    .I0(n397bar),
    .I1(n183bar)
  );
  //OR U468
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U468 (
    .O(n398),
    .I0(n184),
    .I1(key[36])
  );
  //AND U468bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U468bar (
    .O(n398bar),
    .I0(n184bar),
    .I1(keybar[36])
  );
  //AND U469
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U469 (
    .O(n397),
    .I0(key[36]),
    .I1(n184)
  );
  //OR U469bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U469bar (
    .O(n397bar),
    .I0(keybar[36]),
    .I1(n184bar)
  );
  //OR U470
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U470 (
    .O(out[35]),
    .I0(n399),
    .I1(n185)
  );
  //AND U470bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U470bar (
    .O(outbar[35]),
    .I0(n399bar),
    .I1(n185bar)
  );
  //OR U471
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U471 (
    .O(n400),
    .I0(n186),
    .I1(key[35])
  );
  //AND U471bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U471bar (
    .O(n400bar),
    .I0(n186bar),
    .I1(keybar[35])
  );
  //AND U472
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U472 (
    .O(n399),
    .I0(key[35]),
    .I1(n186)
  );
  //OR U472bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U472bar (
    .O(n399bar),
    .I0(keybar[35]),
    .I1(n186bar)
  );
  //OR U473
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U473 (
    .O(out[34]),
    .I0(n401),
    .I1(n187)
  );
  //AND U473bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U473bar (
    .O(outbar[34]),
    .I0(n401bar),
    .I1(n187bar)
  );
  //OR U474
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U474 (
    .O(n402),
    .I0(n188),
    .I1(key[34])
  );
  //AND U474bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U474bar (
    .O(n402bar),
    .I0(n188bar),
    .I1(keybar[34])
  );
  //AND U475
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U475 (
    .O(n401),
    .I0(key[34]),
    .I1(n188)
  );
  //OR U475bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U475bar (
    .O(n401bar),
    .I0(keybar[34]),
    .I1(n188bar)
  );
  //OR U476
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U476 (
    .O(out[33]),
    .I0(n403),
    .I1(n189)
  );
  //AND U476bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U476bar (
    .O(outbar[33]),
    .I0(n403bar),
    .I1(n189bar)
  );
  //OR U477
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U477 (
    .O(n404),
    .I0(n190),
    .I1(key[33])
  );
  //AND U477bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U477bar (
    .O(n404bar),
    .I0(n190bar),
    .I1(keybar[33])
  );
  //AND U478
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U478 (
    .O(n403),
    .I0(key[33]),
    .I1(n190)
  );
  //OR U478bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U478bar (
    .O(n403bar),
    .I0(keybar[33]),
    .I1(n190bar)
  );
  //OR U479
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U479 (
    .O(out[32]),
    .I0(n405),
    .I1(n191)
  );
  //AND U479bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U479bar (
    .O(outbar[32]),
    .I0(n405bar),
    .I1(n191bar)
  );
  //OR U480
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U480 (
    .O(n406),
    .I0(n192),
    .I1(key[32])
  );
  //AND U480bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U480bar (
    .O(n406bar),
    .I0(n192bar),
    .I1(keybar[32])
  );
  //AND U481
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U481 (
    .O(n405),
    .I0(key[32]),
    .I1(n192)
  );
  //OR U481bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U481bar (
    .O(n405bar),
    .I0(keybar[32]),
    .I1(n192bar)
  );
  //OR U482
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U482 (
    .O(out[31]),
    .I0(n407),
    .I1(n193)
  );
  //AND U482bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U482bar (
    .O(outbar[31]),
    .I0(n407bar),
    .I1(n193bar)
  );
  //OR U483
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U483 (
    .O(n408),
    .I0(n194),
    .I1(key[31])
  );
  //AND U483bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U483bar (
    .O(n408bar),
    .I0(n194bar),
    .I1(keybar[31])
  );
  //AND U484
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U484 (
    .O(n407),
    .I0(key[31]),
    .I1(n194)
  );
  //OR U484bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U484bar (
    .O(n407bar),
    .I0(keybar[31]),
    .I1(n194bar)
  );
  //OR U485
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U485 (
    .O(out[30]),
    .I0(n409),
    .I1(n195)
  );
  //AND U485bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U485bar (
    .O(outbar[30]),
    .I0(n409bar),
    .I1(n195bar)
  );
  //OR U486
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U486 (
    .O(n410),
    .I0(n196),
    .I1(key[30])
  );
  //AND U486bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U486bar (
    .O(n410bar),
    .I0(n196bar),
    .I1(keybar[30])
  );
  //AND U487
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U487 (
    .O(n409),
    .I0(key[30]),
    .I1(n196)
  );
  //OR U487bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U487bar (
    .O(n409bar),
    .I0(keybar[30]),
    .I1(n196bar)
  );
  //OR U488
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U488 (
    .O(out[2]),
    .I0(n411),
    .I1(n251)
  );
  //AND U488bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U488bar (
    .O(outbar[2]),
    .I0(n411bar),
    .I1(n251bar)
  );
  //OR U489
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U489 (
    .O(n412),
    .I0(n252),
    .I1(key[2])
  );
  //AND U489bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U489bar (
    .O(n412bar),
    .I0(n252bar),
    .I1(keybar[2])
  );
  //AND U490
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U490 (
    .O(n411),
    .I0(key[2]),
    .I1(n252)
  );
  //OR U490bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U490bar (
    .O(n411bar),
    .I0(keybar[2]),
    .I1(n252bar)
  );
  //OR U491
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U491 (
    .O(out[29]),
    .I0(n413),
    .I1(n197)
  );
  //AND U491bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U491bar (
    .O(outbar[29]),
    .I0(n413bar),
    .I1(n197bar)
  );
  //OR U492
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U492 (
    .O(n414),
    .I0(n198),
    .I1(key[29])
  );
  //AND U492bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U492bar (
    .O(n414bar),
    .I0(n198bar),
    .I1(keybar[29])
  );
  //AND U493
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U493 (
    .O(n413),
    .I0(key[29]),
    .I1(n198)
  );
  //OR U493bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U493bar (
    .O(n413bar),
    .I0(keybar[29]),
    .I1(n198bar)
  );
  //OR U494
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U494 (
    .O(out[28]),
    .I0(n415),
    .I1(n199)
  );
  //AND U494bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U494bar (
    .O(outbar[28]),
    .I0(n415bar),
    .I1(n199bar)
  );
  //OR U495
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U495 (
    .O(n416),
    .I0(n200),
    .I1(key[28])
  );
  //AND U495bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U495bar (
    .O(n416bar),
    .I0(n200bar),
    .I1(keybar[28])
  );
  //AND U496
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U496 (
    .O(n415),
    .I0(key[28]),
    .I1(n200)
  );
  //OR U496bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U496bar (
    .O(n415bar),
    .I0(keybar[28]),
    .I1(n200bar)
  );
  //OR U497
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U497 (
    .O(out[27]),
    .I0(n417),
    .I1(n201)
  );
  //AND U497bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U497bar (
    .O(outbar[27]),
    .I0(n417bar),
    .I1(n201bar)
  );
  //OR U498
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U498 (
    .O(n418),
    .I0(n202),
    .I1(key[27])
  );
  //AND U498bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U498bar (
    .O(n418bar),
    .I0(n202bar),
    .I1(keybar[27])
  );
  //AND U499
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U499 (
    .O(n417),
    .I0(key[27]),
    .I1(n202)
  );
  //OR U499bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U499bar (
    .O(n417bar),
    .I0(keybar[27]),
    .I1(n202bar)
  );
  //OR U500
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U500 (
    .O(out[26]),
    .I0(n419),
    .I1(n203)
  );
  //AND U500bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U500bar (
    .O(outbar[26]),
    .I0(n419bar),
    .I1(n203bar)
  );
  //OR U501
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U501 (
    .O(n420),
    .I0(n204),
    .I1(key[26])
  );
  //AND U501bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U501bar (
    .O(n420bar),
    .I0(n204bar),
    .I1(keybar[26])
  );
  //AND U502
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U502 (
    .O(n419),
    .I0(key[26]),
    .I1(n204)
  );
  //OR U502bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U502bar (
    .O(n419bar),
    .I0(keybar[26]),
    .I1(n204bar)
  );
  //OR U503
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U503 (
    .O(out[25]),
    .I0(n421),
    .I1(n205)
  );
  //AND U503bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U503bar (
    .O(outbar[25]),
    .I0(n421bar),
    .I1(n205bar)
  );
  //OR U504
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U504 (
    .O(n422),
    .I0(n206),
    .I1(key[25])
  );
  //AND U504bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U504bar (
    .O(n422bar),
    .I0(n206bar),
    .I1(keybar[25])
  );
  //AND U505
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U505 (
    .O(n421),
    .I0(key[25]),
    .I1(n206)
  );
  //OR U505bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U505bar (
    .O(n421bar),
    .I0(keybar[25]),
    .I1(n206bar)
  );
  //OR U506
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U506 (
    .O(out[24]),
    .I0(n423),
    .I1(n207)
  );
  //AND U506bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U506bar (
    .O(outbar[24]),
    .I0(n423bar),
    .I1(n207bar)
  );
  //OR U507
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U507 (
    .O(n424),
    .I0(n208),
    .I1(key[24])
  );
  //AND U507bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U507bar (
    .O(n424bar),
    .I0(n208bar),
    .I1(keybar[24])
  );
  //AND U508
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U508 (
    .O(n423),
    .I0(key[24]),
    .I1(n208)
  );
  //OR U508bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U508bar (
    .O(n423bar),
    .I0(keybar[24]),
    .I1(n208bar)
  );
  //OR U509
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U509 (
    .O(out[23]),
    .I0(n425),
    .I1(n209)
  );
  //AND U509bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U509bar (
    .O(outbar[23]),
    .I0(n425bar),
    .I1(n209bar)
  );
  //OR U510
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U510 (
    .O(n426),
    .I0(n210),
    .I1(key[23])
  );
  //AND U510bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U510bar (
    .O(n426bar),
    .I0(n210bar),
    .I1(keybar[23])
  );
  //AND U511
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U511 (
    .O(n425),
    .I0(key[23]),
    .I1(n210)
  );
  //OR U511bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U511bar (
    .O(n425bar),
    .I0(keybar[23]),
    .I1(n210bar)
  );
  //OR U512
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U512 (
    .O(out[22]),
    .I0(n427),
    .I1(n211)
  );
  //AND U512bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U512bar (
    .O(outbar[22]),
    .I0(n427bar),
    .I1(n211bar)
  );
  //OR U513
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U513 (
    .O(n428),
    .I0(n212),
    .I1(key[22])
  );
  //AND U513bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U513bar (
    .O(n428bar),
    .I0(n212bar),
    .I1(keybar[22])
  );
  //AND U514
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U514 (
    .O(n427),
    .I0(key[22]),
    .I1(n212)
  );
  //OR U514bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U514bar (
    .O(n427bar),
    .I0(keybar[22]),
    .I1(n212bar)
  );
  //OR U515
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U515 (
    .O(out[21]),
    .I0(n429),
    .I1(n213)
  );
  //AND U515bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U515bar (
    .O(outbar[21]),
    .I0(n429bar),
    .I1(n213bar)
  );
  //OR U516
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U516 (
    .O(n430),
    .I0(n214),
    .I1(key[21])
  );
  //AND U516bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U516bar (
    .O(n430bar),
    .I0(n214bar),
    .I1(keybar[21])
  );
  //AND U517
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U517 (
    .O(n429),
    .I0(key[21]),
    .I1(n214)
  );
  //OR U517bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U517bar (
    .O(n429bar),
    .I0(keybar[21]),
    .I1(n214bar)
  );
  //OR U518
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U518 (
    .O(out[20]),
    .I0(n431),
    .I1(n215)
  );
  //AND U518bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U518bar (
    .O(outbar[20]),
    .I0(n431bar),
    .I1(n215bar)
  );
  //OR U519
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U519 (
    .O(n432),
    .I0(n216),
    .I1(key[20])
  );
  //AND U519bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U519bar (
    .O(n432bar),
    .I0(n216bar),
    .I1(keybar[20])
  );
  //AND U520
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U520 (
    .O(n431),
    .I0(key[20]),
    .I1(n216)
  );
  //OR U520bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U520bar (
    .O(n431bar),
    .I0(keybar[20]),
    .I1(n216bar)
  );
  //OR U521
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U521 (
    .O(out[1]),
    .I0(n433),
    .I1(n253)
  );
  //AND U521bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U521bar (
    .O(outbar[1]),
    .I0(n433bar),
    .I1(n253bar)
  );
  //OR U522
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U522 (
    .O(n434),
    .I0(n254),
    .I1(key[1])
  );
  //AND U522bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U522bar (
    .O(n434bar),
    .I0(n254bar),
    .I1(keybar[1])
  );
  //AND U523
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U523 (
    .O(n433),
    .I0(key[1]),
    .I1(n254)
  );
  //OR U523bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U523bar (
    .O(n433bar),
    .I0(keybar[1]),
    .I1(n254bar)
  );
  //OR U524
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U524 (
    .O(out[19]),
    .I0(n435),
    .I1(n217)
  );
  //AND U524bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U524bar (
    .O(outbar[19]),
    .I0(n435bar),
    .I1(n217bar)
  );
  //OR U525
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U525 (
    .O(n436),
    .I0(n218),
    .I1(key[19])
  );
  //AND U525bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U525bar (
    .O(n436bar),
    .I0(n218bar),
    .I1(keybar[19])
  );
  //AND U526
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U526 (
    .O(n435),
    .I0(key[19]),
    .I1(n218)
  );
  //OR U526bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U526bar (
    .O(n435bar),
    .I0(keybar[19]),
    .I1(n218bar)
  );
  //OR U527
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U527 (
    .O(out[18]),
    .I0(n437),
    .I1(n219)
  );
  //AND U527bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U527bar (
    .O(outbar[18]),
    .I0(n437bar),
    .I1(n219bar)
  );
  //OR U528
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U528 (
    .O(n438),
    .I0(n220),
    .I1(key[18])
  );
  //AND U528bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U528bar (
    .O(n438bar),
    .I0(n220bar),
    .I1(keybar[18])
  );
  //AND U529
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U529 (
    .O(n437),
    .I0(key[18]),
    .I1(n220)
  );
  //OR U529bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U529bar (
    .O(n437bar),
    .I0(keybar[18]),
    .I1(n220bar)
  );
  //OR U530
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U530 (
    .O(out[17]),
    .I0(n439),
    .I1(n221)
  );
  //AND U530bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U530bar (
    .O(outbar[17]),
    .I0(n439bar),
    .I1(n221bar)
  );
  //OR U531
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U531 (
    .O(n440),
    .I0(n222),
    .I1(key[17])
  );
  //AND U531bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U531bar (
    .O(n440bar),
    .I0(n222bar),
    .I1(keybar[17])
  );
  //AND U532
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U532 (
    .O(n439),
    .I0(key[17]),
    .I1(n222)
  );
  //OR U532bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U532bar (
    .O(n439bar),
    .I0(keybar[17]),
    .I1(n222bar)
  );
  //OR U533
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U533 (
    .O(out[16]),
    .I0(n441),
    .I1(n223)
  );
  //AND U533bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U533bar (
    .O(outbar[16]),
    .I0(n441bar),
    .I1(n223bar)
  );
  //OR U534
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U534 (
    .O(n442),
    .I0(n224),
    .I1(key[16])
  );
  //AND U534bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U534bar (
    .O(n442bar),
    .I0(n224bar),
    .I1(keybar[16])
  );
  //AND U535
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U535 (
    .O(n441),
    .I0(key[16]),
    .I1(n224)
  );
  //OR U535bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U535bar (
    .O(n441bar),
    .I0(keybar[16]),
    .I1(n224bar)
  );
  //OR U536
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U536 (
    .O(out[15]),
    .I0(n443),
    .I1(n225)
  );
  //AND U536bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U536bar (
    .O(outbar[15]),
    .I0(n443bar),
    .I1(n225bar)
  );
  //OR U537
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U537 (
    .O(n444),
    .I0(n226),
    .I1(key[15])
  );
  //AND U537bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U537bar (
    .O(n444bar),
    .I0(n226bar),
    .I1(keybar[15])
  );
  //AND U538
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U538 (
    .O(n443),
    .I0(key[15]),
    .I1(n226)
  );
  //OR U538bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U538bar (
    .O(n443bar),
    .I0(keybar[15]),
    .I1(n226bar)
  );
  //OR U539
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U539 (
    .O(out[14]),
    .I0(n445),
    .I1(n227)
  );
  //AND U539bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U539bar (
    .O(outbar[14]),
    .I0(n445bar),
    .I1(n227bar)
  );
  //OR U540
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U540 (
    .O(n446),
    .I0(n228),
    .I1(key[14])
  );
  //AND U540bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U540bar (
    .O(n446bar),
    .I0(n228bar),
    .I1(keybar[14])
  );
  //AND U541
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U541 (
    .O(n445),
    .I0(key[14]),
    .I1(n228)
  );
  //OR U541bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U541bar (
    .O(n445bar),
    .I0(keybar[14]),
    .I1(n228bar)
  );
  //OR U542
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U542 (
    .O(out[13]),
    .I0(n447),
    .I1(n229)
  );
  //AND U542bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U542bar (
    .O(outbar[13]),
    .I0(n447bar),
    .I1(n229bar)
  );
  //OR U543
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U543 (
    .O(n448),
    .I0(n230),
    .I1(key[13])
  );
  //AND U543bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U543bar (
    .O(n448bar),
    .I0(n230bar),
    .I1(keybar[13])
  );
  //AND U544
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U544 (
    .O(n447),
    .I0(key[13]),
    .I1(n230)
  );
  //OR U544bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U544bar (
    .O(n447bar),
    .I0(keybar[13]),
    .I1(n230bar)
  );
  //OR U545
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U545 (
    .O(out[12]),
    .I0(n449),
    .I1(n231)
  );
  //AND U545bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U545bar (
    .O(outbar[12]),
    .I0(n449bar),
    .I1(n231bar)
  );
  //OR U546
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U546 (
    .O(n450),
    .I0(n232),
    .I1(key[12])
  );
  //AND U546bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U546bar (
    .O(n450bar),
    .I0(n232bar),
    .I1(keybar[12])
  );
  //AND U547
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U547 (
    .O(n449),
    .I0(key[12]),
    .I1(n232)
  );
  //OR U547bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U547bar (
    .O(n449bar),
    .I0(keybar[12]),
    .I1(n232bar)
  );
  //OR U548
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U548 (
    .O(out[127]),
    .I0(n451),
    .I1(n1)
  );
  //AND U548bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U548bar (
    .O(outbar[127]),
    .I0(n451bar),
    .I1(n1bar)
  );
  //OR U549
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U549 (
    .O(n452),
    .I0(n2),
    .I1(key[127])
  );
  //AND U549bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U549bar (
    .O(n452bar),
    .I0(n2bar),
    .I1(keybar[127])
  );
  //AND U550
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U550 (
    .O(n451),
    .I0(key[127]),
    .I1(n2)
  );
  //OR U550bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U550bar (
    .O(n451bar),
    .I0(keybar[127]),
    .I1(n2bar)
  );
  //OR U551
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U551 (
    .O(out[126]),
    .I0(n453),
    .I1(n3)
  );
  //AND U551bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U551bar (
    .O(outbar[126]),
    .I0(n453bar),
    .I1(n3bar)
  );
  //OR U552
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U552 (
    .O(n454),
    .I0(n4),
    .I1(key[126])
  );
  //AND U552bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U552bar (
    .O(n454bar),
    .I0(n4bar),
    .I1(keybar[126])
  );
  //AND U553
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U553 (
    .O(n453),
    .I0(key[126]),
    .I1(n4)
  );
  //OR U553bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U553bar (
    .O(n453bar),
    .I0(keybar[126]),
    .I1(n4bar)
  );
  //OR U554
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U554 (
    .O(out[125]),
    .I0(n455),
    .I1(n5)
  );
  //AND U554bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U554bar (
    .O(outbar[125]),
    .I0(n455bar),
    .I1(n5bar)
  );
  //OR U555
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U555 (
    .O(n456),
    .I0(n6),
    .I1(key[125])
  );
  //AND U555bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U555bar (
    .O(n456bar),
    .I0(n6bar),
    .I1(keybar[125])
  );
  //AND U556
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U556 (
    .O(n455),
    .I0(key[125]),
    .I1(n6)
  );
  //OR U556bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U556bar (
    .O(n455bar),
    .I0(keybar[125]),
    .I1(n6bar)
  );
  //OR U557
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U557 (
    .O(out[124]),
    .I0(n457),
    .I1(n7)
  );
  //AND U557bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U557bar (
    .O(outbar[124]),
    .I0(n457bar),
    .I1(n7bar)
  );
  //OR U558
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U558 (
    .O(n458),
    .I0(n8),
    .I1(key[124])
  );
  //AND U558bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U558bar (
    .O(n458bar),
    .I0(n8bar),
    .I1(keybar[124])
  );
  //AND U559
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U559 (
    .O(n457),
    .I0(key[124]),
    .I1(n8)
  );
  //OR U559bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U559bar (
    .O(n457bar),
    .I0(keybar[124]),
    .I1(n8bar)
  );
  //OR U560
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U560 (
    .O(out[123]),
    .I0(n459),
    .I1(n9)
  );
  //AND U560bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U560bar (
    .O(outbar[123]),
    .I0(n459bar),
    .I1(n9bar)
  );
  //OR U561
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U561 (
    .O(n460),
    .I0(n10),
    .I1(key[123])
  );
  //AND U561bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U561bar (
    .O(n460bar),
    .I0(n10bar),
    .I1(keybar[123])
  );
  //AND U562
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U562 (
    .O(n459),
    .I0(key[123]),
    .I1(n10)
  );
  //OR U562bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U562bar (
    .O(n459bar),
    .I0(keybar[123]),
    .I1(n10bar)
  );
  //OR U563
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U563 (
    .O(out[122]),
    .I0(n461),
    .I1(n11)
  );
  //AND U563bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U563bar (
    .O(outbar[122]),
    .I0(n461bar),
    .I1(n11bar)
  );
  //OR U564
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U564 (
    .O(n462),
    .I0(n12),
    .I1(key[122])
  );
  //AND U564bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U564bar (
    .O(n462bar),
    .I0(n12bar),
    .I1(keybar[122])
  );
  //AND U565
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U565 (
    .O(n461),
    .I0(key[122]),
    .I1(n12)
  );
  //OR U565bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U565bar (
    .O(n461bar),
    .I0(keybar[122]),
    .I1(n12bar)
  );
  //OR U566
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U566 (
    .O(out[121]),
    .I0(n463),
    .I1(n13)
  );
  //AND U566bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U566bar (
    .O(outbar[121]),
    .I0(n463bar),
    .I1(n13bar)
  );
  //OR U567
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U567 (
    .O(n464),
    .I0(n14),
    .I1(key[121])
  );
  //AND U567bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U567bar (
    .O(n464bar),
    .I0(n14bar),
    .I1(keybar[121])
  );
  //AND U568
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U568 (
    .O(n463),
    .I0(key[121]),
    .I1(n14)
  );
  //OR U568bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U568bar (
    .O(n463bar),
    .I0(keybar[121]),
    .I1(n14bar)
  );
  //OR U569
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U569 (
    .O(out[120]),
    .I0(n465),
    .I1(n15)
  );
  //AND U569bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U569bar (
    .O(outbar[120]),
    .I0(n465bar),
    .I1(n15bar)
  );
  //OR U570
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U570 (
    .O(n466),
    .I0(n16),
    .I1(key[120])
  );
  //AND U570bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U570bar (
    .O(n466bar),
    .I0(n16bar),
    .I1(keybar[120])
  );
  //AND U571
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U571 (
    .O(n465),
    .I0(key[120]),
    .I1(n16)
  );
  //OR U571bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U571bar (
    .O(n465bar),
    .I0(keybar[120]),
    .I1(n16bar)
  );
  //OR U572
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U572 (
    .O(out[11]),
    .I0(n467),
    .I1(n233)
  );
  //AND U572bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U572bar (
    .O(outbar[11]),
    .I0(n467bar),
    .I1(n233bar)
  );
  //OR U573
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U573 (
    .O(n468),
    .I0(n234),
    .I1(key[11])
  );
  //AND U573bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U573bar (
    .O(n468bar),
    .I0(n234bar),
    .I1(keybar[11])
  );
  //AND U574
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U574 (
    .O(n467),
    .I0(key[11]),
    .I1(n234)
  );
  //OR U574bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U574bar (
    .O(n467bar),
    .I0(keybar[11]),
    .I1(n234bar)
  );
  //OR U575
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U575 (
    .O(out[119]),
    .I0(n469),
    .I1(n17)
  );
  //AND U575bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U575bar (
    .O(outbar[119]),
    .I0(n469bar),
    .I1(n17bar)
  );
  //OR U576
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U576 (
    .O(n470),
    .I0(n18),
    .I1(key[119])
  );
  //AND U576bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U576bar (
    .O(n470bar),
    .I0(n18bar),
    .I1(keybar[119])
  );
  //AND U577
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U577 (
    .O(n469),
    .I0(key[119]),
    .I1(n18)
  );
  //OR U577bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U577bar (
    .O(n469bar),
    .I0(keybar[119]),
    .I1(n18bar)
  );
  //OR U578
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U578 (
    .O(out[118]),
    .I0(n471),
    .I1(n19)
  );
  //AND U578bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U578bar (
    .O(outbar[118]),
    .I0(n471bar),
    .I1(n19bar)
  );
  //OR U579
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U579 (
    .O(n472),
    .I0(n20),
    .I1(key[118])
  );
  //AND U579bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U579bar (
    .O(n472bar),
    .I0(n20bar),
    .I1(keybar[118])
  );
  //AND U580
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U580 (
    .O(n471),
    .I0(key[118]),
    .I1(n20)
  );
  //OR U580bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U580bar (
    .O(n471bar),
    .I0(keybar[118]),
    .I1(n20bar)
  );
  //OR U581
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U581 (
    .O(out[117]),
    .I0(n473),
    .I1(n21)
  );
  //AND U581bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U581bar (
    .O(outbar[117]),
    .I0(n473bar),
    .I1(n21bar)
  );
  //OR U582
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U582 (
    .O(n474),
    .I0(n22),
    .I1(key[117])
  );
  //AND U582bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U582bar (
    .O(n474bar),
    .I0(n22bar),
    .I1(keybar[117])
  );
  //AND U583
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U583 (
    .O(n473),
    .I0(key[117]),
    .I1(n22)
  );
  //OR U583bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U583bar (
    .O(n473bar),
    .I0(keybar[117]),
    .I1(n22bar)
  );
  //OR U584
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U584 (
    .O(out[116]),
    .I0(n475),
    .I1(n23)
  );
  //AND U584bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U584bar (
    .O(outbar[116]),
    .I0(n475bar),
    .I1(n23bar)
  );
  //OR U585
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U585 (
    .O(n476),
    .I0(n24),
    .I1(key[116])
  );
  //AND U585bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U585bar (
    .O(n476bar),
    .I0(n24bar),
    .I1(keybar[116])
  );
  //AND U586
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U586 (
    .O(n475),
    .I0(key[116]),
    .I1(n24)
  );
  //OR U586bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U586bar (
    .O(n475bar),
    .I0(keybar[116]),
    .I1(n24bar)
  );
  //OR U587
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U587 (
    .O(out[115]),
    .I0(n477),
    .I1(n25)
  );
  //AND U587bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U587bar (
    .O(outbar[115]),
    .I0(n477bar),
    .I1(n25bar)
  );
  //OR U588
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U588 (
    .O(n478),
    .I0(n26),
    .I1(key[115])
  );
  //AND U588bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U588bar (
    .O(n478bar),
    .I0(n26bar),
    .I1(keybar[115])
  );
  //AND U589
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U589 (
    .O(n477),
    .I0(key[115]),
    .I1(n26)
  );
  //OR U589bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U589bar (
    .O(n477bar),
    .I0(keybar[115]),
    .I1(n26bar)
  );
  //OR U590
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U590 (
    .O(out[114]),
    .I0(n479),
    .I1(n27)
  );
  //AND U590bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U590bar (
    .O(outbar[114]),
    .I0(n479bar),
    .I1(n27bar)
  );
  //OR U591
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U591 (
    .O(n480),
    .I0(n28),
    .I1(key[114])
  );
  //AND U591bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U591bar (
    .O(n480bar),
    .I0(n28bar),
    .I1(keybar[114])
  );
  //AND U592
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U592 (
    .O(n479),
    .I0(key[114]),
    .I1(n28)
  );
  //OR U592bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U592bar (
    .O(n479bar),
    .I0(keybar[114]),
    .I1(n28bar)
  );
  //OR U593
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U593 (
    .O(out[113]),
    .I0(n481),
    .I1(n29)
  );
  //AND U593bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U593bar (
    .O(outbar[113]),
    .I0(n481bar),
    .I1(n29bar)
  );
  //OR U594
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U594 (
    .O(n482),
    .I0(n30),
    .I1(key[113])
  );
  //AND U594bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U594bar (
    .O(n482bar),
    .I0(n30bar),
    .I1(keybar[113])
  );
  //AND U595
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U595 (
    .O(n481),
    .I0(key[113]),
    .I1(n30)
  );
  //OR U595bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U595bar (
    .O(n481bar),
    .I0(keybar[113]),
    .I1(n30bar)
  );
  //OR U596
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U596 (
    .O(out[112]),
    .I0(n483),
    .I1(n31)
  );
  //AND U596bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U596bar (
    .O(outbar[112]),
    .I0(n483bar),
    .I1(n31bar)
  );
  //OR U597
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U597 (
    .O(n484),
    .I0(n32),
    .I1(key[112])
  );
  //AND U597bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U597bar (
    .O(n484bar),
    .I0(n32bar),
    .I1(keybar[112])
  );
  //AND U598
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U598 (
    .O(n483),
    .I0(key[112]),
    .I1(n32)
  );
  //OR U598bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U598bar (
    .O(n483bar),
    .I0(keybar[112]),
    .I1(n32bar)
  );
  //OR U599
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U599 (
    .O(out[111]),
    .I0(n485),
    .I1(n33)
  );
  //AND U599bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U599bar (
    .O(outbar[111]),
    .I0(n485bar),
    .I1(n33bar)
  );
  //OR U600
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U600 (
    .O(n486),
    .I0(n34),
    .I1(key[111])
  );
  //AND U600bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U600bar (
    .O(n486bar),
    .I0(n34bar),
    .I1(keybar[111])
  );
  //AND U601
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U601 (
    .O(n485),
    .I0(key[111]),
    .I1(n34)
  );
  //OR U601bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U601bar (
    .O(n485bar),
    .I0(keybar[111]),
    .I1(n34bar)
  );
  //OR U602
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U602 (
    .O(out[110]),
    .I0(n487),
    .I1(n35)
  );
  //AND U602bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U602bar (
    .O(outbar[110]),
    .I0(n487bar),
    .I1(n35bar)
  );
  //OR U603
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U603 (
    .O(n488),
    .I0(n36),
    .I1(key[110])
  );
  //AND U603bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U603bar (
    .O(n488bar),
    .I0(n36bar),
    .I1(keybar[110])
  );
  //AND U604
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U604 (
    .O(n487),
    .I0(key[110]),
    .I1(n36)
  );
  //OR U604bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U604bar (
    .O(n487bar),
    .I0(keybar[110]),
    .I1(n36bar)
  );
  //OR U605
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U605 (
    .O(out[10]),
    .I0(n489),
    .I1(n235)
  );
  //AND U605bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U605bar (
    .O(outbar[10]),
    .I0(n489bar),
    .I1(n235bar)
  );
  //OR U606
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U606 (
    .O(n490),
    .I0(n236),
    .I1(key[10])
  );
  //AND U606bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U606bar (
    .O(n490bar),
    .I0(n236bar),
    .I1(keybar[10])
  );
  //AND U607
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U607 (
    .O(n489),
    .I0(key[10]),
    .I1(n236)
  );
  //OR U607bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U607bar (
    .O(n489bar),
    .I0(keybar[10]),
    .I1(n236bar)
  );
  //OR U608
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U608 (
    .O(out[109]),
    .I0(n491),
    .I1(n37)
  );
  //AND U608bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U608bar (
    .O(outbar[109]),
    .I0(n491bar),
    .I1(n37bar)
  );
  //OR U609
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U609 (
    .O(n492),
    .I0(n38),
    .I1(key[109])
  );
  //AND U609bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U609bar (
    .O(n492bar),
    .I0(n38bar),
    .I1(keybar[109])
  );
  //AND U610
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U610 (
    .O(n491),
    .I0(key[109]),
    .I1(n38)
  );
  //OR U610bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U610bar (
    .O(n491bar),
    .I0(keybar[109]),
    .I1(n38bar)
  );
  //OR U611
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U611 (
    .O(out[108]),
    .I0(n493),
    .I1(n39)
  );
  //AND U611bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U611bar (
    .O(outbar[108]),
    .I0(n493bar),
    .I1(n39bar)
  );
  //OR U612
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U612 (
    .O(n494),
    .I0(n40),
    .I1(key[108])
  );
  //AND U612bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U612bar (
    .O(n494bar),
    .I0(n40bar),
    .I1(keybar[108])
  );
  //AND U613
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U613 (
    .O(n493),
    .I0(key[108]),
    .I1(n40)
  );
  //OR U613bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U613bar (
    .O(n493bar),
    .I0(keybar[108]),
    .I1(n40bar)
  );
  //OR U614
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U614 (
    .O(out[107]),
    .I0(n495),
    .I1(n41)
  );
  //AND U614bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U614bar (
    .O(outbar[107]),
    .I0(n495bar),
    .I1(n41bar)
  );
  //OR U615
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U615 (
    .O(n496),
    .I0(n42),
    .I1(key[107])
  );
  //AND U615bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U615bar (
    .O(n496bar),
    .I0(n42bar),
    .I1(keybar[107])
  );
  //AND U616
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U616 (
    .O(n495),
    .I0(key[107]),
    .I1(n42)
  );
  //OR U616bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U616bar (
    .O(n495bar),
    .I0(keybar[107]),
    .I1(n42bar)
  );
  //OR U617
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U617 (
    .O(out[106]),
    .I0(n497),
    .I1(n43)
  );
  //AND U617bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U617bar (
    .O(outbar[106]),
    .I0(n497bar),
    .I1(n43bar)
  );
  //OR U618
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U618 (
    .O(n498),
    .I0(n44),
    .I1(key[106])
  );
  //AND U618bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U618bar (
    .O(n498bar),
    .I0(n44bar),
    .I1(keybar[106])
  );
  //AND U619
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U619 (
    .O(n497),
    .I0(key[106]),
    .I1(n44)
  );
  //OR U619bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U619bar (
    .O(n497bar),
    .I0(keybar[106]),
    .I1(n44bar)
  );
  //OR U620
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U620 (
    .O(out[105]),
    .I0(n499),
    .I1(n45)
  );
  //AND U620bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U620bar (
    .O(outbar[105]),
    .I0(n499bar),
    .I1(n45bar)
  );
  //OR U621
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U621 (
    .O(n500),
    .I0(n46),
    .I1(key[105])
  );
  //AND U621bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U621bar (
    .O(n500bar),
    .I0(n46bar),
    .I1(keybar[105])
  );
  //AND U622
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U622 (
    .O(n499),
    .I0(key[105]),
    .I1(n46)
  );
  //OR U622bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U622bar (
    .O(n499bar),
    .I0(keybar[105]),
    .I1(n46bar)
  );
  //OR U623
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U623 (
    .O(out[104]),
    .I0(n501),
    .I1(n47)
  );
  //AND U623bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U623bar (
    .O(outbar[104]),
    .I0(n501bar),
    .I1(n47bar)
  );
  //OR U624
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U624 (
    .O(n502),
    .I0(n48),
    .I1(key[104])
  );
  //AND U624bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U624bar (
    .O(n502bar),
    .I0(n48bar),
    .I1(keybar[104])
  );
  //AND U625
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U625 (
    .O(n501),
    .I0(key[104]),
    .I1(n48)
  );
  //OR U625bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U625bar (
    .O(n501bar),
    .I0(keybar[104]),
    .I1(n48bar)
  );
  //OR U626
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U626 (
    .O(out[103]),
    .I0(n503),
    .I1(n49)
  );
  //AND U626bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U626bar (
    .O(outbar[103]),
    .I0(n503bar),
    .I1(n49bar)
  );
  //OR U627
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U627 (
    .O(n504),
    .I0(n50),
    .I1(key[103])
  );
  //AND U627bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U627bar (
    .O(n504bar),
    .I0(n50bar),
    .I1(keybar[103])
  );
  //AND U628
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U628 (
    .O(n503),
    .I0(key[103]),
    .I1(n50)
  );
  //OR U628bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U628bar (
    .O(n503bar),
    .I0(keybar[103]),
    .I1(n50bar)
  );
  //OR U629
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U629 (
    .O(out[102]),
    .I0(n505),
    .I1(n51)
  );
  //AND U629bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U629bar (
    .O(outbar[102]),
    .I0(n505bar),
    .I1(n51bar)
  );
  //OR U630
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U630 (
    .O(n506),
    .I0(n52),
    .I1(key[102])
  );
  //AND U630bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U630bar (
    .O(n506bar),
    .I0(n52bar),
    .I1(keybar[102])
  );
  //AND U631
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U631 (
    .O(n505),
    .I0(key[102]),
    .I1(n52)
  );
  //OR U631bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U631bar (
    .O(n505bar),
    .I0(keybar[102]),
    .I1(n52bar)
  );
  //OR U632
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U632 (
    .O(out[101]),
    .I0(n507),
    .I1(n53)
  );
  //AND U632bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U632bar (
    .O(outbar[101]),
    .I0(n507bar),
    .I1(n53bar)
  );
  //OR U633
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U633 (
    .O(n508),
    .I0(n54),
    .I1(key[101])
  );
  //AND U633bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U633bar (
    .O(n508bar),
    .I0(n54bar),
    .I1(keybar[101])
  );
  //AND U634
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U634 (
    .O(n507),
    .I0(key[101]),
    .I1(n54)
  );
  //OR U634bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U634bar (
    .O(n507bar),
    .I0(keybar[101]),
    .I1(n54bar)
  );
  //OR U635
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U635 (
    .O(out[100]),
    .I0(n509),
    .I1(n55)
  );
  //AND U635bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U635bar (
    .O(outbar[100]),
    .I0(n509bar),
    .I1(n55bar)
  );
  //OR U636
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U636 (
    .O(n510),
    .I0(n56),
    .I1(key[100])
  );
  //AND U636bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U636bar (
    .O(n510bar),
    .I0(n56bar),
    .I1(keybar[100])
  );
  //AND U637
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U637 (
    .O(n509),
    .I0(key[100]),
    .I1(n56)
  );
  //OR U637bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U637bar (
    .O(n509bar),
    .I0(keybar[100]),
    .I1(n56bar)
  );
  //OR U638
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U638 (
    .O(out[0]),
    .I0(n511),
    .I1(n255)
  );
  //AND U638bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U638bar (
    .O(outbar[0]),
    .I0(n511bar),
    .I1(n255bar)
  );
  //OR U639
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U639 (
    .O(n512),
    .I0(n256),
    .I1(key[0])
  );
  //AND U639bar
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U639bar (
    .O(n512bar),
    .I0(n256bar),
    .I1(keybar[0])
  );
  //AND U640
  LUT2 #(
    .INIT(4'h8)
  ) LUT2_U640 (
    .O(n511),
    .I0(key[0]),
    .I1(n256)
  );
  //OR U640bar
  LUT2 #(
    .INIT(4'he)
  ) LUT2_U640bar (
    .O(n511bar),
    .I0(keybar[0]),
    .I1(n256bar)
  );
endmodule

//done
