module sample_circuit ( a, b, c, d, out );
  input a;
  input b;
  input c;
  input d;
  output out;
