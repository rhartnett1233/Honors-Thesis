`timescale 1ns / 1ps

module AND2_X1( A1, A2, ZN );
  input wire A1;
  input wire A2;
  //input_done

  output wire ZN;
  //output_done

  //wire_done

  assign ZN = A1 & A2;
endmodule


module OR2_X1( A1, A2, ZN );
  input wire A1;
  input wire A2;
  //input_done

  output wire ZN;
  //output_done

  //wire_done

  assign ZN = A1 | A2;
endmodule


module addRoundKey_Precharge ( data, databar, key, out, outbar );

  input wire [127:0] data;
  input wire [127:0] key;
  input wire [127:0] databar;
  wire [127:0] keybar;
  assign keybar[0] = ~key[0];
  assign keybar[1] = ~key[1];
  assign keybar[2] = ~key[2];
  assign keybar[3] = ~key[3];
  assign keybar[4] = ~key[4];
  assign keybar[5] = ~key[5];
  assign keybar[6] = ~key[6];
  assign keybar[7] = ~key[7];
  assign keybar[8] = ~key[8];
  assign keybar[9] = ~key[9];
  assign keybar[10] = ~key[10];
  assign keybar[11] = ~key[11];
  assign keybar[12] = ~key[12];
  assign keybar[13] = ~key[13];
  assign keybar[14] = ~key[14];
  assign keybar[15] = ~key[15];
  assign keybar[16] = ~key[16];
  assign keybar[17] = ~key[17];
  assign keybar[18] = ~key[18];
  assign keybar[19] = ~key[19];
  assign keybar[20] = ~key[20];
  assign keybar[21] = ~key[21];
  assign keybar[22] = ~key[22];
  assign keybar[23] = ~key[23];
  assign keybar[24] = ~key[24];
  assign keybar[25] = ~key[25];
  assign keybar[26] = ~key[26];
  assign keybar[27] = ~key[27];
  assign keybar[28] = ~key[28];
  assign keybar[29] = ~key[29];
  assign keybar[30] = ~key[30];
  assign keybar[31] = ~key[31];
  assign keybar[32] = ~key[32];
  assign keybar[33] = ~key[33];
  assign keybar[34] = ~key[34];
  assign keybar[35] = ~key[35];
  assign keybar[36] = ~key[36];
  assign keybar[37] = ~key[37];
  assign keybar[38] = ~key[38];
  assign keybar[39] = ~key[39];
  assign keybar[40] = ~key[40];
  assign keybar[41] = ~key[41];
  assign keybar[42] = ~key[42];
  assign keybar[43] = ~key[43];
  assign keybar[44] = ~key[44];
  assign keybar[45] = ~key[45];
  assign keybar[46] = ~key[46];
  assign keybar[47] = ~key[47];
  assign keybar[48] = ~key[48];
  assign keybar[49] = ~key[49];
  assign keybar[50] = ~key[50];
  assign keybar[51] = ~key[51];
  assign keybar[52] = ~key[52];
  assign keybar[53] = ~key[53];
  assign keybar[54] = ~key[54];
  assign keybar[55] = ~key[55];
  assign keybar[56] = ~key[56];
  assign keybar[57] = ~key[57];
  assign keybar[58] = ~key[58];
  assign keybar[59] = ~key[59];
  assign keybar[60] = ~key[60];
  assign keybar[61] = ~key[61];
  assign keybar[62] = ~key[62];
  assign keybar[63] = ~key[63];
  assign keybar[64] = ~key[64];
  assign keybar[65] = ~key[65];
  assign keybar[66] = ~key[66];
  assign keybar[67] = ~key[67];
  assign keybar[68] = ~key[68];
  assign keybar[69] = ~key[69];
  assign keybar[70] = ~key[70];
  assign keybar[71] = ~key[71];
  assign keybar[72] = ~key[72];
  assign keybar[73] = ~key[73];
  assign keybar[74] = ~key[74];
  assign keybar[75] = ~key[75];
  assign keybar[76] = ~key[76];
  assign keybar[77] = ~key[77];
  assign keybar[78] = ~key[78];
  assign keybar[79] = ~key[79];
  assign keybar[80] = ~key[80];
  assign keybar[81] = ~key[81];
  assign keybar[82] = ~key[82];
  assign keybar[83] = ~key[83];
  assign keybar[84] = ~key[84];
  assign keybar[85] = ~key[85];
  assign keybar[86] = ~key[86];
  assign keybar[87] = ~key[87];
  assign keybar[88] = ~key[88];
  assign keybar[89] = ~key[89];
  assign keybar[90] = ~key[90];
  assign keybar[91] = ~key[91];
  assign keybar[92] = ~key[92];
  assign keybar[93] = ~key[93];
  assign keybar[94] = ~key[94];
  assign keybar[95] = ~key[95];
  assign keybar[96] = ~key[96];
  assign keybar[97] = ~key[97];
  assign keybar[98] = ~key[98];
  assign keybar[99] = ~key[99];
  assign keybar[100] = ~key[100];
  assign keybar[101] = ~key[101];
  assign keybar[102] = ~key[102];
  assign keybar[103] = ~key[103];
  assign keybar[104] = ~key[104];
  assign keybar[105] = ~key[105];
  assign keybar[106] = ~key[106];
  assign keybar[107] = ~key[107];
  assign keybar[108] = ~key[108];
  assign keybar[109] = ~key[109];
  assign keybar[110] = ~key[110];
  assign keybar[111] = ~key[111];
  assign keybar[112] = ~key[112];
  assign keybar[113] = ~key[113];
  assign keybar[114] = ~key[114];
  assign keybar[115] = ~key[115];
  assign keybar[116] = ~key[116];
  assign keybar[117] = ~key[117];
  assign keybar[118] = ~key[118];
  assign keybar[119] = ~key[119];
  assign keybar[120] = ~key[120];
  assign keybar[121] = ~key[121];
  assign keybar[122] = ~key[122];
  assign keybar[123] = ~key[123];
  assign keybar[124] = ~key[124];
  assign keybar[125] = ~key[125];
  assign keybar[126] = ~key[126];
  assign keybar[127] = ~key[127];
//input_done

  output wire [127:0] out;
  output wire [127:0] outbar;
//output_done

  wire n1;
  wire n2;
  wire n3;
  wire n4;
  wire n5;
  wire n6;
  wire n7;
  wire n8;
  wire n9;
  wire n10;
  wire n11;
  wire n12;
  wire n13;
  wire n14;
  wire n15;
  wire n16;
  wire n17;
  wire n18;
  wire n19;
  wire n20;
  wire n21;
  wire n22;
  wire n23;
  wire n24;
  wire n25;
  wire n26;
  wire n27;
  wire n28;
  wire n29;
  wire n30;
  wire n31;
  wire n32;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n1bar;
  wire n2bar;
  wire n3bar;
  wire n4bar;
  wire n5bar;
  wire n6bar;
  wire n7bar;
  wire n8bar;
  wire n9bar;
  wire n10bar;
  wire n11bar;
  wire n12bar;
  wire n13bar;
  wire n14bar;
  wire n15bar;
  wire n16bar;
  wire n17bar;
  wire n18bar;
  wire n19bar;
  wire n20bar;
  wire n21bar;
  wire n22bar;
  wire n23bar;
  wire n24bar;
  wire n25bar;
  wire n26bar;
  wire n27bar;
  wire n28bar;
  wire n29bar;
  wire n30bar;
  wire n31bar;
  wire n32bar;
  wire n33bar;
  wire n34bar;
  wire n35bar;
  wire n36bar;
  wire n37bar;
  wire n38bar;
  wire n39bar;
  wire n40bar;
  wire n41bar;
  wire n42bar;
  wire n43bar;
  wire n44bar;
  wire n45bar;
  wire n46bar;
  wire n47bar;
  wire n48bar;
  wire n49bar;
  wire n50bar;
  wire n51bar;
  wire n52bar;
  wire n53bar;
  wire n54bar;
  wire n55bar;
  wire n56bar;
  wire n57bar;
  wire n58bar;
  wire n59bar;
  wire n60bar;
  wire n61bar;
  wire n62bar;
  wire n63bar;
  wire n64bar;
  wire n65bar;
  wire n66bar;
  wire n67bar;
  wire n68bar;
  wire n69bar;
  wire n70bar;
  wire n71bar;
  wire n72bar;
  wire n73bar;
  wire n74bar;
  wire n75bar;
  wire n76bar;
  wire n77bar;
  wire n78bar;
  wire n79bar;
  wire n80bar;
  wire n81bar;
  wire n82bar;
  wire n83bar;
  wire n84bar;
  wire n85bar;
  wire n86bar;
  wire n87bar;
  wire n88bar;
  wire n89bar;
  wire n90bar;
  wire n91bar;
  wire n92bar;
  wire n93bar;
  wire n94bar;
  wire n95bar;
  wire n96bar;
  wire n97bar;
  wire n98bar;
  wire n99bar;
  wire n100bar;
  wire n101bar;
  wire n102bar;
  wire n103bar;
  wire n104bar;
  wire n105bar;
  wire n106bar;
  wire n107bar;
  wire n108bar;
  wire n109bar;
  wire n110bar;
  wire n111bar;
  wire n112bar;
  wire n113bar;
  wire n114bar;
  wire n115bar;
  wire n116bar;
  wire n117bar;
  wire n118bar;
  wire n119bar;
  wire n120bar;
  wire n121bar;
  wire n122bar;
  wire n123bar;
  wire n124bar;
  wire n125bar;
  wire n126bar;
  wire n127bar;
  wire n128bar;
  wire n129bar;
  wire n130bar;
  wire n131bar;
  wire n132bar;
  wire n133bar;
  wire n134bar;
  wire n135bar;
  wire n136bar;
  wire n137bar;
  wire n138bar;
  wire n139bar;
  wire n140bar;
  wire n141bar;
  wire n142bar;
  wire n143bar;
  wire n144bar;
  wire n145bar;
  wire n146bar;
  wire n147bar;
  wire n148bar;
  wire n149bar;
  wire n150bar;
  wire n151bar;
  wire n152bar;
  wire n153bar;
  wire n154bar;
  wire n155bar;
  wire n156bar;
  wire n157bar;
  wire n158bar;
  wire n159bar;
  wire n160bar;
  wire n161bar;
  wire n162bar;
  wire n163bar;
  wire n164bar;
  wire n165bar;
  wire n166bar;
  wire n167bar;
  wire n168bar;
  wire n169bar;
  wire n170bar;
  wire n171bar;
  wire n172bar;
  wire n173bar;
  wire n174bar;
  wire n175bar;
  wire n176bar;
  wire n177bar;
  wire n178bar;
  wire n179bar;
  wire n180bar;
  wire n181bar;
  wire n182bar;
  wire n183bar;
  wire n184bar;
  wire n185bar;
  wire n186bar;
  wire n187bar;
  wire n188bar;
  wire n189bar;
  wire n190bar;
  wire n191bar;
  wire n192bar;
  wire n193bar;
  wire n194bar;
  wire n195bar;
  wire n196bar;
  wire n197bar;
  wire n198bar;
  wire n199bar;
  wire n200bar;
  wire n201bar;
  wire n202bar;
  wire n203bar;
  wire n204bar;
  wire n205bar;
  wire n206bar;
  wire n207bar;
  wire n208bar;
  wire n209bar;
  wire n210bar;
  wire n211bar;
  wire n212bar;
  wire n213bar;
  wire n214bar;
  wire n215bar;
  wire n216bar;
  wire n217bar;
  wire n218bar;
  wire n219bar;
  wire n220bar;
  wire n221bar;
  wire n222bar;
  wire n223bar;
  wire n224bar;
  wire n225bar;
  wire n226bar;
  wire n227bar;
  wire n228bar;
  wire n229bar;
  wire n230bar;
  wire n231bar;
  wire n232bar;
  wire n233bar;
  wire n234bar;
  wire n235bar;
  wire n236bar;
  wire n237bar;
  wire n238bar;
  wire n239bar;
  wire n240bar;
  wire n241bar;
  wire n242bar;
  wire n243bar;
  wire n244bar;
  wire n245bar;
  wire n246bar;
  wire n247bar;
  wire n248bar;
  wire n249bar;
  wire n250bar;
  wire n251bar;
  wire n252bar;
  wire n253bar;
  wire n254bar;
  wire n255bar;
  wire n256bar;
  wire n257bar;
  wire n258bar;
  wire n259bar;
  wire n260bar;
  wire n261bar;
  wire n262bar;
  wire n263bar;
  wire n264bar;
  wire n265bar;
  wire n266bar;
  wire n267bar;
  wire n268bar;
  wire n269bar;
  wire n270bar;
  wire n271bar;
  wire n272bar;
  wire n273bar;
  wire n274bar;
  wire n275bar;
  wire n276bar;
  wire n277bar;
  wire n278bar;
  wire n279bar;
  wire n280bar;
  wire n281bar;
  wire n282bar;
  wire n283bar;
  wire n284bar;
  wire n285bar;
  wire n286bar;
  wire n287bar;
  wire n288bar;
  wire n289bar;
  wire n290bar;
  wire n291bar;
  wire n292bar;
  wire n293bar;
  wire n294bar;
  wire n295bar;
  wire n296bar;
  wire n297bar;
  wire n298bar;
  wire n299bar;
  wire n300bar;
  wire n301bar;
  wire n302bar;
  wire n303bar;
  wire n304bar;
  wire n305bar;
  wire n306bar;
  wire n307bar;
  wire n308bar;
  wire n309bar;
  wire n310bar;
  wire n311bar;
  wire n312bar;
  wire n313bar;
  wire n314bar;
  wire n315bar;
  wire n316bar;
  wire n317bar;
  wire n318bar;
  wire n319bar;
  wire n320bar;
  wire n321bar;
  wire n322bar;
  wire n323bar;
  wire n324bar;
  wire n325bar;
  wire n326bar;
  wire n327bar;
  wire n328bar;
  wire n329bar;
  wire n330bar;
  wire n331bar;
  wire n332bar;
  wire n333bar;
  wire n334bar;
  wire n335bar;
  wire n336bar;
  wire n337bar;
  wire n338bar;
  wire n339bar;
  wire n340bar;
  wire n341bar;
  wire n342bar;
  wire n343bar;
  wire n344bar;
  wire n345bar;
  wire n346bar;
  wire n347bar;
  wire n348bar;
  wire n349bar;
  wire n350bar;
  wire n351bar;
  wire n352bar;
  wire n353bar;
  wire n354bar;
  wire n355bar;
  wire n356bar;
  wire n357bar;
  wire n358bar;
  wire n359bar;
  wire n360bar;
  wire n361bar;
  wire n362bar;
  wire n363bar;
  wire n364bar;
  wire n365bar;
  wire n366bar;
  wire n367bar;
  wire n368bar;
  wire n369bar;
  wire n370bar;
  wire n371bar;
  wire n372bar;
  wire n373bar;
  wire n374bar;
  wire n375bar;
  wire n376bar;
  wire n377bar;
  wire n378bar;
  wire n379bar;
  wire n380bar;
  wire n381bar;
  wire n382bar;
  wire n383bar;
  wire n384bar;
  wire n385bar;
  wire n386bar;
  wire n387bar;
  wire n388bar;
  wire n389bar;
  wire n390bar;
  wire n391bar;
  wire n392bar;
  wire n393bar;
  wire n394bar;
  wire n395bar;
  wire n396bar;
  wire n397bar;
  wire n398bar;
  wire n399bar;
  wire n400bar;
  wire n401bar;
  wire n402bar;
  wire n403bar;
  wire n404bar;
  wire n405bar;
  wire n406bar;
  wire n407bar;
  wire n408bar;
  wire n409bar;
  wire n410bar;
  wire n411bar;
  wire n412bar;
  wire n413bar;
  wire n414bar;
  wire n415bar;
  wire n416bar;
  wire n417bar;
  wire n418bar;
  wire n419bar;
  wire n420bar;
  wire n421bar;
  wire n422bar;
  wire n423bar;
  wire n424bar;
  wire n425bar;
  wire n426bar;
  wire n427bar;
  wire n428bar;
  wire n429bar;
  wire n430bar;
  wire n431bar;
  wire n432bar;
  wire n433bar;
  wire n434bar;
  wire n435bar;
  wire n436bar;
  wire n437bar;
  wire n438bar;
  wire n439bar;
  wire n440bar;
  wire n441bar;
  wire n442bar;
  wire n443bar;
  wire n444bar;
  wire n445bar;
  wire n446bar;
  wire n447bar;
  wire n448bar;
  wire n449bar;
  wire n450bar;
  wire n451bar;
  wire n452bar;
  wire n453bar;
  wire n454bar;
  wire n455bar;
  wire n456bar;
  wire n457bar;
  wire n458bar;
  wire n459bar;
  wire n460bar;
  wire n461bar;
  wire n462bar;
  wire n463bar;
  wire n464bar;
  wire n465bar;
  wire n466bar;
  wire n467bar;
  wire n468bar;
  wire n469bar;
  wire n470bar;
  wire n471bar;
  wire n472bar;
  wire n473bar;
  wire n474bar;
  wire n475bar;
  wire n476bar;
  wire n477bar;
  wire n478bar;
  wire n479bar;
  wire n480bar;
  wire n481bar;
  wire n482bar;
  wire n483bar;
  wire n484bar;
  wire n485bar;
  wire n486bar;
  wire n487bar;
  wire n488bar;
  wire n489bar;
  wire n490bar;
  wire n491bar;
  wire n492bar;
  wire n493bar;
  wire n494bar;
  wire n495bar;
  wire n496bar;
  wire n497bar;
  wire n498bar;
  wire n499bar;
  wire n500bar;
  wire n501bar;
  wire n502bar;
  wire n503bar;
  wire n504bar;
  wire n505bar;
  wire n506bar;
  wire n507bar;
  wire n508bar;
  wire n509bar;
  wire n510bar;
  wire n511bar;
  wire n512bar;
//wire_done

 //assign_done

  assign n1bar = n452;
  assign n1 = n452bar;
  assign n2bar = data[127];
  assign n2 = databar[127];
  assign n3bar = n454;
  assign n3 = n454bar;
  assign n4bar = data[126];
  assign n4 = databar[126];
  assign n5bar = n456;
  assign n5 = n456bar;
  assign n6bar = data[125];
  assign n6 = databar[125];
  assign n7bar = n458;
  assign n7 = n458bar;
  assign n8bar = data[124];
  assign n8 = databar[124];
  assign n9bar = n460;
  assign n9 = n460bar;
  assign n10bar = data[123];
  assign n10 = databar[123];
  assign n11bar = n462;
  assign n11 = n462bar;
  assign n12bar = data[122];
  assign n12 = databar[122];
  assign n13bar = n464;
  assign n13 = n464bar;
  assign n14bar = data[121];
  assign n14 = databar[121];
  assign n15bar = n466;
  assign n15 = n466bar;
  assign n16bar = data[120];
  assign n16 = databar[120];
  assign n17bar = n470;
  assign n17 = n470bar;
  assign n18bar = data[119];
  assign n18 = databar[119];
  assign n19bar = n472;
  assign n19 = n472bar;
  assign n20bar = data[118];
  assign n20 = databar[118];
  assign n21bar = n474;
  assign n21 = n474bar;
  assign n22bar = data[117];
  assign n22 = databar[117];
  assign n23bar = n476;
  assign n23 = n476bar;
  assign n24bar = data[116];
  assign n24 = databar[116];
  assign n25bar = n478;
  assign n25 = n478bar;
  assign n26bar = data[115];
  assign n26 = databar[115];
  assign n27bar = n480;
  assign n27 = n480bar;
  assign n28bar = data[114];
  assign n28 = databar[114];
  assign n29bar = n482;
  assign n29 = n482bar;
  assign n30bar = data[113];
  assign n30 = databar[113];
  assign n31bar = n484;
  assign n31 = n484bar;
  assign n32bar = data[112];
  assign n32 = databar[112];
  assign n33bar = n486;
  assign n33 = n486bar;
  assign n34bar = data[111];
  assign n34 = databar[111];
  assign n35bar = n488;
  assign n35 = n488bar;
  assign n36bar = data[110];
  assign n36 = databar[110];
  assign n37bar = n492;
  assign n37 = n492bar;
  assign n38bar = data[109];
  assign n38 = databar[109];
  assign n39bar = n494;
  assign n39 = n494bar;
  assign n40bar = data[108];
  assign n40 = databar[108];
  assign n41bar = n496;
  assign n41 = n496bar;
  assign n42bar = data[107];
  assign n42 = databar[107];
  assign n43bar = n498;
  assign n43 = n498bar;
  assign n44bar = data[106];
  assign n44 = databar[106];
  assign n45bar = n500;
  assign n45 = n500bar;
  assign n46bar = data[105];
  assign n46 = databar[105];
  assign n47bar = n502;
  assign n47 = n502bar;
  assign n48bar = data[104];
  assign n48 = databar[104];
  assign n49bar = n504;
  assign n49 = n504bar;
  assign n50bar = data[103];
  assign n50 = databar[103];
  assign n51bar = n506;
  assign n51 = n506bar;
  assign n52bar = data[102];
  assign n52 = databar[102];
  assign n53bar = n508;
  assign n53 = n508bar;
  assign n54bar = data[101];
  assign n54 = databar[101];
  assign n55bar = n510;
  assign n55 = n510bar;
  assign n56bar = data[100];
  assign n56 = databar[100];
  assign n57bar = n260;
  assign n57 = n260bar;
  assign n58bar = data[99];
  assign n58 = databar[99];
  assign n59bar = n262;
  assign n59 = n262bar;
  assign n60bar = data[98];
  assign n60 = databar[98];
  assign n61bar = n264;
  assign n61 = n264bar;
  assign n62bar = data[97];
  assign n62 = databar[97];
  assign n63bar = n266;
  assign n63 = n266bar;
  assign n64bar = data[96];
  assign n64 = databar[96];
  assign n65bar = n268;
  assign n65 = n268bar;
  assign n66bar = data[95];
  assign n66 = databar[95];
  assign n67bar = n270;
  assign n67 = n270bar;
  assign n68bar = data[94];
  assign n68 = databar[94];
  assign n69bar = n272;
  assign n69 = n272bar;
  assign n70bar = data[93];
  assign n70 = databar[93];
  assign n71bar = n274;
  assign n71 = n274bar;
  assign n72bar = data[92];
  assign n72 = databar[92];
  assign n73bar = n276;
  assign n73 = n276bar;
  assign n74bar = data[91];
  assign n74 = databar[91];
  assign n75bar = n278;
  assign n75 = n278bar;
  assign n76bar = data[90];
  assign n76 = databar[90];
  assign n77bar = n282;
  assign n77 = n282bar;
  assign n78bar = data[89];
  assign n78 = databar[89];
  assign n79bar = n284;
  assign n79 = n284bar;
  assign n80bar = data[88];
  assign n80 = databar[88];
  assign n81bar = n286;
  assign n81 = n286bar;
  assign n82bar = data[87];
  assign n82 = databar[87];
  assign n83bar = n288;
  assign n83 = n288bar;
  assign n84bar = data[86];
  assign n84 = databar[86];
  assign n85bar = n290;
  assign n85 = n290bar;
  assign n86bar = data[85];
  assign n86 = databar[85];
  assign n87bar = n292;
  assign n87 = n292bar;
  assign n88bar = data[84];
  assign n88 = databar[84];
  assign n89bar = n294;
  assign n89 = n294bar;
  assign n90bar = data[83];
  assign n90 = databar[83];
  assign n91bar = n296;
  assign n91 = n296bar;
  assign n92bar = data[82];
  assign n92 = databar[82];
  assign n93bar = n298;
  assign n93 = n298bar;
  assign n94bar = data[81];
  assign n94 = databar[81];
  assign n95bar = n300;
  assign n95 = n300bar;
  assign n96bar = data[80];
  assign n96 = databar[80];
  assign n97bar = n304;
  assign n97 = n304bar;
  assign n98bar = data[79];
  assign n98 = databar[79];
  assign n99bar = n306;
  assign n99 = n306bar;
  assign n100bar = data[78];
  assign n100 = databar[78];
  assign n101bar = n308;
  assign n101 = n308bar;
  assign n102bar = data[77];
  assign n102 = databar[77];
  assign n103bar = n310;
  assign n103 = n310bar;
  assign n104bar = data[76];
  assign n104 = databar[76];
  assign n105bar = n312;
  assign n105 = n312bar;
  assign n106bar = data[75];
  assign n106 = databar[75];
  assign n107bar = n314;
  assign n107 = n314bar;
  assign n108bar = data[74];
  assign n108 = databar[74];
  assign n109bar = n316;
  assign n109 = n316bar;
  assign n110bar = data[73];
  assign n110 = databar[73];
  assign n111bar = n318;
  assign n111 = n318bar;
  assign n112bar = data[72];
  assign n112 = databar[72];
  assign n113bar = n320;
  assign n113 = n320bar;
  assign n114bar = data[71];
  assign n114 = databar[71];
  assign n115bar = n322;
  assign n115 = n322bar;
  assign n116bar = data[70];
  assign n116 = databar[70];
  assign n117bar = n326;
  assign n117 = n326bar;
  assign n118bar = data[69];
  assign n118 = databar[69];
  assign n119bar = n328;
  assign n119 = n328bar;
  assign n120bar = data[68];
  assign n120 = databar[68];
  assign n121bar = n330;
  assign n121 = n330bar;
  assign n122bar = data[67];
  assign n122 = databar[67];
  assign n123bar = n332;
  assign n123 = n332bar;
  assign n124bar = data[66];
  assign n124 = databar[66];
  assign n125bar = n334;
  assign n125 = n334bar;
  assign n126bar = data[65];
  assign n126 = databar[65];
  assign n127bar = n336;
  assign n127 = n336bar;
  assign n128bar = data[64];
  assign n128 = databar[64];
  assign n129bar = n338;
  assign n129 = n338bar;
  assign n130bar = data[63];
  assign n130 = databar[63];
  assign n131bar = n340;
  assign n131 = n340bar;
  assign n132bar = data[62];
  assign n132 = databar[62];
  assign n133bar = n342;
  assign n133 = n342bar;
  assign n134bar = data[61];
  assign n134 = databar[61];
  assign n135bar = n344;
  assign n135 = n344bar;
  assign n136bar = data[60];
  assign n136 = databar[60];
  assign n137bar = n348;
  assign n137 = n348bar;
  assign n138bar = data[59];
  assign n138 = databar[59];
  assign n139bar = n350;
  assign n139 = n350bar;
  assign n140bar = data[58];
  assign n140 = databar[58];
  assign n141bar = n352;
  assign n141 = n352bar;
  assign n142bar = data[57];
  assign n142 = databar[57];
  assign n143bar = n354;
  assign n143 = n354bar;
  assign n144bar = data[56];
  assign n144 = databar[56];
  assign n145bar = n356;
  assign n145 = n356bar;
  assign n146bar = data[55];
  assign n146 = databar[55];
  assign n147bar = n358;
  assign n147 = n358bar;
  assign n148bar = data[54];
  assign n148 = databar[54];
  assign n149bar = n360;
  assign n149 = n360bar;
  assign n150bar = data[53];
  assign n150 = databar[53];
  assign n151bar = n362;
  assign n151 = n362bar;
  assign n152bar = data[52];
  assign n152 = databar[52];
  assign n153bar = n364;
  assign n153 = n364bar;
  assign n154bar = data[51];
  assign n154 = databar[51];
  assign n155bar = n366;
  assign n155 = n366bar;
  assign n156bar = data[50];
  assign n156 = databar[50];
  assign n157bar = n370;
  assign n157 = n370bar;
  assign n158bar = data[49];
  assign n158 = databar[49];
  assign n159bar = n372;
  assign n159 = n372bar;
  assign n160bar = data[48];
  assign n160 = databar[48];
  assign n161bar = n374;
  assign n161 = n374bar;
  assign n162bar = data[47];
  assign n162 = databar[47];
  assign n163bar = n376;
  assign n163 = n376bar;
  assign n164bar = data[46];
  assign n164 = databar[46];
  assign n165bar = n378;
  assign n165 = n378bar;
  assign n166bar = data[45];
  assign n166 = databar[45];
  assign n167bar = n380;
  assign n167 = n380bar;
  assign n168bar = data[44];
  assign n168 = databar[44];
  assign n169bar = n382;
  assign n169 = n382bar;
  assign n170bar = data[43];
  assign n170 = databar[43];
  assign n171bar = n384;
  assign n171 = n384bar;
  assign n172bar = data[42];
  assign n172 = databar[42];
  assign n173bar = n386;
  assign n173 = n386bar;
  assign n174bar = data[41];
  assign n174 = databar[41];
  assign n175bar = n388;
  assign n175 = n388bar;
  assign n176bar = data[40];
  assign n176 = databar[40];
  assign n177bar = n392;
  assign n177 = n392bar;
  assign n178bar = data[39];
  assign n178 = databar[39];
  assign n179bar = n394;
  assign n179 = n394bar;
  assign n180bar = data[38];
  assign n180 = databar[38];
  assign n181bar = n396;
  assign n181 = n396bar;
  assign n182bar = data[37];
  assign n182 = databar[37];
  assign n183bar = n398;
  assign n183 = n398bar;
  assign n184bar = data[36];
  assign n184 = databar[36];
  assign n185bar = n400;
  assign n185 = n400bar;
  assign n186bar = data[35];
  assign n186 = databar[35];
  assign n187bar = n402;
  assign n187 = n402bar;
  assign n188bar = data[34];
  assign n188 = databar[34];
  assign n189bar = n404;
  assign n189 = n404bar;
  assign n190bar = data[33];
  assign n190 = databar[33];
  assign n191bar = n406;
  assign n191 = n406bar;
  assign n192bar = data[32];
  assign n192 = databar[32];
  assign n193bar = n408;
  assign n193 = n408bar;
  assign n194bar = data[31];
  assign n194 = databar[31];
  assign n195bar = n410;
  assign n195 = n410bar;
  assign n196bar = data[30];
  assign n196 = databar[30];
  assign n197bar = n414;
  assign n197 = n414bar;
  assign n198bar = data[29];
  assign n198 = databar[29];
  assign n199bar = n416;
  assign n199 = n416bar;
  assign n200bar = data[28];
  assign n200 = databar[28];
  assign n201bar = n418;
  assign n201 = n418bar;
  assign n202bar = data[27];
  assign n202 = databar[27];
  assign n203bar = n420;
  assign n203 = n420bar;
  assign n204bar = data[26];
  assign n204 = databar[26];
  assign n205bar = n422;
  assign n205 = n422bar;
  assign n206bar = data[25];
  assign n206 = databar[25];
  assign n207bar = n424;
  assign n207 = n424bar;
  assign n208bar = data[24];
  assign n208 = databar[24];
  assign n209bar = n426;
  assign n209 = n426bar;
  assign n210bar = data[23];
  assign n210 = databar[23];
  assign n211bar = n428;
  assign n211 = n428bar;
  assign n212bar = data[22];
  assign n212 = databar[22];
  assign n213bar = n430;
  assign n213 = n430bar;
  assign n214bar = data[21];
  assign n214 = databar[21];
  assign n215bar = n432;
  assign n215 = n432bar;
  assign n216bar = data[20];
  assign n216 = databar[20];
  assign n217bar = n436;
  assign n217 = n436bar;
  assign n218bar = data[19];
  assign n218 = databar[19];
  assign n219bar = n438;
  assign n219 = n438bar;
  assign n220bar = data[18];
  assign n220 = databar[18];
  assign n221bar = n440;
  assign n221 = n440bar;
  assign n222bar = data[17];
  assign n222 = databar[17];
  assign n223bar = n442;
  assign n223 = n442bar;
  assign n224bar = data[16];
  assign n224 = databar[16];
  assign n225bar = n444;
  assign n225 = n444bar;
  assign n226bar = data[15];
  assign n226 = databar[15];
  assign n227bar = n446;
  assign n227 = n446bar;
  assign n228bar = data[14];
  assign n228 = databar[14];
  assign n229bar = n448;
  assign n229 = n448bar;
  assign n230bar = data[13];
  assign n230 = databar[13];
  assign n231bar = n450;
  assign n231 = n450bar;
  assign n232bar = data[12];
  assign n232 = databar[12];
  assign n233bar = n468;
  assign n233 = n468bar;
  assign n234bar = data[11];
  assign n234 = databar[11];
  assign n235bar = n490;
  assign n235 = n490bar;
  assign n236bar = data[10];
  assign n236 = databar[10];
  assign n237bar = n258;
  assign n237 = n258bar;
  assign n238bar = data[9];
  assign n238 = databar[9];
  assign n239bar = n280;
  assign n239 = n280bar;
  assign n240bar = data[8];
  assign n240 = databar[8];
  assign n241bar = n302;
  assign n241 = n302bar;
  assign n242bar = data[7];
  assign n242 = databar[7];
  assign n243bar = n324;
  assign n243 = n324bar;
  assign n244bar = data[6];
  assign n244 = databar[6];
  assign n245bar = n346;
  assign n245 = n346bar;
  assign n246bar = data[5];
  assign n246 = databar[5];
  assign n247bar = n368;
  assign n247 = n368bar;
  assign n248bar = data[4];
  assign n248 = databar[4];
  assign n249bar = n390;
  assign n249 = n390bar;
  assign n250bar = data[3];
  assign n250 = databar[3];
  assign n251bar = n412;
  assign n251 = n412bar;
  assign n252bar = data[2];
  assign n252 = databar[2];
  assign n253bar = n434;
  assign n253 = n434bar;
  assign n254bar = data[1];
  assign n254 = databar[1];
  assign n255bar = n512;
  assign n255 = n512bar;
  assign n256bar = data[0];
  assign n256 = databar[0];
  OR2_X1 U257 ( .A1(n257), .A2(n237), .ZN(out[9]) );
  AND2_X1 U257bar ( .A1(n257bar), .A2(n237bar), .ZN(outbar[9]) );
  OR2_X1 U258 ( .A1(n238), .A2(key[9]), .ZN(n258) );
  AND2_X1 U258bar ( .A1(n238bar), .A2(keybar[9]), .ZN(n258bar) );
  AND2_X1 U259 ( .A1(key[9]), .A2(n238), .ZN(n257) );
  OR2_X1 U259bar ( .A1(keybar[9]), .A2(n238bar), .ZN(n257bar) );
  OR2_X1 U260 ( .A1(n259), .A2(n57), .ZN(out[99]) );
  AND2_X1 U260bar ( .A1(n259bar), .A2(n57bar), .ZN(outbar[99]) );
  OR2_X1 U261 ( .A1(n58), .A2(key[99]), .ZN(n260) );
  AND2_X1 U261bar ( .A1(n58bar), .A2(keybar[99]), .ZN(n260bar) );
  AND2_X1 U262 ( .A1(key[99]), .A2(n58), .ZN(n259) );
  OR2_X1 U262bar ( .A1(keybar[99]), .A2(n58bar), .ZN(n259bar) );
  OR2_X1 U263 ( .A1(n261), .A2(n59), .ZN(out[98]) );
  AND2_X1 U263bar ( .A1(n261bar), .A2(n59bar), .ZN(outbar[98]) );
  OR2_X1 U264 ( .A1(n60), .A2(key[98]), .ZN(n262) );
  AND2_X1 U264bar ( .A1(n60bar), .A2(keybar[98]), .ZN(n262bar) );
  AND2_X1 U265 ( .A1(key[98]), .A2(n60), .ZN(n261) );
  OR2_X1 U265bar ( .A1(keybar[98]), .A2(n60bar), .ZN(n261bar) );
  OR2_X1 U266 ( .A1(n263), .A2(n61), .ZN(out[97]) );
  AND2_X1 U266bar ( .A1(n263bar), .A2(n61bar), .ZN(outbar[97]) );
  OR2_X1 U267 ( .A1(n62), .A2(key[97]), .ZN(n264) );
  AND2_X1 U267bar ( .A1(n62bar), .A2(keybar[97]), .ZN(n264bar) );
  AND2_X1 U268 ( .A1(key[97]), .A2(n62), .ZN(n263) );
  OR2_X1 U268bar ( .A1(keybar[97]), .A2(n62bar), .ZN(n263bar) );
  OR2_X1 U269 ( .A1(n265), .A2(n63), .ZN(out[96]) );
  AND2_X1 U269bar ( .A1(n265bar), .A2(n63bar), .ZN(outbar[96]) );
  OR2_X1 U270 ( .A1(n64), .A2(key[96]), .ZN(n266) );
  AND2_X1 U270bar ( .A1(n64bar), .A2(keybar[96]), .ZN(n266bar) );
  AND2_X1 U271 ( .A1(key[96]), .A2(n64), .ZN(n265) );
  OR2_X1 U271bar ( .A1(keybar[96]), .A2(n64bar), .ZN(n265bar) );
  OR2_X1 U272 ( .A1(n267), .A2(n65), .ZN(out[95]) );
  AND2_X1 U272bar ( .A1(n267bar), .A2(n65bar), .ZN(outbar[95]) );
  OR2_X1 U273 ( .A1(n66), .A2(key[95]), .ZN(n268) );
  AND2_X1 U273bar ( .A1(n66bar), .A2(keybar[95]), .ZN(n268bar) );
  AND2_X1 U274 ( .A1(key[95]), .A2(n66), .ZN(n267) );
  OR2_X1 U274bar ( .A1(keybar[95]), .A2(n66bar), .ZN(n267bar) );
  OR2_X1 U275 ( .A1(n269), .A2(n67), .ZN(out[94]) );
  AND2_X1 U275bar ( .A1(n269bar), .A2(n67bar), .ZN(outbar[94]) );
  OR2_X1 U276 ( .A1(n68), .A2(key[94]), .ZN(n270) );
  AND2_X1 U276bar ( .A1(n68bar), .A2(keybar[94]), .ZN(n270bar) );
  AND2_X1 U277 ( .A1(key[94]), .A2(n68), .ZN(n269) );
  OR2_X1 U277bar ( .A1(keybar[94]), .A2(n68bar), .ZN(n269bar) );
  OR2_X1 U278 ( .A1(n271), .A2(n69), .ZN(out[93]) );
  AND2_X1 U278bar ( .A1(n271bar), .A2(n69bar), .ZN(outbar[93]) );
  OR2_X1 U279 ( .A1(n70), .A2(key[93]), .ZN(n272) );
  AND2_X1 U279bar ( .A1(n70bar), .A2(keybar[93]), .ZN(n272bar) );
  AND2_X1 U280 ( .A1(key[93]), .A2(n70), .ZN(n271) );
  OR2_X1 U280bar ( .A1(keybar[93]), .A2(n70bar), .ZN(n271bar) );
  OR2_X1 U281 ( .A1(n273), .A2(n71), .ZN(out[92]) );
  AND2_X1 U281bar ( .A1(n273bar), .A2(n71bar), .ZN(outbar[92]) );
  OR2_X1 U282 ( .A1(n72), .A2(key[92]), .ZN(n274) );
  AND2_X1 U282bar ( .A1(n72bar), .A2(keybar[92]), .ZN(n274bar) );
  AND2_X1 U283 ( .A1(key[92]), .A2(n72), .ZN(n273) );
  OR2_X1 U283bar ( .A1(keybar[92]), .A2(n72bar), .ZN(n273bar) );
  OR2_X1 U284 ( .A1(n275), .A2(n73), .ZN(out[91]) );
  AND2_X1 U284bar ( .A1(n275bar), .A2(n73bar), .ZN(outbar[91]) );
  OR2_X1 U285 ( .A1(n74), .A2(key[91]), .ZN(n276) );
  AND2_X1 U285bar ( .A1(n74bar), .A2(keybar[91]), .ZN(n276bar) );
  AND2_X1 U286 ( .A1(key[91]), .A2(n74), .ZN(n275) );
  OR2_X1 U286bar ( .A1(keybar[91]), .A2(n74bar), .ZN(n275bar) );
  OR2_X1 U287 ( .A1(n277), .A2(n75), .ZN(out[90]) );
  AND2_X1 U287bar ( .A1(n277bar), .A2(n75bar), .ZN(outbar[90]) );
  OR2_X1 U288 ( .A1(n76), .A2(key[90]), .ZN(n278) );
  AND2_X1 U288bar ( .A1(n76bar), .A2(keybar[90]), .ZN(n278bar) );
  AND2_X1 U289 ( .A1(key[90]), .A2(n76), .ZN(n277) );
  OR2_X1 U289bar ( .A1(keybar[90]), .A2(n76bar), .ZN(n277bar) );
  OR2_X1 U290 ( .A1(n279), .A2(n239), .ZN(out[8]) );
  AND2_X1 U290bar ( .A1(n279bar), .A2(n239bar), .ZN(outbar[8]) );
  OR2_X1 U291 ( .A1(n240), .A2(key[8]), .ZN(n280) );
  AND2_X1 U291bar ( .A1(n240bar), .A2(keybar[8]), .ZN(n280bar) );
  AND2_X1 U292 ( .A1(key[8]), .A2(n240), .ZN(n279) );
  OR2_X1 U292bar ( .A1(keybar[8]), .A2(n240bar), .ZN(n279bar) );
  OR2_X1 U293 ( .A1(n281), .A2(n77), .ZN(out[89]) );
  AND2_X1 U293bar ( .A1(n281bar), .A2(n77bar), .ZN(outbar[89]) );
  OR2_X1 U294 ( .A1(n78), .A2(key[89]), .ZN(n282) );
  AND2_X1 U294bar ( .A1(n78bar), .A2(keybar[89]), .ZN(n282bar) );
  AND2_X1 U295 ( .A1(key[89]), .A2(n78), .ZN(n281) );
  OR2_X1 U295bar ( .A1(keybar[89]), .A2(n78bar), .ZN(n281bar) );
  OR2_X1 U296 ( .A1(n283), .A2(n79), .ZN(out[88]) );
  AND2_X1 U296bar ( .A1(n283bar), .A2(n79bar), .ZN(outbar[88]) );
  OR2_X1 U297 ( .A1(n80), .A2(key[88]), .ZN(n284) );
  AND2_X1 U297bar ( .A1(n80bar), .A2(keybar[88]), .ZN(n284bar) );
  AND2_X1 U298 ( .A1(key[88]), .A2(n80), .ZN(n283) );
  OR2_X1 U298bar ( .A1(keybar[88]), .A2(n80bar), .ZN(n283bar) );
  OR2_X1 U299 ( .A1(n285), .A2(n81), .ZN(out[87]) );
  AND2_X1 U299bar ( .A1(n285bar), .A2(n81bar), .ZN(outbar[87]) );
  OR2_X1 U300 ( .A1(n82), .A2(key[87]), .ZN(n286) );
  AND2_X1 U300bar ( .A1(n82bar), .A2(keybar[87]), .ZN(n286bar) );
  AND2_X1 U301 ( .A1(key[87]), .A2(n82), .ZN(n285) );
  OR2_X1 U301bar ( .A1(keybar[87]), .A2(n82bar), .ZN(n285bar) );
  OR2_X1 U302 ( .A1(n287), .A2(n83), .ZN(out[86]) );
  AND2_X1 U302bar ( .A1(n287bar), .A2(n83bar), .ZN(outbar[86]) );
  OR2_X1 U303 ( .A1(n84), .A2(key[86]), .ZN(n288) );
  AND2_X1 U303bar ( .A1(n84bar), .A2(keybar[86]), .ZN(n288bar) );
  AND2_X1 U304 ( .A1(key[86]), .A2(n84), .ZN(n287) );
  OR2_X1 U304bar ( .A1(keybar[86]), .A2(n84bar), .ZN(n287bar) );
  OR2_X1 U305 ( .A1(n289), .A2(n85), .ZN(out[85]) );
  AND2_X1 U305bar ( .A1(n289bar), .A2(n85bar), .ZN(outbar[85]) );
  OR2_X1 U306 ( .A1(n86), .A2(key[85]), .ZN(n290) );
  AND2_X1 U306bar ( .A1(n86bar), .A2(keybar[85]), .ZN(n290bar) );
  AND2_X1 U307 ( .A1(key[85]), .A2(n86), .ZN(n289) );
  OR2_X1 U307bar ( .A1(keybar[85]), .A2(n86bar), .ZN(n289bar) );
  OR2_X1 U308 ( .A1(n291), .A2(n87), .ZN(out[84]) );
  AND2_X1 U308bar ( .A1(n291bar), .A2(n87bar), .ZN(outbar[84]) );
  OR2_X1 U309 ( .A1(n88), .A2(key[84]), .ZN(n292) );
  AND2_X1 U309bar ( .A1(n88bar), .A2(keybar[84]), .ZN(n292bar) );
  AND2_X1 U310 ( .A1(key[84]), .A2(n88), .ZN(n291) );
  OR2_X1 U310bar ( .A1(keybar[84]), .A2(n88bar), .ZN(n291bar) );
  OR2_X1 U311 ( .A1(n293), .A2(n89), .ZN(out[83]) );
  AND2_X1 U311bar ( .A1(n293bar), .A2(n89bar), .ZN(outbar[83]) );
  OR2_X1 U312 ( .A1(n90), .A2(key[83]), .ZN(n294) );
  AND2_X1 U312bar ( .A1(n90bar), .A2(keybar[83]), .ZN(n294bar) );
  AND2_X1 U313 ( .A1(key[83]), .A2(n90), .ZN(n293) );
  OR2_X1 U313bar ( .A1(keybar[83]), .A2(n90bar), .ZN(n293bar) );
  OR2_X1 U314 ( .A1(n295), .A2(n91), .ZN(out[82]) );
  AND2_X1 U314bar ( .A1(n295bar), .A2(n91bar), .ZN(outbar[82]) );
  OR2_X1 U315 ( .A1(n92), .A2(key[82]), .ZN(n296) );
  AND2_X1 U315bar ( .A1(n92bar), .A2(keybar[82]), .ZN(n296bar) );
  AND2_X1 U316 ( .A1(key[82]), .A2(n92), .ZN(n295) );
  OR2_X1 U316bar ( .A1(keybar[82]), .A2(n92bar), .ZN(n295bar) );
  OR2_X1 U317 ( .A1(n297), .A2(n93), .ZN(out[81]) );
  AND2_X1 U317bar ( .A1(n297bar), .A2(n93bar), .ZN(outbar[81]) );
  OR2_X1 U318 ( .A1(n94), .A2(key[81]), .ZN(n298) );
  AND2_X1 U318bar ( .A1(n94bar), .A2(keybar[81]), .ZN(n298bar) );
  AND2_X1 U319 ( .A1(key[81]), .A2(n94), .ZN(n297) );
  OR2_X1 U319bar ( .A1(keybar[81]), .A2(n94bar), .ZN(n297bar) );
  OR2_X1 U320 ( .A1(n299), .A2(n95), .ZN(out[80]) );
  AND2_X1 U320bar ( .A1(n299bar), .A2(n95bar), .ZN(outbar[80]) );
  OR2_X1 U321 ( .A1(n96), .A2(key[80]), .ZN(n300) );
  AND2_X1 U321bar ( .A1(n96bar), .A2(keybar[80]), .ZN(n300bar) );
  AND2_X1 U322 ( .A1(key[80]), .A2(n96), .ZN(n299) );
  OR2_X1 U322bar ( .A1(keybar[80]), .A2(n96bar), .ZN(n299bar) );
  OR2_X1 U323 ( .A1(n301), .A2(n241), .ZN(out[7]) );
  AND2_X1 U323bar ( .A1(n301bar), .A2(n241bar), .ZN(outbar[7]) );
  OR2_X1 U324 ( .A1(n242), .A2(key[7]), .ZN(n302) );
  AND2_X1 U324bar ( .A1(n242bar), .A2(keybar[7]), .ZN(n302bar) );
  AND2_X1 U325 ( .A1(key[7]), .A2(n242), .ZN(n301) );
  OR2_X1 U325bar ( .A1(keybar[7]), .A2(n242bar), .ZN(n301bar) );
  OR2_X1 U326 ( .A1(n303), .A2(n97), .ZN(out[79]) );
  AND2_X1 U326bar ( .A1(n303bar), .A2(n97bar), .ZN(outbar[79]) );
  OR2_X1 U327 ( .A1(n98), .A2(key[79]), .ZN(n304) );
  AND2_X1 U327bar ( .A1(n98bar), .A2(keybar[79]), .ZN(n304bar) );
  AND2_X1 U328 ( .A1(key[79]), .A2(n98), .ZN(n303) );
  OR2_X1 U328bar ( .A1(keybar[79]), .A2(n98bar), .ZN(n303bar) );
  OR2_X1 U329 ( .A1(n305), .A2(n99), .ZN(out[78]) );
  AND2_X1 U329bar ( .A1(n305bar), .A2(n99bar), .ZN(outbar[78]) );
  OR2_X1 U330 ( .A1(n100), .A2(key[78]), .ZN(n306) );
  AND2_X1 U330bar ( .A1(n100bar), .A2(keybar[78]), .ZN(n306bar) );
  AND2_X1 U331 ( .A1(key[78]), .A2(n100), .ZN(n305) );
  OR2_X1 U331bar ( .A1(keybar[78]), .A2(n100bar), .ZN(n305bar) );
  OR2_X1 U332 ( .A1(n307), .A2(n101), .ZN(out[77]) );
  AND2_X1 U332bar ( .A1(n307bar), .A2(n101bar), .ZN(outbar[77]) );
  OR2_X1 U333 ( .A1(n102), .A2(key[77]), .ZN(n308) );
  AND2_X1 U333bar ( .A1(n102bar), .A2(keybar[77]), .ZN(n308bar) );
  AND2_X1 U334 ( .A1(key[77]), .A2(n102), .ZN(n307) );
  OR2_X1 U334bar ( .A1(keybar[77]), .A2(n102bar), .ZN(n307bar) );
  OR2_X1 U335 ( .A1(n309), .A2(n103), .ZN(out[76]) );
  AND2_X1 U335bar ( .A1(n309bar), .A2(n103bar), .ZN(outbar[76]) );
  OR2_X1 U336 ( .A1(n104), .A2(key[76]), .ZN(n310) );
  AND2_X1 U336bar ( .A1(n104bar), .A2(keybar[76]), .ZN(n310bar) );
  AND2_X1 U337 ( .A1(key[76]), .A2(n104), .ZN(n309) );
  OR2_X1 U337bar ( .A1(keybar[76]), .A2(n104bar), .ZN(n309bar) );
  OR2_X1 U338 ( .A1(n311), .A2(n105), .ZN(out[75]) );
  AND2_X1 U338bar ( .A1(n311bar), .A2(n105bar), .ZN(outbar[75]) );
  OR2_X1 U339 ( .A1(n106), .A2(key[75]), .ZN(n312) );
  AND2_X1 U339bar ( .A1(n106bar), .A2(keybar[75]), .ZN(n312bar) );
  AND2_X1 U340 ( .A1(key[75]), .A2(n106), .ZN(n311) );
  OR2_X1 U340bar ( .A1(keybar[75]), .A2(n106bar), .ZN(n311bar) );
  OR2_X1 U341 ( .A1(n313), .A2(n107), .ZN(out[74]) );
  AND2_X1 U341bar ( .A1(n313bar), .A2(n107bar), .ZN(outbar[74]) );
  OR2_X1 U342 ( .A1(n108), .A2(key[74]), .ZN(n314) );
  AND2_X1 U342bar ( .A1(n108bar), .A2(keybar[74]), .ZN(n314bar) );
  AND2_X1 U343 ( .A1(key[74]), .A2(n108), .ZN(n313) );
  OR2_X1 U343bar ( .A1(keybar[74]), .A2(n108bar), .ZN(n313bar) );
  OR2_X1 U344 ( .A1(n315), .A2(n109), .ZN(out[73]) );
  AND2_X1 U344bar ( .A1(n315bar), .A2(n109bar), .ZN(outbar[73]) );
  OR2_X1 U345 ( .A1(n110), .A2(key[73]), .ZN(n316) );
  AND2_X1 U345bar ( .A1(n110bar), .A2(keybar[73]), .ZN(n316bar) );
  AND2_X1 U346 ( .A1(key[73]), .A2(n110), .ZN(n315) );
  OR2_X1 U346bar ( .A1(keybar[73]), .A2(n110bar), .ZN(n315bar) );
  OR2_X1 U347 ( .A1(n317), .A2(n111), .ZN(out[72]) );
  AND2_X1 U347bar ( .A1(n317bar), .A2(n111bar), .ZN(outbar[72]) );
  OR2_X1 U348 ( .A1(n112), .A2(key[72]), .ZN(n318) );
  AND2_X1 U348bar ( .A1(n112bar), .A2(keybar[72]), .ZN(n318bar) );
  AND2_X1 U349 ( .A1(key[72]), .A2(n112), .ZN(n317) );
  OR2_X1 U349bar ( .A1(keybar[72]), .A2(n112bar), .ZN(n317bar) );
  OR2_X1 U350 ( .A1(n319), .A2(n113), .ZN(out[71]) );
  AND2_X1 U350bar ( .A1(n319bar), .A2(n113bar), .ZN(outbar[71]) );
  OR2_X1 U351 ( .A1(n114), .A2(key[71]), .ZN(n320) );
  AND2_X1 U351bar ( .A1(n114bar), .A2(keybar[71]), .ZN(n320bar) );
  AND2_X1 U352 ( .A1(key[71]), .A2(n114), .ZN(n319) );
  OR2_X1 U352bar ( .A1(keybar[71]), .A2(n114bar), .ZN(n319bar) );
  OR2_X1 U353 ( .A1(n321), .A2(n115), .ZN(out[70]) );
  AND2_X1 U353bar ( .A1(n321bar), .A2(n115bar), .ZN(outbar[70]) );
  OR2_X1 U354 ( .A1(n116), .A2(key[70]), .ZN(n322) );
  AND2_X1 U354bar ( .A1(n116bar), .A2(keybar[70]), .ZN(n322bar) );
  AND2_X1 U355 ( .A1(key[70]), .A2(n116), .ZN(n321) );
  OR2_X1 U355bar ( .A1(keybar[70]), .A2(n116bar), .ZN(n321bar) );
  OR2_X1 U356 ( .A1(n323), .A2(n243), .ZN(out[6]) );
  AND2_X1 U356bar ( .A1(n323bar), .A2(n243bar), .ZN(outbar[6]) );
  OR2_X1 U357 ( .A1(n244), .A2(key[6]), .ZN(n324) );
  AND2_X1 U357bar ( .A1(n244bar), .A2(keybar[6]), .ZN(n324bar) );
  AND2_X1 U358 ( .A1(key[6]), .A2(n244), .ZN(n323) );
  OR2_X1 U358bar ( .A1(keybar[6]), .A2(n244bar), .ZN(n323bar) );
  OR2_X1 U359 ( .A1(n325), .A2(n117), .ZN(out[69]) );
  AND2_X1 U359bar ( .A1(n325bar), .A2(n117bar), .ZN(outbar[69]) );
  OR2_X1 U360 ( .A1(n118), .A2(key[69]), .ZN(n326) );
  AND2_X1 U360bar ( .A1(n118bar), .A2(keybar[69]), .ZN(n326bar) );
  AND2_X1 U361 ( .A1(key[69]), .A2(n118), .ZN(n325) );
  OR2_X1 U361bar ( .A1(keybar[69]), .A2(n118bar), .ZN(n325bar) );
  OR2_X1 U362 ( .A1(n327), .A2(n119), .ZN(out[68]) );
  AND2_X1 U362bar ( .A1(n327bar), .A2(n119bar), .ZN(outbar[68]) );
  OR2_X1 U363 ( .A1(n120), .A2(key[68]), .ZN(n328) );
  AND2_X1 U363bar ( .A1(n120bar), .A2(keybar[68]), .ZN(n328bar) );
  AND2_X1 U364 ( .A1(key[68]), .A2(n120), .ZN(n327) );
  OR2_X1 U364bar ( .A1(keybar[68]), .A2(n120bar), .ZN(n327bar) );
  OR2_X1 U365 ( .A1(n329), .A2(n121), .ZN(out[67]) );
  AND2_X1 U365bar ( .A1(n329bar), .A2(n121bar), .ZN(outbar[67]) );
  OR2_X1 U366 ( .A1(n122), .A2(key[67]), .ZN(n330) );
  AND2_X1 U366bar ( .A1(n122bar), .A2(keybar[67]), .ZN(n330bar) );
  AND2_X1 U367 ( .A1(key[67]), .A2(n122), .ZN(n329) );
  OR2_X1 U367bar ( .A1(keybar[67]), .A2(n122bar), .ZN(n329bar) );
  OR2_X1 U368 ( .A1(n331), .A2(n123), .ZN(out[66]) );
  AND2_X1 U368bar ( .A1(n331bar), .A2(n123bar), .ZN(outbar[66]) );
  OR2_X1 U369 ( .A1(n124), .A2(key[66]), .ZN(n332) );
  AND2_X1 U369bar ( .A1(n124bar), .A2(keybar[66]), .ZN(n332bar) );
  AND2_X1 U370 ( .A1(key[66]), .A2(n124), .ZN(n331) );
  OR2_X1 U370bar ( .A1(keybar[66]), .A2(n124bar), .ZN(n331bar) );
  OR2_X1 U371 ( .A1(n333), .A2(n125), .ZN(out[65]) );
  AND2_X1 U371bar ( .A1(n333bar), .A2(n125bar), .ZN(outbar[65]) );
  OR2_X1 U372 ( .A1(n126), .A2(key[65]), .ZN(n334) );
  AND2_X1 U372bar ( .A1(n126bar), .A2(keybar[65]), .ZN(n334bar) );
  AND2_X1 U373 ( .A1(key[65]), .A2(n126), .ZN(n333) );
  OR2_X1 U373bar ( .A1(keybar[65]), .A2(n126bar), .ZN(n333bar) );
  OR2_X1 U374 ( .A1(n335), .A2(n127), .ZN(out[64]) );
  AND2_X1 U374bar ( .A1(n335bar), .A2(n127bar), .ZN(outbar[64]) );
  OR2_X1 U375 ( .A1(n128), .A2(key[64]), .ZN(n336) );
  AND2_X1 U375bar ( .A1(n128bar), .A2(keybar[64]), .ZN(n336bar) );
  AND2_X1 U376 ( .A1(key[64]), .A2(n128), .ZN(n335) );
  OR2_X1 U376bar ( .A1(keybar[64]), .A2(n128bar), .ZN(n335bar) );
  OR2_X1 U377 ( .A1(n337), .A2(n129), .ZN(out[63]) );
  AND2_X1 U377bar ( .A1(n337bar), .A2(n129bar), .ZN(outbar[63]) );
  OR2_X1 U378 ( .A1(n130), .A2(key[63]), .ZN(n338) );
  AND2_X1 U378bar ( .A1(n130bar), .A2(keybar[63]), .ZN(n338bar) );
  AND2_X1 U379 ( .A1(key[63]), .A2(n130), .ZN(n337) );
  OR2_X1 U379bar ( .A1(keybar[63]), .A2(n130bar), .ZN(n337bar) );
  OR2_X1 U380 ( .A1(n339), .A2(n131), .ZN(out[62]) );
  AND2_X1 U380bar ( .A1(n339bar), .A2(n131bar), .ZN(outbar[62]) );
  OR2_X1 U381 ( .A1(n132), .A2(key[62]), .ZN(n340) );
  AND2_X1 U381bar ( .A1(n132bar), .A2(keybar[62]), .ZN(n340bar) );
  AND2_X1 U382 ( .A1(key[62]), .A2(n132), .ZN(n339) );
  OR2_X1 U382bar ( .A1(keybar[62]), .A2(n132bar), .ZN(n339bar) );
  OR2_X1 U383 ( .A1(n341), .A2(n133), .ZN(out[61]) );
  AND2_X1 U383bar ( .A1(n341bar), .A2(n133bar), .ZN(outbar[61]) );
  OR2_X1 U384 ( .A1(n134), .A2(key[61]), .ZN(n342) );
  AND2_X1 U384bar ( .A1(n134bar), .A2(keybar[61]), .ZN(n342bar) );
  AND2_X1 U385 ( .A1(key[61]), .A2(n134), .ZN(n341) );
  OR2_X1 U385bar ( .A1(keybar[61]), .A2(n134bar), .ZN(n341bar) );
  OR2_X1 U386 ( .A1(n343), .A2(n135), .ZN(out[60]) );
  AND2_X1 U386bar ( .A1(n343bar), .A2(n135bar), .ZN(outbar[60]) );
  OR2_X1 U387 ( .A1(n136), .A2(key[60]), .ZN(n344) );
  AND2_X1 U387bar ( .A1(n136bar), .A2(keybar[60]), .ZN(n344bar) );
  AND2_X1 U388 ( .A1(key[60]), .A2(n136), .ZN(n343) );
  OR2_X1 U388bar ( .A1(keybar[60]), .A2(n136bar), .ZN(n343bar) );
  OR2_X1 U389 ( .A1(n345), .A2(n245), .ZN(out[5]) );
  AND2_X1 U389bar ( .A1(n345bar), .A2(n245bar), .ZN(outbar[5]) );
  OR2_X1 U390 ( .A1(n246), .A2(key[5]), .ZN(n346) );
  AND2_X1 U390bar ( .A1(n246bar), .A2(keybar[5]), .ZN(n346bar) );
  AND2_X1 U391 ( .A1(key[5]), .A2(n246), .ZN(n345) );
  OR2_X1 U391bar ( .A1(keybar[5]), .A2(n246bar), .ZN(n345bar) );
  OR2_X1 U392 ( .A1(n347), .A2(n137), .ZN(out[59]) );
  AND2_X1 U392bar ( .A1(n347bar), .A2(n137bar), .ZN(outbar[59]) );
  OR2_X1 U393 ( .A1(n138), .A2(key[59]), .ZN(n348) );
  AND2_X1 U393bar ( .A1(n138bar), .A2(keybar[59]), .ZN(n348bar) );
  AND2_X1 U394 ( .A1(key[59]), .A2(n138), .ZN(n347) );
  OR2_X1 U394bar ( .A1(keybar[59]), .A2(n138bar), .ZN(n347bar) );
  OR2_X1 U395 ( .A1(n349), .A2(n139), .ZN(out[58]) );
  AND2_X1 U395bar ( .A1(n349bar), .A2(n139bar), .ZN(outbar[58]) );
  OR2_X1 U396 ( .A1(n140), .A2(key[58]), .ZN(n350) );
  AND2_X1 U396bar ( .A1(n140bar), .A2(keybar[58]), .ZN(n350bar) );
  AND2_X1 U397 ( .A1(key[58]), .A2(n140), .ZN(n349) );
  OR2_X1 U397bar ( .A1(keybar[58]), .A2(n140bar), .ZN(n349bar) );
  OR2_X1 U398 ( .A1(n351), .A2(n141), .ZN(out[57]) );
  AND2_X1 U398bar ( .A1(n351bar), .A2(n141bar), .ZN(outbar[57]) );
  OR2_X1 U399 ( .A1(n142), .A2(key[57]), .ZN(n352) );
  AND2_X1 U399bar ( .A1(n142bar), .A2(keybar[57]), .ZN(n352bar) );
  AND2_X1 U400 ( .A1(key[57]), .A2(n142), .ZN(n351) );
  OR2_X1 U400bar ( .A1(keybar[57]), .A2(n142bar), .ZN(n351bar) );
  OR2_X1 U401 ( .A1(n353), .A2(n143), .ZN(out[56]) );
  AND2_X1 U401bar ( .A1(n353bar), .A2(n143bar), .ZN(outbar[56]) );
  OR2_X1 U402 ( .A1(n144), .A2(key[56]), .ZN(n354) );
  AND2_X1 U402bar ( .A1(n144bar), .A2(keybar[56]), .ZN(n354bar) );
  AND2_X1 U403 ( .A1(key[56]), .A2(n144), .ZN(n353) );
  OR2_X1 U403bar ( .A1(keybar[56]), .A2(n144bar), .ZN(n353bar) );
  OR2_X1 U404 ( .A1(n355), .A2(n145), .ZN(out[55]) );
  AND2_X1 U404bar ( .A1(n355bar), .A2(n145bar), .ZN(outbar[55]) );
  OR2_X1 U405 ( .A1(n146), .A2(key[55]), .ZN(n356) );
  AND2_X1 U405bar ( .A1(n146bar), .A2(keybar[55]), .ZN(n356bar) );
  AND2_X1 U406 ( .A1(key[55]), .A2(n146), .ZN(n355) );
  OR2_X1 U406bar ( .A1(keybar[55]), .A2(n146bar), .ZN(n355bar) );
  OR2_X1 U407 ( .A1(n357), .A2(n147), .ZN(out[54]) );
  AND2_X1 U407bar ( .A1(n357bar), .A2(n147bar), .ZN(outbar[54]) );
  OR2_X1 U408 ( .A1(n148), .A2(key[54]), .ZN(n358) );
  AND2_X1 U408bar ( .A1(n148bar), .A2(keybar[54]), .ZN(n358bar) );
  AND2_X1 U409 ( .A1(key[54]), .A2(n148), .ZN(n357) );
  OR2_X1 U409bar ( .A1(keybar[54]), .A2(n148bar), .ZN(n357bar) );
  OR2_X1 U410 ( .A1(n359), .A2(n149), .ZN(out[53]) );
  AND2_X1 U410bar ( .A1(n359bar), .A2(n149bar), .ZN(outbar[53]) );
  OR2_X1 U411 ( .A1(n150), .A2(key[53]), .ZN(n360) );
  AND2_X1 U411bar ( .A1(n150bar), .A2(keybar[53]), .ZN(n360bar) );
  AND2_X1 U412 ( .A1(key[53]), .A2(n150), .ZN(n359) );
  OR2_X1 U412bar ( .A1(keybar[53]), .A2(n150bar), .ZN(n359bar) );
  OR2_X1 U413 ( .A1(n361), .A2(n151), .ZN(out[52]) );
  AND2_X1 U413bar ( .A1(n361bar), .A2(n151bar), .ZN(outbar[52]) );
  OR2_X1 U414 ( .A1(n152), .A2(key[52]), .ZN(n362) );
  AND2_X1 U414bar ( .A1(n152bar), .A2(keybar[52]), .ZN(n362bar) );
  AND2_X1 U415 ( .A1(key[52]), .A2(n152), .ZN(n361) );
  OR2_X1 U415bar ( .A1(keybar[52]), .A2(n152bar), .ZN(n361bar) );
  OR2_X1 U416 ( .A1(n363), .A2(n153), .ZN(out[51]) );
  AND2_X1 U416bar ( .A1(n363bar), .A2(n153bar), .ZN(outbar[51]) );
  OR2_X1 U417 ( .A1(n154), .A2(key[51]), .ZN(n364) );
  AND2_X1 U417bar ( .A1(n154bar), .A2(keybar[51]), .ZN(n364bar) );
  AND2_X1 U418 ( .A1(key[51]), .A2(n154), .ZN(n363) );
  OR2_X1 U418bar ( .A1(keybar[51]), .A2(n154bar), .ZN(n363bar) );
  OR2_X1 U419 ( .A1(n365), .A2(n155), .ZN(out[50]) );
  AND2_X1 U419bar ( .A1(n365bar), .A2(n155bar), .ZN(outbar[50]) );
  OR2_X1 U420 ( .A1(n156), .A2(key[50]), .ZN(n366) );
  AND2_X1 U420bar ( .A1(n156bar), .A2(keybar[50]), .ZN(n366bar) );
  AND2_X1 U421 ( .A1(key[50]), .A2(n156), .ZN(n365) );
  OR2_X1 U421bar ( .A1(keybar[50]), .A2(n156bar), .ZN(n365bar) );
  OR2_X1 U422 ( .A1(n367), .A2(n247), .ZN(out[4]) );
  AND2_X1 U422bar ( .A1(n367bar), .A2(n247bar), .ZN(outbar[4]) );
  OR2_X1 U423 ( .A1(n248), .A2(key[4]), .ZN(n368) );
  AND2_X1 U423bar ( .A1(n248bar), .A2(keybar[4]), .ZN(n368bar) );
  AND2_X1 U424 ( .A1(key[4]), .A2(n248), .ZN(n367) );
  OR2_X1 U424bar ( .A1(keybar[4]), .A2(n248bar), .ZN(n367bar) );
  OR2_X1 U425 ( .A1(n369), .A2(n157), .ZN(out[49]) );
  AND2_X1 U425bar ( .A1(n369bar), .A2(n157bar), .ZN(outbar[49]) );
  OR2_X1 U426 ( .A1(n158), .A2(key[49]), .ZN(n370) );
  AND2_X1 U426bar ( .A1(n158bar), .A2(keybar[49]), .ZN(n370bar) );
  AND2_X1 U427 ( .A1(key[49]), .A2(n158), .ZN(n369) );
  OR2_X1 U427bar ( .A1(keybar[49]), .A2(n158bar), .ZN(n369bar) );
  OR2_X1 U428 ( .A1(n371), .A2(n159), .ZN(out[48]) );
  AND2_X1 U428bar ( .A1(n371bar), .A2(n159bar), .ZN(outbar[48]) );
  OR2_X1 U429 ( .A1(n160), .A2(key[48]), .ZN(n372) );
  AND2_X1 U429bar ( .A1(n160bar), .A2(keybar[48]), .ZN(n372bar) );
  AND2_X1 U430 ( .A1(key[48]), .A2(n160), .ZN(n371) );
  OR2_X1 U430bar ( .A1(keybar[48]), .A2(n160bar), .ZN(n371bar) );
  OR2_X1 U431 ( .A1(n373), .A2(n161), .ZN(out[47]) );
  AND2_X1 U431bar ( .A1(n373bar), .A2(n161bar), .ZN(outbar[47]) );
  OR2_X1 U432 ( .A1(n162), .A2(key[47]), .ZN(n374) );
  AND2_X1 U432bar ( .A1(n162bar), .A2(keybar[47]), .ZN(n374bar) );
  AND2_X1 U433 ( .A1(key[47]), .A2(n162), .ZN(n373) );
  OR2_X1 U433bar ( .A1(keybar[47]), .A2(n162bar), .ZN(n373bar) );
  OR2_X1 U434 ( .A1(n375), .A2(n163), .ZN(out[46]) );
  AND2_X1 U434bar ( .A1(n375bar), .A2(n163bar), .ZN(outbar[46]) );
  OR2_X1 U435 ( .A1(n164), .A2(key[46]), .ZN(n376) );
  AND2_X1 U435bar ( .A1(n164bar), .A2(keybar[46]), .ZN(n376bar) );
  AND2_X1 U436 ( .A1(key[46]), .A2(n164), .ZN(n375) );
  OR2_X1 U436bar ( .A1(keybar[46]), .A2(n164bar), .ZN(n375bar) );
  OR2_X1 U437 ( .A1(n377), .A2(n165), .ZN(out[45]) );
  AND2_X1 U437bar ( .A1(n377bar), .A2(n165bar), .ZN(outbar[45]) );
  OR2_X1 U438 ( .A1(n166), .A2(key[45]), .ZN(n378) );
  AND2_X1 U438bar ( .A1(n166bar), .A2(keybar[45]), .ZN(n378bar) );
  AND2_X1 U439 ( .A1(key[45]), .A2(n166), .ZN(n377) );
  OR2_X1 U439bar ( .A1(keybar[45]), .A2(n166bar), .ZN(n377bar) );
  OR2_X1 U440 ( .A1(n379), .A2(n167), .ZN(out[44]) );
  AND2_X1 U440bar ( .A1(n379bar), .A2(n167bar), .ZN(outbar[44]) );
  OR2_X1 U441 ( .A1(n168), .A2(key[44]), .ZN(n380) );
  AND2_X1 U441bar ( .A1(n168bar), .A2(keybar[44]), .ZN(n380bar) );
  AND2_X1 U442 ( .A1(key[44]), .A2(n168), .ZN(n379) );
  OR2_X1 U442bar ( .A1(keybar[44]), .A2(n168bar), .ZN(n379bar) );
  OR2_X1 U443 ( .A1(n381), .A2(n169), .ZN(out[43]) );
  AND2_X1 U443bar ( .A1(n381bar), .A2(n169bar), .ZN(outbar[43]) );
  OR2_X1 U444 ( .A1(n170), .A2(key[43]), .ZN(n382) );
  AND2_X1 U444bar ( .A1(n170bar), .A2(keybar[43]), .ZN(n382bar) );
  AND2_X1 U445 ( .A1(key[43]), .A2(n170), .ZN(n381) );
  OR2_X1 U445bar ( .A1(keybar[43]), .A2(n170bar), .ZN(n381bar) );
  OR2_X1 U446 ( .A1(n383), .A2(n171), .ZN(out[42]) );
  AND2_X1 U446bar ( .A1(n383bar), .A2(n171bar), .ZN(outbar[42]) );
  OR2_X1 U447 ( .A1(n172), .A2(key[42]), .ZN(n384) );
  AND2_X1 U447bar ( .A1(n172bar), .A2(keybar[42]), .ZN(n384bar) );
  AND2_X1 U448 ( .A1(key[42]), .A2(n172), .ZN(n383) );
  OR2_X1 U448bar ( .A1(keybar[42]), .A2(n172bar), .ZN(n383bar) );
  OR2_X1 U449 ( .A1(n385), .A2(n173), .ZN(out[41]) );
  AND2_X1 U449bar ( .A1(n385bar), .A2(n173bar), .ZN(outbar[41]) );
  OR2_X1 U450 ( .A1(n174), .A2(key[41]), .ZN(n386) );
  AND2_X1 U450bar ( .A1(n174bar), .A2(keybar[41]), .ZN(n386bar) );
  AND2_X1 U451 ( .A1(key[41]), .A2(n174), .ZN(n385) );
  OR2_X1 U451bar ( .A1(keybar[41]), .A2(n174bar), .ZN(n385bar) );
  OR2_X1 U452 ( .A1(n387), .A2(n175), .ZN(out[40]) );
  AND2_X1 U452bar ( .A1(n387bar), .A2(n175bar), .ZN(outbar[40]) );
  OR2_X1 U453 ( .A1(n176), .A2(key[40]), .ZN(n388) );
  AND2_X1 U453bar ( .A1(n176bar), .A2(keybar[40]), .ZN(n388bar) );
  AND2_X1 U454 ( .A1(key[40]), .A2(n176), .ZN(n387) );
  OR2_X1 U454bar ( .A1(keybar[40]), .A2(n176bar), .ZN(n387bar) );
  OR2_X1 U455 ( .A1(n389), .A2(n249), .ZN(out[3]) );
  AND2_X1 U455bar ( .A1(n389bar), .A2(n249bar), .ZN(outbar[3]) );
  OR2_X1 U456 ( .A1(n250), .A2(key[3]), .ZN(n390) );
  AND2_X1 U456bar ( .A1(n250bar), .A2(keybar[3]), .ZN(n390bar) );
  AND2_X1 U457 ( .A1(key[3]), .A2(n250), .ZN(n389) );
  OR2_X1 U457bar ( .A1(keybar[3]), .A2(n250bar), .ZN(n389bar) );
  OR2_X1 U458 ( .A1(n391), .A2(n177), .ZN(out[39]) );
  AND2_X1 U458bar ( .A1(n391bar), .A2(n177bar), .ZN(outbar[39]) );
  OR2_X1 U459 ( .A1(n178), .A2(key[39]), .ZN(n392) );
  AND2_X1 U459bar ( .A1(n178bar), .A2(keybar[39]), .ZN(n392bar) );
  AND2_X1 U460 ( .A1(key[39]), .A2(n178), .ZN(n391) );
  OR2_X1 U460bar ( .A1(keybar[39]), .A2(n178bar), .ZN(n391bar) );
  OR2_X1 U461 ( .A1(n393), .A2(n179), .ZN(out[38]) );
  AND2_X1 U461bar ( .A1(n393bar), .A2(n179bar), .ZN(outbar[38]) );
  OR2_X1 U462 ( .A1(n180), .A2(key[38]), .ZN(n394) );
  AND2_X1 U462bar ( .A1(n180bar), .A2(keybar[38]), .ZN(n394bar) );
  AND2_X1 U463 ( .A1(key[38]), .A2(n180), .ZN(n393) );
  OR2_X1 U463bar ( .A1(keybar[38]), .A2(n180bar), .ZN(n393bar) );
  OR2_X1 U464 ( .A1(n395), .A2(n181), .ZN(out[37]) );
  AND2_X1 U464bar ( .A1(n395bar), .A2(n181bar), .ZN(outbar[37]) );
  OR2_X1 U465 ( .A1(n182), .A2(key[37]), .ZN(n396) );
  AND2_X1 U465bar ( .A1(n182bar), .A2(keybar[37]), .ZN(n396bar) );
  AND2_X1 U466 ( .A1(key[37]), .A2(n182), .ZN(n395) );
  OR2_X1 U466bar ( .A1(keybar[37]), .A2(n182bar), .ZN(n395bar) );
  OR2_X1 U467 ( .A1(n397), .A2(n183), .ZN(out[36]) );
  AND2_X1 U467bar ( .A1(n397bar), .A2(n183bar), .ZN(outbar[36]) );
  OR2_X1 U468 ( .A1(n184), .A2(key[36]), .ZN(n398) );
  AND2_X1 U468bar ( .A1(n184bar), .A2(keybar[36]), .ZN(n398bar) );
  AND2_X1 U469 ( .A1(key[36]), .A2(n184), .ZN(n397) );
  OR2_X1 U469bar ( .A1(keybar[36]), .A2(n184bar), .ZN(n397bar) );
  OR2_X1 U470 ( .A1(n399), .A2(n185), .ZN(out[35]) );
  AND2_X1 U470bar ( .A1(n399bar), .A2(n185bar), .ZN(outbar[35]) );
  OR2_X1 U471 ( .A1(n186), .A2(key[35]), .ZN(n400) );
  AND2_X1 U471bar ( .A1(n186bar), .A2(keybar[35]), .ZN(n400bar) );
  AND2_X1 U472 ( .A1(key[35]), .A2(n186), .ZN(n399) );
  OR2_X1 U472bar ( .A1(keybar[35]), .A2(n186bar), .ZN(n399bar) );
  OR2_X1 U473 ( .A1(n401), .A2(n187), .ZN(out[34]) );
  AND2_X1 U473bar ( .A1(n401bar), .A2(n187bar), .ZN(outbar[34]) );
  OR2_X1 U474 ( .A1(n188), .A2(key[34]), .ZN(n402) );
  AND2_X1 U474bar ( .A1(n188bar), .A2(keybar[34]), .ZN(n402bar) );
  AND2_X1 U475 ( .A1(key[34]), .A2(n188), .ZN(n401) );
  OR2_X1 U475bar ( .A1(keybar[34]), .A2(n188bar), .ZN(n401bar) );
  OR2_X1 U476 ( .A1(n403), .A2(n189), .ZN(out[33]) );
  AND2_X1 U476bar ( .A1(n403bar), .A2(n189bar), .ZN(outbar[33]) );
  OR2_X1 U477 ( .A1(n190), .A2(key[33]), .ZN(n404) );
  AND2_X1 U477bar ( .A1(n190bar), .A2(keybar[33]), .ZN(n404bar) );
  AND2_X1 U478 ( .A1(key[33]), .A2(n190), .ZN(n403) );
  OR2_X1 U478bar ( .A1(keybar[33]), .A2(n190bar), .ZN(n403bar) );
  OR2_X1 U479 ( .A1(n405), .A2(n191), .ZN(out[32]) );
  AND2_X1 U479bar ( .A1(n405bar), .A2(n191bar), .ZN(outbar[32]) );
  OR2_X1 U480 ( .A1(n192), .A2(key[32]), .ZN(n406) );
  AND2_X1 U480bar ( .A1(n192bar), .A2(keybar[32]), .ZN(n406bar) );
  AND2_X1 U481 ( .A1(key[32]), .A2(n192), .ZN(n405) );
  OR2_X1 U481bar ( .A1(keybar[32]), .A2(n192bar), .ZN(n405bar) );
  OR2_X1 U482 ( .A1(n407), .A2(n193), .ZN(out[31]) );
  AND2_X1 U482bar ( .A1(n407bar), .A2(n193bar), .ZN(outbar[31]) );
  OR2_X1 U483 ( .A1(n194), .A2(key[31]), .ZN(n408) );
  AND2_X1 U483bar ( .A1(n194bar), .A2(keybar[31]), .ZN(n408bar) );
  AND2_X1 U484 ( .A1(key[31]), .A2(n194), .ZN(n407) );
  OR2_X1 U484bar ( .A1(keybar[31]), .A2(n194bar), .ZN(n407bar) );
  OR2_X1 U485 ( .A1(n409), .A2(n195), .ZN(out[30]) );
  AND2_X1 U485bar ( .A1(n409bar), .A2(n195bar), .ZN(outbar[30]) );
  OR2_X1 U486 ( .A1(n196), .A2(key[30]), .ZN(n410) );
  AND2_X1 U486bar ( .A1(n196bar), .A2(keybar[30]), .ZN(n410bar) );
  AND2_X1 U487 ( .A1(key[30]), .A2(n196), .ZN(n409) );
  OR2_X1 U487bar ( .A1(keybar[30]), .A2(n196bar), .ZN(n409bar) );
  OR2_X1 U488 ( .A1(n411), .A2(n251), .ZN(out[2]) );
  AND2_X1 U488bar ( .A1(n411bar), .A2(n251bar), .ZN(outbar[2]) );
  OR2_X1 U489 ( .A1(n252), .A2(key[2]), .ZN(n412) );
  AND2_X1 U489bar ( .A1(n252bar), .A2(keybar[2]), .ZN(n412bar) );
  AND2_X1 U490 ( .A1(key[2]), .A2(n252), .ZN(n411) );
  OR2_X1 U490bar ( .A1(keybar[2]), .A2(n252bar), .ZN(n411bar) );
  OR2_X1 U491 ( .A1(n413), .A2(n197), .ZN(out[29]) );
  AND2_X1 U491bar ( .A1(n413bar), .A2(n197bar), .ZN(outbar[29]) );
  OR2_X1 U492 ( .A1(n198), .A2(key[29]), .ZN(n414) );
  AND2_X1 U492bar ( .A1(n198bar), .A2(keybar[29]), .ZN(n414bar) );
  AND2_X1 U493 ( .A1(key[29]), .A2(n198), .ZN(n413) );
  OR2_X1 U493bar ( .A1(keybar[29]), .A2(n198bar), .ZN(n413bar) );
  OR2_X1 U494 ( .A1(n415), .A2(n199), .ZN(out[28]) );
  AND2_X1 U494bar ( .A1(n415bar), .A2(n199bar), .ZN(outbar[28]) );
  OR2_X1 U495 ( .A1(n200), .A2(key[28]), .ZN(n416) );
  AND2_X1 U495bar ( .A1(n200bar), .A2(keybar[28]), .ZN(n416bar) );
  AND2_X1 U496 ( .A1(key[28]), .A2(n200), .ZN(n415) );
  OR2_X1 U496bar ( .A1(keybar[28]), .A2(n200bar), .ZN(n415bar) );
  OR2_X1 U497 ( .A1(n417), .A2(n201), .ZN(out[27]) );
  AND2_X1 U497bar ( .A1(n417bar), .A2(n201bar), .ZN(outbar[27]) );
  OR2_X1 U498 ( .A1(n202), .A2(key[27]), .ZN(n418) );
  AND2_X1 U498bar ( .A1(n202bar), .A2(keybar[27]), .ZN(n418bar) );
  AND2_X1 U499 ( .A1(key[27]), .A2(n202), .ZN(n417) );
  OR2_X1 U499bar ( .A1(keybar[27]), .A2(n202bar), .ZN(n417bar) );
  OR2_X1 U500 ( .A1(n419), .A2(n203), .ZN(out[26]) );
  AND2_X1 U500bar ( .A1(n419bar), .A2(n203bar), .ZN(outbar[26]) );
  OR2_X1 U501 ( .A1(n204), .A2(key[26]), .ZN(n420) );
  AND2_X1 U501bar ( .A1(n204bar), .A2(keybar[26]), .ZN(n420bar) );
  AND2_X1 U502 ( .A1(key[26]), .A2(n204), .ZN(n419) );
  OR2_X1 U502bar ( .A1(keybar[26]), .A2(n204bar), .ZN(n419bar) );
  OR2_X1 U503 ( .A1(n421), .A2(n205), .ZN(out[25]) );
  AND2_X1 U503bar ( .A1(n421bar), .A2(n205bar), .ZN(outbar[25]) );
  OR2_X1 U504 ( .A1(n206), .A2(key[25]), .ZN(n422) );
  AND2_X1 U504bar ( .A1(n206bar), .A2(keybar[25]), .ZN(n422bar) );
  AND2_X1 U505 ( .A1(key[25]), .A2(n206), .ZN(n421) );
  OR2_X1 U505bar ( .A1(keybar[25]), .A2(n206bar), .ZN(n421bar) );
  OR2_X1 U506 ( .A1(n423), .A2(n207), .ZN(out[24]) );
  AND2_X1 U506bar ( .A1(n423bar), .A2(n207bar), .ZN(outbar[24]) );
  OR2_X1 U507 ( .A1(n208), .A2(key[24]), .ZN(n424) );
  AND2_X1 U507bar ( .A1(n208bar), .A2(keybar[24]), .ZN(n424bar) );
  AND2_X1 U508 ( .A1(key[24]), .A2(n208), .ZN(n423) );
  OR2_X1 U508bar ( .A1(keybar[24]), .A2(n208bar), .ZN(n423bar) );
  OR2_X1 U509 ( .A1(n425), .A2(n209), .ZN(out[23]) );
  AND2_X1 U509bar ( .A1(n425bar), .A2(n209bar), .ZN(outbar[23]) );
  OR2_X1 U510 ( .A1(n210), .A2(key[23]), .ZN(n426) );
  AND2_X1 U510bar ( .A1(n210bar), .A2(keybar[23]), .ZN(n426bar) );
  AND2_X1 U511 ( .A1(key[23]), .A2(n210), .ZN(n425) );
  OR2_X1 U511bar ( .A1(keybar[23]), .A2(n210bar), .ZN(n425bar) );
  OR2_X1 U512 ( .A1(n427), .A2(n211), .ZN(out[22]) );
  AND2_X1 U512bar ( .A1(n427bar), .A2(n211bar), .ZN(outbar[22]) );
  OR2_X1 U513 ( .A1(n212), .A2(key[22]), .ZN(n428) );
  AND2_X1 U513bar ( .A1(n212bar), .A2(keybar[22]), .ZN(n428bar) );
  AND2_X1 U514 ( .A1(key[22]), .A2(n212), .ZN(n427) );
  OR2_X1 U514bar ( .A1(keybar[22]), .A2(n212bar), .ZN(n427bar) );
  OR2_X1 U515 ( .A1(n429), .A2(n213), .ZN(out[21]) );
  AND2_X1 U515bar ( .A1(n429bar), .A2(n213bar), .ZN(outbar[21]) );
  OR2_X1 U516 ( .A1(n214), .A2(key[21]), .ZN(n430) );
  AND2_X1 U516bar ( .A1(n214bar), .A2(keybar[21]), .ZN(n430bar) );
  AND2_X1 U517 ( .A1(key[21]), .A2(n214), .ZN(n429) );
  OR2_X1 U517bar ( .A1(keybar[21]), .A2(n214bar), .ZN(n429bar) );
  OR2_X1 U518 ( .A1(n431), .A2(n215), .ZN(out[20]) );
  AND2_X1 U518bar ( .A1(n431bar), .A2(n215bar), .ZN(outbar[20]) );
  OR2_X1 U519 ( .A1(n216), .A2(key[20]), .ZN(n432) );
  AND2_X1 U519bar ( .A1(n216bar), .A2(keybar[20]), .ZN(n432bar) );
  AND2_X1 U520 ( .A1(key[20]), .A2(n216), .ZN(n431) );
  OR2_X1 U520bar ( .A1(keybar[20]), .A2(n216bar), .ZN(n431bar) );
  OR2_X1 U521 ( .A1(n433), .A2(n253), .ZN(out[1]) );
  AND2_X1 U521bar ( .A1(n433bar), .A2(n253bar), .ZN(outbar[1]) );
  OR2_X1 U522 ( .A1(n254), .A2(key[1]), .ZN(n434) );
  AND2_X1 U522bar ( .A1(n254bar), .A2(keybar[1]), .ZN(n434bar) );
  AND2_X1 U523 ( .A1(key[1]), .A2(n254), .ZN(n433) );
  OR2_X1 U523bar ( .A1(keybar[1]), .A2(n254bar), .ZN(n433bar) );
  OR2_X1 U524 ( .A1(n435), .A2(n217), .ZN(out[19]) );
  AND2_X1 U524bar ( .A1(n435bar), .A2(n217bar), .ZN(outbar[19]) );
  OR2_X1 U525 ( .A1(n218), .A2(key[19]), .ZN(n436) );
  AND2_X1 U525bar ( .A1(n218bar), .A2(keybar[19]), .ZN(n436bar) );
  AND2_X1 U526 ( .A1(key[19]), .A2(n218), .ZN(n435) );
  OR2_X1 U526bar ( .A1(keybar[19]), .A2(n218bar), .ZN(n435bar) );
  OR2_X1 U527 ( .A1(n437), .A2(n219), .ZN(out[18]) );
  AND2_X1 U527bar ( .A1(n437bar), .A2(n219bar), .ZN(outbar[18]) );
  OR2_X1 U528 ( .A1(n220), .A2(key[18]), .ZN(n438) );
  AND2_X1 U528bar ( .A1(n220bar), .A2(keybar[18]), .ZN(n438bar) );
  AND2_X1 U529 ( .A1(key[18]), .A2(n220), .ZN(n437) );
  OR2_X1 U529bar ( .A1(keybar[18]), .A2(n220bar), .ZN(n437bar) );
  OR2_X1 U530 ( .A1(n439), .A2(n221), .ZN(out[17]) );
  AND2_X1 U530bar ( .A1(n439bar), .A2(n221bar), .ZN(outbar[17]) );
  OR2_X1 U531 ( .A1(n222), .A2(key[17]), .ZN(n440) );
  AND2_X1 U531bar ( .A1(n222bar), .A2(keybar[17]), .ZN(n440bar) );
  AND2_X1 U532 ( .A1(key[17]), .A2(n222), .ZN(n439) );
  OR2_X1 U532bar ( .A1(keybar[17]), .A2(n222bar), .ZN(n439bar) );
  OR2_X1 U533 ( .A1(n441), .A2(n223), .ZN(out[16]) );
  AND2_X1 U533bar ( .A1(n441bar), .A2(n223bar), .ZN(outbar[16]) );
  OR2_X1 U534 ( .A1(n224), .A2(key[16]), .ZN(n442) );
  AND2_X1 U534bar ( .A1(n224bar), .A2(keybar[16]), .ZN(n442bar) );
  AND2_X1 U535 ( .A1(key[16]), .A2(n224), .ZN(n441) );
  OR2_X1 U535bar ( .A1(keybar[16]), .A2(n224bar), .ZN(n441bar) );
  OR2_X1 U536 ( .A1(n443), .A2(n225), .ZN(out[15]) );
  AND2_X1 U536bar ( .A1(n443bar), .A2(n225bar), .ZN(outbar[15]) );
  OR2_X1 U537 ( .A1(n226), .A2(key[15]), .ZN(n444) );
  AND2_X1 U537bar ( .A1(n226bar), .A2(keybar[15]), .ZN(n444bar) );
  AND2_X1 U538 ( .A1(key[15]), .A2(n226), .ZN(n443) );
  OR2_X1 U538bar ( .A1(keybar[15]), .A2(n226bar), .ZN(n443bar) );
  OR2_X1 U539 ( .A1(n445), .A2(n227), .ZN(out[14]) );
  AND2_X1 U539bar ( .A1(n445bar), .A2(n227bar), .ZN(outbar[14]) );
  OR2_X1 U540 ( .A1(n228), .A2(key[14]), .ZN(n446) );
  AND2_X1 U540bar ( .A1(n228bar), .A2(keybar[14]), .ZN(n446bar) );
  AND2_X1 U541 ( .A1(key[14]), .A2(n228), .ZN(n445) );
  OR2_X1 U541bar ( .A1(keybar[14]), .A2(n228bar), .ZN(n445bar) );
  OR2_X1 U542 ( .A1(n447), .A2(n229), .ZN(out[13]) );
  AND2_X1 U542bar ( .A1(n447bar), .A2(n229bar), .ZN(outbar[13]) );
  OR2_X1 U543 ( .A1(n230), .A2(key[13]), .ZN(n448) );
  AND2_X1 U543bar ( .A1(n230bar), .A2(keybar[13]), .ZN(n448bar) );
  AND2_X1 U544 ( .A1(key[13]), .A2(n230), .ZN(n447) );
  OR2_X1 U544bar ( .A1(keybar[13]), .A2(n230bar), .ZN(n447bar) );
  OR2_X1 U545 ( .A1(n449), .A2(n231), .ZN(out[12]) );
  AND2_X1 U545bar ( .A1(n449bar), .A2(n231bar), .ZN(outbar[12]) );
  OR2_X1 U546 ( .A1(n232), .A2(key[12]), .ZN(n450) );
  AND2_X1 U546bar ( .A1(n232bar), .A2(keybar[12]), .ZN(n450bar) );
  AND2_X1 U547 ( .A1(key[12]), .A2(n232), .ZN(n449) );
  OR2_X1 U547bar ( .A1(keybar[12]), .A2(n232bar), .ZN(n449bar) );
  OR2_X1 U548 ( .A1(n451), .A2(n1), .ZN(out[127]) );
  AND2_X1 U548bar ( .A1(n451bar), .A2(n1bar), .ZN(outbar[127]) );
  OR2_X1 U549 ( .A1(n2), .A2(key[127]), .ZN(n452) );
  AND2_X1 U549bar ( .A1(n2bar), .A2(keybar[127]), .ZN(n452bar) );
  AND2_X1 U550 ( .A1(key[127]), .A2(n2), .ZN(n451) );
  OR2_X1 U550bar ( .A1(keybar[127]), .A2(n2bar), .ZN(n451bar) );
  OR2_X1 U551 ( .A1(n453), .A2(n3), .ZN(out[126]) );
  AND2_X1 U551bar ( .A1(n453bar), .A2(n3bar), .ZN(outbar[126]) );
  OR2_X1 U552 ( .A1(n4), .A2(key[126]), .ZN(n454) );
  AND2_X1 U552bar ( .A1(n4bar), .A2(keybar[126]), .ZN(n454bar) );
  AND2_X1 U553 ( .A1(key[126]), .A2(n4), .ZN(n453) );
  OR2_X1 U553bar ( .A1(keybar[126]), .A2(n4bar), .ZN(n453bar) );
  OR2_X1 U554 ( .A1(n455), .A2(n5), .ZN(out[125]) );
  AND2_X1 U554bar ( .A1(n455bar), .A2(n5bar), .ZN(outbar[125]) );
  OR2_X1 U555 ( .A1(n6), .A2(key[125]), .ZN(n456) );
  AND2_X1 U555bar ( .A1(n6bar), .A2(keybar[125]), .ZN(n456bar) );
  AND2_X1 U556 ( .A1(key[125]), .A2(n6), .ZN(n455) );
  OR2_X1 U556bar ( .A1(keybar[125]), .A2(n6bar), .ZN(n455bar) );
  OR2_X1 U557 ( .A1(n457), .A2(n7), .ZN(out[124]) );
  AND2_X1 U557bar ( .A1(n457bar), .A2(n7bar), .ZN(outbar[124]) );
  OR2_X1 U558 ( .A1(n8), .A2(key[124]), .ZN(n458) );
  AND2_X1 U558bar ( .A1(n8bar), .A2(keybar[124]), .ZN(n458bar) );
  AND2_X1 U559 ( .A1(key[124]), .A2(n8), .ZN(n457) );
  OR2_X1 U559bar ( .A1(keybar[124]), .A2(n8bar), .ZN(n457bar) );
  OR2_X1 U560 ( .A1(n459), .A2(n9), .ZN(out[123]) );
  AND2_X1 U560bar ( .A1(n459bar), .A2(n9bar), .ZN(outbar[123]) );
  OR2_X1 U561 ( .A1(n10), .A2(key[123]), .ZN(n460) );
  AND2_X1 U561bar ( .A1(n10bar), .A2(keybar[123]), .ZN(n460bar) );
  AND2_X1 U562 ( .A1(key[123]), .A2(n10), .ZN(n459) );
  OR2_X1 U562bar ( .A1(keybar[123]), .A2(n10bar), .ZN(n459bar) );
  OR2_X1 U563 ( .A1(n461), .A2(n11), .ZN(out[122]) );
  AND2_X1 U563bar ( .A1(n461bar), .A2(n11bar), .ZN(outbar[122]) );
  OR2_X1 U564 ( .A1(n12), .A2(key[122]), .ZN(n462) );
  AND2_X1 U564bar ( .A1(n12bar), .A2(keybar[122]), .ZN(n462bar) );
  AND2_X1 U565 ( .A1(key[122]), .A2(n12), .ZN(n461) );
  OR2_X1 U565bar ( .A1(keybar[122]), .A2(n12bar), .ZN(n461bar) );
  OR2_X1 U566 ( .A1(n463), .A2(n13), .ZN(out[121]) );
  AND2_X1 U566bar ( .A1(n463bar), .A2(n13bar), .ZN(outbar[121]) );
  OR2_X1 U567 ( .A1(n14), .A2(key[121]), .ZN(n464) );
  AND2_X1 U567bar ( .A1(n14bar), .A2(keybar[121]), .ZN(n464bar) );
  AND2_X1 U568 ( .A1(key[121]), .A2(n14), .ZN(n463) );
  OR2_X1 U568bar ( .A1(keybar[121]), .A2(n14bar), .ZN(n463bar) );
  OR2_X1 U569 ( .A1(n465), .A2(n15), .ZN(out[120]) );
  AND2_X1 U569bar ( .A1(n465bar), .A2(n15bar), .ZN(outbar[120]) );
  OR2_X1 U570 ( .A1(n16), .A2(key[120]), .ZN(n466) );
  AND2_X1 U570bar ( .A1(n16bar), .A2(keybar[120]), .ZN(n466bar) );
  AND2_X1 U571 ( .A1(key[120]), .A2(n16), .ZN(n465) );
  OR2_X1 U571bar ( .A1(keybar[120]), .A2(n16bar), .ZN(n465bar) );
  OR2_X1 U572 ( .A1(n467), .A2(n233), .ZN(out[11]) );
  AND2_X1 U572bar ( .A1(n467bar), .A2(n233bar), .ZN(outbar[11]) );
  OR2_X1 U573 ( .A1(n234), .A2(key[11]), .ZN(n468) );
  AND2_X1 U573bar ( .A1(n234bar), .A2(keybar[11]), .ZN(n468bar) );
  AND2_X1 U574 ( .A1(key[11]), .A2(n234), .ZN(n467) );
  OR2_X1 U574bar ( .A1(keybar[11]), .A2(n234bar), .ZN(n467bar) );
  OR2_X1 U575 ( .A1(n469), .A2(n17), .ZN(out[119]) );
  AND2_X1 U575bar ( .A1(n469bar), .A2(n17bar), .ZN(outbar[119]) );
  OR2_X1 U576 ( .A1(n18), .A2(key[119]), .ZN(n470) );
  AND2_X1 U576bar ( .A1(n18bar), .A2(keybar[119]), .ZN(n470bar) );
  AND2_X1 U577 ( .A1(key[119]), .A2(n18), .ZN(n469) );
  OR2_X1 U577bar ( .A1(keybar[119]), .A2(n18bar), .ZN(n469bar) );
  OR2_X1 U578 ( .A1(n471), .A2(n19), .ZN(out[118]) );
  AND2_X1 U578bar ( .A1(n471bar), .A2(n19bar), .ZN(outbar[118]) );
  OR2_X1 U579 ( .A1(n20), .A2(key[118]), .ZN(n472) );
  AND2_X1 U579bar ( .A1(n20bar), .A2(keybar[118]), .ZN(n472bar) );
  AND2_X1 U580 ( .A1(key[118]), .A2(n20), .ZN(n471) );
  OR2_X1 U580bar ( .A1(keybar[118]), .A2(n20bar), .ZN(n471bar) );
  OR2_X1 U581 ( .A1(n473), .A2(n21), .ZN(out[117]) );
  AND2_X1 U581bar ( .A1(n473bar), .A2(n21bar), .ZN(outbar[117]) );
  OR2_X1 U582 ( .A1(n22), .A2(key[117]), .ZN(n474) );
  AND2_X1 U582bar ( .A1(n22bar), .A2(keybar[117]), .ZN(n474bar) );
  AND2_X1 U583 ( .A1(key[117]), .A2(n22), .ZN(n473) );
  OR2_X1 U583bar ( .A1(keybar[117]), .A2(n22bar), .ZN(n473bar) );
  OR2_X1 U584 ( .A1(n475), .A2(n23), .ZN(out[116]) );
  AND2_X1 U584bar ( .A1(n475bar), .A2(n23bar), .ZN(outbar[116]) );
  OR2_X1 U585 ( .A1(n24), .A2(key[116]), .ZN(n476) );
  AND2_X1 U585bar ( .A1(n24bar), .A2(keybar[116]), .ZN(n476bar) );
  AND2_X1 U586 ( .A1(key[116]), .A2(n24), .ZN(n475) );
  OR2_X1 U586bar ( .A1(keybar[116]), .A2(n24bar), .ZN(n475bar) );
  OR2_X1 U587 ( .A1(n477), .A2(n25), .ZN(out[115]) );
  AND2_X1 U587bar ( .A1(n477bar), .A2(n25bar), .ZN(outbar[115]) );
  OR2_X1 U588 ( .A1(n26), .A2(key[115]), .ZN(n478) );
  AND2_X1 U588bar ( .A1(n26bar), .A2(keybar[115]), .ZN(n478bar) );
  AND2_X1 U589 ( .A1(key[115]), .A2(n26), .ZN(n477) );
  OR2_X1 U589bar ( .A1(keybar[115]), .A2(n26bar), .ZN(n477bar) );
  OR2_X1 U590 ( .A1(n479), .A2(n27), .ZN(out[114]) );
  AND2_X1 U590bar ( .A1(n479bar), .A2(n27bar), .ZN(outbar[114]) );
  OR2_X1 U591 ( .A1(n28), .A2(key[114]), .ZN(n480) );
  AND2_X1 U591bar ( .A1(n28bar), .A2(keybar[114]), .ZN(n480bar) );
  AND2_X1 U592 ( .A1(key[114]), .A2(n28), .ZN(n479) );
  OR2_X1 U592bar ( .A1(keybar[114]), .A2(n28bar), .ZN(n479bar) );
  OR2_X1 U593 ( .A1(n481), .A2(n29), .ZN(out[113]) );
  AND2_X1 U593bar ( .A1(n481bar), .A2(n29bar), .ZN(outbar[113]) );
  OR2_X1 U594 ( .A1(n30), .A2(key[113]), .ZN(n482) );
  AND2_X1 U594bar ( .A1(n30bar), .A2(keybar[113]), .ZN(n482bar) );
  AND2_X1 U595 ( .A1(key[113]), .A2(n30), .ZN(n481) );
  OR2_X1 U595bar ( .A1(keybar[113]), .A2(n30bar), .ZN(n481bar) );
  OR2_X1 U596 ( .A1(n483), .A2(n31), .ZN(out[112]) );
  AND2_X1 U596bar ( .A1(n483bar), .A2(n31bar), .ZN(outbar[112]) );
  OR2_X1 U597 ( .A1(n32), .A2(key[112]), .ZN(n484) );
  AND2_X1 U597bar ( .A1(n32bar), .A2(keybar[112]), .ZN(n484bar) );
  AND2_X1 U598 ( .A1(key[112]), .A2(n32), .ZN(n483) );
  OR2_X1 U598bar ( .A1(keybar[112]), .A2(n32bar), .ZN(n483bar) );
  OR2_X1 U599 ( .A1(n485), .A2(n33), .ZN(out[111]) );
  AND2_X1 U599bar ( .A1(n485bar), .A2(n33bar), .ZN(outbar[111]) );
  OR2_X1 U600 ( .A1(n34), .A2(key[111]), .ZN(n486) );
  AND2_X1 U600bar ( .A1(n34bar), .A2(keybar[111]), .ZN(n486bar) );
  AND2_X1 U601 ( .A1(key[111]), .A2(n34), .ZN(n485) );
  OR2_X1 U601bar ( .A1(keybar[111]), .A2(n34bar), .ZN(n485bar) );
  OR2_X1 U602 ( .A1(n487), .A2(n35), .ZN(out[110]) );
  AND2_X1 U602bar ( .A1(n487bar), .A2(n35bar), .ZN(outbar[110]) );
  OR2_X1 U603 ( .A1(n36), .A2(key[110]), .ZN(n488) );
  AND2_X1 U603bar ( .A1(n36bar), .A2(keybar[110]), .ZN(n488bar) );
  AND2_X1 U604 ( .A1(key[110]), .A2(n36), .ZN(n487) );
  OR2_X1 U604bar ( .A1(keybar[110]), .A2(n36bar), .ZN(n487bar) );
  OR2_X1 U605 ( .A1(n489), .A2(n235), .ZN(out[10]) );
  AND2_X1 U605bar ( .A1(n489bar), .A2(n235bar), .ZN(outbar[10]) );
  OR2_X1 U606 ( .A1(n236), .A2(key[10]), .ZN(n490) );
  AND2_X1 U606bar ( .A1(n236bar), .A2(keybar[10]), .ZN(n490bar) );
  AND2_X1 U607 ( .A1(key[10]), .A2(n236), .ZN(n489) );
  OR2_X1 U607bar ( .A1(keybar[10]), .A2(n236bar), .ZN(n489bar) );
  OR2_X1 U608 ( .A1(n491), .A2(n37), .ZN(out[109]) );
  AND2_X1 U608bar ( .A1(n491bar), .A2(n37bar), .ZN(outbar[109]) );
  OR2_X1 U609 ( .A1(n38), .A2(key[109]), .ZN(n492) );
  AND2_X1 U609bar ( .A1(n38bar), .A2(keybar[109]), .ZN(n492bar) );
  AND2_X1 U610 ( .A1(key[109]), .A2(n38), .ZN(n491) );
  OR2_X1 U610bar ( .A1(keybar[109]), .A2(n38bar), .ZN(n491bar) );
  OR2_X1 U611 ( .A1(n493), .A2(n39), .ZN(out[108]) );
  AND2_X1 U611bar ( .A1(n493bar), .A2(n39bar), .ZN(outbar[108]) );
  OR2_X1 U612 ( .A1(n40), .A2(key[108]), .ZN(n494) );
  AND2_X1 U612bar ( .A1(n40bar), .A2(keybar[108]), .ZN(n494bar) );
  AND2_X1 U613 ( .A1(key[108]), .A2(n40), .ZN(n493) );
  OR2_X1 U613bar ( .A1(keybar[108]), .A2(n40bar), .ZN(n493bar) );
  OR2_X1 U614 ( .A1(n495), .A2(n41), .ZN(out[107]) );
  AND2_X1 U614bar ( .A1(n495bar), .A2(n41bar), .ZN(outbar[107]) );
  OR2_X1 U615 ( .A1(n42), .A2(key[107]), .ZN(n496) );
  AND2_X1 U615bar ( .A1(n42bar), .A2(keybar[107]), .ZN(n496bar) );
  AND2_X1 U616 ( .A1(key[107]), .A2(n42), .ZN(n495) );
  OR2_X1 U616bar ( .A1(keybar[107]), .A2(n42bar), .ZN(n495bar) );
  OR2_X1 U617 ( .A1(n497), .A2(n43), .ZN(out[106]) );
  AND2_X1 U617bar ( .A1(n497bar), .A2(n43bar), .ZN(outbar[106]) );
  OR2_X1 U618 ( .A1(n44), .A2(key[106]), .ZN(n498) );
  AND2_X1 U618bar ( .A1(n44bar), .A2(keybar[106]), .ZN(n498bar) );
  AND2_X1 U619 ( .A1(key[106]), .A2(n44), .ZN(n497) );
  OR2_X1 U619bar ( .A1(keybar[106]), .A2(n44bar), .ZN(n497bar) );
  OR2_X1 U620 ( .A1(n499), .A2(n45), .ZN(out[105]) );
  AND2_X1 U620bar ( .A1(n499bar), .A2(n45bar), .ZN(outbar[105]) );
  OR2_X1 U621 ( .A1(n46), .A2(key[105]), .ZN(n500) );
  AND2_X1 U621bar ( .A1(n46bar), .A2(keybar[105]), .ZN(n500bar) );
  AND2_X1 U622 ( .A1(key[105]), .A2(n46), .ZN(n499) );
  OR2_X1 U622bar ( .A1(keybar[105]), .A2(n46bar), .ZN(n499bar) );
  OR2_X1 U623 ( .A1(n501), .A2(n47), .ZN(out[104]) );
  AND2_X1 U623bar ( .A1(n501bar), .A2(n47bar), .ZN(outbar[104]) );
  OR2_X1 U624 ( .A1(n48), .A2(key[104]), .ZN(n502) );
  AND2_X1 U624bar ( .A1(n48bar), .A2(keybar[104]), .ZN(n502bar) );
  AND2_X1 U625 ( .A1(key[104]), .A2(n48), .ZN(n501) );
  OR2_X1 U625bar ( .A1(keybar[104]), .A2(n48bar), .ZN(n501bar) );
  OR2_X1 U626 ( .A1(n503), .A2(n49), .ZN(out[103]) );
  AND2_X1 U626bar ( .A1(n503bar), .A2(n49bar), .ZN(outbar[103]) );
  OR2_X1 U627 ( .A1(n50), .A2(key[103]), .ZN(n504) );
  AND2_X1 U627bar ( .A1(n50bar), .A2(keybar[103]), .ZN(n504bar) );
  AND2_X1 U628 ( .A1(key[103]), .A2(n50), .ZN(n503) );
  OR2_X1 U628bar ( .A1(keybar[103]), .A2(n50bar), .ZN(n503bar) );
  OR2_X1 U629 ( .A1(n505), .A2(n51), .ZN(out[102]) );
  AND2_X1 U629bar ( .A1(n505bar), .A2(n51bar), .ZN(outbar[102]) );
  OR2_X1 U630 ( .A1(n52), .A2(key[102]), .ZN(n506) );
  AND2_X1 U630bar ( .A1(n52bar), .A2(keybar[102]), .ZN(n506bar) );
  AND2_X1 U631 ( .A1(key[102]), .A2(n52), .ZN(n505) );
  OR2_X1 U631bar ( .A1(keybar[102]), .A2(n52bar), .ZN(n505bar) );
  OR2_X1 U632 ( .A1(n507), .A2(n53), .ZN(out[101]) );
  AND2_X1 U632bar ( .A1(n507bar), .A2(n53bar), .ZN(outbar[101]) );
  OR2_X1 U633 ( .A1(n54), .A2(key[101]), .ZN(n508) );
  AND2_X1 U633bar ( .A1(n54bar), .A2(keybar[101]), .ZN(n508bar) );
  AND2_X1 U634 ( .A1(key[101]), .A2(n54), .ZN(n507) );
  OR2_X1 U634bar ( .A1(keybar[101]), .A2(n54bar), .ZN(n507bar) );
  OR2_X1 U635 ( .A1(n509), .A2(n55), .ZN(out[100]) );
  AND2_X1 U635bar ( .A1(n509bar), .A2(n55bar), .ZN(outbar[100]) );
  OR2_X1 U636 ( .A1(n56), .A2(key[100]), .ZN(n510) );
  AND2_X1 U636bar ( .A1(n56bar), .A2(keybar[100]), .ZN(n510bar) );
  AND2_X1 U637 ( .A1(key[100]), .A2(n56), .ZN(n509) );
  OR2_X1 U637bar ( .A1(keybar[100]), .A2(n56bar), .ZN(n509bar) );
  OR2_X1 U638 ( .A1(n511), .A2(n255), .ZN(out[0]) );
  AND2_X1 U638bar ( .A1(n511bar), .A2(n255bar), .ZN(outbar[0]) );
  OR2_X1 U639 ( .A1(n256), .A2(key[0]), .ZN(n512) );
  AND2_X1 U639bar ( .A1(n256bar), .A2(keybar[0]), .ZN(n512bar) );
  AND2_X1 U640 ( .A1(key[0]), .A2(n256), .ZN(n511) );
  OR2_X1 U640bar ( .A1(keybar[0]), .A2(n256bar), .ZN(n511bar) );
endmodule

//done
