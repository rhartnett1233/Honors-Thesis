
module sample_circuit ( in, out );
  input [255:0] in;
  //input_done

  output [7:0] out;
  //output_done

  wire   in_81, in_80, in_79, in_78, in_77, in_76, in_75, in_74, in_73, in_72,
         in_71, in_70, in_69, in_68, in_67, in_66, in_65, in_64, in_63, in_62,
         in_61, in_60, in_59, in_58, in_57, in_56, in_55, in_54, in_53, in_52,
         in_51, in_50, in_49, in_48, in_47, in_46, in_45, in_44, in_43, in_42,
         in_41, in_40, in_39, in_38, in_37, in_36, in_35, in_34, in_33, in_32,
         in_31, in_30, in_29, in_28, in_27, in_26, in_25, in_24, in_23, in_22,
         in_21, in_20, in_19, in_18, in_17, in_16, in_15, in_14, in_13, in_12,
         in_11, in_10, in_9, in_8, in_7, in_6, in_5, in_4, in_3, in_2, in_1,
         in_0, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972;
  //wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];

  OR2_X1 U1 ( .A1(n972), .A2(n971), .ZN(out[7]) );
  OR2_X1 U2 ( .A1(n970), .A2(n969), .ZN(n971) );
  OR2_X1 U3 ( .A1(n968), .A2(n967), .ZN(n969) );
  OR2_X1 U4 ( .A1(n966), .A2(n965), .ZN(n967) );
  OR2_X1 U5 ( .A1(n964), .A2(n963), .ZN(n968) );
  OR2_X1 U6 ( .A1(in[116]), .A2(n962), .ZN(n963) );
  OR2_X1 U7 ( .A1(n961), .A2(n960), .ZN(n970) );
  OR2_X1 U8 ( .A1(in[150]), .A2(in[127]), .ZN(n960) );
  OR2_X1 U9 ( .A1(in[160]), .A2(n959), .ZN(n961) );
  OR2_X1 U10 ( .A1(in[252]), .A2(in[168]), .ZN(n959) );
  OR2_X1 U11 ( .A1(n958), .A2(n957), .ZN(n972) );
  OR2_X1 U12 ( .A1(n956), .A2(n955), .ZN(n957) );
  OR2_X1 U13 ( .A1(in_17), .A2(in[96]), .ZN(n955) );
  OR2_X1 U14 ( .A1(in_23), .A2(n954), .ZN(n956) );
  OR2_X1 U15 ( .A1(in_31), .A2(in_26), .ZN(n954) );
  OR2_X1 U16 ( .A1(n953), .A2(n952), .ZN(n958) );
  OR2_X1 U17 ( .A1(in_58), .A2(in_4), .ZN(n952) );
  OR2_X1 U18 ( .A1(in_59), .A2(n951), .ZN(n953) );
  OR2_X1 U19 ( .A1(in_71), .A2(in_62), .ZN(n951) );
  OR2_X1 U20 ( .A1(n950), .A2(n949), .ZN(out[6]) );
  OR2_X1 U21 ( .A1(n948), .A2(n947), .ZN(n949) );
  OR2_X1 U22 ( .A1(n946), .A2(n945), .ZN(n947) );
  OR2_X1 U23 ( .A1(n944), .A2(n943), .ZN(n945) );
  OR2_X1 U24 ( .A1(n942), .A2(n941), .ZN(n946) );
  OR2_X1 U25 ( .A1(in[101]), .A2(n940), .ZN(n941) );
  OR2_X1 U26 ( .A1(n939), .A2(n938), .ZN(n948) );
  OR2_X1 U27 ( .A1(in[114]), .A2(in[104]), .ZN(n938) );
  OR2_X1 U28 ( .A1(in[128]), .A2(n937), .ZN(n939) );
  OR2_X1 U29 ( .A1(in[136]), .A2(in[134]), .ZN(n937) );
  OR2_X1 U30 ( .A1(n936), .A2(n935), .ZN(n950) );
  OR2_X1 U31 ( .A1(n934), .A2(n933), .ZN(n935) );
  OR2_X1 U32 ( .A1(in[177]), .A2(in[164]), .ZN(n933) );
  OR2_X1 U33 ( .A1(in[212]), .A2(n932), .ZN(n934) );
  OR2_X1 U34 ( .A1(in[248]), .A2(in[221]), .ZN(n932) );
  OR2_X1 U35 ( .A1(n931), .A2(n930), .ZN(n936) );
  OR2_X1 U36 ( .A1(in_18), .A2(in[93]), .ZN(n930) );
  OR2_X1 U37 ( .A1(in_31), .A2(n929), .ZN(n931) );
  OR2_X1 U38 ( .A1(in_7), .A2(in_39), .ZN(n929) );
  OR2_X1 U39 ( .A1(n928), .A2(n927), .ZN(out[5]) );
  OR2_X1 U40 ( .A1(n926), .A2(n925), .ZN(n927) );
  OR2_X1 U41 ( .A1(n924), .A2(n923), .ZN(n925) );
  OR2_X1 U42 ( .A1(n922), .A2(n921), .ZN(n923) );
  OR2_X1 U43 ( .A1(n940), .A2(n920), .ZN(n924) );
  OR2_X1 U44 ( .A1(in[111]), .A2(n919), .ZN(n920) );
  OR2_X1 U45 ( .A1(n918), .A2(n917), .ZN(n940) );
  OR2_X1 U46 ( .A1(n916), .A2(n915), .ZN(n917) );
  OR2_X1 U47 ( .A1(n914), .A2(n913), .ZN(n915) );
  OR2_X1 U48 ( .A1(in[140]), .A2(in[131]), .ZN(n913) );
  OR2_X1 U49 ( .A1(in[160]), .A2(in[144]), .ZN(n914) );
  OR2_X1 U50 ( .A1(n912), .A2(n911), .ZN(n916) );
  OR2_X1 U51 ( .A1(in[179]), .A2(in[174]), .ZN(n911) );
  OR2_X1 U52 ( .A1(in[188]), .A2(in[184]), .ZN(n912) );
  OR2_X1 U53 ( .A1(n910), .A2(n909), .ZN(n918) );
  OR2_X1 U54 ( .A1(n908), .A2(n907), .ZN(n909) );
  OR2_X1 U55 ( .A1(in[216]), .A2(in[200]), .ZN(n907) );
  OR2_X1 U56 ( .A1(in[228]), .A2(in[224]), .ZN(n908) );
  OR2_X1 U57 ( .A1(n906), .A2(n905), .ZN(n910) );
  OR2_X1 U58 ( .A1(in[247]), .A2(in[235]), .ZN(n905) );
  OR2_X1 U59 ( .A1(in_42), .A2(in[83]), .ZN(n906) );
  OR2_X1 U60 ( .A1(n904), .A2(n903), .ZN(n926) );
  OR2_X1 U61 ( .A1(in[166]), .A2(in[123]), .ZN(n903) );
  OR2_X1 U62 ( .A1(in[170]), .A2(n902), .ZN(n904) );
  OR2_X1 U63 ( .A1(in[194]), .A2(in[183]), .ZN(n902) );
  OR2_X1 U64 ( .A1(n901), .A2(n900), .ZN(n928) );
  OR2_X1 U65 ( .A1(n899), .A2(n898), .ZN(n900) );
  OR2_X1 U66 ( .A1(in[241]), .A2(in[238]), .ZN(n898) );
  OR2_X1 U67 ( .A1(in[250]), .A2(n897), .ZN(n899) );
  OR2_X1 U68 ( .A1(in_24), .A2(in[84]), .ZN(n897) );
  OR2_X1 U69 ( .A1(n896), .A2(n895), .ZN(n901) );
  OR2_X1 U70 ( .A1(in_41), .A2(in_29), .ZN(n895) );
  OR2_X1 U71 ( .A1(in_66), .A2(n894), .ZN(n896) );
  OR2_X1 U72 ( .A1(in_76), .A2(in_71), .ZN(n894) );
  OR2_X1 U73 ( .A1(n893), .A2(n892), .ZN(out[4]) );
  OR2_X1 U74 ( .A1(n891), .A2(n890), .ZN(n892) );
  OR2_X1 U75 ( .A1(n889), .A2(n888), .ZN(n890) );
  OR2_X1 U76 ( .A1(n922), .A2(n887), .ZN(n888) );
  OR2_X1 U77 ( .A1(n886), .A2(n885), .ZN(n922) );
  OR2_X1 U78 ( .A1(n884), .A2(n883), .ZN(n885) );
  OR2_X1 U79 ( .A1(n882), .A2(n881), .ZN(n883) );
  OR2_X1 U80 ( .A1(in[118]), .A2(in[109]), .ZN(n881) );
  OR2_X1 U81 ( .A1(in[139]), .A2(in[120]), .ZN(n882) );
  OR2_X1 U82 ( .A1(n880), .A2(n879), .ZN(n884) );
  OR2_X1 U83 ( .A1(in[198]), .A2(in[154]), .ZN(n879) );
  OR2_X1 U84 ( .A1(in[210]), .A2(in[205]), .ZN(n880) );
  OR2_X1 U85 ( .A1(n878), .A2(n877), .ZN(n886) );
  OR2_X1 U86 ( .A1(n876), .A2(n875), .ZN(n877) );
  OR2_X1 U87 ( .A1(in[219]), .A2(in[217]), .ZN(n875) );
  OR2_X1 U88 ( .A1(in[86]), .A2(in[252]), .ZN(n876) );
  OR2_X1 U89 ( .A1(n874), .A2(n873), .ZN(n878) );
  OR2_X1 U90 ( .A1(in_40), .A2(in[91]), .ZN(n873) );
  OR2_X1 U91 ( .A1(in_8), .A2(in_46), .ZN(n874) );
  OR2_X1 U92 ( .A1(n872), .A2(n871), .ZN(n889) );
  OR2_X1 U93 ( .A1(in[117]), .A2(n943), .ZN(n871) );
  OR2_X1 U94 ( .A1(n870), .A2(n869), .ZN(n943) );
  OR2_X1 U95 ( .A1(n868), .A2(n867), .ZN(n869) );
  OR2_X1 U96 ( .A1(n866), .A2(n865), .ZN(n867) );
  OR2_X1 U97 ( .A1(n864), .A2(n863), .ZN(n865) );
  OR2_X1 U98 ( .A1(in[108]), .A2(n919), .ZN(n866) );
  OR2_X1 U99 ( .A1(n862), .A2(n861), .ZN(n919) );
  OR2_X1 U100 ( .A1(n860), .A2(n859), .ZN(n861) );
  OR2_X1 U101 ( .A1(n858), .A2(n857), .ZN(n859) );
  OR2_X1 U102 ( .A1(in[119]), .A2(in[105]), .ZN(n857) );
  OR2_X1 U103 ( .A1(in[186]), .A2(in[175]), .ZN(n858) );
  OR2_X1 U104 ( .A1(n856), .A2(n855), .ZN(n860) );
  OR2_X1 U105 ( .A1(in[202]), .A2(in[193]), .ZN(n855) );
  OR2_X1 U106 ( .A1(in[225]), .A2(in[208]), .ZN(n856) );
  OR2_X1 U107 ( .A1(n854), .A2(n853), .ZN(n862) );
  OR2_X1 U108 ( .A1(n852), .A2(n851), .ZN(n853) );
  OR2_X1 U109 ( .A1(in_1), .A2(in[85]), .ZN(n851) );
  OR2_X1 U110 ( .A1(in_23), .A2(in_19), .ZN(n852) );
  OR2_X1 U111 ( .A1(n850), .A2(n849), .ZN(n854) );
  OR2_X1 U112 ( .A1(in_43), .A2(in_33), .ZN(n849) );
  OR2_X1 U113 ( .A1(in_63), .A2(in_44), .ZN(n850) );
  OR2_X1 U114 ( .A1(n848), .A2(n847), .ZN(n868) );
  OR2_X1 U115 ( .A1(in[141]), .A2(in[112]), .ZN(n847) );
  OR2_X1 U116 ( .A1(in[147]), .A2(n846), .ZN(n848) );
  OR2_X1 U117 ( .A1(in[181]), .A2(in[167]), .ZN(n846) );
  OR2_X1 U118 ( .A1(n845), .A2(n844), .ZN(n870) );
  OR2_X1 U119 ( .A1(n843), .A2(n842), .ZN(n844) );
  OR2_X1 U120 ( .A1(in[229]), .A2(in[201]), .ZN(n842) );
  OR2_X1 U121 ( .A1(in[237]), .A2(n841), .ZN(n843) );
  OR2_X1 U122 ( .A1(in[94]), .A2(in[253]), .ZN(n841) );
  OR2_X1 U123 ( .A1(n840), .A2(n839), .ZN(n845) );
  OR2_X1 U124 ( .A1(in_21), .A2(in[96]), .ZN(n839) );
  OR2_X1 U125 ( .A1(in_25), .A2(n838), .ZN(n840) );
  OR2_X1 U126 ( .A1(in_81), .A2(in_45), .ZN(n838) );
  OR2_X1 U127 ( .A1(n837), .A2(n836), .ZN(n891) );
  OR2_X1 U128 ( .A1(in[142]), .A2(in[124]), .ZN(n836) );
  OR2_X1 U129 ( .A1(in[150]), .A2(n835), .ZN(n837) );
  OR2_X1 U130 ( .A1(in[172]), .A2(in[155]), .ZN(n835) );
  OR2_X1 U131 ( .A1(n834), .A2(n833), .ZN(n893) );
  OR2_X1 U132 ( .A1(n832), .A2(n831), .ZN(n833) );
  OR2_X1 U133 ( .A1(in[196]), .A2(in[173]), .ZN(n831) );
  OR2_X1 U134 ( .A1(in[222]), .A2(n830), .ZN(n832) );
  OR2_X1 U135 ( .A1(in[227]), .A2(in[226]), .ZN(n830) );
  OR2_X1 U136 ( .A1(n829), .A2(n828), .ZN(n834) );
  OR2_X1 U137 ( .A1(in[249]), .A2(in[231]), .ZN(n828) );
  OR2_X1 U138 ( .A1(in_28), .A2(n827), .ZN(n829) );
  OR2_X1 U139 ( .A1(in_52), .A2(in_47), .ZN(n827) );
  OR2_X1 U140 ( .A1(n826), .A2(n825), .ZN(out[3]) );
  OR2_X1 U141 ( .A1(n824), .A2(n823), .ZN(n825) );
  OR2_X1 U142 ( .A1(n822), .A2(n821), .ZN(n823) );
  OR2_X1 U143 ( .A1(n820), .A2(n819), .ZN(n821) );
  OR2_X1 U144 ( .A1(n964), .A2(n818), .ZN(n822) );
  OR2_X1 U145 ( .A1(in[118]), .A2(n817), .ZN(n818) );
  OR2_X1 U146 ( .A1(n816), .A2(n815), .ZN(n964) );
  OR2_X1 U147 ( .A1(n814), .A2(n813), .ZN(n815) );
  OR2_X1 U148 ( .A1(n812), .A2(n811), .ZN(n813) );
  OR2_X1 U149 ( .A1(in[122]), .A2(in[111]), .ZN(n811) );
  OR2_X1 U150 ( .A1(in[154]), .A2(in[151]), .ZN(n812) );
  OR2_X1 U151 ( .A1(n810), .A2(n809), .ZN(n814) );
  OR2_X1 U152 ( .A1(in[187]), .A2(in[177]), .ZN(n809) );
  OR2_X1 U153 ( .A1(in[200]), .A2(in[192]), .ZN(n810) );
  OR2_X1 U154 ( .A1(n808), .A2(n807), .ZN(n816) );
  OR2_X1 U155 ( .A1(n806), .A2(n805), .ZN(n807) );
  OR2_X1 U156 ( .A1(in[225]), .A2(in[207]), .ZN(n805) );
  OR2_X1 U157 ( .A1(in[98]), .A2(in[226]), .ZN(n806) );
  OR2_X1 U158 ( .A1(n804), .A2(n803), .ZN(n808) );
  OR2_X1 U159 ( .A1(in_20), .A2(in_16), .ZN(n803) );
  OR2_X1 U160 ( .A1(in_55), .A2(in_45), .ZN(n804) );
  OR2_X1 U161 ( .A1(n802), .A2(n801), .ZN(n824) );
  OR2_X1 U162 ( .A1(in[162]), .A2(in[149]), .ZN(n801) );
  OR2_X1 U163 ( .A1(in[163]), .A2(n800), .ZN(n802) );
  OR2_X1 U164 ( .A1(in[191]), .A2(in[189]), .ZN(n800) );
  OR2_X1 U165 ( .A1(n799), .A2(n798), .ZN(n826) );
  OR2_X1 U166 ( .A1(n797), .A2(n796), .ZN(n798) );
  OR2_X1 U167 ( .A1(in[212]), .A2(in[193]), .ZN(n796) );
  OR2_X1 U168 ( .A1(in[238]), .A2(n795), .ZN(n797) );
  OR2_X1 U169 ( .A1(in[88]), .A2(in[247]), .ZN(n795) );
  OR2_X1 U170 ( .A1(n794), .A2(n793), .ZN(n799) );
  OR2_X1 U171 ( .A1(in[94]), .A2(in[92]), .ZN(n793) );
  OR2_X1 U172 ( .A1(in_52), .A2(n792), .ZN(n794) );
  OR2_X1 U173 ( .A1(in_70), .A2(in_67), .ZN(n792) );
  OR2_X1 U174 ( .A1(n791), .A2(n790), .ZN(out[2]) );
  OR2_X1 U175 ( .A1(n789), .A2(n788), .ZN(n790) );
  OR2_X1 U176 ( .A1(n787), .A2(n786), .ZN(n788) );
  OR2_X1 U177 ( .A1(n819), .A2(n785), .ZN(n786) );
  OR2_X1 U178 ( .A1(n784), .A2(n783), .ZN(n819) );
  OR2_X1 U179 ( .A1(n782), .A2(n781), .ZN(n783) );
  OR2_X1 U180 ( .A1(n780), .A2(n779), .ZN(n781) );
  OR2_X1 U181 ( .A1(n962), .A2(n778), .ZN(n779) );
  OR2_X1 U182 ( .A1(n777), .A2(n776), .ZN(n962) );
  OR2_X1 U183 ( .A1(n775), .A2(n774), .ZN(n776) );
  OR2_X1 U184 ( .A1(n773), .A2(n772), .ZN(n774) );
  OR2_X1 U185 ( .A1(in[131]), .A2(in[120]), .ZN(n772) );
  OR2_X1 U186 ( .A1(in[153]), .A2(in[147]), .ZN(n773) );
  OR2_X1 U187 ( .A1(n771), .A2(n770), .ZN(n775) );
  OR2_X1 U188 ( .A1(in[170]), .A2(in[156]), .ZN(n770) );
  OR2_X1 U189 ( .A1(in[223]), .A2(in[190]), .ZN(n771) );
  OR2_X1 U190 ( .A1(n769), .A2(n768), .ZN(n777) );
  OR2_X1 U191 ( .A1(n767), .A2(n766), .ZN(n768) );
  OR2_X1 U192 ( .A1(in[236]), .A2(in[230]), .ZN(n766) );
  OR2_X1 U193 ( .A1(in[85]), .A2(in[240]), .ZN(n767) );
  OR2_X1 U194 ( .A1(n765), .A2(n764), .ZN(n769) );
  OR2_X1 U195 ( .A1(in_12), .A2(in[90]), .ZN(n764) );
  OR2_X1 U196 ( .A1(in_39), .A2(in_28), .ZN(n765) );
  OR2_X1 U197 ( .A1(in[109]), .A2(n763), .ZN(n780) );
  OR2_X1 U198 ( .A1(n762), .A2(n761), .ZN(n782) );
  OR2_X1 U199 ( .A1(in[138]), .A2(in[129]), .ZN(n761) );
  OR2_X1 U200 ( .A1(in[157]), .A2(n760), .ZN(n762) );
  OR2_X1 U201 ( .A1(in[182]), .A2(in[167]), .ZN(n760) );
  OR2_X1 U202 ( .A1(n759), .A2(n758), .ZN(n784) );
  OR2_X1 U203 ( .A1(n757), .A2(n756), .ZN(n758) );
  OR2_X1 U204 ( .A1(in[195]), .A2(in[184]), .ZN(n756) );
  OR2_X1 U205 ( .A1(in[196]), .A2(n755), .ZN(n757) );
  OR2_X1 U206 ( .A1(in[215]), .A2(in[209]), .ZN(n755) );
  OR2_X1 U207 ( .A1(n754), .A2(n753), .ZN(n759) );
  OR2_X1 U208 ( .A1(in[93]), .A2(in[233]), .ZN(n753) );
  OR2_X1 U209 ( .A1(in_1), .A2(n752), .ZN(n754) );
  OR2_X1 U210 ( .A1(in_69), .A2(in_66), .ZN(n752) );
  OR2_X1 U211 ( .A1(n966), .A2(n751), .ZN(n787) );
  OR2_X1 U212 ( .A1(in[134]), .A2(n750), .ZN(n751) );
  OR2_X1 U213 ( .A1(n749), .A2(n748), .ZN(n966) );
  OR2_X1 U214 ( .A1(n747), .A2(n746), .ZN(n748) );
  OR2_X1 U215 ( .A1(n745), .A2(n744), .ZN(n746) );
  OR2_X1 U216 ( .A1(in[136]), .A2(in[121]), .ZN(n744) );
  OR2_X1 U217 ( .A1(in[186]), .A2(in[174]), .ZN(n745) );
  OR2_X1 U218 ( .A1(n743), .A2(n742), .ZN(n747) );
  OR2_X1 U219 ( .A1(in[198]), .A2(in[197]), .ZN(n742) );
  OR2_X1 U220 ( .A1(in[214]), .A2(in[199]), .ZN(n743) );
  OR2_X1 U221 ( .A1(n741), .A2(n740), .ZN(n749) );
  OR2_X1 U222 ( .A1(n739), .A2(n738), .ZN(n740) );
  OR2_X1 U223 ( .A1(in[231]), .A2(in[220]), .ZN(n738) );
  OR2_X1 U224 ( .A1(in_25), .A2(in[245]), .ZN(n739) );
  OR2_X1 U225 ( .A1(n737), .A2(n736), .ZN(n741) );
  OR2_X1 U226 ( .A1(in_53), .A2(in_29), .ZN(n736) );
  OR2_X1 U227 ( .A1(in_79), .A2(in_74), .ZN(n737) );
  OR2_X1 U228 ( .A1(n735), .A2(n734), .ZN(n789) );
  OR2_X1 U229 ( .A1(in[152]), .A2(in[140]), .ZN(n734) );
  OR2_X1 U230 ( .A1(in[155]), .A2(n733), .ZN(n735) );
  OR2_X1 U231 ( .A1(in[166]), .A2(in[165]), .ZN(n733) );
  OR2_X1 U232 ( .A1(n732), .A2(n731), .ZN(n791) );
  OR2_X1 U233 ( .A1(n730), .A2(n729), .ZN(n731) );
  OR2_X1 U234 ( .A1(in[202]), .A2(in[185]), .ZN(n729) );
  OR2_X1 U235 ( .A1(in[211]), .A2(n728), .ZN(n730) );
  OR2_X1 U236 ( .A1(in[255]), .A2(in[253]), .ZN(n728) );
  OR2_X1 U237 ( .A1(n727), .A2(n726), .ZN(n732) );
  OR2_X1 U238 ( .A1(in_35), .A2(in_15), .ZN(n726) );
  OR2_X1 U239 ( .A1(in_36), .A2(n725), .ZN(n727) );
  OR2_X1 U240 ( .A1(in_48), .A2(in_40), .ZN(n725) );
  OR2_X1 U241 ( .A1(n724), .A2(n723), .ZN(out[1]) );
  OR2_X1 U242 ( .A1(n722), .A2(n721), .ZN(n723) );
  OR2_X1 U243 ( .A1(n720), .A2(n719), .ZN(n721) );
  OR2_X1 U244 ( .A1(n921), .A2(n887), .ZN(n719) );
  OR2_X1 U245 ( .A1(n718), .A2(n717), .ZN(n887) );
  OR2_X1 U246 ( .A1(n716), .A2(n715), .ZN(n717) );
  OR2_X1 U247 ( .A1(n714), .A2(n713), .ZN(n715) );
  OR2_X1 U248 ( .A1(in[116]), .A2(in[110]), .ZN(n713) );
  OR2_X1 U249 ( .A1(in[133]), .A2(in[130]), .ZN(n714) );
  OR2_X1 U250 ( .A1(n712), .A2(n711), .ZN(n716) );
  OR2_X1 U251 ( .A1(in[203]), .A2(in[135]), .ZN(n711) );
  OR2_X1 U252 ( .A1(in[232]), .A2(in[223]), .ZN(n712) );
  OR2_X1 U253 ( .A1(n710), .A2(n709), .ZN(n718) );
  OR2_X1 U254 ( .A1(n708), .A2(n707), .ZN(n709) );
  OR2_X1 U255 ( .A1(in[255]), .A2(in[233]), .ZN(n707) );
  OR2_X1 U256 ( .A1(in_53), .A2(in_34), .ZN(n708) );
  OR2_X1 U257 ( .A1(n706), .A2(n705), .ZN(n710) );
  OR2_X1 U258 ( .A1(in_57), .A2(in_55), .ZN(n705) );
  OR2_X1 U259 ( .A1(in_68), .A2(in_67), .ZN(n706) );
  OR2_X1 U260 ( .A1(n704), .A2(n703), .ZN(n921) );
  OR2_X1 U261 ( .A1(n702), .A2(n701), .ZN(n703) );
  OR2_X1 U262 ( .A1(n700), .A2(n699), .ZN(n701) );
  OR2_X1 U263 ( .A1(n944), .A2(n872), .ZN(n699) );
  OR2_X1 U264 ( .A1(n698), .A2(n697), .ZN(n872) );
  OR2_X1 U265 ( .A1(n696), .A2(n695), .ZN(n697) );
  OR2_X1 U266 ( .A1(n694), .A2(n693), .ZN(n695) );
  OR2_X1 U267 ( .A1(in[121]), .A2(in[102]), .ZN(n693) );
  OR2_X1 U268 ( .A1(in[162]), .A2(in[161]), .ZN(n694) );
  OR2_X1 U269 ( .A1(n692), .A2(n691), .ZN(n696) );
  OR2_X1 U270 ( .A1(in[192]), .A2(in[178]), .ZN(n691) );
  OR2_X1 U271 ( .A1(in[244]), .A2(in[209]), .ZN(n692) );
  OR2_X1 U272 ( .A1(n690), .A2(n689), .ZN(n698) );
  OR2_X1 U273 ( .A1(n688), .A2(n687), .ZN(n689) );
  OR2_X1 U274 ( .A1(in[90]), .A2(in[254]), .ZN(n687) );
  OR2_X1 U275 ( .A1(in_36), .A2(in_32), .ZN(n688) );
  OR2_X1 U276 ( .A1(n686), .A2(n685), .ZN(n690) );
  OR2_X1 U277 ( .A1(in_62), .A2(in_37), .ZN(n685) );
  OR2_X1 U278 ( .A1(in_75), .A2(in_73), .ZN(n686) );
  OR2_X1 U279 ( .A1(n684), .A2(n683), .ZN(n944) );
  OR2_X1 U280 ( .A1(n682), .A2(n681), .ZN(n683) );
  OR2_X1 U281 ( .A1(n680), .A2(n679), .ZN(n681) );
  OR2_X1 U282 ( .A1(in[171]), .A2(in[153]), .ZN(n679) );
  OR2_X1 U283 ( .A1(in[187]), .A2(in[176]), .ZN(n680) );
  OR2_X1 U284 ( .A1(n678), .A2(n677), .ZN(n682) );
  OR2_X1 U285 ( .A1(in[245]), .A2(in[211]), .ZN(n677) );
  OR2_X1 U286 ( .A1(in[97]), .A2(in[88]), .ZN(n678) );
  OR2_X1 U287 ( .A1(n676), .A2(n675), .ZN(n684) );
  OR2_X1 U288 ( .A1(n674), .A2(n673), .ZN(n675) );
  OR2_X1 U289 ( .A1(in_10), .A2(in_0), .ZN(n673) );
  OR2_X1 U290 ( .A1(in_59), .A2(in_5), .ZN(n674) );
  OR2_X1 U291 ( .A1(n672), .A2(n671), .ZN(n676) );
  OR2_X1 U292 ( .A1(in_60), .A2(in_6), .ZN(n671) );
  OR2_X1 U293 ( .A1(in_77), .A2(in_69), .ZN(n672) );
  OR2_X1 U294 ( .A1(in[113]), .A2(n864), .ZN(n700) );
  OR2_X1 U295 ( .A1(n670), .A2(n669), .ZN(n864) );
  OR2_X1 U296 ( .A1(n668), .A2(n667), .ZN(n669) );
  OR2_X1 U297 ( .A1(n666), .A2(n665), .ZN(n667) );
  OR2_X1 U298 ( .A1(in[125]), .A2(in[107]), .ZN(n665) );
  OR2_X1 U299 ( .A1(in[138]), .A2(in[126]), .ZN(n666) );
  OR2_X1 U300 ( .A1(n664), .A2(n663), .ZN(n668) );
  OR2_X1 U301 ( .A1(in[189]), .A2(in[143]), .ZN(n663) );
  OR2_X1 U302 ( .A1(in[99]), .A2(in[214]), .ZN(n664) );
  OR2_X1 U303 ( .A1(n662), .A2(n661), .ZN(n670) );
  OR2_X1 U304 ( .A1(n660), .A2(n659), .ZN(n661) );
  OR2_X1 U305 ( .A1(in_15), .A2(in_12), .ZN(n659) );
  OR2_X1 U306 ( .A1(in_20), .A2(in_2), .ZN(n660) );
  OR2_X1 U307 ( .A1(n658), .A2(n657), .ZN(n662) );
  OR2_X1 U308 ( .A1(in_30), .A2(in_3), .ZN(n657) );
  OR2_X1 U309 ( .A1(in_4), .A2(in_38), .ZN(n658) );
  OR2_X1 U310 ( .A1(n656), .A2(n655), .ZN(n702) );
  OR2_X1 U311 ( .A1(in[148]), .A2(in[137]), .ZN(n655) );
  OR2_X1 U312 ( .A1(in[149]), .A2(n654), .ZN(n656) );
  OR2_X1 U313 ( .A1(in[195]), .A2(in[190]), .ZN(n654) );
  OR2_X1 U314 ( .A1(n653), .A2(n652), .ZN(n704) );
  OR2_X1 U315 ( .A1(n651), .A2(n650), .ZN(n652) );
  OR2_X1 U316 ( .A1(in[98]), .A2(in[197]), .ZN(n650) );
  OR2_X1 U317 ( .A1(in_11), .A2(n649), .ZN(n651) );
  OR2_X1 U318 ( .A1(in_26), .A2(in_14), .ZN(n649) );
  OR2_X1 U319 ( .A1(n648), .A2(n647), .ZN(n653) );
  OR2_X1 U320 ( .A1(in_35), .A2(in_27), .ZN(n647) );
  OR2_X1 U321 ( .A1(in_50), .A2(n646), .ZN(n648) );
  OR2_X1 U322 ( .A1(in_78), .A2(in_61), .ZN(n646) );
  OR2_X1 U323 ( .A1(n942), .A2(n645), .ZN(n720) );
  OR2_X1 U324 ( .A1(in[106]), .A2(n863), .ZN(n645) );
  OR2_X1 U325 ( .A1(n644), .A2(n643), .ZN(n863) );
  OR2_X1 U326 ( .A1(n642), .A2(n641), .ZN(n643) );
  OR2_X1 U327 ( .A1(n640), .A2(n639), .ZN(n641) );
  OR2_X1 U328 ( .A1(in[127]), .A2(in[122]), .ZN(n639) );
  OR2_X1 U329 ( .A1(in[156]), .A2(in[132]), .ZN(n640) );
  OR2_X1 U330 ( .A1(n638), .A2(n637), .ZN(n642) );
  OR2_X1 U331 ( .A1(in[159]), .A2(in[157]), .ZN(n637) );
  OR2_X1 U332 ( .A1(in[185]), .A2(in[169]), .ZN(n638) );
  OR2_X1 U333 ( .A1(n636), .A2(n635), .ZN(n644) );
  OR2_X1 U334 ( .A1(n634), .A2(n633), .ZN(n635) );
  OR2_X1 U335 ( .A1(in[239]), .A2(in[218]), .ZN(n633) );
  OR2_X1 U336 ( .A1(in_13), .A2(in[87]), .ZN(n634) );
  OR2_X1 U337 ( .A1(n632), .A2(n631), .ZN(n636) );
  OR2_X1 U338 ( .A1(in_72), .A2(in_70), .ZN(n631) );
  OR2_X1 U339 ( .A1(in_80), .A2(in_74), .ZN(n632) );
  OR2_X1 U340 ( .A1(n630), .A2(n629), .ZN(n942) );
  OR2_X1 U341 ( .A1(n628), .A2(n627), .ZN(n629) );
  OR2_X1 U342 ( .A1(n626), .A2(n625), .ZN(n627) );
  OR2_X1 U343 ( .A1(in[146]), .A2(in[100]), .ZN(n625) );
  OR2_X1 U344 ( .A1(in[168]), .A2(in[152]), .ZN(n626) );
  OR2_X1 U345 ( .A1(n624), .A2(n623), .ZN(n628) );
  OR2_X1 U346 ( .A1(in[199]), .A2(in[182]), .ZN(n623) );
  OR2_X1 U347 ( .A1(in[236]), .A2(in[204]), .ZN(n624) );
  OR2_X1 U348 ( .A1(n622), .A2(n621), .ZN(n630) );
  OR2_X1 U349 ( .A1(n620), .A2(n619), .ZN(n621) );
  OR2_X1 U350 ( .A1(in[89]), .A2(in[246]), .ZN(n619) );
  OR2_X1 U351 ( .A1(in[95]), .A2(in[92]), .ZN(n620) );
  OR2_X1 U352 ( .A1(n618), .A2(n617), .ZN(n622) );
  OR2_X1 U353 ( .A1(in_22), .A2(in_16), .ZN(n617) );
  OR2_X1 U354 ( .A1(in_51), .A2(in_49), .ZN(n618) );
  OR2_X1 U355 ( .A1(n616), .A2(n615), .ZN(n722) );
  OR2_X1 U356 ( .A1(in[158]), .A2(in[115]), .ZN(n615) );
  OR2_X1 U357 ( .A1(in[163]), .A2(n614), .ZN(n616) );
  OR2_X1 U358 ( .A1(in[206]), .A2(in[165]), .ZN(n614) );
  OR2_X1 U359 ( .A1(n613), .A2(n612), .ZN(n724) );
  OR2_X1 U360 ( .A1(n611), .A2(n610), .ZN(n612) );
  OR2_X1 U361 ( .A1(in[213]), .A2(in[207]), .ZN(n610) );
  OR2_X1 U362 ( .A1(in[215]), .A2(n609), .ZN(n611) );
  OR2_X1 U363 ( .A1(in[230]), .A2(in[220]), .ZN(n609) );
  OR2_X1 U364 ( .A1(n608), .A2(n607), .ZN(n613) );
  OR2_X1 U365 ( .A1(in[251]), .A2(in[234]), .ZN(n607) );
  OR2_X1 U366 ( .A1(in_17), .A2(n606), .ZN(n608) );
  OR2_X1 U367 ( .A1(in_65), .A2(in_56), .ZN(n606) );
  OR2_X1 U368 ( .A1(n605), .A2(n604), .ZN(out[0]) );
  OR2_X1 U369 ( .A1(n603), .A2(n602), .ZN(n604) );
  OR2_X1 U370 ( .A1(n601), .A2(n600), .ZN(n602) );
  OR2_X1 U371 ( .A1(n820), .A2(n785), .ZN(n600) );
  OR2_X1 U372 ( .A1(n599), .A2(n598), .ZN(n785) );
  OR2_X1 U373 ( .A1(n597), .A2(n596), .ZN(n598) );
  OR2_X1 U374 ( .A1(n595), .A2(n594), .ZN(n596) );
  OR2_X1 U375 ( .A1(in[135]), .A2(in[104]), .ZN(n594) );
  OR2_X1 U376 ( .A1(in[188]), .A2(in[178]), .ZN(n595) );
  OR2_X1 U377 ( .A1(n593), .A2(n592), .ZN(n597) );
  OR2_X1 U378 ( .A1(in[217]), .A2(in[194]), .ZN(n592) );
  OR2_X1 U379 ( .A1(in[237]), .A2(in[218]), .ZN(n593) );
  OR2_X1 U380 ( .A1(n591), .A2(n590), .ZN(n599) );
  OR2_X1 U381 ( .A1(n589), .A2(n588), .ZN(n590) );
  OR2_X1 U382 ( .A1(in_2), .A2(in_10), .ZN(n588) );
  OR2_X1 U383 ( .A1(in_47), .A2(in_22), .ZN(n589) );
  OR2_X1 U384 ( .A1(n587), .A2(n586), .ZN(n591) );
  OR2_X1 U385 ( .A1(in_56), .A2(in_54), .ZN(n586) );
  OR2_X1 U386 ( .A1(in_63), .A2(in_61), .ZN(n587) );
  OR2_X1 U387 ( .A1(n585), .A2(n584), .ZN(n820) );
  OR2_X1 U388 ( .A1(n583), .A2(n582), .ZN(n584) );
  OR2_X1 U389 ( .A1(n581), .A2(n580), .ZN(n582) );
  OR2_X1 U390 ( .A1(in[158]), .A2(in[142]), .ZN(n580) );
  OR2_X1 U391 ( .A1(in[175]), .A2(in[164]), .ZN(n581) );
  OR2_X1 U392 ( .A1(n579), .A2(n578), .ZN(n583) );
  OR2_X1 U393 ( .A1(in[228]), .A2(in[204]), .ZN(n578) );
  OR2_X1 U394 ( .A1(in[91]), .A2(in[87]), .ZN(n579) );
  OR2_X1 U395 ( .A1(n577), .A2(n576), .ZN(n585) );
  OR2_X1 U396 ( .A1(n575), .A2(n574), .ZN(n576) );
  OR2_X1 U397 ( .A1(in_21), .A2(in_11), .ZN(n574) );
  OR2_X1 U398 ( .A1(in_5), .A2(in_3), .ZN(n575) );
  OR2_X1 U399 ( .A1(n573), .A2(n572), .ZN(n577) );
  OR2_X1 U400 ( .A1(in_68), .A2(in_64), .ZN(n572) );
  OR2_X1 U401 ( .A1(in_76), .A2(in_73), .ZN(n573) );
  OR2_X1 U402 ( .A1(n778), .A2(n571), .ZN(n601) );
  OR2_X1 U403 ( .A1(in[100]), .A2(n965), .ZN(n571) );
  OR2_X1 U404 ( .A1(n570), .A2(n569), .ZN(n965) );
  OR2_X1 U405 ( .A1(n568), .A2(n567), .ZN(n569) );
  OR2_X1 U406 ( .A1(n566), .A2(n565), .ZN(n567) );
  OR2_X1 U407 ( .A1(n817), .A2(n750), .ZN(n565) );
  OR2_X1 U408 ( .A1(n564), .A2(n563), .ZN(n750) );
  OR2_X1 U409 ( .A1(n562), .A2(n561), .ZN(n563) );
  OR2_X1 U410 ( .A1(n560), .A2(n559), .ZN(n561) );
  OR2_X1 U411 ( .A1(in[119]), .A2(in[103]), .ZN(n559) );
  OR2_X1 U412 ( .A1(in[137]), .A2(in[133]), .ZN(n560) );
  OR2_X1 U413 ( .A1(n558), .A2(n557), .ZN(n562) );
  OR2_X1 U414 ( .A1(in[176]), .A2(in[173]), .ZN(n557) );
  OR2_X1 U415 ( .A1(in[210]), .A2(in[181]), .ZN(n558) );
  OR2_X1 U416 ( .A1(n556), .A2(n555), .ZN(n564) );
  OR2_X1 U417 ( .A1(n554), .A2(n553), .ZN(n555) );
  OR2_X1 U418 ( .A1(in_13), .A2(in[234]), .ZN(n553) );
  OR2_X1 U419 ( .A1(in_38), .A2(in_32), .ZN(n554) );
  OR2_X1 U420 ( .A1(n552), .A2(n551), .ZN(n556) );
  OR2_X1 U421 ( .A1(in_42), .A2(in_41), .ZN(n551) );
  OR2_X1 U422 ( .A1(in_7), .A2(in_49), .ZN(n552) );
  OR2_X1 U423 ( .A1(n550), .A2(n549), .ZN(n817) );
  OR2_X1 U424 ( .A1(n548), .A2(n547), .ZN(n549) );
  OR2_X1 U425 ( .A1(n546), .A2(n545), .ZN(n547) );
  OR2_X1 U426 ( .A1(in[159]), .A2(in[105]), .ZN(n545) );
  OR2_X1 U427 ( .A1(in[206]), .A2(in[183]), .ZN(n546) );
  OR2_X1 U428 ( .A1(n544), .A2(n543), .ZN(n548) );
  OR2_X1 U429 ( .A1(in[229]), .A2(in[219]), .ZN(n543) );
  OR2_X1 U430 ( .A1(in[235]), .A2(in[232]), .ZN(n544) );
  OR2_X1 U431 ( .A1(n542), .A2(n541), .ZN(n550) );
  OR2_X1 U432 ( .A1(n540), .A2(n539), .ZN(n541) );
  OR2_X1 U433 ( .A1(in[249]), .A2(in[242]), .ZN(n539) );
  OR2_X1 U434 ( .A1(in[89]), .A2(in[254]), .ZN(n540) );
  OR2_X1 U435 ( .A1(n538), .A2(n537), .ZN(n542) );
  OR2_X1 U436 ( .A1(in_14), .A2(in[99]), .ZN(n537) );
  OR2_X1 U437 ( .A1(in_60), .A2(in_18), .ZN(n538) );
  OR2_X1 U438 ( .A1(in[113]), .A2(n763), .ZN(n566) );
  OR2_X1 U439 ( .A1(n536), .A2(n535), .ZN(n763) );
  OR2_X1 U440 ( .A1(n534), .A2(n533), .ZN(n535) );
  OR2_X1 U441 ( .A1(n532), .A2(n531), .ZN(n533) );
  OR2_X1 U442 ( .A1(in[115]), .A2(in[110]), .ZN(n531) );
  OR2_X1 U443 ( .A1(in[125]), .A2(in[117]), .ZN(n532) );
  OR2_X1 U444 ( .A1(n530), .A2(n529), .ZN(n534) );
  OR2_X1 U445 ( .A1(in[180]), .A2(in[128]), .ZN(n529) );
  OR2_X1 U446 ( .A1(in[205]), .A2(in[201]), .ZN(n530) );
  OR2_X1 U447 ( .A1(n528), .A2(n527), .ZN(n536) );
  OR2_X1 U448 ( .A1(n526), .A2(n525), .ZN(n527) );
  OR2_X1 U449 ( .A1(in[244]), .A2(in[239]), .ZN(n525) );
  OR2_X1 U450 ( .A1(in[95]), .A2(in[83]), .ZN(n526) );
  OR2_X1 U451 ( .A1(n524), .A2(n523), .ZN(n528) );
  OR2_X1 U452 ( .A1(in_24), .A2(in[97]), .ZN(n523) );
  OR2_X1 U453 ( .A1(in_33), .A2(in_27), .ZN(n524) );
  OR2_X1 U454 ( .A1(n522), .A2(n521), .ZN(n568) );
  OR2_X1 U455 ( .A1(in[145]), .A2(in[126]), .ZN(n521) );
  OR2_X1 U456 ( .A1(in[169]), .A2(n520), .ZN(n522) );
  OR2_X1 U457 ( .A1(in[221]), .A2(in[172]), .ZN(n520) );
  OR2_X1 U458 ( .A1(n519), .A2(n518), .ZN(n570) );
  OR2_X1 U459 ( .A1(n517), .A2(n516), .ZN(n518) );
  OR2_X1 U460 ( .A1(in[241]), .A2(in[224]), .ZN(n516) );
  OR2_X1 U461 ( .A1(in[86]), .A2(n515), .ZN(n517) );
  OR2_X1 U462 ( .A1(in_43), .A2(in_34), .ZN(n515) );
  OR2_X1 U463 ( .A1(n514), .A2(n513), .ZN(n519) );
  OR2_X1 U464 ( .A1(in_65), .A2(in_51), .ZN(n513) );
  OR2_X1 U465 ( .A1(in_75), .A2(n512), .ZN(n514) );
  OR2_X1 U466 ( .A1(in_81), .A2(in_77), .ZN(n512) );
  OR2_X1 U467 ( .A1(n511), .A2(n510), .ZN(n778) );
  OR2_X1 U468 ( .A1(n509), .A2(n508), .ZN(n510) );
  OR2_X1 U469 ( .A1(n507), .A2(n506), .ZN(n508) );
  OR2_X1 U470 ( .A1(in[107]), .A2(in[101]), .ZN(n506) );
  OR2_X1 U471 ( .A1(in[139]), .A2(in[132]), .ZN(n507) );
  OR2_X1 U472 ( .A1(n505), .A2(n504), .ZN(n509) );
  OR2_X1 U473 ( .A1(in[146]), .A2(in[141]), .ZN(n504) );
  OR2_X1 U474 ( .A1(in[203]), .A2(in[179]), .ZN(n505) );
  OR2_X1 U475 ( .A1(n503), .A2(n502), .ZN(n511) );
  OR2_X1 U476 ( .A1(n501), .A2(n500), .ZN(n502) );
  OR2_X1 U477 ( .A1(in[243]), .A2(in[222]), .ZN(n500) );
  OR2_X1 U478 ( .A1(in[251]), .A2(in[250]), .ZN(n501) );
  OR2_X1 U479 ( .A1(n499), .A2(n498), .ZN(n503) );
  OR2_X1 U480 ( .A1(in_37), .A2(in_19), .ZN(n498) );
  OR2_X1 U481 ( .A1(in_78), .A2(in_6), .ZN(n499) );
  OR2_X1 U482 ( .A1(n497), .A2(n496), .ZN(n603) );
  OR2_X1 U483 ( .A1(in[112]), .A2(in[102]), .ZN(n496) );
  OR2_X1 U484 ( .A1(in[123]), .A2(n495), .ZN(n497) );
  OR2_X1 U485 ( .A1(in[143]), .A2(in[130]), .ZN(n495) );
  OR2_X1 U486 ( .A1(n494), .A2(n493), .ZN(n605) );
  OR2_X1 U487 ( .A1(n492), .A2(n491), .ZN(n493) );
  OR2_X1 U488 ( .A1(in[216]), .A2(in[213]), .ZN(n491) );
  OR2_X1 U489 ( .A1(in[227]), .A2(n490), .ZN(n492) );
  OR2_X1 U490 ( .A1(in_0), .A2(in[248]), .ZN(n490) );
  OR2_X1 U491 ( .A1(n489), .A2(n488), .ZN(n494) );
  OR2_X1 U492 ( .A1(in_46), .A2(in_44), .ZN(n488) );
  OR2_X1 U493 ( .A1(in_50), .A2(n487), .ZN(n489) );
  OR2_X1 U494 ( .A1(in_9), .A2(in_80), .ZN(n487) );
endmodule
//done