`timescale 1ns / 1ps

module AND2_X1( A1, A2, ZN );
  input wire A1;
  input wire A2;
  //input_done

  output wire ZN;
  //output_done

  //wire_done

  assign ZN = A1 & A2;
endmodule


module OR2_X1( A1, A2, ZN );
  input wire A1;
  input wire A2;
  //input_done

  output wire ZN;
  //output_done

  //wire_done

  assign ZN = A1 | A2;
endmodule

module CD2_0 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD4_0 ( a, abar, b, bbar, y, ybar );

  input wire [3:0] a;
  input wire [3:0] b;
  input wire [3:0] abar;
  input wire [3:0] bbar;
//input_done

  output wire [15:0] y;
  output wire [15:0] ybar;
//output_done

//wire_done

  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]) );
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]) );
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]) );
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]) );
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]) );
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]) );
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]) );
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]) );
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]) );
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]) );
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]) );
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]) );
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]) );
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]) );
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]) );
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]) );
endmodule

module CD16_0 ( a, abar, b, bbar, y, ybar );

  input wire [15:0] a;
  input wire [15:0] b;
  input wire [15:0] abar;
  input wire [15:0] bbar;
//input_done

  output wire [255:0] y;
  output wire [255:0] ybar;
//output_done

//wire_done

  AND2_X1 U1 ( .A1(b[9]), .A2(a[0]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[9]), .A2(abar[0]), .ZN(ybar[9]) );
  AND2_X1 U2 ( .A1(b[3]), .A2(a[6]), .ZN(y[99]) );
  OR2_X1 U2bar ( .A1(bbar[3]), .A2(abar[6]), .ZN(ybar[99]) );
  AND2_X1 U3 ( .A1(b[2]), .A2(a[6]), .ZN(y[98]) );
  OR2_X1 U3bar ( .A1(bbar[2]), .A2(abar[6]), .ZN(ybar[98]) );
  AND2_X1 U4 ( .A1(b[1]), .A2(a[6]), .ZN(y[97]) );
  OR2_X1 U4bar ( .A1(bbar[1]), .A2(abar[6]), .ZN(ybar[97]) );
  AND2_X1 U5 ( .A1(b[0]), .A2(a[6]), .ZN(y[96]) );
  OR2_X1 U5bar ( .A1(bbar[0]), .A2(abar[6]), .ZN(ybar[96]) );
  AND2_X1 U6 ( .A1(b[15]), .A2(a[5]), .ZN(y[95]) );
  OR2_X1 U6bar ( .A1(bbar[15]), .A2(abar[5]), .ZN(ybar[95]) );
  AND2_X1 U7 ( .A1(b[14]), .A2(a[5]), .ZN(y[94]) );
  OR2_X1 U7bar ( .A1(bbar[14]), .A2(abar[5]), .ZN(ybar[94]) );
  AND2_X1 U8 ( .A1(b[13]), .A2(a[5]), .ZN(y[93]) );
  OR2_X1 U8bar ( .A1(bbar[13]), .A2(abar[5]), .ZN(ybar[93]) );
  AND2_X1 U9 ( .A1(b[12]), .A2(a[5]), .ZN(y[92]) );
  OR2_X1 U9bar ( .A1(bbar[12]), .A2(abar[5]), .ZN(ybar[92]) );
  AND2_X1 U10 ( .A1(b[11]), .A2(a[5]), .ZN(y[91]) );
  OR2_X1 U10bar ( .A1(bbar[11]), .A2(abar[5]), .ZN(ybar[91]) );
  AND2_X1 U11 ( .A1(b[10]), .A2(a[5]), .ZN(y[90]) );
  OR2_X1 U11bar ( .A1(bbar[10]), .A2(abar[5]), .ZN(ybar[90]) );
  AND2_X1 U12 ( .A1(b[8]), .A2(a[0]), .ZN(y[8]) );
  OR2_X1 U12bar ( .A1(bbar[8]), .A2(abar[0]), .ZN(ybar[8]) );
  AND2_X1 U13 ( .A1(a[5]), .A2(b[9]), .ZN(y[89]) );
  OR2_X1 U13bar ( .A1(abar[5]), .A2(bbar[9]), .ZN(ybar[89]) );
  AND2_X1 U14 ( .A1(b[8]), .A2(a[5]), .ZN(y[88]) );
  OR2_X1 U14bar ( .A1(bbar[8]), .A2(abar[5]), .ZN(ybar[88]) );
  AND2_X1 U15 ( .A1(b[7]), .A2(a[5]), .ZN(y[87]) );
  OR2_X1 U15bar ( .A1(bbar[7]), .A2(abar[5]), .ZN(ybar[87]) );
  AND2_X1 U16 ( .A1(b[6]), .A2(a[5]), .ZN(y[86]) );
  OR2_X1 U16bar ( .A1(bbar[6]), .A2(abar[5]), .ZN(ybar[86]) );
  AND2_X1 U17 ( .A1(b[5]), .A2(a[5]), .ZN(y[85]) );
  OR2_X1 U17bar ( .A1(bbar[5]), .A2(abar[5]), .ZN(ybar[85]) );
  AND2_X1 U18 ( .A1(b[4]), .A2(a[5]), .ZN(y[84]) );
  OR2_X1 U18bar ( .A1(bbar[4]), .A2(abar[5]), .ZN(ybar[84]) );
  AND2_X1 U19 ( .A1(a[5]), .A2(b[3]), .ZN(y[83]) );
  OR2_X1 U19bar ( .A1(abar[5]), .A2(bbar[3]), .ZN(ybar[83]) );
  AND2_X1 U20 ( .A1(a[5]), .A2(b[2]), .ZN(y[82]) );
  OR2_X1 U20bar ( .A1(abar[5]), .A2(bbar[2]), .ZN(ybar[82]) );
  AND2_X1 U21 ( .A1(a[5]), .A2(b[1]), .ZN(y[81]) );
  OR2_X1 U21bar ( .A1(abar[5]), .A2(bbar[1]), .ZN(ybar[81]) );
  AND2_X1 U22 ( .A1(a[5]), .A2(b[0]), .ZN(y[80]) );
  OR2_X1 U22bar ( .A1(abar[5]), .A2(bbar[0]), .ZN(ybar[80]) );
  AND2_X1 U23 ( .A1(b[7]), .A2(a[0]), .ZN(y[7]) );
  OR2_X1 U23bar ( .A1(bbar[7]), .A2(abar[0]), .ZN(ybar[7]) );
  AND2_X1 U24 ( .A1(a[4]), .A2(b[15]), .ZN(y[79]) );
  OR2_X1 U24bar ( .A1(abar[4]), .A2(bbar[15]), .ZN(ybar[79]) );
  AND2_X1 U25 ( .A1(a[4]), .A2(b[14]), .ZN(y[78]) );
  OR2_X1 U25bar ( .A1(abar[4]), .A2(bbar[14]), .ZN(ybar[78]) );
  AND2_X1 U26 ( .A1(a[4]), .A2(b[13]), .ZN(y[77]) );
  OR2_X1 U26bar ( .A1(abar[4]), .A2(bbar[13]), .ZN(ybar[77]) );
  AND2_X1 U27 ( .A1(a[4]), .A2(b[12]), .ZN(y[76]) );
  OR2_X1 U27bar ( .A1(abar[4]), .A2(bbar[12]), .ZN(ybar[76]) );
  AND2_X1 U28 ( .A1(a[4]), .A2(b[11]), .ZN(y[75]) );
  OR2_X1 U28bar ( .A1(abar[4]), .A2(bbar[11]), .ZN(ybar[75]) );
  AND2_X1 U29 ( .A1(a[4]), .A2(b[10]), .ZN(y[74]) );
  OR2_X1 U29bar ( .A1(abar[4]), .A2(bbar[10]), .ZN(ybar[74]) );
  AND2_X1 U30 ( .A1(a[4]), .A2(b[9]), .ZN(y[73]) );
  OR2_X1 U30bar ( .A1(abar[4]), .A2(bbar[9]), .ZN(ybar[73]) );
  AND2_X1 U31 ( .A1(a[4]), .A2(b[8]), .ZN(y[72]) );
  OR2_X1 U31bar ( .A1(abar[4]), .A2(bbar[8]), .ZN(ybar[72]) );
  AND2_X1 U32 ( .A1(a[4]), .A2(b[7]), .ZN(y[71]) );
  OR2_X1 U32bar ( .A1(abar[4]), .A2(bbar[7]), .ZN(ybar[71]) );
  AND2_X1 U33 ( .A1(a[4]), .A2(b[6]), .ZN(y[70]) );
  OR2_X1 U33bar ( .A1(abar[4]), .A2(bbar[6]), .ZN(ybar[70]) );
  AND2_X1 U34 ( .A1(b[6]), .A2(a[0]), .ZN(y[6]) );
  OR2_X1 U34bar ( .A1(bbar[6]), .A2(abar[0]), .ZN(ybar[6]) );
  AND2_X1 U35 ( .A1(a[4]), .A2(b[5]), .ZN(y[69]) );
  OR2_X1 U35bar ( .A1(abar[4]), .A2(bbar[5]), .ZN(ybar[69]) );
  AND2_X1 U36 ( .A1(a[4]), .A2(b[4]), .ZN(y[68]) );
  OR2_X1 U36bar ( .A1(abar[4]), .A2(bbar[4]), .ZN(ybar[68]) );
  AND2_X1 U37 ( .A1(a[4]), .A2(b[3]), .ZN(y[67]) );
  OR2_X1 U37bar ( .A1(abar[4]), .A2(bbar[3]), .ZN(ybar[67]) );
  AND2_X1 U38 ( .A1(a[4]), .A2(b[2]), .ZN(y[66]) );
  OR2_X1 U38bar ( .A1(abar[4]), .A2(bbar[2]), .ZN(ybar[66]) );
  AND2_X1 U39 ( .A1(a[4]), .A2(b[1]), .ZN(y[65]) );
  OR2_X1 U39bar ( .A1(abar[4]), .A2(bbar[1]), .ZN(ybar[65]) );
  AND2_X1 U40 ( .A1(a[4]), .A2(b[0]), .ZN(y[64]) );
  OR2_X1 U40bar ( .A1(abar[4]), .A2(bbar[0]), .ZN(ybar[64]) );
  AND2_X1 U41 ( .A1(a[3]), .A2(b[15]), .ZN(y[63]) );
  OR2_X1 U41bar ( .A1(abar[3]), .A2(bbar[15]), .ZN(ybar[63]) );
  AND2_X1 U42 ( .A1(a[3]), .A2(b[14]), .ZN(y[62]) );
  OR2_X1 U42bar ( .A1(abar[3]), .A2(bbar[14]), .ZN(ybar[62]) );
  AND2_X1 U43 ( .A1(a[3]), .A2(b[13]), .ZN(y[61]) );
  OR2_X1 U43bar ( .A1(abar[3]), .A2(bbar[13]), .ZN(ybar[61]) );
  AND2_X1 U44 ( .A1(a[3]), .A2(b[12]), .ZN(y[60]) );
  OR2_X1 U44bar ( .A1(abar[3]), .A2(bbar[12]), .ZN(ybar[60]) );
  AND2_X1 U45 ( .A1(b[5]), .A2(a[0]), .ZN(y[5]) );
  OR2_X1 U45bar ( .A1(bbar[5]), .A2(abar[0]), .ZN(ybar[5]) );
  AND2_X1 U46 ( .A1(a[3]), .A2(b[11]), .ZN(y[59]) );
  OR2_X1 U46bar ( .A1(abar[3]), .A2(bbar[11]), .ZN(ybar[59]) );
  AND2_X1 U47 ( .A1(a[3]), .A2(b[10]), .ZN(y[58]) );
  OR2_X1 U47bar ( .A1(abar[3]), .A2(bbar[10]), .ZN(ybar[58]) );
  AND2_X1 U48 ( .A1(a[3]), .A2(b[9]), .ZN(y[57]) );
  OR2_X1 U48bar ( .A1(abar[3]), .A2(bbar[9]), .ZN(ybar[57]) );
  AND2_X1 U49 ( .A1(a[3]), .A2(b[8]), .ZN(y[56]) );
  OR2_X1 U49bar ( .A1(abar[3]), .A2(bbar[8]), .ZN(ybar[56]) );
  AND2_X1 U50 ( .A1(a[3]), .A2(b[7]), .ZN(y[55]) );
  OR2_X1 U50bar ( .A1(abar[3]), .A2(bbar[7]), .ZN(ybar[55]) );
  AND2_X1 U51 ( .A1(a[3]), .A2(b[6]), .ZN(y[54]) );
  OR2_X1 U51bar ( .A1(abar[3]), .A2(bbar[6]), .ZN(ybar[54]) );
  AND2_X1 U52 ( .A1(a[3]), .A2(b[5]), .ZN(y[53]) );
  OR2_X1 U52bar ( .A1(abar[3]), .A2(bbar[5]), .ZN(ybar[53]) );
  AND2_X1 U53 ( .A1(a[3]), .A2(b[4]), .ZN(y[52]) );
  OR2_X1 U53bar ( .A1(abar[3]), .A2(bbar[4]), .ZN(ybar[52]) );
  AND2_X1 U54 ( .A1(a[3]), .A2(b[3]), .ZN(y[51]) );
  OR2_X1 U54bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[51]) );
  AND2_X1 U55 ( .A1(a[3]), .A2(b[2]), .ZN(y[50]) );
  OR2_X1 U55bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[50]) );
  AND2_X1 U56 ( .A1(b[4]), .A2(a[0]), .ZN(y[4]) );
  OR2_X1 U56bar ( .A1(bbar[4]), .A2(abar[0]), .ZN(ybar[4]) );
  AND2_X1 U57 ( .A1(a[3]), .A2(b[1]), .ZN(y[49]) );
  OR2_X1 U57bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[49]) );
  AND2_X1 U58 ( .A1(a[3]), .A2(b[0]), .ZN(y[48]) );
  OR2_X1 U58bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[48]) );
  AND2_X1 U59 ( .A1(a[2]), .A2(b[15]), .ZN(y[47]) );
  OR2_X1 U59bar ( .A1(abar[2]), .A2(bbar[15]), .ZN(ybar[47]) );
  AND2_X1 U60 ( .A1(a[2]), .A2(b[14]), .ZN(y[46]) );
  OR2_X1 U60bar ( .A1(abar[2]), .A2(bbar[14]), .ZN(ybar[46]) );
  AND2_X1 U61 ( .A1(a[2]), .A2(b[13]), .ZN(y[45]) );
  OR2_X1 U61bar ( .A1(abar[2]), .A2(bbar[13]), .ZN(ybar[45]) );
  AND2_X1 U62 ( .A1(a[2]), .A2(b[12]), .ZN(y[44]) );
  OR2_X1 U62bar ( .A1(abar[2]), .A2(bbar[12]), .ZN(ybar[44]) );
  AND2_X1 U63 ( .A1(a[2]), .A2(b[11]), .ZN(y[43]) );
  OR2_X1 U63bar ( .A1(abar[2]), .A2(bbar[11]), .ZN(ybar[43]) );
  AND2_X1 U64 ( .A1(a[2]), .A2(b[10]), .ZN(y[42]) );
  OR2_X1 U64bar ( .A1(abar[2]), .A2(bbar[10]), .ZN(ybar[42]) );
  AND2_X1 U65 ( .A1(a[2]), .A2(b[9]), .ZN(y[41]) );
  OR2_X1 U65bar ( .A1(abar[2]), .A2(bbar[9]), .ZN(ybar[41]) );
  AND2_X1 U66 ( .A1(a[2]), .A2(b[8]), .ZN(y[40]) );
  OR2_X1 U66bar ( .A1(abar[2]), .A2(bbar[8]), .ZN(ybar[40]) );
  AND2_X1 U67 ( .A1(b[3]), .A2(a[0]), .ZN(y[3]) );
  OR2_X1 U67bar ( .A1(bbar[3]), .A2(abar[0]), .ZN(ybar[3]) );
  AND2_X1 U68 ( .A1(a[2]), .A2(b[7]), .ZN(y[39]) );
  OR2_X1 U68bar ( .A1(abar[2]), .A2(bbar[7]), .ZN(ybar[39]) );
  AND2_X1 U69 ( .A1(a[2]), .A2(b[6]), .ZN(y[38]) );
  OR2_X1 U69bar ( .A1(abar[2]), .A2(bbar[6]), .ZN(ybar[38]) );
  AND2_X1 U70 ( .A1(a[2]), .A2(b[5]), .ZN(y[37]) );
  OR2_X1 U70bar ( .A1(abar[2]), .A2(bbar[5]), .ZN(ybar[37]) );
  AND2_X1 U71 ( .A1(a[2]), .A2(b[4]), .ZN(y[36]) );
  OR2_X1 U71bar ( .A1(abar[2]), .A2(bbar[4]), .ZN(ybar[36]) );
  AND2_X1 U72 ( .A1(a[2]), .A2(b[3]), .ZN(y[35]) );
  OR2_X1 U72bar ( .A1(abar[2]), .A2(bbar[3]), .ZN(ybar[35]) );
  AND2_X1 U73 ( .A1(a[2]), .A2(b[2]), .ZN(y[34]) );
  OR2_X1 U73bar ( .A1(abar[2]), .A2(bbar[2]), .ZN(ybar[34]) );
  AND2_X1 U74 ( .A1(a[2]), .A2(b[1]), .ZN(y[33]) );
  OR2_X1 U74bar ( .A1(abar[2]), .A2(bbar[1]), .ZN(ybar[33]) );
  AND2_X1 U75 ( .A1(a[2]), .A2(b[0]), .ZN(y[32]) );
  OR2_X1 U75bar ( .A1(abar[2]), .A2(bbar[0]), .ZN(ybar[32]) );
  AND2_X1 U76 ( .A1(a[1]), .A2(b[15]), .ZN(y[31]) );
  OR2_X1 U76bar ( .A1(abar[1]), .A2(bbar[15]), .ZN(ybar[31]) );
  AND2_X1 U77 ( .A1(a[1]), .A2(b[14]), .ZN(y[30]) );
  OR2_X1 U77bar ( .A1(abar[1]), .A2(bbar[14]), .ZN(ybar[30]) );
  AND2_X1 U78 ( .A1(b[2]), .A2(a[0]), .ZN(y[2]) );
  OR2_X1 U78bar ( .A1(bbar[2]), .A2(abar[0]), .ZN(ybar[2]) );
  AND2_X1 U79 ( .A1(a[1]), .A2(b[13]), .ZN(y[29]) );
  OR2_X1 U79bar ( .A1(abar[1]), .A2(bbar[13]), .ZN(ybar[29]) );
  AND2_X1 U80 ( .A1(a[1]), .A2(b[12]), .ZN(y[28]) );
  OR2_X1 U80bar ( .A1(abar[1]), .A2(bbar[12]), .ZN(ybar[28]) );
  AND2_X1 U81 ( .A1(a[1]), .A2(b[11]), .ZN(y[27]) );
  OR2_X1 U81bar ( .A1(abar[1]), .A2(bbar[11]), .ZN(ybar[27]) );
  AND2_X1 U82 ( .A1(a[1]), .A2(b[10]), .ZN(y[26]) );
  OR2_X1 U82bar ( .A1(abar[1]), .A2(bbar[10]), .ZN(ybar[26]) );
  AND2_X1 U83 ( .A1(a[1]), .A2(b[9]), .ZN(y[25]) );
  OR2_X1 U83bar ( .A1(abar[1]), .A2(bbar[9]), .ZN(ybar[25]) );
  AND2_X1 U84 ( .A1(a[15]), .A2(b[15]), .ZN(y[255]) );
  OR2_X1 U84bar ( .A1(abar[15]), .A2(bbar[15]), .ZN(ybar[255]) );
  AND2_X1 U85 ( .A1(a[15]), .A2(b[14]), .ZN(y[254]) );
  OR2_X1 U85bar ( .A1(abar[15]), .A2(bbar[14]), .ZN(ybar[254]) );
  AND2_X1 U86 ( .A1(a[15]), .A2(b[13]), .ZN(y[253]) );
  OR2_X1 U86bar ( .A1(abar[15]), .A2(bbar[13]), .ZN(ybar[253]) );
  AND2_X1 U87 ( .A1(a[15]), .A2(b[12]), .ZN(y[252]) );
  OR2_X1 U87bar ( .A1(abar[15]), .A2(bbar[12]), .ZN(ybar[252]) );
  AND2_X1 U88 ( .A1(a[15]), .A2(b[11]), .ZN(y[251]) );
  OR2_X1 U88bar ( .A1(abar[15]), .A2(bbar[11]), .ZN(ybar[251]) );
  AND2_X1 U89 ( .A1(a[15]), .A2(b[10]), .ZN(y[250]) );
  OR2_X1 U89bar ( .A1(abar[15]), .A2(bbar[10]), .ZN(ybar[250]) );
  AND2_X1 U90 ( .A1(a[1]), .A2(b[8]), .ZN(y[24]) );
  OR2_X1 U90bar ( .A1(abar[1]), .A2(bbar[8]), .ZN(ybar[24]) );
  AND2_X1 U91 ( .A1(a[15]), .A2(b[9]), .ZN(y[249]) );
  OR2_X1 U91bar ( .A1(abar[15]), .A2(bbar[9]), .ZN(ybar[249]) );
  AND2_X1 U92 ( .A1(a[15]), .A2(b[8]), .ZN(y[248]) );
  OR2_X1 U92bar ( .A1(abar[15]), .A2(bbar[8]), .ZN(ybar[248]) );
  AND2_X1 U93 ( .A1(a[15]), .A2(b[7]), .ZN(y[247]) );
  OR2_X1 U93bar ( .A1(abar[15]), .A2(bbar[7]), .ZN(ybar[247]) );
  AND2_X1 U94 ( .A1(a[15]), .A2(b[6]), .ZN(y[246]) );
  OR2_X1 U94bar ( .A1(abar[15]), .A2(bbar[6]), .ZN(ybar[246]) );
  AND2_X1 U95 ( .A1(a[15]), .A2(b[5]), .ZN(y[245]) );
  OR2_X1 U95bar ( .A1(abar[15]), .A2(bbar[5]), .ZN(ybar[245]) );
  AND2_X1 U96 ( .A1(a[15]), .A2(b[4]), .ZN(y[244]) );
  OR2_X1 U96bar ( .A1(abar[15]), .A2(bbar[4]), .ZN(ybar[244]) );
  AND2_X1 U97 ( .A1(a[15]), .A2(b[3]), .ZN(y[243]) );
  OR2_X1 U97bar ( .A1(abar[15]), .A2(bbar[3]), .ZN(ybar[243]) );
  AND2_X1 U98 ( .A1(a[15]), .A2(b[2]), .ZN(y[242]) );
  OR2_X1 U98bar ( .A1(abar[15]), .A2(bbar[2]), .ZN(ybar[242]) );
  AND2_X1 U99 ( .A1(a[15]), .A2(b[1]), .ZN(y[241]) );
  OR2_X1 U99bar ( .A1(abar[15]), .A2(bbar[1]), .ZN(ybar[241]) );
  AND2_X1 U100 ( .A1(a[15]), .A2(b[0]), .ZN(y[240]) );
  OR2_X1 U100bar ( .A1(abar[15]), .A2(bbar[0]), .ZN(ybar[240]) );
  AND2_X1 U101 ( .A1(a[1]), .A2(b[7]), .ZN(y[23]) );
  OR2_X1 U101bar ( .A1(abar[1]), .A2(bbar[7]), .ZN(ybar[23]) );
  AND2_X1 U102 ( .A1(a[14]), .A2(b[15]), .ZN(y[239]) );
  OR2_X1 U102bar ( .A1(abar[14]), .A2(bbar[15]), .ZN(ybar[239]) );
  AND2_X1 U103 ( .A1(a[14]), .A2(b[14]), .ZN(y[238]) );
  OR2_X1 U103bar ( .A1(abar[14]), .A2(bbar[14]), .ZN(ybar[238]) );
  AND2_X1 U104 ( .A1(a[14]), .A2(b[13]), .ZN(y[237]) );
  OR2_X1 U104bar ( .A1(abar[14]), .A2(bbar[13]), .ZN(ybar[237]) );
  AND2_X1 U105 ( .A1(a[14]), .A2(b[12]), .ZN(y[236]) );
  OR2_X1 U105bar ( .A1(abar[14]), .A2(bbar[12]), .ZN(ybar[236]) );
  AND2_X1 U106 ( .A1(a[14]), .A2(b[11]), .ZN(y[235]) );
  OR2_X1 U106bar ( .A1(abar[14]), .A2(bbar[11]), .ZN(ybar[235]) );
  AND2_X1 U107 ( .A1(a[14]), .A2(b[10]), .ZN(y[234]) );
  OR2_X1 U107bar ( .A1(abar[14]), .A2(bbar[10]), .ZN(ybar[234]) );
  AND2_X1 U108 ( .A1(a[14]), .A2(b[9]), .ZN(y[233]) );
  OR2_X1 U108bar ( .A1(abar[14]), .A2(bbar[9]), .ZN(ybar[233]) );
  AND2_X1 U109 ( .A1(a[14]), .A2(b[8]), .ZN(y[232]) );
  OR2_X1 U109bar ( .A1(abar[14]), .A2(bbar[8]), .ZN(ybar[232]) );
  AND2_X1 U110 ( .A1(a[14]), .A2(b[7]), .ZN(y[231]) );
  OR2_X1 U110bar ( .A1(abar[14]), .A2(bbar[7]), .ZN(ybar[231]) );
  AND2_X1 U111 ( .A1(a[14]), .A2(b[6]), .ZN(y[230]) );
  OR2_X1 U111bar ( .A1(abar[14]), .A2(bbar[6]), .ZN(ybar[230]) );
  AND2_X1 U112 ( .A1(a[1]), .A2(b[6]), .ZN(y[22]) );
  OR2_X1 U112bar ( .A1(abar[1]), .A2(bbar[6]), .ZN(ybar[22]) );
  AND2_X1 U113 ( .A1(a[14]), .A2(b[5]), .ZN(y[229]) );
  OR2_X1 U113bar ( .A1(abar[14]), .A2(bbar[5]), .ZN(ybar[229]) );
  AND2_X1 U114 ( .A1(a[14]), .A2(b[4]), .ZN(y[228]) );
  OR2_X1 U114bar ( .A1(abar[14]), .A2(bbar[4]), .ZN(ybar[228]) );
  AND2_X1 U115 ( .A1(a[14]), .A2(b[3]), .ZN(y[227]) );
  OR2_X1 U115bar ( .A1(abar[14]), .A2(bbar[3]), .ZN(ybar[227]) );
  AND2_X1 U116 ( .A1(a[14]), .A2(b[2]), .ZN(y[226]) );
  OR2_X1 U116bar ( .A1(abar[14]), .A2(bbar[2]), .ZN(ybar[226]) );
  AND2_X1 U117 ( .A1(a[14]), .A2(b[1]), .ZN(y[225]) );
  OR2_X1 U117bar ( .A1(abar[14]), .A2(bbar[1]), .ZN(ybar[225]) );
  AND2_X1 U118 ( .A1(a[14]), .A2(b[0]), .ZN(y[224]) );
  OR2_X1 U118bar ( .A1(abar[14]), .A2(bbar[0]), .ZN(ybar[224]) );
  AND2_X1 U119 ( .A1(a[13]), .A2(b[15]), .ZN(y[223]) );
  OR2_X1 U119bar ( .A1(abar[13]), .A2(bbar[15]), .ZN(ybar[223]) );
  AND2_X1 U120 ( .A1(a[13]), .A2(b[14]), .ZN(y[222]) );
  OR2_X1 U120bar ( .A1(abar[13]), .A2(bbar[14]), .ZN(ybar[222]) );
  AND2_X1 U121 ( .A1(a[13]), .A2(b[13]), .ZN(y[221]) );
  OR2_X1 U121bar ( .A1(abar[13]), .A2(bbar[13]), .ZN(ybar[221]) );
  AND2_X1 U122 ( .A1(a[13]), .A2(b[12]), .ZN(y[220]) );
  OR2_X1 U122bar ( .A1(abar[13]), .A2(bbar[12]), .ZN(ybar[220]) );
  AND2_X1 U123 ( .A1(a[1]), .A2(b[5]), .ZN(y[21]) );
  OR2_X1 U123bar ( .A1(abar[1]), .A2(bbar[5]), .ZN(ybar[21]) );
  AND2_X1 U124 ( .A1(a[13]), .A2(b[11]), .ZN(y[219]) );
  OR2_X1 U124bar ( .A1(abar[13]), .A2(bbar[11]), .ZN(ybar[219]) );
  AND2_X1 U125 ( .A1(a[13]), .A2(b[10]), .ZN(y[218]) );
  OR2_X1 U125bar ( .A1(abar[13]), .A2(bbar[10]), .ZN(ybar[218]) );
  AND2_X1 U126 ( .A1(a[13]), .A2(b[9]), .ZN(y[217]) );
  OR2_X1 U126bar ( .A1(abar[13]), .A2(bbar[9]), .ZN(ybar[217]) );
  AND2_X1 U127 ( .A1(a[13]), .A2(b[8]), .ZN(y[216]) );
  OR2_X1 U127bar ( .A1(abar[13]), .A2(bbar[8]), .ZN(ybar[216]) );
  AND2_X1 U128 ( .A1(a[13]), .A2(b[7]), .ZN(y[215]) );
  OR2_X1 U128bar ( .A1(abar[13]), .A2(bbar[7]), .ZN(ybar[215]) );
  AND2_X1 U129 ( .A1(a[13]), .A2(b[6]), .ZN(y[214]) );
  OR2_X1 U129bar ( .A1(abar[13]), .A2(bbar[6]), .ZN(ybar[214]) );
  AND2_X1 U130 ( .A1(a[13]), .A2(b[5]), .ZN(y[213]) );
  OR2_X1 U130bar ( .A1(abar[13]), .A2(bbar[5]), .ZN(ybar[213]) );
  AND2_X1 U131 ( .A1(a[13]), .A2(b[4]), .ZN(y[212]) );
  OR2_X1 U131bar ( .A1(abar[13]), .A2(bbar[4]), .ZN(ybar[212]) );
  AND2_X1 U132 ( .A1(a[13]), .A2(b[3]), .ZN(y[211]) );
  OR2_X1 U132bar ( .A1(abar[13]), .A2(bbar[3]), .ZN(ybar[211]) );
  AND2_X1 U133 ( .A1(a[13]), .A2(b[2]), .ZN(y[210]) );
  OR2_X1 U133bar ( .A1(abar[13]), .A2(bbar[2]), .ZN(ybar[210]) );
  AND2_X1 U134 ( .A1(a[1]), .A2(b[4]), .ZN(y[20]) );
  OR2_X1 U134bar ( .A1(abar[1]), .A2(bbar[4]), .ZN(ybar[20]) );
  AND2_X1 U135 ( .A1(a[13]), .A2(b[1]), .ZN(y[209]) );
  OR2_X1 U135bar ( .A1(abar[13]), .A2(bbar[1]), .ZN(ybar[209]) );
  AND2_X1 U136 ( .A1(a[13]), .A2(b[0]), .ZN(y[208]) );
  OR2_X1 U136bar ( .A1(abar[13]), .A2(bbar[0]), .ZN(ybar[208]) );
  AND2_X1 U137 ( .A1(a[12]), .A2(b[15]), .ZN(y[207]) );
  OR2_X1 U137bar ( .A1(abar[12]), .A2(bbar[15]), .ZN(ybar[207]) );
  AND2_X1 U138 ( .A1(a[12]), .A2(b[14]), .ZN(y[206]) );
  OR2_X1 U138bar ( .A1(abar[12]), .A2(bbar[14]), .ZN(ybar[206]) );
  AND2_X1 U139 ( .A1(a[12]), .A2(b[13]), .ZN(y[205]) );
  OR2_X1 U139bar ( .A1(abar[12]), .A2(bbar[13]), .ZN(ybar[205]) );
  AND2_X1 U140 ( .A1(a[12]), .A2(b[12]), .ZN(y[204]) );
  OR2_X1 U140bar ( .A1(abar[12]), .A2(bbar[12]), .ZN(ybar[204]) );
  AND2_X1 U141 ( .A1(a[12]), .A2(b[11]), .ZN(y[203]) );
  OR2_X1 U141bar ( .A1(abar[12]), .A2(bbar[11]), .ZN(ybar[203]) );
  AND2_X1 U142 ( .A1(a[12]), .A2(b[10]), .ZN(y[202]) );
  OR2_X1 U142bar ( .A1(abar[12]), .A2(bbar[10]), .ZN(ybar[202]) );
  AND2_X1 U143 ( .A1(a[12]), .A2(b[9]), .ZN(y[201]) );
  OR2_X1 U143bar ( .A1(abar[12]), .A2(bbar[9]), .ZN(ybar[201]) );
  AND2_X1 U144 ( .A1(a[12]), .A2(b[8]), .ZN(y[200]) );
  OR2_X1 U144bar ( .A1(abar[12]), .A2(bbar[8]), .ZN(ybar[200]) );
  AND2_X1 U145 ( .A1(b[1]), .A2(a[0]), .ZN(y[1]) );
  OR2_X1 U145bar ( .A1(bbar[1]), .A2(abar[0]), .ZN(ybar[1]) );
  AND2_X1 U146 ( .A1(a[1]), .A2(b[3]), .ZN(y[19]) );
  OR2_X1 U146bar ( .A1(abar[1]), .A2(bbar[3]), .ZN(ybar[19]) );
  AND2_X1 U147 ( .A1(a[12]), .A2(b[7]), .ZN(y[199]) );
  OR2_X1 U147bar ( .A1(abar[12]), .A2(bbar[7]), .ZN(ybar[199]) );
  AND2_X1 U148 ( .A1(a[12]), .A2(b[6]), .ZN(y[198]) );
  OR2_X1 U148bar ( .A1(abar[12]), .A2(bbar[6]), .ZN(ybar[198]) );
  AND2_X1 U149 ( .A1(a[12]), .A2(b[5]), .ZN(y[197]) );
  OR2_X1 U149bar ( .A1(abar[12]), .A2(bbar[5]), .ZN(ybar[197]) );
  AND2_X1 U150 ( .A1(a[12]), .A2(b[4]), .ZN(y[196]) );
  OR2_X1 U150bar ( .A1(abar[12]), .A2(bbar[4]), .ZN(ybar[196]) );
  AND2_X1 U151 ( .A1(a[12]), .A2(b[3]), .ZN(y[195]) );
  OR2_X1 U151bar ( .A1(abar[12]), .A2(bbar[3]), .ZN(ybar[195]) );
  AND2_X1 U152 ( .A1(a[12]), .A2(b[2]), .ZN(y[194]) );
  OR2_X1 U152bar ( .A1(abar[12]), .A2(bbar[2]), .ZN(ybar[194]) );
  AND2_X1 U153 ( .A1(a[12]), .A2(b[1]), .ZN(y[193]) );
  OR2_X1 U153bar ( .A1(abar[12]), .A2(bbar[1]), .ZN(ybar[193]) );
  AND2_X1 U154 ( .A1(a[12]), .A2(b[0]), .ZN(y[192]) );
  OR2_X1 U154bar ( .A1(abar[12]), .A2(bbar[0]), .ZN(ybar[192]) );
  AND2_X1 U155 ( .A1(a[11]), .A2(b[15]), .ZN(y[191]) );
  OR2_X1 U155bar ( .A1(abar[11]), .A2(bbar[15]), .ZN(ybar[191]) );
  AND2_X1 U156 ( .A1(a[11]), .A2(b[14]), .ZN(y[190]) );
  OR2_X1 U156bar ( .A1(abar[11]), .A2(bbar[14]), .ZN(ybar[190]) );
  AND2_X1 U157 ( .A1(a[1]), .A2(b[2]), .ZN(y[18]) );
  OR2_X1 U157bar ( .A1(abar[1]), .A2(bbar[2]), .ZN(ybar[18]) );
  AND2_X1 U158 ( .A1(a[11]), .A2(b[13]), .ZN(y[189]) );
  OR2_X1 U158bar ( .A1(abar[11]), .A2(bbar[13]), .ZN(ybar[189]) );
  AND2_X1 U159 ( .A1(a[11]), .A2(b[12]), .ZN(y[188]) );
  OR2_X1 U159bar ( .A1(abar[11]), .A2(bbar[12]), .ZN(ybar[188]) );
  AND2_X1 U160 ( .A1(a[11]), .A2(b[11]), .ZN(y[187]) );
  OR2_X1 U160bar ( .A1(abar[11]), .A2(bbar[11]), .ZN(ybar[187]) );
  AND2_X1 U161 ( .A1(a[11]), .A2(b[10]), .ZN(y[186]) );
  OR2_X1 U161bar ( .A1(abar[11]), .A2(bbar[10]), .ZN(ybar[186]) );
  AND2_X1 U162 ( .A1(a[11]), .A2(b[9]), .ZN(y[185]) );
  OR2_X1 U162bar ( .A1(abar[11]), .A2(bbar[9]), .ZN(ybar[185]) );
  AND2_X1 U163 ( .A1(a[11]), .A2(b[8]), .ZN(y[184]) );
  OR2_X1 U163bar ( .A1(abar[11]), .A2(bbar[8]), .ZN(ybar[184]) );
  AND2_X1 U164 ( .A1(a[11]), .A2(b[7]), .ZN(y[183]) );
  OR2_X1 U164bar ( .A1(abar[11]), .A2(bbar[7]), .ZN(ybar[183]) );
  AND2_X1 U165 ( .A1(a[11]), .A2(b[6]), .ZN(y[182]) );
  OR2_X1 U165bar ( .A1(abar[11]), .A2(bbar[6]), .ZN(ybar[182]) );
  AND2_X1 U166 ( .A1(a[11]), .A2(b[5]), .ZN(y[181]) );
  OR2_X1 U166bar ( .A1(abar[11]), .A2(bbar[5]), .ZN(ybar[181]) );
  AND2_X1 U167 ( .A1(a[11]), .A2(b[4]), .ZN(y[180]) );
  OR2_X1 U167bar ( .A1(abar[11]), .A2(bbar[4]), .ZN(ybar[180]) );
  AND2_X1 U168 ( .A1(a[1]), .A2(b[1]), .ZN(y[17]) );
  OR2_X1 U168bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[17]) );
  AND2_X1 U169 ( .A1(a[11]), .A2(b[3]), .ZN(y[179]) );
  OR2_X1 U169bar ( .A1(abar[11]), .A2(bbar[3]), .ZN(ybar[179]) );
  AND2_X1 U170 ( .A1(a[11]), .A2(b[2]), .ZN(y[178]) );
  OR2_X1 U170bar ( .A1(abar[11]), .A2(bbar[2]), .ZN(ybar[178]) );
  AND2_X1 U171 ( .A1(a[11]), .A2(b[1]), .ZN(y[177]) );
  OR2_X1 U171bar ( .A1(abar[11]), .A2(bbar[1]), .ZN(ybar[177]) );
  AND2_X1 U172 ( .A1(a[11]), .A2(b[0]), .ZN(y[176]) );
  OR2_X1 U172bar ( .A1(abar[11]), .A2(bbar[0]), .ZN(ybar[176]) );
  AND2_X1 U173 ( .A1(a[10]), .A2(b[15]), .ZN(y[175]) );
  OR2_X1 U173bar ( .A1(abar[10]), .A2(bbar[15]), .ZN(ybar[175]) );
  AND2_X1 U174 ( .A1(a[10]), .A2(b[14]), .ZN(y[174]) );
  OR2_X1 U174bar ( .A1(abar[10]), .A2(bbar[14]), .ZN(ybar[174]) );
  AND2_X1 U175 ( .A1(a[10]), .A2(b[13]), .ZN(y[173]) );
  OR2_X1 U175bar ( .A1(abar[10]), .A2(bbar[13]), .ZN(ybar[173]) );
  AND2_X1 U176 ( .A1(a[10]), .A2(b[12]), .ZN(y[172]) );
  OR2_X1 U176bar ( .A1(abar[10]), .A2(bbar[12]), .ZN(ybar[172]) );
  AND2_X1 U177 ( .A1(a[10]), .A2(b[11]), .ZN(y[171]) );
  OR2_X1 U177bar ( .A1(abar[10]), .A2(bbar[11]), .ZN(ybar[171]) );
  AND2_X1 U178 ( .A1(a[10]), .A2(b[10]), .ZN(y[170]) );
  OR2_X1 U178bar ( .A1(abar[10]), .A2(bbar[10]), .ZN(ybar[170]) );
  AND2_X1 U179 ( .A1(a[1]), .A2(b[0]), .ZN(y[16]) );
  OR2_X1 U179bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[16]) );
  AND2_X1 U180 ( .A1(a[10]), .A2(b[9]), .ZN(y[169]) );
  OR2_X1 U180bar ( .A1(abar[10]), .A2(bbar[9]), .ZN(ybar[169]) );
  AND2_X1 U181 ( .A1(a[10]), .A2(b[8]), .ZN(y[168]) );
  OR2_X1 U181bar ( .A1(abar[10]), .A2(bbar[8]), .ZN(ybar[168]) );
  AND2_X1 U182 ( .A1(a[10]), .A2(b[7]), .ZN(y[167]) );
  OR2_X1 U182bar ( .A1(abar[10]), .A2(bbar[7]), .ZN(ybar[167]) );
  AND2_X1 U183 ( .A1(a[10]), .A2(b[6]), .ZN(y[166]) );
  OR2_X1 U183bar ( .A1(abar[10]), .A2(bbar[6]), .ZN(ybar[166]) );
  AND2_X1 U184 ( .A1(a[10]), .A2(b[5]), .ZN(y[165]) );
  OR2_X1 U184bar ( .A1(abar[10]), .A2(bbar[5]), .ZN(ybar[165]) );
  AND2_X1 U185 ( .A1(a[10]), .A2(b[4]), .ZN(y[164]) );
  OR2_X1 U185bar ( .A1(abar[10]), .A2(bbar[4]), .ZN(ybar[164]) );
  AND2_X1 U186 ( .A1(a[10]), .A2(b[3]), .ZN(y[163]) );
  OR2_X1 U186bar ( .A1(abar[10]), .A2(bbar[3]), .ZN(ybar[163]) );
  AND2_X1 U187 ( .A1(a[10]), .A2(b[2]), .ZN(y[162]) );
  OR2_X1 U187bar ( .A1(abar[10]), .A2(bbar[2]), .ZN(ybar[162]) );
  AND2_X1 U188 ( .A1(a[10]), .A2(b[1]), .ZN(y[161]) );
  OR2_X1 U188bar ( .A1(abar[10]), .A2(bbar[1]), .ZN(ybar[161]) );
  AND2_X1 U189 ( .A1(a[10]), .A2(b[0]), .ZN(y[160]) );
  OR2_X1 U189bar ( .A1(abar[10]), .A2(bbar[0]), .ZN(ybar[160]) );
  AND2_X1 U190 ( .A1(b[15]), .A2(a[0]), .ZN(y[15]) );
  OR2_X1 U190bar ( .A1(bbar[15]), .A2(abar[0]), .ZN(ybar[15]) );
  AND2_X1 U191 ( .A1(a[9]), .A2(b[15]), .ZN(y[159]) );
  OR2_X1 U191bar ( .A1(abar[9]), .A2(bbar[15]), .ZN(ybar[159]) );
  AND2_X1 U192 ( .A1(a[9]), .A2(b[14]), .ZN(y[158]) );
  OR2_X1 U192bar ( .A1(abar[9]), .A2(bbar[14]), .ZN(ybar[158]) );
  AND2_X1 U193 ( .A1(a[9]), .A2(b[13]), .ZN(y[157]) );
  OR2_X1 U193bar ( .A1(abar[9]), .A2(bbar[13]), .ZN(ybar[157]) );
  AND2_X1 U194 ( .A1(a[9]), .A2(b[12]), .ZN(y[156]) );
  OR2_X1 U194bar ( .A1(abar[9]), .A2(bbar[12]), .ZN(ybar[156]) );
  AND2_X1 U195 ( .A1(a[9]), .A2(b[11]), .ZN(y[155]) );
  OR2_X1 U195bar ( .A1(abar[9]), .A2(bbar[11]), .ZN(ybar[155]) );
  AND2_X1 U196 ( .A1(a[9]), .A2(b[10]), .ZN(y[154]) );
  OR2_X1 U196bar ( .A1(abar[9]), .A2(bbar[10]), .ZN(ybar[154]) );
  AND2_X1 U197 ( .A1(a[9]), .A2(b[9]), .ZN(y[153]) );
  OR2_X1 U197bar ( .A1(abar[9]), .A2(bbar[9]), .ZN(ybar[153]) );
  AND2_X1 U198 ( .A1(a[9]), .A2(b[8]), .ZN(y[152]) );
  OR2_X1 U198bar ( .A1(abar[9]), .A2(bbar[8]), .ZN(ybar[152]) );
  AND2_X1 U199 ( .A1(a[9]), .A2(b[7]), .ZN(y[151]) );
  OR2_X1 U199bar ( .A1(abar[9]), .A2(bbar[7]), .ZN(ybar[151]) );
  AND2_X1 U200 ( .A1(a[9]), .A2(b[6]), .ZN(y[150]) );
  OR2_X1 U200bar ( .A1(abar[9]), .A2(bbar[6]), .ZN(ybar[150]) );
  AND2_X1 U201 ( .A1(b[14]), .A2(a[0]), .ZN(y[14]) );
  OR2_X1 U201bar ( .A1(bbar[14]), .A2(abar[0]), .ZN(ybar[14]) );
  AND2_X1 U202 ( .A1(a[9]), .A2(b[5]), .ZN(y[149]) );
  OR2_X1 U202bar ( .A1(abar[9]), .A2(bbar[5]), .ZN(ybar[149]) );
  AND2_X1 U203 ( .A1(a[9]), .A2(b[4]), .ZN(y[148]) );
  OR2_X1 U203bar ( .A1(abar[9]), .A2(bbar[4]), .ZN(ybar[148]) );
  AND2_X1 U204 ( .A1(a[9]), .A2(b[3]), .ZN(y[147]) );
  OR2_X1 U204bar ( .A1(abar[9]), .A2(bbar[3]), .ZN(ybar[147]) );
  AND2_X1 U205 ( .A1(a[9]), .A2(b[2]), .ZN(y[146]) );
  OR2_X1 U205bar ( .A1(abar[9]), .A2(bbar[2]), .ZN(ybar[146]) );
  AND2_X1 U206 ( .A1(a[9]), .A2(b[1]), .ZN(y[145]) );
  OR2_X1 U206bar ( .A1(abar[9]), .A2(bbar[1]), .ZN(ybar[145]) );
  AND2_X1 U207 ( .A1(a[9]), .A2(b[0]), .ZN(y[144]) );
  OR2_X1 U207bar ( .A1(abar[9]), .A2(bbar[0]), .ZN(ybar[144]) );
  AND2_X1 U208 ( .A1(a[8]), .A2(b[15]), .ZN(y[143]) );
  OR2_X1 U208bar ( .A1(abar[8]), .A2(bbar[15]), .ZN(ybar[143]) );
  AND2_X1 U209 ( .A1(a[8]), .A2(b[14]), .ZN(y[142]) );
  OR2_X1 U209bar ( .A1(abar[8]), .A2(bbar[14]), .ZN(ybar[142]) );
  AND2_X1 U210 ( .A1(a[8]), .A2(b[13]), .ZN(y[141]) );
  OR2_X1 U210bar ( .A1(abar[8]), .A2(bbar[13]), .ZN(ybar[141]) );
  AND2_X1 U211 ( .A1(a[8]), .A2(b[12]), .ZN(y[140]) );
  OR2_X1 U211bar ( .A1(abar[8]), .A2(bbar[12]), .ZN(ybar[140]) );
  AND2_X1 U212 ( .A1(b[13]), .A2(a[0]), .ZN(y[13]) );
  OR2_X1 U212bar ( .A1(bbar[13]), .A2(abar[0]), .ZN(ybar[13]) );
  AND2_X1 U213 ( .A1(a[8]), .A2(b[11]), .ZN(y[139]) );
  OR2_X1 U213bar ( .A1(abar[8]), .A2(bbar[11]), .ZN(ybar[139]) );
  AND2_X1 U214 ( .A1(a[8]), .A2(b[10]), .ZN(y[138]) );
  OR2_X1 U214bar ( .A1(abar[8]), .A2(bbar[10]), .ZN(ybar[138]) );
  AND2_X1 U215 ( .A1(a[8]), .A2(b[9]), .ZN(y[137]) );
  OR2_X1 U215bar ( .A1(abar[8]), .A2(bbar[9]), .ZN(ybar[137]) );
  AND2_X1 U216 ( .A1(a[8]), .A2(b[8]), .ZN(y[136]) );
  OR2_X1 U216bar ( .A1(abar[8]), .A2(bbar[8]), .ZN(ybar[136]) );
  AND2_X1 U217 ( .A1(a[8]), .A2(b[7]), .ZN(y[135]) );
  OR2_X1 U217bar ( .A1(abar[8]), .A2(bbar[7]), .ZN(ybar[135]) );
  AND2_X1 U218 ( .A1(a[8]), .A2(b[6]), .ZN(y[134]) );
  OR2_X1 U218bar ( .A1(abar[8]), .A2(bbar[6]), .ZN(ybar[134]) );
  AND2_X1 U219 ( .A1(a[8]), .A2(b[5]), .ZN(y[133]) );
  OR2_X1 U219bar ( .A1(abar[8]), .A2(bbar[5]), .ZN(ybar[133]) );
  AND2_X1 U220 ( .A1(a[8]), .A2(b[4]), .ZN(y[132]) );
  OR2_X1 U220bar ( .A1(abar[8]), .A2(bbar[4]), .ZN(ybar[132]) );
  AND2_X1 U221 ( .A1(a[8]), .A2(b[3]), .ZN(y[131]) );
  OR2_X1 U221bar ( .A1(abar[8]), .A2(bbar[3]), .ZN(ybar[131]) );
  AND2_X1 U222 ( .A1(a[8]), .A2(b[2]), .ZN(y[130]) );
  OR2_X1 U222bar ( .A1(abar[8]), .A2(bbar[2]), .ZN(ybar[130]) );
  AND2_X1 U223 ( .A1(b[12]), .A2(a[0]), .ZN(y[12]) );
  OR2_X1 U223bar ( .A1(bbar[12]), .A2(abar[0]), .ZN(ybar[12]) );
  AND2_X1 U224 ( .A1(a[8]), .A2(b[1]), .ZN(y[129]) );
  OR2_X1 U224bar ( .A1(abar[8]), .A2(bbar[1]), .ZN(ybar[129]) );
  AND2_X1 U225 ( .A1(a[8]), .A2(b[0]), .ZN(y[128]) );
  OR2_X1 U225bar ( .A1(abar[8]), .A2(bbar[0]), .ZN(ybar[128]) );
  AND2_X1 U226 ( .A1(a[7]), .A2(b[15]), .ZN(y[127]) );
  OR2_X1 U226bar ( .A1(abar[7]), .A2(bbar[15]), .ZN(ybar[127]) );
  AND2_X1 U227 ( .A1(a[7]), .A2(b[14]), .ZN(y[126]) );
  OR2_X1 U227bar ( .A1(abar[7]), .A2(bbar[14]), .ZN(ybar[126]) );
  AND2_X1 U228 ( .A1(a[7]), .A2(b[13]), .ZN(y[125]) );
  OR2_X1 U228bar ( .A1(abar[7]), .A2(bbar[13]), .ZN(ybar[125]) );
  AND2_X1 U229 ( .A1(a[7]), .A2(b[12]), .ZN(y[124]) );
  OR2_X1 U229bar ( .A1(abar[7]), .A2(bbar[12]), .ZN(ybar[124]) );
  AND2_X1 U230 ( .A1(a[7]), .A2(b[11]), .ZN(y[123]) );
  OR2_X1 U230bar ( .A1(abar[7]), .A2(bbar[11]), .ZN(ybar[123]) );
  AND2_X1 U231 ( .A1(a[7]), .A2(b[10]), .ZN(y[122]) );
  OR2_X1 U231bar ( .A1(abar[7]), .A2(bbar[10]), .ZN(ybar[122]) );
  AND2_X1 U232 ( .A1(a[7]), .A2(b[9]), .ZN(y[121]) );
  OR2_X1 U232bar ( .A1(abar[7]), .A2(bbar[9]), .ZN(ybar[121]) );
  AND2_X1 U233 ( .A1(a[7]), .A2(b[8]), .ZN(y[120]) );
  OR2_X1 U233bar ( .A1(abar[7]), .A2(bbar[8]), .ZN(ybar[120]) );
  AND2_X1 U234 ( .A1(b[11]), .A2(a[0]), .ZN(y[11]) );
  OR2_X1 U234bar ( .A1(bbar[11]), .A2(abar[0]), .ZN(ybar[11]) );
  AND2_X1 U235 ( .A1(a[7]), .A2(b[7]), .ZN(y[119]) );
  OR2_X1 U235bar ( .A1(abar[7]), .A2(bbar[7]), .ZN(ybar[119]) );
  AND2_X1 U236 ( .A1(a[7]), .A2(b[6]), .ZN(y[118]) );
  OR2_X1 U236bar ( .A1(abar[7]), .A2(bbar[6]), .ZN(ybar[118]) );
  AND2_X1 U237 ( .A1(a[7]), .A2(b[5]), .ZN(y[117]) );
  OR2_X1 U237bar ( .A1(abar[7]), .A2(bbar[5]), .ZN(ybar[117]) );
  AND2_X1 U238 ( .A1(a[7]), .A2(b[4]), .ZN(y[116]) );
  OR2_X1 U238bar ( .A1(abar[7]), .A2(bbar[4]), .ZN(ybar[116]) );
  AND2_X1 U239 ( .A1(a[7]), .A2(b[3]), .ZN(y[115]) );
  OR2_X1 U239bar ( .A1(abar[7]), .A2(bbar[3]), .ZN(ybar[115]) );
  AND2_X1 U240 ( .A1(a[7]), .A2(b[2]), .ZN(y[114]) );
  OR2_X1 U240bar ( .A1(abar[7]), .A2(bbar[2]), .ZN(ybar[114]) );
  AND2_X1 U241 ( .A1(a[7]), .A2(b[1]), .ZN(y[113]) );
  OR2_X1 U241bar ( .A1(abar[7]), .A2(bbar[1]), .ZN(ybar[113]) );
  AND2_X1 U242 ( .A1(a[7]), .A2(b[0]), .ZN(y[112]) );
  OR2_X1 U242bar ( .A1(abar[7]), .A2(bbar[0]), .ZN(ybar[112]) );
  AND2_X1 U243 ( .A1(b[15]), .A2(a[6]), .ZN(y[111]) );
  OR2_X1 U243bar ( .A1(bbar[15]), .A2(abar[6]), .ZN(ybar[111]) );
  AND2_X1 U244 ( .A1(b[14]), .A2(a[6]), .ZN(y[110]) );
  OR2_X1 U244bar ( .A1(bbar[14]), .A2(abar[6]), .ZN(ybar[110]) );
  AND2_X1 U245 ( .A1(b[10]), .A2(a[0]), .ZN(y[10]) );
  OR2_X1 U245bar ( .A1(bbar[10]), .A2(abar[0]), .ZN(ybar[10]) );
  AND2_X1 U246 ( .A1(b[13]), .A2(a[6]), .ZN(y[109]) );
  OR2_X1 U246bar ( .A1(bbar[13]), .A2(abar[6]), .ZN(ybar[109]) );
  AND2_X1 U247 ( .A1(b[12]), .A2(a[6]), .ZN(y[108]) );
  OR2_X1 U247bar ( .A1(bbar[12]), .A2(abar[6]), .ZN(ybar[108]) );
  AND2_X1 U248 ( .A1(b[11]), .A2(a[6]), .ZN(y[107]) );
  OR2_X1 U248bar ( .A1(bbar[11]), .A2(abar[6]), .ZN(ybar[107]) );
  AND2_X1 U249 ( .A1(b[10]), .A2(a[6]), .ZN(y[106]) );
  OR2_X1 U249bar ( .A1(bbar[10]), .A2(abar[6]), .ZN(ybar[106]) );
  AND2_X1 U250 ( .A1(a[6]), .A2(b[9]), .ZN(y[105]) );
  OR2_X1 U250bar ( .A1(abar[6]), .A2(bbar[9]), .ZN(ybar[105]) );
  AND2_X1 U251 ( .A1(b[8]), .A2(a[6]), .ZN(y[104]) );
  OR2_X1 U251bar ( .A1(bbar[8]), .A2(abar[6]), .ZN(ybar[104]) );
  AND2_X1 U252 ( .A1(b[7]), .A2(a[6]), .ZN(y[103]) );
  OR2_X1 U252bar ( .A1(bbar[7]), .A2(abar[6]), .ZN(ybar[103]) );
  AND2_X1 U253 ( .A1(b[6]), .A2(a[6]), .ZN(y[102]) );
  OR2_X1 U253bar ( .A1(bbar[6]), .A2(abar[6]), .ZN(ybar[102]) );
  AND2_X1 U254 ( .A1(b[5]), .A2(a[6]), .ZN(y[101]) );
  OR2_X1 U254bar ( .A1(bbar[5]), .A2(abar[6]), .ZN(ybar[101]) );
  AND2_X1 U255 ( .A1(b[4]), .A2(a[6]), .ZN(y[100]) );
  OR2_X1 U255bar ( .A1(bbar[4]), .A2(abar[6]), .ZN(ybar[100]) );
  AND2_X1 U256 ( .A1(b[0]), .A2(a[0]), .ZN(y[0]) );
  OR2_X1 U256bar ( .A1(bbar[0]), .A2(abar[0]), .ZN(ybar[0]) );
endmodule

module CD2_77 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD2_78 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD2_79 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD4_39 ( a, abar, b, bbar, y, ybar );

  input wire [3:0] a;
  input wire [3:0] b;
  input wire [3:0] abar;
  input wire [3:0] bbar;
//input_done

  output wire [15:0] y;
  output wire [15:0] ybar;
//output_done

//wire_done

  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]) );
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]) );
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]) );
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]) );
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]) );
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]) );
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]) );
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]) );
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]) );
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]) );
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]) );
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]) );
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]) );
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]) );
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]) );
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]) );
endmodule

module decode_0 ( in, inbar, out, outbar );

  input wire [7:0] in;
  input wire [7:0] inbar;
//input_done

  output wire [255:0] out;
  output wire [255:0] outbar;
//output_done

  wire [15:0] level1;
  wire [31:0] level2;
  wire [15:0] level1bar;
  wire [31:0] level2bar;
//wire_done

  CD2_0 cd_l1_1 ( .a(in[1]), .abar(inbar[1]), .b(in[0]), .bbar(inbar[0]), .y(level1[3:0]), .ybar(level1bar[3:0]) );
  CD2_79 cd_l1_2 ( .a(in[3]), .abar(inbar[3]), .b(in[2]), .bbar(inbar[2]), .y(level1[7:4]), .ybar(level1bar[7:4]) );
  CD2_78 cd_l1_3 ( .a(in[5]), .abar(inbar[5]), .b(in[4]), .bbar(inbar[4]), .y(level1[11:8]), .ybar(level1bar[11:8]) );
  CD2_77 cd_l1_4 ( .a(in[7]), .abar(inbar[7]), .b(in[6]), .bbar(inbar[6]), .y(level1[15:12]), .ybar(level1bar[15:12]) );

  CD4_0 cd_l2_1 ( .a(level1[7:4]), .abar(level1bar[7:4]), .b(level1[3:0]), .bbar(level1bar[3:0]), 
        .y(level2[15:0]), .ybar(level2bar[15:0]) );
  CD4_39 cd_l2_2 ( .a(level1[15:12]), .abar(level1bar[15:12]), .b(level1[11:8]), .bbar(level1bar[11:8]), 
        .y(level2[31:16]), .ybar(level2bar[31:16]) );
  CD16_0 cd_l3 ( .a(level2[31:16]), .abar(level2bar[31:16]), .b(level2[15:0]), .bbar(level2bar[15:0]), 
        .y(out), .ybar(outbar) );
endmodule

module encode_0 ( in, inbar, out, outbar );

  input wire [255:0] in;
  input wire [255:0] inbar;
//input_done

  output wire [7:0] out;
  output wire [7:0] outbar;
//output_done

  wire in_81;
  wire in_80;
  wire in_79;
  wire in_78;
  wire in_77;
  wire in_76;
  wire in_75;
  wire in_74;
  wire in_73;
  wire in_72;
  wire in_71;
  wire in_70;
  wire in_69;
  wire in_68;
  wire in_67;
  wire in_66;
  wire in_65;
  wire in_64;
  wire in_63;
  wire in_62;
  wire in_61;
  wire in_60;
  wire in_59;
  wire in_58;
  wire in_57;
  wire in_56;
  wire in_55;
  wire in_54;
  wire in_53;
  wire in_52;
  wire in_51;
  wire in_50;
  wire in_49;
  wire in_48;
  wire in_47;
  wire in_46;
  wire in_45;
  wire in_44;
  wire in_43;
  wire in_42;
  wire in_41;
  wire in_40;
  wire in_39;
  wire in_38;
  wire in_37;
  wire in_36;
  wire in_35;
  wire in_34;
  wire in_33;
  wire in_32;
  wire in_31;
  wire in_30;
  wire in_29;
  wire in_28;
  wire in_27;
  wire in_26;
  wire in_25;
  wire in_24;
  wire in_23;
  wire in_22;
  wire in_21;
  wire in_20;
  wire in_19;
  wire in_18;
  wire in_17;
  wire in_16;
  wire in_15;
  wire in_14;
  wire in_13;
  wire in_12;
  wire in_11;
  wire in_10;
  wire in_9;
  wire in_8;
  wire in_7;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_3;
  wire in_2;
  wire in_1;
  wire in_0;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire in_81bar;
  wire in_80bar;
  wire in_79bar;
  wire in_78bar;
  wire in_77bar;
  wire in_76bar;
  wire in_75bar;
  wire in_74bar;
  wire in_73bar;
  wire in_72bar;
  wire in_71bar;
  wire in_70bar;
  wire in_69bar;
  wire in_68bar;
  wire in_67bar;
  wire in_66bar;
  wire in_65bar;
  wire in_64bar;
  wire in_63bar;
  wire in_62bar;
  wire in_61bar;
  wire in_60bar;
  wire in_59bar;
  wire in_58bar;
  wire in_57bar;
  wire in_56bar;
  wire in_55bar;
  wire in_54bar;
  wire in_53bar;
  wire in_52bar;
  wire in_51bar;
  wire in_50bar;
  wire in_49bar;
  wire in_48bar;
  wire in_47bar;
  wire in_46bar;
  wire in_45bar;
  wire in_44bar;
  wire in_43bar;
  wire in_42bar;
  wire in_41bar;
  wire in_40bar;
  wire in_39bar;
  wire in_38bar;
  wire in_37bar;
  wire in_36bar;
  wire in_35bar;
  wire in_34bar;
  wire in_33bar;
  wire in_32bar;
  wire in_31bar;
  wire in_30bar;
  wire in_29bar;
  wire in_28bar;
  wire in_27bar;
  wire in_26bar;
  wire in_25bar;
  wire in_24bar;
  wire in_23bar;
  wire in_22bar;
  wire in_21bar;
  wire in_20bar;
  wire in_19bar;
  wire in_18bar;
  wire in_17bar;
  wire in_16bar;
  wire in_15bar;
  wire in_14bar;
  wire in_13bar;
  wire in_12bar;
  wire in_11bar;
  wire in_10bar;
  wire in_9bar;
  wire in_8bar;
  wire in_7bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_3bar;
  wire in_2bar;
  wire in_1bar;
  wire in_0bar;
  wire n487bar;
  wire n488bar;
  wire n489bar;
  wire n490bar;
  wire n491bar;
  wire n492bar;
  wire n493bar;
  wire n494bar;
  wire n495bar;
  wire n496bar;
  wire n497bar;
  wire n498bar;
  wire n499bar;
  wire n500bar;
  wire n501bar;
  wire n502bar;
  wire n503bar;
  wire n504bar;
  wire n505bar;
  wire n506bar;
  wire n507bar;
  wire n508bar;
  wire n509bar;
  wire n510bar;
  wire n511bar;
  wire n512bar;
  wire n513bar;
  wire n514bar;
  wire n515bar;
  wire n516bar;
  wire n517bar;
  wire n518bar;
  wire n519bar;
  wire n520bar;
  wire n521bar;
  wire n522bar;
  wire n523bar;
  wire n524bar;
  wire n525bar;
  wire n526bar;
  wire n527bar;
  wire n528bar;
  wire n529bar;
  wire n530bar;
  wire n531bar;
  wire n532bar;
  wire n533bar;
  wire n534bar;
  wire n535bar;
  wire n536bar;
  wire n537bar;
  wire n538bar;
  wire n539bar;
  wire n540bar;
  wire n541bar;
  wire n542bar;
  wire n543bar;
  wire n544bar;
  wire n545bar;
  wire n546bar;
  wire n547bar;
  wire n548bar;
  wire n549bar;
  wire n550bar;
  wire n551bar;
  wire n552bar;
  wire n553bar;
  wire n554bar;
  wire n555bar;
  wire n556bar;
  wire n557bar;
  wire n558bar;
  wire n559bar;
  wire n560bar;
  wire n561bar;
  wire n562bar;
  wire n563bar;
  wire n564bar;
  wire n565bar;
  wire n566bar;
  wire n567bar;
  wire n568bar;
  wire n569bar;
  wire n570bar;
  wire n571bar;
  wire n572bar;
  wire n573bar;
  wire n574bar;
  wire n575bar;
  wire n576bar;
  wire n577bar;
  wire n578bar;
  wire n579bar;
  wire n580bar;
  wire n581bar;
  wire n582bar;
  wire n583bar;
  wire n584bar;
  wire n585bar;
  wire n586bar;
  wire n587bar;
  wire n588bar;
  wire n589bar;
  wire n590bar;
  wire n591bar;
  wire n592bar;
  wire n593bar;
  wire n594bar;
  wire n595bar;
  wire n596bar;
  wire n597bar;
  wire n598bar;
  wire n599bar;
  wire n600bar;
  wire n601bar;
  wire n602bar;
  wire n603bar;
  wire n604bar;
  wire n605bar;
  wire n606bar;
  wire n607bar;
  wire n608bar;
  wire n609bar;
  wire n610bar;
  wire n611bar;
  wire n612bar;
  wire n613bar;
  wire n614bar;
  wire n615bar;
  wire n616bar;
  wire n617bar;
  wire n618bar;
  wire n619bar;
  wire n620bar;
  wire n621bar;
  wire n622bar;
  wire n623bar;
  wire n624bar;
  wire n625bar;
  wire n626bar;
  wire n627bar;
  wire n628bar;
  wire n629bar;
  wire n630bar;
  wire n631bar;
  wire n632bar;
  wire n633bar;
  wire n634bar;
  wire n635bar;
  wire n636bar;
  wire n637bar;
  wire n638bar;
  wire n639bar;
  wire n640bar;
  wire n641bar;
  wire n642bar;
  wire n643bar;
  wire n644bar;
  wire n645bar;
  wire n646bar;
  wire n647bar;
  wire n648bar;
  wire n649bar;
  wire n650bar;
  wire n651bar;
  wire n652bar;
  wire n653bar;
  wire n654bar;
  wire n655bar;
  wire n656bar;
  wire n657bar;
  wire n658bar;
  wire n659bar;
  wire n660bar;
  wire n661bar;
  wire n662bar;
  wire n663bar;
  wire n664bar;
  wire n665bar;
  wire n666bar;
  wire n667bar;
  wire n668bar;
  wire n669bar;
  wire n670bar;
  wire n671bar;
  wire n672bar;
  wire n673bar;
  wire n674bar;
  wire n675bar;
  wire n676bar;
  wire n677bar;
  wire n678bar;
  wire n679bar;
  wire n680bar;
  wire n681bar;
  wire n682bar;
  wire n683bar;
  wire n684bar;
  wire n685bar;
  wire n686bar;
  wire n687bar;
  wire n688bar;
  wire n689bar;
  wire n690bar;
  wire n691bar;
  wire n692bar;
  wire n693bar;
  wire n694bar;
  wire n695bar;
  wire n696bar;
  wire n697bar;
  wire n698bar;
  wire n699bar;
  wire n700bar;
  wire n701bar;
  wire n702bar;
  wire n703bar;
  wire n704bar;
  wire n705bar;
  wire n706bar;
  wire n707bar;
  wire n708bar;
  wire n709bar;
  wire n710bar;
  wire n711bar;
  wire n712bar;
  wire n713bar;
  wire n714bar;
  wire n715bar;
  wire n716bar;
  wire n717bar;
  wire n718bar;
  wire n719bar;
  wire n720bar;
  wire n721bar;
  wire n722bar;
  wire n723bar;
  wire n724bar;
  wire n725bar;
  wire n726bar;
  wire n727bar;
  wire n728bar;
  wire n729bar;
  wire n730bar;
  wire n731bar;
  wire n732bar;
  wire n733bar;
  wire n734bar;
  wire n735bar;
  wire n736bar;
  wire n737bar;
  wire n738bar;
  wire n739bar;
  wire n740bar;
  wire n741bar;
  wire n742bar;
  wire n743bar;
  wire n744bar;
  wire n745bar;
  wire n746bar;
  wire n747bar;
  wire n748bar;
  wire n749bar;
  wire n750bar;
  wire n751bar;
  wire n752bar;
  wire n753bar;
  wire n754bar;
  wire n755bar;
  wire n756bar;
  wire n757bar;
  wire n758bar;
  wire n759bar;
  wire n760bar;
  wire n761bar;
  wire n762bar;
  wire n763bar;
  wire n764bar;
  wire n765bar;
  wire n766bar;
  wire n767bar;
  wire n768bar;
  wire n769bar;
  wire n770bar;
  wire n771bar;
  wire n772bar;
  wire n773bar;
  wire n774bar;
  wire n775bar;
  wire n776bar;
  wire n777bar;
  wire n778bar;
  wire n779bar;
  wire n780bar;
  wire n781bar;
  wire n782bar;
  wire n783bar;
  wire n784bar;
  wire n785bar;
  wire n786bar;
  wire n787bar;
  wire n788bar;
  wire n789bar;
  wire n790bar;
  wire n791bar;
  wire n792bar;
  wire n793bar;
  wire n794bar;
  wire n795bar;
  wire n796bar;
  wire n797bar;
  wire n798bar;
  wire n799bar;
  wire n800bar;
  wire n801bar;
  wire n802bar;
  wire n803bar;
  wire n804bar;
  wire n805bar;
  wire n806bar;
  wire n807bar;
  wire n808bar;
  wire n809bar;
  wire n810bar;
  wire n811bar;
  wire n812bar;
  wire n813bar;
  wire n814bar;
  wire n815bar;
  wire n816bar;
  wire n817bar;
  wire n818bar;
  wire n819bar;
  wire n820bar;
  wire n821bar;
  wire n822bar;
  wire n823bar;
  wire n824bar;
  wire n825bar;
  wire n826bar;
  wire n827bar;
  wire n828bar;
  wire n829bar;
  wire n830bar;
  wire n831bar;
  wire n832bar;
  wire n833bar;
  wire n834bar;
  wire n835bar;
  wire n836bar;
  wire n837bar;
  wire n838bar;
  wire n839bar;
  wire n840bar;
  wire n841bar;
  wire n842bar;
  wire n843bar;
  wire n844bar;
  wire n845bar;
  wire n846bar;
  wire n847bar;
  wire n848bar;
  wire n849bar;
  wire n850bar;
  wire n851bar;
  wire n852bar;
  wire n853bar;
  wire n854bar;
  wire n855bar;
  wire n856bar;
  wire n857bar;
  wire n858bar;
  wire n859bar;
  wire n860bar;
  wire n861bar;
  wire n862bar;
  wire n863bar;
  wire n864bar;
  wire n865bar;
  wire n866bar;
  wire n867bar;
  wire n868bar;
  wire n869bar;
  wire n870bar;
  wire n871bar;
  wire n872bar;
  wire n873bar;
  wire n874bar;
  wire n875bar;
  wire n876bar;
  wire n877bar;
  wire n878bar;
  wire n879bar;
  wire n880bar;
  wire n881bar;
  wire n882bar;
  wire n883bar;
  wire n884bar;
  wire n885bar;
  wire n886bar;
  wire n887bar;
  wire n888bar;
  wire n889bar;
  wire n890bar;
  wire n891bar;
  wire n892bar;
  wire n893bar;
  wire n894bar;
  wire n895bar;
  wire n896bar;
  wire n897bar;
  wire n898bar;
  wire n899bar;
  wire n900bar;
  wire n901bar;
  wire n902bar;
  wire n903bar;
  wire n904bar;
  wire n905bar;
  wire n906bar;
  wire n907bar;
  wire n908bar;
  wire n909bar;
  wire n910bar;
  wire n911bar;
  wire n912bar;
  wire n913bar;
  wire n914bar;
  wire n915bar;
  wire n916bar;
  wire n917bar;
  wire n918bar;
  wire n919bar;
  wire n920bar;
  wire n921bar;
  wire n922bar;
  wire n923bar;
  wire n924bar;
  wire n925bar;
  wire n926bar;
  wire n927bar;
  wire n928bar;
  wire n929bar;
  wire n930bar;
  wire n931bar;
  wire n932bar;
  wire n933bar;
  wire n934bar;
  wire n935bar;
  wire n936bar;
  wire n937bar;
  wire n938bar;
  wire n939bar;
  wire n940bar;
  wire n941bar;
  wire n942bar;
  wire n943bar;
  wire n944bar;
  wire n945bar;
  wire n946bar;
  wire n947bar;
  wire n948bar;
  wire n949bar;
  wire n950bar;
  wire n951bar;
  wire n952bar;
  wire n953bar;
  wire n954bar;
  wire n955bar;
  wire n956bar;
  wire n957bar;
  wire n958bar;
  wire n959bar;
  wire n960bar;
  wire n961bar;
  wire n962bar;
  wire n963bar;
  wire n964bar;
  wire n965bar;
  wire n966bar;
  wire n967bar;
  wire n968bar;
  wire n969bar;
  wire n970bar;
  wire n971bar;
  wire n972bar;
//wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];
  assign in_81bar = inbar[81];
  assign in_80bar = inbar[80];
  assign in_79bar = inbar[79];
  assign in_78bar = inbar[78];
  assign in_77bar = inbar[77];
  assign in_76bar = inbar[76];
  assign in_75bar = inbar[75];
  assign in_74bar = inbar[74];
  assign in_73bar = inbar[73];
  assign in_72bar = inbar[72];
  assign in_71bar = inbar[71];
  assign in_70bar = inbar[70];
  assign in_69bar = inbar[69];
  assign in_68bar = inbar[68];
  assign in_67bar = inbar[67];
  assign in_66bar = inbar[66];
  assign in_65bar = inbar[65];
  assign in_64bar = inbar[64];
  assign in_63bar = inbar[63];
  assign in_62bar = inbar[62];
  assign in_61bar = inbar[61];
  assign in_60bar = inbar[60];
  assign in_59bar = inbar[59];
  assign in_58bar = inbar[58];
  assign in_57bar = inbar[57];
  assign in_56bar = inbar[56];
  assign in_55bar = inbar[55];
  assign in_54bar = inbar[54];
  assign in_53bar = inbar[53];
  assign in_52bar = inbar[52];
  assign in_51bar = inbar[51];
  assign in_50bar = inbar[50];
  assign in_49bar = inbar[49];
  assign in_48bar = inbar[48];
  assign in_47bar = inbar[47];
  assign in_46bar = inbar[46];
  assign in_45bar = inbar[45];
  assign in_44bar = inbar[44];
  assign in_43bar = inbar[43];
  assign in_42bar = inbar[42];
  assign in_41bar = inbar[41];
  assign in_40bar = inbar[40];
  assign in_39bar = inbar[39];
  assign in_38bar = inbar[38];
  assign in_37bar = inbar[37];
  assign in_36bar = inbar[36];
  assign in_35bar = inbar[35];
  assign in_34bar = inbar[34];
  assign in_33bar = inbar[33];
  assign in_32bar = inbar[32];
  assign in_31bar = inbar[31];
  assign in_30bar = inbar[30];
  assign in_29bar = inbar[29];
  assign in_28bar = inbar[28];
  assign in_27bar = inbar[27];
  assign in_26bar = inbar[26];
  assign in_25bar = inbar[25];
  assign in_24bar = inbar[24];
  assign in_23bar = inbar[23];
  assign in_22bar = inbar[22];
  assign in_21bar = inbar[21];
  assign in_20bar = inbar[20];
  assign in_19bar = inbar[19];
  assign in_18bar = inbar[18];
  assign in_17bar = inbar[17];
  assign in_16bar = inbar[16];
  assign in_15bar = inbar[15];
  assign in_14bar = inbar[14];
  assign in_13bar = inbar[13];
  assign in_12bar = inbar[12];
  assign in_11bar = inbar[11];
  assign in_10bar = inbar[10];
  assign in_9bar = inbar[9];
  assign in_8bar = inbar[8];
  assign in_7bar = inbar[7];
  assign in_6bar = inbar[6];
  assign in_5bar = inbar[5];
  assign in_4bar = inbar[4];
  assign in_3bar = inbar[3];
  assign in_2bar = inbar[2];
  assign in_1bar = inbar[1];
  assign in_0bar = inbar[0];
//assign_done

  OR2_X1 U1 ( .A1(n972), .A2(n971), .ZN(out[7]) );
  AND2_X1 U1bar ( .A1(n972bar), .A2(n971bar), .ZN(outbar[7]) );
  OR2_X1 U2 ( .A1(n970), .A2(n969), .ZN(n971) );
  AND2_X1 U2bar ( .A1(n970bar), .A2(n969bar), .ZN(n971bar) );
  OR2_X1 U3 ( .A1(n968), .A2(n967), .ZN(n969) );
  AND2_X1 U3bar ( .A1(n968bar), .A2(n967bar), .ZN(n969bar) );
  OR2_X1 U4 ( .A1(n966), .A2(n965), .ZN(n967) );
  AND2_X1 U4bar ( .A1(n966bar), .A2(n965bar), .ZN(n967bar) );
  OR2_X1 U5 ( .A1(n964), .A2(n963), .ZN(n968) );
  AND2_X1 U5bar ( .A1(n964bar), .A2(n963bar), .ZN(n968bar) );
  OR2_X1 U6 ( .A1(in[116]), .A2(n962), .ZN(n963) );
  AND2_X1 U6bar ( .A1(inbar[116]), .A2(n962bar), .ZN(n963bar) );
  OR2_X1 U7 ( .A1(n961), .A2(n960), .ZN(n970) );
  AND2_X1 U7bar ( .A1(n961bar), .A2(n960bar), .ZN(n970bar) );
  OR2_X1 U8 ( .A1(in[150]), .A2(in[127]), .ZN(n960) );
  AND2_X1 U8bar ( .A1(inbar[150]), .A2(inbar[127]), .ZN(n960bar) );
  OR2_X1 U9 ( .A1(in[160]), .A2(n959), .ZN(n961) );
  AND2_X1 U9bar ( .A1(inbar[160]), .A2(n959bar), .ZN(n961bar) );
  OR2_X1 U10 ( .A1(in[252]), .A2(in[168]), .ZN(n959) );
  AND2_X1 U10bar ( .A1(inbar[252]), .A2(inbar[168]), .ZN(n959bar) );
  OR2_X1 U11 ( .A1(n958), .A2(n957), .ZN(n972) );
  AND2_X1 U11bar ( .A1(n958bar), .A2(n957bar), .ZN(n972bar) );
  OR2_X1 U12 ( .A1(n956), .A2(n955), .ZN(n957) );
  AND2_X1 U12bar ( .A1(n956bar), .A2(n955bar), .ZN(n957bar) );
  OR2_X1 U13 ( .A1(in_17), .A2(in[96]), .ZN(n955) );
  AND2_X1 U13bar ( .A1(in_17bar), .A2(inbar[96]), .ZN(n955bar) );
  OR2_X1 U14 ( .A1(in_23), .A2(n954), .ZN(n956) );
  AND2_X1 U14bar ( .A1(in_23bar), .A2(n954bar), .ZN(n956bar) );
  OR2_X1 U15 ( .A1(in_31), .A2(in_26), .ZN(n954) );
  AND2_X1 U15bar ( .A1(in_31bar), .A2(in_26bar), .ZN(n954bar) );
  OR2_X1 U16 ( .A1(n953), .A2(n952), .ZN(n958) );
  AND2_X1 U16bar ( .A1(n953bar), .A2(n952bar), .ZN(n958bar) );
  OR2_X1 U17 ( .A1(in_58), .A2(in_4), .ZN(n952) );
  AND2_X1 U17bar ( .A1(in_58bar), .A2(in_4bar), .ZN(n952bar) );
  OR2_X1 U18 ( .A1(in_59), .A2(n951), .ZN(n953) );
  AND2_X1 U18bar ( .A1(in_59bar), .A2(n951bar), .ZN(n953bar) );
  OR2_X1 U19 ( .A1(in_71), .A2(in_62), .ZN(n951) );
  AND2_X1 U19bar ( .A1(in_71bar), .A2(in_62bar), .ZN(n951bar) );
  OR2_X1 U20 ( .A1(n950), .A2(n949), .ZN(out[6]) );
  AND2_X1 U20bar ( .A1(n950bar), .A2(n949bar), .ZN(outbar[6]) );
  OR2_X1 U21 ( .A1(n948), .A2(n947), .ZN(n949) );
  AND2_X1 U21bar ( .A1(n948bar), .A2(n947bar), .ZN(n949bar) );
  OR2_X1 U22 ( .A1(n946), .A2(n945), .ZN(n947) );
  AND2_X1 U22bar ( .A1(n946bar), .A2(n945bar), .ZN(n947bar) );
  OR2_X1 U23 ( .A1(n944), .A2(n943), .ZN(n945) );
  AND2_X1 U23bar ( .A1(n944bar), .A2(n943bar), .ZN(n945bar) );
  OR2_X1 U24 ( .A1(n942), .A2(n941), .ZN(n946) );
  AND2_X1 U24bar ( .A1(n942bar), .A2(n941bar), .ZN(n946bar) );
  OR2_X1 U25 ( .A1(in[101]), .A2(n940), .ZN(n941) );
  AND2_X1 U25bar ( .A1(inbar[101]), .A2(n940bar), .ZN(n941bar) );
  OR2_X1 U26 ( .A1(n939), .A2(n938), .ZN(n948) );
  AND2_X1 U26bar ( .A1(n939bar), .A2(n938bar), .ZN(n948bar) );
  OR2_X1 U27 ( .A1(in[114]), .A2(in[104]), .ZN(n938) );
  AND2_X1 U27bar ( .A1(inbar[114]), .A2(inbar[104]), .ZN(n938bar) );
  OR2_X1 U28 ( .A1(in[128]), .A2(n937), .ZN(n939) );
  AND2_X1 U28bar ( .A1(inbar[128]), .A2(n937bar), .ZN(n939bar) );
  OR2_X1 U29 ( .A1(in[136]), .A2(in[134]), .ZN(n937) );
  AND2_X1 U29bar ( .A1(inbar[136]), .A2(inbar[134]), .ZN(n937bar) );
  OR2_X1 U30 ( .A1(n936), .A2(n935), .ZN(n950) );
  AND2_X1 U30bar ( .A1(n936bar), .A2(n935bar), .ZN(n950bar) );
  OR2_X1 U31 ( .A1(n934), .A2(n933), .ZN(n935) );
  AND2_X1 U31bar ( .A1(n934bar), .A2(n933bar), .ZN(n935bar) );
  OR2_X1 U32 ( .A1(in[177]), .A2(in[164]), .ZN(n933) );
  AND2_X1 U32bar ( .A1(inbar[177]), .A2(inbar[164]), .ZN(n933bar) );
  OR2_X1 U33 ( .A1(in[212]), .A2(n932), .ZN(n934) );
  AND2_X1 U33bar ( .A1(inbar[212]), .A2(n932bar), .ZN(n934bar) );
  OR2_X1 U34 ( .A1(in[248]), .A2(in[221]), .ZN(n932) );
  AND2_X1 U34bar ( .A1(inbar[248]), .A2(inbar[221]), .ZN(n932bar) );
  OR2_X1 U35 ( .A1(n931), .A2(n930), .ZN(n936) );
  AND2_X1 U35bar ( .A1(n931bar), .A2(n930bar), .ZN(n936bar) );
  OR2_X1 U36 ( .A1(in_18), .A2(in[93]), .ZN(n930) );
  AND2_X1 U36bar ( .A1(in_18bar), .A2(inbar[93]), .ZN(n930bar) );
  OR2_X1 U37 ( .A1(in_31), .A2(n929), .ZN(n931) );
  AND2_X1 U37bar ( .A1(in_31bar), .A2(n929bar), .ZN(n931bar) );
  OR2_X1 U38 ( .A1(in_7), .A2(in_39), .ZN(n929) );
  AND2_X1 U38bar ( .A1(in_7bar), .A2(in_39bar), .ZN(n929bar) );
  OR2_X1 U39 ( .A1(n928), .A2(n927), .ZN(out[5]) );
  AND2_X1 U39bar ( .A1(n928bar), .A2(n927bar), .ZN(outbar[5]) );
  OR2_X1 U40 ( .A1(n926), .A2(n925), .ZN(n927) );
  AND2_X1 U40bar ( .A1(n926bar), .A2(n925bar), .ZN(n927bar) );
  OR2_X1 U41 ( .A1(n924), .A2(n923), .ZN(n925) );
  AND2_X1 U41bar ( .A1(n924bar), .A2(n923bar), .ZN(n925bar) );
  OR2_X1 U42 ( .A1(n922), .A2(n921), .ZN(n923) );
  AND2_X1 U42bar ( .A1(n922bar), .A2(n921bar), .ZN(n923bar) );
  OR2_X1 U43 ( .A1(n940), .A2(n920), .ZN(n924) );
  AND2_X1 U43bar ( .A1(n940bar), .A2(n920bar), .ZN(n924bar) );
  OR2_X1 U44 ( .A1(in[111]), .A2(n919), .ZN(n920) );
  AND2_X1 U44bar ( .A1(inbar[111]), .A2(n919bar), .ZN(n920bar) );
  OR2_X1 U45 ( .A1(n918), .A2(n917), .ZN(n940) );
  AND2_X1 U45bar ( .A1(n918bar), .A2(n917bar), .ZN(n940bar) );
  OR2_X1 U46 ( .A1(n916), .A2(n915), .ZN(n917) );
  AND2_X1 U46bar ( .A1(n916bar), .A2(n915bar), .ZN(n917bar) );
  OR2_X1 U47 ( .A1(n914), .A2(n913), .ZN(n915) );
  AND2_X1 U47bar ( .A1(n914bar), .A2(n913bar), .ZN(n915bar) );
  OR2_X1 U48 ( .A1(in[140]), .A2(in[131]), .ZN(n913) );
  AND2_X1 U48bar ( .A1(inbar[140]), .A2(inbar[131]), .ZN(n913bar) );
  OR2_X1 U49 ( .A1(in[160]), .A2(in[144]), .ZN(n914) );
  AND2_X1 U49bar ( .A1(inbar[160]), .A2(inbar[144]), .ZN(n914bar) );
  OR2_X1 U50 ( .A1(n912), .A2(n911), .ZN(n916) );
  AND2_X1 U50bar ( .A1(n912bar), .A2(n911bar), .ZN(n916bar) );
  OR2_X1 U51 ( .A1(in[179]), .A2(in[174]), .ZN(n911) );
  AND2_X1 U51bar ( .A1(inbar[179]), .A2(inbar[174]), .ZN(n911bar) );
  OR2_X1 U52 ( .A1(in[188]), .A2(in[184]), .ZN(n912) );
  AND2_X1 U52bar ( .A1(inbar[188]), .A2(inbar[184]), .ZN(n912bar) );
  OR2_X1 U53 ( .A1(n910), .A2(n909), .ZN(n918) );
  AND2_X1 U53bar ( .A1(n910bar), .A2(n909bar), .ZN(n918bar) );
  OR2_X1 U54 ( .A1(n908), .A2(n907), .ZN(n909) );
  AND2_X1 U54bar ( .A1(n908bar), .A2(n907bar), .ZN(n909bar) );
  OR2_X1 U55 ( .A1(in[216]), .A2(in[200]), .ZN(n907) );
  AND2_X1 U55bar ( .A1(inbar[216]), .A2(inbar[200]), .ZN(n907bar) );
  OR2_X1 U56 ( .A1(in[228]), .A2(in[224]), .ZN(n908) );
  AND2_X1 U56bar ( .A1(inbar[228]), .A2(inbar[224]), .ZN(n908bar) );
  OR2_X1 U57 ( .A1(n906), .A2(n905), .ZN(n910) );
  AND2_X1 U57bar ( .A1(n906bar), .A2(n905bar), .ZN(n910bar) );
  OR2_X1 U58 ( .A1(in[247]), .A2(in[235]), .ZN(n905) );
  AND2_X1 U58bar ( .A1(inbar[247]), .A2(inbar[235]), .ZN(n905bar) );
  OR2_X1 U59 ( .A1(in_42), .A2(in[83]), .ZN(n906) );
  AND2_X1 U59bar ( .A1(in_42bar), .A2(inbar[83]), .ZN(n906bar) );
  OR2_X1 U60 ( .A1(n904), .A2(n903), .ZN(n926) );
  AND2_X1 U60bar ( .A1(n904bar), .A2(n903bar), .ZN(n926bar) );
  OR2_X1 U61 ( .A1(in[166]), .A2(in[123]), .ZN(n903) );
  AND2_X1 U61bar ( .A1(inbar[166]), .A2(inbar[123]), .ZN(n903bar) );
  OR2_X1 U62 ( .A1(in[170]), .A2(n902), .ZN(n904) );
  AND2_X1 U62bar ( .A1(inbar[170]), .A2(n902bar), .ZN(n904bar) );
  OR2_X1 U63 ( .A1(in[194]), .A2(in[183]), .ZN(n902) );
  AND2_X1 U63bar ( .A1(inbar[194]), .A2(inbar[183]), .ZN(n902bar) );
  OR2_X1 U64 ( .A1(n901), .A2(n900), .ZN(n928) );
  AND2_X1 U64bar ( .A1(n901bar), .A2(n900bar), .ZN(n928bar) );
  OR2_X1 U65 ( .A1(n899), .A2(n898), .ZN(n900) );
  AND2_X1 U65bar ( .A1(n899bar), .A2(n898bar), .ZN(n900bar) );
  OR2_X1 U66 ( .A1(in[241]), .A2(in[238]), .ZN(n898) );
  AND2_X1 U66bar ( .A1(inbar[241]), .A2(inbar[238]), .ZN(n898bar) );
  OR2_X1 U67 ( .A1(in[250]), .A2(n897), .ZN(n899) );
  AND2_X1 U67bar ( .A1(inbar[250]), .A2(n897bar), .ZN(n899bar) );
  OR2_X1 U68 ( .A1(in_24), .A2(in[84]), .ZN(n897) );
  AND2_X1 U68bar ( .A1(in_24bar), .A2(inbar[84]), .ZN(n897bar) );
  OR2_X1 U69 ( .A1(n896), .A2(n895), .ZN(n901) );
  AND2_X1 U69bar ( .A1(n896bar), .A2(n895bar), .ZN(n901bar) );
  OR2_X1 U70 ( .A1(in_41), .A2(in_29), .ZN(n895) );
  AND2_X1 U70bar ( .A1(in_41bar), .A2(in_29bar), .ZN(n895bar) );
  OR2_X1 U71 ( .A1(in_66), .A2(n894), .ZN(n896) );
  AND2_X1 U71bar ( .A1(in_66bar), .A2(n894bar), .ZN(n896bar) );
  OR2_X1 U72 ( .A1(in_76), .A2(in_71), .ZN(n894) );
  AND2_X1 U72bar ( .A1(in_76bar), .A2(in_71bar), .ZN(n894bar) );
  OR2_X1 U73 ( .A1(n893), .A2(n892), .ZN(out[4]) );
  AND2_X1 U73bar ( .A1(n893bar), .A2(n892bar), .ZN(outbar[4]) );
  OR2_X1 U74 ( .A1(n891), .A2(n890), .ZN(n892) );
  AND2_X1 U74bar ( .A1(n891bar), .A2(n890bar), .ZN(n892bar) );
  OR2_X1 U75 ( .A1(n889), .A2(n888), .ZN(n890) );
  AND2_X1 U75bar ( .A1(n889bar), .A2(n888bar), .ZN(n890bar) );
  OR2_X1 U76 ( .A1(n922), .A2(n887), .ZN(n888) );
  AND2_X1 U76bar ( .A1(n922bar), .A2(n887bar), .ZN(n888bar) );
  OR2_X1 U77 ( .A1(n886), .A2(n885), .ZN(n922) );
  AND2_X1 U77bar ( .A1(n886bar), .A2(n885bar), .ZN(n922bar) );
  OR2_X1 U78 ( .A1(n884), .A2(n883), .ZN(n885) );
  AND2_X1 U78bar ( .A1(n884bar), .A2(n883bar), .ZN(n885bar) );
  OR2_X1 U79 ( .A1(n882), .A2(n881), .ZN(n883) );
  AND2_X1 U79bar ( .A1(n882bar), .A2(n881bar), .ZN(n883bar) );
  OR2_X1 U80 ( .A1(in[118]), .A2(in[109]), .ZN(n881) );
  AND2_X1 U80bar ( .A1(inbar[118]), .A2(inbar[109]), .ZN(n881bar) );
  OR2_X1 U81 ( .A1(in[139]), .A2(in[120]), .ZN(n882) );
  AND2_X1 U81bar ( .A1(inbar[139]), .A2(inbar[120]), .ZN(n882bar) );
  OR2_X1 U82 ( .A1(n880), .A2(n879), .ZN(n884) );
  AND2_X1 U82bar ( .A1(n880bar), .A2(n879bar), .ZN(n884bar) );
  OR2_X1 U83 ( .A1(in[198]), .A2(in[154]), .ZN(n879) );
  AND2_X1 U83bar ( .A1(inbar[198]), .A2(inbar[154]), .ZN(n879bar) );
  OR2_X1 U84 ( .A1(in[210]), .A2(in[205]), .ZN(n880) );
  AND2_X1 U84bar ( .A1(inbar[210]), .A2(inbar[205]), .ZN(n880bar) );
  OR2_X1 U85 ( .A1(n878), .A2(n877), .ZN(n886) );
  AND2_X1 U85bar ( .A1(n878bar), .A2(n877bar), .ZN(n886bar) );
  OR2_X1 U86 ( .A1(n876), .A2(n875), .ZN(n877) );
  AND2_X1 U86bar ( .A1(n876bar), .A2(n875bar), .ZN(n877bar) );
  OR2_X1 U87 ( .A1(in[219]), .A2(in[217]), .ZN(n875) );
  AND2_X1 U87bar ( .A1(inbar[219]), .A2(inbar[217]), .ZN(n875bar) );
  OR2_X1 U88 ( .A1(in[86]), .A2(in[252]), .ZN(n876) );
  AND2_X1 U88bar ( .A1(inbar[86]), .A2(inbar[252]), .ZN(n876bar) );
  OR2_X1 U89 ( .A1(n874), .A2(n873), .ZN(n878) );
  AND2_X1 U89bar ( .A1(n874bar), .A2(n873bar), .ZN(n878bar) );
  OR2_X1 U90 ( .A1(in_40), .A2(in[91]), .ZN(n873) );
  AND2_X1 U90bar ( .A1(in_40bar), .A2(inbar[91]), .ZN(n873bar) );
  OR2_X1 U91 ( .A1(in_8), .A2(in_46), .ZN(n874) );
  AND2_X1 U91bar ( .A1(in_8bar), .A2(in_46bar), .ZN(n874bar) );
  OR2_X1 U92 ( .A1(n872), .A2(n871), .ZN(n889) );
  AND2_X1 U92bar ( .A1(n872bar), .A2(n871bar), .ZN(n889bar) );
  OR2_X1 U93 ( .A1(in[117]), .A2(n943), .ZN(n871) );
  AND2_X1 U93bar ( .A1(inbar[117]), .A2(n943bar), .ZN(n871bar) );
  OR2_X1 U94 ( .A1(n870), .A2(n869), .ZN(n943) );
  AND2_X1 U94bar ( .A1(n870bar), .A2(n869bar), .ZN(n943bar) );
  OR2_X1 U95 ( .A1(n868), .A2(n867), .ZN(n869) );
  AND2_X1 U95bar ( .A1(n868bar), .A2(n867bar), .ZN(n869bar) );
  OR2_X1 U96 ( .A1(n866), .A2(n865), .ZN(n867) );
  AND2_X1 U96bar ( .A1(n866bar), .A2(n865bar), .ZN(n867bar) );
  OR2_X1 U97 ( .A1(n864), .A2(n863), .ZN(n865) );
  AND2_X1 U97bar ( .A1(n864bar), .A2(n863bar), .ZN(n865bar) );
  OR2_X1 U98 ( .A1(in[108]), .A2(n919), .ZN(n866) );
  AND2_X1 U98bar ( .A1(inbar[108]), .A2(n919bar), .ZN(n866bar) );
  OR2_X1 U99 ( .A1(n862), .A2(n861), .ZN(n919) );
  AND2_X1 U99bar ( .A1(n862bar), .A2(n861bar), .ZN(n919bar) );
  OR2_X1 U100 ( .A1(n860), .A2(n859), .ZN(n861) );
  AND2_X1 U100bar ( .A1(n860bar), .A2(n859bar), .ZN(n861bar) );
  OR2_X1 U101 ( .A1(n858), .A2(n857), .ZN(n859) );
  AND2_X1 U101bar ( .A1(n858bar), .A2(n857bar), .ZN(n859bar) );
  OR2_X1 U102 ( .A1(in[119]), .A2(in[105]), .ZN(n857) );
  AND2_X1 U102bar ( .A1(inbar[119]), .A2(inbar[105]), .ZN(n857bar) );
  OR2_X1 U103 ( .A1(in[186]), .A2(in[175]), .ZN(n858) );
  AND2_X1 U103bar ( .A1(inbar[186]), .A2(inbar[175]), .ZN(n858bar) );
  OR2_X1 U104 ( .A1(n856), .A2(n855), .ZN(n860) );
  AND2_X1 U104bar ( .A1(n856bar), .A2(n855bar), .ZN(n860bar) );
  OR2_X1 U105 ( .A1(in[202]), .A2(in[193]), .ZN(n855) );
  AND2_X1 U105bar ( .A1(inbar[202]), .A2(inbar[193]), .ZN(n855bar) );
  OR2_X1 U106 ( .A1(in[225]), .A2(in[208]), .ZN(n856) );
  AND2_X1 U106bar ( .A1(inbar[225]), .A2(inbar[208]), .ZN(n856bar) );
  OR2_X1 U107 ( .A1(n854), .A2(n853), .ZN(n862) );
  AND2_X1 U107bar ( .A1(n854bar), .A2(n853bar), .ZN(n862bar) );
  OR2_X1 U108 ( .A1(n852), .A2(n851), .ZN(n853) );
  AND2_X1 U108bar ( .A1(n852bar), .A2(n851bar), .ZN(n853bar) );
  OR2_X1 U109 ( .A1(in_1), .A2(in[85]), .ZN(n851) );
  AND2_X1 U109bar ( .A1(in_1bar), .A2(inbar[85]), .ZN(n851bar) );
  OR2_X1 U110 ( .A1(in_23), .A2(in_19), .ZN(n852) );
  AND2_X1 U110bar ( .A1(in_23bar), .A2(in_19bar), .ZN(n852bar) );
  OR2_X1 U111 ( .A1(n850), .A2(n849), .ZN(n854) );
  AND2_X1 U111bar ( .A1(n850bar), .A2(n849bar), .ZN(n854bar) );
  OR2_X1 U112 ( .A1(in_43), .A2(in_33), .ZN(n849) );
  AND2_X1 U112bar ( .A1(in_43bar), .A2(in_33bar), .ZN(n849bar) );
  OR2_X1 U113 ( .A1(in_63), .A2(in_44), .ZN(n850) );
  AND2_X1 U113bar ( .A1(in_63bar), .A2(in_44bar), .ZN(n850bar) );
  OR2_X1 U114 ( .A1(n848), .A2(n847), .ZN(n868) );
  AND2_X1 U114bar ( .A1(n848bar), .A2(n847bar), .ZN(n868bar) );
  OR2_X1 U115 ( .A1(in[141]), .A2(in[112]), .ZN(n847) );
  AND2_X1 U115bar ( .A1(inbar[141]), .A2(inbar[112]), .ZN(n847bar) );
  OR2_X1 U116 ( .A1(in[147]), .A2(n846), .ZN(n848) );
  AND2_X1 U116bar ( .A1(inbar[147]), .A2(n846bar), .ZN(n848bar) );
  OR2_X1 U117 ( .A1(in[181]), .A2(in[167]), .ZN(n846) );
  AND2_X1 U117bar ( .A1(inbar[181]), .A2(inbar[167]), .ZN(n846bar) );
  OR2_X1 U118 ( .A1(n845), .A2(n844), .ZN(n870) );
  AND2_X1 U118bar ( .A1(n845bar), .A2(n844bar), .ZN(n870bar) );
  OR2_X1 U119 ( .A1(n843), .A2(n842), .ZN(n844) );
  AND2_X1 U119bar ( .A1(n843bar), .A2(n842bar), .ZN(n844bar) );
  OR2_X1 U120 ( .A1(in[229]), .A2(in[201]), .ZN(n842) );
  AND2_X1 U120bar ( .A1(inbar[229]), .A2(inbar[201]), .ZN(n842bar) );
  OR2_X1 U121 ( .A1(in[237]), .A2(n841), .ZN(n843) );
  AND2_X1 U121bar ( .A1(inbar[237]), .A2(n841bar), .ZN(n843bar) );
  OR2_X1 U122 ( .A1(in[94]), .A2(in[253]), .ZN(n841) );
  AND2_X1 U122bar ( .A1(inbar[94]), .A2(inbar[253]), .ZN(n841bar) );
  OR2_X1 U123 ( .A1(n840), .A2(n839), .ZN(n845) );
  AND2_X1 U123bar ( .A1(n840bar), .A2(n839bar), .ZN(n845bar) );
  OR2_X1 U124 ( .A1(in_21), .A2(in[96]), .ZN(n839) );
  AND2_X1 U124bar ( .A1(in_21bar), .A2(inbar[96]), .ZN(n839bar) );
  OR2_X1 U125 ( .A1(in_25), .A2(n838), .ZN(n840) );
  AND2_X1 U125bar ( .A1(in_25bar), .A2(n838bar), .ZN(n840bar) );
  OR2_X1 U126 ( .A1(in_81), .A2(in_45), .ZN(n838) );
  AND2_X1 U126bar ( .A1(in_81bar), .A2(in_45bar), .ZN(n838bar) );
  OR2_X1 U127 ( .A1(n837), .A2(n836), .ZN(n891) );
  AND2_X1 U127bar ( .A1(n837bar), .A2(n836bar), .ZN(n891bar) );
  OR2_X1 U128 ( .A1(in[142]), .A2(in[124]), .ZN(n836) );
  AND2_X1 U128bar ( .A1(inbar[142]), .A2(inbar[124]), .ZN(n836bar) );
  OR2_X1 U129 ( .A1(in[150]), .A2(n835), .ZN(n837) );
  AND2_X1 U129bar ( .A1(inbar[150]), .A2(n835bar), .ZN(n837bar) );
  OR2_X1 U130 ( .A1(in[172]), .A2(in[155]), .ZN(n835) );
  AND2_X1 U130bar ( .A1(inbar[172]), .A2(inbar[155]), .ZN(n835bar) );
  OR2_X1 U131 ( .A1(n834), .A2(n833), .ZN(n893) );
  AND2_X1 U131bar ( .A1(n834bar), .A2(n833bar), .ZN(n893bar) );
  OR2_X1 U132 ( .A1(n832), .A2(n831), .ZN(n833) );
  AND2_X1 U132bar ( .A1(n832bar), .A2(n831bar), .ZN(n833bar) );
  OR2_X1 U133 ( .A1(in[196]), .A2(in[173]), .ZN(n831) );
  AND2_X1 U133bar ( .A1(inbar[196]), .A2(inbar[173]), .ZN(n831bar) );
  OR2_X1 U134 ( .A1(in[222]), .A2(n830), .ZN(n832) );
  AND2_X1 U134bar ( .A1(inbar[222]), .A2(n830bar), .ZN(n832bar) );
  OR2_X1 U135 ( .A1(in[227]), .A2(in[226]), .ZN(n830) );
  AND2_X1 U135bar ( .A1(inbar[227]), .A2(inbar[226]), .ZN(n830bar) );
  OR2_X1 U136 ( .A1(n829), .A2(n828), .ZN(n834) );
  AND2_X1 U136bar ( .A1(n829bar), .A2(n828bar), .ZN(n834bar) );
  OR2_X1 U137 ( .A1(in[249]), .A2(in[231]), .ZN(n828) );
  AND2_X1 U137bar ( .A1(inbar[249]), .A2(inbar[231]), .ZN(n828bar) );
  OR2_X1 U138 ( .A1(in_28), .A2(n827), .ZN(n829) );
  AND2_X1 U138bar ( .A1(in_28bar), .A2(n827bar), .ZN(n829bar) );
  OR2_X1 U139 ( .A1(in_52), .A2(in_47), .ZN(n827) );
  AND2_X1 U139bar ( .A1(in_52bar), .A2(in_47bar), .ZN(n827bar) );
  OR2_X1 U140 ( .A1(n826), .A2(n825), .ZN(out[3]) );
  AND2_X1 U140bar ( .A1(n826bar), .A2(n825bar), .ZN(outbar[3]) );
  OR2_X1 U141 ( .A1(n824), .A2(n823), .ZN(n825) );
  AND2_X1 U141bar ( .A1(n824bar), .A2(n823bar), .ZN(n825bar) );
  OR2_X1 U142 ( .A1(n822), .A2(n821), .ZN(n823) );
  AND2_X1 U142bar ( .A1(n822bar), .A2(n821bar), .ZN(n823bar) );
  OR2_X1 U143 ( .A1(n820), .A2(n819), .ZN(n821) );
  AND2_X1 U143bar ( .A1(n820bar), .A2(n819bar), .ZN(n821bar) );
  OR2_X1 U144 ( .A1(n964), .A2(n818), .ZN(n822) );
  AND2_X1 U144bar ( .A1(n964bar), .A2(n818bar), .ZN(n822bar) );
  OR2_X1 U145 ( .A1(in[118]), .A2(n817), .ZN(n818) );
  AND2_X1 U145bar ( .A1(inbar[118]), .A2(n817bar), .ZN(n818bar) );
  OR2_X1 U146 ( .A1(n816), .A2(n815), .ZN(n964) );
  AND2_X1 U146bar ( .A1(n816bar), .A2(n815bar), .ZN(n964bar) );
  OR2_X1 U147 ( .A1(n814), .A2(n813), .ZN(n815) );
  AND2_X1 U147bar ( .A1(n814bar), .A2(n813bar), .ZN(n815bar) );
  OR2_X1 U148 ( .A1(n812), .A2(n811), .ZN(n813) );
  AND2_X1 U148bar ( .A1(n812bar), .A2(n811bar), .ZN(n813bar) );
  OR2_X1 U149 ( .A1(in[122]), .A2(in[111]), .ZN(n811) );
  AND2_X1 U149bar ( .A1(inbar[122]), .A2(inbar[111]), .ZN(n811bar) );
  OR2_X1 U150 ( .A1(in[154]), .A2(in[151]), .ZN(n812) );
  AND2_X1 U150bar ( .A1(inbar[154]), .A2(inbar[151]), .ZN(n812bar) );
  OR2_X1 U151 ( .A1(n810), .A2(n809), .ZN(n814) );
  AND2_X1 U151bar ( .A1(n810bar), .A2(n809bar), .ZN(n814bar) );
  OR2_X1 U152 ( .A1(in[187]), .A2(in[177]), .ZN(n809) );
  AND2_X1 U152bar ( .A1(inbar[187]), .A2(inbar[177]), .ZN(n809bar) );
  OR2_X1 U153 ( .A1(in[200]), .A2(in[192]), .ZN(n810) );
  AND2_X1 U153bar ( .A1(inbar[200]), .A2(inbar[192]), .ZN(n810bar) );
  OR2_X1 U154 ( .A1(n808), .A2(n807), .ZN(n816) );
  AND2_X1 U154bar ( .A1(n808bar), .A2(n807bar), .ZN(n816bar) );
  OR2_X1 U155 ( .A1(n806), .A2(n805), .ZN(n807) );
  AND2_X1 U155bar ( .A1(n806bar), .A2(n805bar), .ZN(n807bar) );
  OR2_X1 U156 ( .A1(in[225]), .A2(in[207]), .ZN(n805) );
  AND2_X1 U156bar ( .A1(inbar[225]), .A2(inbar[207]), .ZN(n805bar) );
  OR2_X1 U157 ( .A1(in[98]), .A2(in[226]), .ZN(n806) );
  AND2_X1 U157bar ( .A1(inbar[98]), .A2(inbar[226]), .ZN(n806bar) );
  OR2_X1 U158 ( .A1(n804), .A2(n803), .ZN(n808) );
  AND2_X1 U158bar ( .A1(n804bar), .A2(n803bar), .ZN(n808bar) );
  OR2_X1 U159 ( .A1(in_20), .A2(in_16), .ZN(n803) );
  AND2_X1 U159bar ( .A1(in_20bar), .A2(in_16bar), .ZN(n803bar) );
  OR2_X1 U160 ( .A1(in_55), .A2(in_45), .ZN(n804) );
  AND2_X1 U160bar ( .A1(in_55bar), .A2(in_45bar), .ZN(n804bar) );
  OR2_X1 U161 ( .A1(n802), .A2(n801), .ZN(n824) );
  AND2_X1 U161bar ( .A1(n802bar), .A2(n801bar), .ZN(n824bar) );
  OR2_X1 U162 ( .A1(in[162]), .A2(in[149]), .ZN(n801) );
  AND2_X1 U162bar ( .A1(inbar[162]), .A2(inbar[149]), .ZN(n801bar) );
  OR2_X1 U163 ( .A1(in[163]), .A2(n800), .ZN(n802) );
  AND2_X1 U163bar ( .A1(inbar[163]), .A2(n800bar), .ZN(n802bar) );
  OR2_X1 U164 ( .A1(in[191]), .A2(in[189]), .ZN(n800) );
  AND2_X1 U164bar ( .A1(inbar[191]), .A2(inbar[189]), .ZN(n800bar) );
  OR2_X1 U165 ( .A1(n799), .A2(n798), .ZN(n826) );
  AND2_X1 U165bar ( .A1(n799bar), .A2(n798bar), .ZN(n826bar) );
  OR2_X1 U166 ( .A1(n797), .A2(n796), .ZN(n798) );
  AND2_X1 U166bar ( .A1(n797bar), .A2(n796bar), .ZN(n798bar) );
  OR2_X1 U167 ( .A1(in[212]), .A2(in[193]), .ZN(n796) );
  AND2_X1 U167bar ( .A1(inbar[212]), .A2(inbar[193]), .ZN(n796bar) );
  OR2_X1 U168 ( .A1(in[238]), .A2(n795), .ZN(n797) );
  AND2_X1 U168bar ( .A1(inbar[238]), .A2(n795bar), .ZN(n797bar) );
  OR2_X1 U169 ( .A1(in[88]), .A2(in[247]), .ZN(n795) );
  AND2_X1 U169bar ( .A1(inbar[88]), .A2(inbar[247]), .ZN(n795bar) );
  OR2_X1 U170 ( .A1(n794), .A2(n793), .ZN(n799) );
  AND2_X1 U170bar ( .A1(n794bar), .A2(n793bar), .ZN(n799bar) );
  OR2_X1 U171 ( .A1(in[94]), .A2(in[92]), .ZN(n793) );
  AND2_X1 U171bar ( .A1(inbar[94]), .A2(inbar[92]), .ZN(n793bar) );
  OR2_X1 U172 ( .A1(in_52), .A2(n792), .ZN(n794) );
  AND2_X1 U172bar ( .A1(in_52bar), .A2(n792bar), .ZN(n794bar) );
  OR2_X1 U173 ( .A1(in_70), .A2(in_67), .ZN(n792) );
  AND2_X1 U173bar ( .A1(in_70bar), .A2(in_67bar), .ZN(n792bar) );
  OR2_X1 U174 ( .A1(n791), .A2(n790), .ZN(out[2]) );
  AND2_X1 U174bar ( .A1(n791bar), .A2(n790bar), .ZN(outbar[2]) );
  OR2_X1 U175 ( .A1(n789), .A2(n788), .ZN(n790) );
  AND2_X1 U175bar ( .A1(n789bar), .A2(n788bar), .ZN(n790bar) );
  OR2_X1 U176 ( .A1(n787), .A2(n786), .ZN(n788) );
  AND2_X1 U176bar ( .A1(n787bar), .A2(n786bar), .ZN(n788bar) );
  OR2_X1 U177 ( .A1(n819), .A2(n785), .ZN(n786) );
  AND2_X1 U177bar ( .A1(n819bar), .A2(n785bar), .ZN(n786bar) );
  OR2_X1 U178 ( .A1(n784), .A2(n783), .ZN(n819) );
  AND2_X1 U178bar ( .A1(n784bar), .A2(n783bar), .ZN(n819bar) );
  OR2_X1 U179 ( .A1(n782), .A2(n781), .ZN(n783) );
  AND2_X1 U179bar ( .A1(n782bar), .A2(n781bar), .ZN(n783bar) );
  OR2_X1 U180 ( .A1(n780), .A2(n779), .ZN(n781) );
  AND2_X1 U180bar ( .A1(n780bar), .A2(n779bar), .ZN(n781bar) );
  OR2_X1 U181 ( .A1(n962), .A2(n778), .ZN(n779) );
  AND2_X1 U181bar ( .A1(n962bar), .A2(n778bar), .ZN(n779bar) );
  OR2_X1 U182 ( .A1(n777), .A2(n776), .ZN(n962) );
  AND2_X1 U182bar ( .A1(n777bar), .A2(n776bar), .ZN(n962bar) );
  OR2_X1 U183 ( .A1(n775), .A2(n774), .ZN(n776) );
  AND2_X1 U183bar ( .A1(n775bar), .A2(n774bar), .ZN(n776bar) );
  OR2_X1 U184 ( .A1(n773), .A2(n772), .ZN(n774) );
  AND2_X1 U184bar ( .A1(n773bar), .A2(n772bar), .ZN(n774bar) );
  OR2_X1 U185 ( .A1(in[131]), .A2(in[120]), .ZN(n772) );
  AND2_X1 U185bar ( .A1(inbar[131]), .A2(inbar[120]), .ZN(n772bar) );
  OR2_X1 U186 ( .A1(in[153]), .A2(in[147]), .ZN(n773) );
  AND2_X1 U186bar ( .A1(inbar[153]), .A2(inbar[147]), .ZN(n773bar) );
  OR2_X1 U187 ( .A1(n771), .A2(n770), .ZN(n775) );
  AND2_X1 U187bar ( .A1(n771bar), .A2(n770bar), .ZN(n775bar) );
  OR2_X1 U188 ( .A1(in[170]), .A2(in[156]), .ZN(n770) );
  AND2_X1 U188bar ( .A1(inbar[170]), .A2(inbar[156]), .ZN(n770bar) );
  OR2_X1 U189 ( .A1(in[223]), .A2(in[190]), .ZN(n771) );
  AND2_X1 U189bar ( .A1(inbar[223]), .A2(inbar[190]), .ZN(n771bar) );
  OR2_X1 U190 ( .A1(n769), .A2(n768), .ZN(n777) );
  AND2_X1 U190bar ( .A1(n769bar), .A2(n768bar), .ZN(n777bar) );
  OR2_X1 U191 ( .A1(n767), .A2(n766), .ZN(n768) );
  AND2_X1 U191bar ( .A1(n767bar), .A2(n766bar), .ZN(n768bar) );
  OR2_X1 U192 ( .A1(in[236]), .A2(in[230]), .ZN(n766) );
  AND2_X1 U192bar ( .A1(inbar[236]), .A2(inbar[230]), .ZN(n766bar) );
  OR2_X1 U193 ( .A1(in[85]), .A2(in[240]), .ZN(n767) );
  AND2_X1 U193bar ( .A1(inbar[85]), .A2(inbar[240]), .ZN(n767bar) );
  OR2_X1 U194 ( .A1(n765), .A2(n764), .ZN(n769) );
  AND2_X1 U194bar ( .A1(n765bar), .A2(n764bar), .ZN(n769bar) );
  OR2_X1 U195 ( .A1(in_12), .A2(in[90]), .ZN(n764) );
  AND2_X1 U195bar ( .A1(in_12bar), .A2(inbar[90]), .ZN(n764bar) );
  OR2_X1 U196 ( .A1(in_39), .A2(in_28), .ZN(n765) );
  AND2_X1 U196bar ( .A1(in_39bar), .A2(in_28bar), .ZN(n765bar) );
  OR2_X1 U197 ( .A1(in[109]), .A2(n763), .ZN(n780) );
  AND2_X1 U197bar ( .A1(inbar[109]), .A2(n763bar), .ZN(n780bar) );
  OR2_X1 U198 ( .A1(n762), .A2(n761), .ZN(n782) );
  AND2_X1 U198bar ( .A1(n762bar), .A2(n761bar), .ZN(n782bar) );
  OR2_X1 U199 ( .A1(in[138]), .A2(in[129]), .ZN(n761) );
  AND2_X1 U199bar ( .A1(inbar[138]), .A2(inbar[129]), .ZN(n761bar) );
  OR2_X1 U200 ( .A1(in[157]), .A2(n760), .ZN(n762) );
  AND2_X1 U200bar ( .A1(inbar[157]), .A2(n760bar), .ZN(n762bar) );
  OR2_X1 U201 ( .A1(in[182]), .A2(in[167]), .ZN(n760) );
  AND2_X1 U201bar ( .A1(inbar[182]), .A2(inbar[167]), .ZN(n760bar) );
  OR2_X1 U202 ( .A1(n759), .A2(n758), .ZN(n784) );
  AND2_X1 U202bar ( .A1(n759bar), .A2(n758bar), .ZN(n784bar) );
  OR2_X1 U203 ( .A1(n757), .A2(n756), .ZN(n758) );
  AND2_X1 U203bar ( .A1(n757bar), .A2(n756bar), .ZN(n758bar) );
  OR2_X1 U204 ( .A1(in[195]), .A2(in[184]), .ZN(n756) );
  AND2_X1 U204bar ( .A1(inbar[195]), .A2(inbar[184]), .ZN(n756bar) );
  OR2_X1 U205 ( .A1(in[196]), .A2(n755), .ZN(n757) );
  AND2_X1 U205bar ( .A1(inbar[196]), .A2(n755bar), .ZN(n757bar) );
  OR2_X1 U206 ( .A1(in[215]), .A2(in[209]), .ZN(n755) );
  AND2_X1 U206bar ( .A1(inbar[215]), .A2(inbar[209]), .ZN(n755bar) );
  OR2_X1 U207 ( .A1(n754), .A2(n753), .ZN(n759) );
  AND2_X1 U207bar ( .A1(n754bar), .A2(n753bar), .ZN(n759bar) );
  OR2_X1 U208 ( .A1(in[93]), .A2(in[233]), .ZN(n753) );
  AND2_X1 U208bar ( .A1(inbar[93]), .A2(inbar[233]), .ZN(n753bar) );
  OR2_X1 U209 ( .A1(in_1), .A2(n752), .ZN(n754) );
  AND2_X1 U209bar ( .A1(in_1bar), .A2(n752bar), .ZN(n754bar) );
  OR2_X1 U210 ( .A1(in_69), .A2(in_66), .ZN(n752) );
  AND2_X1 U210bar ( .A1(in_69bar), .A2(in_66bar), .ZN(n752bar) );
  OR2_X1 U211 ( .A1(n966), .A2(n751), .ZN(n787) );
  AND2_X1 U211bar ( .A1(n966bar), .A2(n751bar), .ZN(n787bar) );
  OR2_X1 U212 ( .A1(in[134]), .A2(n750), .ZN(n751) );
  AND2_X1 U212bar ( .A1(inbar[134]), .A2(n750bar), .ZN(n751bar) );
  OR2_X1 U213 ( .A1(n749), .A2(n748), .ZN(n966) );
  AND2_X1 U213bar ( .A1(n749bar), .A2(n748bar), .ZN(n966bar) );
  OR2_X1 U214 ( .A1(n747), .A2(n746), .ZN(n748) );
  AND2_X1 U214bar ( .A1(n747bar), .A2(n746bar), .ZN(n748bar) );
  OR2_X1 U215 ( .A1(n745), .A2(n744), .ZN(n746) );
  AND2_X1 U215bar ( .A1(n745bar), .A2(n744bar), .ZN(n746bar) );
  OR2_X1 U216 ( .A1(in[136]), .A2(in[121]), .ZN(n744) );
  AND2_X1 U216bar ( .A1(inbar[136]), .A2(inbar[121]), .ZN(n744bar) );
  OR2_X1 U217 ( .A1(in[186]), .A2(in[174]), .ZN(n745) );
  AND2_X1 U217bar ( .A1(inbar[186]), .A2(inbar[174]), .ZN(n745bar) );
  OR2_X1 U218 ( .A1(n743), .A2(n742), .ZN(n747) );
  AND2_X1 U218bar ( .A1(n743bar), .A2(n742bar), .ZN(n747bar) );
  OR2_X1 U219 ( .A1(in[198]), .A2(in[197]), .ZN(n742) );
  AND2_X1 U219bar ( .A1(inbar[198]), .A2(inbar[197]), .ZN(n742bar) );
  OR2_X1 U220 ( .A1(in[214]), .A2(in[199]), .ZN(n743) );
  AND2_X1 U220bar ( .A1(inbar[214]), .A2(inbar[199]), .ZN(n743bar) );
  OR2_X1 U221 ( .A1(n741), .A2(n740), .ZN(n749) );
  AND2_X1 U221bar ( .A1(n741bar), .A2(n740bar), .ZN(n749bar) );
  OR2_X1 U222 ( .A1(n739), .A2(n738), .ZN(n740) );
  AND2_X1 U222bar ( .A1(n739bar), .A2(n738bar), .ZN(n740bar) );
  OR2_X1 U223 ( .A1(in[231]), .A2(in[220]), .ZN(n738) );
  AND2_X1 U223bar ( .A1(inbar[231]), .A2(inbar[220]), .ZN(n738bar) );
  OR2_X1 U224 ( .A1(in_25), .A2(in[245]), .ZN(n739) );
  AND2_X1 U224bar ( .A1(in_25bar), .A2(inbar[245]), .ZN(n739bar) );
  OR2_X1 U225 ( .A1(n737), .A2(n736), .ZN(n741) );
  AND2_X1 U225bar ( .A1(n737bar), .A2(n736bar), .ZN(n741bar) );
  OR2_X1 U226 ( .A1(in_53), .A2(in_29), .ZN(n736) );
  AND2_X1 U226bar ( .A1(in_53bar), .A2(in_29bar), .ZN(n736bar) );
  OR2_X1 U227 ( .A1(in_79), .A2(in_74), .ZN(n737) );
  AND2_X1 U227bar ( .A1(in_79bar), .A2(in_74bar), .ZN(n737bar) );
  OR2_X1 U228 ( .A1(n735), .A2(n734), .ZN(n789) );
  AND2_X1 U228bar ( .A1(n735bar), .A2(n734bar), .ZN(n789bar) );
  OR2_X1 U229 ( .A1(in[152]), .A2(in[140]), .ZN(n734) );
  AND2_X1 U229bar ( .A1(inbar[152]), .A2(inbar[140]), .ZN(n734bar) );
  OR2_X1 U230 ( .A1(in[155]), .A2(n733), .ZN(n735) );
  AND2_X1 U230bar ( .A1(inbar[155]), .A2(n733bar), .ZN(n735bar) );
  OR2_X1 U231 ( .A1(in[166]), .A2(in[165]), .ZN(n733) );
  AND2_X1 U231bar ( .A1(inbar[166]), .A2(inbar[165]), .ZN(n733bar) );
  OR2_X1 U232 ( .A1(n732), .A2(n731), .ZN(n791) );
  AND2_X1 U232bar ( .A1(n732bar), .A2(n731bar), .ZN(n791bar) );
  OR2_X1 U233 ( .A1(n730), .A2(n729), .ZN(n731) );
  AND2_X1 U233bar ( .A1(n730bar), .A2(n729bar), .ZN(n731bar) );
  OR2_X1 U234 ( .A1(in[202]), .A2(in[185]), .ZN(n729) );
  AND2_X1 U234bar ( .A1(inbar[202]), .A2(inbar[185]), .ZN(n729bar) );
  OR2_X1 U235 ( .A1(in[211]), .A2(n728), .ZN(n730) );
  AND2_X1 U235bar ( .A1(inbar[211]), .A2(n728bar), .ZN(n730bar) );
  OR2_X1 U236 ( .A1(in[255]), .A2(in[253]), .ZN(n728) );
  AND2_X1 U236bar ( .A1(inbar[255]), .A2(inbar[253]), .ZN(n728bar) );
  OR2_X1 U237 ( .A1(n727), .A2(n726), .ZN(n732) );
  AND2_X1 U237bar ( .A1(n727bar), .A2(n726bar), .ZN(n732bar) );
  OR2_X1 U238 ( .A1(in_35), .A2(in_15), .ZN(n726) );
  AND2_X1 U238bar ( .A1(in_35bar), .A2(in_15bar), .ZN(n726bar) );
  OR2_X1 U239 ( .A1(in_36), .A2(n725), .ZN(n727) );
  AND2_X1 U239bar ( .A1(in_36bar), .A2(n725bar), .ZN(n727bar) );
  OR2_X1 U240 ( .A1(in_48), .A2(in_40), .ZN(n725) );
  AND2_X1 U240bar ( .A1(in_48bar), .A2(in_40bar), .ZN(n725bar) );
  OR2_X1 U241 ( .A1(n724), .A2(n723), .ZN(out[1]) );
  AND2_X1 U241bar ( .A1(n724bar), .A2(n723bar), .ZN(outbar[1]) );
  OR2_X1 U242 ( .A1(n722), .A2(n721), .ZN(n723) );
  AND2_X1 U242bar ( .A1(n722bar), .A2(n721bar), .ZN(n723bar) );
  OR2_X1 U243 ( .A1(n720), .A2(n719), .ZN(n721) );
  AND2_X1 U243bar ( .A1(n720bar), .A2(n719bar), .ZN(n721bar) );
  OR2_X1 U244 ( .A1(n921), .A2(n887), .ZN(n719) );
  AND2_X1 U244bar ( .A1(n921bar), .A2(n887bar), .ZN(n719bar) );
  OR2_X1 U245 ( .A1(n718), .A2(n717), .ZN(n887) );
  AND2_X1 U245bar ( .A1(n718bar), .A2(n717bar), .ZN(n887bar) );
  OR2_X1 U246 ( .A1(n716), .A2(n715), .ZN(n717) );
  AND2_X1 U246bar ( .A1(n716bar), .A2(n715bar), .ZN(n717bar) );
  OR2_X1 U247 ( .A1(n714), .A2(n713), .ZN(n715) );
  AND2_X1 U247bar ( .A1(n714bar), .A2(n713bar), .ZN(n715bar) );
  OR2_X1 U248 ( .A1(in[116]), .A2(in[110]), .ZN(n713) );
  AND2_X1 U248bar ( .A1(inbar[116]), .A2(inbar[110]), .ZN(n713bar) );
  OR2_X1 U249 ( .A1(in[133]), .A2(in[130]), .ZN(n714) );
  AND2_X1 U249bar ( .A1(inbar[133]), .A2(inbar[130]), .ZN(n714bar) );
  OR2_X1 U250 ( .A1(n712), .A2(n711), .ZN(n716) );
  AND2_X1 U250bar ( .A1(n712bar), .A2(n711bar), .ZN(n716bar) );
  OR2_X1 U251 ( .A1(in[203]), .A2(in[135]), .ZN(n711) );
  AND2_X1 U251bar ( .A1(inbar[203]), .A2(inbar[135]), .ZN(n711bar) );
  OR2_X1 U252 ( .A1(in[232]), .A2(in[223]), .ZN(n712) );
  AND2_X1 U252bar ( .A1(inbar[232]), .A2(inbar[223]), .ZN(n712bar) );
  OR2_X1 U253 ( .A1(n710), .A2(n709), .ZN(n718) );
  AND2_X1 U253bar ( .A1(n710bar), .A2(n709bar), .ZN(n718bar) );
  OR2_X1 U254 ( .A1(n708), .A2(n707), .ZN(n709) );
  AND2_X1 U254bar ( .A1(n708bar), .A2(n707bar), .ZN(n709bar) );
  OR2_X1 U255 ( .A1(in[255]), .A2(in[233]), .ZN(n707) );
  AND2_X1 U255bar ( .A1(inbar[255]), .A2(inbar[233]), .ZN(n707bar) );
  OR2_X1 U256 ( .A1(in_53), .A2(in_34), .ZN(n708) );
  AND2_X1 U256bar ( .A1(in_53bar), .A2(in_34bar), .ZN(n708bar) );
  OR2_X1 U257 ( .A1(n706), .A2(n705), .ZN(n710) );
  AND2_X1 U257bar ( .A1(n706bar), .A2(n705bar), .ZN(n710bar) );
  OR2_X1 U258 ( .A1(in_57), .A2(in_55), .ZN(n705) );
  AND2_X1 U258bar ( .A1(in_57bar), .A2(in_55bar), .ZN(n705bar) );
  OR2_X1 U259 ( .A1(in_68), .A2(in_67), .ZN(n706) );
  AND2_X1 U259bar ( .A1(in_68bar), .A2(in_67bar), .ZN(n706bar) );
  OR2_X1 U260 ( .A1(n704), .A2(n703), .ZN(n921) );
  AND2_X1 U260bar ( .A1(n704bar), .A2(n703bar), .ZN(n921bar) );
  OR2_X1 U261 ( .A1(n702), .A2(n701), .ZN(n703) );
  AND2_X1 U261bar ( .A1(n702bar), .A2(n701bar), .ZN(n703bar) );
  OR2_X1 U262 ( .A1(n700), .A2(n699), .ZN(n701) );
  AND2_X1 U262bar ( .A1(n700bar), .A2(n699bar), .ZN(n701bar) );
  OR2_X1 U263 ( .A1(n944), .A2(n872), .ZN(n699) );
  AND2_X1 U263bar ( .A1(n944bar), .A2(n872bar), .ZN(n699bar) );
  OR2_X1 U264 ( .A1(n698), .A2(n697), .ZN(n872) );
  AND2_X1 U264bar ( .A1(n698bar), .A2(n697bar), .ZN(n872bar) );
  OR2_X1 U265 ( .A1(n696), .A2(n695), .ZN(n697) );
  AND2_X1 U265bar ( .A1(n696bar), .A2(n695bar), .ZN(n697bar) );
  OR2_X1 U266 ( .A1(n694), .A2(n693), .ZN(n695) );
  AND2_X1 U266bar ( .A1(n694bar), .A2(n693bar), .ZN(n695bar) );
  OR2_X1 U267 ( .A1(in[121]), .A2(in[102]), .ZN(n693) );
  AND2_X1 U267bar ( .A1(inbar[121]), .A2(inbar[102]), .ZN(n693bar) );
  OR2_X1 U268 ( .A1(in[162]), .A2(in[161]), .ZN(n694) );
  AND2_X1 U268bar ( .A1(inbar[162]), .A2(inbar[161]), .ZN(n694bar) );
  OR2_X1 U269 ( .A1(n692), .A2(n691), .ZN(n696) );
  AND2_X1 U269bar ( .A1(n692bar), .A2(n691bar), .ZN(n696bar) );
  OR2_X1 U270 ( .A1(in[192]), .A2(in[178]), .ZN(n691) );
  AND2_X1 U270bar ( .A1(inbar[192]), .A2(inbar[178]), .ZN(n691bar) );
  OR2_X1 U271 ( .A1(in[244]), .A2(in[209]), .ZN(n692) );
  AND2_X1 U271bar ( .A1(inbar[244]), .A2(inbar[209]), .ZN(n692bar) );
  OR2_X1 U272 ( .A1(n690), .A2(n689), .ZN(n698) );
  AND2_X1 U272bar ( .A1(n690bar), .A2(n689bar), .ZN(n698bar) );
  OR2_X1 U273 ( .A1(n688), .A2(n687), .ZN(n689) );
  AND2_X1 U273bar ( .A1(n688bar), .A2(n687bar), .ZN(n689bar) );
  OR2_X1 U274 ( .A1(in[90]), .A2(in[254]), .ZN(n687) );
  AND2_X1 U274bar ( .A1(inbar[90]), .A2(inbar[254]), .ZN(n687bar) );
  OR2_X1 U275 ( .A1(in_36), .A2(in_32), .ZN(n688) );
  AND2_X1 U275bar ( .A1(in_36bar), .A2(in_32bar), .ZN(n688bar) );
  OR2_X1 U276 ( .A1(n686), .A2(n685), .ZN(n690) );
  AND2_X1 U276bar ( .A1(n686bar), .A2(n685bar), .ZN(n690bar) );
  OR2_X1 U277 ( .A1(in_62), .A2(in_37), .ZN(n685) );
  AND2_X1 U277bar ( .A1(in_62bar), .A2(in_37bar), .ZN(n685bar) );
  OR2_X1 U278 ( .A1(in_75), .A2(in_73), .ZN(n686) );
  AND2_X1 U278bar ( .A1(in_75bar), .A2(in_73bar), .ZN(n686bar) );
  OR2_X1 U279 ( .A1(n684), .A2(n683), .ZN(n944) );
  AND2_X1 U279bar ( .A1(n684bar), .A2(n683bar), .ZN(n944bar) );
  OR2_X1 U280 ( .A1(n682), .A2(n681), .ZN(n683) );
  AND2_X1 U280bar ( .A1(n682bar), .A2(n681bar), .ZN(n683bar) );
  OR2_X1 U281 ( .A1(n680), .A2(n679), .ZN(n681) );
  AND2_X1 U281bar ( .A1(n680bar), .A2(n679bar), .ZN(n681bar) );
  OR2_X1 U282 ( .A1(in[171]), .A2(in[153]), .ZN(n679) );
  AND2_X1 U282bar ( .A1(inbar[171]), .A2(inbar[153]), .ZN(n679bar) );
  OR2_X1 U283 ( .A1(in[187]), .A2(in[176]), .ZN(n680) );
  AND2_X1 U283bar ( .A1(inbar[187]), .A2(inbar[176]), .ZN(n680bar) );
  OR2_X1 U284 ( .A1(n678), .A2(n677), .ZN(n682) );
  AND2_X1 U284bar ( .A1(n678bar), .A2(n677bar), .ZN(n682bar) );
  OR2_X1 U285 ( .A1(in[245]), .A2(in[211]), .ZN(n677) );
  AND2_X1 U285bar ( .A1(inbar[245]), .A2(inbar[211]), .ZN(n677bar) );
  OR2_X1 U286 ( .A1(in[97]), .A2(in[88]), .ZN(n678) );
  AND2_X1 U286bar ( .A1(inbar[97]), .A2(inbar[88]), .ZN(n678bar) );
  OR2_X1 U287 ( .A1(n676), .A2(n675), .ZN(n684) );
  AND2_X1 U287bar ( .A1(n676bar), .A2(n675bar), .ZN(n684bar) );
  OR2_X1 U288 ( .A1(n674), .A2(n673), .ZN(n675) );
  AND2_X1 U288bar ( .A1(n674bar), .A2(n673bar), .ZN(n675bar) );
  OR2_X1 U289 ( .A1(in_10), .A2(in_0), .ZN(n673) );
  AND2_X1 U289bar ( .A1(in_10bar), .A2(in_0bar), .ZN(n673bar) );
  OR2_X1 U290 ( .A1(in_59), .A2(in_5), .ZN(n674) );
  AND2_X1 U290bar ( .A1(in_59bar), .A2(in_5bar), .ZN(n674bar) );
  OR2_X1 U291 ( .A1(n672), .A2(n671), .ZN(n676) );
  AND2_X1 U291bar ( .A1(n672bar), .A2(n671bar), .ZN(n676bar) );
  OR2_X1 U292 ( .A1(in_60), .A2(in_6), .ZN(n671) );
  AND2_X1 U292bar ( .A1(in_60bar), .A2(in_6bar), .ZN(n671bar) );
  OR2_X1 U293 ( .A1(in_77), .A2(in_69), .ZN(n672) );
  AND2_X1 U293bar ( .A1(in_77bar), .A2(in_69bar), .ZN(n672bar) );
  OR2_X1 U294 ( .A1(in[113]), .A2(n864), .ZN(n700) );
  AND2_X1 U294bar ( .A1(inbar[113]), .A2(n864bar), .ZN(n700bar) );
  OR2_X1 U295 ( .A1(n670), .A2(n669), .ZN(n864) );
  AND2_X1 U295bar ( .A1(n670bar), .A2(n669bar), .ZN(n864bar) );
  OR2_X1 U296 ( .A1(n668), .A2(n667), .ZN(n669) );
  AND2_X1 U296bar ( .A1(n668bar), .A2(n667bar), .ZN(n669bar) );
  OR2_X1 U297 ( .A1(n666), .A2(n665), .ZN(n667) );
  AND2_X1 U297bar ( .A1(n666bar), .A2(n665bar), .ZN(n667bar) );
  OR2_X1 U298 ( .A1(in[125]), .A2(in[107]), .ZN(n665) );
  AND2_X1 U298bar ( .A1(inbar[125]), .A2(inbar[107]), .ZN(n665bar) );
  OR2_X1 U299 ( .A1(in[138]), .A2(in[126]), .ZN(n666) );
  AND2_X1 U299bar ( .A1(inbar[138]), .A2(inbar[126]), .ZN(n666bar) );
  OR2_X1 U300 ( .A1(n664), .A2(n663), .ZN(n668) );
  AND2_X1 U300bar ( .A1(n664bar), .A2(n663bar), .ZN(n668bar) );
  OR2_X1 U301 ( .A1(in[189]), .A2(in[143]), .ZN(n663) );
  AND2_X1 U301bar ( .A1(inbar[189]), .A2(inbar[143]), .ZN(n663bar) );
  OR2_X1 U302 ( .A1(in[99]), .A2(in[214]), .ZN(n664) );
  AND2_X1 U302bar ( .A1(inbar[99]), .A2(inbar[214]), .ZN(n664bar) );
  OR2_X1 U303 ( .A1(n662), .A2(n661), .ZN(n670) );
  AND2_X1 U303bar ( .A1(n662bar), .A2(n661bar), .ZN(n670bar) );
  OR2_X1 U304 ( .A1(n660), .A2(n659), .ZN(n661) );
  AND2_X1 U304bar ( .A1(n660bar), .A2(n659bar), .ZN(n661bar) );
  OR2_X1 U305 ( .A1(in_15), .A2(in_12), .ZN(n659) );
  AND2_X1 U305bar ( .A1(in_15bar), .A2(in_12bar), .ZN(n659bar) );
  OR2_X1 U306 ( .A1(in_20), .A2(in_2), .ZN(n660) );
  AND2_X1 U306bar ( .A1(in_20bar), .A2(in_2bar), .ZN(n660bar) );
  OR2_X1 U307 ( .A1(n658), .A2(n657), .ZN(n662) );
  AND2_X1 U307bar ( .A1(n658bar), .A2(n657bar), .ZN(n662bar) );
  OR2_X1 U308 ( .A1(in_30), .A2(in_3), .ZN(n657) );
  AND2_X1 U308bar ( .A1(in_30bar), .A2(in_3bar), .ZN(n657bar) );
  OR2_X1 U309 ( .A1(in_4), .A2(in_38), .ZN(n658) );
  AND2_X1 U309bar ( .A1(in_4bar), .A2(in_38bar), .ZN(n658bar) );
  OR2_X1 U310 ( .A1(n656), .A2(n655), .ZN(n702) );
  AND2_X1 U310bar ( .A1(n656bar), .A2(n655bar), .ZN(n702bar) );
  OR2_X1 U311 ( .A1(in[148]), .A2(in[137]), .ZN(n655) );
  AND2_X1 U311bar ( .A1(inbar[148]), .A2(inbar[137]), .ZN(n655bar) );
  OR2_X1 U312 ( .A1(in[149]), .A2(n654), .ZN(n656) );
  AND2_X1 U312bar ( .A1(inbar[149]), .A2(n654bar), .ZN(n656bar) );
  OR2_X1 U313 ( .A1(in[195]), .A2(in[190]), .ZN(n654) );
  AND2_X1 U313bar ( .A1(inbar[195]), .A2(inbar[190]), .ZN(n654bar) );
  OR2_X1 U314 ( .A1(n653), .A2(n652), .ZN(n704) );
  AND2_X1 U314bar ( .A1(n653bar), .A2(n652bar), .ZN(n704bar) );
  OR2_X1 U315 ( .A1(n651), .A2(n650), .ZN(n652) );
  AND2_X1 U315bar ( .A1(n651bar), .A2(n650bar), .ZN(n652bar) );
  OR2_X1 U316 ( .A1(in[98]), .A2(in[197]), .ZN(n650) );
  AND2_X1 U316bar ( .A1(inbar[98]), .A2(inbar[197]), .ZN(n650bar) );
  OR2_X1 U317 ( .A1(in_11), .A2(n649), .ZN(n651) );
  AND2_X1 U317bar ( .A1(in_11bar), .A2(n649bar), .ZN(n651bar) );
  OR2_X1 U318 ( .A1(in_26), .A2(in_14), .ZN(n649) );
  AND2_X1 U318bar ( .A1(in_26bar), .A2(in_14bar), .ZN(n649bar) );
  OR2_X1 U319 ( .A1(n648), .A2(n647), .ZN(n653) );
  AND2_X1 U319bar ( .A1(n648bar), .A2(n647bar), .ZN(n653bar) );
  OR2_X1 U320 ( .A1(in_35), .A2(in_27), .ZN(n647) );
  AND2_X1 U320bar ( .A1(in_35bar), .A2(in_27bar), .ZN(n647bar) );
  OR2_X1 U321 ( .A1(in_50), .A2(n646), .ZN(n648) );
  AND2_X1 U321bar ( .A1(in_50bar), .A2(n646bar), .ZN(n648bar) );
  OR2_X1 U322 ( .A1(in_78), .A2(in_61), .ZN(n646) );
  AND2_X1 U322bar ( .A1(in_78bar), .A2(in_61bar), .ZN(n646bar) );
  OR2_X1 U323 ( .A1(n942), .A2(n645), .ZN(n720) );
  AND2_X1 U323bar ( .A1(n942bar), .A2(n645bar), .ZN(n720bar) );
  OR2_X1 U324 ( .A1(in[106]), .A2(n863), .ZN(n645) );
  AND2_X1 U324bar ( .A1(inbar[106]), .A2(n863bar), .ZN(n645bar) );
  OR2_X1 U325 ( .A1(n644), .A2(n643), .ZN(n863) );
  AND2_X1 U325bar ( .A1(n644bar), .A2(n643bar), .ZN(n863bar) );
  OR2_X1 U326 ( .A1(n642), .A2(n641), .ZN(n643) );
  AND2_X1 U326bar ( .A1(n642bar), .A2(n641bar), .ZN(n643bar) );
  OR2_X1 U327 ( .A1(n640), .A2(n639), .ZN(n641) );
  AND2_X1 U327bar ( .A1(n640bar), .A2(n639bar), .ZN(n641bar) );
  OR2_X1 U328 ( .A1(in[127]), .A2(in[122]), .ZN(n639) );
  AND2_X1 U328bar ( .A1(inbar[127]), .A2(inbar[122]), .ZN(n639bar) );
  OR2_X1 U329 ( .A1(in[156]), .A2(in[132]), .ZN(n640) );
  AND2_X1 U329bar ( .A1(inbar[156]), .A2(inbar[132]), .ZN(n640bar) );
  OR2_X1 U330 ( .A1(n638), .A2(n637), .ZN(n642) );
  AND2_X1 U330bar ( .A1(n638bar), .A2(n637bar), .ZN(n642bar) );
  OR2_X1 U331 ( .A1(in[159]), .A2(in[157]), .ZN(n637) );
  AND2_X1 U331bar ( .A1(inbar[159]), .A2(inbar[157]), .ZN(n637bar) );
  OR2_X1 U332 ( .A1(in[185]), .A2(in[169]), .ZN(n638) );
  AND2_X1 U332bar ( .A1(inbar[185]), .A2(inbar[169]), .ZN(n638bar) );
  OR2_X1 U333 ( .A1(n636), .A2(n635), .ZN(n644) );
  AND2_X1 U333bar ( .A1(n636bar), .A2(n635bar), .ZN(n644bar) );
  OR2_X1 U334 ( .A1(n634), .A2(n633), .ZN(n635) );
  AND2_X1 U334bar ( .A1(n634bar), .A2(n633bar), .ZN(n635bar) );
  OR2_X1 U335 ( .A1(in[239]), .A2(in[218]), .ZN(n633) );
  AND2_X1 U335bar ( .A1(inbar[239]), .A2(inbar[218]), .ZN(n633bar) );
  OR2_X1 U336 ( .A1(in_13), .A2(in[87]), .ZN(n634) );
  AND2_X1 U336bar ( .A1(in_13bar), .A2(inbar[87]), .ZN(n634bar) );
  OR2_X1 U337 ( .A1(n632), .A2(n631), .ZN(n636) );
  AND2_X1 U337bar ( .A1(n632bar), .A2(n631bar), .ZN(n636bar) );
  OR2_X1 U338 ( .A1(in_72), .A2(in_70), .ZN(n631) );
  AND2_X1 U338bar ( .A1(in_72bar), .A2(in_70bar), .ZN(n631bar) );
  OR2_X1 U339 ( .A1(in_80), .A2(in_74), .ZN(n632) );
  AND2_X1 U339bar ( .A1(in_80bar), .A2(in_74bar), .ZN(n632bar) );
  OR2_X1 U340 ( .A1(n630), .A2(n629), .ZN(n942) );
  AND2_X1 U340bar ( .A1(n630bar), .A2(n629bar), .ZN(n942bar) );
  OR2_X1 U341 ( .A1(n628), .A2(n627), .ZN(n629) );
  AND2_X1 U341bar ( .A1(n628bar), .A2(n627bar), .ZN(n629bar) );
  OR2_X1 U342 ( .A1(n626), .A2(n625), .ZN(n627) );
  AND2_X1 U342bar ( .A1(n626bar), .A2(n625bar), .ZN(n627bar) );
  OR2_X1 U343 ( .A1(in[146]), .A2(in[100]), .ZN(n625) );
  AND2_X1 U343bar ( .A1(inbar[146]), .A2(inbar[100]), .ZN(n625bar) );
  OR2_X1 U344 ( .A1(in[168]), .A2(in[152]), .ZN(n626) );
  AND2_X1 U344bar ( .A1(inbar[168]), .A2(inbar[152]), .ZN(n626bar) );
  OR2_X1 U345 ( .A1(n624), .A2(n623), .ZN(n628) );
  AND2_X1 U345bar ( .A1(n624bar), .A2(n623bar), .ZN(n628bar) );
  OR2_X1 U346 ( .A1(in[199]), .A2(in[182]), .ZN(n623) );
  AND2_X1 U346bar ( .A1(inbar[199]), .A2(inbar[182]), .ZN(n623bar) );
  OR2_X1 U347 ( .A1(in[236]), .A2(in[204]), .ZN(n624) );
  AND2_X1 U347bar ( .A1(inbar[236]), .A2(inbar[204]), .ZN(n624bar) );
  OR2_X1 U348 ( .A1(n622), .A2(n621), .ZN(n630) );
  AND2_X1 U348bar ( .A1(n622bar), .A2(n621bar), .ZN(n630bar) );
  OR2_X1 U349 ( .A1(n620), .A2(n619), .ZN(n621) );
  AND2_X1 U349bar ( .A1(n620bar), .A2(n619bar), .ZN(n621bar) );
  OR2_X1 U350 ( .A1(in[89]), .A2(in[246]), .ZN(n619) );
  AND2_X1 U350bar ( .A1(inbar[89]), .A2(inbar[246]), .ZN(n619bar) );
  OR2_X1 U351 ( .A1(in[95]), .A2(in[92]), .ZN(n620) );
  AND2_X1 U351bar ( .A1(inbar[95]), .A2(inbar[92]), .ZN(n620bar) );
  OR2_X1 U352 ( .A1(n618), .A2(n617), .ZN(n622) );
  AND2_X1 U352bar ( .A1(n618bar), .A2(n617bar), .ZN(n622bar) );
  OR2_X1 U353 ( .A1(in_22), .A2(in_16), .ZN(n617) );
  AND2_X1 U353bar ( .A1(in_22bar), .A2(in_16bar), .ZN(n617bar) );
  OR2_X1 U354 ( .A1(in_51), .A2(in_49), .ZN(n618) );
  AND2_X1 U354bar ( .A1(in_51bar), .A2(in_49bar), .ZN(n618bar) );
  OR2_X1 U355 ( .A1(n616), .A2(n615), .ZN(n722) );
  AND2_X1 U355bar ( .A1(n616bar), .A2(n615bar), .ZN(n722bar) );
  OR2_X1 U356 ( .A1(in[158]), .A2(in[115]), .ZN(n615) );
  AND2_X1 U356bar ( .A1(inbar[158]), .A2(inbar[115]), .ZN(n615bar) );
  OR2_X1 U357 ( .A1(in[163]), .A2(n614), .ZN(n616) );
  AND2_X1 U357bar ( .A1(inbar[163]), .A2(n614bar), .ZN(n616bar) );
  OR2_X1 U358 ( .A1(in[206]), .A2(in[165]), .ZN(n614) );
  AND2_X1 U358bar ( .A1(inbar[206]), .A2(inbar[165]), .ZN(n614bar) );
  OR2_X1 U359 ( .A1(n613), .A2(n612), .ZN(n724) );
  AND2_X1 U359bar ( .A1(n613bar), .A2(n612bar), .ZN(n724bar) );
  OR2_X1 U360 ( .A1(n611), .A2(n610), .ZN(n612) );
  AND2_X1 U360bar ( .A1(n611bar), .A2(n610bar), .ZN(n612bar) );
  OR2_X1 U361 ( .A1(in[213]), .A2(in[207]), .ZN(n610) );
  AND2_X1 U361bar ( .A1(inbar[213]), .A2(inbar[207]), .ZN(n610bar) );
  OR2_X1 U362 ( .A1(in[215]), .A2(n609), .ZN(n611) );
  AND2_X1 U362bar ( .A1(inbar[215]), .A2(n609bar), .ZN(n611bar) );
  OR2_X1 U363 ( .A1(in[230]), .A2(in[220]), .ZN(n609) );
  AND2_X1 U363bar ( .A1(inbar[230]), .A2(inbar[220]), .ZN(n609bar) );
  OR2_X1 U364 ( .A1(n608), .A2(n607), .ZN(n613) );
  AND2_X1 U364bar ( .A1(n608bar), .A2(n607bar), .ZN(n613bar) );
  OR2_X1 U365 ( .A1(in[251]), .A2(in[234]), .ZN(n607) );
  AND2_X1 U365bar ( .A1(inbar[251]), .A2(inbar[234]), .ZN(n607bar) );
  OR2_X1 U366 ( .A1(in_17), .A2(n606), .ZN(n608) );
  AND2_X1 U366bar ( .A1(in_17bar), .A2(n606bar), .ZN(n608bar) );
  OR2_X1 U367 ( .A1(in_65), .A2(in_56), .ZN(n606) );
  AND2_X1 U367bar ( .A1(in_65bar), .A2(in_56bar), .ZN(n606bar) );
  OR2_X1 U368 ( .A1(n605), .A2(n604), .ZN(out[0]) );
  AND2_X1 U368bar ( .A1(n605bar), .A2(n604bar), .ZN(outbar[0]) );
  OR2_X1 U369 ( .A1(n603), .A2(n602), .ZN(n604) );
  AND2_X1 U369bar ( .A1(n603bar), .A2(n602bar), .ZN(n604bar) );
  OR2_X1 U370 ( .A1(n601), .A2(n600), .ZN(n602) );
  AND2_X1 U370bar ( .A1(n601bar), .A2(n600bar), .ZN(n602bar) );
  OR2_X1 U371 ( .A1(n820), .A2(n785), .ZN(n600) );
  AND2_X1 U371bar ( .A1(n820bar), .A2(n785bar), .ZN(n600bar) );
  OR2_X1 U372 ( .A1(n599), .A2(n598), .ZN(n785) );
  AND2_X1 U372bar ( .A1(n599bar), .A2(n598bar), .ZN(n785bar) );
  OR2_X1 U373 ( .A1(n597), .A2(n596), .ZN(n598) );
  AND2_X1 U373bar ( .A1(n597bar), .A2(n596bar), .ZN(n598bar) );
  OR2_X1 U374 ( .A1(n595), .A2(n594), .ZN(n596) );
  AND2_X1 U374bar ( .A1(n595bar), .A2(n594bar), .ZN(n596bar) );
  OR2_X1 U375 ( .A1(in[135]), .A2(in[104]), .ZN(n594) );
  AND2_X1 U375bar ( .A1(inbar[135]), .A2(inbar[104]), .ZN(n594bar) );
  OR2_X1 U376 ( .A1(in[188]), .A2(in[178]), .ZN(n595) );
  AND2_X1 U376bar ( .A1(inbar[188]), .A2(inbar[178]), .ZN(n595bar) );
  OR2_X1 U377 ( .A1(n593), .A2(n592), .ZN(n597) );
  AND2_X1 U377bar ( .A1(n593bar), .A2(n592bar), .ZN(n597bar) );
  OR2_X1 U378 ( .A1(in[217]), .A2(in[194]), .ZN(n592) );
  AND2_X1 U378bar ( .A1(inbar[217]), .A2(inbar[194]), .ZN(n592bar) );
  OR2_X1 U379 ( .A1(in[237]), .A2(in[218]), .ZN(n593) );
  AND2_X1 U379bar ( .A1(inbar[237]), .A2(inbar[218]), .ZN(n593bar) );
  OR2_X1 U380 ( .A1(n591), .A2(n590), .ZN(n599) );
  AND2_X1 U380bar ( .A1(n591bar), .A2(n590bar), .ZN(n599bar) );
  OR2_X1 U381 ( .A1(n589), .A2(n588), .ZN(n590) );
  AND2_X1 U381bar ( .A1(n589bar), .A2(n588bar), .ZN(n590bar) );
  OR2_X1 U382 ( .A1(in_2), .A2(in_10), .ZN(n588) );
  AND2_X1 U382bar ( .A1(in_2bar), .A2(in_10bar), .ZN(n588bar) );
  OR2_X1 U383 ( .A1(in_47), .A2(in_22), .ZN(n589) );
  AND2_X1 U383bar ( .A1(in_47bar), .A2(in_22bar), .ZN(n589bar) );
  OR2_X1 U384 ( .A1(n587), .A2(n586), .ZN(n591) );
  AND2_X1 U384bar ( .A1(n587bar), .A2(n586bar), .ZN(n591bar) );
  OR2_X1 U385 ( .A1(in_56), .A2(in_54), .ZN(n586) );
  AND2_X1 U385bar ( .A1(in_56bar), .A2(in_54bar), .ZN(n586bar) );
  OR2_X1 U386 ( .A1(in_63), .A2(in_61), .ZN(n587) );
  AND2_X1 U386bar ( .A1(in_63bar), .A2(in_61bar), .ZN(n587bar) );
  OR2_X1 U387 ( .A1(n585), .A2(n584), .ZN(n820) );
  AND2_X1 U387bar ( .A1(n585bar), .A2(n584bar), .ZN(n820bar) );
  OR2_X1 U388 ( .A1(n583), .A2(n582), .ZN(n584) );
  AND2_X1 U388bar ( .A1(n583bar), .A2(n582bar), .ZN(n584bar) );
  OR2_X1 U389 ( .A1(n581), .A2(n580), .ZN(n582) );
  AND2_X1 U389bar ( .A1(n581bar), .A2(n580bar), .ZN(n582bar) );
  OR2_X1 U390 ( .A1(in[158]), .A2(in[142]), .ZN(n580) );
  AND2_X1 U390bar ( .A1(inbar[158]), .A2(inbar[142]), .ZN(n580bar) );
  OR2_X1 U391 ( .A1(in[175]), .A2(in[164]), .ZN(n581) );
  AND2_X1 U391bar ( .A1(inbar[175]), .A2(inbar[164]), .ZN(n581bar) );
  OR2_X1 U392 ( .A1(n579), .A2(n578), .ZN(n583) );
  AND2_X1 U392bar ( .A1(n579bar), .A2(n578bar), .ZN(n583bar) );
  OR2_X1 U393 ( .A1(in[228]), .A2(in[204]), .ZN(n578) );
  AND2_X1 U393bar ( .A1(inbar[228]), .A2(inbar[204]), .ZN(n578bar) );
  OR2_X1 U394 ( .A1(in[91]), .A2(in[87]), .ZN(n579) );
  AND2_X1 U394bar ( .A1(inbar[91]), .A2(inbar[87]), .ZN(n579bar) );
  OR2_X1 U395 ( .A1(n577), .A2(n576), .ZN(n585) );
  AND2_X1 U395bar ( .A1(n577bar), .A2(n576bar), .ZN(n585bar) );
  OR2_X1 U396 ( .A1(n575), .A2(n574), .ZN(n576) );
  AND2_X1 U396bar ( .A1(n575bar), .A2(n574bar), .ZN(n576bar) );
  OR2_X1 U397 ( .A1(in_21), .A2(in_11), .ZN(n574) );
  AND2_X1 U397bar ( .A1(in_21bar), .A2(in_11bar), .ZN(n574bar) );
  OR2_X1 U398 ( .A1(in_5), .A2(in_3), .ZN(n575) );
  AND2_X1 U398bar ( .A1(in_5bar), .A2(in_3bar), .ZN(n575bar) );
  OR2_X1 U399 ( .A1(n573), .A2(n572), .ZN(n577) );
  AND2_X1 U399bar ( .A1(n573bar), .A2(n572bar), .ZN(n577bar) );
  OR2_X1 U400 ( .A1(in_68), .A2(in_64), .ZN(n572) );
  AND2_X1 U400bar ( .A1(in_68bar), .A2(in_64bar), .ZN(n572bar) );
  OR2_X1 U401 ( .A1(in_76), .A2(in_73), .ZN(n573) );
  AND2_X1 U401bar ( .A1(in_76bar), .A2(in_73bar), .ZN(n573bar) );
  OR2_X1 U402 ( .A1(n778), .A2(n571), .ZN(n601) );
  AND2_X1 U402bar ( .A1(n778bar), .A2(n571bar), .ZN(n601bar) );
  OR2_X1 U403 ( .A1(in[100]), .A2(n965), .ZN(n571) );
  AND2_X1 U403bar ( .A1(inbar[100]), .A2(n965bar), .ZN(n571bar) );
  OR2_X1 U404 ( .A1(n570), .A2(n569), .ZN(n965) );
  AND2_X1 U404bar ( .A1(n570bar), .A2(n569bar), .ZN(n965bar) );
  OR2_X1 U405 ( .A1(n568), .A2(n567), .ZN(n569) );
  AND2_X1 U405bar ( .A1(n568bar), .A2(n567bar), .ZN(n569bar) );
  OR2_X1 U406 ( .A1(n566), .A2(n565), .ZN(n567) );
  AND2_X1 U406bar ( .A1(n566bar), .A2(n565bar), .ZN(n567bar) );
  OR2_X1 U407 ( .A1(n817), .A2(n750), .ZN(n565) );
  AND2_X1 U407bar ( .A1(n817bar), .A2(n750bar), .ZN(n565bar) );
  OR2_X1 U408 ( .A1(n564), .A2(n563), .ZN(n750) );
  AND2_X1 U408bar ( .A1(n564bar), .A2(n563bar), .ZN(n750bar) );
  OR2_X1 U409 ( .A1(n562), .A2(n561), .ZN(n563) );
  AND2_X1 U409bar ( .A1(n562bar), .A2(n561bar), .ZN(n563bar) );
  OR2_X1 U410 ( .A1(n560), .A2(n559), .ZN(n561) );
  AND2_X1 U410bar ( .A1(n560bar), .A2(n559bar), .ZN(n561bar) );
  OR2_X1 U411 ( .A1(in[119]), .A2(in[103]), .ZN(n559) );
  AND2_X1 U411bar ( .A1(inbar[119]), .A2(inbar[103]), .ZN(n559bar) );
  OR2_X1 U412 ( .A1(in[137]), .A2(in[133]), .ZN(n560) );
  AND2_X1 U412bar ( .A1(inbar[137]), .A2(inbar[133]), .ZN(n560bar) );
  OR2_X1 U413 ( .A1(n558), .A2(n557), .ZN(n562) );
  AND2_X1 U413bar ( .A1(n558bar), .A2(n557bar), .ZN(n562bar) );
  OR2_X1 U414 ( .A1(in[176]), .A2(in[173]), .ZN(n557) );
  AND2_X1 U414bar ( .A1(inbar[176]), .A2(inbar[173]), .ZN(n557bar) );
  OR2_X1 U415 ( .A1(in[210]), .A2(in[181]), .ZN(n558) );
  AND2_X1 U415bar ( .A1(inbar[210]), .A2(inbar[181]), .ZN(n558bar) );
  OR2_X1 U416 ( .A1(n556), .A2(n555), .ZN(n564) );
  AND2_X1 U416bar ( .A1(n556bar), .A2(n555bar), .ZN(n564bar) );
  OR2_X1 U417 ( .A1(n554), .A2(n553), .ZN(n555) );
  AND2_X1 U417bar ( .A1(n554bar), .A2(n553bar), .ZN(n555bar) );
  OR2_X1 U418 ( .A1(in_13), .A2(in[234]), .ZN(n553) );
  AND2_X1 U418bar ( .A1(in_13bar), .A2(inbar[234]), .ZN(n553bar) );
  OR2_X1 U419 ( .A1(in_38), .A2(in_32), .ZN(n554) );
  AND2_X1 U419bar ( .A1(in_38bar), .A2(in_32bar), .ZN(n554bar) );
  OR2_X1 U420 ( .A1(n552), .A2(n551), .ZN(n556) );
  AND2_X1 U420bar ( .A1(n552bar), .A2(n551bar), .ZN(n556bar) );
  OR2_X1 U421 ( .A1(in_42), .A2(in_41), .ZN(n551) );
  AND2_X1 U421bar ( .A1(in_42bar), .A2(in_41bar), .ZN(n551bar) );
  OR2_X1 U422 ( .A1(in_7), .A2(in_49), .ZN(n552) );
  AND2_X1 U422bar ( .A1(in_7bar), .A2(in_49bar), .ZN(n552bar) );
  OR2_X1 U423 ( .A1(n550), .A2(n549), .ZN(n817) );
  AND2_X1 U423bar ( .A1(n550bar), .A2(n549bar), .ZN(n817bar) );
  OR2_X1 U424 ( .A1(n548), .A2(n547), .ZN(n549) );
  AND2_X1 U424bar ( .A1(n548bar), .A2(n547bar), .ZN(n549bar) );
  OR2_X1 U425 ( .A1(n546), .A2(n545), .ZN(n547) );
  AND2_X1 U425bar ( .A1(n546bar), .A2(n545bar), .ZN(n547bar) );
  OR2_X1 U426 ( .A1(in[159]), .A2(in[105]), .ZN(n545) );
  AND2_X1 U426bar ( .A1(inbar[159]), .A2(inbar[105]), .ZN(n545bar) );
  OR2_X1 U427 ( .A1(in[206]), .A2(in[183]), .ZN(n546) );
  AND2_X1 U427bar ( .A1(inbar[206]), .A2(inbar[183]), .ZN(n546bar) );
  OR2_X1 U428 ( .A1(n544), .A2(n543), .ZN(n548) );
  AND2_X1 U428bar ( .A1(n544bar), .A2(n543bar), .ZN(n548bar) );
  OR2_X1 U429 ( .A1(in[229]), .A2(in[219]), .ZN(n543) );
  AND2_X1 U429bar ( .A1(inbar[229]), .A2(inbar[219]), .ZN(n543bar) );
  OR2_X1 U430 ( .A1(in[235]), .A2(in[232]), .ZN(n544) );
  AND2_X1 U430bar ( .A1(inbar[235]), .A2(inbar[232]), .ZN(n544bar) );
  OR2_X1 U431 ( .A1(n542), .A2(n541), .ZN(n550) );
  AND2_X1 U431bar ( .A1(n542bar), .A2(n541bar), .ZN(n550bar) );
  OR2_X1 U432 ( .A1(n540), .A2(n539), .ZN(n541) );
  AND2_X1 U432bar ( .A1(n540bar), .A2(n539bar), .ZN(n541bar) );
  OR2_X1 U433 ( .A1(in[249]), .A2(in[242]), .ZN(n539) );
  AND2_X1 U433bar ( .A1(inbar[249]), .A2(inbar[242]), .ZN(n539bar) );
  OR2_X1 U434 ( .A1(in[89]), .A2(in[254]), .ZN(n540) );
  AND2_X1 U434bar ( .A1(inbar[89]), .A2(inbar[254]), .ZN(n540bar) );
  OR2_X1 U435 ( .A1(n538), .A2(n537), .ZN(n542) );
  AND2_X1 U435bar ( .A1(n538bar), .A2(n537bar), .ZN(n542bar) );
  OR2_X1 U436 ( .A1(in_14), .A2(in[99]), .ZN(n537) );
  AND2_X1 U436bar ( .A1(in_14bar), .A2(inbar[99]), .ZN(n537bar) );
  OR2_X1 U437 ( .A1(in_60), .A2(in_18), .ZN(n538) );
  AND2_X1 U437bar ( .A1(in_60bar), .A2(in_18bar), .ZN(n538bar) );
  OR2_X1 U438 ( .A1(in[113]), .A2(n763), .ZN(n566) );
  AND2_X1 U438bar ( .A1(inbar[113]), .A2(n763bar), .ZN(n566bar) );
  OR2_X1 U439 ( .A1(n536), .A2(n535), .ZN(n763) );
  AND2_X1 U439bar ( .A1(n536bar), .A2(n535bar), .ZN(n763bar) );
  OR2_X1 U440 ( .A1(n534), .A2(n533), .ZN(n535) );
  AND2_X1 U440bar ( .A1(n534bar), .A2(n533bar), .ZN(n535bar) );
  OR2_X1 U441 ( .A1(n532), .A2(n531), .ZN(n533) );
  AND2_X1 U441bar ( .A1(n532bar), .A2(n531bar), .ZN(n533bar) );
  OR2_X1 U442 ( .A1(in[115]), .A2(in[110]), .ZN(n531) );
  AND2_X1 U442bar ( .A1(inbar[115]), .A2(inbar[110]), .ZN(n531bar) );
  OR2_X1 U443 ( .A1(in[125]), .A2(in[117]), .ZN(n532) );
  AND2_X1 U443bar ( .A1(inbar[125]), .A2(inbar[117]), .ZN(n532bar) );
  OR2_X1 U444 ( .A1(n530), .A2(n529), .ZN(n534) );
  AND2_X1 U444bar ( .A1(n530bar), .A2(n529bar), .ZN(n534bar) );
  OR2_X1 U445 ( .A1(in[180]), .A2(in[128]), .ZN(n529) );
  AND2_X1 U445bar ( .A1(inbar[180]), .A2(inbar[128]), .ZN(n529bar) );
  OR2_X1 U446 ( .A1(in[205]), .A2(in[201]), .ZN(n530) );
  AND2_X1 U446bar ( .A1(inbar[205]), .A2(inbar[201]), .ZN(n530bar) );
  OR2_X1 U447 ( .A1(n528), .A2(n527), .ZN(n536) );
  AND2_X1 U447bar ( .A1(n528bar), .A2(n527bar), .ZN(n536bar) );
  OR2_X1 U448 ( .A1(n526), .A2(n525), .ZN(n527) );
  AND2_X1 U448bar ( .A1(n526bar), .A2(n525bar), .ZN(n527bar) );
  OR2_X1 U449 ( .A1(in[244]), .A2(in[239]), .ZN(n525) );
  AND2_X1 U449bar ( .A1(inbar[244]), .A2(inbar[239]), .ZN(n525bar) );
  OR2_X1 U450 ( .A1(in[95]), .A2(in[83]), .ZN(n526) );
  AND2_X1 U450bar ( .A1(inbar[95]), .A2(inbar[83]), .ZN(n526bar) );
  OR2_X1 U451 ( .A1(n524), .A2(n523), .ZN(n528) );
  AND2_X1 U451bar ( .A1(n524bar), .A2(n523bar), .ZN(n528bar) );
  OR2_X1 U452 ( .A1(in_24), .A2(in[97]), .ZN(n523) );
  AND2_X1 U452bar ( .A1(in_24bar), .A2(inbar[97]), .ZN(n523bar) );
  OR2_X1 U453 ( .A1(in_33), .A2(in_27), .ZN(n524) );
  AND2_X1 U453bar ( .A1(in_33bar), .A2(in_27bar), .ZN(n524bar) );
  OR2_X1 U454 ( .A1(n522), .A2(n521), .ZN(n568) );
  AND2_X1 U454bar ( .A1(n522bar), .A2(n521bar), .ZN(n568bar) );
  OR2_X1 U455 ( .A1(in[145]), .A2(in[126]), .ZN(n521) );
  AND2_X1 U455bar ( .A1(inbar[145]), .A2(inbar[126]), .ZN(n521bar) );
  OR2_X1 U456 ( .A1(in[169]), .A2(n520), .ZN(n522) );
  AND2_X1 U456bar ( .A1(inbar[169]), .A2(n520bar), .ZN(n522bar) );
  OR2_X1 U457 ( .A1(in[221]), .A2(in[172]), .ZN(n520) );
  AND2_X1 U457bar ( .A1(inbar[221]), .A2(inbar[172]), .ZN(n520bar) );
  OR2_X1 U458 ( .A1(n519), .A2(n518), .ZN(n570) );
  AND2_X1 U458bar ( .A1(n519bar), .A2(n518bar), .ZN(n570bar) );
  OR2_X1 U459 ( .A1(n517), .A2(n516), .ZN(n518) );
  AND2_X1 U459bar ( .A1(n517bar), .A2(n516bar), .ZN(n518bar) );
  OR2_X1 U460 ( .A1(in[241]), .A2(in[224]), .ZN(n516) );
  AND2_X1 U460bar ( .A1(inbar[241]), .A2(inbar[224]), .ZN(n516bar) );
  OR2_X1 U461 ( .A1(in[86]), .A2(n515), .ZN(n517) );
  AND2_X1 U461bar ( .A1(inbar[86]), .A2(n515bar), .ZN(n517bar) );
  OR2_X1 U462 ( .A1(in_43), .A2(in_34), .ZN(n515) );
  AND2_X1 U462bar ( .A1(in_43bar), .A2(in_34bar), .ZN(n515bar) );
  OR2_X1 U463 ( .A1(n514), .A2(n513), .ZN(n519) );
  AND2_X1 U463bar ( .A1(n514bar), .A2(n513bar), .ZN(n519bar) );
  OR2_X1 U464 ( .A1(in_65), .A2(in_51), .ZN(n513) );
  AND2_X1 U464bar ( .A1(in_65bar), .A2(in_51bar), .ZN(n513bar) );
  OR2_X1 U465 ( .A1(in_75), .A2(n512), .ZN(n514) );
  AND2_X1 U465bar ( .A1(in_75bar), .A2(n512bar), .ZN(n514bar) );
  OR2_X1 U466 ( .A1(in_81), .A2(in_77), .ZN(n512) );
  AND2_X1 U466bar ( .A1(in_81bar), .A2(in_77bar), .ZN(n512bar) );
  OR2_X1 U467 ( .A1(n511), .A2(n510), .ZN(n778) );
  AND2_X1 U467bar ( .A1(n511bar), .A2(n510bar), .ZN(n778bar) );
  OR2_X1 U468 ( .A1(n509), .A2(n508), .ZN(n510) );
  AND2_X1 U468bar ( .A1(n509bar), .A2(n508bar), .ZN(n510bar) );
  OR2_X1 U469 ( .A1(n507), .A2(n506), .ZN(n508) );
  AND2_X1 U469bar ( .A1(n507bar), .A2(n506bar), .ZN(n508bar) );
  OR2_X1 U470 ( .A1(in[107]), .A2(in[101]), .ZN(n506) );
  AND2_X1 U470bar ( .A1(inbar[107]), .A2(inbar[101]), .ZN(n506bar) );
  OR2_X1 U471 ( .A1(in[139]), .A2(in[132]), .ZN(n507) );
  AND2_X1 U471bar ( .A1(inbar[139]), .A2(inbar[132]), .ZN(n507bar) );
  OR2_X1 U472 ( .A1(n505), .A2(n504), .ZN(n509) );
  AND2_X1 U472bar ( .A1(n505bar), .A2(n504bar), .ZN(n509bar) );
  OR2_X1 U473 ( .A1(in[146]), .A2(in[141]), .ZN(n504) );
  AND2_X1 U473bar ( .A1(inbar[146]), .A2(inbar[141]), .ZN(n504bar) );
  OR2_X1 U474 ( .A1(in[203]), .A2(in[179]), .ZN(n505) );
  AND2_X1 U474bar ( .A1(inbar[203]), .A2(inbar[179]), .ZN(n505bar) );
  OR2_X1 U475 ( .A1(n503), .A2(n502), .ZN(n511) );
  AND2_X1 U475bar ( .A1(n503bar), .A2(n502bar), .ZN(n511bar) );
  OR2_X1 U476 ( .A1(n501), .A2(n500), .ZN(n502) );
  AND2_X1 U476bar ( .A1(n501bar), .A2(n500bar), .ZN(n502bar) );
  OR2_X1 U477 ( .A1(in[243]), .A2(in[222]), .ZN(n500) );
  AND2_X1 U477bar ( .A1(inbar[243]), .A2(inbar[222]), .ZN(n500bar) );
  OR2_X1 U478 ( .A1(in[251]), .A2(in[250]), .ZN(n501) );
  AND2_X1 U478bar ( .A1(inbar[251]), .A2(inbar[250]), .ZN(n501bar) );
  OR2_X1 U479 ( .A1(n499), .A2(n498), .ZN(n503) );
  AND2_X1 U479bar ( .A1(n499bar), .A2(n498bar), .ZN(n503bar) );
  OR2_X1 U480 ( .A1(in_37), .A2(in_19), .ZN(n498) );
  AND2_X1 U480bar ( .A1(in_37bar), .A2(in_19bar), .ZN(n498bar) );
  OR2_X1 U481 ( .A1(in_78), .A2(in_6), .ZN(n499) );
  AND2_X1 U481bar ( .A1(in_78bar), .A2(in_6bar), .ZN(n499bar) );
  OR2_X1 U482 ( .A1(n497), .A2(n496), .ZN(n603) );
  AND2_X1 U482bar ( .A1(n497bar), .A2(n496bar), .ZN(n603bar) );
  OR2_X1 U483 ( .A1(in[112]), .A2(in[102]), .ZN(n496) );
  AND2_X1 U483bar ( .A1(inbar[112]), .A2(inbar[102]), .ZN(n496bar) );
  OR2_X1 U484 ( .A1(in[123]), .A2(n495), .ZN(n497) );
  AND2_X1 U484bar ( .A1(inbar[123]), .A2(n495bar), .ZN(n497bar) );
  OR2_X1 U485 ( .A1(in[143]), .A2(in[130]), .ZN(n495) );
  AND2_X1 U485bar ( .A1(inbar[143]), .A2(inbar[130]), .ZN(n495bar) );
  OR2_X1 U486 ( .A1(n494), .A2(n493), .ZN(n605) );
  AND2_X1 U486bar ( .A1(n494bar), .A2(n493bar), .ZN(n605bar) );
  OR2_X1 U487 ( .A1(n492), .A2(n491), .ZN(n493) );
  AND2_X1 U487bar ( .A1(n492bar), .A2(n491bar), .ZN(n493bar) );
  OR2_X1 U488 ( .A1(in[216]), .A2(in[213]), .ZN(n491) );
  AND2_X1 U488bar ( .A1(inbar[216]), .A2(inbar[213]), .ZN(n491bar) );
  OR2_X1 U489 ( .A1(in[227]), .A2(n490), .ZN(n492) );
  AND2_X1 U489bar ( .A1(inbar[227]), .A2(n490bar), .ZN(n492bar) );
  OR2_X1 U490 ( .A1(in_0), .A2(in[248]), .ZN(n490) );
  AND2_X1 U490bar ( .A1(in_0bar), .A2(inbar[248]), .ZN(n490bar) );
  OR2_X1 U491 ( .A1(n489), .A2(n488), .ZN(n494) );
  AND2_X1 U491bar ( .A1(n489bar), .A2(n488bar), .ZN(n494bar) );
  OR2_X1 U492 ( .A1(in_46), .A2(in_44), .ZN(n488) );
  AND2_X1 U492bar ( .A1(in_46bar), .A2(in_44bar), .ZN(n488bar) );
  OR2_X1 U493 ( .A1(in_50), .A2(n487), .ZN(n489) );
  AND2_X1 U493bar ( .A1(in_50bar), .A2(n487bar), .ZN(n489bar) );
  OR2_X1 U494 ( .A1(in_9), .A2(in_80), .ZN(n487) );
  AND2_X1 U494bar ( .A1(in_9bar), .A2(in_80bar), .ZN(n487bar) );
endmodule

module sBox_0 ( in, inbar, out, outbar );

  input wire [7:0] in;
  input wire [7:0] inbar;
//input_done

  output wire [7:0] out;
  output wire [7:0] outbar;
//output_done

  wire [255:0] decodeOut;
  wire [255:0] decodeOutbar;
//wire_done

  decode_0 dec ( .in(in), .inbar(inbar), .out(decodeOut), .outbar(decodeOutbar) );
  encode_0 enc ( .in(decodeOut), .inbar(decodeOutbar), .out(out), .outbar(outbar) );
endmodule

module CD2_1 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD2_2 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD2_3 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD2_4 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD4_1 ( a, abar, b, bbar, y, ybar );

  input wire [3:0] a;
  input wire [3:0] b;
  input wire [3:0] abar;
  input wire [3:0] bbar;
//input_done

  output wire [15:0] y;
  output wire [15:0] ybar;
//output_done

//wire_done

  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]) );
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]) );
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]) );
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]) );
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]) );
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]) );
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]) );
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]) );
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]) );
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]) );
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]) );
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]) );
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]) );
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]) );
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]) );
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]) );
endmodule

module CD4_2 ( a, abar, b, bbar, y, ybar );

  input wire [3:0] a;
  input wire [3:0] b;
  input wire [3:0] abar;
  input wire [3:0] bbar;
//input_done

  output wire [15:0] y;
  output wire [15:0] ybar;
//output_done

//wire_done

  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]) );
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]) );
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]) );
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]) );
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]) );
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]) );
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]) );
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]) );
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]) );
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]) );
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]) );
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]) );
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]) );
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]) );
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]) );
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]) );
endmodule

module CD16_1 ( a, abar, b, bbar, y, ybar );

  input wire [15:0] a;
  input wire [15:0] b;
  input wire [15:0] abar;
  input wire [15:0] bbar;
//input_done

  output wire [255:0] y;
  output wire [255:0] ybar;
//output_done

//wire_done

  AND2_X1 U1 ( .A1(b[9]), .A2(a[0]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[9]), .A2(abar[0]), .ZN(ybar[9]) );
  AND2_X1 U2 ( .A1(b[3]), .A2(a[6]), .ZN(y[99]) );
  OR2_X1 U2bar ( .A1(bbar[3]), .A2(abar[6]), .ZN(ybar[99]) );
  AND2_X1 U3 ( .A1(b[2]), .A2(a[6]), .ZN(y[98]) );
  OR2_X1 U3bar ( .A1(bbar[2]), .A2(abar[6]), .ZN(ybar[98]) );
  AND2_X1 U4 ( .A1(b[1]), .A2(a[6]), .ZN(y[97]) );
  OR2_X1 U4bar ( .A1(bbar[1]), .A2(abar[6]), .ZN(ybar[97]) );
  AND2_X1 U5 ( .A1(b[0]), .A2(a[6]), .ZN(y[96]) );
  OR2_X1 U5bar ( .A1(bbar[0]), .A2(abar[6]), .ZN(ybar[96]) );
  AND2_X1 U6 ( .A1(b[15]), .A2(a[5]), .ZN(y[95]) );
  OR2_X1 U6bar ( .A1(bbar[15]), .A2(abar[5]), .ZN(ybar[95]) );
  AND2_X1 U7 ( .A1(b[14]), .A2(a[5]), .ZN(y[94]) );
  OR2_X1 U7bar ( .A1(bbar[14]), .A2(abar[5]), .ZN(ybar[94]) );
  AND2_X1 U8 ( .A1(b[13]), .A2(a[5]), .ZN(y[93]) );
  OR2_X1 U8bar ( .A1(bbar[13]), .A2(abar[5]), .ZN(ybar[93]) );
  AND2_X1 U9 ( .A1(b[12]), .A2(a[5]), .ZN(y[92]) );
  OR2_X1 U9bar ( .A1(bbar[12]), .A2(abar[5]), .ZN(ybar[92]) );
  AND2_X1 U10 ( .A1(b[11]), .A2(a[5]), .ZN(y[91]) );
  OR2_X1 U10bar ( .A1(bbar[11]), .A2(abar[5]), .ZN(ybar[91]) );
  AND2_X1 U11 ( .A1(b[10]), .A2(a[5]), .ZN(y[90]) );
  OR2_X1 U11bar ( .A1(bbar[10]), .A2(abar[5]), .ZN(ybar[90]) );
  AND2_X1 U12 ( .A1(b[8]), .A2(a[0]), .ZN(y[8]) );
  OR2_X1 U12bar ( .A1(bbar[8]), .A2(abar[0]), .ZN(ybar[8]) );
  AND2_X1 U13 ( .A1(a[5]), .A2(b[9]), .ZN(y[89]) );
  OR2_X1 U13bar ( .A1(abar[5]), .A2(bbar[9]), .ZN(ybar[89]) );
  AND2_X1 U14 ( .A1(b[8]), .A2(a[5]), .ZN(y[88]) );
  OR2_X1 U14bar ( .A1(bbar[8]), .A2(abar[5]), .ZN(ybar[88]) );
  AND2_X1 U15 ( .A1(b[7]), .A2(a[5]), .ZN(y[87]) );
  OR2_X1 U15bar ( .A1(bbar[7]), .A2(abar[5]), .ZN(ybar[87]) );
  AND2_X1 U16 ( .A1(b[6]), .A2(a[5]), .ZN(y[86]) );
  OR2_X1 U16bar ( .A1(bbar[6]), .A2(abar[5]), .ZN(ybar[86]) );
  AND2_X1 U17 ( .A1(b[5]), .A2(a[5]), .ZN(y[85]) );
  OR2_X1 U17bar ( .A1(bbar[5]), .A2(abar[5]), .ZN(ybar[85]) );
  AND2_X1 U18 ( .A1(b[4]), .A2(a[5]), .ZN(y[84]) );
  OR2_X1 U18bar ( .A1(bbar[4]), .A2(abar[5]), .ZN(ybar[84]) );
  AND2_X1 U19 ( .A1(a[5]), .A2(b[3]), .ZN(y[83]) );
  OR2_X1 U19bar ( .A1(abar[5]), .A2(bbar[3]), .ZN(ybar[83]) );
  AND2_X1 U20 ( .A1(a[5]), .A2(b[2]), .ZN(y[82]) );
  OR2_X1 U20bar ( .A1(abar[5]), .A2(bbar[2]), .ZN(ybar[82]) );
  AND2_X1 U21 ( .A1(a[5]), .A2(b[1]), .ZN(y[81]) );
  OR2_X1 U21bar ( .A1(abar[5]), .A2(bbar[1]), .ZN(ybar[81]) );
  AND2_X1 U22 ( .A1(a[5]), .A2(b[0]), .ZN(y[80]) );
  OR2_X1 U22bar ( .A1(abar[5]), .A2(bbar[0]), .ZN(ybar[80]) );
  AND2_X1 U23 ( .A1(b[7]), .A2(a[0]), .ZN(y[7]) );
  OR2_X1 U23bar ( .A1(bbar[7]), .A2(abar[0]), .ZN(ybar[7]) );
  AND2_X1 U24 ( .A1(a[4]), .A2(b[15]), .ZN(y[79]) );
  OR2_X1 U24bar ( .A1(abar[4]), .A2(bbar[15]), .ZN(ybar[79]) );
  AND2_X1 U25 ( .A1(a[4]), .A2(b[14]), .ZN(y[78]) );
  OR2_X1 U25bar ( .A1(abar[4]), .A2(bbar[14]), .ZN(ybar[78]) );
  AND2_X1 U26 ( .A1(a[4]), .A2(b[13]), .ZN(y[77]) );
  OR2_X1 U26bar ( .A1(abar[4]), .A2(bbar[13]), .ZN(ybar[77]) );
  AND2_X1 U27 ( .A1(a[4]), .A2(b[12]), .ZN(y[76]) );
  OR2_X1 U27bar ( .A1(abar[4]), .A2(bbar[12]), .ZN(ybar[76]) );
  AND2_X1 U28 ( .A1(a[4]), .A2(b[11]), .ZN(y[75]) );
  OR2_X1 U28bar ( .A1(abar[4]), .A2(bbar[11]), .ZN(ybar[75]) );
  AND2_X1 U29 ( .A1(a[4]), .A2(b[10]), .ZN(y[74]) );
  OR2_X1 U29bar ( .A1(abar[4]), .A2(bbar[10]), .ZN(ybar[74]) );
  AND2_X1 U30 ( .A1(a[4]), .A2(b[9]), .ZN(y[73]) );
  OR2_X1 U30bar ( .A1(abar[4]), .A2(bbar[9]), .ZN(ybar[73]) );
  AND2_X1 U31 ( .A1(a[4]), .A2(b[8]), .ZN(y[72]) );
  OR2_X1 U31bar ( .A1(abar[4]), .A2(bbar[8]), .ZN(ybar[72]) );
  AND2_X1 U32 ( .A1(a[4]), .A2(b[7]), .ZN(y[71]) );
  OR2_X1 U32bar ( .A1(abar[4]), .A2(bbar[7]), .ZN(ybar[71]) );
  AND2_X1 U33 ( .A1(a[4]), .A2(b[6]), .ZN(y[70]) );
  OR2_X1 U33bar ( .A1(abar[4]), .A2(bbar[6]), .ZN(ybar[70]) );
  AND2_X1 U34 ( .A1(b[6]), .A2(a[0]), .ZN(y[6]) );
  OR2_X1 U34bar ( .A1(bbar[6]), .A2(abar[0]), .ZN(ybar[6]) );
  AND2_X1 U35 ( .A1(a[4]), .A2(b[5]), .ZN(y[69]) );
  OR2_X1 U35bar ( .A1(abar[4]), .A2(bbar[5]), .ZN(ybar[69]) );
  AND2_X1 U36 ( .A1(a[4]), .A2(b[4]), .ZN(y[68]) );
  OR2_X1 U36bar ( .A1(abar[4]), .A2(bbar[4]), .ZN(ybar[68]) );
  AND2_X1 U37 ( .A1(a[4]), .A2(b[3]), .ZN(y[67]) );
  OR2_X1 U37bar ( .A1(abar[4]), .A2(bbar[3]), .ZN(ybar[67]) );
  AND2_X1 U38 ( .A1(a[4]), .A2(b[2]), .ZN(y[66]) );
  OR2_X1 U38bar ( .A1(abar[4]), .A2(bbar[2]), .ZN(ybar[66]) );
  AND2_X1 U39 ( .A1(a[4]), .A2(b[1]), .ZN(y[65]) );
  OR2_X1 U39bar ( .A1(abar[4]), .A2(bbar[1]), .ZN(ybar[65]) );
  AND2_X1 U40 ( .A1(a[4]), .A2(b[0]), .ZN(y[64]) );
  OR2_X1 U40bar ( .A1(abar[4]), .A2(bbar[0]), .ZN(ybar[64]) );
  AND2_X1 U41 ( .A1(a[3]), .A2(b[15]), .ZN(y[63]) );
  OR2_X1 U41bar ( .A1(abar[3]), .A2(bbar[15]), .ZN(ybar[63]) );
  AND2_X1 U42 ( .A1(a[3]), .A2(b[14]), .ZN(y[62]) );
  OR2_X1 U42bar ( .A1(abar[3]), .A2(bbar[14]), .ZN(ybar[62]) );
  AND2_X1 U43 ( .A1(a[3]), .A2(b[13]), .ZN(y[61]) );
  OR2_X1 U43bar ( .A1(abar[3]), .A2(bbar[13]), .ZN(ybar[61]) );
  AND2_X1 U44 ( .A1(a[3]), .A2(b[12]), .ZN(y[60]) );
  OR2_X1 U44bar ( .A1(abar[3]), .A2(bbar[12]), .ZN(ybar[60]) );
  AND2_X1 U45 ( .A1(b[5]), .A2(a[0]), .ZN(y[5]) );
  OR2_X1 U45bar ( .A1(bbar[5]), .A2(abar[0]), .ZN(ybar[5]) );
  AND2_X1 U46 ( .A1(a[3]), .A2(b[11]), .ZN(y[59]) );
  OR2_X1 U46bar ( .A1(abar[3]), .A2(bbar[11]), .ZN(ybar[59]) );
  AND2_X1 U47 ( .A1(a[3]), .A2(b[10]), .ZN(y[58]) );
  OR2_X1 U47bar ( .A1(abar[3]), .A2(bbar[10]), .ZN(ybar[58]) );
  AND2_X1 U48 ( .A1(a[3]), .A2(b[9]), .ZN(y[57]) );
  OR2_X1 U48bar ( .A1(abar[3]), .A2(bbar[9]), .ZN(ybar[57]) );
  AND2_X1 U49 ( .A1(a[3]), .A2(b[8]), .ZN(y[56]) );
  OR2_X1 U49bar ( .A1(abar[3]), .A2(bbar[8]), .ZN(ybar[56]) );
  AND2_X1 U50 ( .A1(a[3]), .A2(b[7]), .ZN(y[55]) );
  OR2_X1 U50bar ( .A1(abar[3]), .A2(bbar[7]), .ZN(ybar[55]) );
  AND2_X1 U51 ( .A1(a[3]), .A2(b[6]), .ZN(y[54]) );
  OR2_X1 U51bar ( .A1(abar[3]), .A2(bbar[6]), .ZN(ybar[54]) );
  AND2_X1 U52 ( .A1(a[3]), .A2(b[5]), .ZN(y[53]) );
  OR2_X1 U52bar ( .A1(abar[3]), .A2(bbar[5]), .ZN(ybar[53]) );
  AND2_X1 U53 ( .A1(a[3]), .A2(b[4]), .ZN(y[52]) );
  OR2_X1 U53bar ( .A1(abar[3]), .A2(bbar[4]), .ZN(ybar[52]) );
  AND2_X1 U54 ( .A1(a[3]), .A2(b[3]), .ZN(y[51]) );
  OR2_X1 U54bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[51]) );
  AND2_X1 U55 ( .A1(a[3]), .A2(b[2]), .ZN(y[50]) );
  OR2_X1 U55bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[50]) );
  AND2_X1 U56 ( .A1(b[4]), .A2(a[0]), .ZN(y[4]) );
  OR2_X1 U56bar ( .A1(bbar[4]), .A2(abar[0]), .ZN(ybar[4]) );
  AND2_X1 U57 ( .A1(a[3]), .A2(b[1]), .ZN(y[49]) );
  OR2_X1 U57bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[49]) );
  AND2_X1 U58 ( .A1(a[3]), .A2(b[0]), .ZN(y[48]) );
  OR2_X1 U58bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[48]) );
  AND2_X1 U59 ( .A1(a[2]), .A2(b[15]), .ZN(y[47]) );
  OR2_X1 U59bar ( .A1(abar[2]), .A2(bbar[15]), .ZN(ybar[47]) );
  AND2_X1 U60 ( .A1(a[2]), .A2(b[14]), .ZN(y[46]) );
  OR2_X1 U60bar ( .A1(abar[2]), .A2(bbar[14]), .ZN(ybar[46]) );
  AND2_X1 U61 ( .A1(a[2]), .A2(b[13]), .ZN(y[45]) );
  OR2_X1 U61bar ( .A1(abar[2]), .A2(bbar[13]), .ZN(ybar[45]) );
  AND2_X1 U62 ( .A1(a[2]), .A2(b[12]), .ZN(y[44]) );
  OR2_X1 U62bar ( .A1(abar[2]), .A2(bbar[12]), .ZN(ybar[44]) );
  AND2_X1 U63 ( .A1(a[2]), .A2(b[11]), .ZN(y[43]) );
  OR2_X1 U63bar ( .A1(abar[2]), .A2(bbar[11]), .ZN(ybar[43]) );
  AND2_X1 U64 ( .A1(a[2]), .A2(b[10]), .ZN(y[42]) );
  OR2_X1 U64bar ( .A1(abar[2]), .A2(bbar[10]), .ZN(ybar[42]) );
  AND2_X1 U65 ( .A1(a[2]), .A2(b[9]), .ZN(y[41]) );
  OR2_X1 U65bar ( .A1(abar[2]), .A2(bbar[9]), .ZN(ybar[41]) );
  AND2_X1 U66 ( .A1(a[2]), .A2(b[8]), .ZN(y[40]) );
  OR2_X1 U66bar ( .A1(abar[2]), .A2(bbar[8]), .ZN(ybar[40]) );
  AND2_X1 U67 ( .A1(b[3]), .A2(a[0]), .ZN(y[3]) );
  OR2_X1 U67bar ( .A1(bbar[3]), .A2(abar[0]), .ZN(ybar[3]) );
  AND2_X1 U68 ( .A1(a[2]), .A2(b[7]), .ZN(y[39]) );
  OR2_X1 U68bar ( .A1(abar[2]), .A2(bbar[7]), .ZN(ybar[39]) );
  AND2_X1 U69 ( .A1(a[2]), .A2(b[6]), .ZN(y[38]) );
  OR2_X1 U69bar ( .A1(abar[2]), .A2(bbar[6]), .ZN(ybar[38]) );
  AND2_X1 U70 ( .A1(a[2]), .A2(b[5]), .ZN(y[37]) );
  OR2_X1 U70bar ( .A1(abar[2]), .A2(bbar[5]), .ZN(ybar[37]) );
  AND2_X1 U71 ( .A1(a[2]), .A2(b[4]), .ZN(y[36]) );
  OR2_X1 U71bar ( .A1(abar[2]), .A2(bbar[4]), .ZN(ybar[36]) );
  AND2_X1 U72 ( .A1(a[2]), .A2(b[3]), .ZN(y[35]) );
  OR2_X1 U72bar ( .A1(abar[2]), .A2(bbar[3]), .ZN(ybar[35]) );
  AND2_X1 U73 ( .A1(a[2]), .A2(b[2]), .ZN(y[34]) );
  OR2_X1 U73bar ( .A1(abar[2]), .A2(bbar[2]), .ZN(ybar[34]) );
  AND2_X1 U74 ( .A1(a[2]), .A2(b[1]), .ZN(y[33]) );
  OR2_X1 U74bar ( .A1(abar[2]), .A2(bbar[1]), .ZN(ybar[33]) );
  AND2_X1 U75 ( .A1(a[2]), .A2(b[0]), .ZN(y[32]) );
  OR2_X1 U75bar ( .A1(abar[2]), .A2(bbar[0]), .ZN(ybar[32]) );
  AND2_X1 U76 ( .A1(a[1]), .A2(b[15]), .ZN(y[31]) );
  OR2_X1 U76bar ( .A1(abar[1]), .A2(bbar[15]), .ZN(ybar[31]) );
  AND2_X1 U77 ( .A1(a[1]), .A2(b[14]), .ZN(y[30]) );
  OR2_X1 U77bar ( .A1(abar[1]), .A2(bbar[14]), .ZN(ybar[30]) );
  AND2_X1 U78 ( .A1(b[2]), .A2(a[0]), .ZN(y[2]) );
  OR2_X1 U78bar ( .A1(bbar[2]), .A2(abar[0]), .ZN(ybar[2]) );
  AND2_X1 U79 ( .A1(a[1]), .A2(b[13]), .ZN(y[29]) );
  OR2_X1 U79bar ( .A1(abar[1]), .A2(bbar[13]), .ZN(ybar[29]) );
  AND2_X1 U80 ( .A1(a[1]), .A2(b[12]), .ZN(y[28]) );
  OR2_X1 U80bar ( .A1(abar[1]), .A2(bbar[12]), .ZN(ybar[28]) );
  AND2_X1 U81 ( .A1(a[1]), .A2(b[11]), .ZN(y[27]) );
  OR2_X1 U81bar ( .A1(abar[1]), .A2(bbar[11]), .ZN(ybar[27]) );
  AND2_X1 U82 ( .A1(a[1]), .A2(b[10]), .ZN(y[26]) );
  OR2_X1 U82bar ( .A1(abar[1]), .A2(bbar[10]), .ZN(ybar[26]) );
  AND2_X1 U83 ( .A1(a[1]), .A2(b[9]), .ZN(y[25]) );
  OR2_X1 U83bar ( .A1(abar[1]), .A2(bbar[9]), .ZN(ybar[25]) );
  AND2_X1 U84 ( .A1(a[15]), .A2(b[15]), .ZN(y[255]) );
  OR2_X1 U84bar ( .A1(abar[15]), .A2(bbar[15]), .ZN(ybar[255]) );
  AND2_X1 U85 ( .A1(a[15]), .A2(b[14]), .ZN(y[254]) );
  OR2_X1 U85bar ( .A1(abar[15]), .A2(bbar[14]), .ZN(ybar[254]) );
  AND2_X1 U86 ( .A1(a[15]), .A2(b[13]), .ZN(y[253]) );
  OR2_X1 U86bar ( .A1(abar[15]), .A2(bbar[13]), .ZN(ybar[253]) );
  AND2_X1 U87 ( .A1(a[15]), .A2(b[12]), .ZN(y[252]) );
  OR2_X1 U87bar ( .A1(abar[15]), .A2(bbar[12]), .ZN(ybar[252]) );
  AND2_X1 U88 ( .A1(a[15]), .A2(b[11]), .ZN(y[251]) );
  OR2_X1 U88bar ( .A1(abar[15]), .A2(bbar[11]), .ZN(ybar[251]) );
  AND2_X1 U89 ( .A1(a[15]), .A2(b[10]), .ZN(y[250]) );
  OR2_X1 U89bar ( .A1(abar[15]), .A2(bbar[10]), .ZN(ybar[250]) );
  AND2_X1 U90 ( .A1(a[1]), .A2(b[8]), .ZN(y[24]) );
  OR2_X1 U90bar ( .A1(abar[1]), .A2(bbar[8]), .ZN(ybar[24]) );
  AND2_X1 U91 ( .A1(a[15]), .A2(b[9]), .ZN(y[249]) );
  OR2_X1 U91bar ( .A1(abar[15]), .A2(bbar[9]), .ZN(ybar[249]) );
  AND2_X1 U92 ( .A1(a[15]), .A2(b[8]), .ZN(y[248]) );
  OR2_X1 U92bar ( .A1(abar[15]), .A2(bbar[8]), .ZN(ybar[248]) );
  AND2_X1 U93 ( .A1(a[15]), .A2(b[7]), .ZN(y[247]) );
  OR2_X1 U93bar ( .A1(abar[15]), .A2(bbar[7]), .ZN(ybar[247]) );
  AND2_X1 U94 ( .A1(a[15]), .A2(b[6]), .ZN(y[246]) );
  OR2_X1 U94bar ( .A1(abar[15]), .A2(bbar[6]), .ZN(ybar[246]) );
  AND2_X1 U95 ( .A1(a[15]), .A2(b[5]), .ZN(y[245]) );
  OR2_X1 U95bar ( .A1(abar[15]), .A2(bbar[5]), .ZN(ybar[245]) );
  AND2_X1 U96 ( .A1(a[15]), .A2(b[4]), .ZN(y[244]) );
  OR2_X1 U96bar ( .A1(abar[15]), .A2(bbar[4]), .ZN(ybar[244]) );
  AND2_X1 U97 ( .A1(a[15]), .A2(b[3]), .ZN(y[243]) );
  OR2_X1 U97bar ( .A1(abar[15]), .A2(bbar[3]), .ZN(ybar[243]) );
  AND2_X1 U98 ( .A1(a[15]), .A2(b[2]), .ZN(y[242]) );
  OR2_X1 U98bar ( .A1(abar[15]), .A2(bbar[2]), .ZN(ybar[242]) );
  AND2_X1 U99 ( .A1(a[15]), .A2(b[1]), .ZN(y[241]) );
  OR2_X1 U99bar ( .A1(abar[15]), .A2(bbar[1]), .ZN(ybar[241]) );
  AND2_X1 U100 ( .A1(a[15]), .A2(b[0]), .ZN(y[240]) );
  OR2_X1 U100bar ( .A1(abar[15]), .A2(bbar[0]), .ZN(ybar[240]) );
  AND2_X1 U101 ( .A1(a[1]), .A2(b[7]), .ZN(y[23]) );
  OR2_X1 U101bar ( .A1(abar[1]), .A2(bbar[7]), .ZN(ybar[23]) );
  AND2_X1 U102 ( .A1(a[14]), .A2(b[15]), .ZN(y[239]) );
  OR2_X1 U102bar ( .A1(abar[14]), .A2(bbar[15]), .ZN(ybar[239]) );
  AND2_X1 U103 ( .A1(a[14]), .A2(b[14]), .ZN(y[238]) );
  OR2_X1 U103bar ( .A1(abar[14]), .A2(bbar[14]), .ZN(ybar[238]) );
  AND2_X1 U104 ( .A1(a[14]), .A2(b[13]), .ZN(y[237]) );
  OR2_X1 U104bar ( .A1(abar[14]), .A2(bbar[13]), .ZN(ybar[237]) );
  AND2_X1 U105 ( .A1(a[14]), .A2(b[12]), .ZN(y[236]) );
  OR2_X1 U105bar ( .A1(abar[14]), .A2(bbar[12]), .ZN(ybar[236]) );
  AND2_X1 U106 ( .A1(a[14]), .A2(b[11]), .ZN(y[235]) );
  OR2_X1 U106bar ( .A1(abar[14]), .A2(bbar[11]), .ZN(ybar[235]) );
  AND2_X1 U107 ( .A1(a[14]), .A2(b[10]), .ZN(y[234]) );
  OR2_X1 U107bar ( .A1(abar[14]), .A2(bbar[10]), .ZN(ybar[234]) );
  AND2_X1 U108 ( .A1(a[14]), .A2(b[9]), .ZN(y[233]) );
  OR2_X1 U108bar ( .A1(abar[14]), .A2(bbar[9]), .ZN(ybar[233]) );
  AND2_X1 U109 ( .A1(a[14]), .A2(b[8]), .ZN(y[232]) );
  OR2_X1 U109bar ( .A1(abar[14]), .A2(bbar[8]), .ZN(ybar[232]) );
  AND2_X1 U110 ( .A1(a[14]), .A2(b[7]), .ZN(y[231]) );
  OR2_X1 U110bar ( .A1(abar[14]), .A2(bbar[7]), .ZN(ybar[231]) );
  AND2_X1 U111 ( .A1(a[14]), .A2(b[6]), .ZN(y[230]) );
  OR2_X1 U111bar ( .A1(abar[14]), .A2(bbar[6]), .ZN(ybar[230]) );
  AND2_X1 U112 ( .A1(a[1]), .A2(b[6]), .ZN(y[22]) );
  OR2_X1 U112bar ( .A1(abar[1]), .A2(bbar[6]), .ZN(ybar[22]) );
  AND2_X1 U113 ( .A1(a[14]), .A2(b[5]), .ZN(y[229]) );
  OR2_X1 U113bar ( .A1(abar[14]), .A2(bbar[5]), .ZN(ybar[229]) );
  AND2_X1 U114 ( .A1(a[14]), .A2(b[4]), .ZN(y[228]) );
  OR2_X1 U114bar ( .A1(abar[14]), .A2(bbar[4]), .ZN(ybar[228]) );
  AND2_X1 U115 ( .A1(a[14]), .A2(b[3]), .ZN(y[227]) );
  OR2_X1 U115bar ( .A1(abar[14]), .A2(bbar[3]), .ZN(ybar[227]) );
  AND2_X1 U116 ( .A1(a[14]), .A2(b[2]), .ZN(y[226]) );
  OR2_X1 U116bar ( .A1(abar[14]), .A2(bbar[2]), .ZN(ybar[226]) );
  AND2_X1 U117 ( .A1(a[14]), .A2(b[1]), .ZN(y[225]) );
  OR2_X1 U117bar ( .A1(abar[14]), .A2(bbar[1]), .ZN(ybar[225]) );
  AND2_X1 U118 ( .A1(a[14]), .A2(b[0]), .ZN(y[224]) );
  OR2_X1 U118bar ( .A1(abar[14]), .A2(bbar[0]), .ZN(ybar[224]) );
  AND2_X1 U119 ( .A1(a[13]), .A2(b[15]), .ZN(y[223]) );
  OR2_X1 U119bar ( .A1(abar[13]), .A2(bbar[15]), .ZN(ybar[223]) );
  AND2_X1 U120 ( .A1(a[13]), .A2(b[14]), .ZN(y[222]) );
  OR2_X1 U120bar ( .A1(abar[13]), .A2(bbar[14]), .ZN(ybar[222]) );
  AND2_X1 U121 ( .A1(a[13]), .A2(b[13]), .ZN(y[221]) );
  OR2_X1 U121bar ( .A1(abar[13]), .A2(bbar[13]), .ZN(ybar[221]) );
  AND2_X1 U122 ( .A1(a[13]), .A2(b[12]), .ZN(y[220]) );
  OR2_X1 U122bar ( .A1(abar[13]), .A2(bbar[12]), .ZN(ybar[220]) );
  AND2_X1 U123 ( .A1(a[1]), .A2(b[5]), .ZN(y[21]) );
  OR2_X1 U123bar ( .A1(abar[1]), .A2(bbar[5]), .ZN(ybar[21]) );
  AND2_X1 U124 ( .A1(a[13]), .A2(b[11]), .ZN(y[219]) );
  OR2_X1 U124bar ( .A1(abar[13]), .A2(bbar[11]), .ZN(ybar[219]) );
  AND2_X1 U125 ( .A1(a[13]), .A2(b[10]), .ZN(y[218]) );
  OR2_X1 U125bar ( .A1(abar[13]), .A2(bbar[10]), .ZN(ybar[218]) );
  AND2_X1 U126 ( .A1(a[13]), .A2(b[9]), .ZN(y[217]) );
  OR2_X1 U126bar ( .A1(abar[13]), .A2(bbar[9]), .ZN(ybar[217]) );
  AND2_X1 U127 ( .A1(a[13]), .A2(b[8]), .ZN(y[216]) );
  OR2_X1 U127bar ( .A1(abar[13]), .A2(bbar[8]), .ZN(ybar[216]) );
  AND2_X1 U128 ( .A1(a[13]), .A2(b[7]), .ZN(y[215]) );
  OR2_X1 U128bar ( .A1(abar[13]), .A2(bbar[7]), .ZN(ybar[215]) );
  AND2_X1 U129 ( .A1(a[13]), .A2(b[6]), .ZN(y[214]) );
  OR2_X1 U129bar ( .A1(abar[13]), .A2(bbar[6]), .ZN(ybar[214]) );
  AND2_X1 U130 ( .A1(a[13]), .A2(b[5]), .ZN(y[213]) );
  OR2_X1 U130bar ( .A1(abar[13]), .A2(bbar[5]), .ZN(ybar[213]) );
  AND2_X1 U131 ( .A1(a[13]), .A2(b[4]), .ZN(y[212]) );
  OR2_X1 U131bar ( .A1(abar[13]), .A2(bbar[4]), .ZN(ybar[212]) );
  AND2_X1 U132 ( .A1(a[13]), .A2(b[3]), .ZN(y[211]) );
  OR2_X1 U132bar ( .A1(abar[13]), .A2(bbar[3]), .ZN(ybar[211]) );
  AND2_X1 U133 ( .A1(a[13]), .A2(b[2]), .ZN(y[210]) );
  OR2_X1 U133bar ( .A1(abar[13]), .A2(bbar[2]), .ZN(ybar[210]) );
  AND2_X1 U134 ( .A1(a[1]), .A2(b[4]), .ZN(y[20]) );
  OR2_X1 U134bar ( .A1(abar[1]), .A2(bbar[4]), .ZN(ybar[20]) );
  AND2_X1 U135 ( .A1(a[13]), .A2(b[1]), .ZN(y[209]) );
  OR2_X1 U135bar ( .A1(abar[13]), .A2(bbar[1]), .ZN(ybar[209]) );
  AND2_X1 U136 ( .A1(a[13]), .A2(b[0]), .ZN(y[208]) );
  OR2_X1 U136bar ( .A1(abar[13]), .A2(bbar[0]), .ZN(ybar[208]) );
  AND2_X1 U137 ( .A1(a[12]), .A2(b[15]), .ZN(y[207]) );
  OR2_X1 U137bar ( .A1(abar[12]), .A2(bbar[15]), .ZN(ybar[207]) );
  AND2_X1 U138 ( .A1(a[12]), .A2(b[14]), .ZN(y[206]) );
  OR2_X1 U138bar ( .A1(abar[12]), .A2(bbar[14]), .ZN(ybar[206]) );
  AND2_X1 U139 ( .A1(a[12]), .A2(b[13]), .ZN(y[205]) );
  OR2_X1 U139bar ( .A1(abar[12]), .A2(bbar[13]), .ZN(ybar[205]) );
  AND2_X1 U140 ( .A1(a[12]), .A2(b[12]), .ZN(y[204]) );
  OR2_X1 U140bar ( .A1(abar[12]), .A2(bbar[12]), .ZN(ybar[204]) );
  AND2_X1 U141 ( .A1(a[12]), .A2(b[11]), .ZN(y[203]) );
  OR2_X1 U141bar ( .A1(abar[12]), .A2(bbar[11]), .ZN(ybar[203]) );
  AND2_X1 U142 ( .A1(a[12]), .A2(b[10]), .ZN(y[202]) );
  OR2_X1 U142bar ( .A1(abar[12]), .A2(bbar[10]), .ZN(ybar[202]) );
  AND2_X1 U143 ( .A1(a[12]), .A2(b[9]), .ZN(y[201]) );
  OR2_X1 U143bar ( .A1(abar[12]), .A2(bbar[9]), .ZN(ybar[201]) );
  AND2_X1 U144 ( .A1(a[12]), .A2(b[8]), .ZN(y[200]) );
  OR2_X1 U144bar ( .A1(abar[12]), .A2(bbar[8]), .ZN(ybar[200]) );
  AND2_X1 U145 ( .A1(b[1]), .A2(a[0]), .ZN(y[1]) );
  OR2_X1 U145bar ( .A1(bbar[1]), .A2(abar[0]), .ZN(ybar[1]) );
  AND2_X1 U146 ( .A1(a[1]), .A2(b[3]), .ZN(y[19]) );
  OR2_X1 U146bar ( .A1(abar[1]), .A2(bbar[3]), .ZN(ybar[19]) );
  AND2_X1 U147 ( .A1(a[12]), .A2(b[7]), .ZN(y[199]) );
  OR2_X1 U147bar ( .A1(abar[12]), .A2(bbar[7]), .ZN(ybar[199]) );
  AND2_X1 U148 ( .A1(a[12]), .A2(b[6]), .ZN(y[198]) );
  OR2_X1 U148bar ( .A1(abar[12]), .A2(bbar[6]), .ZN(ybar[198]) );
  AND2_X1 U149 ( .A1(a[12]), .A2(b[5]), .ZN(y[197]) );
  OR2_X1 U149bar ( .A1(abar[12]), .A2(bbar[5]), .ZN(ybar[197]) );
  AND2_X1 U150 ( .A1(a[12]), .A2(b[4]), .ZN(y[196]) );
  OR2_X1 U150bar ( .A1(abar[12]), .A2(bbar[4]), .ZN(ybar[196]) );
  AND2_X1 U151 ( .A1(a[12]), .A2(b[3]), .ZN(y[195]) );
  OR2_X1 U151bar ( .A1(abar[12]), .A2(bbar[3]), .ZN(ybar[195]) );
  AND2_X1 U152 ( .A1(a[12]), .A2(b[2]), .ZN(y[194]) );
  OR2_X1 U152bar ( .A1(abar[12]), .A2(bbar[2]), .ZN(ybar[194]) );
  AND2_X1 U153 ( .A1(a[12]), .A2(b[1]), .ZN(y[193]) );
  OR2_X1 U153bar ( .A1(abar[12]), .A2(bbar[1]), .ZN(ybar[193]) );
  AND2_X1 U154 ( .A1(a[12]), .A2(b[0]), .ZN(y[192]) );
  OR2_X1 U154bar ( .A1(abar[12]), .A2(bbar[0]), .ZN(ybar[192]) );
  AND2_X1 U155 ( .A1(a[11]), .A2(b[15]), .ZN(y[191]) );
  OR2_X1 U155bar ( .A1(abar[11]), .A2(bbar[15]), .ZN(ybar[191]) );
  AND2_X1 U156 ( .A1(a[11]), .A2(b[14]), .ZN(y[190]) );
  OR2_X1 U156bar ( .A1(abar[11]), .A2(bbar[14]), .ZN(ybar[190]) );
  AND2_X1 U157 ( .A1(a[1]), .A2(b[2]), .ZN(y[18]) );
  OR2_X1 U157bar ( .A1(abar[1]), .A2(bbar[2]), .ZN(ybar[18]) );
  AND2_X1 U158 ( .A1(a[11]), .A2(b[13]), .ZN(y[189]) );
  OR2_X1 U158bar ( .A1(abar[11]), .A2(bbar[13]), .ZN(ybar[189]) );
  AND2_X1 U159 ( .A1(a[11]), .A2(b[12]), .ZN(y[188]) );
  OR2_X1 U159bar ( .A1(abar[11]), .A2(bbar[12]), .ZN(ybar[188]) );
  AND2_X1 U160 ( .A1(a[11]), .A2(b[11]), .ZN(y[187]) );
  OR2_X1 U160bar ( .A1(abar[11]), .A2(bbar[11]), .ZN(ybar[187]) );
  AND2_X1 U161 ( .A1(a[11]), .A2(b[10]), .ZN(y[186]) );
  OR2_X1 U161bar ( .A1(abar[11]), .A2(bbar[10]), .ZN(ybar[186]) );
  AND2_X1 U162 ( .A1(a[11]), .A2(b[9]), .ZN(y[185]) );
  OR2_X1 U162bar ( .A1(abar[11]), .A2(bbar[9]), .ZN(ybar[185]) );
  AND2_X1 U163 ( .A1(a[11]), .A2(b[8]), .ZN(y[184]) );
  OR2_X1 U163bar ( .A1(abar[11]), .A2(bbar[8]), .ZN(ybar[184]) );
  AND2_X1 U164 ( .A1(a[11]), .A2(b[7]), .ZN(y[183]) );
  OR2_X1 U164bar ( .A1(abar[11]), .A2(bbar[7]), .ZN(ybar[183]) );
  AND2_X1 U165 ( .A1(a[11]), .A2(b[6]), .ZN(y[182]) );
  OR2_X1 U165bar ( .A1(abar[11]), .A2(bbar[6]), .ZN(ybar[182]) );
  AND2_X1 U166 ( .A1(a[11]), .A2(b[5]), .ZN(y[181]) );
  OR2_X1 U166bar ( .A1(abar[11]), .A2(bbar[5]), .ZN(ybar[181]) );
  AND2_X1 U167 ( .A1(a[11]), .A2(b[4]), .ZN(y[180]) );
  OR2_X1 U167bar ( .A1(abar[11]), .A2(bbar[4]), .ZN(ybar[180]) );
  AND2_X1 U168 ( .A1(a[1]), .A2(b[1]), .ZN(y[17]) );
  OR2_X1 U168bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[17]) );
  AND2_X1 U169 ( .A1(a[11]), .A2(b[3]), .ZN(y[179]) );
  OR2_X1 U169bar ( .A1(abar[11]), .A2(bbar[3]), .ZN(ybar[179]) );
  AND2_X1 U170 ( .A1(a[11]), .A2(b[2]), .ZN(y[178]) );
  OR2_X1 U170bar ( .A1(abar[11]), .A2(bbar[2]), .ZN(ybar[178]) );
  AND2_X1 U171 ( .A1(a[11]), .A2(b[1]), .ZN(y[177]) );
  OR2_X1 U171bar ( .A1(abar[11]), .A2(bbar[1]), .ZN(ybar[177]) );
  AND2_X1 U172 ( .A1(a[11]), .A2(b[0]), .ZN(y[176]) );
  OR2_X1 U172bar ( .A1(abar[11]), .A2(bbar[0]), .ZN(ybar[176]) );
  AND2_X1 U173 ( .A1(a[10]), .A2(b[15]), .ZN(y[175]) );
  OR2_X1 U173bar ( .A1(abar[10]), .A2(bbar[15]), .ZN(ybar[175]) );
  AND2_X1 U174 ( .A1(a[10]), .A2(b[14]), .ZN(y[174]) );
  OR2_X1 U174bar ( .A1(abar[10]), .A2(bbar[14]), .ZN(ybar[174]) );
  AND2_X1 U175 ( .A1(a[10]), .A2(b[13]), .ZN(y[173]) );
  OR2_X1 U175bar ( .A1(abar[10]), .A2(bbar[13]), .ZN(ybar[173]) );
  AND2_X1 U176 ( .A1(a[10]), .A2(b[12]), .ZN(y[172]) );
  OR2_X1 U176bar ( .A1(abar[10]), .A2(bbar[12]), .ZN(ybar[172]) );
  AND2_X1 U177 ( .A1(a[10]), .A2(b[11]), .ZN(y[171]) );
  OR2_X1 U177bar ( .A1(abar[10]), .A2(bbar[11]), .ZN(ybar[171]) );
  AND2_X1 U178 ( .A1(a[10]), .A2(b[10]), .ZN(y[170]) );
  OR2_X1 U178bar ( .A1(abar[10]), .A2(bbar[10]), .ZN(ybar[170]) );
  AND2_X1 U179 ( .A1(a[1]), .A2(b[0]), .ZN(y[16]) );
  OR2_X1 U179bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[16]) );
  AND2_X1 U180 ( .A1(a[10]), .A2(b[9]), .ZN(y[169]) );
  OR2_X1 U180bar ( .A1(abar[10]), .A2(bbar[9]), .ZN(ybar[169]) );
  AND2_X1 U181 ( .A1(a[10]), .A2(b[8]), .ZN(y[168]) );
  OR2_X1 U181bar ( .A1(abar[10]), .A2(bbar[8]), .ZN(ybar[168]) );
  AND2_X1 U182 ( .A1(a[10]), .A2(b[7]), .ZN(y[167]) );
  OR2_X1 U182bar ( .A1(abar[10]), .A2(bbar[7]), .ZN(ybar[167]) );
  AND2_X1 U183 ( .A1(a[10]), .A2(b[6]), .ZN(y[166]) );
  OR2_X1 U183bar ( .A1(abar[10]), .A2(bbar[6]), .ZN(ybar[166]) );
  AND2_X1 U184 ( .A1(a[10]), .A2(b[5]), .ZN(y[165]) );
  OR2_X1 U184bar ( .A1(abar[10]), .A2(bbar[5]), .ZN(ybar[165]) );
  AND2_X1 U185 ( .A1(a[10]), .A2(b[4]), .ZN(y[164]) );
  OR2_X1 U185bar ( .A1(abar[10]), .A2(bbar[4]), .ZN(ybar[164]) );
  AND2_X1 U186 ( .A1(a[10]), .A2(b[3]), .ZN(y[163]) );
  OR2_X1 U186bar ( .A1(abar[10]), .A2(bbar[3]), .ZN(ybar[163]) );
  AND2_X1 U187 ( .A1(a[10]), .A2(b[2]), .ZN(y[162]) );
  OR2_X1 U187bar ( .A1(abar[10]), .A2(bbar[2]), .ZN(ybar[162]) );
  AND2_X1 U188 ( .A1(a[10]), .A2(b[1]), .ZN(y[161]) );
  OR2_X1 U188bar ( .A1(abar[10]), .A2(bbar[1]), .ZN(ybar[161]) );
  AND2_X1 U189 ( .A1(a[10]), .A2(b[0]), .ZN(y[160]) );
  OR2_X1 U189bar ( .A1(abar[10]), .A2(bbar[0]), .ZN(ybar[160]) );
  AND2_X1 U190 ( .A1(b[15]), .A2(a[0]), .ZN(y[15]) );
  OR2_X1 U190bar ( .A1(bbar[15]), .A2(abar[0]), .ZN(ybar[15]) );
  AND2_X1 U191 ( .A1(a[9]), .A2(b[15]), .ZN(y[159]) );
  OR2_X1 U191bar ( .A1(abar[9]), .A2(bbar[15]), .ZN(ybar[159]) );
  AND2_X1 U192 ( .A1(a[9]), .A2(b[14]), .ZN(y[158]) );
  OR2_X1 U192bar ( .A1(abar[9]), .A2(bbar[14]), .ZN(ybar[158]) );
  AND2_X1 U193 ( .A1(a[9]), .A2(b[13]), .ZN(y[157]) );
  OR2_X1 U193bar ( .A1(abar[9]), .A2(bbar[13]), .ZN(ybar[157]) );
  AND2_X1 U194 ( .A1(a[9]), .A2(b[12]), .ZN(y[156]) );
  OR2_X1 U194bar ( .A1(abar[9]), .A2(bbar[12]), .ZN(ybar[156]) );
  AND2_X1 U195 ( .A1(a[9]), .A2(b[11]), .ZN(y[155]) );
  OR2_X1 U195bar ( .A1(abar[9]), .A2(bbar[11]), .ZN(ybar[155]) );
  AND2_X1 U196 ( .A1(a[9]), .A2(b[10]), .ZN(y[154]) );
  OR2_X1 U196bar ( .A1(abar[9]), .A2(bbar[10]), .ZN(ybar[154]) );
  AND2_X1 U197 ( .A1(a[9]), .A2(b[9]), .ZN(y[153]) );
  OR2_X1 U197bar ( .A1(abar[9]), .A2(bbar[9]), .ZN(ybar[153]) );
  AND2_X1 U198 ( .A1(a[9]), .A2(b[8]), .ZN(y[152]) );
  OR2_X1 U198bar ( .A1(abar[9]), .A2(bbar[8]), .ZN(ybar[152]) );
  AND2_X1 U199 ( .A1(a[9]), .A2(b[7]), .ZN(y[151]) );
  OR2_X1 U199bar ( .A1(abar[9]), .A2(bbar[7]), .ZN(ybar[151]) );
  AND2_X1 U200 ( .A1(a[9]), .A2(b[6]), .ZN(y[150]) );
  OR2_X1 U200bar ( .A1(abar[9]), .A2(bbar[6]), .ZN(ybar[150]) );
  AND2_X1 U201 ( .A1(b[14]), .A2(a[0]), .ZN(y[14]) );
  OR2_X1 U201bar ( .A1(bbar[14]), .A2(abar[0]), .ZN(ybar[14]) );
  AND2_X1 U202 ( .A1(a[9]), .A2(b[5]), .ZN(y[149]) );
  OR2_X1 U202bar ( .A1(abar[9]), .A2(bbar[5]), .ZN(ybar[149]) );
  AND2_X1 U203 ( .A1(a[9]), .A2(b[4]), .ZN(y[148]) );
  OR2_X1 U203bar ( .A1(abar[9]), .A2(bbar[4]), .ZN(ybar[148]) );
  AND2_X1 U204 ( .A1(a[9]), .A2(b[3]), .ZN(y[147]) );
  OR2_X1 U204bar ( .A1(abar[9]), .A2(bbar[3]), .ZN(ybar[147]) );
  AND2_X1 U205 ( .A1(a[9]), .A2(b[2]), .ZN(y[146]) );
  OR2_X1 U205bar ( .A1(abar[9]), .A2(bbar[2]), .ZN(ybar[146]) );
  AND2_X1 U206 ( .A1(a[9]), .A2(b[1]), .ZN(y[145]) );
  OR2_X1 U206bar ( .A1(abar[9]), .A2(bbar[1]), .ZN(ybar[145]) );
  AND2_X1 U207 ( .A1(a[9]), .A2(b[0]), .ZN(y[144]) );
  OR2_X1 U207bar ( .A1(abar[9]), .A2(bbar[0]), .ZN(ybar[144]) );
  AND2_X1 U208 ( .A1(a[8]), .A2(b[15]), .ZN(y[143]) );
  OR2_X1 U208bar ( .A1(abar[8]), .A2(bbar[15]), .ZN(ybar[143]) );
  AND2_X1 U209 ( .A1(a[8]), .A2(b[14]), .ZN(y[142]) );
  OR2_X1 U209bar ( .A1(abar[8]), .A2(bbar[14]), .ZN(ybar[142]) );
  AND2_X1 U210 ( .A1(a[8]), .A2(b[13]), .ZN(y[141]) );
  OR2_X1 U210bar ( .A1(abar[8]), .A2(bbar[13]), .ZN(ybar[141]) );
  AND2_X1 U211 ( .A1(a[8]), .A2(b[12]), .ZN(y[140]) );
  OR2_X1 U211bar ( .A1(abar[8]), .A2(bbar[12]), .ZN(ybar[140]) );
  AND2_X1 U212 ( .A1(b[13]), .A2(a[0]), .ZN(y[13]) );
  OR2_X1 U212bar ( .A1(bbar[13]), .A2(abar[0]), .ZN(ybar[13]) );
  AND2_X1 U213 ( .A1(a[8]), .A2(b[11]), .ZN(y[139]) );
  OR2_X1 U213bar ( .A1(abar[8]), .A2(bbar[11]), .ZN(ybar[139]) );
  AND2_X1 U214 ( .A1(a[8]), .A2(b[10]), .ZN(y[138]) );
  OR2_X1 U214bar ( .A1(abar[8]), .A2(bbar[10]), .ZN(ybar[138]) );
  AND2_X1 U215 ( .A1(a[8]), .A2(b[9]), .ZN(y[137]) );
  OR2_X1 U215bar ( .A1(abar[8]), .A2(bbar[9]), .ZN(ybar[137]) );
  AND2_X1 U216 ( .A1(a[8]), .A2(b[8]), .ZN(y[136]) );
  OR2_X1 U216bar ( .A1(abar[8]), .A2(bbar[8]), .ZN(ybar[136]) );
  AND2_X1 U217 ( .A1(a[8]), .A2(b[7]), .ZN(y[135]) );
  OR2_X1 U217bar ( .A1(abar[8]), .A2(bbar[7]), .ZN(ybar[135]) );
  AND2_X1 U218 ( .A1(a[8]), .A2(b[6]), .ZN(y[134]) );
  OR2_X1 U218bar ( .A1(abar[8]), .A2(bbar[6]), .ZN(ybar[134]) );
  AND2_X1 U219 ( .A1(a[8]), .A2(b[5]), .ZN(y[133]) );
  OR2_X1 U219bar ( .A1(abar[8]), .A2(bbar[5]), .ZN(ybar[133]) );
  AND2_X1 U220 ( .A1(a[8]), .A2(b[4]), .ZN(y[132]) );
  OR2_X1 U220bar ( .A1(abar[8]), .A2(bbar[4]), .ZN(ybar[132]) );
  AND2_X1 U221 ( .A1(a[8]), .A2(b[3]), .ZN(y[131]) );
  OR2_X1 U221bar ( .A1(abar[8]), .A2(bbar[3]), .ZN(ybar[131]) );
  AND2_X1 U222 ( .A1(a[8]), .A2(b[2]), .ZN(y[130]) );
  OR2_X1 U222bar ( .A1(abar[8]), .A2(bbar[2]), .ZN(ybar[130]) );
  AND2_X1 U223 ( .A1(b[12]), .A2(a[0]), .ZN(y[12]) );
  OR2_X1 U223bar ( .A1(bbar[12]), .A2(abar[0]), .ZN(ybar[12]) );
  AND2_X1 U224 ( .A1(a[8]), .A2(b[1]), .ZN(y[129]) );
  OR2_X1 U224bar ( .A1(abar[8]), .A2(bbar[1]), .ZN(ybar[129]) );
  AND2_X1 U225 ( .A1(a[8]), .A2(b[0]), .ZN(y[128]) );
  OR2_X1 U225bar ( .A1(abar[8]), .A2(bbar[0]), .ZN(ybar[128]) );
  AND2_X1 U226 ( .A1(a[7]), .A2(b[15]), .ZN(y[127]) );
  OR2_X1 U226bar ( .A1(abar[7]), .A2(bbar[15]), .ZN(ybar[127]) );
  AND2_X1 U227 ( .A1(a[7]), .A2(b[14]), .ZN(y[126]) );
  OR2_X1 U227bar ( .A1(abar[7]), .A2(bbar[14]), .ZN(ybar[126]) );
  AND2_X1 U228 ( .A1(a[7]), .A2(b[13]), .ZN(y[125]) );
  OR2_X1 U228bar ( .A1(abar[7]), .A2(bbar[13]), .ZN(ybar[125]) );
  AND2_X1 U229 ( .A1(a[7]), .A2(b[12]), .ZN(y[124]) );
  OR2_X1 U229bar ( .A1(abar[7]), .A2(bbar[12]), .ZN(ybar[124]) );
  AND2_X1 U230 ( .A1(a[7]), .A2(b[11]), .ZN(y[123]) );
  OR2_X1 U230bar ( .A1(abar[7]), .A2(bbar[11]), .ZN(ybar[123]) );
  AND2_X1 U231 ( .A1(a[7]), .A2(b[10]), .ZN(y[122]) );
  OR2_X1 U231bar ( .A1(abar[7]), .A2(bbar[10]), .ZN(ybar[122]) );
  AND2_X1 U232 ( .A1(a[7]), .A2(b[9]), .ZN(y[121]) );
  OR2_X1 U232bar ( .A1(abar[7]), .A2(bbar[9]), .ZN(ybar[121]) );
  AND2_X1 U233 ( .A1(a[7]), .A2(b[8]), .ZN(y[120]) );
  OR2_X1 U233bar ( .A1(abar[7]), .A2(bbar[8]), .ZN(ybar[120]) );
  AND2_X1 U234 ( .A1(b[11]), .A2(a[0]), .ZN(y[11]) );
  OR2_X1 U234bar ( .A1(bbar[11]), .A2(abar[0]), .ZN(ybar[11]) );
  AND2_X1 U235 ( .A1(a[7]), .A2(b[7]), .ZN(y[119]) );
  OR2_X1 U235bar ( .A1(abar[7]), .A2(bbar[7]), .ZN(ybar[119]) );
  AND2_X1 U236 ( .A1(a[7]), .A2(b[6]), .ZN(y[118]) );
  OR2_X1 U236bar ( .A1(abar[7]), .A2(bbar[6]), .ZN(ybar[118]) );
  AND2_X1 U237 ( .A1(a[7]), .A2(b[5]), .ZN(y[117]) );
  OR2_X1 U237bar ( .A1(abar[7]), .A2(bbar[5]), .ZN(ybar[117]) );
  AND2_X1 U238 ( .A1(a[7]), .A2(b[4]), .ZN(y[116]) );
  OR2_X1 U238bar ( .A1(abar[7]), .A2(bbar[4]), .ZN(ybar[116]) );
  AND2_X1 U239 ( .A1(a[7]), .A2(b[3]), .ZN(y[115]) );
  OR2_X1 U239bar ( .A1(abar[7]), .A2(bbar[3]), .ZN(ybar[115]) );
  AND2_X1 U240 ( .A1(a[7]), .A2(b[2]), .ZN(y[114]) );
  OR2_X1 U240bar ( .A1(abar[7]), .A2(bbar[2]), .ZN(ybar[114]) );
  AND2_X1 U241 ( .A1(a[7]), .A2(b[1]), .ZN(y[113]) );
  OR2_X1 U241bar ( .A1(abar[7]), .A2(bbar[1]), .ZN(ybar[113]) );
  AND2_X1 U242 ( .A1(a[7]), .A2(b[0]), .ZN(y[112]) );
  OR2_X1 U242bar ( .A1(abar[7]), .A2(bbar[0]), .ZN(ybar[112]) );
  AND2_X1 U243 ( .A1(b[15]), .A2(a[6]), .ZN(y[111]) );
  OR2_X1 U243bar ( .A1(bbar[15]), .A2(abar[6]), .ZN(ybar[111]) );
  AND2_X1 U244 ( .A1(b[14]), .A2(a[6]), .ZN(y[110]) );
  OR2_X1 U244bar ( .A1(bbar[14]), .A2(abar[6]), .ZN(ybar[110]) );
  AND2_X1 U245 ( .A1(b[10]), .A2(a[0]), .ZN(y[10]) );
  OR2_X1 U245bar ( .A1(bbar[10]), .A2(abar[0]), .ZN(ybar[10]) );
  AND2_X1 U246 ( .A1(b[13]), .A2(a[6]), .ZN(y[109]) );
  OR2_X1 U246bar ( .A1(bbar[13]), .A2(abar[6]), .ZN(ybar[109]) );
  AND2_X1 U247 ( .A1(b[12]), .A2(a[6]), .ZN(y[108]) );
  OR2_X1 U247bar ( .A1(bbar[12]), .A2(abar[6]), .ZN(ybar[108]) );
  AND2_X1 U248 ( .A1(b[11]), .A2(a[6]), .ZN(y[107]) );
  OR2_X1 U248bar ( .A1(bbar[11]), .A2(abar[6]), .ZN(ybar[107]) );
  AND2_X1 U249 ( .A1(b[10]), .A2(a[6]), .ZN(y[106]) );
  OR2_X1 U249bar ( .A1(bbar[10]), .A2(abar[6]), .ZN(ybar[106]) );
  AND2_X1 U250 ( .A1(a[6]), .A2(b[9]), .ZN(y[105]) );
  OR2_X1 U250bar ( .A1(abar[6]), .A2(bbar[9]), .ZN(ybar[105]) );
  AND2_X1 U251 ( .A1(b[8]), .A2(a[6]), .ZN(y[104]) );
  OR2_X1 U251bar ( .A1(bbar[8]), .A2(abar[6]), .ZN(ybar[104]) );
  AND2_X1 U252 ( .A1(b[7]), .A2(a[6]), .ZN(y[103]) );
  OR2_X1 U252bar ( .A1(bbar[7]), .A2(abar[6]), .ZN(ybar[103]) );
  AND2_X1 U253 ( .A1(b[6]), .A2(a[6]), .ZN(y[102]) );
  OR2_X1 U253bar ( .A1(bbar[6]), .A2(abar[6]), .ZN(ybar[102]) );
  AND2_X1 U254 ( .A1(b[5]), .A2(a[6]), .ZN(y[101]) );
  OR2_X1 U254bar ( .A1(bbar[5]), .A2(abar[6]), .ZN(ybar[101]) );
  AND2_X1 U255 ( .A1(b[4]), .A2(a[6]), .ZN(y[100]) );
  OR2_X1 U255bar ( .A1(bbar[4]), .A2(abar[6]), .ZN(ybar[100]) );
  AND2_X1 U256 ( .A1(b[0]), .A2(a[0]), .ZN(y[0]) );
  OR2_X1 U256bar ( .A1(bbar[0]), .A2(abar[0]), .ZN(ybar[0]) );
endmodule

module decode_1 ( in, inbar, out, outbar );

  input wire [7:0] in;
  input wire [7:0] inbar;
//input_done

  output wire [255:0] out;
  output wire [255:0] outbar;
//output_done

  wire [15:0] level1;
  wire [31:0] level2;
  wire [15:0] level1bar;
  wire [31:0] level2bar;
//wire_done

  CD2_4 cd_l1_1 ( .a(in[1]), .abar(inbar[1]), .b(in[0]), .bbar(inbar[0]), .y(level1[3:0]), .ybar(level1bar[3:0]) );
  CD2_3 cd_l1_2 ( .a(in[3]), .abar(inbar[3]), .b(in[2]), .bbar(inbar[2]), .y(level1[7:4]), .ybar(level1bar[7:4]) );
  CD2_2 cd_l1_3 ( .a(in[5]), .abar(inbar[5]), .b(in[4]), .bbar(inbar[4]), .y(level1[11:8]), .ybar(level1bar[11:8]) );
  CD2_1 cd_l1_4 ( .a(in[7]), .abar(inbar[7]), .b(in[6]), .bbar(inbar[6]), .y(level1[15:12]), .ybar(level1bar[15:12]) );

  CD4_2 cd_l2_1 ( .a(level1[7:4]), .abar(level1bar[7:4]), .b(level1[3:0]), .bbar(level1bar[3:0]), 
        .y(level2[15:0]), .ybar(level2bar[15:0]) );
  CD4_1 cd_l2_2 ( .a(level1[15:12]), .abar(level1bar[15:12]), .b(level1[11:8]), .bbar(level1bar[11:8]), 
        .y(level2[31:16]), .ybar(level2bar[31:16]) );
  CD16_1 cd_l3 ( .a(level2[31:16]), .abar(level2bar[31:16]), .b(level2[15:0]), .bbar(level2bar[15:0]), 
        .y(out), .ybar(outbar) );
endmodule

module encode_1 ( in, inbar, out, outbar );

  input wire [255:0] in;
  input wire [255:0] inbar;
//input_done

  output wire [7:0] out;
  output wire [7:0] outbar;
//output_done

  wire in_81;
  wire in_80;
  wire in_79;
  wire in_78;
  wire in_77;
  wire in_76;
  wire in_75;
  wire in_74;
  wire in_73;
  wire in_72;
  wire in_71;
  wire in_70;
  wire in_69;
  wire in_68;
  wire in_67;
  wire in_66;
  wire in_65;
  wire in_64;
  wire in_63;
  wire in_62;
  wire in_61;
  wire in_60;
  wire in_59;
  wire in_58;
  wire in_57;
  wire in_56;
  wire in_55;
  wire in_54;
  wire in_53;
  wire in_52;
  wire in_51;
  wire in_50;
  wire in_49;
  wire in_48;
  wire in_47;
  wire in_46;
  wire in_45;
  wire in_44;
  wire in_43;
  wire in_42;
  wire in_41;
  wire in_40;
  wire in_39;
  wire in_38;
  wire in_37;
  wire in_36;
  wire in_35;
  wire in_34;
  wire in_33;
  wire in_32;
  wire in_31;
  wire in_30;
  wire in_29;
  wire in_28;
  wire in_27;
  wire in_26;
  wire in_25;
  wire in_24;
  wire in_23;
  wire in_22;
  wire in_21;
  wire in_20;
  wire in_19;
  wire in_18;
  wire in_17;
  wire in_16;
  wire in_15;
  wire in_14;
  wire in_13;
  wire in_12;
  wire in_11;
  wire in_10;
  wire in_9;
  wire in_8;
  wire in_7;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_3;
  wire in_2;
  wire in_1;
  wire in_0;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire in_81bar;
  wire in_80bar;
  wire in_79bar;
  wire in_78bar;
  wire in_77bar;
  wire in_76bar;
  wire in_75bar;
  wire in_74bar;
  wire in_73bar;
  wire in_72bar;
  wire in_71bar;
  wire in_70bar;
  wire in_69bar;
  wire in_68bar;
  wire in_67bar;
  wire in_66bar;
  wire in_65bar;
  wire in_64bar;
  wire in_63bar;
  wire in_62bar;
  wire in_61bar;
  wire in_60bar;
  wire in_59bar;
  wire in_58bar;
  wire in_57bar;
  wire in_56bar;
  wire in_55bar;
  wire in_54bar;
  wire in_53bar;
  wire in_52bar;
  wire in_51bar;
  wire in_50bar;
  wire in_49bar;
  wire in_48bar;
  wire in_47bar;
  wire in_46bar;
  wire in_45bar;
  wire in_44bar;
  wire in_43bar;
  wire in_42bar;
  wire in_41bar;
  wire in_40bar;
  wire in_39bar;
  wire in_38bar;
  wire in_37bar;
  wire in_36bar;
  wire in_35bar;
  wire in_34bar;
  wire in_33bar;
  wire in_32bar;
  wire in_31bar;
  wire in_30bar;
  wire in_29bar;
  wire in_28bar;
  wire in_27bar;
  wire in_26bar;
  wire in_25bar;
  wire in_24bar;
  wire in_23bar;
  wire in_22bar;
  wire in_21bar;
  wire in_20bar;
  wire in_19bar;
  wire in_18bar;
  wire in_17bar;
  wire in_16bar;
  wire in_15bar;
  wire in_14bar;
  wire in_13bar;
  wire in_12bar;
  wire in_11bar;
  wire in_10bar;
  wire in_9bar;
  wire in_8bar;
  wire in_7bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_3bar;
  wire in_2bar;
  wire in_1bar;
  wire in_0bar;
  wire n487bar;
  wire n488bar;
  wire n489bar;
  wire n490bar;
  wire n491bar;
  wire n492bar;
  wire n493bar;
  wire n494bar;
  wire n495bar;
  wire n496bar;
  wire n497bar;
  wire n498bar;
  wire n499bar;
  wire n500bar;
  wire n501bar;
  wire n502bar;
  wire n503bar;
  wire n504bar;
  wire n505bar;
  wire n506bar;
  wire n507bar;
  wire n508bar;
  wire n509bar;
  wire n510bar;
  wire n511bar;
  wire n512bar;
  wire n513bar;
  wire n514bar;
  wire n515bar;
  wire n516bar;
  wire n517bar;
  wire n518bar;
  wire n519bar;
  wire n520bar;
  wire n521bar;
  wire n522bar;
  wire n523bar;
  wire n524bar;
  wire n525bar;
  wire n526bar;
  wire n527bar;
  wire n528bar;
  wire n529bar;
  wire n530bar;
  wire n531bar;
  wire n532bar;
  wire n533bar;
  wire n534bar;
  wire n535bar;
  wire n536bar;
  wire n537bar;
  wire n538bar;
  wire n539bar;
  wire n540bar;
  wire n541bar;
  wire n542bar;
  wire n543bar;
  wire n544bar;
  wire n545bar;
  wire n546bar;
  wire n547bar;
  wire n548bar;
  wire n549bar;
  wire n550bar;
  wire n551bar;
  wire n552bar;
  wire n553bar;
  wire n554bar;
  wire n555bar;
  wire n556bar;
  wire n557bar;
  wire n558bar;
  wire n559bar;
  wire n560bar;
  wire n561bar;
  wire n562bar;
  wire n563bar;
  wire n564bar;
  wire n565bar;
  wire n566bar;
  wire n567bar;
  wire n568bar;
  wire n569bar;
  wire n570bar;
  wire n571bar;
  wire n572bar;
  wire n573bar;
  wire n574bar;
  wire n575bar;
  wire n576bar;
  wire n577bar;
  wire n578bar;
  wire n579bar;
  wire n580bar;
  wire n581bar;
  wire n582bar;
  wire n583bar;
  wire n584bar;
  wire n585bar;
  wire n586bar;
  wire n587bar;
  wire n588bar;
  wire n589bar;
  wire n590bar;
  wire n591bar;
  wire n592bar;
  wire n593bar;
  wire n594bar;
  wire n595bar;
  wire n596bar;
  wire n597bar;
  wire n598bar;
  wire n599bar;
  wire n600bar;
  wire n601bar;
  wire n602bar;
  wire n603bar;
  wire n604bar;
  wire n605bar;
  wire n606bar;
  wire n607bar;
  wire n608bar;
  wire n609bar;
  wire n610bar;
  wire n611bar;
  wire n612bar;
  wire n613bar;
  wire n614bar;
  wire n615bar;
  wire n616bar;
  wire n617bar;
  wire n618bar;
  wire n619bar;
  wire n620bar;
  wire n621bar;
  wire n622bar;
  wire n623bar;
  wire n624bar;
  wire n625bar;
  wire n626bar;
  wire n627bar;
  wire n628bar;
  wire n629bar;
  wire n630bar;
  wire n631bar;
  wire n632bar;
  wire n633bar;
  wire n634bar;
  wire n635bar;
  wire n636bar;
  wire n637bar;
  wire n638bar;
  wire n639bar;
  wire n640bar;
  wire n641bar;
  wire n642bar;
  wire n643bar;
  wire n644bar;
  wire n645bar;
  wire n646bar;
  wire n647bar;
  wire n648bar;
  wire n649bar;
  wire n650bar;
  wire n651bar;
  wire n652bar;
  wire n653bar;
  wire n654bar;
  wire n655bar;
  wire n656bar;
  wire n657bar;
  wire n658bar;
  wire n659bar;
  wire n660bar;
  wire n661bar;
  wire n662bar;
  wire n663bar;
  wire n664bar;
  wire n665bar;
  wire n666bar;
  wire n667bar;
  wire n668bar;
  wire n669bar;
  wire n670bar;
  wire n671bar;
  wire n672bar;
  wire n673bar;
  wire n674bar;
  wire n675bar;
  wire n676bar;
  wire n677bar;
  wire n678bar;
  wire n679bar;
  wire n680bar;
  wire n681bar;
  wire n682bar;
  wire n683bar;
  wire n684bar;
  wire n685bar;
  wire n686bar;
  wire n687bar;
  wire n688bar;
  wire n689bar;
  wire n690bar;
  wire n691bar;
  wire n692bar;
  wire n693bar;
  wire n694bar;
  wire n695bar;
  wire n696bar;
  wire n697bar;
  wire n698bar;
  wire n699bar;
  wire n700bar;
  wire n701bar;
  wire n702bar;
  wire n703bar;
  wire n704bar;
  wire n705bar;
  wire n706bar;
  wire n707bar;
  wire n708bar;
  wire n709bar;
  wire n710bar;
  wire n711bar;
  wire n712bar;
  wire n713bar;
  wire n714bar;
  wire n715bar;
  wire n716bar;
  wire n717bar;
  wire n718bar;
  wire n719bar;
  wire n720bar;
  wire n721bar;
  wire n722bar;
  wire n723bar;
  wire n724bar;
  wire n725bar;
  wire n726bar;
  wire n727bar;
  wire n728bar;
  wire n729bar;
  wire n730bar;
  wire n731bar;
  wire n732bar;
  wire n733bar;
  wire n734bar;
  wire n735bar;
  wire n736bar;
  wire n737bar;
  wire n738bar;
  wire n739bar;
  wire n740bar;
  wire n741bar;
  wire n742bar;
  wire n743bar;
  wire n744bar;
  wire n745bar;
  wire n746bar;
  wire n747bar;
  wire n748bar;
  wire n749bar;
  wire n750bar;
  wire n751bar;
  wire n752bar;
  wire n753bar;
  wire n754bar;
  wire n755bar;
  wire n756bar;
  wire n757bar;
  wire n758bar;
  wire n759bar;
  wire n760bar;
  wire n761bar;
  wire n762bar;
  wire n763bar;
  wire n764bar;
  wire n765bar;
  wire n766bar;
  wire n767bar;
  wire n768bar;
  wire n769bar;
  wire n770bar;
  wire n771bar;
  wire n772bar;
  wire n773bar;
  wire n774bar;
  wire n775bar;
  wire n776bar;
  wire n777bar;
  wire n778bar;
  wire n779bar;
  wire n780bar;
  wire n781bar;
  wire n782bar;
  wire n783bar;
  wire n784bar;
  wire n785bar;
  wire n786bar;
  wire n787bar;
  wire n788bar;
  wire n789bar;
  wire n790bar;
  wire n791bar;
  wire n792bar;
  wire n793bar;
  wire n794bar;
  wire n795bar;
  wire n796bar;
  wire n797bar;
  wire n798bar;
  wire n799bar;
  wire n800bar;
  wire n801bar;
  wire n802bar;
  wire n803bar;
  wire n804bar;
  wire n805bar;
  wire n806bar;
  wire n807bar;
  wire n808bar;
  wire n809bar;
  wire n810bar;
  wire n811bar;
  wire n812bar;
  wire n813bar;
  wire n814bar;
  wire n815bar;
  wire n816bar;
  wire n817bar;
  wire n818bar;
  wire n819bar;
  wire n820bar;
  wire n821bar;
  wire n822bar;
  wire n823bar;
  wire n824bar;
  wire n825bar;
  wire n826bar;
  wire n827bar;
  wire n828bar;
  wire n829bar;
  wire n830bar;
  wire n831bar;
  wire n832bar;
  wire n833bar;
  wire n834bar;
  wire n835bar;
  wire n836bar;
  wire n837bar;
  wire n838bar;
  wire n839bar;
  wire n840bar;
  wire n841bar;
  wire n842bar;
  wire n843bar;
  wire n844bar;
  wire n845bar;
  wire n846bar;
  wire n847bar;
  wire n848bar;
  wire n849bar;
  wire n850bar;
  wire n851bar;
  wire n852bar;
  wire n853bar;
  wire n854bar;
  wire n855bar;
  wire n856bar;
  wire n857bar;
  wire n858bar;
  wire n859bar;
  wire n860bar;
  wire n861bar;
  wire n862bar;
  wire n863bar;
  wire n864bar;
  wire n865bar;
  wire n866bar;
  wire n867bar;
  wire n868bar;
  wire n869bar;
  wire n870bar;
  wire n871bar;
  wire n872bar;
  wire n873bar;
  wire n874bar;
  wire n875bar;
  wire n876bar;
  wire n877bar;
  wire n878bar;
  wire n879bar;
  wire n880bar;
  wire n881bar;
  wire n882bar;
  wire n883bar;
  wire n884bar;
  wire n885bar;
  wire n886bar;
  wire n887bar;
  wire n888bar;
  wire n889bar;
  wire n890bar;
  wire n891bar;
  wire n892bar;
  wire n893bar;
  wire n894bar;
  wire n895bar;
  wire n896bar;
  wire n897bar;
  wire n898bar;
  wire n899bar;
  wire n900bar;
  wire n901bar;
  wire n902bar;
  wire n903bar;
  wire n904bar;
  wire n905bar;
  wire n906bar;
  wire n907bar;
  wire n908bar;
  wire n909bar;
  wire n910bar;
  wire n911bar;
  wire n912bar;
  wire n913bar;
  wire n914bar;
  wire n915bar;
  wire n916bar;
  wire n917bar;
  wire n918bar;
  wire n919bar;
  wire n920bar;
  wire n921bar;
  wire n922bar;
  wire n923bar;
  wire n924bar;
  wire n925bar;
  wire n926bar;
  wire n927bar;
  wire n928bar;
  wire n929bar;
  wire n930bar;
  wire n931bar;
  wire n932bar;
  wire n933bar;
  wire n934bar;
  wire n935bar;
  wire n936bar;
  wire n937bar;
  wire n938bar;
  wire n939bar;
  wire n940bar;
  wire n941bar;
  wire n942bar;
  wire n943bar;
  wire n944bar;
  wire n945bar;
  wire n946bar;
  wire n947bar;
  wire n948bar;
  wire n949bar;
  wire n950bar;
  wire n951bar;
  wire n952bar;
  wire n953bar;
  wire n954bar;
  wire n955bar;
  wire n956bar;
  wire n957bar;
  wire n958bar;
  wire n959bar;
  wire n960bar;
  wire n961bar;
  wire n962bar;
  wire n963bar;
  wire n964bar;
  wire n965bar;
  wire n966bar;
  wire n967bar;
  wire n968bar;
  wire n969bar;
  wire n970bar;
  wire n971bar;
  wire n972bar;
//wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];
  assign in_81bar = inbar[81];
  assign in_80bar = inbar[80];
  assign in_79bar = inbar[79];
  assign in_78bar = inbar[78];
  assign in_77bar = inbar[77];
  assign in_76bar = inbar[76];
  assign in_75bar = inbar[75];
  assign in_74bar = inbar[74];
  assign in_73bar = inbar[73];
  assign in_72bar = inbar[72];
  assign in_71bar = inbar[71];
  assign in_70bar = inbar[70];
  assign in_69bar = inbar[69];
  assign in_68bar = inbar[68];
  assign in_67bar = inbar[67];
  assign in_66bar = inbar[66];
  assign in_65bar = inbar[65];
  assign in_64bar = inbar[64];
  assign in_63bar = inbar[63];
  assign in_62bar = inbar[62];
  assign in_61bar = inbar[61];
  assign in_60bar = inbar[60];
  assign in_59bar = inbar[59];
  assign in_58bar = inbar[58];
  assign in_57bar = inbar[57];
  assign in_56bar = inbar[56];
  assign in_55bar = inbar[55];
  assign in_54bar = inbar[54];
  assign in_53bar = inbar[53];
  assign in_52bar = inbar[52];
  assign in_51bar = inbar[51];
  assign in_50bar = inbar[50];
  assign in_49bar = inbar[49];
  assign in_48bar = inbar[48];
  assign in_47bar = inbar[47];
  assign in_46bar = inbar[46];
  assign in_45bar = inbar[45];
  assign in_44bar = inbar[44];
  assign in_43bar = inbar[43];
  assign in_42bar = inbar[42];
  assign in_41bar = inbar[41];
  assign in_40bar = inbar[40];
  assign in_39bar = inbar[39];
  assign in_38bar = inbar[38];
  assign in_37bar = inbar[37];
  assign in_36bar = inbar[36];
  assign in_35bar = inbar[35];
  assign in_34bar = inbar[34];
  assign in_33bar = inbar[33];
  assign in_32bar = inbar[32];
  assign in_31bar = inbar[31];
  assign in_30bar = inbar[30];
  assign in_29bar = inbar[29];
  assign in_28bar = inbar[28];
  assign in_27bar = inbar[27];
  assign in_26bar = inbar[26];
  assign in_25bar = inbar[25];
  assign in_24bar = inbar[24];
  assign in_23bar = inbar[23];
  assign in_22bar = inbar[22];
  assign in_21bar = inbar[21];
  assign in_20bar = inbar[20];
  assign in_19bar = inbar[19];
  assign in_18bar = inbar[18];
  assign in_17bar = inbar[17];
  assign in_16bar = inbar[16];
  assign in_15bar = inbar[15];
  assign in_14bar = inbar[14];
  assign in_13bar = inbar[13];
  assign in_12bar = inbar[12];
  assign in_11bar = inbar[11];
  assign in_10bar = inbar[10];
  assign in_9bar = inbar[9];
  assign in_8bar = inbar[8];
  assign in_7bar = inbar[7];
  assign in_6bar = inbar[6];
  assign in_5bar = inbar[5];
  assign in_4bar = inbar[4];
  assign in_3bar = inbar[3];
  assign in_2bar = inbar[2];
  assign in_1bar = inbar[1];
  assign in_0bar = inbar[0];
//assign_done

  OR2_X1 U1 ( .A1(n972), .A2(n971), .ZN(out[7]) );
  AND2_X1 U1bar ( .A1(n972bar), .A2(n971bar), .ZN(outbar[7]) );
  OR2_X1 U2 ( .A1(n970), .A2(n969), .ZN(n971) );
  AND2_X1 U2bar ( .A1(n970bar), .A2(n969bar), .ZN(n971bar) );
  OR2_X1 U3 ( .A1(n968), .A2(n967), .ZN(n969) );
  AND2_X1 U3bar ( .A1(n968bar), .A2(n967bar), .ZN(n969bar) );
  OR2_X1 U4 ( .A1(n966), .A2(n965), .ZN(n967) );
  AND2_X1 U4bar ( .A1(n966bar), .A2(n965bar), .ZN(n967bar) );
  OR2_X1 U5 ( .A1(n964), .A2(n963), .ZN(n968) );
  AND2_X1 U5bar ( .A1(n964bar), .A2(n963bar), .ZN(n968bar) );
  OR2_X1 U6 ( .A1(in[116]), .A2(n962), .ZN(n963) );
  AND2_X1 U6bar ( .A1(inbar[116]), .A2(n962bar), .ZN(n963bar) );
  OR2_X1 U7 ( .A1(n961), .A2(n960), .ZN(n970) );
  AND2_X1 U7bar ( .A1(n961bar), .A2(n960bar), .ZN(n970bar) );
  OR2_X1 U8 ( .A1(in[150]), .A2(in[127]), .ZN(n960) );
  AND2_X1 U8bar ( .A1(inbar[150]), .A2(inbar[127]), .ZN(n960bar) );
  OR2_X1 U9 ( .A1(in[160]), .A2(n959), .ZN(n961) );
  AND2_X1 U9bar ( .A1(inbar[160]), .A2(n959bar), .ZN(n961bar) );
  OR2_X1 U10 ( .A1(in[252]), .A2(in[168]), .ZN(n959) );
  AND2_X1 U10bar ( .A1(inbar[252]), .A2(inbar[168]), .ZN(n959bar) );
  OR2_X1 U11 ( .A1(n958), .A2(n957), .ZN(n972) );
  AND2_X1 U11bar ( .A1(n958bar), .A2(n957bar), .ZN(n972bar) );
  OR2_X1 U12 ( .A1(n956), .A2(n955), .ZN(n957) );
  AND2_X1 U12bar ( .A1(n956bar), .A2(n955bar), .ZN(n957bar) );
  OR2_X1 U13 ( .A1(in_17), .A2(in[96]), .ZN(n955) );
  AND2_X1 U13bar ( .A1(in_17bar), .A2(inbar[96]), .ZN(n955bar) );
  OR2_X1 U14 ( .A1(in_23), .A2(n954), .ZN(n956) );
  AND2_X1 U14bar ( .A1(in_23bar), .A2(n954bar), .ZN(n956bar) );
  OR2_X1 U15 ( .A1(in_31), .A2(in_26), .ZN(n954) );
  AND2_X1 U15bar ( .A1(in_31bar), .A2(in_26bar), .ZN(n954bar) );
  OR2_X1 U16 ( .A1(n953), .A2(n952), .ZN(n958) );
  AND2_X1 U16bar ( .A1(n953bar), .A2(n952bar), .ZN(n958bar) );
  OR2_X1 U17 ( .A1(in_58), .A2(in_4), .ZN(n952) );
  AND2_X1 U17bar ( .A1(in_58bar), .A2(in_4bar), .ZN(n952bar) );
  OR2_X1 U18 ( .A1(in_59), .A2(n951), .ZN(n953) );
  AND2_X1 U18bar ( .A1(in_59bar), .A2(n951bar), .ZN(n953bar) );
  OR2_X1 U19 ( .A1(in_71), .A2(in_62), .ZN(n951) );
  AND2_X1 U19bar ( .A1(in_71bar), .A2(in_62bar), .ZN(n951bar) );
  OR2_X1 U20 ( .A1(n950), .A2(n949), .ZN(out[6]) );
  AND2_X1 U20bar ( .A1(n950bar), .A2(n949bar), .ZN(outbar[6]) );
  OR2_X1 U21 ( .A1(n948), .A2(n947), .ZN(n949) );
  AND2_X1 U21bar ( .A1(n948bar), .A2(n947bar), .ZN(n949bar) );
  OR2_X1 U22 ( .A1(n946), .A2(n945), .ZN(n947) );
  AND2_X1 U22bar ( .A1(n946bar), .A2(n945bar), .ZN(n947bar) );
  OR2_X1 U23 ( .A1(n944), .A2(n943), .ZN(n945) );
  AND2_X1 U23bar ( .A1(n944bar), .A2(n943bar), .ZN(n945bar) );
  OR2_X1 U24 ( .A1(n942), .A2(n941), .ZN(n946) );
  AND2_X1 U24bar ( .A1(n942bar), .A2(n941bar), .ZN(n946bar) );
  OR2_X1 U25 ( .A1(in[101]), .A2(n940), .ZN(n941) );
  AND2_X1 U25bar ( .A1(inbar[101]), .A2(n940bar), .ZN(n941bar) );
  OR2_X1 U26 ( .A1(n939), .A2(n938), .ZN(n948) );
  AND2_X1 U26bar ( .A1(n939bar), .A2(n938bar), .ZN(n948bar) );
  OR2_X1 U27 ( .A1(in[114]), .A2(in[104]), .ZN(n938) );
  AND2_X1 U27bar ( .A1(inbar[114]), .A2(inbar[104]), .ZN(n938bar) );
  OR2_X1 U28 ( .A1(in[128]), .A2(n937), .ZN(n939) );
  AND2_X1 U28bar ( .A1(inbar[128]), .A2(n937bar), .ZN(n939bar) );
  OR2_X1 U29 ( .A1(in[136]), .A2(in[134]), .ZN(n937) );
  AND2_X1 U29bar ( .A1(inbar[136]), .A2(inbar[134]), .ZN(n937bar) );
  OR2_X1 U30 ( .A1(n936), .A2(n935), .ZN(n950) );
  AND2_X1 U30bar ( .A1(n936bar), .A2(n935bar), .ZN(n950bar) );
  OR2_X1 U31 ( .A1(n934), .A2(n933), .ZN(n935) );
  AND2_X1 U31bar ( .A1(n934bar), .A2(n933bar), .ZN(n935bar) );
  OR2_X1 U32 ( .A1(in[177]), .A2(in[164]), .ZN(n933) );
  AND2_X1 U32bar ( .A1(inbar[177]), .A2(inbar[164]), .ZN(n933bar) );
  OR2_X1 U33 ( .A1(in[212]), .A2(n932), .ZN(n934) );
  AND2_X1 U33bar ( .A1(inbar[212]), .A2(n932bar), .ZN(n934bar) );
  OR2_X1 U34 ( .A1(in[248]), .A2(in[221]), .ZN(n932) );
  AND2_X1 U34bar ( .A1(inbar[248]), .A2(inbar[221]), .ZN(n932bar) );
  OR2_X1 U35 ( .A1(n931), .A2(n930), .ZN(n936) );
  AND2_X1 U35bar ( .A1(n931bar), .A2(n930bar), .ZN(n936bar) );
  OR2_X1 U36 ( .A1(in_18), .A2(in[93]), .ZN(n930) );
  AND2_X1 U36bar ( .A1(in_18bar), .A2(inbar[93]), .ZN(n930bar) );
  OR2_X1 U37 ( .A1(in_31), .A2(n929), .ZN(n931) );
  AND2_X1 U37bar ( .A1(in_31bar), .A2(n929bar), .ZN(n931bar) );
  OR2_X1 U38 ( .A1(in_7), .A2(in_39), .ZN(n929) );
  AND2_X1 U38bar ( .A1(in_7bar), .A2(in_39bar), .ZN(n929bar) );
  OR2_X1 U39 ( .A1(n928), .A2(n927), .ZN(out[5]) );
  AND2_X1 U39bar ( .A1(n928bar), .A2(n927bar), .ZN(outbar[5]) );
  OR2_X1 U40 ( .A1(n926), .A2(n925), .ZN(n927) );
  AND2_X1 U40bar ( .A1(n926bar), .A2(n925bar), .ZN(n927bar) );
  OR2_X1 U41 ( .A1(n924), .A2(n923), .ZN(n925) );
  AND2_X1 U41bar ( .A1(n924bar), .A2(n923bar), .ZN(n925bar) );
  OR2_X1 U42 ( .A1(n922), .A2(n921), .ZN(n923) );
  AND2_X1 U42bar ( .A1(n922bar), .A2(n921bar), .ZN(n923bar) );
  OR2_X1 U43 ( .A1(n940), .A2(n920), .ZN(n924) );
  AND2_X1 U43bar ( .A1(n940bar), .A2(n920bar), .ZN(n924bar) );
  OR2_X1 U44 ( .A1(in[111]), .A2(n919), .ZN(n920) );
  AND2_X1 U44bar ( .A1(inbar[111]), .A2(n919bar), .ZN(n920bar) );
  OR2_X1 U45 ( .A1(n918), .A2(n917), .ZN(n940) );
  AND2_X1 U45bar ( .A1(n918bar), .A2(n917bar), .ZN(n940bar) );
  OR2_X1 U46 ( .A1(n916), .A2(n915), .ZN(n917) );
  AND2_X1 U46bar ( .A1(n916bar), .A2(n915bar), .ZN(n917bar) );
  OR2_X1 U47 ( .A1(n914), .A2(n913), .ZN(n915) );
  AND2_X1 U47bar ( .A1(n914bar), .A2(n913bar), .ZN(n915bar) );
  OR2_X1 U48 ( .A1(in[140]), .A2(in[131]), .ZN(n913) );
  AND2_X1 U48bar ( .A1(inbar[140]), .A2(inbar[131]), .ZN(n913bar) );
  OR2_X1 U49 ( .A1(in[160]), .A2(in[144]), .ZN(n914) );
  AND2_X1 U49bar ( .A1(inbar[160]), .A2(inbar[144]), .ZN(n914bar) );
  OR2_X1 U50 ( .A1(n912), .A2(n911), .ZN(n916) );
  AND2_X1 U50bar ( .A1(n912bar), .A2(n911bar), .ZN(n916bar) );
  OR2_X1 U51 ( .A1(in[179]), .A2(in[174]), .ZN(n911) );
  AND2_X1 U51bar ( .A1(inbar[179]), .A2(inbar[174]), .ZN(n911bar) );
  OR2_X1 U52 ( .A1(in[188]), .A2(in[184]), .ZN(n912) );
  AND2_X1 U52bar ( .A1(inbar[188]), .A2(inbar[184]), .ZN(n912bar) );
  OR2_X1 U53 ( .A1(n910), .A2(n909), .ZN(n918) );
  AND2_X1 U53bar ( .A1(n910bar), .A2(n909bar), .ZN(n918bar) );
  OR2_X1 U54 ( .A1(n908), .A2(n907), .ZN(n909) );
  AND2_X1 U54bar ( .A1(n908bar), .A2(n907bar), .ZN(n909bar) );
  OR2_X1 U55 ( .A1(in[216]), .A2(in[200]), .ZN(n907) );
  AND2_X1 U55bar ( .A1(inbar[216]), .A2(inbar[200]), .ZN(n907bar) );
  OR2_X1 U56 ( .A1(in[228]), .A2(in[224]), .ZN(n908) );
  AND2_X1 U56bar ( .A1(inbar[228]), .A2(inbar[224]), .ZN(n908bar) );
  OR2_X1 U57 ( .A1(n906), .A2(n905), .ZN(n910) );
  AND2_X1 U57bar ( .A1(n906bar), .A2(n905bar), .ZN(n910bar) );
  OR2_X1 U58 ( .A1(in[247]), .A2(in[235]), .ZN(n905) );
  AND2_X1 U58bar ( .A1(inbar[247]), .A2(inbar[235]), .ZN(n905bar) );
  OR2_X1 U59 ( .A1(in_42), .A2(in[83]), .ZN(n906) );
  AND2_X1 U59bar ( .A1(in_42bar), .A2(inbar[83]), .ZN(n906bar) );
  OR2_X1 U60 ( .A1(n904), .A2(n903), .ZN(n926) );
  AND2_X1 U60bar ( .A1(n904bar), .A2(n903bar), .ZN(n926bar) );
  OR2_X1 U61 ( .A1(in[166]), .A2(in[123]), .ZN(n903) );
  AND2_X1 U61bar ( .A1(inbar[166]), .A2(inbar[123]), .ZN(n903bar) );
  OR2_X1 U62 ( .A1(in[170]), .A2(n902), .ZN(n904) );
  AND2_X1 U62bar ( .A1(inbar[170]), .A2(n902bar), .ZN(n904bar) );
  OR2_X1 U63 ( .A1(in[194]), .A2(in[183]), .ZN(n902) );
  AND2_X1 U63bar ( .A1(inbar[194]), .A2(inbar[183]), .ZN(n902bar) );
  OR2_X1 U64 ( .A1(n901), .A2(n900), .ZN(n928) );
  AND2_X1 U64bar ( .A1(n901bar), .A2(n900bar), .ZN(n928bar) );
  OR2_X1 U65 ( .A1(n899), .A2(n898), .ZN(n900) );
  AND2_X1 U65bar ( .A1(n899bar), .A2(n898bar), .ZN(n900bar) );
  OR2_X1 U66 ( .A1(in[241]), .A2(in[238]), .ZN(n898) );
  AND2_X1 U66bar ( .A1(inbar[241]), .A2(inbar[238]), .ZN(n898bar) );
  OR2_X1 U67 ( .A1(in[250]), .A2(n897), .ZN(n899) );
  AND2_X1 U67bar ( .A1(inbar[250]), .A2(n897bar), .ZN(n899bar) );
  OR2_X1 U68 ( .A1(in_24), .A2(in[84]), .ZN(n897) );
  AND2_X1 U68bar ( .A1(in_24bar), .A2(inbar[84]), .ZN(n897bar) );
  OR2_X1 U69 ( .A1(n896), .A2(n895), .ZN(n901) );
  AND2_X1 U69bar ( .A1(n896bar), .A2(n895bar), .ZN(n901bar) );
  OR2_X1 U70 ( .A1(in_41), .A2(in_29), .ZN(n895) );
  AND2_X1 U70bar ( .A1(in_41bar), .A2(in_29bar), .ZN(n895bar) );
  OR2_X1 U71 ( .A1(in_66), .A2(n894), .ZN(n896) );
  AND2_X1 U71bar ( .A1(in_66bar), .A2(n894bar), .ZN(n896bar) );
  OR2_X1 U72 ( .A1(in_76), .A2(in_71), .ZN(n894) );
  AND2_X1 U72bar ( .A1(in_76bar), .A2(in_71bar), .ZN(n894bar) );
  OR2_X1 U73 ( .A1(n893), .A2(n892), .ZN(out[4]) );
  AND2_X1 U73bar ( .A1(n893bar), .A2(n892bar), .ZN(outbar[4]) );
  OR2_X1 U74 ( .A1(n891), .A2(n890), .ZN(n892) );
  AND2_X1 U74bar ( .A1(n891bar), .A2(n890bar), .ZN(n892bar) );
  OR2_X1 U75 ( .A1(n889), .A2(n888), .ZN(n890) );
  AND2_X1 U75bar ( .A1(n889bar), .A2(n888bar), .ZN(n890bar) );
  OR2_X1 U76 ( .A1(n922), .A2(n887), .ZN(n888) );
  AND2_X1 U76bar ( .A1(n922bar), .A2(n887bar), .ZN(n888bar) );
  OR2_X1 U77 ( .A1(n886), .A2(n885), .ZN(n922) );
  AND2_X1 U77bar ( .A1(n886bar), .A2(n885bar), .ZN(n922bar) );
  OR2_X1 U78 ( .A1(n884), .A2(n883), .ZN(n885) );
  AND2_X1 U78bar ( .A1(n884bar), .A2(n883bar), .ZN(n885bar) );
  OR2_X1 U79 ( .A1(n882), .A2(n881), .ZN(n883) );
  AND2_X1 U79bar ( .A1(n882bar), .A2(n881bar), .ZN(n883bar) );
  OR2_X1 U80 ( .A1(in[118]), .A2(in[109]), .ZN(n881) );
  AND2_X1 U80bar ( .A1(inbar[118]), .A2(inbar[109]), .ZN(n881bar) );
  OR2_X1 U81 ( .A1(in[139]), .A2(in[120]), .ZN(n882) );
  AND2_X1 U81bar ( .A1(inbar[139]), .A2(inbar[120]), .ZN(n882bar) );
  OR2_X1 U82 ( .A1(n880), .A2(n879), .ZN(n884) );
  AND2_X1 U82bar ( .A1(n880bar), .A2(n879bar), .ZN(n884bar) );
  OR2_X1 U83 ( .A1(in[198]), .A2(in[154]), .ZN(n879) );
  AND2_X1 U83bar ( .A1(inbar[198]), .A2(inbar[154]), .ZN(n879bar) );
  OR2_X1 U84 ( .A1(in[210]), .A2(in[205]), .ZN(n880) );
  AND2_X1 U84bar ( .A1(inbar[210]), .A2(inbar[205]), .ZN(n880bar) );
  OR2_X1 U85 ( .A1(n878), .A2(n877), .ZN(n886) );
  AND2_X1 U85bar ( .A1(n878bar), .A2(n877bar), .ZN(n886bar) );
  OR2_X1 U86 ( .A1(n876), .A2(n875), .ZN(n877) );
  AND2_X1 U86bar ( .A1(n876bar), .A2(n875bar), .ZN(n877bar) );
  OR2_X1 U87 ( .A1(in[219]), .A2(in[217]), .ZN(n875) );
  AND2_X1 U87bar ( .A1(inbar[219]), .A2(inbar[217]), .ZN(n875bar) );
  OR2_X1 U88 ( .A1(in[86]), .A2(in[252]), .ZN(n876) );
  AND2_X1 U88bar ( .A1(inbar[86]), .A2(inbar[252]), .ZN(n876bar) );
  OR2_X1 U89 ( .A1(n874), .A2(n873), .ZN(n878) );
  AND2_X1 U89bar ( .A1(n874bar), .A2(n873bar), .ZN(n878bar) );
  OR2_X1 U90 ( .A1(in_40), .A2(in[91]), .ZN(n873) );
  AND2_X1 U90bar ( .A1(in_40bar), .A2(inbar[91]), .ZN(n873bar) );
  OR2_X1 U91 ( .A1(in_8), .A2(in_46), .ZN(n874) );
  AND2_X1 U91bar ( .A1(in_8bar), .A2(in_46bar), .ZN(n874bar) );
  OR2_X1 U92 ( .A1(n872), .A2(n871), .ZN(n889) );
  AND2_X1 U92bar ( .A1(n872bar), .A2(n871bar), .ZN(n889bar) );
  OR2_X1 U93 ( .A1(in[117]), .A2(n943), .ZN(n871) );
  AND2_X1 U93bar ( .A1(inbar[117]), .A2(n943bar), .ZN(n871bar) );
  OR2_X1 U94 ( .A1(n870), .A2(n869), .ZN(n943) );
  AND2_X1 U94bar ( .A1(n870bar), .A2(n869bar), .ZN(n943bar) );
  OR2_X1 U95 ( .A1(n868), .A2(n867), .ZN(n869) );
  AND2_X1 U95bar ( .A1(n868bar), .A2(n867bar), .ZN(n869bar) );
  OR2_X1 U96 ( .A1(n866), .A2(n865), .ZN(n867) );
  AND2_X1 U96bar ( .A1(n866bar), .A2(n865bar), .ZN(n867bar) );
  OR2_X1 U97 ( .A1(n864), .A2(n863), .ZN(n865) );
  AND2_X1 U97bar ( .A1(n864bar), .A2(n863bar), .ZN(n865bar) );
  OR2_X1 U98 ( .A1(in[108]), .A2(n919), .ZN(n866) );
  AND2_X1 U98bar ( .A1(inbar[108]), .A2(n919bar), .ZN(n866bar) );
  OR2_X1 U99 ( .A1(n862), .A2(n861), .ZN(n919) );
  AND2_X1 U99bar ( .A1(n862bar), .A2(n861bar), .ZN(n919bar) );
  OR2_X1 U100 ( .A1(n860), .A2(n859), .ZN(n861) );
  AND2_X1 U100bar ( .A1(n860bar), .A2(n859bar), .ZN(n861bar) );
  OR2_X1 U101 ( .A1(n858), .A2(n857), .ZN(n859) );
  AND2_X1 U101bar ( .A1(n858bar), .A2(n857bar), .ZN(n859bar) );
  OR2_X1 U102 ( .A1(in[119]), .A2(in[105]), .ZN(n857) );
  AND2_X1 U102bar ( .A1(inbar[119]), .A2(inbar[105]), .ZN(n857bar) );
  OR2_X1 U103 ( .A1(in[186]), .A2(in[175]), .ZN(n858) );
  AND2_X1 U103bar ( .A1(inbar[186]), .A2(inbar[175]), .ZN(n858bar) );
  OR2_X1 U104 ( .A1(n856), .A2(n855), .ZN(n860) );
  AND2_X1 U104bar ( .A1(n856bar), .A2(n855bar), .ZN(n860bar) );
  OR2_X1 U105 ( .A1(in[202]), .A2(in[193]), .ZN(n855) );
  AND2_X1 U105bar ( .A1(inbar[202]), .A2(inbar[193]), .ZN(n855bar) );
  OR2_X1 U106 ( .A1(in[225]), .A2(in[208]), .ZN(n856) );
  AND2_X1 U106bar ( .A1(inbar[225]), .A2(inbar[208]), .ZN(n856bar) );
  OR2_X1 U107 ( .A1(n854), .A2(n853), .ZN(n862) );
  AND2_X1 U107bar ( .A1(n854bar), .A2(n853bar), .ZN(n862bar) );
  OR2_X1 U108 ( .A1(n852), .A2(n851), .ZN(n853) );
  AND2_X1 U108bar ( .A1(n852bar), .A2(n851bar), .ZN(n853bar) );
  OR2_X1 U109 ( .A1(in_1), .A2(in[85]), .ZN(n851) );
  AND2_X1 U109bar ( .A1(in_1bar), .A2(inbar[85]), .ZN(n851bar) );
  OR2_X1 U110 ( .A1(in_23), .A2(in_19), .ZN(n852) );
  AND2_X1 U110bar ( .A1(in_23bar), .A2(in_19bar), .ZN(n852bar) );
  OR2_X1 U111 ( .A1(n850), .A2(n849), .ZN(n854) );
  AND2_X1 U111bar ( .A1(n850bar), .A2(n849bar), .ZN(n854bar) );
  OR2_X1 U112 ( .A1(in_43), .A2(in_33), .ZN(n849) );
  AND2_X1 U112bar ( .A1(in_43bar), .A2(in_33bar), .ZN(n849bar) );
  OR2_X1 U113 ( .A1(in_63), .A2(in_44), .ZN(n850) );
  AND2_X1 U113bar ( .A1(in_63bar), .A2(in_44bar), .ZN(n850bar) );
  OR2_X1 U114 ( .A1(n848), .A2(n847), .ZN(n868) );
  AND2_X1 U114bar ( .A1(n848bar), .A2(n847bar), .ZN(n868bar) );
  OR2_X1 U115 ( .A1(in[141]), .A2(in[112]), .ZN(n847) );
  AND2_X1 U115bar ( .A1(inbar[141]), .A2(inbar[112]), .ZN(n847bar) );
  OR2_X1 U116 ( .A1(in[147]), .A2(n846), .ZN(n848) );
  AND2_X1 U116bar ( .A1(inbar[147]), .A2(n846bar), .ZN(n848bar) );
  OR2_X1 U117 ( .A1(in[181]), .A2(in[167]), .ZN(n846) );
  AND2_X1 U117bar ( .A1(inbar[181]), .A2(inbar[167]), .ZN(n846bar) );
  OR2_X1 U118 ( .A1(n845), .A2(n844), .ZN(n870) );
  AND2_X1 U118bar ( .A1(n845bar), .A2(n844bar), .ZN(n870bar) );
  OR2_X1 U119 ( .A1(n843), .A2(n842), .ZN(n844) );
  AND2_X1 U119bar ( .A1(n843bar), .A2(n842bar), .ZN(n844bar) );
  OR2_X1 U120 ( .A1(in[229]), .A2(in[201]), .ZN(n842) );
  AND2_X1 U120bar ( .A1(inbar[229]), .A2(inbar[201]), .ZN(n842bar) );
  OR2_X1 U121 ( .A1(in[237]), .A2(n841), .ZN(n843) );
  AND2_X1 U121bar ( .A1(inbar[237]), .A2(n841bar), .ZN(n843bar) );
  OR2_X1 U122 ( .A1(in[94]), .A2(in[253]), .ZN(n841) );
  AND2_X1 U122bar ( .A1(inbar[94]), .A2(inbar[253]), .ZN(n841bar) );
  OR2_X1 U123 ( .A1(n840), .A2(n839), .ZN(n845) );
  AND2_X1 U123bar ( .A1(n840bar), .A2(n839bar), .ZN(n845bar) );
  OR2_X1 U124 ( .A1(in_21), .A2(in[96]), .ZN(n839) );
  AND2_X1 U124bar ( .A1(in_21bar), .A2(inbar[96]), .ZN(n839bar) );
  OR2_X1 U125 ( .A1(in_25), .A2(n838), .ZN(n840) );
  AND2_X1 U125bar ( .A1(in_25bar), .A2(n838bar), .ZN(n840bar) );
  OR2_X1 U126 ( .A1(in_81), .A2(in_45), .ZN(n838) );
  AND2_X1 U126bar ( .A1(in_81bar), .A2(in_45bar), .ZN(n838bar) );
  OR2_X1 U127 ( .A1(n837), .A2(n836), .ZN(n891) );
  AND2_X1 U127bar ( .A1(n837bar), .A2(n836bar), .ZN(n891bar) );
  OR2_X1 U128 ( .A1(in[142]), .A2(in[124]), .ZN(n836) );
  AND2_X1 U128bar ( .A1(inbar[142]), .A2(inbar[124]), .ZN(n836bar) );
  OR2_X1 U129 ( .A1(in[150]), .A2(n835), .ZN(n837) );
  AND2_X1 U129bar ( .A1(inbar[150]), .A2(n835bar), .ZN(n837bar) );
  OR2_X1 U130 ( .A1(in[172]), .A2(in[155]), .ZN(n835) );
  AND2_X1 U130bar ( .A1(inbar[172]), .A2(inbar[155]), .ZN(n835bar) );
  OR2_X1 U131 ( .A1(n834), .A2(n833), .ZN(n893) );
  AND2_X1 U131bar ( .A1(n834bar), .A2(n833bar), .ZN(n893bar) );
  OR2_X1 U132 ( .A1(n832), .A2(n831), .ZN(n833) );
  AND2_X1 U132bar ( .A1(n832bar), .A2(n831bar), .ZN(n833bar) );
  OR2_X1 U133 ( .A1(in[196]), .A2(in[173]), .ZN(n831) );
  AND2_X1 U133bar ( .A1(inbar[196]), .A2(inbar[173]), .ZN(n831bar) );
  OR2_X1 U134 ( .A1(in[222]), .A2(n830), .ZN(n832) );
  AND2_X1 U134bar ( .A1(inbar[222]), .A2(n830bar), .ZN(n832bar) );
  OR2_X1 U135 ( .A1(in[227]), .A2(in[226]), .ZN(n830) );
  AND2_X1 U135bar ( .A1(inbar[227]), .A2(inbar[226]), .ZN(n830bar) );
  OR2_X1 U136 ( .A1(n829), .A2(n828), .ZN(n834) );
  AND2_X1 U136bar ( .A1(n829bar), .A2(n828bar), .ZN(n834bar) );
  OR2_X1 U137 ( .A1(in[249]), .A2(in[231]), .ZN(n828) );
  AND2_X1 U137bar ( .A1(inbar[249]), .A2(inbar[231]), .ZN(n828bar) );
  OR2_X1 U138 ( .A1(in_28), .A2(n827), .ZN(n829) );
  AND2_X1 U138bar ( .A1(in_28bar), .A2(n827bar), .ZN(n829bar) );
  OR2_X1 U139 ( .A1(in_52), .A2(in_47), .ZN(n827) );
  AND2_X1 U139bar ( .A1(in_52bar), .A2(in_47bar), .ZN(n827bar) );
  OR2_X1 U140 ( .A1(n826), .A2(n825), .ZN(out[3]) );
  AND2_X1 U140bar ( .A1(n826bar), .A2(n825bar), .ZN(outbar[3]) );
  OR2_X1 U141 ( .A1(n824), .A2(n823), .ZN(n825) );
  AND2_X1 U141bar ( .A1(n824bar), .A2(n823bar), .ZN(n825bar) );
  OR2_X1 U142 ( .A1(n822), .A2(n821), .ZN(n823) );
  AND2_X1 U142bar ( .A1(n822bar), .A2(n821bar), .ZN(n823bar) );
  OR2_X1 U143 ( .A1(n820), .A2(n819), .ZN(n821) );
  AND2_X1 U143bar ( .A1(n820bar), .A2(n819bar), .ZN(n821bar) );
  OR2_X1 U144 ( .A1(n964), .A2(n818), .ZN(n822) );
  AND2_X1 U144bar ( .A1(n964bar), .A2(n818bar), .ZN(n822bar) );
  OR2_X1 U145 ( .A1(in[118]), .A2(n817), .ZN(n818) );
  AND2_X1 U145bar ( .A1(inbar[118]), .A2(n817bar), .ZN(n818bar) );
  OR2_X1 U146 ( .A1(n816), .A2(n815), .ZN(n964) );
  AND2_X1 U146bar ( .A1(n816bar), .A2(n815bar), .ZN(n964bar) );
  OR2_X1 U147 ( .A1(n814), .A2(n813), .ZN(n815) );
  AND2_X1 U147bar ( .A1(n814bar), .A2(n813bar), .ZN(n815bar) );
  OR2_X1 U148 ( .A1(n812), .A2(n811), .ZN(n813) );
  AND2_X1 U148bar ( .A1(n812bar), .A2(n811bar), .ZN(n813bar) );
  OR2_X1 U149 ( .A1(in[122]), .A2(in[111]), .ZN(n811) );
  AND2_X1 U149bar ( .A1(inbar[122]), .A2(inbar[111]), .ZN(n811bar) );
  OR2_X1 U150 ( .A1(in[154]), .A2(in[151]), .ZN(n812) );
  AND2_X1 U150bar ( .A1(inbar[154]), .A2(inbar[151]), .ZN(n812bar) );
  OR2_X1 U151 ( .A1(n810), .A2(n809), .ZN(n814) );
  AND2_X1 U151bar ( .A1(n810bar), .A2(n809bar), .ZN(n814bar) );
  OR2_X1 U152 ( .A1(in[187]), .A2(in[177]), .ZN(n809) );
  AND2_X1 U152bar ( .A1(inbar[187]), .A2(inbar[177]), .ZN(n809bar) );
  OR2_X1 U153 ( .A1(in[200]), .A2(in[192]), .ZN(n810) );
  AND2_X1 U153bar ( .A1(inbar[200]), .A2(inbar[192]), .ZN(n810bar) );
  OR2_X1 U154 ( .A1(n808), .A2(n807), .ZN(n816) );
  AND2_X1 U154bar ( .A1(n808bar), .A2(n807bar), .ZN(n816bar) );
  OR2_X1 U155 ( .A1(n806), .A2(n805), .ZN(n807) );
  AND2_X1 U155bar ( .A1(n806bar), .A2(n805bar), .ZN(n807bar) );
  OR2_X1 U156 ( .A1(in[225]), .A2(in[207]), .ZN(n805) );
  AND2_X1 U156bar ( .A1(inbar[225]), .A2(inbar[207]), .ZN(n805bar) );
  OR2_X1 U157 ( .A1(in[98]), .A2(in[226]), .ZN(n806) );
  AND2_X1 U157bar ( .A1(inbar[98]), .A2(inbar[226]), .ZN(n806bar) );
  OR2_X1 U158 ( .A1(n804), .A2(n803), .ZN(n808) );
  AND2_X1 U158bar ( .A1(n804bar), .A2(n803bar), .ZN(n808bar) );
  OR2_X1 U159 ( .A1(in_20), .A2(in_16), .ZN(n803) );
  AND2_X1 U159bar ( .A1(in_20bar), .A2(in_16bar), .ZN(n803bar) );
  OR2_X1 U160 ( .A1(in_55), .A2(in_45), .ZN(n804) );
  AND2_X1 U160bar ( .A1(in_55bar), .A2(in_45bar), .ZN(n804bar) );
  OR2_X1 U161 ( .A1(n802), .A2(n801), .ZN(n824) );
  AND2_X1 U161bar ( .A1(n802bar), .A2(n801bar), .ZN(n824bar) );
  OR2_X1 U162 ( .A1(in[162]), .A2(in[149]), .ZN(n801) );
  AND2_X1 U162bar ( .A1(inbar[162]), .A2(inbar[149]), .ZN(n801bar) );
  OR2_X1 U163 ( .A1(in[163]), .A2(n800), .ZN(n802) );
  AND2_X1 U163bar ( .A1(inbar[163]), .A2(n800bar), .ZN(n802bar) );
  OR2_X1 U164 ( .A1(in[191]), .A2(in[189]), .ZN(n800) );
  AND2_X1 U164bar ( .A1(inbar[191]), .A2(inbar[189]), .ZN(n800bar) );
  OR2_X1 U165 ( .A1(n799), .A2(n798), .ZN(n826) );
  AND2_X1 U165bar ( .A1(n799bar), .A2(n798bar), .ZN(n826bar) );
  OR2_X1 U166 ( .A1(n797), .A2(n796), .ZN(n798) );
  AND2_X1 U166bar ( .A1(n797bar), .A2(n796bar), .ZN(n798bar) );
  OR2_X1 U167 ( .A1(in[212]), .A2(in[193]), .ZN(n796) );
  AND2_X1 U167bar ( .A1(inbar[212]), .A2(inbar[193]), .ZN(n796bar) );
  OR2_X1 U168 ( .A1(in[238]), .A2(n795), .ZN(n797) );
  AND2_X1 U168bar ( .A1(inbar[238]), .A2(n795bar), .ZN(n797bar) );
  OR2_X1 U169 ( .A1(in[88]), .A2(in[247]), .ZN(n795) );
  AND2_X1 U169bar ( .A1(inbar[88]), .A2(inbar[247]), .ZN(n795bar) );
  OR2_X1 U170 ( .A1(n794), .A2(n793), .ZN(n799) );
  AND2_X1 U170bar ( .A1(n794bar), .A2(n793bar), .ZN(n799bar) );
  OR2_X1 U171 ( .A1(in[94]), .A2(in[92]), .ZN(n793) );
  AND2_X1 U171bar ( .A1(inbar[94]), .A2(inbar[92]), .ZN(n793bar) );
  OR2_X1 U172 ( .A1(in_52), .A2(n792), .ZN(n794) );
  AND2_X1 U172bar ( .A1(in_52bar), .A2(n792bar), .ZN(n794bar) );
  OR2_X1 U173 ( .A1(in_70), .A2(in_67), .ZN(n792) );
  AND2_X1 U173bar ( .A1(in_70bar), .A2(in_67bar), .ZN(n792bar) );
  OR2_X1 U174 ( .A1(n791), .A2(n790), .ZN(out[2]) );
  AND2_X1 U174bar ( .A1(n791bar), .A2(n790bar), .ZN(outbar[2]) );
  OR2_X1 U175 ( .A1(n789), .A2(n788), .ZN(n790) );
  AND2_X1 U175bar ( .A1(n789bar), .A2(n788bar), .ZN(n790bar) );
  OR2_X1 U176 ( .A1(n787), .A2(n786), .ZN(n788) );
  AND2_X1 U176bar ( .A1(n787bar), .A2(n786bar), .ZN(n788bar) );
  OR2_X1 U177 ( .A1(n819), .A2(n785), .ZN(n786) );
  AND2_X1 U177bar ( .A1(n819bar), .A2(n785bar), .ZN(n786bar) );
  OR2_X1 U178 ( .A1(n784), .A2(n783), .ZN(n819) );
  AND2_X1 U178bar ( .A1(n784bar), .A2(n783bar), .ZN(n819bar) );
  OR2_X1 U179 ( .A1(n782), .A2(n781), .ZN(n783) );
  AND2_X1 U179bar ( .A1(n782bar), .A2(n781bar), .ZN(n783bar) );
  OR2_X1 U180 ( .A1(n780), .A2(n779), .ZN(n781) );
  AND2_X1 U180bar ( .A1(n780bar), .A2(n779bar), .ZN(n781bar) );
  OR2_X1 U181 ( .A1(n962), .A2(n778), .ZN(n779) );
  AND2_X1 U181bar ( .A1(n962bar), .A2(n778bar), .ZN(n779bar) );
  OR2_X1 U182 ( .A1(n777), .A2(n776), .ZN(n962) );
  AND2_X1 U182bar ( .A1(n777bar), .A2(n776bar), .ZN(n962bar) );
  OR2_X1 U183 ( .A1(n775), .A2(n774), .ZN(n776) );
  AND2_X1 U183bar ( .A1(n775bar), .A2(n774bar), .ZN(n776bar) );
  OR2_X1 U184 ( .A1(n773), .A2(n772), .ZN(n774) );
  AND2_X1 U184bar ( .A1(n773bar), .A2(n772bar), .ZN(n774bar) );
  OR2_X1 U185 ( .A1(in[131]), .A2(in[120]), .ZN(n772) );
  AND2_X1 U185bar ( .A1(inbar[131]), .A2(inbar[120]), .ZN(n772bar) );
  OR2_X1 U186 ( .A1(in[153]), .A2(in[147]), .ZN(n773) );
  AND2_X1 U186bar ( .A1(inbar[153]), .A2(inbar[147]), .ZN(n773bar) );
  OR2_X1 U187 ( .A1(n771), .A2(n770), .ZN(n775) );
  AND2_X1 U187bar ( .A1(n771bar), .A2(n770bar), .ZN(n775bar) );
  OR2_X1 U188 ( .A1(in[170]), .A2(in[156]), .ZN(n770) );
  AND2_X1 U188bar ( .A1(inbar[170]), .A2(inbar[156]), .ZN(n770bar) );
  OR2_X1 U189 ( .A1(in[223]), .A2(in[190]), .ZN(n771) );
  AND2_X1 U189bar ( .A1(inbar[223]), .A2(inbar[190]), .ZN(n771bar) );
  OR2_X1 U190 ( .A1(n769), .A2(n768), .ZN(n777) );
  AND2_X1 U190bar ( .A1(n769bar), .A2(n768bar), .ZN(n777bar) );
  OR2_X1 U191 ( .A1(n767), .A2(n766), .ZN(n768) );
  AND2_X1 U191bar ( .A1(n767bar), .A2(n766bar), .ZN(n768bar) );
  OR2_X1 U192 ( .A1(in[236]), .A2(in[230]), .ZN(n766) );
  AND2_X1 U192bar ( .A1(inbar[236]), .A2(inbar[230]), .ZN(n766bar) );
  OR2_X1 U193 ( .A1(in[85]), .A2(in[240]), .ZN(n767) );
  AND2_X1 U193bar ( .A1(inbar[85]), .A2(inbar[240]), .ZN(n767bar) );
  OR2_X1 U194 ( .A1(n765), .A2(n764), .ZN(n769) );
  AND2_X1 U194bar ( .A1(n765bar), .A2(n764bar), .ZN(n769bar) );
  OR2_X1 U195 ( .A1(in_12), .A2(in[90]), .ZN(n764) );
  AND2_X1 U195bar ( .A1(in_12bar), .A2(inbar[90]), .ZN(n764bar) );
  OR2_X1 U196 ( .A1(in_39), .A2(in_28), .ZN(n765) );
  AND2_X1 U196bar ( .A1(in_39bar), .A2(in_28bar), .ZN(n765bar) );
  OR2_X1 U197 ( .A1(in[109]), .A2(n763), .ZN(n780) );
  AND2_X1 U197bar ( .A1(inbar[109]), .A2(n763bar), .ZN(n780bar) );
  OR2_X1 U198 ( .A1(n762), .A2(n761), .ZN(n782) );
  AND2_X1 U198bar ( .A1(n762bar), .A2(n761bar), .ZN(n782bar) );
  OR2_X1 U199 ( .A1(in[138]), .A2(in[129]), .ZN(n761) );
  AND2_X1 U199bar ( .A1(inbar[138]), .A2(inbar[129]), .ZN(n761bar) );
  OR2_X1 U200 ( .A1(in[157]), .A2(n760), .ZN(n762) );
  AND2_X1 U200bar ( .A1(inbar[157]), .A2(n760bar), .ZN(n762bar) );
  OR2_X1 U201 ( .A1(in[182]), .A2(in[167]), .ZN(n760) );
  AND2_X1 U201bar ( .A1(inbar[182]), .A2(inbar[167]), .ZN(n760bar) );
  OR2_X1 U202 ( .A1(n759), .A2(n758), .ZN(n784) );
  AND2_X1 U202bar ( .A1(n759bar), .A2(n758bar), .ZN(n784bar) );
  OR2_X1 U203 ( .A1(n757), .A2(n756), .ZN(n758) );
  AND2_X1 U203bar ( .A1(n757bar), .A2(n756bar), .ZN(n758bar) );
  OR2_X1 U204 ( .A1(in[195]), .A2(in[184]), .ZN(n756) );
  AND2_X1 U204bar ( .A1(inbar[195]), .A2(inbar[184]), .ZN(n756bar) );
  OR2_X1 U205 ( .A1(in[196]), .A2(n755), .ZN(n757) );
  AND2_X1 U205bar ( .A1(inbar[196]), .A2(n755bar), .ZN(n757bar) );
  OR2_X1 U206 ( .A1(in[215]), .A2(in[209]), .ZN(n755) );
  AND2_X1 U206bar ( .A1(inbar[215]), .A2(inbar[209]), .ZN(n755bar) );
  OR2_X1 U207 ( .A1(n754), .A2(n753), .ZN(n759) );
  AND2_X1 U207bar ( .A1(n754bar), .A2(n753bar), .ZN(n759bar) );
  OR2_X1 U208 ( .A1(in[93]), .A2(in[233]), .ZN(n753) );
  AND2_X1 U208bar ( .A1(inbar[93]), .A2(inbar[233]), .ZN(n753bar) );
  OR2_X1 U209 ( .A1(in_1), .A2(n752), .ZN(n754) );
  AND2_X1 U209bar ( .A1(in_1bar), .A2(n752bar), .ZN(n754bar) );
  OR2_X1 U210 ( .A1(in_69), .A2(in_66), .ZN(n752) );
  AND2_X1 U210bar ( .A1(in_69bar), .A2(in_66bar), .ZN(n752bar) );
  OR2_X1 U211 ( .A1(n966), .A2(n751), .ZN(n787) );
  AND2_X1 U211bar ( .A1(n966bar), .A2(n751bar), .ZN(n787bar) );
  OR2_X1 U212 ( .A1(in[134]), .A2(n750), .ZN(n751) );
  AND2_X1 U212bar ( .A1(inbar[134]), .A2(n750bar), .ZN(n751bar) );
  OR2_X1 U213 ( .A1(n749), .A2(n748), .ZN(n966) );
  AND2_X1 U213bar ( .A1(n749bar), .A2(n748bar), .ZN(n966bar) );
  OR2_X1 U214 ( .A1(n747), .A2(n746), .ZN(n748) );
  AND2_X1 U214bar ( .A1(n747bar), .A2(n746bar), .ZN(n748bar) );
  OR2_X1 U215 ( .A1(n745), .A2(n744), .ZN(n746) );
  AND2_X1 U215bar ( .A1(n745bar), .A2(n744bar), .ZN(n746bar) );
  OR2_X1 U216 ( .A1(in[136]), .A2(in[121]), .ZN(n744) );
  AND2_X1 U216bar ( .A1(inbar[136]), .A2(inbar[121]), .ZN(n744bar) );
  OR2_X1 U217 ( .A1(in[186]), .A2(in[174]), .ZN(n745) );
  AND2_X1 U217bar ( .A1(inbar[186]), .A2(inbar[174]), .ZN(n745bar) );
  OR2_X1 U218 ( .A1(n743), .A2(n742), .ZN(n747) );
  AND2_X1 U218bar ( .A1(n743bar), .A2(n742bar), .ZN(n747bar) );
  OR2_X1 U219 ( .A1(in[198]), .A2(in[197]), .ZN(n742) );
  AND2_X1 U219bar ( .A1(inbar[198]), .A2(inbar[197]), .ZN(n742bar) );
  OR2_X1 U220 ( .A1(in[214]), .A2(in[199]), .ZN(n743) );
  AND2_X1 U220bar ( .A1(inbar[214]), .A2(inbar[199]), .ZN(n743bar) );
  OR2_X1 U221 ( .A1(n741), .A2(n740), .ZN(n749) );
  AND2_X1 U221bar ( .A1(n741bar), .A2(n740bar), .ZN(n749bar) );
  OR2_X1 U222 ( .A1(n739), .A2(n738), .ZN(n740) );
  AND2_X1 U222bar ( .A1(n739bar), .A2(n738bar), .ZN(n740bar) );
  OR2_X1 U223 ( .A1(in[231]), .A2(in[220]), .ZN(n738) );
  AND2_X1 U223bar ( .A1(inbar[231]), .A2(inbar[220]), .ZN(n738bar) );
  OR2_X1 U224 ( .A1(in_25), .A2(in[245]), .ZN(n739) );
  AND2_X1 U224bar ( .A1(in_25bar), .A2(inbar[245]), .ZN(n739bar) );
  OR2_X1 U225 ( .A1(n737), .A2(n736), .ZN(n741) );
  AND2_X1 U225bar ( .A1(n737bar), .A2(n736bar), .ZN(n741bar) );
  OR2_X1 U226 ( .A1(in_53), .A2(in_29), .ZN(n736) );
  AND2_X1 U226bar ( .A1(in_53bar), .A2(in_29bar), .ZN(n736bar) );
  OR2_X1 U227 ( .A1(in_79), .A2(in_74), .ZN(n737) );
  AND2_X1 U227bar ( .A1(in_79bar), .A2(in_74bar), .ZN(n737bar) );
  OR2_X1 U228 ( .A1(n735), .A2(n734), .ZN(n789) );
  AND2_X1 U228bar ( .A1(n735bar), .A2(n734bar), .ZN(n789bar) );
  OR2_X1 U229 ( .A1(in[152]), .A2(in[140]), .ZN(n734) );
  AND2_X1 U229bar ( .A1(inbar[152]), .A2(inbar[140]), .ZN(n734bar) );
  OR2_X1 U230 ( .A1(in[155]), .A2(n733), .ZN(n735) );
  AND2_X1 U230bar ( .A1(inbar[155]), .A2(n733bar), .ZN(n735bar) );
  OR2_X1 U231 ( .A1(in[166]), .A2(in[165]), .ZN(n733) );
  AND2_X1 U231bar ( .A1(inbar[166]), .A2(inbar[165]), .ZN(n733bar) );
  OR2_X1 U232 ( .A1(n732), .A2(n731), .ZN(n791) );
  AND2_X1 U232bar ( .A1(n732bar), .A2(n731bar), .ZN(n791bar) );
  OR2_X1 U233 ( .A1(n730), .A2(n729), .ZN(n731) );
  AND2_X1 U233bar ( .A1(n730bar), .A2(n729bar), .ZN(n731bar) );
  OR2_X1 U234 ( .A1(in[202]), .A2(in[185]), .ZN(n729) );
  AND2_X1 U234bar ( .A1(inbar[202]), .A2(inbar[185]), .ZN(n729bar) );
  OR2_X1 U235 ( .A1(in[211]), .A2(n728), .ZN(n730) );
  AND2_X1 U235bar ( .A1(inbar[211]), .A2(n728bar), .ZN(n730bar) );
  OR2_X1 U236 ( .A1(in[255]), .A2(in[253]), .ZN(n728) );
  AND2_X1 U236bar ( .A1(inbar[255]), .A2(inbar[253]), .ZN(n728bar) );
  OR2_X1 U237 ( .A1(n727), .A2(n726), .ZN(n732) );
  AND2_X1 U237bar ( .A1(n727bar), .A2(n726bar), .ZN(n732bar) );
  OR2_X1 U238 ( .A1(in_35), .A2(in_15), .ZN(n726) );
  AND2_X1 U238bar ( .A1(in_35bar), .A2(in_15bar), .ZN(n726bar) );
  OR2_X1 U239 ( .A1(in_36), .A2(n725), .ZN(n727) );
  AND2_X1 U239bar ( .A1(in_36bar), .A2(n725bar), .ZN(n727bar) );
  OR2_X1 U240 ( .A1(in_48), .A2(in_40), .ZN(n725) );
  AND2_X1 U240bar ( .A1(in_48bar), .A2(in_40bar), .ZN(n725bar) );
  OR2_X1 U241 ( .A1(n724), .A2(n723), .ZN(out[1]) );
  AND2_X1 U241bar ( .A1(n724bar), .A2(n723bar), .ZN(outbar[1]) );
  OR2_X1 U242 ( .A1(n722), .A2(n721), .ZN(n723) );
  AND2_X1 U242bar ( .A1(n722bar), .A2(n721bar), .ZN(n723bar) );
  OR2_X1 U243 ( .A1(n720), .A2(n719), .ZN(n721) );
  AND2_X1 U243bar ( .A1(n720bar), .A2(n719bar), .ZN(n721bar) );
  OR2_X1 U244 ( .A1(n921), .A2(n887), .ZN(n719) );
  AND2_X1 U244bar ( .A1(n921bar), .A2(n887bar), .ZN(n719bar) );
  OR2_X1 U245 ( .A1(n718), .A2(n717), .ZN(n887) );
  AND2_X1 U245bar ( .A1(n718bar), .A2(n717bar), .ZN(n887bar) );
  OR2_X1 U246 ( .A1(n716), .A2(n715), .ZN(n717) );
  AND2_X1 U246bar ( .A1(n716bar), .A2(n715bar), .ZN(n717bar) );
  OR2_X1 U247 ( .A1(n714), .A2(n713), .ZN(n715) );
  AND2_X1 U247bar ( .A1(n714bar), .A2(n713bar), .ZN(n715bar) );
  OR2_X1 U248 ( .A1(in[116]), .A2(in[110]), .ZN(n713) );
  AND2_X1 U248bar ( .A1(inbar[116]), .A2(inbar[110]), .ZN(n713bar) );
  OR2_X1 U249 ( .A1(in[133]), .A2(in[130]), .ZN(n714) );
  AND2_X1 U249bar ( .A1(inbar[133]), .A2(inbar[130]), .ZN(n714bar) );
  OR2_X1 U250 ( .A1(n712), .A2(n711), .ZN(n716) );
  AND2_X1 U250bar ( .A1(n712bar), .A2(n711bar), .ZN(n716bar) );
  OR2_X1 U251 ( .A1(in[203]), .A2(in[135]), .ZN(n711) );
  AND2_X1 U251bar ( .A1(inbar[203]), .A2(inbar[135]), .ZN(n711bar) );
  OR2_X1 U252 ( .A1(in[232]), .A2(in[223]), .ZN(n712) );
  AND2_X1 U252bar ( .A1(inbar[232]), .A2(inbar[223]), .ZN(n712bar) );
  OR2_X1 U253 ( .A1(n710), .A2(n709), .ZN(n718) );
  AND2_X1 U253bar ( .A1(n710bar), .A2(n709bar), .ZN(n718bar) );
  OR2_X1 U254 ( .A1(n708), .A2(n707), .ZN(n709) );
  AND2_X1 U254bar ( .A1(n708bar), .A2(n707bar), .ZN(n709bar) );
  OR2_X1 U255 ( .A1(in[255]), .A2(in[233]), .ZN(n707) );
  AND2_X1 U255bar ( .A1(inbar[255]), .A2(inbar[233]), .ZN(n707bar) );
  OR2_X1 U256 ( .A1(in_53), .A2(in_34), .ZN(n708) );
  AND2_X1 U256bar ( .A1(in_53bar), .A2(in_34bar), .ZN(n708bar) );
  OR2_X1 U257 ( .A1(n706), .A2(n705), .ZN(n710) );
  AND2_X1 U257bar ( .A1(n706bar), .A2(n705bar), .ZN(n710bar) );
  OR2_X1 U258 ( .A1(in_57), .A2(in_55), .ZN(n705) );
  AND2_X1 U258bar ( .A1(in_57bar), .A2(in_55bar), .ZN(n705bar) );
  OR2_X1 U259 ( .A1(in_68), .A2(in_67), .ZN(n706) );
  AND2_X1 U259bar ( .A1(in_68bar), .A2(in_67bar), .ZN(n706bar) );
  OR2_X1 U260 ( .A1(n704), .A2(n703), .ZN(n921) );
  AND2_X1 U260bar ( .A1(n704bar), .A2(n703bar), .ZN(n921bar) );
  OR2_X1 U261 ( .A1(n702), .A2(n701), .ZN(n703) );
  AND2_X1 U261bar ( .A1(n702bar), .A2(n701bar), .ZN(n703bar) );
  OR2_X1 U262 ( .A1(n700), .A2(n699), .ZN(n701) );
  AND2_X1 U262bar ( .A1(n700bar), .A2(n699bar), .ZN(n701bar) );
  OR2_X1 U263 ( .A1(n944), .A2(n872), .ZN(n699) );
  AND2_X1 U263bar ( .A1(n944bar), .A2(n872bar), .ZN(n699bar) );
  OR2_X1 U264 ( .A1(n698), .A2(n697), .ZN(n872) );
  AND2_X1 U264bar ( .A1(n698bar), .A2(n697bar), .ZN(n872bar) );
  OR2_X1 U265 ( .A1(n696), .A2(n695), .ZN(n697) );
  AND2_X1 U265bar ( .A1(n696bar), .A2(n695bar), .ZN(n697bar) );
  OR2_X1 U266 ( .A1(n694), .A2(n693), .ZN(n695) );
  AND2_X1 U266bar ( .A1(n694bar), .A2(n693bar), .ZN(n695bar) );
  OR2_X1 U267 ( .A1(in[121]), .A2(in[102]), .ZN(n693) );
  AND2_X1 U267bar ( .A1(inbar[121]), .A2(inbar[102]), .ZN(n693bar) );
  OR2_X1 U268 ( .A1(in[162]), .A2(in[161]), .ZN(n694) );
  AND2_X1 U268bar ( .A1(inbar[162]), .A2(inbar[161]), .ZN(n694bar) );
  OR2_X1 U269 ( .A1(n692), .A2(n691), .ZN(n696) );
  AND2_X1 U269bar ( .A1(n692bar), .A2(n691bar), .ZN(n696bar) );
  OR2_X1 U270 ( .A1(in[192]), .A2(in[178]), .ZN(n691) );
  AND2_X1 U270bar ( .A1(inbar[192]), .A2(inbar[178]), .ZN(n691bar) );
  OR2_X1 U271 ( .A1(in[244]), .A2(in[209]), .ZN(n692) );
  AND2_X1 U271bar ( .A1(inbar[244]), .A2(inbar[209]), .ZN(n692bar) );
  OR2_X1 U272 ( .A1(n690), .A2(n689), .ZN(n698) );
  AND2_X1 U272bar ( .A1(n690bar), .A2(n689bar), .ZN(n698bar) );
  OR2_X1 U273 ( .A1(n688), .A2(n687), .ZN(n689) );
  AND2_X1 U273bar ( .A1(n688bar), .A2(n687bar), .ZN(n689bar) );
  OR2_X1 U274 ( .A1(in[90]), .A2(in[254]), .ZN(n687) );
  AND2_X1 U274bar ( .A1(inbar[90]), .A2(inbar[254]), .ZN(n687bar) );
  OR2_X1 U275 ( .A1(in_36), .A2(in_32), .ZN(n688) );
  AND2_X1 U275bar ( .A1(in_36bar), .A2(in_32bar), .ZN(n688bar) );
  OR2_X1 U276 ( .A1(n686), .A2(n685), .ZN(n690) );
  AND2_X1 U276bar ( .A1(n686bar), .A2(n685bar), .ZN(n690bar) );
  OR2_X1 U277 ( .A1(in_62), .A2(in_37), .ZN(n685) );
  AND2_X1 U277bar ( .A1(in_62bar), .A2(in_37bar), .ZN(n685bar) );
  OR2_X1 U278 ( .A1(in_75), .A2(in_73), .ZN(n686) );
  AND2_X1 U278bar ( .A1(in_75bar), .A2(in_73bar), .ZN(n686bar) );
  OR2_X1 U279 ( .A1(n684), .A2(n683), .ZN(n944) );
  AND2_X1 U279bar ( .A1(n684bar), .A2(n683bar), .ZN(n944bar) );
  OR2_X1 U280 ( .A1(n682), .A2(n681), .ZN(n683) );
  AND2_X1 U280bar ( .A1(n682bar), .A2(n681bar), .ZN(n683bar) );
  OR2_X1 U281 ( .A1(n680), .A2(n679), .ZN(n681) );
  AND2_X1 U281bar ( .A1(n680bar), .A2(n679bar), .ZN(n681bar) );
  OR2_X1 U282 ( .A1(in[171]), .A2(in[153]), .ZN(n679) );
  AND2_X1 U282bar ( .A1(inbar[171]), .A2(inbar[153]), .ZN(n679bar) );
  OR2_X1 U283 ( .A1(in[187]), .A2(in[176]), .ZN(n680) );
  AND2_X1 U283bar ( .A1(inbar[187]), .A2(inbar[176]), .ZN(n680bar) );
  OR2_X1 U284 ( .A1(n678), .A2(n677), .ZN(n682) );
  AND2_X1 U284bar ( .A1(n678bar), .A2(n677bar), .ZN(n682bar) );
  OR2_X1 U285 ( .A1(in[245]), .A2(in[211]), .ZN(n677) );
  AND2_X1 U285bar ( .A1(inbar[245]), .A2(inbar[211]), .ZN(n677bar) );
  OR2_X1 U286 ( .A1(in[97]), .A2(in[88]), .ZN(n678) );
  AND2_X1 U286bar ( .A1(inbar[97]), .A2(inbar[88]), .ZN(n678bar) );
  OR2_X1 U287 ( .A1(n676), .A2(n675), .ZN(n684) );
  AND2_X1 U287bar ( .A1(n676bar), .A2(n675bar), .ZN(n684bar) );
  OR2_X1 U288 ( .A1(n674), .A2(n673), .ZN(n675) );
  AND2_X1 U288bar ( .A1(n674bar), .A2(n673bar), .ZN(n675bar) );
  OR2_X1 U289 ( .A1(in_10), .A2(in_0), .ZN(n673) );
  AND2_X1 U289bar ( .A1(in_10bar), .A2(in_0bar), .ZN(n673bar) );
  OR2_X1 U290 ( .A1(in_59), .A2(in_5), .ZN(n674) );
  AND2_X1 U290bar ( .A1(in_59bar), .A2(in_5bar), .ZN(n674bar) );
  OR2_X1 U291 ( .A1(n672), .A2(n671), .ZN(n676) );
  AND2_X1 U291bar ( .A1(n672bar), .A2(n671bar), .ZN(n676bar) );
  OR2_X1 U292 ( .A1(in_60), .A2(in_6), .ZN(n671) );
  AND2_X1 U292bar ( .A1(in_60bar), .A2(in_6bar), .ZN(n671bar) );
  OR2_X1 U293 ( .A1(in_77), .A2(in_69), .ZN(n672) );
  AND2_X1 U293bar ( .A1(in_77bar), .A2(in_69bar), .ZN(n672bar) );
  OR2_X1 U294 ( .A1(in[113]), .A2(n864), .ZN(n700) );
  AND2_X1 U294bar ( .A1(inbar[113]), .A2(n864bar), .ZN(n700bar) );
  OR2_X1 U295 ( .A1(n670), .A2(n669), .ZN(n864) );
  AND2_X1 U295bar ( .A1(n670bar), .A2(n669bar), .ZN(n864bar) );
  OR2_X1 U296 ( .A1(n668), .A2(n667), .ZN(n669) );
  AND2_X1 U296bar ( .A1(n668bar), .A2(n667bar), .ZN(n669bar) );
  OR2_X1 U297 ( .A1(n666), .A2(n665), .ZN(n667) );
  AND2_X1 U297bar ( .A1(n666bar), .A2(n665bar), .ZN(n667bar) );
  OR2_X1 U298 ( .A1(in[125]), .A2(in[107]), .ZN(n665) );
  AND2_X1 U298bar ( .A1(inbar[125]), .A2(inbar[107]), .ZN(n665bar) );
  OR2_X1 U299 ( .A1(in[138]), .A2(in[126]), .ZN(n666) );
  AND2_X1 U299bar ( .A1(inbar[138]), .A2(inbar[126]), .ZN(n666bar) );
  OR2_X1 U300 ( .A1(n664), .A2(n663), .ZN(n668) );
  AND2_X1 U300bar ( .A1(n664bar), .A2(n663bar), .ZN(n668bar) );
  OR2_X1 U301 ( .A1(in[189]), .A2(in[143]), .ZN(n663) );
  AND2_X1 U301bar ( .A1(inbar[189]), .A2(inbar[143]), .ZN(n663bar) );
  OR2_X1 U302 ( .A1(in[99]), .A2(in[214]), .ZN(n664) );
  AND2_X1 U302bar ( .A1(inbar[99]), .A2(inbar[214]), .ZN(n664bar) );
  OR2_X1 U303 ( .A1(n662), .A2(n661), .ZN(n670) );
  AND2_X1 U303bar ( .A1(n662bar), .A2(n661bar), .ZN(n670bar) );
  OR2_X1 U304 ( .A1(n660), .A2(n659), .ZN(n661) );
  AND2_X1 U304bar ( .A1(n660bar), .A2(n659bar), .ZN(n661bar) );
  OR2_X1 U305 ( .A1(in_15), .A2(in_12), .ZN(n659) );
  AND2_X1 U305bar ( .A1(in_15bar), .A2(in_12bar), .ZN(n659bar) );
  OR2_X1 U306 ( .A1(in_20), .A2(in_2), .ZN(n660) );
  AND2_X1 U306bar ( .A1(in_20bar), .A2(in_2bar), .ZN(n660bar) );
  OR2_X1 U307 ( .A1(n658), .A2(n657), .ZN(n662) );
  AND2_X1 U307bar ( .A1(n658bar), .A2(n657bar), .ZN(n662bar) );
  OR2_X1 U308 ( .A1(in_30), .A2(in_3), .ZN(n657) );
  AND2_X1 U308bar ( .A1(in_30bar), .A2(in_3bar), .ZN(n657bar) );
  OR2_X1 U309 ( .A1(in_4), .A2(in_38), .ZN(n658) );
  AND2_X1 U309bar ( .A1(in_4bar), .A2(in_38bar), .ZN(n658bar) );
  OR2_X1 U310 ( .A1(n656), .A2(n655), .ZN(n702) );
  AND2_X1 U310bar ( .A1(n656bar), .A2(n655bar), .ZN(n702bar) );
  OR2_X1 U311 ( .A1(in[148]), .A2(in[137]), .ZN(n655) );
  AND2_X1 U311bar ( .A1(inbar[148]), .A2(inbar[137]), .ZN(n655bar) );
  OR2_X1 U312 ( .A1(in[149]), .A2(n654), .ZN(n656) );
  AND2_X1 U312bar ( .A1(inbar[149]), .A2(n654bar), .ZN(n656bar) );
  OR2_X1 U313 ( .A1(in[195]), .A2(in[190]), .ZN(n654) );
  AND2_X1 U313bar ( .A1(inbar[195]), .A2(inbar[190]), .ZN(n654bar) );
  OR2_X1 U314 ( .A1(n653), .A2(n652), .ZN(n704) );
  AND2_X1 U314bar ( .A1(n653bar), .A2(n652bar), .ZN(n704bar) );
  OR2_X1 U315 ( .A1(n651), .A2(n650), .ZN(n652) );
  AND2_X1 U315bar ( .A1(n651bar), .A2(n650bar), .ZN(n652bar) );
  OR2_X1 U316 ( .A1(in[98]), .A2(in[197]), .ZN(n650) );
  AND2_X1 U316bar ( .A1(inbar[98]), .A2(inbar[197]), .ZN(n650bar) );
  OR2_X1 U317 ( .A1(in_11), .A2(n649), .ZN(n651) );
  AND2_X1 U317bar ( .A1(in_11bar), .A2(n649bar), .ZN(n651bar) );
  OR2_X1 U318 ( .A1(in_26), .A2(in_14), .ZN(n649) );
  AND2_X1 U318bar ( .A1(in_26bar), .A2(in_14bar), .ZN(n649bar) );
  OR2_X1 U319 ( .A1(n648), .A2(n647), .ZN(n653) );
  AND2_X1 U319bar ( .A1(n648bar), .A2(n647bar), .ZN(n653bar) );
  OR2_X1 U320 ( .A1(in_35), .A2(in_27), .ZN(n647) );
  AND2_X1 U320bar ( .A1(in_35bar), .A2(in_27bar), .ZN(n647bar) );
  OR2_X1 U321 ( .A1(in_50), .A2(n646), .ZN(n648) );
  AND2_X1 U321bar ( .A1(in_50bar), .A2(n646bar), .ZN(n648bar) );
  OR2_X1 U322 ( .A1(in_78), .A2(in_61), .ZN(n646) );
  AND2_X1 U322bar ( .A1(in_78bar), .A2(in_61bar), .ZN(n646bar) );
  OR2_X1 U323 ( .A1(n942), .A2(n645), .ZN(n720) );
  AND2_X1 U323bar ( .A1(n942bar), .A2(n645bar), .ZN(n720bar) );
  OR2_X1 U324 ( .A1(in[106]), .A2(n863), .ZN(n645) );
  AND2_X1 U324bar ( .A1(inbar[106]), .A2(n863bar), .ZN(n645bar) );
  OR2_X1 U325 ( .A1(n644), .A2(n643), .ZN(n863) );
  AND2_X1 U325bar ( .A1(n644bar), .A2(n643bar), .ZN(n863bar) );
  OR2_X1 U326 ( .A1(n642), .A2(n641), .ZN(n643) );
  AND2_X1 U326bar ( .A1(n642bar), .A2(n641bar), .ZN(n643bar) );
  OR2_X1 U327 ( .A1(n640), .A2(n639), .ZN(n641) );
  AND2_X1 U327bar ( .A1(n640bar), .A2(n639bar), .ZN(n641bar) );
  OR2_X1 U328 ( .A1(in[127]), .A2(in[122]), .ZN(n639) );
  AND2_X1 U328bar ( .A1(inbar[127]), .A2(inbar[122]), .ZN(n639bar) );
  OR2_X1 U329 ( .A1(in[156]), .A2(in[132]), .ZN(n640) );
  AND2_X1 U329bar ( .A1(inbar[156]), .A2(inbar[132]), .ZN(n640bar) );
  OR2_X1 U330 ( .A1(n638), .A2(n637), .ZN(n642) );
  AND2_X1 U330bar ( .A1(n638bar), .A2(n637bar), .ZN(n642bar) );
  OR2_X1 U331 ( .A1(in[159]), .A2(in[157]), .ZN(n637) );
  AND2_X1 U331bar ( .A1(inbar[159]), .A2(inbar[157]), .ZN(n637bar) );
  OR2_X1 U332 ( .A1(in[185]), .A2(in[169]), .ZN(n638) );
  AND2_X1 U332bar ( .A1(inbar[185]), .A2(inbar[169]), .ZN(n638bar) );
  OR2_X1 U333 ( .A1(n636), .A2(n635), .ZN(n644) );
  AND2_X1 U333bar ( .A1(n636bar), .A2(n635bar), .ZN(n644bar) );
  OR2_X1 U334 ( .A1(n634), .A2(n633), .ZN(n635) );
  AND2_X1 U334bar ( .A1(n634bar), .A2(n633bar), .ZN(n635bar) );
  OR2_X1 U335 ( .A1(in[239]), .A2(in[218]), .ZN(n633) );
  AND2_X1 U335bar ( .A1(inbar[239]), .A2(inbar[218]), .ZN(n633bar) );
  OR2_X1 U336 ( .A1(in_13), .A2(in[87]), .ZN(n634) );
  AND2_X1 U336bar ( .A1(in_13bar), .A2(inbar[87]), .ZN(n634bar) );
  OR2_X1 U337 ( .A1(n632), .A2(n631), .ZN(n636) );
  AND2_X1 U337bar ( .A1(n632bar), .A2(n631bar), .ZN(n636bar) );
  OR2_X1 U338 ( .A1(in_72), .A2(in_70), .ZN(n631) );
  AND2_X1 U338bar ( .A1(in_72bar), .A2(in_70bar), .ZN(n631bar) );
  OR2_X1 U339 ( .A1(in_80), .A2(in_74), .ZN(n632) );
  AND2_X1 U339bar ( .A1(in_80bar), .A2(in_74bar), .ZN(n632bar) );
  OR2_X1 U340 ( .A1(n630), .A2(n629), .ZN(n942) );
  AND2_X1 U340bar ( .A1(n630bar), .A2(n629bar), .ZN(n942bar) );
  OR2_X1 U341 ( .A1(n628), .A2(n627), .ZN(n629) );
  AND2_X1 U341bar ( .A1(n628bar), .A2(n627bar), .ZN(n629bar) );
  OR2_X1 U342 ( .A1(n626), .A2(n625), .ZN(n627) );
  AND2_X1 U342bar ( .A1(n626bar), .A2(n625bar), .ZN(n627bar) );
  OR2_X1 U343 ( .A1(in[146]), .A2(in[100]), .ZN(n625) );
  AND2_X1 U343bar ( .A1(inbar[146]), .A2(inbar[100]), .ZN(n625bar) );
  OR2_X1 U344 ( .A1(in[168]), .A2(in[152]), .ZN(n626) );
  AND2_X1 U344bar ( .A1(inbar[168]), .A2(inbar[152]), .ZN(n626bar) );
  OR2_X1 U345 ( .A1(n624), .A2(n623), .ZN(n628) );
  AND2_X1 U345bar ( .A1(n624bar), .A2(n623bar), .ZN(n628bar) );
  OR2_X1 U346 ( .A1(in[199]), .A2(in[182]), .ZN(n623) );
  AND2_X1 U346bar ( .A1(inbar[199]), .A2(inbar[182]), .ZN(n623bar) );
  OR2_X1 U347 ( .A1(in[236]), .A2(in[204]), .ZN(n624) );
  AND2_X1 U347bar ( .A1(inbar[236]), .A2(inbar[204]), .ZN(n624bar) );
  OR2_X1 U348 ( .A1(n622), .A2(n621), .ZN(n630) );
  AND2_X1 U348bar ( .A1(n622bar), .A2(n621bar), .ZN(n630bar) );
  OR2_X1 U349 ( .A1(n620), .A2(n619), .ZN(n621) );
  AND2_X1 U349bar ( .A1(n620bar), .A2(n619bar), .ZN(n621bar) );
  OR2_X1 U350 ( .A1(in[89]), .A2(in[246]), .ZN(n619) );
  AND2_X1 U350bar ( .A1(inbar[89]), .A2(inbar[246]), .ZN(n619bar) );
  OR2_X1 U351 ( .A1(in[95]), .A2(in[92]), .ZN(n620) );
  AND2_X1 U351bar ( .A1(inbar[95]), .A2(inbar[92]), .ZN(n620bar) );
  OR2_X1 U352 ( .A1(n618), .A2(n617), .ZN(n622) );
  AND2_X1 U352bar ( .A1(n618bar), .A2(n617bar), .ZN(n622bar) );
  OR2_X1 U353 ( .A1(in_22), .A2(in_16), .ZN(n617) );
  AND2_X1 U353bar ( .A1(in_22bar), .A2(in_16bar), .ZN(n617bar) );
  OR2_X1 U354 ( .A1(in_51), .A2(in_49), .ZN(n618) );
  AND2_X1 U354bar ( .A1(in_51bar), .A2(in_49bar), .ZN(n618bar) );
  OR2_X1 U355 ( .A1(n616), .A2(n615), .ZN(n722) );
  AND2_X1 U355bar ( .A1(n616bar), .A2(n615bar), .ZN(n722bar) );
  OR2_X1 U356 ( .A1(in[158]), .A2(in[115]), .ZN(n615) );
  AND2_X1 U356bar ( .A1(inbar[158]), .A2(inbar[115]), .ZN(n615bar) );
  OR2_X1 U357 ( .A1(in[163]), .A2(n614), .ZN(n616) );
  AND2_X1 U357bar ( .A1(inbar[163]), .A2(n614bar), .ZN(n616bar) );
  OR2_X1 U358 ( .A1(in[206]), .A2(in[165]), .ZN(n614) );
  AND2_X1 U358bar ( .A1(inbar[206]), .A2(inbar[165]), .ZN(n614bar) );
  OR2_X1 U359 ( .A1(n613), .A2(n612), .ZN(n724) );
  AND2_X1 U359bar ( .A1(n613bar), .A2(n612bar), .ZN(n724bar) );
  OR2_X1 U360 ( .A1(n611), .A2(n610), .ZN(n612) );
  AND2_X1 U360bar ( .A1(n611bar), .A2(n610bar), .ZN(n612bar) );
  OR2_X1 U361 ( .A1(in[213]), .A2(in[207]), .ZN(n610) );
  AND2_X1 U361bar ( .A1(inbar[213]), .A2(inbar[207]), .ZN(n610bar) );
  OR2_X1 U362 ( .A1(in[215]), .A2(n609), .ZN(n611) );
  AND2_X1 U362bar ( .A1(inbar[215]), .A2(n609bar), .ZN(n611bar) );
  OR2_X1 U363 ( .A1(in[230]), .A2(in[220]), .ZN(n609) );
  AND2_X1 U363bar ( .A1(inbar[230]), .A2(inbar[220]), .ZN(n609bar) );
  OR2_X1 U364 ( .A1(n608), .A2(n607), .ZN(n613) );
  AND2_X1 U364bar ( .A1(n608bar), .A2(n607bar), .ZN(n613bar) );
  OR2_X1 U365 ( .A1(in[251]), .A2(in[234]), .ZN(n607) );
  AND2_X1 U365bar ( .A1(inbar[251]), .A2(inbar[234]), .ZN(n607bar) );
  OR2_X1 U366 ( .A1(in_17), .A2(n606), .ZN(n608) );
  AND2_X1 U366bar ( .A1(in_17bar), .A2(n606bar), .ZN(n608bar) );
  OR2_X1 U367 ( .A1(in_65), .A2(in_56), .ZN(n606) );
  AND2_X1 U367bar ( .A1(in_65bar), .A2(in_56bar), .ZN(n606bar) );
  OR2_X1 U368 ( .A1(n605), .A2(n604), .ZN(out[0]) );
  AND2_X1 U368bar ( .A1(n605bar), .A2(n604bar), .ZN(outbar[0]) );
  OR2_X1 U369 ( .A1(n603), .A2(n602), .ZN(n604) );
  AND2_X1 U369bar ( .A1(n603bar), .A2(n602bar), .ZN(n604bar) );
  OR2_X1 U370 ( .A1(n601), .A2(n600), .ZN(n602) );
  AND2_X1 U370bar ( .A1(n601bar), .A2(n600bar), .ZN(n602bar) );
  OR2_X1 U371 ( .A1(n820), .A2(n785), .ZN(n600) );
  AND2_X1 U371bar ( .A1(n820bar), .A2(n785bar), .ZN(n600bar) );
  OR2_X1 U372 ( .A1(n599), .A2(n598), .ZN(n785) );
  AND2_X1 U372bar ( .A1(n599bar), .A2(n598bar), .ZN(n785bar) );
  OR2_X1 U373 ( .A1(n597), .A2(n596), .ZN(n598) );
  AND2_X1 U373bar ( .A1(n597bar), .A2(n596bar), .ZN(n598bar) );
  OR2_X1 U374 ( .A1(n595), .A2(n594), .ZN(n596) );
  AND2_X1 U374bar ( .A1(n595bar), .A2(n594bar), .ZN(n596bar) );
  OR2_X1 U375 ( .A1(in[135]), .A2(in[104]), .ZN(n594) );
  AND2_X1 U375bar ( .A1(inbar[135]), .A2(inbar[104]), .ZN(n594bar) );
  OR2_X1 U376 ( .A1(in[188]), .A2(in[178]), .ZN(n595) );
  AND2_X1 U376bar ( .A1(inbar[188]), .A2(inbar[178]), .ZN(n595bar) );
  OR2_X1 U377 ( .A1(n593), .A2(n592), .ZN(n597) );
  AND2_X1 U377bar ( .A1(n593bar), .A2(n592bar), .ZN(n597bar) );
  OR2_X1 U378 ( .A1(in[217]), .A2(in[194]), .ZN(n592) );
  AND2_X1 U378bar ( .A1(inbar[217]), .A2(inbar[194]), .ZN(n592bar) );
  OR2_X1 U379 ( .A1(in[237]), .A2(in[218]), .ZN(n593) );
  AND2_X1 U379bar ( .A1(inbar[237]), .A2(inbar[218]), .ZN(n593bar) );
  OR2_X1 U380 ( .A1(n591), .A2(n590), .ZN(n599) );
  AND2_X1 U380bar ( .A1(n591bar), .A2(n590bar), .ZN(n599bar) );
  OR2_X1 U381 ( .A1(n589), .A2(n588), .ZN(n590) );
  AND2_X1 U381bar ( .A1(n589bar), .A2(n588bar), .ZN(n590bar) );
  OR2_X1 U382 ( .A1(in_2), .A2(in_10), .ZN(n588) );
  AND2_X1 U382bar ( .A1(in_2bar), .A2(in_10bar), .ZN(n588bar) );
  OR2_X1 U383 ( .A1(in_47), .A2(in_22), .ZN(n589) );
  AND2_X1 U383bar ( .A1(in_47bar), .A2(in_22bar), .ZN(n589bar) );
  OR2_X1 U384 ( .A1(n587), .A2(n586), .ZN(n591) );
  AND2_X1 U384bar ( .A1(n587bar), .A2(n586bar), .ZN(n591bar) );
  OR2_X1 U385 ( .A1(in_56), .A2(in_54), .ZN(n586) );
  AND2_X1 U385bar ( .A1(in_56bar), .A2(in_54bar), .ZN(n586bar) );
  OR2_X1 U386 ( .A1(in_63), .A2(in_61), .ZN(n587) );
  AND2_X1 U386bar ( .A1(in_63bar), .A2(in_61bar), .ZN(n587bar) );
  OR2_X1 U387 ( .A1(n585), .A2(n584), .ZN(n820) );
  AND2_X1 U387bar ( .A1(n585bar), .A2(n584bar), .ZN(n820bar) );
  OR2_X1 U388 ( .A1(n583), .A2(n582), .ZN(n584) );
  AND2_X1 U388bar ( .A1(n583bar), .A2(n582bar), .ZN(n584bar) );
  OR2_X1 U389 ( .A1(n581), .A2(n580), .ZN(n582) );
  AND2_X1 U389bar ( .A1(n581bar), .A2(n580bar), .ZN(n582bar) );
  OR2_X1 U390 ( .A1(in[158]), .A2(in[142]), .ZN(n580) );
  AND2_X1 U390bar ( .A1(inbar[158]), .A2(inbar[142]), .ZN(n580bar) );
  OR2_X1 U391 ( .A1(in[175]), .A2(in[164]), .ZN(n581) );
  AND2_X1 U391bar ( .A1(inbar[175]), .A2(inbar[164]), .ZN(n581bar) );
  OR2_X1 U392 ( .A1(n579), .A2(n578), .ZN(n583) );
  AND2_X1 U392bar ( .A1(n579bar), .A2(n578bar), .ZN(n583bar) );
  OR2_X1 U393 ( .A1(in[228]), .A2(in[204]), .ZN(n578) );
  AND2_X1 U393bar ( .A1(inbar[228]), .A2(inbar[204]), .ZN(n578bar) );
  OR2_X1 U394 ( .A1(in[91]), .A2(in[87]), .ZN(n579) );
  AND2_X1 U394bar ( .A1(inbar[91]), .A2(inbar[87]), .ZN(n579bar) );
  OR2_X1 U395 ( .A1(n577), .A2(n576), .ZN(n585) );
  AND2_X1 U395bar ( .A1(n577bar), .A2(n576bar), .ZN(n585bar) );
  OR2_X1 U396 ( .A1(n575), .A2(n574), .ZN(n576) );
  AND2_X1 U396bar ( .A1(n575bar), .A2(n574bar), .ZN(n576bar) );
  OR2_X1 U397 ( .A1(in_21), .A2(in_11), .ZN(n574) );
  AND2_X1 U397bar ( .A1(in_21bar), .A2(in_11bar), .ZN(n574bar) );
  OR2_X1 U398 ( .A1(in_5), .A2(in_3), .ZN(n575) );
  AND2_X1 U398bar ( .A1(in_5bar), .A2(in_3bar), .ZN(n575bar) );
  OR2_X1 U399 ( .A1(n573), .A2(n572), .ZN(n577) );
  AND2_X1 U399bar ( .A1(n573bar), .A2(n572bar), .ZN(n577bar) );
  OR2_X1 U400 ( .A1(in_68), .A2(in_64), .ZN(n572) );
  AND2_X1 U400bar ( .A1(in_68bar), .A2(in_64bar), .ZN(n572bar) );
  OR2_X1 U401 ( .A1(in_76), .A2(in_73), .ZN(n573) );
  AND2_X1 U401bar ( .A1(in_76bar), .A2(in_73bar), .ZN(n573bar) );
  OR2_X1 U402 ( .A1(n778), .A2(n571), .ZN(n601) );
  AND2_X1 U402bar ( .A1(n778bar), .A2(n571bar), .ZN(n601bar) );
  OR2_X1 U403 ( .A1(in[100]), .A2(n965), .ZN(n571) );
  AND2_X1 U403bar ( .A1(inbar[100]), .A2(n965bar), .ZN(n571bar) );
  OR2_X1 U404 ( .A1(n570), .A2(n569), .ZN(n965) );
  AND2_X1 U404bar ( .A1(n570bar), .A2(n569bar), .ZN(n965bar) );
  OR2_X1 U405 ( .A1(n568), .A2(n567), .ZN(n569) );
  AND2_X1 U405bar ( .A1(n568bar), .A2(n567bar), .ZN(n569bar) );
  OR2_X1 U406 ( .A1(n566), .A2(n565), .ZN(n567) );
  AND2_X1 U406bar ( .A1(n566bar), .A2(n565bar), .ZN(n567bar) );
  OR2_X1 U407 ( .A1(n817), .A2(n750), .ZN(n565) );
  AND2_X1 U407bar ( .A1(n817bar), .A2(n750bar), .ZN(n565bar) );
  OR2_X1 U408 ( .A1(n564), .A2(n563), .ZN(n750) );
  AND2_X1 U408bar ( .A1(n564bar), .A2(n563bar), .ZN(n750bar) );
  OR2_X1 U409 ( .A1(n562), .A2(n561), .ZN(n563) );
  AND2_X1 U409bar ( .A1(n562bar), .A2(n561bar), .ZN(n563bar) );
  OR2_X1 U410 ( .A1(n560), .A2(n559), .ZN(n561) );
  AND2_X1 U410bar ( .A1(n560bar), .A2(n559bar), .ZN(n561bar) );
  OR2_X1 U411 ( .A1(in[119]), .A2(in[103]), .ZN(n559) );
  AND2_X1 U411bar ( .A1(inbar[119]), .A2(inbar[103]), .ZN(n559bar) );
  OR2_X1 U412 ( .A1(in[137]), .A2(in[133]), .ZN(n560) );
  AND2_X1 U412bar ( .A1(inbar[137]), .A2(inbar[133]), .ZN(n560bar) );
  OR2_X1 U413 ( .A1(n558), .A2(n557), .ZN(n562) );
  AND2_X1 U413bar ( .A1(n558bar), .A2(n557bar), .ZN(n562bar) );
  OR2_X1 U414 ( .A1(in[176]), .A2(in[173]), .ZN(n557) );
  AND2_X1 U414bar ( .A1(inbar[176]), .A2(inbar[173]), .ZN(n557bar) );
  OR2_X1 U415 ( .A1(in[210]), .A2(in[181]), .ZN(n558) );
  AND2_X1 U415bar ( .A1(inbar[210]), .A2(inbar[181]), .ZN(n558bar) );
  OR2_X1 U416 ( .A1(n556), .A2(n555), .ZN(n564) );
  AND2_X1 U416bar ( .A1(n556bar), .A2(n555bar), .ZN(n564bar) );
  OR2_X1 U417 ( .A1(n554), .A2(n553), .ZN(n555) );
  AND2_X1 U417bar ( .A1(n554bar), .A2(n553bar), .ZN(n555bar) );
  OR2_X1 U418 ( .A1(in_13), .A2(in[234]), .ZN(n553) );
  AND2_X1 U418bar ( .A1(in_13bar), .A2(inbar[234]), .ZN(n553bar) );
  OR2_X1 U419 ( .A1(in_38), .A2(in_32), .ZN(n554) );
  AND2_X1 U419bar ( .A1(in_38bar), .A2(in_32bar), .ZN(n554bar) );
  OR2_X1 U420 ( .A1(n552), .A2(n551), .ZN(n556) );
  AND2_X1 U420bar ( .A1(n552bar), .A2(n551bar), .ZN(n556bar) );
  OR2_X1 U421 ( .A1(in_42), .A2(in_41), .ZN(n551) );
  AND2_X1 U421bar ( .A1(in_42bar), .A2(in_41bar), .ZN(n551bar) );
  OR2_X1 U422 ( .A1(in_7), .A2(in_49), .ZN(n552) );
  AND2_X1 U422bar ( .A1(in_7bar), .A2(in_49bar), .ZN(n552bar) );
  OR2_X1 U423 ( .A1(n550), .A2(n549), .ZN(n817) );
  AND2_X1 U423bar ( .A1(n550bar), .A2(n549bar), .ZN(n817bar) );
  OR2_X1 U424 ( .A1(n548), .A2(n547), .ZN(n549) );
  AND2_X1 U424bar ( .A1(n548bar), .A2(n547bar), .ZN(n549bar) );
  OR2_X1 U425 ( .A1(n546), .A2(n545), .ZN(n547) );
  AND2_X1 U425bar ( .A1(n546bar), .A2(n545bar), .ZN(n547bar) );
  OR2_X1 U426 ( .A1(in[159]), .A2(in[105]), .ZN(n545) );
  AND2_X1 U426bar ( .A1(inbar[159]), .A2(inbar[105]), .ZN(n545bar) );
  OR2_X1 U427 ( .A1(in[206]), .A2(in[183]), .ZN(n546) );
  AND2_X1 U427bar ( .A1(inbar[206]), .A2(inbar[183]), .ZN(n546bar) );
  OR2_X1 U428 ( .A1(n544), .A2(n543), .ZN(n548) );
  AND2_X1 U428bar ( .A1(n544bar), .A2(n543bar), .ZN(n548bar) );
  OR2_X1 U429 ( .A1(in[229]), .A2(in[219]), .ZN(n543) );
  AND2_X1 U429bar ( .A1(inbar[229]), .A2(inbar[219]), .ZN(n543bar) );
  OR2_X1 U430 ( .A1(in[235]), .A2(in[232]), .ZN(n544) );
  AND2_X1 U430bar ( .A1(inbar[235]), .A2(inbar[232]), .ZN(n544bar) );
  OR2_X1 U431 ( .A1(n542), .A2(n541), .ZN(n550) );
  AND2_X1 U431bar ( .A1(n542bar), .A2(n541bar), .ZN(n550bar) );
  OR2_X1 U432 ( .A1(n540), .A2(n539), .ZN(n541) );
  AND2_X1 U432bar ( .A1(n540bar), .A2(n539bar), .ZN(n541bar) );
  OR2_X1 U433 ( .A1(in[249]), .A2(in[242]), .ZN(n539) );
  AND2_X1 U433bar ( .A1(inbar[249]), .A2(inbar[242]), .ZN(n539bar) );
  OR2_X1 U434 ( .A1(in[89]), .A2(in[254]), .ZN(n540) );
  AND2_X1 U434bar ( .A1(inbar[89]), .A2(inbar[254]), .ZN(n540bar) );
  OR2_X1 U435 ( .A1(n538), .A2(n537), .ZN(n542) );
  AND2_X1 U435bar ( .A1(n538bar), .A2(n537bar), .ZN(n542bar) );
  OR2_X1 U436 ( .A1(in_14), .A2(in[99]), .ZN(n537) );
  AND2_X1 U436bar ( .A1(in_14bar), .A2(inbar[99]), .ZN(n537bar) );
  OR2_X1 U437 ( .A1(in_60), .A2(in_18), .ZN(n538) );
  AND2_X1 U437bar ( .A1(in_60bar), .A2(in_18bar), .ZN(n538bar) );
  OR2_X1 U438 ( .A1(in[113]), .A2(n763), .ZN(n566) );
  AND2_X1 U438bar ( .A1(inbar[113]), .A2(n763bar), .ZN(n566bar) );
  OR2_X1 U439 ( .A1(n536), .A2(n535), .ZN(n763) );
  AND2_X1 U439bar ( .A1(n536bar), .A2(n535bar), .ZN(n763bar) );
  OR2_X1 U440 ( .A1(n534), .A2(n533), .ZN(n535) );
  AND2_X1 U440bar ( .A1(n534bar), .A2(n533bar), .ZN(n535bar) );
  OR2_X1 U441 ( .A1(n532), .A2(n531), .ZN(n533) );
  AND2_X1 U441bar ( .A1(n532bar), .A2(n531bar), .ZN(n533bar) );
  OR2_X1 U442 ( .A1(in[115]), .A2(in[110]), .ZN(n531) );
  AND2_X1 U442bar ( .A1(inbar[115]), .A2(inbar[110]), .ZN(n531bar) );
  OR2_X1 U443 ( .A1(in[125]), .A2(in[117]), .ZN(n532) );
  AND2_X1 U443bar ( .A1(inbar[125]), .A2(inbar[117]), .ZN(n532bar) );
  OR2_X1 U444 ( .A1(n530), .A2(n529), .ZN(n534) );
  AND2_X1 U444bar ( .A1(n530bar), .A2(n529bar), .ZN(n534bar) );
  OR2_X1 U445 ( .A1(in[180]), .A2(in[128]), .ZN(n529) );
  AND2_X1 U445bar ( .A1(inbar[180]), .A2(inbar[128]), .ZN(n529bar) );
  OR2_X1 U446 ( .A1(in[205]), .A2(in[201]), .ZN(n530) );
  AND2_X1 U446bar ( .A1(inbar[205]), .A2(inbar[201]), .ZN(n530bar) );
  OR2_X1 U447 ( .A1(n528), .A2(n527), .ZN(n536) );
  AND2_X1 U447bar ( .A1(n528bar), .A2(n527bar), .ZN(n536bar) );
  OR2_X1 U448 ( .A1(n526), .A2(n525), .ZN(n527) );
  AND2_X1 U448bar ( .A1(n526bar), .A2(n525bar), .ZN(n527bar) );
  OR2_X1 U449 ( .A1(in[244]), .A2(in[239]), .ZN(n525) );
  AND2_X1 U449bar ( .A1(inbar[244]), .A2(inbar[239]), .ZN(n525bar) );
  OR2_X1 U450 ( .A1(in[95]), .A2(in[83]), .ZN(n526) );
  AND2_X1 U450bar ( .A1(inbar[95]), .A2(inbar[83]), .ZN(n526bar) );
  OR2_X1 U451 ( .A1(n524), .A2(n523), .ZN(n528) );
  AND2_X1 U451bar ( .A1(n524bar), .A2(n523bar), .ZN(n528bar) );
  OR2_X1 U452 ( .A1(in_24), .A2(in[97]), .ZN(n523) );
  AND2_X1 U452bar ( .A1(in_24bar), .A2(inbar[97]), .ZN(n523bar) );
  OR2_X1 U453 ( .A1(in_33), .A2(in_27), .ZN(n524) );
  AND2_X1 U453bar ( .A1(in_33bar), .A2(in_27bar), .ZN(n524bar) );
  OR2_X1 U454 ( .A1(n522), .A2(n521), .ZN(n568) );
  AND2_X1 U454bar ( .A1(n522bar), .A2(n521bar), .ZN(n568bar) );
  OR2_X1 U455 ( .A1(in[145]), .A2(in[126]), .ZN(n521) );
  AND2_X1 U455bar ( .A1(inbar[145]), .A2(inbar[126]), .ZN(n521bar) );
  OR2_X1 U456 ( .A1(in[169]), .A2(n520), .ZN(n522) );
  AND2_X1 U456bar ( .A1(inbar[169]), .A2(n520bar), .ZN(n522bar) );
  OR2_X1 U457 ( .A1(in[221]), .A2(in[172]), .ZN(n520) );
  AND2_X1 U457bar ( .A1(inbar[221]), .A2(inbar[172]), .ZN(n520bar) );
  OR2_X1 U458 ( .A1(n519), .A2(n518), .ZN(n570) );
  AND2_X1 U458bar ( .A1(n519bar), .A2(n518bar), .ZN(n570bar) );
  OR2_X1 U459 ( .A1(n517), .A2(n516), .ZN(n518) );
  AND2_X1 U459bar ( .A1(n517bar), .A2(n516bar), .ZN(n518bar) );
  OR2_X1 U460 ( .A1(in[241]), .A2(in[224]), .ZN(n516) );
  AND2_X1 U460bar ( .A1(inbar[241]), .A2(inbar[224]), .ZN(n516bar) );
  OR2_X1 U461 ( .A1(in[86]), .A2(n515), .ZN(n517) );
  AND2_X1 U461bar ( .A1(inbar[86]), .A2(n515bar), .ZN(n517bar) );
  OR2_X1 U462 ( .A1(in_43), .A2(in_34), .ZN(n515) );
  AND2_X1 U462bar ( .A1(in_43bar), .A2(in_34bar), .ZN(n515bar) );
  OR2_X1 U463 ( .A1(n514), .A2(n513), .ZN(n519) );
  AND2_X1 U463bar ( .A1(n514bar), .A2(n513bar), .ZN(n519bar) );
  OR2_X1 U464 ( .A1(in_65), .A2(in_51), .ZN(n513) );
  AND2_X1 U464bar ( .A1(in_65bar), .A2(in_51bar), .ZN(n513bar) );
  OR2_X1 U465 ( .A1(in_75), .A2(n512), .ZN(n514) );
  AND2_X1 U465bar ( .A1(in_75bar), .A2(n512bar), .ZN(n514bar) );
  OR2_X1 U466 ( .A1(in_81), .A2(in_77), .ZN(n512) );
  AND2_X1 U466bar ( .A1(in_81bar), .A2(in_77bar), .ZN(n512bar) );
  OR2_X1 U467 ( .A1(n511), .A2(n510), .ZN(n778) );
  AND2_X1 U467bar ( .A1(n511bar), .A2(n510bar), .ZN(n778bar) );
  OR2_X1 U468 ( .A1(n509), .A2(n508), .ZN(n510) );
  AND2_X1 U468bar ( .A1(n509bar), .A2(n508bar), .ZN(n510bar) );
  OR2_X1 U469 ( .A1(n507), .A2(n506), .ZN(n508) );
  AND2_X1 U469bar ( .A1(n507bar), .A2(n506bar), .ZN(n508bar) );
  OR2_X1 U470 ( .A1(in[107]), .A2(in[101]), .ZN(n506) );
  AND2_X1 U470bar ( .A1(inbar[107]), .A2(inbar[101]), .ZN(n506bar) );
  OR2_X1 U471 ( .A1(in[139]), .A2(in[132]), .ZN(n507) );
  AND2_X1 U471bar ( .A1(inbar[139]), .A2(inbar[132]), .ZN(n507bar) );
  OR2_X1 U472 ( .A1(n505), .A2(n504), .ZN(n509) );
  AND2_X1 U472bar ( .A1(n505bar), .A2(n504bar), .ZN(n509bar) );
  OR2_X1 U473 ( .A1(in[146]), .A2(in[141]), .ZN(n504) );
  AND2_X1 U473bar ( .A1(inbar[146]), .A2(inbar[141]), .ZN(n504bar) );
  OR2_X1 U474 ( .A1(in[203]), .A2(in[179]), .ZN(n505) );
  AND2_X1 U474bar ( .A1(inbar[203]), .A2(inbar[179]), .ZN(n505bar) );
  OR2_X1 U475 ( .A1(n503), .A2(n502), .ZN(n511) );
  AND2_X1 U475bar ( .A1(n503bar), .A2(n502bar), .ZN(n511bar) );
  OR2_X1 U476 ( .A1(n501), .A2(n500), .ZN(n502) );
  AND2_X1 U476bar ( .A1(n501bar), .A2(n500bar), .ZN(n502bar) );
  OR2_X1 U477 ( .A1(in[243]), .A2(in[222]), .ZN(n500) );
  AND2_X1 U477bar ( .A1(inbar[243]), .A2(inbar[222]), .ZN(n500bar) );
  OR2_X1 U478 ( .A1(in[251]), .A2(in[250]), .ZN(n501) );
  AND2_X1 U478bar ( .A1(inbar[251]), .A2(inbar[250]), .ZN(n501bar) );
  OR2_X1 U479 ( .A1(n499), .A2(n498), .ZN(n503) );
  AND2_X1 U479bar ( .A1(n499bar), .A2(n498bar), .ZN(n503bar) );
  OR2_X1 U480 ( .A1(in_37), .A2(in_19), .ZN(n498) );
  AND2_X1 U480bar ( .A1(in_37bar), .A2(in_19bar), .ZN(n498bar) );
  OR2_X1 U481 ( .A1(in_78), .A2(in_6), .ZN(n499) );
  AND2_X1 U481bar ( .A1(in_78bar), .A2(in_6bar), .ZN(n499bar) );
  OR2_X1 U482 ( .A1(n497), .A2(n496), .ZN(n603) );
  AND2_X1 U482bar ( .A1(n497bar), .A2(n496bar), .ZN(n603bar) );
  OR2_X1 U483 ( .A1(in[112]), .A2(in[102]), .ZN(n496) );
  AND2_X1 U483bar ( .A1(inbar[112]), .A2(inbar[102]), .ZN(n496bar) );
  OR2_X1 U484 ( .A1(in[123]), .A2(n495), .ZN(n497) );
  AND2_X1 U484bar ( .A1(inbar[123]), .A2(n495bar), .ZN(n497bar) );
  OR2_X1 U485 ( .A1(in[143]), .A2(in[130]), .ZN(n495) );
  AND2_X1 U485bar ( .A1(inbar[143]), .A2(inbar[130]), .ZN(n495bar) );
  OR2_X1 U486 ( .A1(n494), .A2(n493), .ZN(n605) );
  AND2_X1 U486bar ( .A1(n494bar), .A2(n493bar), .ZN(n605bar) );
  OR2_X1 U487 ( .A1(n492), .A2(n491), .ZN(n493) );
  AND2_X1 U487bar ( .A1(n492bar), .A2(n491bar), .ZN(n493bar) );
  OR2_X1 U488 ( .A1(in[216]), .A2(in[213]), .ZN(n491) );
  AND2_X1 U488bar ( .A1(inbar[216]), .A2(inbar[213]), .ZN(n491bar) );
  OR2_X1 U489 ( .A1(in[227]), .A2(n490), .ZN(n492) );
  AND2_X1 U489bar ( .A1(inbar[227]), .A2(n490bar), .ZN(n492bar) );
  OR2_X1 U490 ( .A1(in_0), .A2(in[248]), .ZN(n490) );
  AND2_X1 U490bar ( .A1(in_0bar), .A2(inbar[248]), .ZN(n490bar) );
  OR2_X1 U491 ( .A1(n489), .A2(n488), .ZN(n494) );
  AND2_X1 U491bar ( .A1(n489bar), .A2(n488bar), .ZN(n494bar) );
  OR2_X1 U492 ( .A1(in_46), .A2(in_44), .ZN(n488) );
  AND2_X1 U492bar ( .A1(in_46bar), .A2(in_44bar), .ZN(n488bar) );
  OR2_X1 U493 ( .A1(in_50), .A2(n487), .ZN(n489) );
  AND2_X1 U493bar ( .A1(in_50bar), .A2(n487bar), .ZN(n489bar) );
  OR2_X1 U494 ( .A1(in_9), .A2(in_80), .ZN(n487) );
  AND2_X1 U494bar ( .A1(in_9bar), .A2(in_80bar), .ZN(n487bar) );
endmodule

module sBox_1 ( in, inbar, out, outbar );

  input wire [7:0] in;
  input wire [7:0] inbar;
//input_done

  output wire [7:0] out;
  output wire [7:0] outbar;
//output_done

  wire [255:0] decodeOut;
  wire [255:0] decodeOutbar;
//wire_done

  decode_1 dec ( .in(in), .inbar(inbar), .out(decodeOut), .outbar(decodeOutbar) );
  encode_1 enc ( .in(decodeOut), .inbar(decodeOutbar), .out(out), .outbar(outbar) );
endmodule

module CD2_5 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD2_6 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD2_7 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD2_8 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD4_3 ( a, abar, b, bbar, y, ybar );

  input wire [3:0] a;
  input wire [3:0] b;
  input wire [3:0] abar;
  input wire [3:0] bbar;
//input_done

  output wire [15:0] y;
  output wire [15:0] ybar;
//output_done

//wire_done

  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]) );
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]) );
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]) );
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]) );
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]) );
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]) );
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]) );
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]) );
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]) );
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]) );
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]) );
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]) );
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]) );
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]) );
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]) );
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]) );
endmodule

module CD4_4 ( a, abar, b, bbar, y, ybar );

  input wire [3:0] a;
  input wire [3:0] b;
  input wire [3:0] abar;
  input wire [3:0] bbar;
//input_done

  output wire [15:0] y;
  output wire [15:0] ybar;
//output_done

//wire_done

  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]) );
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]) );
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]) );
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]) );
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]) );
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]) );
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]) );
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]) );
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]) );
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]) );
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]) );
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]) );
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]) );
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]) );
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]) );
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]) );
endmodule

module CD16_2 ( a, abar, b, bbar, y, ybar );

  input wire [15:0] a;
  input wire [15:0] b;
  input wire [15:0] abar;
  input wire [15:0] bbar;
//input_done

  output wire [255:0] y;
  output wire [255:0] ybar;
//output_done

//wire_done

  AND2_X1 U1 ( .A1(b[9]), .A2(a[0]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[9]), .A2(abar[0]), .ZN(ybar[9]) );
  AND2_X1 U2 ( .A1(b[3]), .A2(a[6]), .ZN(y[99]) );
  OR2_X1 U2bar ( .A1(bbar[3]), .A2(abar[6]), .ZN(ybar[99]) );
  AND2_X1 U3 ( .A1(b[2]), .A2(a[6]), .ZN(y[98]) );
  OR2_X1 U3bar ( .A1(bbar[2]), .A2(abar[6]), .ZN(ybar[98]) );
  AND2_X1 U4 ( .A1(b[1]), .A2(a[6]), .ZN(y[97]) );
  OR2_X1 U4bar ( .A1(bbar[1]), .A2(abar[6]), .ZN(ybar[97]) );
  AND2_X1 U5 ( .A1(b[0]), .A2(a[6]), .ZN(y[96]) );
  OR2_X1 U5bar ( .A1(bbar[0]), .A2(abar[6]), .ZN(ybar[96]) );
  AND2_X1 U6 ( .A1(b[15]), .A2(a[5]), .ZN(y[95]) );
  OR2_X1 U6bar ( .A1(bbar[15]), .A2(abar[5]), .ZN(ybar[95]) );
  AND2_X1 U7 ( .A1(b[14]), .A2(a[5]), .ZN(y[94]) );
  OR2_X1 U7bar ( .A1(bbar[14]), .A2(abar[5]), .ZN(ybar[94]) );
  AND2_X1 U8 ( .A1(b[13]), .A2(a[5]), .ZN(y[93]) );
  OR2_X1 U8bar ( .A1(bbar[13]), .A2(abar[5]), .ZN(ybar[93]) );
  AND2_X1 U9 ( .A1(b[12]), .A2(a[5]), .ZN(y[92]) );
  OR2_X1 U9bar ( .A1(bbar[12]), .A2(abar[5]), .ZN(ybar[92]) );
  AND2_X1 U10 ( .A1(b[11]), .A2(a[5]), .ZN(y[91]) );
  OR2_X1 U10bar ( .A1(bbar[11]), .A2(abar[5]), .ZN(ybar[91]) );
  AND2_X1 U11 ( .A1(b[10]), .A2(a[5]), .ZN(y[90]) );
  OR2_X1 U11bar ( .A1(bbar[10]), .A2(abar[5]), .ZN(ybar[90]) );
  AND2_X1 U12 ( .A1(b[8]), .A2(a[0]), .ZN(y[8]) );
  OR2_X1 U12bar ( .A1(bbar[8]), .A2(abar[0]), .ZN(ybar[8]) );
  AND2_X1 U13 ( .A1(a[5]), .A2(b[9]), .ZN(y[89]) );
  OR2_X1 U13bar ( .A1(abar[5]), .A2(bbar[9]), .ZN(ybar[89]) );
  AND2_X1 U14 ( .A1(b[8]), .A2(a[5]), .ZN(y[88]) );
  OR2_X1 U14bar ( .A1(bbar[8]), .A2(abar[5]), .ZN(ybar[88]) );
  AND2_X1 U15 ( .A1(b[7]), .A2(a[5]), .ZN(y[87]) );
  OR2_X1 U15bar ( .A1(bbar[7]), .A2(abar[5]), .ZN(ybar[87]) );
  AND2_X1 U16 ( .A1(b[6]), .A2(a[5]), .ZN(y[86]) );
  OR2_X1 U16bar ( .A1(bbar[6]), .A2(abar[5]), .ZN(ybar[86]) );
  AND2_X1 U17 ( .A1(b[5]), .A2(a[5]), .ZN(y[85]) );
  OR2_X1 U17bar ( .A1(bbar[5]), .A2(abar[5]), .ZN(ybar[85]) );
  AND2_X1 U18 ( .A1(b[4]), .A2(a[5]), .ZN(y[84]) );
  OR2_X1 U18bar ( .A1(bbar[4]), .A2(abar[5]), .ZN(ybar[84]) );
  AND2_X1 U19 ( .A1(a[5]), .A2(b[3]), .ZN(y[83]) );
  OR2_X1 U19bar ( .A1(abar[5]), .A2(bbar[3]), .ZN(ybar[83]) );
  AND2_X1 U20 ( .A1(a[5]), .A2(b[2]), .ZN(y[82]) );
  OR2_X1 U20bar ( .A1(abar[5]), .A2(bbar[2]), .ZN(ybar[82]) );
  AND2_X1 U21 ( .A1(a[5]), .A2(b[1]), .ZN(y[81]) );
  OR2_X1 U21bar ( .A1(abar[5]), .A2(bbar[1]), .ZN(ybar[81]) );
  AND2_X1 U22 ( .A1(a[5]), .A2(b[0]), .ZN(y[80]) );
  OR2_X1 U22bar ( .A1(abar[5]), .A2(bbar[0]), .ZN(ybar[80]) );
  AND2_X1 U23 ( .A1(b[7]), .A2(a[0]), .ZN(y[7]) );
  OR2_X1 U23bar ( .A1(bbar[7]), .A2(abar[0]), .ZN(ybar[7]) );
  AND2_X1 U24 ( .A1(a[4]), .A2(b[15]), .ZN(y[79]) );
  OR2_X1 U24bar ( .A1(abar[4]), .A2(bbar[15]), .ZN(ybar[79]) );
  AND2_X1 U25 ( .A1(a[4]), .A2(b[14]), .ZN(y[78]) );
  OR2_X1 U25bar ( .A1(abar[4]), .A2(bbar[14]), .ZN(ybar[78]) );
  AND2_X1 U26 ( .A1(a[4]), .A2(b[13]), .ZN(y[77]) );
  OR2_X1 U26bar ( .A1(abar[4]), .A2(bbar[13]), .ZN(ybar[77]) );
  AND2_X1 U27 ( .A1(a[4]), .A2(b[12]), .ZN(y[76]) );
  OR2_X1 U27bar ( .A1(abar[4]), .A2(bbar[12]), .ZN(ybar[76]) );
  AND2_X1 U28 ( .A1(a[4]), .A2(b[11]), .ZN(y[75]) );
  OR2_X1 U28bar ( .A1(abar[4]), .A2(bbar[11]), .ZN(ybar[75]) );
  AND2_X1 U29 ( .A1(a[4]), .A2(b[10]), .ZN(y[74]) );
  OR2_X1 U29bar ( .A1(abar[4]), .A2(bbar[10]), .ZN(ybar[74]) );
  AND2_X1 U30 ( .A1(a[4]), .A2(b[9]), .ZN(y[73]) );
  OR2_X1 U30bar ( .A1(abar[4]), .A2(bbar[9]), .ZN(ybar[73]) );
  AND2_X1 U31 ( .A1(a[4]), .A2(b[8]), .ZN(y[72]) );
  OR2_X1 U31bar ( .A1(abar[4]), .A2(bbar[8]), .ZN(ybar[72]) );
  AND2_X1 U32 ( .A1(a[4]), .A2(b[7]), .ZN(y[71]) );
  OR2_X1 U32bar ( .A1(abar[4]), .A2(bbar[7]), .ZN(ybar[71]) );
  AND2_X1 U33 ( .A1(a[4]), .A2(b[6]), .ZN(y[70]) );
  OR2_X1 U33bar ( .A1(abar[4]), .A2(bbar[6]), .ZN(ybar[70]) );
  AND2_X1 U34 ( .A1(b[6]), .A2(a[0]), .ZN(y[6]) );
  OR2_X1 U34bar ( .A1(bbar[6]), .A2(abar[0]), .ZN(ybar[6]) );
  AND2_X1 U35 ( .A1(a[4]), .A2(b[5]), .ZN(y[69]) );
  OR2_X1 U35bar ( .A1(abar[4]), .A2(bbar[5]), .ZN(ybar[69]) );
  AND2_X1 U36 ( .A1(a[4]), .A2(b[4]), .ZN(y[68]) );
  OR2_X1 U36bar ( .A1(abar[4]), .A2(bbar[4]), .ZN(ybar[68]) );
  AND2_X1 U37 ( .A1(a[4]), .A2(b[3]), .ZN(y[67]) );
  OR2_X1 U37bar ( .A1(abar[4]), .A2(bbar[3]), .ZN(ybar[67]) );
  AND2_X1 U38 ( .A1(a[4]), .A2(b[2]), .ZN(y[66]) );
  OR2_X1 U38bar ( .A1(abar[4]), .A2(bbar[2]), .ZN(ybar[66]) );
  AND2_X1 U39 ( .A1(a[4]), .A2(b[1]), .ZN(y[65]) );
  OR2_X1 U39bar ( .A1(abar[4]), .A2(bbar[1]), .ZN(ybar[65]) );
  AND2_X1 U40 ( .A1(a[4]), .A2(b[0]), .ZN(y[64]) );
  OR2_X1 U40bar ( .A1(abar[4]), .A2(bbar[0]), .ZN(ybar[64]) );
  AND2_X1 U41 ( .A1(a[3]), .A2(b[15]), .ZN(y[63]) );
  OR2_X1 U41bar ( .A1(abar[3]), .A2(bbar[15]), .ZN(ybar[63]) );
  AND2_X1 U42 ( .A1(a[3]), .A2(b[14]), .ZN(y[62]) );
  OR2_X1 U42bar ( .A1(abar[3]), .A2(bbar[14]), .ZN(ybar[62]) );
  AND2_X1 U43 ( .A1(a[3]), .A2(b[13]), .ZN(y[61]) );
  OR2_X1 U43bar ( .A1(abar[3]), .A2(bbar[13]), .ZN(ybar[61]) );
  AND2_X1 U44 ( .A1(a[3]), .A2(b[12]), .ZN(y[60]) );
  OR2_X1 U44bar ( .A1(abar[3]), .A2(bbar[12]), .ZN(ybar[60]) );
  AND2_X1 U45 ( .A1(b[5]), .A2(a[0]), .ZN(y[5]) );
  OR2_X1 U45bar ( .A1(bbar[5]), .A2(abar[0]), .ZN(ybar[5]) );
  AND2_X1 U46 ( .A1(a[3]), .A2(b[11]), .ZN(y[59]) );
  OR2_X1 U46bar ( .A1(abar[3]), .A2(bbar[11]), .ZN(ybar[59]) );
  AND2_X1 U47 ( .A1(a[3]), .A2(b[10]), .ZN(y[58]) );
  OR2_X1 U47bar ( .A1(abar[3]), .A2(bbar[10]), .ZN(ybar[58]) );
  AND2_X1 U48 ( .A1(a[3]), .A2(b[9]), .ZN(y[57]) );
  OR2_X1 U48bar ( .A1(abar[3]), .A2(bbar[9]), .ZN(ybar[57]) );
  AND2_X1 U49 ( .A1(a[3]), .A2(b[8]), .ZN(y[56]) );
  OR2_X1 U49bar ( .A1(abar[3]), .A2(bbar[8]), .ZN(ybar[56]) );
  AND2_X1 U50 ( .A1(a[3]), .A2(b[7]), .ZN(y[55]) );
  OR2_X1 U50bar ( .A1(abar[3]), .A2(bbar[7]), .ZN(ybar[55]) );
  AND2_X1 U51 ( .A1(a[3]), .A2(b[6]), .ZN(y[54]) );
  OR2_X1 U51bar ( .A1(abar[3]), .A2(bbar[6]), .ZN(ybar[54]) );
  AND2_X1 U52 ( .A1(a[3]), .A2(b[5]), .ZN(y[53]) );
  OR2_X1 U52bar ( .A1(abar[3]), .A2(bbar[5]), .ZN(ybar[53]) );
  AND2_X1 U53 ( .A1(a[3]), .A2(b[4]), .ZN(y[52]) );
  OR2_X1 U53bar ( .A1(abar[3]), .A2(bbar[4]), .ZN(ybar[52]) );
  AND2_X1 U54 ( .A1(a[3]), .A2(b[3]), .ZN(y[51]) );
  OR2_X1 U54bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[51]) );
  AND2_X1 U55 ( .A1(a[3]), .A2(b[2]), .ZN(y[50]) );
  OR2_X1 U55bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[50]) );
  AND2_X1 U56 ( .A1(b[4]), .A2(a[0]), .ZN(y[4]) );
  OR2_X1 U56bar ( .A1(bbar[4]), .A2(abar[0]), .ZN(ybar[4]) );
  AND2_X1 U57 ( .A1(a[3]), .A2(b[1]), .ZN(y[49]) );
  OR2_X1 U57bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[49]) );
  AND2_X1 U58 ( .A1(a[3]), .A2(b[0]), .ZN(y[48]) );
  OR2_X1 U58bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[48]) );
  AND2_X1 U59 ( .A1(a[2]), .A2(b[15]), .ZN(y[47]) );
  OR2_X1 U59bar ( .A1(abar[2]), .A2(bbar[15]), .ZN(ybar[47]) );
  AND2_X1 U60 ( .A1(a[2]), .A2(b[14]), .ZN(y[46]) );
  OR2_X1 U60bar ( .A1(abar[2]), .A2(bbar[14]), .ZN(ybar[46]) );
  AND2_X1 U61 ( .A1(a[2]), .A2(b[13]), .ZN(y[45]) );
  OR2_X1 U61bar ( .A1(abar[2]), .A2(bbar[13]), .ZN(ybar[45]) );
  AND2_X1 U62 ( .A1(a[2]), .A2(b[12]), .ZN(y[44]) );
  OR2_X1 U62bar ( .A1(abar[2]), .A2(bbar[12]), .ZN(ybar[44]) );
  AND2_X1 U63 ( .A1(a[2]), .A2(b[11]), .ZN(y[43]) );
  OR2_X1 U63bar ( .A1(abar[2]), .A2(bbar[11]), .ZN(ybar[43]) );
  AND2_X1 U64 ( .A1(a[2]), .A2(b[10]), .ZN(y[42]) );
  OR2_X1 U64bar ( .A1(abar[2]), .A2(bbar[10]), .ZN(ybar[42]) );
  AND2_X1 U65 ( .A1(a[2]), .A2(b[9]), .ZN(y[41]) );
  OR2_X1 U65bar ( .A1(abar[2]), .A2(bbar[9]), .ZN(ybar[41]) );
  AND2_X1 U66 ( .A1(a[2]), .A2(b[8]), .ZN(y[40]) );
  OR2_X1 U66bar ( .A1(abar[2]), .A2(bbar[8]), .ZN(ybar[40]) );
  AND2_X1 U67 ( .A1(b[3]), .A2(a[0]), .ZN(y[3]) );
  OR2_X1 U67bar ( .A1(bbar[3]), .A2(abar[0]), .ZN(ybar[3]) );
  AND2_X1 U68 ( .A1(a[2]), .A2(b[7]), .ZN(y[39]) );
  OR2_X1 U68bar ( .A1(abar[2]), .A2(bbar[7]), .ZN(ybar[39]) );
  AND2_X1 U69 ( .A1(a[2]), .A2(b[6]), .ZN(y[38]) );
  OR2_X1 U69bar ( .A1(abar[2]), .A2(bbar[6]), .ZN(ybar[38]) );
  AND2_X1 U70 ( .A1(a[2]), .A2(b[5]), .ZN(y[37]) );
  OR2_X1 U70bar ( .A1(abar[2]), .A2(bbar[5]), .ZN(ybar[37]) );
  AND2_X1 U71 ( .A1(a[2]), .A2(b[4]), .ZN(y[36]) );
  OR2_X1 U71bar ( .A1(abar[2]), .A2(bbar[4]), .ZN(ybar[36]) );
  AND2_X1 U72 ( .A1(a[2]), .A2(b[3]), .ZN(y[35]) );
  OR2_X1 U72bar ( .A1(abar[2]), .A2(bbar[3]), .ZN(ybar[35]) );
  AND2_X1 U73 ( .A1(a[2]), .A2(b[2]), .ZN(y[34]) );
  OR2_X1 U73bar ( .A1(abar[2]), .A2(bbar[2]), .ZN(ybar[34]) );
  AND2_X1 U74 ( .A1(a[2]), .A2(b[1]), .ZN(y[33]) );
  OR2_X1 U74bar ( .A1(abar[2]), .A2(bbar[1]), .ZN(ybar[33]) );
  AND2_X1 U75 ( .A1(a[2]), .A2(b[0]), .ZN(y[32]) );
  OR2_X1 U75bar ( .A1(abar[2]), .A2(bbar[0]), .ZN(ybar[32]) );
  AND2_X1 U76 ( .A1(a[1]), .A2(b[15]), .ZN(y[31]) );
  OR2_X1 U76bar ( .A1(abar[1]), .A2(bbar[15]), .ZN(ybar[31]) );
  AND2_X1 U77 ( .A1(a[1]), .A2(b[14]), .ZN(y[30]) );
  OR2_X1 U77bar ( .A1(abar[1]), .A2(bbar[14]), .ZN(ybar[30]) );
  AND2_X1 U78 ( .A1(b[2]), .A2(a[0]), .ZN(y[2]) );
  OR2_X1 U78bar ( .A1(bbar[2]), .A2(abar[0]), .ZN(ybar[2]) );
  AND2_X1 U79 ( .A1(a[1]), .A2(b[13]), .ZN(y[29]) );
  OR2_X1 U79bar ( .A1(abar[1]), .A2(bbar[13]), .ZN(ybar[29]) );
  AND2_X1 U80 ( .A1(a[1]), .A2(b[12]), .ZN(y[28]) );
  OR2_X1 U80bar ( .A1(abar[1]), .A2(bbar[12]), .ZN(ybar[28]) );
  AND2_X1 U81 ( .A1(a[1]), .A2(b[11]), .ZN(y[27]) );
  OR2_X1 U81bar ( .A1(abar[1]), .A2(bbar[11]), .ZN(ybar[27]) );
  AND2_X1 U82 ( .A1(a[1]), .A2(b[10]), .ZN(y[26]) );
  OR2_X1 U82bar ( .A1(abar[1]), .A2(bbar[10]), .ZN(ybar[26]) );
  AND2_X1 U83 ( .A1(a[1]), .A2(b[9]), .ZN(y[25]) );
  OR2_X1 U83bar ( .A1(abar[1]), .A2(bbar[9]), .ZN(ybar[25]) );
  AND2_X1 U84 ( .A1(a[15]), .A2(b[15]), .ZN(y[255]) );
  OR2_X1 U84bar ( .A1(abar[15]), .A2(bbar[15]), .ZN(ybar[255]) );
  AND2_X1 U85 ( .A1(a[15]), .A2(b[14]), .ZN(y[254]) );
  OR2_X1 U85bar ( .A1(abar[15]), .A2(bbar[14]), .ZN(ybar[254]) );
  AND2_X1 U86 ( .A1(a[15]), .A2(b[13]), .ZN(y[253]) );
  OR2_X1 U86bar ( .A1(abar[15]), .A2(bbar[13]), .ZN(ybar[253]) );
  AND2_X1 U87 ( .A1(a[15]), .A2(b[12]), .ZN(y[252]) );
  OR2_X1 U87bar ( .A1(abar[15]), .A2(bbar[12]), .ZN(ybar[252]) );
  AND2_X1 U88 ( .A1(a[15]), .A2(b[11]), .ZN(y[251]) );
  OR2_X1 U88bar ( .A1(abar[15]), .A2(bbar[11]), .ZN(ybar[251]) );
  AND2_X1 U89 ( .A1(a[15]), .A2(b[10]), .ZN(y[250]) );
  OR2_X1 U89bar ( .A1(abar[15]), .A2(bbar[10]), .ZN(ybar[250]) );
  AND2_X1 U90 ( .A1(a[1]), .A2(b[8]), .ZN(y[24]) );
  OR2_X1 U90bar ( .A1(abar[1]), .A2(bbar[8]), .ZN(ybar[24]) );
  AND2_X1 U91 ( .A1(a[15]), .A2(b[9]), .ZN(y[249]) );
  OR2_X1 U91bar ( .A1(abar[15]), .A2(bbar[9]), .ZN(ybar[249]) );
  AND2_X1 U92 ( .A1(a[15]), .A2(b[8]), .ZN(y[248]) );
  OR2_X1 U92bar ( .A1(abar[15]), .A2(bbar[8]), .ZN(ybar[248]) );
  AND2_X1 U93 ( .A1(a[15]), .A2(b[7]), .ZN(y[247]) );
  OR2_X1 U93bar ( .A1(abar[15]), .A2(bbar[7]), .ZN(ybar[247]) );
  AND2_X1 U94 ( .A1(a[15]), .A2(b[6]), .ZN(y[246]) );
  OR2_X1 U94bar ( .A1(abar[15]), .A2(bbar[6]), .ZN(ybar[246]) );
  AND2_X1 U95 ( .A1(a[15]), .A2(b[5]), .ZN(y[245]) );
  OR2_X1 U95bar ( .A1(abar[15]), .A2(bbar[5]), .ZN(ybar[245]) );
  AND2_X1 U96 ( .A1(a[15]), .A2(b[4]), .ZN(y[244]) );
  OR2_X1 U96bar ( .A1(abar[15]), .A2(bbar[4]), .ZN(ybar[244]) );
  AND2_X1 U97 ( .A1(a[15]), .A2(b[3]), .ZN(y[243]) );
  OR2_X1 U97bar ( .A1(abar[15]), .A2(bbar[3]), .ZN(ybar[243]) );
  AND2_X1 U98 ( .A1(a[15]), .A2(b[2]), .ZN(y[242]) );
  OR2_X1 U98bar ( .A1(abar[15]), .A2(bbar[2]), .ZN(ybar[242]) );
  AND2_X1 U99 ( .A1(a[15]), .A2(b[1]), .ZN(y[241]) );
  OR2_X1 U99bar ( .A1(abar[15]), .A2(bbar[1]), .ZN(ybar[241]) );
  AND2_X1 U100 ( .A1(a[15]), .A2(b[0]), .ZN(y[240]) );
  OR2_X1 U100bar ( .A1(abar[15]), .A2(bbar[0]), .ZN(ybar[240]) );
  AND2_X1 U101 ( .A1(a[1]), .A2(b[7]), .ZN(y[23]) );
  OR2_X1 U101bar ( .A1(abar[1]), .A2(bbar[7]), .ZN(ybar[23]) );
  AND2_X1 U102 ( .A1(a[14]), .A2(b[15]), .ZN(y[239]) );
  OR2_X1 U102bar ( .A1(abar[14]), .A2(bbar[15]), .ZN(ybar[239]) );
  AND2_X1 U103 ( .A1(a[14]), .A2(b[14]), .ZN(y[238]) );
  OR2_X1 U103bar ( .A1(abar[14]), .A2(bbar[14]), .ZN(ybar[238]) );
  AND2_X1 U104 ( .A1(a[14]), .A2(b[13]), .ZN(y[237]) );
  OR2_X1 U104bar ( .A1(abar[14]), .A2(bbar[13]), .ZN(ybar[237]) );
  AND2_X1 U105 ( .A1(a[14]), .A2(b[12]), .ZN(y[236]) );
  OR2_X1 U105bar ( .A1(abar[14]), .A2(bbar[12]), .ZN(ybar[236]) );
  AND2_X1 U106 ( .A1(a[14]), .A2(b[11]), .ZN(y[235]) );
  OR2_X1 U106bar ( .A1(abar[14]), .A2(bbar[11]), .ZN(ybar[235]) );
  AND2_X1 U107 ( .A1(a[14]), .A2(b[10]), .ZN(y[234]) );
  OR2_X1 U107bar ( .A1(abar[14]), .A2(bbar[10]), .ZN(ybar[234]) );
  AND2_X1 U108 ( .A1(a[14]), .A2(b[9]), .ZN(y[233]) );
  OR2_X1 U108bar ( .A1(abar[14]), .A2(bbar[9]), .ZN(ybar[233]) );
  AND2_X1 U109 ( .A1(a[14]), .A2(b[8]), .ZN(y[232]) );
  OR2_X1 U109bar ( .A1(abar[14]), .A2(bbar[8]), .ZN(ybar[232]) );
  AND2_X1 U110 ( .A1(a[14]), .A2(b[7]), .ZN(y[231]) );
  OR2_X1 U110bar ( .A1(abar[14]), .A2(bbar[7]), .ZN(ybar[231]) );
  AND2_X1 U111 ( .A1(a[14]), .A2(b[6]), .ZN(y[230]) );
  OR2_X1 U111bar ( .A1(abar[14]), .A2(bbar[6]), .ZN(ybar[230]) );
  AND2_X1 U112 ( .A1(a[1]), .A2(b[6]), .ZN(y[22]) );
  OR2_X1 U112bar ( .A1(abar[1]), .A2(bbar[6]), .ZN(ybar[22]) );
  AND2_X1 U113 ( .A1(a[14]), .A2(b[5]), .ZN(y[229]) );
  OR2_X1 U113bar ( .A1(abar[14]), .A2(bbar[5]), .ZN(ybar[229]) );
  AND2_X1 U114 ( .A1(a[14]), .A2(b[4]), .ZN(y[228]) );
  OR2_X1 U114bar ( .A1(abar[14]), .A2(bbar[4]), .ZN(ybar[228]) );
  AND2_X1 U115 ( .A1(a[14]), .A2(b[3]), .ZN(y[227]) );
  OR2_X1 U115bar ( .A1(abar[14]), .A2(bbar[3]), .ZN(ybar[227]) );
  AND2_X1 U116 ( .A1(a[14]), .A2(b[2]), .ZN(y[226]) );
  OR2_X1 U116bar ( .A1(abar[14]), .A2(bbar[2]), .ZN(ybar[226]) );
  AND2_X1 U117 ( .A1(a[14]), .A2(b[1]), .ZN(y[225]) );
  OR2_X1 U117bar ( .A1(abar[14]), .A2(bbar[1]), .ZN(ybar[225]) );
  AND2_X1 U118 ( .A1(a[14]), .A2(b[0]), .ZN(y[224]) );
  OR2_X1 U118bar ( .A1(abar[14]), .A2(bbar[0]), .ZN(ybar[224]) );
  AND2_X1 U119 ( .A1(a[13]), .A2(b[15]), .ZN(y[223]) );
  OR2_X1 U119bar ( .A1(abar[13]), .A2(bbar[15]), .ZN(ybar[223]) );
  AND2_X1 U120 ( .A1(a[13]), .A2(b[14]), .ZN(y[222]) );
  OR2_X1 U120bar ( .A1(abar[13]), .A2(bbar[14]), .ZN(ybar[222]) );
  AND2_X1 U121 ( .A1(a[13]), .A2(b[13]), .ZN(y[221]) );
  OR2_X1 U121bar ( .A1(abar[13]), .A2(bbar[13]), .ZN(ybar[221]) );
  AND2_X1 U122 ( .A1(a[13]), .A2(b[12]), .ZN(y[220]) );
  OR2_X1 U122bar ( .A1(abar[13]), .A2(bbar[12]), .ZN(ybar[220]) );
  AND2_X1 U123 ( .A1(a[1]), .A2(b[5]), .ZN(y[21]) );
  OR2_X1 U123bar ( .A1(abar[1]), .A2(bbar[5]), .ZN(ybar[21]) );
  AND2_X1 U124 ( .A1(a[13]), .A2(b[11]), .ZN(y[219]) );
  OR2_X1 U124bar ( .A1(abar[13]), .A2(bbar[11]), .ZN(ybar[219]) );
  AND2_X1 U125 ( .A1(a[13]), .A2(b[10]), .ZN(y[218]) );
  OR2_X1 U125bar ( .A1(abar[13]), .A2(bbar[10]), .ZN(ybar[218]) );
  AND2_X1 U126 ( .A1(a[13]), .A2(b[9]), .ZN(y[217]) );
  OR2_X1 U126bar ( .A1(abar[13]), .A2(bbar[9]), .ZN(ybar[217]) );
  AND2_X1 U127 ( .A1(a[13]), .A2(b[8]), .ZN(y[216]) );
  OR2_X1 U127bar ( .A1(abar[13]), .A2(bbar[8]), .ZN(ybar[216]) );
  AND2_X1 U128 ( .A1(a[13]), .A2(b[7]), .ZN(y[215]) );
  OR2_X1 U128bar ( .A1(abar[13]), .A2(bbar[7]), .ZN(ybar[215]) );
  AND2_X1 U129 ( .A1(a[13]), .A2(b[6]), .ZN(y[214]) );
  OR2_X1 U129bar ( .A1(abar[13]), .A2(bbar[6]), .ZN(ybar[214]) );
  AND2_X1 U130 ( .A1(a[13]), .A2(b[5]), .ZN(y[213]) );
  OR2_X1 U130bar ( .A1(abar[13]), .A2(bbar[5]), .ZN(ybar[213]) );
  AND2_X1 U131 ( .A1(a[13]), .A2(b[4]), .ZN(y[212]) );
  OR2_X1 U131bar ( .A1(abar[13]), .A2(bbar[4]), .ZN(ybar[212]) );
  AND2_X1 U132 ( .A1(a[13]), .A2(b[3]), .ZN(y[211]) );
  OR2_X1 U132bar ( .A1(abar[13]), .A2(bbar[3]), .ZN(ybar[211]) );
  AND2_X1 U133 ( .A1(a[13]), .A2(b[2]), .ZN(y[210]) );
  OR2_X1 U133bar ( .A1(abar[13]), .A2(bbar[2]), .ZN(ybar[210]) );
  AND2_X1 U134 ( .A1(a[1]), .A2(b[4]), .ZN(y[20]) );
  OR2_X1 U134bar ( .A1(abar[1]), .A2(bbar[4]), .ZN(ybar[20]) );
  AND2_X1 U135 ( .A1(a[13]), .A2(b[1]), .ZN(y[209]) );
  OR2_X1 U135bar ( .A1(abar[13]), .A2(bbar[1]), .ZN(ybar[209]) );
  AND2_X1 U136 ( .A1(a[13]), .A2(b[0]), .ZN(y[208]) );
  OR2_X1 U136bar ( .A1(abar[13]), .A2(bbar[0]), .ZN(ybar[208]) );
  AND2_X1 U137 ( .A1(a[12]), .A2(b[15]), .ZN(y[207]) );
  OR2_X1 U137bar ( .A1(abar[12]), .A2(bbar[15]), .ZN(ybar[207]) );
  AND2_X1 U138 ( .A1(a[12]), .A2(b[14]), .ZN(y[206]) );
  OR2_X1 U138bar ( .A1(abar[12]), .A2(bbar[14]), .ZN(ybar[206]) );
  AND2_X1 U139 ( .A1(a[12]), .A2(b[13]), .ZN(y[205]) );
  OR2_X1 U139bar ( .A1(abar[12]), .A2(bbar[13]), .ZN(ybar[205]) );
  AND2_X1 U140 ( .A1(a[12]), .A2(b[12]), .ZN(y[204]) );
  OR2_X1 U140bar ( .A1(abar[12]), .A2(bbar[12]), .ZN(ybar[204]) );
  AND2_X1 U141 ( .A1(a[12]), .A2(b[11]), .ZN(y[203]) );
  OR2_X1 U141bar ( .A1(abar[12]), .A2(bbar[11]), .ZN(ybar[203]) );
  AND2_X1 U142 ( .A1(a[12]), .A2(b[10]), .ZN(y[202]) );
  OR2_X1 U142bar ( .A1(abar[12]), .A2(bbar[10]), .ZN(ybar[202]) );
  AND2_X1 U143 ( .A1(a[12]), .A2(b[9]), .ZN(y[201]) );
  OR2_X1 U143bar ( .A1(abar[12]), .A2(bbar[9]), .ZN(ybar[201]) );
  AND2_X1 U144 ( .A1(a[12]), .A2(b[8]), .ZN(y[200]) );
  OR2_X1 U144bar ( .A1(abar[12]), .A2(bbar[8]), .ZN(ybar[200]) );
  AND2_X1 U145 ( .A1(b[1]), .A2(a[0]), .ZN(y[1]) );
  OR2_X1 U145bar ( .A1(bbar[1]), .A2(abar[0]), .ZN(ybar[1]) );
  AND2_X1 U146 ( .A1(a[1]), .A2(b[3]), .ZN(y[19]) );
  OR2_X1 U146bar ( .A1(abar[1]), .A2(bbar[3]), .ZN(ybar[19]) );
  AND2_X1 U147 ( .A1(a[12]), .A2(b[7]), .ZN(y[199]) );
  OR2_X1 U147bar ( .A1(abar[12]), .A2(bbar[7]), .ZN(ybar[199]) );
  AND2_X1 U148 ( .A1(a[12]), .A2(b[6]), .ZN(y[198]) );
  OR2_X1 U148bar ( .A1(abar[12]), .A2(bbar[6]), .ZN(ybar[198]) );
  AND2_X1 U149 ( .A1(a[12]), .A2(b[5]), .ZN(y[197]) );
  OR2_X1 U149bar ( .A1(abar[12]), .A2(bbar[5]), .ZN(ybar[197]) );
  AND2_X1 U150 ( .A1(a[12]), .A2(b[4]), .ZN(y[196]) );
  OR2_X1 U150bar ( .A1(abar[12]), .A2(bbar[4]), .ZN(ybar[196]) );
  AND2_X1 U151 ( .A1(a[12]), .A2(b[3]), .ZN(y[195]) );
  OR2_X1 U151bar ( .A1(abar[12]), .A2(bbar[3]), .ZN(ybar[195]) );
  AND2_X1 U152 ( .A1(a[12]), .A2(b[2]), .ZN(y[194]) );
  OR2_X1 U152bar ( .A1(abar[12]), .A2(bbar[2]), .ZN(ybar[194]) );
  AND2_X1 U153 ( .A1(a[12]), .A2(b[1]), .ZN(y[193]) );
  OR2_X1 U153bar ( .A1(abar[12]), .A2(bbar[1]), .ZN(ybar[193]) );
  AND2_X1 U154 ( .A1(a[12]), .A2(b[0]), .ZN(y[192]) );
  OR2_X1 U154bar ( .A1(abar[12]), .A2(bbar[0]), .ZN(ybar[192]) );
  AND2_X1 U155 ( .A1(a[11]), .A2(b[15]), .ZN(y[191]) );
  OR2_X1 U155bar ( .A1(abar[11]), .A2(bbar[15]), .ZN(ybar[191]) );
  AND2_X1 U156 ( .A1(a[11]), .A2(b[14]), .ZN(y[190]) );
  OR2_X1 U156bar ( .A1(abar[11]), .A2(bbar[14]), .ZN(ybar[190]) );
  AND2_X1 U157 ( .A1(a[1]), .A2(b[2]), .ZN(y[18]) );
  OR2_X1 U157bar ( .A1(abar[1]), .A2(bbar[2]), .ZN(ybar[18]) );
  AND2_X1 U158 ( .A1(a[11]), .A2(b[13]), .ZN(y[189]) );
  OR2_X1 U158bar ( .A1(abar[11]), .A2(bbar[13]), .ZN(ybar[189]) );
  AND2_X1 U159 ( .A1(a[11]), .A2(b[12]), .ZN(y[188]) );
  OR2_X1 U159bar ( .A1(abar[11]), .A2(bbar[12]), .ZN(ybar[188]) );
  AND2_X1 U160 ( .A1(a[11]), .A2(b[11]), .ZN(y[187]) );
  OR2_X1 U160bar ( .A1(abar[11]), .A2(bbar[11]), .ZN(ybar[187]) );
  AND2_X1 U161 ( .A1(a[11]), .A2(b[10]), .ZN(y[186]) );
  OR2_X1 U161bar ( .A1(abar[11]), .A2(bbar[10]), .ZN(ybar[186]) );
  AND2_X1 U162 ( .A1(a[11]), .A2(b[9]), .ZN(y[185]) );
  OR2_X1 U162bar ( .A1(abar[11]), .A2(bbar[9]), .ZN(ybar[185]) );
  AND2_X1 U163 ( .A1(a[11]), .A2(b[8]), .ZN(y[184]) );
  OR2_X1 U163bar ( .A1(abar[11]), .A2(bbar[8]), .ZN(ybar[184]) );
  AND2_X1 U164 ( .A1(a[11]), .A2(b[7]), .ZN(y[183]) );
  OR2_X1 U164bar ( .A1(abar[11]), .A2(bbar[7]), .ZN(ybar[183]) );
  AND2_X1 U165 ( .A1(a[11]), .A2(b[6]), .ZN(y[182]) );
  OR2_X1 U165bar ( .A1(abar[11]), .A2(bbar[6]), .ZN(ybar[182]) );
  AND2_X1 U166 ( .A1(a[11]), .A2(b[5]), .ZN(y[181]) );
  OR2_X1 U166bar ( .A1(abar[11]), .A2(bbar[5]), .ZN(ybar[181]) );
  AND2_X1 U167 ( .A1(a[11]), .A2(b[4]), .ZN(y[180]) );
  OR2_X1 U167bar ( .A1(abar[11]), .A2(bbar[4]), .ZN(ybar[180]) );
  AND2_X1 U168 ( .A1(a[1]), .A2(b[1]), .ZN(y[17]) );
  OR2_X1 U168bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[17]) );
  AND2_X1 U169 ( .A1(a[11]), .A2(b[3]), .ZN(y[179]) );
  OR2_X1 U169bar ( .A1(abar[11]), .A2(bbar[3]), .ZN(ybar[179]) );
  AND2_X1 U170 ( .A1(a[11]), .A2(b[2]), .ZN(y[178]) );
  OR2_X1 U170bar ( .A1(abar[11]), .A2(bbar[2]), .ZN(ybar[178]) );
  AND2_X1 U171 ( .A1(a[11]), .A2(b[1]), .ZN(y[177]) );
  OR2_X1 U171bar ( .A1(abar[11]), .A2(bbar[1]), .ZN(ybar[177]) );
  AND2_X1 U172 ( .A1(a[11]), .A2(b[0]), .ZN(y[176]) );
  OR2_X1 U172bar ( .A1(abar[11]), .A2(bbar[0]), .ZN(ybar[176]) );
  AND2_X1 U173 ( .A1(a[10]), .A2(b[15]), .ZN(y[175]) );
  OR2_X1 U173bar ( .A1(abar[10]), .A2(bbar[15]), .ZN(ybar[175]) );
  AND2_X1 U174 ( .A1(a[10]), .A2(b[14]), .ZN(y[174]) );
  OR2_X1 U174bar ( .A1(abar[10]), .A2(bbar[14]), .ZN(ybar[174]) );
  AND2_X1 U175 ( .A1(a[10]), .A2(b[13]), .ZN(y[173]) );
  OR2_X1 U175bar ( .A1(abar[10]), .A2(bbar[13]), .ZN(ybar[173]) );
  AND2_X1 U176 ( .A1(a[10]), .A2(b[12]), .ZN(y[172]) );
  OR2_X1 U176bar ( .A1(abar[10]), .A2(bbar[12]), .ZN(ybar[172]) );
  AND2_X1 U177 ( .A1(a[10]), .A2(b[11]), .ZN(y[171]) );
  OR2_X1 U177bar ( .A1(abar[10]), .A2(bbar[11]), .ZN(ybar[171]) );
  AND2_X1 U178 ( .A1(a[10]), .A2(b[10]), .ZN(y[170]) );
  OR2_X1 U178bar ( .A1(abar[10]), .A2(bbar[10]), .ZN(ybar[170]) );
  AND2_X1 U179 ( .A1(a[1]), .A2(b[0]), .ZN(y[16]) );
  OR2_X1 U179bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[16]) );
  AND2_X1 U180 ( .A1(a[10]), .A2(b[9]), .ZN(y[169]) );
  OR2_X1 U180bar ( .A1(abar[10]), .A2(bbar[9]), .ZN(ybar[169]) );
  AND2_X1 U181 ( .A1(a[10]), .A2(b[8]), .ZN(y[168]) );
  OR2_X1 U181bar ( .A1(abar[10]), .A2(bbar[8]), .ZN(ybar[168]) );
  AND2_X1 U182 ( .A1(a[10]), .A2(b[7]), .ZN(y[167]) );
  OR2_X1 U182bar ( .A1(abar[10]), .A2(bbar[7]), .ZN(ybar[167]) );
  AND2_X1 U183 ( .A1(a[10]), .A2(b[6]), .ZN(y[166]) );
  OR2_X1 U183bar ( .A1(abar[10]), .A2(bbar[6]), .ZN(ybar[166]) );
  AND2_X1 U184 ( .A1(a[10]), .A2(b[5]), .ZN(y[165]) );
  OR2_X1 U184bar ( .A1(abar[10]), .A2(bbar[5]), .ZN(ybar[165]) );
  AND2_X1 U185 ( .A1(a[10]), .A2(b[4]), .ZN(y[164]) );
  OR2_X1 U185bar ( .A1(abar[10]), .A2(bbar[4]), .ZN(ybar[164]) );
  AND2_X1 U186 ( .A1(a[10]), .A2(b[3]), .ZN(y[163]) );
  OR2_X1 U186bar ( .A1(abar[10]), .A2(bbar[3]), .ZN(ybar[163]) );
  AND2_X1 U187 ( .A1(a[10]), .A2(b[2]), .ZN(y[162]) );
  OR2_X1 U187bar ( .A1(abar[10]), .A2(bbar[2]), .ZN(ybar[162]) );
  AND2_X1 U188 ( .A1(a[10]), .A2(b[1]), .ZN(y[161]) );
  OR2_X1 U188bar ( .A1(abar[10]), .A2(bbar[1]), .ZN(ybar[161]) );
  AND2_X1 U189 ( .A1(a[10]), .A2(b[0]), .ZN(y[160]) );
  OR2_X1 U189bar ( .A1(abar[10]), .A2(bbar[0]), .ZN(ybar[160]) );
  AND2_X1 U190 ( .A1(b[15]), .A2(a[0]), .ZN(y[15]) );
  OR2_X1 U190bar ( .A1(bbar[15]), .A2(abar[0]), .ZN(ybar[15]) );
  AND2_X1 U191 ( .A1(a[9]), .A2(b[15]), .ZN(y[159]) );
  OR2_X1 U191bar ( .A1(abar[9]), .A2(bbar[15]), .ZN(ybar[159]) );
  AND2_X1 U192 ( .A1(a[9]), .A2(b[14]), .ZN(y[158]) );
  OR2_X1 U192bar ( .A1(abar[9]), .A2(bbar[14]), .ZN(ybar[158]) );
  AND2_X1 U193 ( .A1(a[9]), .A2(b[13]), .ZN(y[157]) );
  OR2_X1 U193bar ( .A1(abar[9]), .A2(bbar[13]), .ZN(ybar[157]) );
  AND2_X1 U194 ( .A1(a[9]), .A2(b[12]), .ZN(y[156]) );
  OR2_X1 U194bar ( .A1(abar[9]), .A2(bbar[12]), .ZN(ybar[156]) );
  AND2_X1 U195 ( .A1(a[9]), .A2(b[11]), .ZN(y[155]) );
  OR2_X1 U195bar ( .A1(abar[9]), .A2(bbar[11]), .ZN(ybar[155]) );
  AND2_X1 U196 ( .A1(a[9]), .A2(b[10]), .ZN(y[154]) );
  OR2_X1 U196bar ( .A1(abar[9]), .A2(bbar[10]), .ZN(ybar[154]) );
  AND2_X1 U197 ( .A1(a[9]), .A2(b[9]), .ZN(y[153]) );
  OR2_X1 U197bar ( .A1(abar[9]), .A2(bbar[9]), .ZN(ybar[153]) );
  AND2_X1 U198 ( .A1(a[9]), .A2(b[8]), .ZN(y[152]) );
  OR2_X1 U198bar ( .A1(abar[9]), .A2(bbar[8]), .ZN(ybar[152]) );
  AND2_X1 U199 ( .A1(a[9]), .A2(b[7]), .ZN(y[151]) );
  OR2_X1 U199bar ( .A1(abar[9]), .A2(bbar[7]), .ZN(ybar[151]) );
  AND2_X1 U200 ( .A1(a[9]), .A2(b[6]), .ZN(y[150]) );
  OR2_X1 U200bar ( .A1(abar[9]), .A2(bbar[6]), .ZN(ybar[150]) );
  AND2_X1 U201 ( .A1(b[14]), .A2(a[0]), .ZN(y[14]) );
  OR2_X1 U201bar ( .A1(bbar[14]), .A2(abar[0]), .ZN(ybar[14]) );
  AND2_X1 U202 ( .A1(a[9]), .A2(b[5]), .ZN(y[149]) );
  OR2_X1 U202bar ( .A1(abar[9]), .A2(bbar[5]), .ZN(ybar[149]) );
  AND2_X1 U203 ( .A1(a[9]), .A2(b[4]), .ZN(y[148]) );
  OR2_X1 U203bar ( .A1(abar[9]), .A2(bbar[4]), .ZN(ybar[148]) );
  AND2_X1 U204 ( .A1(a[9]), .A2(b[3]), .ZN(y[147]) );
  OR2_X1 U204bar ( .A1(abar[9]), .A2(bbar[3]), .ZN(ybar[147]) );
  AND2_X1 U205 ( .A1(a[9]), .A2(b[2]), .ZN(y[146]) );
  OR2_X1 U205bar ( .A1(abar[9]), .A2(bbar[2]), .ZN(ybar[146]) );
  AND2_X1 U206 ( .A1(a[9]), .A2(b[1]), .ZN(y[145]) );
  OR2_X1 U206bar ( .A1(abar[9]), .A2(bbar[1]), .ZN(ybar[145]) );
  AND2_X1 U207 ( .A1(a[9]), .A2(b[0]), .ZN(y[144]) );
  OR2_X1 U207bar ( .A1(abar[9]), .A2(bbar[0]), .ZN(ybar[144]) );
  AND2_X1 U208 ( .A1(a[8]), .A2(b[15]), .ZN(y[143]) );
  OR2_X1 U208bar ( .A1(abar[8]), .A2(bbar[15]), .ZN(ybar[143]) );
  AND2_X1 U209 ( .A1(a[8]), .A2(b[14]), .ZN(y[142]) );
  OR2_X1 U209bar ( .A1(abar[8]), .A2(bbar[14]), .ZN(ybar[142]) );
  AND2_X1 U210 ( .A1(a[8]), .A2(b[13]), .ZN(y[141]) );
  OR2_X1 U210bar ( .A1(abar[8]), .A2(bbar[13]), .ZN(ybar[141]) );
  AND2_X1 U211 ( .A1(a[8]), .A2(b[12]), .ZN(y[140]) );
  OR2_X1 U211bar ( .A1(abar[8]), .A2(bbar[12]), .ZN(ybar[140]) );
  AND2_X1 U212 ( .A1(b[13]), .A2(a[0]), .ZN(y[13]) );
  OR2_X1 U212bar ( .A1(bbar[13]), .A2(abar[0]), .ZN(ybar[13]) );
  AND2_X1 U213 ( .A1(a[8]), .A2(b[11]), .ZN(y[139]) );
  OR2_X1 U213bar ( .A1(abar[8]), .A2(bbar[11]), .ZN(ybar[139]) );
  AND2_X1 U214 ( .A1(a[8]), .A2(b[10]), .ZN(y[138]) );
  OR2_X1 U214bar ( .A1(abar[8]), .A2(bbar[10]), .ZN(ybar[138]) );
  AND2_X1 U215 ( .A1(a[8]), .A2(b[9]), .ZN(y[137]) );
  OR2_X1 U215bar ( .A1(abar[8]), .A2(bbar[9]), .ZN(ybar[137]) );
  AND2_X1 U216 ( .A1(a[8]), .A2(b[8]), .ZN(y[136]) );
  OR2_X1 U216bar ( .A1(abar[8]), .A2(bbar[8]), .ZN(ybar[136]) );
  AND2_X1 U217 ( .A1(a[8]), .A2(b[7]), .ZN(y[135]) );
  OR2_X1 U217bar ( .A1(abar[8]), .A2(bbar[7]), .ZN(ybar[135]) );
  AND2_X1 U218 ( .A1(a[8]), .A2(b[6]), .ZN(y[134]) );
  OR2_X1 U218bar ( .A1(abar[8]), .A2(bbar[6]), .ZN(ybar[134]) );
  AND2_X1 U219 ( .A1(a[8]), .A2(b[5]), .ZN(y[133]) );
  OR2_X1 U219bar ( .A1(abar[8]), .A2(bbar[5]), .ZN(ybar[133]) );
  AND2_X1 U220 ( .A1(a[8]), .A2(b[4]), .ZN(y[132]) );
  OR2_X1 U220bar ( .A1(abar[8]), .A2(bbar[4]), .ZN(ybar[132]) );
  AND2_X1 U221 ( .A1(a[8]), .A2(b[3]), .ZN(y[131]) );
  OR2_X1 U221bar ( .A1(abar[8]), .A2(bbar[3]), .ZN(ybar[131]) );
  AND2_X1 U222 ( .A1(a[8]), .A2(b[2]), .ZN(y[130]) );
  OR2_X1 U222bar ( .A1(abar[8]), .A2(bbar[2]), .ZN(ybar[130]) );
  AND2_X1 U223 ( .A1(b[12]), .A2(a[0]), .ZN(y[12]) );
  OR2_X1 U223bar ( .A1(bbar[12]), .A2(abar[0]), .ZN(ybar[12]) );
  AND2_X1 U224 ( .A1(a[8]), .A2(b[1]), .ZN(y[129]) );
  OR2_X1 U224bar ( .A1(abar[8]), .A2(bbar[1]), .ZN(ybar[129]) );
  AND2_X1 U225 ( .A1(a[8]), .A2(b[0]), .ZN(y[128]) );
  OR2_X1 U225bar ( .A1(abar[8]), .A2(bbar[0]), .ZN(ybar[128]) );
  AND2_X1 U226 ( .A1(a[7]), .A2(b[15]), .ZN(y[127]) );
  OR2_X1 U226bar ( .A1(abar[7]), .A2(bbar[15]), .ZN(ybar[127]) );
  AND2_X1 U227 ( .A1(a[7]), .A2(b[14]), .ZN(y[126]) );
  OR2_X1 U227bar ( .A1(abar[7]), .A2(bbar[14]), .ZN(ybar[126]) );
  AND2_X1 U228 ( .A1(a[7]), .A2(b[13]), .ZN(y[125]) );
  OR2_X1 U228bar ( .A1(abar[7]), .A2(bbar[13]), .ZN(ybar[125]) );
  AND2_X1 U229 ( .A1(a[7]), .A2(b[12]), .ZN(y[124]) );
  OR2_X1 U229bar ( .A1(abar[7]), .A2(bbar[12]), .ZN(ybar[124]) );
  AND2_X1 U230 ( .A1(a[7]), .A2(b[11]), .ZN(y[123]) );
  OR2_X1 U230bar ( .A1(abar[7]), .A2(bbar[11]), .ZN(ybar[123]) );
  AND2_X1 U231 ( .A1(a[7]), .A2(b[10]), .ZN(y[122]) );
  OR2_X1 U231bar ( .A1(abar[7]), .A2(bbar[10]), .ZN(ybar[122]) );
  AND2_X1 U232 ( .A1(a[7]), .A2(b[9]), .ZN(y[121]) );
  OR2_X1 U232bar ( .A1(abar[7]), .A2(bbar[9]), .ZN(ybar[121]) );
  AND2_X1 U233 ( .A1(a[7]), .A2(b[8]), .ZN(y[120]) );
  OR2_X1 U233bar ( .A1(abar[7]), .A2(bbar[8]), .ZN(ybar[120]) );
  AND2_X1 U234 ( .A1(b[11]), .A2(a[0]), .ZN(y[11]) );
  OR2_X1 U234bar ( .A1(bbar[11]), .A2(abar[0]), .ZN(ybar[11]) );
  AND2_X1 U235 ( .A1(a[7]), .A2(b[7]), .ZN(y[119]) );
  OR2_X1 U235bar ( .A1(abar[7]), .A2(bbar[7]), .ZN(ybar[119]) );
  AND2_X1 U236 ( .A1(a[7]), .A2(b[6]), .ZN(y[118]) );
  OR2_X1 U236bar ( .A1(abar[7]), .A2(bbar[6]), .ZN(ybar[118]) );
  AND2_X1 U237 ( .A1(a[7]), .A2(b[5]), .ZN(y[117]) );
  OR2_X1 U237bar ( .A1(abar[7]), .A2(bbar[5]), .ZN(ybar[117]) );
  AND2_X1 U238 ( .A1(a[7]), .A2(b[4]), .ZN(y[116]) );
  OR2_X1 U238bar ( .A1(abar[7]), .A2(bbar[4]), .ZN(ybar[116]) );
  AND2_X1 U239 ( .A1(a[7]), .A2(b[3]), .ZN(y[115]) );
  OR2_X1 U239bar ( .A1(abar[7]), .A2(bbar[3]), .ZN(ybar[115]) );
  AND2_X1 U240 ( .A1(a[7]), .A2(b[2]), .ZN(y[114]) );
  OR2_X1 U240bar ( .A1(abar[7]), .A2(bbar[2]), .ZN(ybar[114]) );
  AND2_X1 U241 ( .A1(a[7]), .A2(b[1]), .ZN(y[113]) );
  OR2_X1 U241bar ( .A1(abar[7]), .A2(bbar[1]), .ZN(ybar[113]) );
  AND2_X1 U242 ( .A1(a[7]), .A2(b[0]), .ZN(y[112]) );
  OR2_X1 U242bar ( .A1(abar[7]), .A2(bbar[0]), .ZN(ybar[112]) );
  AND2_X1 U243 ( .A1(b[15]), .A2(a[6]), .ZN(y[111]) );
  OR2_X1 U243bar ( .A1(bbar[15]), .A2(abar[6]), .ZN(ybar[111]) );
  AND2_X1 U244 ( .A1(b[14]), .A2(a[6]), .ZN(y[110]) );
  OR2_X1 U244bar ( .A1(bbar[14]), .A2(abar[6]), .ZN(ybar[110]) );
  AND2_X1 U245 ( .A1(b[10]), .A2(a[0]), .ZN(y[10]) );
  OR2_X1 U245bar ( .A1(bbar[10]), .A2(abar[0]), .ZN(ybar[10]) );
  AND2_X1 U246 ( .A1(b[13]), .A2(a[6]), .ZN(y[109]) );
  OR2_X1 U246bar ( .A1(bbar[13]), .A2(abar[6]), .ZN(ybar[109]) );
  AND2_X1 U247 ( .A1(b[12]), .A2(a[6]), .ZN(y[108]) );
  OR2_X1 U247bar ( .A1(bbar[12]), .A2(abar[6]), .ZN(ybar[108]) );
  AND2_X1 U248 ( .A1(b[11]), .A2(a[6]), .ZN(y[107]) );
  OR2_X1 U248bar ( .A1(bbar[11]), .A2(abar[6]), .ZN(ybar[107]) );
  AND2_X1 U249 ( .A1(b[10]), .A2(a[6]), .ZN(y[106]) );
  OR2_X1 U249bar ( .A1(bbar[10]), .A2(abar[6]), .ZN(ybar[106]) );
  AND2_X1 U250 ( .A1(a[6]), .A2(b[9]), .ZN(y[105]) );
  OR2_X1 U250bar ( .A1(abar[6]), .A2(bbar[9]), .ZN(ybar[105]) );
  AND2_X1 U251 ( .A1(b[8]), .A2(a[6]), .ZN(y[104]) );
  OR2_X1 U251bar ( .A1(bbar[8]), .A2(abar[6]), .ZN(ybar[104]) );
  AND2_X1 U252 ( .A1(b[7]), .A2(a[6]), .ZN(y[103]) );
  OR2_X1 U252bar ( .A1(bbar[7]), .A2(abar[6]), .ZN(ybar[103]) );
  AND2_X1 U253 ( .A1(b[6]), .A2(a[6]), .ZN(y[102]) );
  OR2_X1 U253bar ( .A1(bbar[6]), .A2(abar[6]), .ZN(ybar[102]) );
  AND2_X1 U254 ( .A1(b[5]), .A2(a[6]), .ZN(y[101]) );
  OR2_X1 U254bar ( .A1(bbar[5]), .A2(abar[6]), .ZN(ybar[101]) );
  AND2_X1 U255 ( .A1(b[4]), .A2(a[6]), .ZN(y[100]) );
  OR2_X1 U255bar ( .A1(bbar[4]), .A2(abar[6]), .ZN(ybar[100]) );
  AND2_X1 U256 ( .A1(b[0]), .A2(a[0]), .ZN(y[0]) );
  OR2_X1 U256bar ( .A1(bbar[0]), .A2(abar[0]), .ZN(ybar[0]) );
endmodule

module decode_2 ( in, inbar, out, outbar );

  input wire [7:0] in;
  input wire [7:0] inbar;
//input_done

  output wire [255:0] out;
  output wire [255:0] outbar;
//output_done

  wire [15:0] level1;
  wire [31:0] level2;
  wire [15:0] level1bar;
  wire [31:0] level2bar;
//wire_done

  CD2_8 cd_l1_1 ( .a(in[1]), .abar(inbar[1]), .b(in[0]), .bbar(inbar[0]), .y(level1[3:0]), .ybar(level1bar[3:0]) );
  CD2_7 cd_l1_2 ( .a(in[3]), .abar(inbar[3]), .b(in[2]), .bbar(inbar[2]), .y(level1[7:4]), .ybar(level1bar[7:4]) );
  CD2_6 cd_l1_3 ( .a(in[5]), .abar(inbar[5]), .b(in[4]), .bbar(inbar[4]), .y(level1[11:8]), .ybar(level1bar[11:8]) );
  CD2_5 cd_l1_4 ( .a(in[7]), .abar(inbar[7]), .b(in[6]), .bbar(inbar[6]), .y(level1[15:12]), .ybar(level1bar[15:12]) );

  CD4_4 cd_l2_1 ( .a(level1[7:4]), .abar(level1bar[7:4]), .b(level1[3:0]), .bbar(level1bar[3:0]), 
        .y(level2[15:0]), .ybar(level2bar[15:0]) );
  CD4_3 cd_l2_2 ( .a(level1[15:12]), .abar(level1bar[15:12]), .b(level1[11:8]), .bbar(level1bar[11:8]), 
        .y(level2[31:16]), .ybar(level2bar[31:16]) );
  CD16_2 cd_l3 ( .a(level2[31:16]), .abar(level2bar[31:16]), .b(level2[15:0]), .bbar(level2bar[15:0]), 
        .y(out), .ybar(outbar) );
endmodule

module encode_2 ( in, inbar, out, outbar );

  input wire [255:0] in;
  input wire [255:0] inbar;
//input_done

  output wire [7:0] out;
  output wire [7:0] outbar;
//output_done

  wire in_81;
  wire in_80;
  wire in_79;
  wire in_78;
  wire in_77;
  wire in_76;
  wire in_75;
  wire in_74;
  wire in_73;
  wire in_72;
  wire in_71;
  wire in_70;
  wire in_69;
  wire in_68;
  wire in_67;
  wire in_66;
  wire in_65;
  wire in_64;
  wire in_63;
  wire in_62;
  wire in_61;
  wire in_60;
  wire in_59;
  wire in_58;
  wire in_57;
  wire in_56;
  wire in_55;
  wire in_54;
  wire in_53;
  wire in_52;
  wire in_51;
  wire in_50;
  wire in_49;
  wire in_48;
  wire in_47;
  wire in_46;
  wire in_45;
  wire in_44;
  wire in_43;
  wire in_42;
  wire in_41;
  wire in_40;
  wire in_39;
  wire in_38;
  wire in_37;
  wire in_36;
  wire in_35;
  wire in_34;
  wire in_33;
  wire in_32;
  wire in_31;
  wire in_30;
  wire in_29;
  wire in_28;
  wire in_27;
  wire in_26;
  wire in_25;
  wire in_24;
  wire in_23;
  wire in_22;
  wire in_21;
  wire in_20;
  wire in_19;
  wire in_18;
  wire in_17;
  wire in_16;
  wire in_15;
  wire in_14;
  wire in_13;
  wire in_12;
  wire in_11;
  wire in_10;
  wire in_9;
  wire in_8;
  wire in_7;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_3;
  wire in_2;
  wire in_1;
  wire in_0;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire in_81bar;
  wire in_80bar;
  wire in_79bar;
  wire in_78bar;
  wire in_77bar;
  wire in_76bar;
  wire in_75bar;
  wire in_74bar;
  wire in_73bar;
  wire in_72bar;
  wire in_71bar;
  wire in_70bar;
  wire in_69bar;
  wire in_68bar;
  wire in_67bar;
  wire in_66bar;
  wire in_65bar;
  wire in_64bar;
  wire in_63bar;
  wire in_62bar;
  wire in_61bar;
  wire in_60bar;
  wire in_59bar;
  wire in_58bar;
  wire in_57bar;
  wire in_56bar;
  wire in_55bar;
  wire in_54bar;
  wire in_53bar;
  wire in_52bar;
  wire in_51bar;
  wire in_50bar;
  wire in_49bar;
  wire in_48bar;
  wire in_47bar;
  wire in_46bar;
  wire in_45bar;
  wire in_44bar;
  wire in_43bar;
  wire in_42bar;
  wire in_41bar;
  wire in_40bar;
  wire in_39bar;
  wire in_38bar;
  wire in_37bar;
  wire in_36bar;
  wire in_35bar;
  wire in_34bar;
  wire in_33bar;
  wire in_32bar;
  wire in_31bar;
  wire in_30bar;
  wire in_29bar;
  wire in_28bar;
  wire in_27bar;
  wire in_26bar;
  wire in_25bar;
  wire in_24bar;
  wire in_23bar;
  wire in_22bar;
  wire in_21bar;
  wire in_20bar;
  wire in_19bar;
  wire in_18bar;
  wire in_17bar;
  wire in_16bar;
  wire in_15bar;
  wire in_14bar;
  wire in_13bar;
  wire in_12bar;
  wire in_11bar;
  wire in_10bar;
  wire in_9bar;
  wire in_8bar;
  wire in_7bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_3bar;
  wire in_2bar;
  wire in_1bar;
  wire in_0bar;
  wire n487bar;
  wire n488bar;
  wire n489bar;
  wire n490bar;
  wire n491bar;
  wire n492bar;
  wire n493bar;
  wire n494bar;
  wire n495bar;
  wire n496bar;
  wire n497bar;
  wire n498bar;
  wire n499bar;
  wire n500bar;
  wire n501bar;
  wire n502bar;
  wire n503bar;
  wire n504bar;
  wire n505bar;
  wire n506bar;
  wire n507bar;
  wire n508bar;
  wire n509bar;
  wire n510bar;
  wire n511bar;
  wire n512bar;
  wire n513bar;
  wire n514bar;
  wire n515bar;
  wire n516bar;
  wire n517bar;
  wire n518bar;
  wire n519bar;
  wire n520bar;
  wire n521bar;
  wire n522bar;
  wire n523bar;
  wire n524bar;
  wire n525bar;
  wire n526bar;
  wire n527bar;
  wire n528bar;
  wire n529bar;
  wire n530bar;
  wire n531bar;
  wire n532bar;
  wire n533bar;
  wire n534bar;
  wire n535bar;
  wire n536bar;
  wire n537bar;
  wire n538bar;
  wire n539bar;
  wire n540bar;
  wire n541bar;
  wire n542bar;
  wire n543bar;
  wire n544bar;
  wire n545bar;
  wire n546bar;
  wire n547bar;
  wire n548bar;
  wire n549bar;
  wire n550bar;
  wire n551bar;
  wire n552bar;
  wire n553bar;
  wire n554bar;
  wire n555bar;
  wire n556bar;
  wire n557bar;
  wire n558bar;
  wire n559bar;
  wire n560bar;
  wire n561bar;
  wire n562bar;
  wire n563bar;
  wire n564bar;
  wire n565bar;
  wire n566bar;
  wire n567bar;
  wire n568bar;
  wire n569bar;
  wire n570bar;
  wire n571bar;
  wire n572bar;
  wire n573bar;
  wire n574bar;
  wire n575bar;
  wire n576bar;
  wire n577bar;
  wire n578bar;
  wire n579bar;
  wire n580bar;
  wire n581bar;
  wire n582bar;
  wire n583bar;
  wire n584bar;
  wire n585bar;
  wire n586bar;
  wire n587bar;
  wire n588bar;
  wire n589bar;
  wire n590bar;
  wire n591bar;
  wire n592bar;
  wire n593bar;
  wire n594bar;
  wire n595bar;
  wire n596bar;
  wire n597bar;
  wire n598bar;
  wire n599bar;
  wire n600bar;
  wire n601bar;
  wire n602bar;
  wire n603bar;
  wire n604bar;
  wire n605bar;
  wire n606bar;
  wire n607bar;
  wire n608bar;
  wire n609bar;
  wire n610bar;
  wire n611bar;
  wire n612bar;
  wire n613bar;
  wire n614bar;
  wire n615bar;
  wire n616bar;
  wire n617bar;
  wire n618bar;
  wire n619bar;
  wire n620bar;
  wire n621bar;
  wire n622bar;
  wire n623bar;
  wire n624bar;
  wire n625bar;
  wire n626bar;
  wire n627bar;
  wire n628bar;
  wire n629bar;
  wire n630bar;
  wire n631bar;
  wire n632bar;
  wire n633bar;
  wire n634bar;
  wire n635bar;
  wire n636bar;
  wire n637bar;
  wire n638bar;
  wire n639bar;
  wire n640bar;
  wire n641bar;
  wire n642bar;
  wire n643bar;
  wire n644bar;
  wire n645bar;
  wire n646bar;
  wire n647bar;
  wire n648bar;
  wire n649bar;
  wire n650bar;
  wire n651bar;
  wire n652bar;
  wire n653bar;
  wire n654bar;
  wire n655bar;
  wire n656bar;
  wire n657bar;
  wire n658bar;
  wire n659bar;
  wire n660bar;
  wire n661bar;
  wire n662bar;
  wire n663bar;
  wire n664bar;
  wire n665bar;
  wire n666bar;
  wire n667bar;
  wire n668bar;
  wire n669bar;
  wire n670bar;
  wire n671bar;
  wire n672bar;
  wire n673bar;
  wire n674bar;
  wire n675bar;
  wire n676bar;
  wire n677bar;
  wire n678bar;
  wire n679bar;
  wire n680bar;
  wire n681bar;
  wire n682bar;
  wire n683bar;
  wire n684bar;
  wire n685bar;
  wire n686bar;
  wire n687bar;
  wire n688bar;
  wire n689bar;
  wire n690bar;
  wire n691bar;
  wire n692bar;
  wire n693bar;
  wire n694bar;
  wire n695bar;
  wire n696bar;
  wire n697bar;
  wire n698bar;
  wire n699bar;
  wire n700bar;
  wire n701bar;
  wire n702bar;
  wire n703bar;
  wire n704bar;
  wire n705bar;
  wire n706bar;
  wire n707bar;
  wire n708bar;
  wire n709bar;
  wire n710bar;
  wire n711bar;
  wire n712bar;
  wire n713bar;
  wire n714bar;
  wire n715bar;
  wire n716bar;
  wire n717bar;
  wire n718bar;
  wire n719bar;
  wire n720bar;
  wire n721bar;
  wire n722bar;
  wire n723bar;
  wire n724bar;
  wire n725bar;
  wire n726bar;
  wire n727bar;
  wire n728bar;
  wire n729bar;
  wire n730bar;
  wire n731bar;
  wire n732bar;
  wire n733bar;
  wire n734bar;
  wire n735bar;
  wire n736bar;
  wire n737bar;
  wire n738bar;
  wire n739bar;
  wire n740bar;
  wire n741bar;
  wire n742bar;
  wire n743bar;
  wire n744bar;
  wire n745bar;
  wire n746bar;
  wire n747bar;
  wire n748bar;
  wire n749bar;
  wire n750bar;
  wire n751bar;
  wire n752bar;
  wire n753bar;
  wire n754bar;
  wire n755bar;
  wire n756bar;
  wire n757bar;
  wire n758bar;
  wire n759bar;
  wire n760bar;
  wire n761bar;
  wire n762bar;
  wire n763bar;
  wire n764bar;
  wire n765bar;
  wire n766bar;
  wire n767bar;
  wire n768bar;
  wire n769bar;
  wire n770bar;
  wire n771bar;
  wire n772bar;
  wire n773bar;
  wire n774bar;
  wire n775bar;
  wire n776bar;
  wire n777bar;
  wire n778bar;
  wire n779bar;
  wire n780bar;
  wire n781bar;
  wire n782bar;
  wire n783bar;
  wire n784bar;
  wire n785bar;
  wire n786bar;
  wire n787bar;
  wire n788bar;
  wire n789bar;
  wire n790bar;
  wire n791bar;
  wire n792bar;
  wire n793bar;
  wire n794bar;
  wire n795bar;
  wire n796bar;
  wire n797bar;
  wire n798bar;
  wire n799bar;
  wire n800bar;
  wire n801bar;
  wire n802bar;
  wire n803bar;
  wire n804bar;
  wire n805bar;
  wire n806bar;
  wire n807bar;
  wire n808bar;
  wire n809bar;
  wire n810bar;
  wire n811bar;
  wire n812bar;
  wire n813bar;
  wire n814bar;
  wire n815bar;
  wire n816bar;
  wire n817bar;
  wire n818bar;
  wire n819bar;
  wire n820bar;
  wire n821bar;
  wire n822bar;
  wire n823bar;
  wire n824bar;
  wire n825bar;
  wire n826bar;
  wire n827bar;
  wire n828bar;
  wire n829bar;
  wire n830bar;
  wire n831bar;
  wire n832bar;
  wire n833bar;
  wire n834bar;
  wire n835bar;
  wire n836bar;
  wire n837bar;
  wire n838bar;
  wire n839bar;
  wire n840bar;
  wire n841bar;
  wire n842bar;
  wire n843bar;
  wire n844bar;
  wire n845bar;
  wire n846bar;
  wire n847bar;
  wire n848bar;
  wire n849bar;
  wire n850bar;
  wire n851bar;
  wire n852bar;
  wire n853bar;
  wire n854bar;
  wire n855bar;
  wire n856bar;
  wire n857bar;
  wire n858bar;
  wire n859bar;
  wire n860bar;
  wire n861bar;
  wire n862bar;
  wire n863bar;
  wire n864bar;
  wire n865bar;
  wire n866bar;
  wire n867bar;
  wire n868bar;
  wire n869bar;
  wire n870bar;
  wire n871bar;
  wire n872bar;
  wire n873bar;
  wire n874bar;
  wire n875bar;
  wire n876bar;
  wire n877bar;
  wire n878bar;
  wire n879bar;
  wire n880bar;
  wire n881bar;
  wire n882bar;
  wire n883bar;
  wire n884bar;
  wire n885bar;
  wire n886bar;
  wire n887bar;
  wire n888bar;
  wire n889bar;
  wire n890bar;
  wire n891bar;
  wire n892bar;
  wire n893bar;
  wire n894bar;
  wire n895bar;
  wire n896bar;
  wire n897bar;
  wire n898bar;
  wire n899bar;
  wire n900bar;
  wire n901bar;
  wire n902bar;
  wire n903bar;
  wire n904bar;
  wire n905bar;
  wire n906bar;
  wire n907bar;
  wire n908bar;
  wire n909bar;
  wire n910bar;
  wire n911bar;
  wire n912bar;
  wire n913bar;
  wire n914bar;
  wire n915bar;
  wire n916bar;
  wire n917bar;
  wire n918bar;
  wire n919bar;
  wire n920bar;
  wire n921bar;
  wire n922bar;
  wire n923bar;
  wire n924bar;
  wire n925bar;
  wire n926bar;
  wire n927bar;
  wire n928bar;
  wire n929bar;
  wire n930bar;
  wire n931bar;
  wire n932bar;
  wire n933bar;
  wire n934bar;
  wire n935bar;
  wire n936bar;
  wire n937bar;
  wire n938bar;
  wire n939bar;
  wire n940bar;
  wire n941bar;
  wire n942bar;
  wire n943bar;
  wire n944bar;
  wire n945bar;
  wire n946bar;
  wire n947bar;
  wire n948bar;
  wire n949bar;
  wire n950bar;
  wire n951bar;
  wire n952bar;
  wire n953bar;
  wire n954bar;
  wire n955bar;
  wire n956bar;
  wire n957bar;
  wire n958bar;
  wire n959bar;
  wire n960bar;
  wire n961bar;
  wire n962bar;
  wire n963bar;
  wire n964bar;
  wire n965bar;
  wire n966bar;
  wire n967bar;
  wire n968bar;
  wire n969bar;
  wire n970bar;
  wire n971bar;
  wire n972bar;
//wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];
  assign in_81bar = inbar[81];
  assign in_80bar = inbar[80];
  assign in_79bar = inbar[79];
  assign in_78bar = inbar[78];
  assign in_77bar = inbar[77];
  assign in_76bar = inbar[76];
  assign in_75bar = inbar[75];
  assign in_74bar = inbar[74];
  assign in_73bar = inbar[73];
  assign in_72bar = inbar[72];
  assign in_71bar = inbar[71];
  assign in_70bar = inbar[70];
  assign in_69bar = inbar[69];
  assign in_68bar = inbar[68];
  assign in_67bar = inbar[67];
  assign in_66bar = inbar[66];
  assign in_65bar = inbar[65];
  assign in_64bar = inbar[64];
  assign in_63bar = inbar[63];
  assign in_62bar = inbar[62];
  assign in_61bar = inbar[61];
  assign in_60bar = inbar[60];
  assign in_59bar = inbar[59];
  assign in_58bar = inbar[58];
  assign in_57bar = inbar[57];
  assign in_56bar = inbar[56];
  assign in_55bar = inbar[55];
  assign in_54bar = inbar[54];
  assign in_53bar = inbar[53];
  assign in_52bar = inbar[52];
  assign in_51bar = inbar[51];
  assign in_50bar = inbar[50];
  assign in_49bar = inbar[49];
  assign in_48bar = inbar[48];
  assign in_47bar = inbar[47];
  assign in_46bar = inbar[46];
  assign in_45bar = inbar[45];
  assign in_44bar = inbar[44];
  assign in_43bar = inbar[43];
  assign in_42bar = inbar[42];
  assign in_41bar = inbar[41];
  assign in_40bar = inbar[40];
  assign in_39bar = inbar[39];
  assign in_38bar = inbar[38];
  assign in_37bar = inbar[37];
  assign in_36bar = inbar[36];
  assign in_35bar = inbar[35];
  assign in_34bar = inbar[34];
  assign in_33bar = inbar[33];
  assign in_32bar = inbar[32];
  assign in_31bar = inbar[31];
  assign in_30bar = inbar[30];
  assign in_29bar = inbar[29];
  assign in_28bar = inbar[28];
  assign in_27bar = inbar[27];
  assign in_26bar = inbar[26];
  assign in_25bar = inbar[25];
  assign in_24bar = inbar[24];
  assign in_23bar = inbar[23];
  assign in_22bar = inbar[22];
  assign in_21bar = inbar[21];
  assign in_20bar = inbar[20];
  assign in_19bar = inbar[19];
  assign in_18bar = inbar[18];
  assign in_17bar = inbar[17];
  assign in_16bar = inbar[16];
  assign in_15bar = inbar[15];
  assign in_14bar = inbar[14];
  assign in_13bar = inbar[13];
  assign in_12bar = inbar[12];
  assign in_11bar = inbar[11];
  assign in_10bar = inbar[10];
  assign in_9bar = inbar[9];
  assign in_8bar = inbar[8];
  assign in_7bar = inbar[7];
  assign in_6bar = inbar[6];
  assign in_5bar = inbar[5];
  assign in_4bar = inbar[4];
  assign in_3bar = inbar[3];
  assign in_2bar = inbar[2];
  assign in_1bar = inbar[1];
  assign in_0bar = inbar[0];
//assign_done

  OR2_X1 U1 ( .A1(n972), .A2(n971), .ZN(out[7]) );
  AND2_X1 U1bar ( .A1(n972bar), .A2(n971bar), .ZN(outbar[7]) );
  OR2_X1 U2 ( .A1(n970), .A2(n969), .ZN(n971) );
  AND2_X1 U2bar ( .A1(n970bar), .A2(n969bar), .ZN(n971bar) );
  OR2_X1 U3 ( .A1(n968), .A2(n967), .ZN(n969) );
  AND2_X1 U3bar ( .A1(n968bar), .A2(n967bar), .ZN(n969bar) );
  OR2_X1 U4 ( .A1(n966), .A2(n965), .ZN(n967) );
  AND2_X1 U4bar ( .A1(n966bar), .A2(n965bar), .ZN(n967bar) );
  OR2_X1 U5 ( .A1(n964), .A2(n963), .ZN(n968) );
  AND2_X1 U5bar ( .A1(n964bar), .A2(n963bar), .ZN(n968bar) );
  OR2_X1 U6 ( .A1(in[116]), .A2(n962), .ZN(n963) );
  AND2_X1 U6bar ( .A1(inbar[116]), .A2(n962bar), .ZN(n963bar) );
  OR2_X1 U7 ( .A1(n961), .A2(n960), .ZN(n970) );
  AND2_X1 U7bar ( .A1(n961bar), .A2(n960bar), .ZN(n970bar) );
  OR2_X1 U8 ( .A1(in[150]), .A2(in[127]), .ZN(n960) );
  AND2_X1 U8bar ( .A1(inbar[150]), .A2(inbar[127]), .ZN(n960bar) );
  OR2_X1 U9 ( .A1(in[160]), .A2(n959), .ZN(n961) );
  AND2_X1 U9bar ( .A1(inbar[160]), .A2(n959bar), .ZN(n961bar) );
  OR2_X1 U10 ( .A1(in[252]), .A2(in[168]), .ZN(n959) );
  AND2_X1 U10bar ( .A1(inbar[252]), .A2(inbar[168]), .ZN(n959bar) );
  OR2_X1 U11 ( .A1(n958), .A2(n957), .ZN(n972) );
  AND2_X1 U11bar ( .A1(n958bar), .A2(n957bar), .ZN(n972bar) );
  OR2_X1 U12 ( .A1(n956), .A2(n955), .ZN(n957) );
  AND2_X1 U12bar ( .A1(n956bar), .A2(n955bar), .ZN(n957bar) );
  OR2_X1 U13 ( .A1(in_17), .A2(in[96]), .ZN(n955) );
  AND2_X1 U13bar ( .A1(in_17bar), .A2(inbar[96]), .ZN(n955bar) );
  OR2_X1 U14 ( .A1(in_23), .A2(n954), .ZN(n956) );
  AND2_X1 U14bar ( .A1(in_23bar), .A2(n954bar), .ZN(n956bar) );
  OR2_X1 U15 ( .A1(in_31), .A2(in_26), .ZN(n954) );
  AND2_X1 U15bar ( .A1(in_31bar), .A2(in_26bar), .ZN(n954bar) );
  OR2_X1 U16 ( .A1(n953), .A2(n952), .ZN(n958) );
  AND2_X1 U16bar ( .A1(n953bar), .A2(n952bar), .ZN(n958bar) );
  OR2_X1 U17 ( .A1(in_58), .A2(in_4), .ZN(n952) );
  AND2_X1 U17bar ( .A1(in_58bar), .A2(in_4bar), .ZN(n952bar) );
  OR2_X1 U18 ( .A1(in_59), .A2(n951), .ZN(n953) );
  AND2_X1 U18bar ( .A1(in_59bar), .A2(n951bar), .ZN(n953bar) );
  OR2_X1 U19 ( .A1(in_71), .A2(in_62), .ZN(n951) );
  AND2_X1 U19bar ( .A1(in_71bar), .A2(in_62bar), .ZN(n951bar) );
  OR2_X1 U20 ( .A1(n950), .A2(n949), .ZN(out[6]) );
  AND2_X1 U20bar ( .A1(n950bar), .A2(n949bar), .ZN(outbar[6]) );
  OR2_X1 U21 ( .A1(n948), .A2(n947), .ZN(n949) );
  AND2_X1 U21bar ( .A1(n948bar), .A2(n947bar), .ZN(n949bar) );
  OR2_X1 U22 ( .A1(n946), .A2(n945), .ZN(n947) );
  AND2_X1 U22bar ( .A1(n946bar), .A2(n945bar), .ZN(n947bar) );
  OR2_X1 U23 ( .A1(n944), .A2(n943), .ZN(n945) );
  AND2_X1 U23bar ( .A1(n944bar), .A2(n943bar), .ZN(n945bar) );
  OR2_X1 U24 ( .A1(n942), .A2(n941), .ZN(n946) );
  AND2_X1 U24bar ( .A1(n942bar), .A2(n941bar), .ZN(n946bar) );
  OR2_X1 U25 ( .A1(in[101]), .A2(n940), .ZN(n941) );
  AND2_X1 U25bar ( .A1(inbar[101]), .A2(n940bar), .ZN(n941bar) );
  OR2_X1 U26 ( .A1(n939), .A2(n938), .ZN(n948) );
  AND2_X1 U26bar ( .A1(n939bar), .A2(n938bar), .ZN(n948bar) );
  OR2_X1 U27 ( .A1(in[114]), .A2(in[104]), .ZN(n938) );
  AND2_X1 U27bar ( .A1(inbar[114]), .A2(inbar[104]), .ZN(n938bar) );
  OR2_X1 U28 ( .A1(in[128]), .A2(n937), .ZN(n939) );
  AND2_X1 U28bar ( .A1(inbar[128]), .A2(n937bar), .ZN(n939bar) );
  OR2_X1 U29 ( .A1(in[136]), .A2(in[134]), .ZN(n937) );
  AND2_X1 U29bar ( .A1(inbar[136]), .A2(inbar[134]), .ZN(n937bar) );
  OR2_X1 U30 ( .A1(n936), .A2(n935), .ZN(n950) );
  AND2_X1 U30bar ( .A1(n936bar), .A2(n935bar), .ZN(n950bar) );
  OR2_X1 U31 ( .A1(n934), .A2(n933), .ZN(n935) );
  AND2_X1 U31bar ( .A1(n934bar), .A2(n933bar), .ZN(n935bar) );
  OR2_X1 U32 ( .A1(in[177]), .A2(in[164]), .ZN(n933) );
  AND2_X1 U32bar ( .A1(inbar[177]), .A2(inbar[164]), .ZN(n933bar) );
  OR2_X1 U33 ( .A1(in[212]), .A2(n932), .ZN(n934) );
  AND2_X1 U33bar ( .A1(inbar[212]), .A2(n932bar), .ZN(n934bar) );
  OR2_X1 U34 ( .A1(in[248]), .A2(in[221]), .ZN(n932) );
  AND2_X1 U34bar ( .A1(inbar[248]), .A2(inbar[221]), .ZN(n932bar) );
  OR2_X1 U35 ( .A1(n931), .A2(n930), .ZN(n936) );
  AND2_X1 U35bar ( .A1(n931bar), .A2(n930bar), .ZN(n936bar) );
  OR2_X1 U36 ( .A1(in_18), .A2(in[93]), .ZN(n930) );
  AND2_X1 U36bar ( .A1(in_18bar), .A2(inbar[93]), .ZN(n930bar) );
  OR2_X1 U37 ( .A1(in_31), .A2(n929), .ZN(n931) );
  AND2_X1 U37bar ( .A1(in_31bar), .A2(n929bar), .ZN(n931bar) );
  OR2_X1 U38 ( .A1(in_7), .A2(in_39), .ZN(n929) );
  AND2_X1 U38bar ( .A1(in_7bar), .A2(in_39bar), .ZN(n929bar) );
  OR2_X1 U39 ( .A1(n928), .A2(n927), .ZN(out[5]) );
  AND2_X1 U39bar ( .A1(n928bar), .A2(n927bar), .ZN(outbar[5]) );
  OR2_X1 U40 ( .A1(n926), .A2(n925), .ZN(n927) );
  AND2_X1 U40bar ( .A1(n926bar), .A2(n925bar), .ZN(n927bar) );
  OR2_X1 U41 ( .A1(n924), .A2(n923), .ZN(n925) );
  AND2_X1 U41bar ( .A1(n924bar), .A2(n923bar), .ZN(n925bar) );
  OR2_X1 U42 ( .A1(n922), .A2(n921), .ZN(n923) );
  AND2_X1 U42bar ( .A1(n922bar), .A2(n921bar), .ZN(n923bar) );
  OR2_X1 U43 ( .A1(n940), .A2(n920), .ZN(n924) );
  AND2_X1 U43bar ( .A1(n940bar), .A2(n920bar), .ZN(n924bar) );
  OR2_X1 U44 ( .A1(in[111]), .A2(n919), .ZN(n920) );
  AND2_X1 U44bar ( .A1(inbar[111]), .A2(n919bar), .ZN(n920bar) );
  OR2_X1 U45 ( .A1(n918), .A2(n917), .ZN(n940) );
  AND2_X1 U45bar ( .A1(n918bar), .A2(n917bar), .ZN(n940bar) );
  OR2_X1 U46 ( .A1(n916), .A2(n915), .ZN(n917) );
  AND2_X1 U46bar ( .A1(n916bar), .A2(n915bar), .ZN(n917bar) );
  OR2_X1 U47 ( .A1(n914), .A2(n913), .ZN(n915) );
  AND2_X1 U47bar ( .A1(n914bar), .A2(n913bar), .ZN(n915bar) );
  OR2_X1 U48 ( .A1(in[140]), .A2(in[131]), .ZN(n913) );
  AND2_X1 U48bar ( .A1(inbar[140]), .A2(inbar[131]), .ZN(n913bar) );
  OR2_X1 U49 ( .A1(in[160]), .A2(in[144]), .ZN(n914) );
  AND2_X1 U49bar ( .A1(inbar[160]), .A2(inbar[144]), .ZN(n914bar) );
  OR2_X1 U50 ( .A1(n912), .A2(n911), .ZN(n916) );
  AND2_X1 U50bar ( .A1(n912bar), .A2(n911bar), .ZN(n916bar) );
  OR2_X1 U51 ( .A1(in[179]), .A2(in[174]), .ZN(n911) );
  AND2_X1 U51bar ( .A1(inbar[179]), .A2(inbar[174]), .ZN(n911bar) );
  OR2_X1 U52 ( .A1(in[188]), .A2(in[184]), .ZN(n912) );
  AND2_X1 U52bar ( .A1(inbar[188]), .A2(inbar[184]), .ZN(n912bar) );
  OR2_X1 U53 ( .A1(n910), .A2(n909), .ZN(n918) );
  AND2_X1 U53bar ( .A1(n910bar), .A2(n909bar), .ZN(n918bar) );
  OR2_X1 U54 ( .A1(n908), .A2(n907), .ZN(n909) );
  AND2_X1 U54bar ( .A1(n908bar), .A2(n907bar), .ZN(n909bar) );
  OR2_X1 U55 ( .A1(in[216]), .A2(in[200]), .ZN(n907) );
  AND2_X1 U55bar ( .A1(inbar[216]), .A2(inbar[200]), .ZN(n907bar) );
  OR2_X1 U56 ( .A1(in[228]), .A2(in[224]), .ZN(n908) );
  AND2_X1 U56bar ( .A1(inbar[228]), .A2(inbar[224]), .ZN(n908bar) );
  OR2_X1 U57 ( .A1(n906), .A2(n905), .ZN(n910) );
  AND2_X1 U57bar ( .A1(n906bar), .A2(n905bar), .ZN(n910bar) );
  OR2_X1 U58 ( .A1(in[247]), .A2(in[235]), .ZN(n905) );
  AND2_X1 U58bar ( .A1(inbar[247]), .A2(inbar[235]), .ZN(n905bar) );
  OR2_X1 U59 ( .A1(in_42), .A2(in[83]), .ZN(n906) );
  AND2_X1 U59bar ( .A1(in_42bar), .A2(inbar[83]), .ZN(n906bar) );
  OR2_X1 U60 ( .A1(n904), .A2(n903), .ZN(n926) );
  AND2_X1 U60bar ( .A1(n904bar), .A2(n903bar), .ZN(n926bar) );
  OR2_X1 U61 ( .A1(in[166]), .A2(in[123]), .ZN(n903) );
  AND2_X1 U61bar ( .A1(inbar[166]), .A2(inbar[123]), .ZN(n903bar) );
  OR2_X1 U62 ( .A1(in[170]), .A2(n902), .ZN(n904) );
  AND2_X1 U62bar ( .A1(inbar[170]), .A2(n902bar), .ZN(n904bar) );
  OR2_X1 U63 ( .A1(in[194]), .A2(in[183]), .ZN(n902) );
  AND2_X1 U63bar ( .A1(inbar[194]), .A2(inbar[183]), .ZN(n902bar) );
  OR2_X1 U64 ( .A1(n901), .A2(n900), .ZN(n928) );
  AND2_X1 U64bar ( .A1(n901bar), .A2(n900bar), .ZN(n928bar) );
  OR2_X1 U65 ( .A1(n899), .A2(n898), .ZN(n900) );
  AND2_X1 U65bar ( .A1(n899bar), .A2(n898bar), .ZN(n900bar) );
  OR2_X1 U66 ( .A1(in[241]), .A2(in[238]), .ZN(n898) );
  AND2_X1 U66bar ( .A1(inbar[241]), .A2(inbar[238]), .ZN(n898bar) );
  OR2_X1 U67 ( .A1(in[250]), .A2(n897), .ZN(n899) );
  AND2_X1 U67bar ( .A1(inbar[250]), .A2(n897bar), .ZN(n899bar) );
  OR2_X1 U68 ( .A1(in_24), .A2(in[84]), .ZN(n897) );
  AND2_X1 U68bar ( .A1(in_24bar), .A2(inbar[84]), .ZN(n897bar) );
  OR2_X1 U69 ( .A1(n896), .A2(n895), .ZN(n901) );
  AND2_X1 U69bar ( .A1(n896bar), .A2(n895bar), .ZN(n901bar) );
  OR2_X1 U70 ( .A1(in_41), .A2(in_29), .ZN(n895) );
  AND2_X1 U70bar ( .A1(in_41bar), .A2(in_29bar), .ZN(n895bar) );
  OR2_X1 U71 ( .A1(in_66), .A2(n894), .ZN(n896) );
  AND2_X1 U71bar ( .A1(in_66bar), .A2(n894bar), .ZN(n896bar) );
  OR2_X1 U72 ( .A1(in_76), .A2(in_71), .ZN(n894) );
  AND2_X1 U72bar ( .A1(in_76bar), .A2(in_71bar), .ZN(n894bar) );
  OR2_X1 U73 ( .A1(n893), .A2(n892), .ZN(out[4]) );
  AND2_X1 U73bar ( .A1(n893bar), .A2(n892bar), .ZN(outbar[4]) );
  OR2_X1 U74 ( .A1(n891), .A2(n890), .ZN(n892) );
  AND2_X1 U74bar ( .A1(n891bar), .A2(n890bar), .ZN(n892bar) );
  OR2_X1 U75 ( .A1(n889), .A2(n888), .ZN(n890) );
  AND2_X1 U75bar ( .A1(n889bar), .A2(n888bar), .ZN(n890bar) );
  OR2_X1 U76 ( .A1(n922), .A2(n887), .ZN(n888) );
  AND2_X1 U76bar ( .A1(n922bar), .A2(n887bar), .ZN(n888bar) );
  OR2_X1 U77 ( .A1(n886), .A2(n885), .ZN(n922) );
  AND2_X1 U77bar ( .A1(n886bar), .A2(n885bar), .ZN(n922bar) );
  OR2_X1 U78 ( .A1(n884), .A2(n883), .ZN(n885) );
  AND2_X1 U78bar ( .A1(n884bar), .A2(n883bar), .ZN(n885bar) );
  OR2_X1 U79 ( .A1(n882), .A2(n881), .ZN(n883) );
  AND2_X1 U79bar ( .A1(n882bar), .A2(n881bar), .ZN(n883bar) );
  OR2_X1 U80 ( .A1(in[118]), .A2(in[109]), .ZN(n881) );
  AND2_X1 U80bar ( .A1(inbar[118]), .A2(inbar[109]), .ZN(n881bar) );
  OR2_X1 U81 ( .A1(in[139]), .A2(in[120]), .ZN(n882) );
  AND2_X1 U81bar ( .A1(inbar[139]), .A2(inbar[120]), .ZN(n882bar) );
  OR2_X1 U82 ( .A1(n880), .A2(n879), .ZN(n884) );
  AND2_X1 U82bar ( .A1(n880bar), .A2(n879bar), .ZN(n884bar) );
  OR2_X1 U83 ( .A1(in[198]), .A2(in[154]), .ZN(n879) );
  AND2_X1 U83bar ( .A1(inbar[198]), .A2(inbar[154]), .ZN(n879bar) );
  OR2_X1 U84 ( .A1(in[210]), .A2(in[205]), .ZN(n880) );
  AND2_X1 U84bar ( .A1(inbar[210]), .A2(inbar[205]), .ZN(n880bar) );
  OR2_X1 U85 ( .A1(n878), .A2(n877), .ZN(n886) );
  AND2_X1 U85bar ( .A1(n878bar), .A2(n877bar), .ZN(n886bar) );
  OR2_X1 U86 ( .A1(n876), .A2(n875), .ZN(n877) );
  AND2_X1 U86bar ( .A1(n876bar), .A2(n875bar), .ZN(n877bar) );
  OR2_X1 U87 ( .A1(in[219]), .A2(in[217]), .ZN(n875) );
  AND2_X1 U87bar ( .A1(inbar[219]), .A2(inbar[217]), .ZN(n875bar) );
  OR2_X1 U88 ( .A1(in[86]), .A2(in[252]), .ZN(n876) );
  AND2_X1 U88bar ( .A1(inbar[86]), .A2(inbar[252]), .ZN(n876bar) );
  OR2_X1 U89 ( .A1(n874), .A2(n873), .ZN(n878) );
  AND2_X1 U89bar ( .A1(n874bar), .A2(n873bar), .ZN(n878bar) );
  OR2_X1 U90 ( .A1(in_40), .A2(in[91]), .ZN(n873) );
  AND2_X1 U90bar ( .A1(in_40bar), .A2(inbar[91]), .ZN(n873bar) );
  OR2_X1 U91 ( .A1(in_8), .A2(in_46), .ZN(n874) );
  AND2_X1 U91bar ( .A1(in_8bar), .A2(in_46bar), .ZN(n874bar) );
  OR2_X1 U92 ( .A1(n872), .A2(n871), .ZN(n889) );
  AND2_X1 U92bar ( .A1(n872bar), .A2(n871bar), .ZN(n889bar) );
  OR2_X1 U93 ( .A1(in[117]), .A2(n943), .ZN(n871) );
  AND2_X1 U93bar ( .A1(inbar[117]), .A2(n943bar), .ZN(n871bar) );
  OR2_X1 U94 ( .A1(n870), .A2(n869), .ZN(n943) );
  AND2_X1 U94bar ( .A1(n870bar), .A2(n869bar), .ZN(n943bar) );
  OR2_X1 U95 ( .A1(n868), .A2(n867), .ZN(n869) );
  AND2_X1 U95bar ( .A1(n868bar), .A2(n867bar), .ZN(n869bar) );
  OR2_X1 U96 ( .A1(n866), .A2(n865), .ZN(n867) );
  AND2_X1 U96bar ( .A1(n866bar), .A2(n865bar), .ZN(n867bar) );
  OR2_X1 U97 ( .A1(n864), .A2(n863), .ZN(n865) );
  AND2_X1 U97bar ( .A1(n864bar), .A2(n863bar), .ZN(n865bar) );
  OR2_X1 U98 ( .A1(in[108]), .A2(n919), .ZN(n866) );
  AND2_X1 U98bar ( .A1(inbar[108]), .A2(n919bar), .ZN(n866bar) );
  OR2_X1 U99 ( .A1(n862), .A2(n861), .ZN(n919) );
  AND2_X1 U99bar ( .A1(n862bar), .A2(n861bar), .ZN(n919bar) );
  OR2_X1 U100 ( .A1(n860), .A2(n859), .ZN(n861) );
  AND2_X1 U100bar ( .A1(n860bar), .A2(n859bar), .ZN(n861bar) );
  OR2_X1 U101 ( .A1(n858), .A2(n857), .ZN(n859) );
  AND2_X1 U101bar ( .A1(n858bar), .A2(n857bar), .ZN(n859bar) );
  OR2_X1 U102 ( .A1(in[119]), .A2(in[105]), .ZN(n857) );
  AND2_X1 U102bar ( .A1(inbar[119]), .A2(inbar[105]), .ZN(n857bar) );
  OR2_X1 U103 ( .A1(in[186]), .A2(in[175]), .ZN(n858) );
  AND2_X1 U103bar ( .A1(inbar[186]), .A2(inbar[175]), .ZN(n858bar) );
  OR2_X1 U104 ( .A1(n856), .A2(n855), .ZN(n860) );
  AND2_X1 U104bar ( .A1(n856bar), .A2(n855bar), .ZN(n860bar) );
  OR2_X1 U105 ( .A1(in[202]), .A2(in[193]), .ZN(n855) );
  AND2_X1 U105bar ( .A1(inbar[202]), .A2(inbar[193]), .ZN(n855bar) );
  OR2_X1 U106 ( .A1(in[225]), .A2(in[208]), .ZN(n856) );
  AND2_X1 U106bar ( .A1(inbar[225]), .A2(inbar[208]), .ZN(n856bar) );
  OR2_X1 U107 ( .A1(n854), .A2(n853), .ZN(n862) );
  AND2_X1 U107bar ( .A1(n854bar), .A2(n853bar), .ZN(n862bar) );
  OR2_X1 U108 ( .A1(n852), .A2(n851), .ZN(n853) );
  AND2_X1 U108bar ( .A1(n852bar), .A2(n851bar), .ZN(n853bar) );
  OR2_X1 U109 ( .A1(in_1), .A2(in[85]), .ZN(n851) );
  AND2_X1 U109bar ( .A1(in_1bar), .A2(inbar[85]), .ZN(n851bar) );
  OR2_X1 U110 ( .A1(in_23), .A2(in_19), .ZN(n852) );
  AND2_X1 U110bar ( .A1(in_23bar), .A2(in_19bar), .ZN(n852bar) );
  OR2_X1 U111 ( .A1(n850), .A2(n849), .ZN(n854) );
  AND2_X1 U111bar ( .A1(n850bar), .A2(n849bar), .ZN(n854bar) );
  OR2_X1 U112 ( .A1(in_43), .A2(in_33), .ZN(n849) );
  AND2_X1 U112bar ( .A1(in_43bar), .A2(in_33bar), .ZN(n849bar) );
  OR2_X1 U113 ( .A1(in_63), .A2(in_44), .ZN(n850) );
  AND2_X1 U113bar ( .A1(in_63bar), .A2(in_44bar), .ZN(n850bar) );
  OR2_X1 U114 ( .A1(n848), .A2(n847), .ZN(n868) );
  AND2_X1 U114bar ( .A1(n848bar), .A2(n847bar), .ZN(n868bar) );
  OR2_X1 U115 ( .A1(in[141]), .A2(in[112]), .ZN(n847) );
  AND2_X1 U115bar ( .A1(inbar[141]), .A2(inbar[112]), .ZN(n847bar) );
  OR2_X1 U116 ( .A1(in[147]), .A2(n846), .ZN(n848) );
  AND2_X1 U116bar ( .A1(inbar[147]), .A2(n846bar), .ZN(n848bar) );
  OR2_X1 U117 ( .A1(in[181]), .A2(in[167]), .ZN(n846) );
  AND2_X1 U117bar ( .A1(inbar[181]), .A2(inbar[167]), .ZN(n846bar) );
  OR2_X1 U118 ( .A1(n845), .A2(n844), .ZN(n870) );
  AND2_X1 U118bar ( .A1(n845bar), .A2(n844bar), .ZN(n870bar) );
  OR2_X1 U119 ( .A1(n843), .A2(n842), .ZN(n844) );
  AND2_X1 U119bar ( .A1(n843bar), .A2(n842bar), .ZN(n844bar) );
  OR2_X1 U120 ( .A1(in[229]), .A2(in[201]), .ZN(n842) );
  AND2_X1 U120bar ( .A1(inbar[229]), .A2(inbar[201]), .ZN(n842bar) );
  OR2_X1 U121 ( .A1(in[237]), .A2(n841), .ZN(n843) );
  AND2_X1 U121bar ( .A1(inbar[237]), .A2(n841bar), .ZN(n843bar) );
  OR2_X1 U122 ( .A1(in[94]), .A2(in[253]), .ZN(n841) );
  AND2_X1 U122bar ( .A1(inbar[94]), .A2(inbar[253]), .ZN(n841bar) );
  OR2_X1 U123 ( .A1(n840), .A2(n839), .ZN(n845) );
  AND2_X1 U123bar ( .A1(n840bar), .A2(n839bar), .ZN(n845bar) );
  OR2_X1 U124 ( .A1(in_21), .A2(in[96]), .ZN(n839) );
  AND2_X1 U124bar ( .A1(in_21bar), .A2(inbar[96]), .ZN(n839bar) );
  OR2_X1 U125 ( .A1(in_25), .A2(n838), .ZN(n840) );
  AND2_X1 U125bar ( .A1(in_25bar), .A2(n838bar), .ZN(n840bar) );
  OR2_X1 U126 ( .A1(in_81), .A2(in_45), .ZN(n838) );
  AND2_X1 U126bar ( .A1(in_81bar), .A2(in_45bar), .ZN(n838bar) );
  OR2_X1 U127 ( .A1(n837), .A2(n836), .ZN(n891) );
  AND2_X1 U127bar ( .A1(n837bar), .A2(n836bar), .ZN(n891bar) );
  OR2_X1 U128 ( .A1(in[142]), .A2(in[124]), .ZN(n836) );
  AND2_X1 U128bar ( .A1(inbar[142]), .A2(inbar[124]), .ZN(n836bar) );
  OR2_X1 U129 ( .A1(in[150]), .A2(n835), .ZN(n837) );
  AND2_X1 U129bar ( .A1(inbar[150]), .A2(n835bar), .ZN(n837bar) );
  OR2_X1 U130 ( .A1(in[172]), .A2(in[155]), .ZN(n835) );
  AND2_X1 U130bar ( .A1(inbar[172]), .A2(inbar[155]), .ZN(n835bar) );
  OR2_X1 U131 ( .A1(n834), .A2(n833), .ZN(n893) );
  AND2_X1 U131bar ( .A1(n834bar), .A2(n833bar), .ZN(n893bar) );
  OR2_X1 U132 ( .A1(n832), .A2(n831), .ZN(n833) );
  AND2_X1 U132bar ( .A1(n832bar), .A2(n831bar), .ZN(n833bar) );
  OR2_X1 U133 ( .A1(in[196]), .A2(in[173]), .ZN(n831) );
  AND2_X1 U133bar ( .A1(inbar[196]), .A2(inbar[173]), .ZN(n831bar) );
  OR2_X1 U134 ( .A1(in[222]), .A2(n830), .ZN(n832) );
  AND2_X1 U134bar ( .A1(inbar[222]), .A2(n830bar), .ZN(n832bar) );
  OR2_X1 U135 ( .A1(in[227]), .A2(in[226]), .ZN(n830) );
  AND2_X1 U135bar ( .A1(inbar[227]), .A2(inbar[226]), .ZN(n830bar) );
  OR2_X1 U136 ( .A1(n829), .A2(n828), .ZN(n834) );
  AND2_X1 U136bar ( .A1(n829bar), .A2(n828bar), .ZN(n834bar) );
  OR2_X1 U137 ( .A1(in[249]), .A2(in[231]), .ZN(n828) );
  AND2_X1 U137bar ( .A1(inbar[249]), .A2(inbar[231]), .ZN(n828bar) );
  OR2_X1 U138 ( .A1(in_28), .A2(n827), .ZN(n829) );
  AND2_X1 U138bar ( .A1(in_28bar), .A2(n827bar), .ZN(n829bar) );
  OR2_X1 U139 ( .A1(in_52), .A2(in_47), .ZN(n827) );
  AND2_X1 U139bar ( .A1(in_52bar), .A2(in_47bar), .ZN(n827bar) );
  OR2_X1 U140 ( .A1(n826), .A2(n825), .ZN(out[3]) );
  AND2_X1 U140bar ( .A1(n826bar), .A2(n825bar), .ZN(outbar[3]) );
  OR2_X1 U141 ( .A1(n824), .A2(n823), .ZN(n825) );
  AND2_X1 U141bar ( .A1(n824bar), .A2(n823bar), .ZN(n825bar) );
  OR2_X1 U142 ( .A1(n822), .A2(n821), .ZN(n823) );
  AND2_X1 U142bar ( .A1(n822bar), .A2(n821bar), .ZN(n823bar) );
  OR2_X1 U143 ( .A1(n820), .A2(n819), .ZN(n821) );
  AND2_X1 U143bar ( .A1(n820bar), .A2(n819bar), .ZN(n821bar) );
  OR2_X1 U144 ( .A1(n964), .A2(n818), .ZN(n822) );
  AND2_X1 U144bar ( .A1(n964bar), .A2(n818bar), .ZN(n822bar) );
  OR2_X1 U145 ( .A1(in[118]), .A2(n817), .ZN(n818) );
  AND2_X1 U145bar ( .A1(inbar[118]), .A2(n817bar), .ZN(n818bar) );
  OR2_X1 U146 ( .A1(n816), .A2(n815), .ZN(n964) );
  AND2_X1 U146bar ( .A1(n816bar), .A2(n815bar), .ZN(n964bar) );
  OR2_X1 U147 ( .A1(n814), .A2(n813), .ZN(n815) );
  AND2_X1 U147bar ( .A1(n814bar), .A2(n813bar), .ZN(n815bar) );
  OR2_X1 U148 ( .A1(n812), .A2(n811), .ZN(n813) );
  AND2_X1 U148bar ( .A1(n812bar), .A2(n811bar), .ZN(n813bar) );
  OR2_X1 U149 ( .A1(in[122]), .A2(in[111]), .ZN(n811) );
  AND2_X1 U149bar ( .A1(inbar[122]), .A2(inbar[111]), .ZN(n811bar) );
  OR2_X1 U150 ( .A1(in[154]), .A2(in[151]), .ZN(n812) );
  AND2_X1 U150bar ( .A1(inbar[154]), .A2(inbar[151]), .ZN(n812bar) );
  OR2_X1 U151 ( .A1(n810), .A2(n809), .ZN(n814) );
  AND2_X1 U151bar ( .A1(n810bar), .A2(n809bar), .ZN(n814bar) );
  OR2_X1 U152 ( .A1(in[187]), .A2(in[177]), .ZN(n809) );
  AND2_X1 U152bar ( .A1(inbar[187]), .A2(inbar[177]), .ZN(n809bar) );
  OR2_X1 U153 ( .A1(in[200]), .A2(in[192]), .ZN(n810) );
  AND2_X1 U153bar ( .A1(inbar[200]), .A2(inbar[192]), .ZN(n810bar) );
  OR2_X1 U154 ( .A1(n808), .A2(n807), .ZN(n816) );
  AND2_X1 U154bar ( .A1(n808bar), .A2(n807bar), .ZN(n816bar) );
  OR2_X1 U155 ( .A1(n806), .A2(n805), .ZN(n807) );
  AND2_X1 U155bar ( .A1(n806bar), .A2(n805bar), .ZN(n807bar) );
  OR2_X1 U156 ( .A1(in[225]), .A2(in[207]), .ZN(n805) );
  AND2_X1 U156bar ( .A1(inbar[225]), .A2(inbar[207]), .ZN(n805bar) );
  OR2_X1 U157 ( .A1(in[98]), .A2(in[226]), .ZN(n806) );
  AND2_X1 U157bar ( .A1(inbar[98]), .A2(inbar[226]), .ZN(n806bar) );
  OR2_X1 U158 ( .A1(n804), .A2(n803), .ZN(n808) );
  AND2_X1 U158bar ( .A1(n804bar), .A2(n803bar), .ZN(n808bar) );
  OR2_X1 U159 ( .A1(in_20), .A2(in_16), .ZN(n803) );
  AND2_X1 U159bar ( .A1(in_20bar), .A2(in_16bar), .ZN(n803bar) );
  OR2_X1 U160 ( .A1(in_55), .A2(in_45), .ZN(n804) );
  AND2_X1 U160bar ( .A1(in_55bar), .A2(in_45bar), .ZN(n804bar) );
  OR2_X1 U161 ( .A1(n802), .A2(n801), .ZN(n824) );
  AND2_X1 U161bar ( .A1(n802bar), .A2(n801bar), .ZN(n824bar) );
  OR2_X1 U162 ( .A1(in[162]), .A2(in[149]), .ZN(n801) );
  AND2_X1 U162bar ( .A1(inbar[162]), .A2(inbar[149]), .ZN(n801bar) );
  OR2_X1 U163 ( .A1(in[163]), .A2(n800), .ZN(n802) );
  AND2_X1 U163bar ( .A1(inbar[163]), .A2(n800bar), .ZN(n802bar) );
  OR2_X1 U164 ( .A1(in[191]), .A2(in[189]), .ZN(n800) );
  AND2_X1 U164bar ( .A1(inbar[191]), .A2(inbar[189]), .ZN(n800bar) );
  OR2_X1 U165 ( .A1(n799), .A2(n798), .ZN(n826) );
  AND2_X1 U165bar ( .A1(n799bar), .A2(n798bar), .ZN(n826bar) );
  OR2_X1 U166 ( .A1(n797), .A2(n796), .ZN(n798) );
  AND2_X1 U166bar ( .A1(n797bar), .A2(n796bar), .ZN(n798bar) );
  OR2_X1 U167 ( .A1(in[212]), .A2(in[193]), .ZN(n796) );
  AND2_X1 U167bar ( .A1(inbar[212]), .A2(inbar[193]), .ZN(n796bar) );
  OR2_X1 U168 ( .A1(in[238]), .A2(n795), .ZN(n797) );
  AND2_X1 U168bar ( .A1(inbar[238]), .A2(n795bar), .ZN(n797bar) );
  OR2_X1 U169 ( .A1(in[88]), .A2(in[247]), .ZN(n795) );
  AND2_X1 U169bar ( .A1(inbar[88]), .A2(inbar[247]), .ZN(n795bar) );
  OR2_X1 U170 ( .A1(n794), .A2(n793), .ZN(n799) );
  AND2_X1 U170bar ( .A1(n794bar), .A2(n793bar), .ZN(n799bar) );
  OR2_X1 U171 ( .A1(in[94]), .A2(in[92]), .ZN(n793) );
  AND2_X1 U171bar ( .A1(inbar[94]), .A2(inbar[92]), .ZN(n793bar) );
  OR2_X1 U172 ( .A1(in_52), .A2(n792), .ZN(n794) );
  AND2_X1 U172bar ( .A1(in_52bar), .A2(n792bar), .ZN(n794bar) );
  OR2_X1 U173 ( .A1(in_70), .A2(in_67), .ZN(n792) );
  AND2_X1 U173bar ( .A1(in_70bar), .A2(in_67bar), .ZN(n792bar) );
  OR2_X1 U174 ( .A1(n791), .A2(n790), .ZN(out[2]) );
  AND2_X1 U174bar ( .A1(n791bar), .A2(n790bar), .ZN(outbar[2]) );
  OR2_X1 U175 ( .A1(n789), .A2(n788), .ZN(n790) );
  AND2_X1 U175bar ( .A1(n789bar), .A2(n788bar), .ZN(n790bar) );
  OR2_X1 U176 ( .A1(n787), .A2(n786), .ZN(n788) );
  AND2_X1 U176bar ( .A1(n787bar), .A2(n786bar), .ZN(n788bar) );
  OR2_X1 U177 ( .A1(n819), .A2(n785), .ZN(n786) );
  AND2_X1 U177bar ( .A1(n819bar), .A2(n785bar), .ZN(n786bar) );
  OR2_X1 U178 ( .A1(n784), .A2(n783), .ZN(n819) );
  AND2_X1 U178bar ( .A1(n784bar), .A2(n783bar), .ZN(n819bar) );
  OR2_X1 U179 ( .A1(n782), .A2(n781), .ZN(n783) );
  AND2_X1 U179bar ( .A1(n782bar), .A2(n781bar), .ZN(n783bar) );
  OR2_X1 U180 ( .A1(n780), .A2(n779), .ZN(n781) );
  AND2_X1 U180bar ( .A1(n780bar), .A2(n779bar), .ZN(n781bar) );
  OR2_X1 U181 ( .A1(n962), .A2(n778), .ZN(n779) );
  AND2_X1 U181bar ( .A1(n962bar), .A2(n778bar), .ZN(n779bar) );
  OR2_X1 U182 ( .A1(n777), .A2(n776), .ZN(n962) );
  AND2_X1 U182bar ( .A1(n777bar), .A2(n776bar), .ZN(n962bar) );
  OR2_X1 U183 ( .A1(n775), .A2(n774), .ZN(n776) );
  AND2_X1 U183bar ( .A1(n775bar), .A2(n774bar), .ZN(n776bar) );
  OR2_X1 U184 ( .A1(n773), .A2(n772), .ZN(n774) );
  AND2_X1 U184bar ( .A1(n773bar), .A2(n772bar), .ZN(n774bar) );
  OR2_X1 U185 ( .A1(in[131]), .A2(in[120]), .ZN(n772) );
  AND2_X1 U185bar ( .A1(inbar[131]), .A2(inbar[120]), .ZN(n772bar) );
  OR2_X1 U186 ( .A1(in[153]), .A2(in[147]), .ZN(n773) );
  AND2_X1 U186bar ( .A1(inbar[153]), .A2(inbar[147]), .ZN(n773bar) );
  OR2_X1 U187 ( .A1(n771), .A2(n770), .ZN(n775) );
  AND2_X1 U187bar ( .A1(n771bar), .A2(n770bar), .ZN(n775bar) );
  OR2_X1 U188 ( .A1(in[170]), .A2(in[156]), .ZN(n770) );
  AND2_X1 U188bar ( .A1(inbar[170]), .A2(inbar[156]), .ZN(n770bar) );
  OR2_X1 U189 ( .A1(in[223]), .A2(in[190]), .ZN(n771) );
  AND2_X1 U189bar ( .A1(inbar[223]), .A2(inbar[190]), .ZN(n771bar) );
  OR2_X1 U190 ( .A1(n769), .A2(n768), .ZN(n777) );
  AND2_X1 U190bar ( .A1(n769bar), .A2(n768bar), .ZN(n777bar) );
  OR2_X1 U191 ( .A1(n767), .A2(n766), .ZN(n768) );
  AND2_X1 U191bar ( .A1(n767bar), .A2(n766bar), .ZN(n768bar) );
  OR2_X1 U192 ( .A1(in[236]), .A2(in[230]), .ZN(n766) );
  AND2_X1 U192bar ( .A1(inbar[236]), .A2(inbar[230]), .ZN(n766bar) );
  OR2_X1 U193 ( .A1(in[85]), .A2(in[240]), .ZN(n767) );
  AND2_X1 U193bar ( .A1(inbar[85]), .A2(inbar[240]), .ZN(n767bar) );
  OR2_X1 U194 ( .A1(n765), .A2(n764), .ZN(n769) );
  AND2_X1 U194bar ( .A1(n765bar), .A2(n764bar), .ZN(n769bar) );
  OR2_X1 U195 ( .A1(in_12), .A2(in[90]), .ZN(n764) );
  AND2_X1 U195bar ( .A1(in_12bar), .A2(inbar[90]), .ZN(n764bar) );
  OR2_X1 U196 ( .A1(in_39), .A2(in_28), .ZN(n765) );
  AND2_X1 U196bar ( .A1(in_39bar), .A2(in_28bar), .ZN(n765bar) );
  OR2_X1 U197 ( .A1(in[109]), .A2(n763), .ZN(n780) );
  AND2_X1 U197bar ( .A1(inbar[109]), .A2(n763bar), .ZN(n780bar) );
  OR2_X1 U198 ( .A1(n762), .A2(n761), .ZN(n782) );
  AND2_X1 U198bar ( .A1(n762bar), .A2(n761bar), .ZN(n782bar) );
  OR2_X1 U199 ( .A1(in[138]), .A2(in[129]), .ZN(n761) );
  AND2_X1 U199bar ( .A1(inbar[138]), .A2(inbar[129]), .ZN(n761bar) );
  OR2_X1 U200 ( .A1(in[157]), .A2(n760), .ZN(n762) );
  AND2_X1 U200bar ( .A1(inbar[157]), .A2(n760bar), .ZN(n762bar) );
  OR2_X1 U201 ( .A1(in[182]), .A2(in[167]), .ZN(n760) );
  AND2_X1 U201bar ( .A1(inbar[182]), .A2(inbar[167]), .ZN(n760bar) );
  OR2_X1 U202 ( .A1(n759), .A2(n758), .ZN(n784) );
  AND2_X1 U202bar ( .A1(n759bar), .A2(n758bar), .ZN(n784bar) );
  OR2_X1 U203 ( .A1(n757), .A2(n756), .ZN(n758) );
  AND2_X1 U203bar ( .A1(n757bar), .A2(n756bar), .ZN(n758bar) );
  OR2_X1 U204 ( .A1(in[195]), .A2(in[184]), .ZN(n756) );
  AND2_X1 U204bar ( .A1(inbar[195]), .A2(inbar[184]), .ZN(n756bar) );
  OR2_X1 U205 ( .A1(in[196]), .A2(n755), .ZN(n757) );
  AND2_X1 U205bar ( .A1(inbar[196]), .A2(n755bar), .ZN(n757bar) );
  OR2_X1 U206 ( .A1(in[215]), .A2(in[209]), .ZN(n755) );
  AND2_X1 U206bar ( .A1(inbar[215]), .A2(inbar[209]), .ZN(n755bar) );
  OR2_X1 U207 ( .A1(n754), .A2(n753), .ZN(n759) );
  AND2_X1 U207bar ( .A1(n754bar), .A2(n753bar), .ZN(n759bar) );
  OR2_X1 U208 ( .A1(in[93]), .A2(in[233]), .ZN(n753) );
  AND2_X1 U208bar ( .A1(inbar[93]), .A2(inbar[233]), .ZN(n753bar) );
  OR2_X1 U209 ( .A1(in_1), .A2(n752), .ZN(n754) );
  AND2_X1 U209bar ( .A1(in_1bar), .A2(n752bar), .ZN(n754bar) );
  OR2_X1 U210 ( .A1(in_69), .A2(in_66), .ZN(n752) );
  AND2_X1 U210bar ( .A1(in_69bar), .A2(in_66bar), .ZN(n752bar) );
  OR2_X1 U211 ( .A1(n966), .A2(n751), .ZN(n787) );
  AND2_X1 U211bar ( .A1(n966bar), .A2(n751bar), .ZN(n787bar) );
  OR2_X1 U212 ( .A1(in[134]), .A2(n750), .ZN(n751) );
  AND2_X1 U212bar ( .A1(inbar[134]), .A2(n750bar), .ZN(n751bar) );
  OR2_X1 U213 ( .A1(n749), .A2(n748), .ZN(n966) );
  AND2_X1 U213bar ( .A1(n749bar), .A2(n748bar), .ZN(n966bar) );
  OR2_X1 U214 ( .A1(n747), .A2(n746), .ZN(n748) );
  AND2_X1 U214bar ( .A1(n747bar), .A2(n746bar), .ZN(n748bar) );
  OR2_X1 U215 ( .A1(n745), .A2(n744), .ZN(n746) );
  AND2_X1 U215bar ( .A1(n745bar), .A2(n744bar), .ZN(n746bar) );
  OR2_X1 U216 ( .A1(in[136]), .A2(in[121]), .ZN(n744) );
  AND2_X1 U216bar ( .A1(inbar[136]), .A2(inbar[121]), .ZN(n744bar) );
  OR2_X1 U217 ( .A1(in[186]), .A2(in[174]), .ZN(n745) );
  AND2_X1 U217bar ( .A1(inbar[186]), .A2(inbar[174]), .ZN(n745bar) );
  OR2_X1 U218 ( .A1(n743), .A2(n742), .ZN(n747) );
  AND2_X1 U218bar ( .A1(n743bar), .A2(n742bar), .ZN(n747bar) );
  OR2_X1 U219 ( .A1(in[198]), .A2(in[197]), .ZN(n742) );
  AND2_X1 U219bar ( .A1(inbar[198]), .A2(inbar[197]), .ZN(n742bar) );
  OR2_X1 U220 ( .A1(in[214]), .A2(in[199]), .ZN(n743) );
  AND2_X1 U220bar ( .A1(inbar[214]), .A2(inbar[199]), .ZN(n743bar) );
  OR2_X1 U221 ( .A1(n741), .A2(n740), .ZN(n749) );
  AND2_X1 U221bar ( .A1(n741bar), .A2(n740bar), .ZN(n749bar) );
  OR2_X1 U222 ( .A1(n739), .A2(n738), .ZN(n740) );
  AND2_X1 U222bar ( .A1(n739bar), .A2(n738bar), .ZN(n740bar) );
  OR2_X1 U223 ( .A1(in[231]), .A2(in[220]), .ZN(n738) );
  AND2_X1 U223bar ( .A1(inbar[231]), .A2(inbar[220]), .ZN(n738bar) );
  OR2_X1 U224 ( .A1(in_25), .A2(in[245]), .ZN(n739) );
  AND2_X1 U224bar ( .A1(in_25bar), .A2(inbar[245]), .ZN(n739bar) );
  OR2_X1 U225 ( .A1(n737), .A2(n736), .ZN(n741) );
  AND2_X1 U225bar ( .A1(n737bar), .A2(n736bar), .ZN(n741bar) );
  OR2_X1 U226 ( .A1(in_53), .A2(in_29), .ZN(n736) );
  AND2_X1 U226bar ( .A1(in_53bar), .A2(in_29bar), .ZN(n736bar) );
  OR2_X1 U227 ( .A1(in_79), .A2(in_74), .ZN(n737) );
  AND2_X1 U227bar ( .A1(in_79bar), .A2(in_74bar), .ZN(n737bar) );
  OR2_X1 U228 ( .A1(n735), .A2(n734), .ZN(n789) );
  AND2_X1 U228bar ( .A1(n735bar), .A2(n734bar), .ZN(n789bar) );
  OR2_X1 U229 ( .A1(in[152]), .A2(in[140]), .ZN(n734) );
  AND2_X1 U229bar ( .A1(inbar[152]), .A2(inbar[140]), .ZN(n734bar) );
  OR2_X1 U230 ( .A1(in[155]), .A2(n733), .ZN(n735) );
  AND2_X1 U230bar ( .A1(inbar[155]), .A2(n733bar), .ZN(n735bar) );
  OR2_X1 U231 ( .A1(in[166]), .A2(in[165]), .ZN(n733) );
  AND2_X1 U231bar ( .A1(inbar[166]), .A2(inbar[165]), .ZN(n733bar) );
  OR2_X1 U232 ( .A1(n732), .A2(n731), .ZN(n791) );
  AND2_X1 U232bar ( .A1(n732bar), .A2(n731bar), .ZN(n791bar) );
  OR2_X1 U233 ( .A1(n730), .A2(n729), .ZN(n731) );
  AND2_X1 U233bar ( .A1(n730bar), .A2(n729bar), .ZN(n731bar) );
  OR2_X1 U234 ( .A1(in[202]), .A2(in[185]), .ZN(n729) );
  AND2_X1 U234bar ( .A1(inbar[202]), .A2(inbar[185]), .ZN(n729bar) );
  OR2_X1 U235 ( .A1(in[211]), .A2(n728), .ZN(n730) );
  AND2_X1 U235bar ( .A1(inbar[211]), .A2(n728bar), .ZN(n730bar) );
  OR2_X1 U236 ( .A1(in[255]), .A2(in[253]), .ZN(n728) );
  AND2_X1 U236bar ( .A1(inbar[255]), .A2(inbar[253]), .ZN(n728bar) );
  OR2_X1 U237 ( .A1(n727), .A2(n726), .ZN(n732) );
  AND2_X1 U237bar ( .A1(n727bar), .A2(n726bar), .ZN(n732bar) );
  OR2_X1 U238 ( .A1(in_35), .A2(in_15), .ZN(n726) );
  AND2_X1 U238bar ( .A1(in_35bar), .A2(in_15bar), .ZN(n726bar) );
  OR2_X1 U239 ( .A1(in_36), .A2(n725), .ZN(n727) );
  AND2_X1 U239bar ( .A1(in_36bar), .A2(n725bar), .ZN(n727bar) );
  OR2_X1 U240 ( .A1(in_48), .A2(in_40), .ZN(n725) );
  AND2_X1 U240bar ( .A1(in_48bar), .A2(in_40bar), .ZN(n725bar) );
  OR2_X1 U241 ( .A1(n724), .A2(n723), .ZN(out[1]) );
  AND2_X1 U241bar ( .A1(n724bar), .A2(n723bar), .ZN(outbar[1]) );
  OR2_X1 U242 ( .A1(n722), .A2(n721), .ZN(n723) );
  AND2_X1 U242bar ( .A1(n722bar), .A2(n721bar), .ZN(n723bar) );
  OR2_X1 U243 ( .A1(n720), .A2(n719), .ZN(n721) );
  AND2_X1 U243bar ( .A1(n720bar), .A2(n719bar), .ZN(n721bar) );
  OR2_X1 U244 ( .A1(n921), .A2(n887), .ZN(n719) );
  AND2_X1 U244bar ( .A1(n921bar), .A2(n887bar), .ZN(n719bar) );
  OR2_X1 U245 ( .A1(n718), .A2(n717), .ZN(n887) );
  AND2_X1 U245bar ( .A1(n718bar), .A2(n717bar), .ZN(n887bar) );
  OR2_X1 U246 ( .A1(n716), .A2(n715), .ZN(n717) );
  AND2_X1 U246bar ( .A1(n716bar), .A2(n715bar), .ZN(n717bar) );
  OR2_X1 U247 ( .A1(n714), .A2(n713), .ZN(n715) );
  AND2_X1 U247bar ( .A1(n714bar), .A2(n713bar), .ZN(n715bar) );
  OR2_X1 U248 ( .A1(in[116]), .A2(in[110]), .ZN(n713) );
  AND2_X1 U248bar ( .A1(inbar[116]), .A2(inbar[110]), .ZN(n713bar) );
  OR2_X1 U249 ( .A1(in[133]), .A2(in[130]), .ZN(n714) );
  AND2_X1 U249bar ( .A1(inbar[133]), .A2(inbar[130]), .ZN(n714bar) );
  OR2_X1 U250 ( .A1(n712), .A2(n711), .ZN(n716) );
  AND2_X1 U250bar ( .A1(n712bar), .A2(n711bar), .ZN(n716bar) );
  OR2_X1 U251 ( .A1(in[203]), .A2(in[135]), .ZN(n711) );
  AND2_X1 U251bar ( .A1(inbar[203]), .A2(inbar[135]), .ZN(n711bar) );
  OR2_X1 U252 ( .A1(in[232]), .A2(in[223]), .ZN(n712) );
  AND2_X1 U252bar ( .A1(inbar[232]), .A2(inbar[223]), .ZN(n712bar) );
  OR2_X1 U253 ( .A1(n710), .A2(n709), .ZN(n718) );
  AND2_X1 U253bar ( .A1(n710bar), .A2(n709bar), .ZN(n718bar) );
  OR2_X1 U254 ( .A1(n708), .A2(n707), .ZN(n709) );
  AND2_X1 U254bar ( .A1(n708bar), .A2(n707bar), .ZN(n709bar) );
  OR2_X1 U255 ( .A1(in[255]), .A2(in[233]), .ZN(n707) );
  AND2_X1 U255bar ( .A1(inbar[255]), .A2(inbar[233]), .ZN(n707bar) );
  OR2_X1 U256 ( .A1(in_53), .A2(in_34), .ZN(n708) );
  AND2_X1 U256bar ( .A1(in_53bar), .A2(in_34bar), .ZN(n708bar) );
  OR2_X1 U257 ( .A1(n706), .A2(n705), .ZN(n710) );
  AND2_X1 U257bar ( .A1(n706bar), .A2(n705bar), .ZN(n710bar) );
  OR2_X1 U258 ( .A1(in_57), .A2(in_55), .ZN(n705) );
  AND2_X1 U258bar ( .A1(in_57bar), .A2(in_55bar), .ZN(n705bar) );
  OR2_X1 U259 ( .A1(in_68), .A2(in_67), .ZN(n706) );
  AND2_X1 U259bar ( .A1(in_68bar), .A2(in_67bar), .ZN(n706bar) );
  OR2_X1 U260 ( .A1(n704), .A2(n703), .ZN(n921) );
  AND2_X1 U260bar ( .A1(n704bar), .A2(n703bar), .ZN(n921bar) );
  OR2_X1 U261 ( .A1(n702), .A2(n701), .ZN(n703) );
  AND2_X1 U261bar ( .A1(n702bar), .A2(n701bar), .ZN(n703bar) );
  OR2_X1 U262 ( .A1(n700), .A2(n699), .ZN(n701) );
  AND2_X1 U262bar ( .A1(n700bar), .A2(n699bar), .ZN(n701bar) );
  OR2_X1 U263 ( .A1(n944), .A2(n872), .ZN(n699) );
  AND2_X1 U263bar ( .A1(n944bar), .A2(n872bar), .ZN(n699bar) );
  OR2_X1 U264 ( .A1(n698), .A2(n697), .ZN(n872) );
  AND2_X1 U264bar ( .A1(n698bar), .A2(n697bar), .ZN(n872bar) );
  OR2_X1 U265 ( .A1(n696), .A2(n695), .ZN(n697) );
  AND2_X1 U265bar ( .A1(n696bar), .A2(n695bar), .ZN(n697bar) );
  OR2_X1 U266 ( .A1(n694), .A2(n693), .ZN(n695) );
  AND2_X1 U266bar ( .A1(n694bar), .A2(n693bar), .ZN(n695bar) );
  OR2_X1 U267 ( .A1(in[121]), .A2(in[102]), .ZN(n693) );
  AND2_X1 U267bar ( .A1(inbar[121]), .A2(inbar[102]), .ZN(n693bar) );
  OR2_X1 U268 ( .A1(in[162]), .A2(in[161]), .ZN(n694) );
  AND2_X1 U268bar ( .A1(inbar[162]), .A2(inbar[161]), .ZN(n694bar) );
  OR2_X1 U269 ( .A1(n692), .A2(n691), .ZN(n696) );
  AND2_X1 U269bar ( .A1(n692bar), .A2(n691bar), .ZN(n696bar) );
  OR2_X1 U270 ( .A1(in[192]), .A2(in[178]), .ZN(n691) );
  AND2_X1 U270bar ( .A1(inbar[192]), .A2(inbar[178]), .ZN(n691bar) );
  OR2_X1 U271 ( .A1(in[244]), .A2(in[209]), .ZN(n692) );
  AND2_X1 U271bar ( .A1(inbar[244]), .A2(inbar[209]), .ZN(n692bar) );
  OR2_X1 U272 ( .A1(n690), .A2(n689), .ZN(n698) );
  AND2_X1 U272bar ( .A1(n690bar), .A2(n689bar), .ZN(n698bar) );
  OR2_X1 U273 ( .A1(n688), .A2(n687), .ZN(n689) );
  AND2_X1 U273bar ( .A1(n688bar), .A2(n687bar), .ZN(n689bar) );
  OR2_X1 U274 ( .A1(in[90]), .A2(in[254]), .ZN(n687) );
  AND2_X1 U274bar ( .A1(inbar[90]), .A2(inbar[254]), .ZN(n687bar) );
  OR2_X1 U275 ( .A1(in_36), .A2(in_32), .ZN(n688) );
  AND2_X1 U275bar ( .A1(in_36bar), .A2(in_32bar), .ZN(n688bar) );
  OR2_X1 U276 ( .A1(n686), .A2(n685), .ZN(n690) );
  AND2_X1 U276bar ( .A1(n686bar), .A2(n685bar), .ZN(n690bar) );
  OR2_X1 U277 ( .A1(in_62), .A2(in_37), .ZN(n685) );
  AND2_X1 U277bar ( .A1(in_62bar), .A2(in_37bar), .ZN(n685bar) );
  OR2_X1 U278 ( .A1(in_75), .A2(in_73), .ZN(n686) );
  AND2_X1 U278bar ( .A1(in_75bar), .A2(in_73bar), .ZN(n686bar) );
  OR2_X1 U279 ( .A1(n684), .A2(n683), .ZN(n944) );
  AND2_X1 U279bar ( .A1(n684bar), .A2(n683bar), .ZN(n944bar) );
  OR2_X1 U280 ( .A1(n682), .A2(n681), .ZN(n683) );
  AND2_X1 U280bar ( .A1(n682bar), .A2(n681bar), .ZN(n683bar) );
  OR2_X1 U281 ( .A1(n680), .A2(n679), .ZN(n681) );
  AND2_X1 U281bar ( .A1(n680bar), .A2(n679bar), .ZN(n681bar) );
  OR2_X1 U282 ( .A1(in[171]), .A2(in[153]), .ZN(n679) );
  AND2_X1 U282bar ( .A1(inbar[171]), .A2(inbar[153]), .ZN(n679bar) );
  OR2_X1 U283 ( .A1(in[187]), .A2(in[176]), .ZN(n680) );
  AND2_X1 U283bar ( .A1(inbar[187]), .A2(inbar[176]), .ZN(n680bar) );
  OR2_X1 U284 ( .A1(n678), .A2(n677), .ZN(n682) );
  AND2_X1 U284bar ( .A1(n678bar), .A2(n677bar), .ZN(n682bar) );
  OR2_X1 U285 ( .A1(in[245]), .A2(in[211]), .ZN(n677) );
  AND2_X1 U285bar ( .A1(inbar[245]), .A2(inbar[211]), .ZN(n677bar) );
  OR2_X1 U286 ( .A1(in[97]), .A2(in[88]), .ZN(n678) );
  AND2_X1 U286bar ( .A1(inbar[97]), .A2(inbar[88]), .ZN(n678bar) );
  OR2_X1 U287 ( .A1(n676), .A2(n675), .ZN(n684) );
  AND2_X1 U287bar ( .A1(n676bar), .A2(n675bar), .ZN(n684bar) );
  OR2_X1 U288 ( .A1(n674), .A2(n673), .ZN(n675) );
  AND2_X1 U288bar ( .A1(n674bar), .A2(n673bar), .ZN(n675bar) );
  OR2_X1 U289 ( .A1(in_10), .A2(in_0), .ZN(n673) );
  AND2_X1 U289bar ( .A1(in_10bar), .A2(in_0bar), .ZN(n673bar) );
  OR2_X1 U290 ( .A1(in_59), .A2(in_5), .ZN(n674) );
  AND2_X1 U290bar ( .A1(in_59bar), .A2(in_5bar), .ZN(n674bar) );
  OR2_X1 U291 ( .A1(n672), .A2(n671), .ZN(n676) );
  AND2_X1 U291bar ( .A1(n672bar), .A2(n671bar), .ZN(n676bar) );
  OR2_X1 U292 ( .A1(in_60), .A2(in_6), .ZN(n671) );
  AND2_X1 U292bar ( .A1(in_60bar), .A2(in_6bar), .ZN(n671bar) );
  OR2_X1 U293 ( .A1(in_77), .A2(in_69), .ZN(n672) );
  AND2_X1 U293bar ( .A1(in_77bar), .A2(in_69bar), .ZN(n672bar) );
  OR2_X1 U294 ( .A1(in[113]), .A2(n864), .ZN(n700) );
  AND2_X1 U294bar ( .A1(inbar[113]), .A2(n864bar), .ZN(n700bar) );
  OR2_X1 U295 ( .A1(n670), .A2(n669), .ZN(n864) );
  AND2_X1 U295bar ( .A1(n670bar), .A2(n669bar), .ZN(n864bar) );
  OR2_X1 U296 ( .A1(n668), .A2(n667), .ZN(n669) );
  AND2_X1 U296bar ( .A1(n668bar), .A2(n667bar), .ZN(n669bar) );
  OR2_X1 U297 ( .A1(n666), .A2(n665), .ZN(n667) );
  AND2_X1 U297bar ( .A1(n666bar), .A2(n665bar), .ZN(n667bar) );
  OR2_X1 U298 ( .A1(in[125]), .A2(in[107]), .ZN(n665) );
  AND2_X1 U298bar ( .A1(inbar[125]), .A2(inbar[107]), .ZN(n665bar) );
  OR2_X1 U299 ( .A1(in[138]), .A2(in[126]), .ZN(n666) );
  AND2_X1 U299bar ( .A1(inbar[138]), .A2(inbar[126]), .ZN(n666bar) );
  OR2_X1 U300 ( .A1(n664), .A2(n663), .ZN(n668) );
  AND2_X1 U300bar ( .A1(n664bar), .A2(n663bar), .ZN(n668bar) );
  OR2_X1 U301 ( .A1(in[189]), .A2(in[143]), .ZN(n663) );
  AND2_X1 U301bar ( .A1(inbar[189]), .A2(inbar[143]), .ZN(n663bar) );
  OR2_X1 U302 ( .A1(in[99]), .A2(in[214]), .ZN(n664) );
  AND2_X1 U302bar ( .A1(inbar[99]), .A2(inbar[214]), .ZN(n664bar) );
  OR2_X1 U303 ( .A1(n662), .A2(n661), .ZN(n670) );
  AND2_X1 U303bar ( .A1(n662bar), .A2(n661bar), .ZN(n670bar) );
  OR2_X1 U304 ( .A1(n660), .A2(n659), .ZN(n661) );
  AND2_X1 U304bar ( .A1(n660bar), .A2(n659bar), .ZN(n661bar) );
  OR2_X1 U305 ( .A1(in_15), .A2(in_12), .ZN(n659) );
  AND2_X1 U305bar ( .A1(in_15bar), .A2(in_12bar), .ZN(n659bar) );
  OR2_X1 U306 ( .A1(in_20), .A2(in_2), .ZN(n660) );
  AND2_X1 U306bar ( .A1(in_20bar), .A2(in_2bar), .ZN(n660bar) );
  OR2_X1 U307 ( .A1(n658), .A2(n657), .ZN(n662) );
  AND2_X1 U307bar ( .A1(n658bar), .A2(n657bar), .ZN(n662bar) );
  OR2_X1 U308 ( .A1(in_30), .A2(in_3), .ZN(n657) );
  AND2_X1 U308bar ( .A1(in_30bar), .A2(in_3bar), .ZN(n657bar) );
  OR2_X1 U309 ( .A1(in_4), .A2(in_38), .ZN(n658) );
  AND2_X1 U309bar ( .A1(in_4bar), .A2(in_38bar), .ZN(n658bar) );
  OR2_X1 U310 ( .A1(n656), .A2(n655), .ZN(n702) );
  AND2_X1 U310bar ( .A1(n656bar), .A2(n655bar), .ZN(n702bar) );
  OR2_X1 U311 ( .A1(in[148]), .A2(in[137]), .ZN(n655) );
  AND2_X1 U311bar ( .A1(inbar[148]), .A2(inbar[137]), .ZN(n655bar) );
  OR2_X1 U312 ( .A1(in[149]), .A2(n654), .ZN(n656) );
  AND2_X1 U312bar ( .A1(inbar[149]), .A2(n654bar), .ZN(n656bar) );
  OR2_X1 U313 ( .A1(in[195]), .A2(in[190]), .ZN(n654) );
  AND2_X1 U313bar ( .A1(inbar[195]), .A2(inbar[190]), .ZN(n654bar) );
  OR2_X1 U314 ( .A1(n653), .A2(n652), .ZN(n704) );
  AND2_X1 U314bar ( .A1(n653bar), .A2(n652bar), .ZN(n704bar) );
  OR2_X1 U315 ( .A1(n651), .A2(n650), .ZN(n652) );
  AND2_X1 U315bar ( .A1(n651bar), .A2(n650bar), .ZN(n652bar) );
  OR2_X1 U316 ( .A1(in[98]), .A2(in[197]), .ZN(n650) );
  AND2_X1 U316bar ( .A1(inbar[98]), .A2(inbar[197]), .ZN(n650bar) );
  OR2_X1 U317 ( .A1(in_11), .A2(n649), .ZN(n651) );
  AND2_X1 U317bar ( .A1(in_11bar), .A2(n649bar), .ZN(n651bar) );
  OR2_X1 U318 ( .A1(in_26), .A2(in_14), .ZN(n649) );
  AND2_X1 U318bar ( .A1(in_26bar), .A2(in_14bar), .ZN(n649bar) );
  OR2_X1 U319 ( .A1(n648), .A2(n647), .ZN(n653) );
  AND2_X1 U319bar ( .A1(n648bar), .A2(n647bar), .ZN(n653bar) );
  OR2_X1 U320 ( .A1(in_35), .A2(in_27), .ZN(n647) );
  AND2_X1 U320bar ( .A1(in_35bar), .A2(in_27bar), .ZN(n647bar) );
  OR2_X1 U321 ( .A1(in_50), .A2(n646), .ZN(n648) );
  AND2_X1 U321bar ( .A1(in_50bar), .A2(n646bar), .ZN(n648bar) );
  OR2_X1 U322 ( .A1(in_78), .A2(in_61), .ZN(n646) );
  AND2_X1 U322bar ( .A1(in_78bar), .A2(in_61bar), .ZN(n646bar) );
  OR2_X1 U323 ( .A1(n942), .A2(n645), .ZN(n720) );
  AND2_X1 U323bar ( .A1(n942bar), .A2(n645bar), .ZN(n720bar) );
  OR2_X1 U324 ( .A1(in[106]), .A2(n863), .ZN(n645) );
  AND2_X1 U324bar ( .A1(inbar[106]), .A2(n863bar), .ZN(n645bar) );
  OR2_X1 U325 ( .A1(n644), .A2(n643), .ZN(n863) );
  AND2_X1 U325bar ( .A1(n644bar), .A2(n643bar), .ZN(n863bar) );
  OR2_X1 U326 ( .A1(n642), .A2(n641), .ZN(n643) );
  AND2_X1 U326bar ( .A1(n642bar), .A2(n641bar), .ZN(n643bar) );
  OR2_X1 U327 ( .A1(n640), .A2(n639), .ZN(n641) );
  AND2_X1 U327bar ( .A1(n640bar), .A2(n639bar), .ZN(n641bar) );
  OR2_X1 U328 ( .A1(in[127]), .A2(in[122]), .ZN(n639) );
  AND2_X1 U328bar ( .A1(inbar[127]), .A2(inbar[122]), .ZN(n639bar) );
  OR2_X1 U329 ( .A1(in[156]), .A2(in[132]), .ZN(n640) );
  AND2_X1 U329bar ( .A1(inbar[156]), .A2(inbar[132]), .ZN(n640bar) );
  OR2_X1 U330 ( .A1(n638), .A2(n637), .ZN(n642) );
  AND2_X1 U330bar ( .A1(n638bar), .A2(n637bar), .ZN(n642bar) );
  OR2_X1 U331 ( .A1(in[159]), .A2(in[157]), .ZN(n637) );
  AND2_X1 U331bar ( .A1(inbar[159]), .A2(inbar[157]), .ZN(n637bar) );
  OR2_X1 U332 ( .A1(in[185]), .A2(in[169]), .ZN(n638) );
  AND2_X1 U332bar ( .A1(inbar[185]), .A2(inbar[169]), .ZN(n638bar) );
  OR2_X1 U333 ( .A1(n636), .A2(n635), .ZN(n644) );
  AND2_X1 U333bar ( .A1(n636bar), .A2(n635bar), .ZN(n644bar) );
  OR2_X1 U334 ( .A1(n634), .A2(n633), .ZN(n635) );
  AND2_X1 U334bar ( .A1(n634bar), .A2(n633bar), .ZN(n635bar) );
  OR2_X1 U335 ( .A1(in[239]), .A2(in[218]), .ZN(n633) );
  AND2_X1 U335bar ( .A1(inbar[239]), .A2(inbar[218]), .ZN(n633bar) );
  OR2_X1 U336 ( .A1(in_13), .A2(in[87]), .ZN(n634) );
  AND2_X1 U336bar ( .A1(in_13bar), .A2(inbar[87]), .ZN(n634bar) );
  OR2_X1 U337 ( .A1(n632), .A2(n631), .ZN(n636) );
  AND2_X1 U337bar ( .A1(n632bar), .A2(n631bar), .ZN(n636bar) );
  OR2_X1 U338 ( .A1(in_72), .A2(in_70), .ZN(n631) );
  AND2_X1 U338bar ( .A1(in_72bar), .A2(in_70bar), .ZN(n631bar) );
  OR2_X1 U339 ( .A1(in_80), .A2(in_74), .ZN(n632) );
  AND2_X1 U339bar ( .A1(in_80bar), .A2(in_74bar), .ZN(n632bar) );
  OR2_X1 U340 ( .A1(n630), .A2(n629), .ZN(n942) );
  AND2_X1 U340bar ( .A1(n630bar), .A2(n629bar), .ZN(n942bar) );
  OR2_X1 U341 ( .A1(n628), .A2(n627), .ZN(n629) );
  AND2_X1 U341bar ( .A1(n628bar), .A2(n627bar), .ZN(n629bar) );
  OR2_X1 U342 ( .A1(n626), .A2(n625), .ZN(n627) );
  AND2_X1 U342bar ( .A1(n626bar), .A2(n625bar), .ZN(n627bar) );
  OR2_X1 U343 ( .A1(in[146]), .A2(in[100]), .ZN(n625) );
  AND2_X1 U343bar ( .A1(inbar[146]), .A2(inbar[100]), .ZN(n625bar) );
  OR2_X1 U344 ( .A1(in[168]), .A2(in[152]), .ZN(n626) );
  AND2_X1 U344bar ( .A1(inbar[168]), .A2(inbar[152]), .ZN(n626bar) );
  OR2_X1 U345 ( .A1(n624), .A2(n623), .ZN(n628) );
  AND2_X1 U345bar ( .A1(n624bar), .A2(n623bar), .ZN(n628bar) );
  OR2_X1 U346 ( .A1(in[199]), .A2(in[182]), .ZN(n623) );
  AND2_X1 U346bar ( .A1(inbar[199]), .A2(inbar[182]), .ZN(n623bar) );
  OR2_X1 U347 ( .A1(in[236]), .A2(in[204]), .ZN(n624) );
  AND2_X1 U347bar ( .A1(inbar[236]), .A2(inbar[204]), .ZN(n624bar) );
  OR2_X1 U348 ( .A1(n622), .A2(n621), .ZN(n630) );
  AND2_X1 U348bar ( .A1(n622bar), .A2(n621bar), .ZN(n630bar) );
  OR2_X1 U349 ( .A1(n620), .A2(n619), .ZN(n621) );
  AND2_X1 U349bar ( .A1(n620bar), .A2(n619bar), .ZN(n621bar) );
  OR2_X1 U350 ( .A1(in[89]), .A2(in[246]), .ZN(n619) );
  AND2_X1 U350bar ( .A1(inbar[89]), .A2(inbar[246]), .ZN(n619bar) );
  OR2_X1 U351 ( .A1(in[95]), .A2(in[92]), .ZN(n620) );
  AND2_X1 U351bar ( .A1(inbar[95]), .A2(inbar[92]), .ZN(n620bar) );
  OR2_X1 U352 ( .A1(n618), .A2(n617), .ZN(n622) );
  AND2_X1 U352bar ( .A1(n618bar), .A2(n617bar), .ZN(n622bar) );
  OR2_X1 U353 ( .A1(in_22), .A2(in_16), .ZN(n617) );
  AND2_X1 U353bar ( .A1(in_22bar), .A2(in_16bar), .ZN(n617bar) );
  OR2_X1 U354 ( .A1(in_51), .A2(in_49), .ZN(n618) );
  AND2_X1 U354bar ( .A1(in_51bar), .A2(in_49bar), .ZN(n618bar) );
  OR2_X1 U355 ( .A1(n616), .A2(n615), .ZN(n722) );
  AND2_X1 U355bar ( .A1(n616bar), .A2(n615bar), .ZN(n722bar) );
  OR2_X1 U356 ( .A1(in[158]), .A2(in[115]), .ZN(n615) );
  AND2_X1 U356bar ( .A1(inbar[158]), .A2(inbar[115]), .ZN(n615bar) );
  OR2_X1 U357 ( .A1(in[163]), .A2(n614), .ZN(n616) );
  AND2_X1 U357bar ( .A1(inbar[163]), .A2(n614bar), .ZN(n616bar) );
  OR2_X1 U358 ( .A1(in[206]), .A2(in[165]), .ZN(n614) );
  AND2_X1 U358bar ( .A1(inbar[206]), .A2(inbar[165]), .ZN(n614bar) );
  OR2_X1 U359 ( .A1(n613), .A2(n612), .ZN(n724) );
  AND2_X1 U359bar ( .A1(n613bar), .A2(n612bar), .ZN(n724bar) );
  OR2_X1 U360 ( .A1(n611), .A2(n610), .ZN(n612) );
  AND2_X1 U360bar ( .A1(n611bar), .A2(n610bar), .ZN(n612bar) );
  OR2_X1 U361 ( .A1(in[213]), .A2(in[207]), .ZN(n610) );
  AND2_X1 U361bar ( .A1(inbar[213]), .A2(inbar[207]), .ZN(n610bar) );
  OR2_X1 U362 ( .A1(in[215]), .A2(n609), .ZN(n611) );
  AND2_X1 U362bar ( .A1(inbar[215]), .A2(n609bar), .ZN(n611bar) );
  OR2_X1 U363 ( .A1(in[230]), .A2(in[220]), .ZN(n609) );
  AND2_X1 U363bar ( .A1(inbar[230]), .A2(inbar[220]), .ZN(n609bar) );
  OR2_X1 U364 ( .A1(n608), .A2(n607), .ZN(n613) );
  AND2_X1 U364bar ( .A1(n608bar), .A2(n607bar), .ZN(n613bar) );
  OR2_X1 U365 ( .A1(in[251]), .A2(in[234]), .ZN(n607) );
  AND2_X1 U365bar ( .A1(inbar[251]), .A2(inbar[234]), .ZN(n607bar) );
  OR2_X1 U366 ( .A1(in_17), .A2(n606), .ZN(n608) );
  AND2_X1 U366bar ( .A1(in_17bar), .A2(n606bar), .ZN(n608bar) );
  OR2_X1 U367 ( .A1(in_65), .A2(in_56), .ZN(n606) );
  AND2_X1 U367bar ( .A1(in_65bar), .A2(in_56bar), .ZN(n606bar) );
  OR2_X1 U368 ( .A1(n605), .A2(n604), .ZN(out[0]) );
  AND2_X1 U368bar ( .A1(n605bar), .A2(n604bar), .ZN(outbar[0]) );
  OR2_X1 U369 ( .A1(n603), .A2(n602), .ZN(n604) );
  AND2_X1 U369bar ( .A1(n603bar), .A2(n602bar), .ZN(n604bar) );
  OR2_X1 U370 ( .A1(n601), .A2(n600), .ZN(n602) );
  AND2_X1 U370bar ( .A1(n601bar), .A2(n600bar), .ZN(n602bar) );
  OR2_X1 U371 ( .A1(n820), .A2(n785), .ZN(n600) );
  AND2_X1 U371bar ( .A1(n820bar), .A2(n785bar), .ZN(n600bar) );
  OR2_X1 U372 ( .A1(n599), .A2(n598), .ZN(n785) );
  AND2_X1 U372bar ( .A1(n599bar), .A2(n598bar), .ZN(n785bar) );
  OR2_X1 U373 ( .A1(n597), .A2(n596), .ZN(n598) );
  AND2_X1 U373bar ( .A1(n597bar), .A2(n596bar), .ZN(n598bar) );
  OR2_X1 U374 ( .A1(n595), .A2(n594), .ZN(n596) );
  AND2_X1 U374bar ( .A1(n595bar), .A2(n594bar), .ZN(n596bar) );
  OR2_X1 U375 ( .A1(in[135]), .A2(in[104]), .ZN(n594) );
  AND2_X1 U375bar ( .A1(inbar[135]), .A2(inbar[104]), .ZN(n594bar) );
  OR2_X1 U376 ( .A1(in[188]), .A2(in[178]), .ZN(n595) );
  AND2_X1 U376bar ( .A1(inbar[188]), .A2(inbar[178]), .ZN(n595bar) );
  OR2_X1 U377 ( .A1(n593), .A2(n592), .ZN(n597) );
  AND2_X1 U377bar ( .A1(n593bar), .A2(n592bar), .ZN(n597bar) );
  OR2_X1 U378 ( .A1(in[217]), .A2(in[194]), .ZN(n592) );
  AND2_X1 U378bar ( .A1(inbar[217]), .A2(inbar[194]), .ZN(n592bar) );
  OR2_X1 U379 ( .A1(in[237]), .A2(in[218]), .ZN(n593) );
  AND2_X1 U379bar ( .A1(inbar[237]), .A2(inbar[218]), .ZN(n593bar) );
  OR2_X1 U380 ( .A1(n591), .A2(n590), .ZN(n599) );
  AND2_X1 U380bar ( .A1(n591bar), .A2(n590bar), .ZN(n599bar) );
  OR2_X1 U381 ( .A1(n589), .A2(n588), .ZN(n590) );
  AND2_X1 U381bar ( .A1(n589bar), .A2(n588bar), .ZN(n590bar) );
  OR2_X1 U382 ( .A1(in_2), .A2(in_10), .ZN(n588) );
  AND2_X1 U382bar ( .A1(in_2bar), .A2(in_10bar), .ZN(n588bar) );
  OR2_X1 U383 ( .A1(in_47), .A2(in_22), .ZN(n589) );
  AND2_X1 U383bar ( .A1(in_47bar), .A2(in_22bar), .ZN(n589bar) );
  OR2_X1 U384 ( .A1(n587), .A2(n586), .ZN(n591) );
  AND2_X1 U384bar ( .A1(n587bar), .A2(n586bar), .ZN(n591bar) );
  OR2_X1 U385 ( .A1(in_56), .A2(in_54), .ZN(n586) );
  AND2_X1 U385bar ( .A1(in_56bar), .A2(in_54bar), .ZN(n586bar) );
  OR2_X1 U386 ( .A1(in_63), .A2(in_61), .ZN(n587) );
  AND2_X1 U386bar ( .A1(in_63bar), .A2(in_61bar), .ZN(n587bar) );
  OR2_X1 U387 ( .A1(n585), .A2(n584), .ZN(n820) );
  AND2_X1 U387bar ( .A1(n585bar), .A2(n584bar), .ZN(n820bar) );
  OR2_X1 U388 ( .A1(n583), .A2(n582), .ZN(n584) );
  AND2_X1 U388bar ( .A1(n583bar), .A2(n582bar), .ZN(n584bar) );
  OR2_X1 U389 ( .A1(n581), .A2(n580), .ZN(n582) );
  AND2_X1 U389bar ( .A1(n581bar), .A2(n580bar), .ZN(n582bar) );
  OR2_X1 U390 ( .A1(in[158]), .A2(in[142]), .ZN(n580) );
  AND2_X1 U390bar ( .A1(inbar[158]), .A2(inbar[142]), .ZN(n580bar) );
  OR2_X1 U391 ( .A1(in[175]), .A2(in[164]), .ZN(n581) );
  AND2_X1 U391bar ( .A1(inbar[175]), .A2(inbar[164]), .ZN(n581bar) );
  OR2_X1 U392 ( .A1(n579), .A2(n578), .ZN(n583) );
  AND2_X1 U392bar ( .A1(n579bar), .A2(n578bar), .ZN(n583bar) );
  OR2_X1 U393 ( .A1(in[228]), .A2(in[204]), .ZN(n578) );
  AND2_X1 U393bar ( .A1(inbar[228]), .A2(inbar[204]), .ZN(n578bar) );
  OR2_X1 U394 ( .A1(in[91]), .A2(in[87]), .ZN(n579) );
  AND2_X1 U394bar ( .A1(inbar[91]), .A2(inbar[87]), .ZN(n579bar) );
  OR2_X1 U395 ( .A1(n577), .A2(n576), .ZN(n585) );
  AND2_X1 U395bar ( .A1(n577bar), .A2(n576bar), .ZN(n585bar) );
  OR2_X1 U396 ( .A1(n575), .A2(n574), .ZN(n576) );
  AND2_X1 U396bar ( .A1(n575bar), .A2(n574bar), .ZN(n576bar) );
  OR2_X1 U397 ( .A1(in_21), .A2(in_11), .ZN(n574) );
  AND2_X1 U397bar ( .A1(in_21bar), .A2(in_11bar), .ZN(n574bar) );
  OR2_X1 U398 ( .A1(in_5), .A2(in_3), .ZN(n575) );
  AND2_X1 U398bar ( .A1(in_5bar), .A2(in_3bar), .ZN(n575bar) );
  OR2_X1 U399 ( .A1(n573), .A2(n572), .ZN(n577) );
  AND2_X1 U399bar ( .A1(n573bar), .A2(n572bar), .ZN(n577bar) );
  OR2_X1 U400 ( .A1(in_68), .A2(in_64), .ZN(n572) );
  AND2_X1 U400bar ( .A1(in_68bar), .A2(in_64bar), .ZN(n572bar) );
  OR2_X1 U401 ( .A1(in_76), .A2(in_73), .ZN(n573) );
  AND2_X1 U401bar ( .A1(in_76bar), .A2(in_73bar), .ZN(n573bar) );
  OR2_X1 U402 ( .A1(n778), .A2(n571), .ZN(n601) );
  AND2_X1 U402bar ( .A1(n778bar), .A2(n571bar), .ZN(n601bar) );
  OR2_X1 U403 ( .A1(in[100]), .A2(n965), .ZN(n571) );
  AND2_X1 U403bar ( .A1(inbar[100]), .A2(n965bar), .ZN(n571bar) );
  OR2_X1 U404 ( .A1(n570), .A2(n569), .ZN(n965) );
  AND2_X1 U404bar ( .A1(n570bar), .A2(n569bar), .ZN(n965bar) );
  OR2_X1 U405 ( .A1(n568), .A2(n567), .ZN(n569) );
  AND2_X1 U405bar ( .A1(n568bar), .A2(n567bar), .ZN(n569bar) );
  OR2_X1 U406 ( .A1(n566), .A2(n565), .ZN(n567) );
  AND2_X1 U406bar ( .A1(n566bar), .A2(n565bar), .ZN(n567bar) );
  OR2_X1 U407 ( .A1(n817), .A2(n750), .ZN(n565) );
  AND2_X1 U407bar ( .A1(n817bar), .A2(n750bar), .ZN(n565bar) );
  OR2_X1 U408 ( .A1(n564), .A2(n563), .ZN(n750) );
  AND2_X1 U408bar ( .A1(n564bar), .A2(n563bar), .ZN(n750bar) );
  OR2_X1 U409 ( .A1(n562), .A2(n561), .ZN(n563) );
  AND2_X1 U409bar ( .A1(n562bar), .A2(n561bar), .ZN(n563bar) );
  OR2_X1 U410 ( .A1(n560), .A2(n559), .ZN(n561) );
  AND2_X1 U410bar ( .A1(n560bar), .A2(n559bar), .ZN(n561bar) );
  OR2_X1 U411 ( .A1(in[119]), .A2(in[103]), .ZN(n559) );
  AND2_X1 U411bar ( .A1(inbar[119]), .A2(inbar[103]), .ZN(n559bar) );
  OR2_X1 U412 ( .A1(in[137]), .A2(in[133]), .ZN(n560) );
  AND2_X1 U412bar ( .A1(inbar[137]), .A2(inbar[133]), .ZN(n560bar) );
  OR2_X1 U413 ( .A1(n558), .A2(n557), .ZN(n562) );
  AND2_X1 U413bar ( .A1(n558bar), .A2(n557bar), .ZN(n562bar) );
  OR2_X1 U414 ( .A1(in[176]), .A2(in[173]), .ZN(n557) );
  AND2_X1 U414bar ( .A1(inbar[176]), .A2(inbar[173]), .ZN(n557bar) );
  OR2_X1 U415 ( .A1(in[210]), .A2(in[181]), .ZN(n558) );
  AND2_X1 U415bar ( .A1(inbar[210]), .A2(inbar[181]), .ZN(n558bar) );
  OR2_X1 U416 ( .A1(n556), .A2(n555), .ZN(n564) );
  AND2_X1 U416bar ( .A1(n556bar), .A2(n555bar), .ZN(n564bar) );
  OR2_X1 U417 ( .A1(n554), .A2(n553), .ZN(n555) );
  AND2_X1 U417bar ( .A1(n554bar), .A2(n553bar), .ZN(n555bar) );
  OR2_X1 U418 ( .A1(in_13), .A2(in[234]), .ZN(n553) );
  AND2_X1 U418bar ( .A1(in_13bar), .A2(inbar[234]), .ZN(n553bar) );
  OR2_X1 U419 ( .A1(in_38), .A2(in_32), .ZN(n554) );
  AND2_X1 U419bar ( .A1(in_38bar), .A2(in_32bar), .ZN(n554bar) );
  OR2_X1 U420 ( .A1(n552), .A2(n551), .ZN(n556) );
  AND2_X1 U420bar ( .A1(n552bar), .A2(n551bar), .ZN(n556bar) );
  OR2_X1 U421 ( .A1(in_42), .A2(in_41), .ZN(n551) );
  AND2_X1 U421bar ( .A1(in_42bar), .A2(in_41bar), .ZN(n551bar) );
  OR2_X1 U422 ( .A1(in_7), .A2(in_49), .ZN(n552) );
  AND2_X1 U422bar ( .A1(in_7bar), .A2(in_49bar), .ZN(n552bar) );
  OR2_X1 U423 ( .A1(n550), .A2(n549), .ZN(n817) );
  AND2_X1 U423bar ( .A1(n550bar), .A2(n549bar), .ZN(n817bar) );
  OR2_X1 U424 ( .A1(n548), .A2(n547), .ZN(n549) );
  AND2_X1 U424bar ( .A1(n548bar), .A2(n547bar), .ZN(n549bar) );
  OR2_X1 U425 ( .A1(n546), .A2(n545), .ZN(n547) );
  AND2_X1 U425bar ( .A1(n546bar), .A2(n545bar), .ZN(n547bar) );
  OR2_X1 U426 ( .A1(in[159]), .A2(in[105]), .ZN(n545) );
  AND2_X1 U426bar ( .A1(inbar[159]), .A2(inbar[105]), .ZN(n545bar) );
  OR2_X1 U427 ( .A1(in[206]), .A2(in[183]), .ZN(n546) );
  AND2_X1 U427bar ( .A1(inbar[206]), .A2(inbar[183]), .ZN(n546bar) );
  OR2_X1 U428 ( .A1(n544), .A2(n543), .ZN(n548) );
  AND2_X1 U428bar ( .A1(n544bar), .A2(n543bar), .ZN(n548bar) );
  OR2_X1 U429 ( .A1(in[229]), .A2(in[219]), .ZN(n543) );
  AND2_X1 U429bar ( .A1(inbar[229]), .A2(inbar[219]), .ZN(n543bar) );
  OR2_X1 U430 ( .A1(in[235]), .A2(in[232]), .ZN(n544) );
  AND2_X1 U430bar ( .A1(inbar[235]), .A2(inbar[232]), .ZN(n544bar) );
  OR2_X1 U431 ( .A1(n542), .A2(n541), .ZN(n550) );
  AND2_X1 U431bar ( .A1(n542bar), .A2(n541bar), .ZN(n550bar) );
  OR2_X1 U432 ( .A1(n540), .A2(n539), .ZN(n541) );
  AND2_X1 U432bar ( .A1(n540bar), .A2(n539bar), .ZN(n541bar) );
  OR2_X1 U433 ( .A1(in[249]), .A2(in[242]), .ZN(n539) );
  AND2_X1 U433bar ( .A1(inbar[249]), .A2(inbar[242]), .ZN(n539bar) );
  OR2_X1 U434 ( .A1(in[89]), .A2(in[254]), .ZN(n540) );
  AND2_X1 U434bar ( .A1(inbar[89]), .A2(inbar[254]), .ZN(n540bar) );
  OR2_X1 U435 ( .A1(n538), .A2(n537), .ZN(n542) );
  AND2_X1 U435bar ( .A1(n538bar), .A2(n537bar), .ZN(n542bar) );
  OR2_X1 U436 ( .A1(in_14), .A2(in[99]), .ZN(n537) );
  AND2_X1 U436bar ( .A1(in_14bar), .A2(inbar[99]), .ZN(n537bar) );
  OR2_X1 U437 ( .A1(in_60), .A2(in_18), .ZN(n538) );
  AND2_X1 U437bar ( .A1(in_60bar), .A2(in_18bar), .ZN(n538bar) );
  OR2_X1 U438 ( .A1(in[113]), .A2(n763), .ZN(n566) );
  AND2_X1 U438bar ( .A1(inbar[113]), .A2(n763bar), .ZN(n566bar) );
  OR2_X1 U439 ( .A1(n536), .A2(n535), .ZN(n763) );
  AND2_X1 U439bar ( .A1(n536bar), .A2(n535bar), .ZN(n763bar) );
  OR2_X1 U440 ( .A1(n534), .A2(n533), .ZN(n535) );
  AND2_X1 U440bar ( .A1(n534bar), .A2(n533bar), .ZN(n535bar) );
  OR2_X1 U441 ( .A1(n532), .A2(n531), .ZN(n533) );
  AND2_X1 U441bar ( .A1(n532bar), .A2(n531bar), .ZN(n533bar) );
  OR2_X1 U442 ( .A1(in[115]), .A2(in[110]), .ZN(n531) );
  AND2_X1 U442bar ( .A1(inbar[115]), .A2(inbar[110]), .ZN(n531bar) );
  OR2_X1 U443 ( .A1(in[125]), .A2(in[117]), .ZN(n532) );
  AND2_X1 U443bar ( .A1(inbar[125]), .A2(inbar[117]), .ZN(n532bar) );
  OR2_X1 U444 ( .A1(n530), .A2(n529), .ZN(n534) );
  AND2_X1 U444bar ( .A1(n530bar), .A2(n529bar), .ZN(n534bar) );
  OR2_X1 U445 ( .A1(in[180]), .A2(in[128]), .ZN(n529) );
  AND2_X1 U445bar ( .A1(inbar[180]), .A2(inbar[128]), .ZN(n529bar) );
  OR2_X1 U446 ( .A1(in[205]), .A2(in[201]), .ZN(n530) );
  AND2_X1 U446bar ( .A1(inbar[205]), .A2(inbar[201]), .ZN(n530bar) );
  OR2_X1 U447 ( .A1(n528), .A2(n527), .ZN(n536) );
  AND2_X1 U447bar ( .A1(n528bar), .A2(n527bar), .ZN(n536bar) );
  OR2_X1 U448 ( .A1(n526), .A2(n525), .ZN(n527) );
  AND2_X1 U448bar ( .A1(n526bar), .A2(n525bar), .ZN(n527bar) );
  OR2_X1 U449 ( .A1(in[244]), .A2(in[239]), .ZN(n525) );
  AND2_X1 U449bar ( .A1(inbar[244]), .A2(inbar[239]), .ZN(n525bar) );
  OR2_X1 U450 ( .A1(in[95]), .A2(in[83]), .ZN(n526) );
  AND2_X1 U450bar ( .A1(inbar[95]), .A2(inbar[83]), .ZN(n526bar) );
  OR2_X1 U451 ( .A1(n524), .A2(n523), .ZN(n528) );
  AND2_X1 U451bar ( .A1(n524bar), .A2(n523bar), .ZN(n528bar) );
  OR2_X1 U452 ( .A1(in_24), .A2(in[97]), .ZN(n523) );
  AND2_X1 U452bar ( .A1(in_24bar), .A2(inbar[97]), .ZN(n523bar) );
  OR2_X1 U453 ( .A1(in_33), .A2(in_27), .ZN(n524) );
  AND2_X1 U453bar ( .A1(in_33bar), .A2(in_27bar), .ZN(n524bar) );
  OR2_X1 U454 ( .A1(n522), .A2(n521), .ZN(n568) );
  AND2_X1 U454bar ( .A1(n522bar), .A2(n521bar), .ZN(n568bar) );
  OR2_X1 U455 ( .A1(in[145]), .A2(in[126]), .ZN(n521) );
  AND2_X1 U455bar ( .A1(inbar[145]), .A2(inbar[126]), .ZN(n521bar) );
  OR2_X1 U456 ( .A1(in[169]), .A2(n520), .ZN(n522) );
  AND2_X1 U456bar ( .A1(inbar[169]), .A2(n520bar), .ZN(n522bar) );
  OR2_X1 U457 ( .A1(in[221]), .A2(in[172]), .ZN(n520) );
  AND2_X1 U457bar ( .A1(inbar[221]), .A2(inbar[172]), .ZN(n520bar) );
  OR2_X1 U458 ( .A1(n519), .A2(n518), .ZN(n570) );
  AND2_X1 U458bar ( .A1(n519bar), .A2(n518bar), .ZN(n570bar) );
  OR2_X1 U459 ( .A1(n517), .A2(n516), .ZN(n518) );
  AND2_X1 U459bar ( .A1(n517bar), .A2(n516bar), .ZN(n518bar) );
  OR2_X1 U460 ( .A1(in[241]), .A2(in[224]), .ZN(n516) );
  AND2_X1 U460bar ( .A1(inbar[241]), .A2(inbar[224]), .ZN(n516bar) );
  OR2_X1 U461 ( .A1(in[86]), .A2(n515), .ZN(n517) );
  AND2_X1 U461bar ( .A1(inbar[86]), .A2(n515bar), .ZN(n517bar) );
  OR2_X1 U462 ( .A1(in_43), .A2(in_34), .ZN(n515) );
  AND2_X1 U462bar ( .A1(in_43bar), .A2(in_34bar), .ZN(n515bar) );
  OR2_X1 U463 ( .A1(n514), .A2(n513), .ZN(n519) );
  AND2_X1 U463bar ( .A1(n514bar), .A2(n513bar), .ZN(n519bar) );
  OR2_X1 U464 ( .A1(in_65), .A2(in_51), .ZN(n513) );
  AND2_X1 U464bar ( .A1(in_65bar), .A2(in_51bar), .ZN(n513bar) );
  OR2_X1 U465 ( .A1(in_75), .A2(n512), .ZN(n514) );
  AND2_X1 U465bar ( .A1(in_75bar), .A2(n512bar), .ZN(n514bar) );
  OR2_X1 U466 ( .A1(in_81), .A2(in_77), .ZN(n512) );
  AND2_X1 U466bar ( .A1(in_81bar), .A2(in_77bar), .ZN(n512bar) );
  OR2_X1 U467 ( .A1(n511), .A2(n510), .ZN(n778) );
  AND2_X1 U467bar ( .A1(n511bar), .A2(n510bar), .ZN(n778bar) );
  OR2_X1 U468 ( .A1(n509), .A2(n508), .ZN(n510) );
  AND2_X1 U468bar ( .A1(n509bar), .A2(n508bar), .ZN(n510bar) );
  OR2_X1 U469 ( .A1(n507), .A2(n506), .ZN(n508) );
  AND2_X1 U469bar ( .A1(n507bar), .A2(n506bar), .ZN(n508bar) );
  OR2_X1 U470 ( .A1(in[107]), .A2(in[101]), .ZN(n506) );
  AND2_X1 U470bar ( .A1(inbar[107]), .A2(inbar[101]), .ZN(n506bar) );
  OR2_X1 U471 ( .A1(in[139]), .A2(in[132]), .ZN(n507) );
  AND2_X1 U471bar ( .A1(inbar[139]), .A2(inbar[132]), .ZN(n507bar) );
  OR2_X1 U472 ( .A1(n505), .A2(n504), .ZN(n509) );
  AND2_X1 U472bar ( .A1(n505bar), .A2(n504bar), .ZN(n509bar) );
  OR2_X1 U473 ( .A1(in[146]), .A2(in[141]), .ZN(n504) );
  AND2_X1 U473bar ( .A1(inbar[146]), .A2(inbar[141]), .ZN(n504bar) );
  OR2_X1 U474 ( .A1(in[203]), .A2(in[179]), .ZN(n505) );
  AND2_X1 U474bar ( .A1(inbar[203]), .A2(inbar[179]), .ZN(n505bar) );
  OR2_X1 U475 ( .A1(n503), .A2(n502), .ZN(n511) );
  AND2_X1 U475bar ( .A1(n503bar), .A2(n502bar), .ZN(n511bar) );
  OR2_X1 U476 ( .A1(n501), .A2(n500), .ZN(n502) );
  AND2_X1 U476bar ( .A1(n501bar), .A2(n500bar), .ZN(n502bar) );
  OR2_X1 U477 ( .A1(in[243]), .A2(in[222]), .ZN(n500) );
  AND2_X1 U477bar ( .A1(inbar[243]), .A2(inbar[222]), .ZN(n500bar) );
  OR2_X1 U478 ( .A1(in[251]), .A2(in[250]), .ZN(n501) );
  AND2_X1 U478bar ( .A1(inbar[251]), .A2(inbar[250]), .ZN(n501bar) );
  OR2_X1 U479 ( .A1(n499), .A2(n498), .ZN(n503) );
  AND2_X1 U479bar ( .A1(n499bar), .A2(n498bar), .ZN(n503bar) );
  OR2_X1 U480 ( .A1(in_37), .A2(in_19), .ZN(n498) );
  AND2_X1 U480bar ( .A1(in_37bar), .A2(in_19bar), .ZN(n498bar) );
  OR2_X1 U481 ( .A1(in_78), .A2(in_6), .ZN(n499) );
  AND2_X1 U481bar ( .A1(in_78bar), .A2(in_6bar), .ZN(n499bar) );
  OR2_X1 U482 ( .A1(n497), .A2(n496), .ZN(n603) );
  AND2_X1 U482bar ( .A1(n497bar), .A2(n496bar), .ZN(n603bar) );
  OR2_X1 U483 ( .A1(in[112]), .A2(in[102]), .ZN(n496) );
  AND2_X1 U483bar ( .A1(inbar[112]), .A2(inbar[102]), .ZN(n496bar) );
  OR2_X1 U484 ( .A1(in[123]), .A2(n495), .ZN(n497) );
  AND2_X1 U484bar ( .A1(inbar[123]), .A2(n495bar), .ZN(n497bar) );
  OR2_X1 U485 ( .A1(in[143]), .A2(in[130]), .ZN(n495) );
  AND2_X1 U485bar ( .A1(inbar[143]), .A2(inbar[130]), .ZN(n495bar) );
  OR2_X1 U486 ( .A1(n494), .A2(n493), .ZN(n605) );
  AND2_X1 U486bar ( .A1(n494bar), .A2(n493bar), .ZN(n605bar) );
  OR2_X1 U487 ( .A1(n492), .A2(n491), .ZN(n493) );
  AND2_X1 U487bar ( .A1(n492bar), .A2(n491bar), .ZN(n493bar) );
  OR2_X1 U488 ( .A1(in[216]), .A2(in[213]), .ZN(n491) );
  AND2_X1 U488bar ( .A1(inbar[216]), .A2(inbar[213]), .ZN(n491bar) );
  OR2_X1 U489 ( .A1(in[227]), .A2(n490), .ZN(n492) );
  AND2_X1 U489bar ( .A1(inbar[227]), .A2(n490bar), .ZN(n492bar) );
  OR2_X1 U490 ( .A1(in_0), .A2(in[248]), .ZN(n490) );
  AND2_X1 U490bar ( .A1(in_0bar), .A2(inbar[248]), .ZN(n490bar) );
  OR2_X1 U491 ( .A1(n489), .A2(n488), .ZN(n494) );
  AND2_X1 U491bar ( .A1(n489bar), .A2(n488bar), .ZN(n494bar) );
  OR2_X1 U492 ( .A1(in_46), .A2(in_44), .ZN(n488) );
  AND2_X1 U492bar ( .A1(in_46bar), .A2(in_44bar), .ZN(n488bar) );
  OR2_X1 U493 ( .A1(in_50), .A2(n487), .ZN(n489) );
  AND2_X1 U493bar ( .A1(in_50bar), .A2(n487bar), .ZN(n489bar) );
  OR2_X1 U494 ( .A1(in_9), .A2(in_80), .ZN(n487) );
  AND2_X1 U494bar ( .A1(in_9bar), .A2(in_80bar), .ZN(n487bar) );
endmodule

module sBox_2 ( in, inbar, out, outbar );

  input wire [7:0] in;
  input wire [7:0] inbar;
//input_done

  output wire [7:0] out;
  output wire [7:0] outbar;
//output_done

  wire [255:0] decodeOut;
  wire [255:0] decodeOutbar;
//wire_done

  decode_2 dec ( .in(in), .inbar(inbar), .out(decodeOut), .outbar(decodeOutbar) );
  encode_2 enc ( .in(decodeOut), .inbar(decodeOutbar), .out(out), .outbar(outbar) );
endmodule

module CD2_9 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD2_10 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD2_11 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD2_12 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD4_5 ( a, abar, b, bbar, y, ybar );

  input wire [3:0] a;
  input wire [3:0] b;
  input wire [3:0] abar;
  input wire [3:0] bbar;
//input_done

  output wire [15:0] y;
  output wire [15:0] ybar;
//output_done

//wire_done

  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]) );
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]) );
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]) );
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]) );
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]) );
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]) );
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]) );
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]) );
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]) );
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]) );
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]) );
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]) );
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]) );
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]) );
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]) );
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]) );
endmodule

module CD4_6 ( a, abar, b, bbar, y, ybar );

  input wire [3:0] a;
  input wire [3:0] b;
  input wire [3:0] abar;
  input wire [3:0] bbar;
//input_done

  output wire [15:0] y;
  output wire [15:0] ybar;
//output_done

//wire_done

  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]) );
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]) );
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]) );
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]) );
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]) );
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]) );
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]) );
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]) );
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]) );
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]) );
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]) );
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]) );
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]) );
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]) );
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]) );
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]) );
endmodule

module CD16_3 ( a, abar, b, bbar, y, ybar );

  input wire [15:0] a;
  input wire [15:0] b;
  input wire [15:0] abar;
  input wire [15:0] bbar;
//input_done

  output wire [255:0] y;
  output wire [255:0] ybar;
//output_done

//wire_done

  AND2_X1 U1 ( .A1(b[9]), .A2(a[0]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[9]), .A2(abar[0]), .ZN(ybar[9]) );
  AND2_X1 U2 ( .A1(b[3]), .A2(a[6]), .ZN(y[99]) );
  OR2_X1 U2bar ( .A1(bbar[3]), .A2(abar[6]), .ZN(ybar[99]) );
  AND2_X1 U3 ( .A1(b[2]), .A2(a[6]), .ZN(y[98]) );
  OR2_X1 U3bar ( .A1(bbar[2]), .A2(abar[6]), .ZN(ybar[98]) );
  AND2_X1 U4 ( .A1(b[1]), .A2(a[6]), .ZN(y[97]) );
  OR2_X1 U4bar ( .A1(bbar[1]), .A2(abar[6]), .ZN(ybar[97]) );
  AND2_X1 U5 ( .A1(b[0]), .A2(a[6]), .ZN(y[96]) );
  OR2_X1 U5bar ( .A1(bbar[0]), .A2(abar[6]), .ZN(ybar[96]) );
  AND2_X1 U6 ( .A1(b[15]), .A2(a[5]), .ZN(y[95]) );
  OR2_X1 U6bar ( .A1(bbar[15]), .A2(abar[5]), .ZN(ybar[95]) );
  AND2_X1 U7 ( .A1(b[14]), .A2(a[5]), .ZN(y[94]) );
  OR2_X1 U7bar ( .A1(bbar[14]), .A2(abar[5]), .ZN(ybar[94]) );
  AND2_X1 U8 ( .A1(b[13]), .A2(a[5]), .ZN(y[93]) );
  OR2_X1 U8bar ( .A1(bbar[13]), .A2(abar[5]), .ZN(ybar[93]) );
  AND2_X1 U9 ( .A1(b[12]), .A2(a[5]), .ZN(y[92]) );
  OR2_X1 U9bar ( .A1(bbar[12]), .A2(abar[5]), .ZN(ybar[92]) );
  AND2_X1 U10 ( .A1(b[11]), .A2(a[5]), .ZN(y[91]) );
  OR2_X1 U10bar ( .A1(bbar[11]), .A2(abar[5]), .ZN(ybar[91]) );
  AND2_X1 U11 ( .A1(b[10]), .A2(a[5]), .ZN(y[90]) );
  OR2_X1 U11bar ( .A1(bbar[10]), .A2(abar[5]), .ZN(ybar[90]) );
  AND2_X1 U12 ( .A1(b[8]), .A2(a[0]), .ZN(y[8]) );
  OR2_X1 U12bar ( .A1(bbar[8]), .A2(abar[0]), .ZN(ybar[8]) );
  AND2_X1 U13 ( .A1(a[5]), .A2(b[9]), .ZN(y[89]) );
  OR2_X1 U13bar ( .A1(abar[5]), .A2(bbar[9]), .ZN(ybar[89]) );
  AND2_X1 U14 ( .A1(b[8]), .A2(a[5]), .ZN(y[88]) );
  OR2_X1 U14bar ( .A1(bbar[8]), .A2(abar[5]), .ZN(ybar[88]) );
  AND2_X1 U15 ( .A1(b[7]), .A2(a[5]), .ZN(y[87]) );
  OR2_X1 U15bar ( .A1(bbar[7]), .A2(abar[5]), .ZN(ybar[87]) );
  AND2_X1 U16 ( .A1(b[6]), .A2(a[5]), .ZN(y[86]) );
  OR2_X1 U16bar ( .A1(bbar[6]), .A2(abar[5]), .ZN(ybar[86]) );
  AND2_X1 U17 ( .A1(b[5]), .A2(a[5]), .ZN(y[85]) );
  OR2_X1 U17bar ( .A1(bbar[5]), .A2(abar[5]), .ZN(ybar[85]) );
  AND2_X1 U18 ( .A1(b[4]), .A2(a[5]), .ZN(y[84]) );
  OR2_X1 U18bar ( .A1(bbar[4]), .A2(abar[5]), .ZN(ybar[84]) );
  AND2_X1 U19 ( .A1(a[5]), .A2(b[3]), .ZN(y[83]) );
  OR2_X1 U19bar ( .A1(abar[5]), .A2(bbar[3]), .ZN(ybar[83]) );
  AND2_X1 U20 ( .A1(a[5]), .A2(b[2]), .ZN(y[82]) );
  OR2_X1 U20bar ( .A1(abar[5]), .A2(bbar[2]), .ZN(ybar[82]) );
  AND2_X1 U21 ( .A1(a[5]), .A2(b[1]), .ZN(y[81]) );
  OR2_X1 U21bar ( .A1(abar[5]), .A2(bbar[1]), .ZN(ybar[81]) );
  AND2_X1 U22 ( .A1(a[5]), .A2(b[0]), .ZN(y[80]) );
  OR2_X1 U22bar ( .A1(abar[5]), .A2(bbar[0]), .ZN(ybar[80]) );
  AND2_X1 U23 ( .A1(b[7]), .A2(a[0]), .ZN(y[7]) );
  OR2_X1 U23bar ( .A1(bbar[7]), .A2(abar[0]), .ZN(ybar[7]) );
  AND2_X1 U24 ( .A1(a[4]), .A2(b[15]), .ZN(y[79]) );
  OR2_X1 U24bar ( .A1(abar[4]), .A2(bbar[15]), .ZN(ybar[79]) );
  AND2_X1 U25 ( .A1(a[4]), .A2(b[14]), .ZN(y[78]) );
  OR2_X1 U25bar ( .A1(abar[4]), .A2(bbar[14]), .ZN(ybar[78]) );
  AND2_X1 U26 ( .A1(a[4]), .A2(b[13]), .ZN(y[77]) );
  OR2_X1 U26bar ( .A1(abar[4]), .A2(bbar[13]), .ZN(ybar[77]) );
  AND2_X1 U27 ( .A1(a[4]), .A2(b[12]), .ZN(y[76]) );
  OR2_X1 U27bar ( .A1(abar[4]), .A2(bbar[12]), .ZN(ybar[76]) );
  AND2_X1 U28 ( .A1(a[4]), .A2(b[11]), .ZN(y[75]) );
  OR2_X1 U28bar ( .A1(abar[4]), .A2(bbar[11]), .ZN(ybar[75]) );
  AND2_X1 U29 ( .A1(a[4]), .A2(b[10]), .ZN(y[74]) );
  OR2_X1 U29bar ( .A1(abar[4]), .A2(bbar[10]), .ZN(ybar[74]) );
  AND2_X1 U30 ( .A1(a[4]), .A2(b[9]), .ZN(y[73]) );
  OR2_X1 U30bar ( .A1(abar[4]), .A2(bbar[9]), .ZN(ybar[73]) );
  AND2_X1 U31 ( .A1(a[4]), .A2(b[8]), .ZN(y[72]) );
  OR2_X1 U31bar ( .A1(abar[4]), .A2(bbar[8]), .ZN(ybar[72]) );
  AND2_X1 U32 ( .A1(a[4]), .A2(b[7]), .ZN(y[71]) );
  OR2_X1 U32bar ( .A1(abar[4]), .A2(bbar[7]), .ZN(ybar[71]) );
  AND2_X1 U33 ( .A1(a[4]), .A2(b[6]), .ZN(y[70]) );
  OR2_X1 U33bar ( .A1(abar[4]), .A2(bbar[6]), .ZN(ybar[70]) );
  AND2_X1 U34 ( .A1(b[6]), .A2(a[0]), .ZN(y[6]) );
  OR2_X1 U34bar ( .A1(bbar[6]), .A2(abar[0]), .ZN(ybar[6]) );
  AND2_X1 U35 ( .A1(a[4]), .A2(b[5]), .ZN(y[69]) );
  OR2_X1 U35bar ( .A1(abar[4]), .A2(bbar[5]), .ZN(ybar[69]) );
  AND2_X1 U36 ( .A1(a[4]), .A2(b[4]), .ZN(y[68]) );
  OR2_X1 U36bar ( .A1(abar[4]), .A2(bbar[4]), .ZN(ybar[68]) );
  AND2_X1 U37 ( .A1(a[4]), .A2(b[3]), .ZN(y[67]) );
  OR2_X1 U37bar ( .A1(abar[4]), .A2(bbar[3]), .ZN(ybar[67]) );
  AND2_X1 U38 ( .A1(a[4]), .A2(b[2]), .ZN(y[66]) );
  OR2_X1 U38bar ( .A1(abar[4]), .A2(bbar[2]), .ZN(ybar[66]) );
  AND2_X1 U39 ( .A1(a[4]), .A2(b[1]), .ZN(y[65]) );
  OR2_X1 U39bar ( .A1(abar[4]), .A2(bbar[1]), .ZN(ybar[65]) );
  AND2_X1 U40 ( .A1(a[4]), .A2(b[0]), .ZN(y[64]) );
  OR2_X1 U40bar ( .A1(abar[4]), .A2(bbar[0]), .ZN(ybar[64]) );
  AND2_X1 U41 ( .A1(a[3]), .A2(b[15]), .ZN(y[63]) );
  OR2_X1 U41bar ( .A1(abar[3]), .A2(bbar[15]), .ZN(ybar[63]) );
  AND2_X1 U42 ( .A1(a[3]), .A2(b[14]), .ZN(y[62]) );
  OR2_X1 U42bar ( .A1(abar[3]), .A2(bbar[14]), .ZN(ybar[62]) );
  AND2_X1 U43 ( .A1(a[3]), .A2(b[13]), .ZN(y[61]) );
  OR2_X1 U43bar ( .A1(abar[3]), .A2(bbar[13]), .ZN(ybar[61]) );
  AND2_X1 U44 ( .A1(a[3]), .A2(b[12]), .ZN(y[60]) );
  OR2_X1 U44bar ( .A1(abar[3]), .A2(bbar[12]), .ZN(ybar[60]) );
  AND2_X1 U45 ( .A1(b[5]), .A2(a[0]), .ZN(y[5]) );
  OR2_X1 U45bar ( .A1(bbar[5]), .A2(abar[0]), .ZN(ybar[5]) );
  AND2_X1 U46 ( .A1(a[3]), .A2(b[11]), .ZN(y[59]) );
  OR2_X1 U46bar ( .A1(abar[3]), .A2(bbar[11]), .ZN(ybar[59]) );
  AND2_X1 U47 ( .A1(a[3]), .A2(b[10]), .ZN(y[58]) );
  OR2_X1 U47bar ( .A1(abar[3]), .A2(bbar[10]), .ZN(ybar[58]) );
  AND2_X1 U48 ( .A1(a[3]), .A2(b[9]), .ZN(y[57]) );
  OR2_X1 U48bar ( .A1(abar[3]), .A2(bbar[9]), .ZN(ybar[57]) );
  AND2_X1 U49 ( .A1(a[3]), .A2(b[8]), .ZN(y[56]) );
  OR2_X1 U49bar ( .A1(abar[3]), .A2(bbar[8]), .ZN(ybar[56]) );
  AND2_X1 U50 ( .A1(a[3]), .A2(b[7]), .ZN(y[55]) );
  OR2_X1 U50bar ( .A1(abar[3]), .A2(bbar[7]), .ZN(ybar[55]) );
  AND2_X1 U51 ( .A1(a[3]), .A2(b[6]), .ZN(y[54]) );
  OR2_X1 U51bar ( .A1(abar[3]), .A2(bbar[6]), .ZN(ybar[54]) );
  AND2_X1 U52 ( .A1(a[3]), .A2(b[5]), .ZN(y[53]) );
  OR2_X1 U52bar ( .A1(abar[3]), .A2(bbar[5]), .ZN(ybar[53]) );
  AND2_X1 U53 ( .A1(a[3]), .A2(b[4]), .ZN(y[52]) );
  OR2_X1 U53bar ( .A1(abar[3]), .A2(bbar[4]), .ZN(ybar[52]) );
  AND2_X1 U54 ( .A1(a[3]), .A2(b[3]), .ZN(y[51]) );
  OR2_X1 U54bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[51]) );
  AND2_X1 U55 ( .A1(a[3]), .A2(b[2]), .ZN(y[50]) );
  OR2_X1 U55bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[50]) );
  AND2_X1 U56 ( .A1(b[4]), .A2(a[0]), .ZN(y[4]) );
  OR2_X1 U56bar ( .A1(bbar[4]), .A2(abar[0]), .ZN(ybar[4]) );
  AND2_X1 U57 ( .A1(a[3]), .A2(b[1]), .ZN(y[49]) );
  OR2_X1 U57bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[49]) );
  AND2_X1 U58 ( .A1(a[3]), .A2(b[0]), .ZN(y[48]) );
  OR2_X1 U58bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[48]) );
  AND2_X1 U59 ( .A1(a[2]), .A2(b[15]), .ZN(y[47]) );
  OR2_X1 U59bar ( .A1(abar[2]), .A2(bbar[15]), .ZN(ybar[47]) );
  AND2_X1 U60 ( .A1(a[2]), .A2(b[14]), .ZN(y[46]) );
  OR2_X1 U60bar ( .A1(abar[2]), .A2(bbar[14]), .ZN(ybar[46]) );
  AND2_X1 U61 ( .A1(a[2]), .A2(b[13]), .ZN(y[45]) );
  OR2_X1 U61bar ( .A1(abar[2]), .A2(bbar[13]), .ZN(ybar[45]) );
  AND2_X1 U62 ( .A1(a[2]), .A2(b[12]), .ZN(y[44]) );
  OR2_X1 U62bar ( .A1(abar[2]), .A2(bbar[12]), .ZN(ybar[44]) );
  AND2_X1 U63 ( .A1(a[2]), .A2(b[11]), .ZN(y[43]) );
  OR2_X1 U63bar ( .A1(abar[2]), .A2(bbar[11]), .ZN(ybar[43]) );
  AND2_X1 U64 ( .A1(a[2]), .A2(b[10]), .ZN(y[42]) );
  OR2_X1 U64bar ( .A1(abar[2]), .A2(bbar[10]), .ZN(ybar[42]) );
  AND2_X1 U65 ( .A1(a[2]), .A2(b[9]), .ZN(y[41]) );
  OR2_X1 U65bar ( .A1(abar[2]), .A2(bbar[9]), .ZN(ybar[41]) );
  AND2_X1 U66 ( .A1(a[2]), .A2(b[8]), .ZN(y[40]) );
  OR2_X1 U66bar ( .A1(abar[2]), .A2(bbar[8]), .ZN(ybar[40]) );
  AND2_X1 U67 ( .A1(b[3]), .A2(a[0]), .ZN(y[3]) );
  OR2_X1 U67bar ( .A1(bbar[3]), .A2(abar[0]), .ZN(ybar[3]) );
  AND2_X1 U68 ( .A1(a[2]), .A2(b[7]), .ZN(y[39]) );
  OR2_X1 U68bar ( .A1(abar[2]), .A2(bbar[7]), .ZN(ybar[39]) );
  AND2_X1 U69 ( .A1(a[2]), .A2(b[6]), .ZN(y[38]) );
  OR2_X1 U69bar ( .A1(abar[2]), .A2(bbar[6]), .ZN(ybar[38]) );
  AND2_X1 U70 ( .A1(a[2]), .A2(b[5]), .ZN(y[37]) );
  OR2_X1 U70bar ( .A1(abar[2]), .A2(bbar[5]), .ZN(ybar[37]) );
  AND2_X1 U71 ( .A1(a[2]), .A2(b[4]), .ZN(y[36]) );
  OR2_X1 U71bar ( .A1(abar[2]), .A2(bbar[4]), .ZN(ybar[36]) );
  AND2_X1 U72 ( .A1(a[2]), .A2(b[3]), .ZN(y[35]) );
  OR2_X1 U72bar ( .A1(abar[2]), .A2(bbar[3]), .ZN(ybar[35]) );
  AND2_X1 U73 ( .A1(a[2]), .A2(b[2]), .ZN(y[34]) );
  OR2_X1 U73bar ( .A1(abar[2]), .A2(bbar[2]), .ZN(ybar[34]) );
  AND2_X1 U74 ( .A1(a[2]), .A2(b[1]), .ZN(y[33]) );
  OR2_X1 U74bar ( .A1(abar[2]), .A2(bbar[1]), .ZN(ybar[33]) );
  AND2_X1 U75 ( .A1(a[2]), .A2(b[0]), .ZN(y[32]) );
  OR2_X1 U75bar ( .A1(abar[2]), .A2(bbar[0]), .ZN(ybar[32]) );
  AND2_X1 U76 ( .A1(a[1]), .A2(b[15]), .ZN(y[31]) );
  OR2_X1 U76bar ( .A1(abar[1]), .A2(bbar[15]), .ZN(ybar[31]) );
  AND2_X1 U77 ( .A1(a[1]), .A2(b[14]), .ZN(y[30]) );
  OR2_X1 U77bar ( .A1(abar[1]), .A2(bbar[14]), .ZN(ybar[30]) );
  AND2_X1 U78 ( .A1(b[2]), .A2(a[0]), .ZN(y[2]) );
  OR2_X1 U78bar ( .A1(bbar[2]), .A2(abar[0]), .ZN(ybar[2]) );
  AND2_X1 U79 ( .A1(a[1]), .A2(b[13]), .ZN(y[29]) );
  OR2_X1 U79bar ( .A1(abar[1]), .A2(bbar[13]), .ZN(ybar[29]) );
  AND2_X1 U80 ( .A1(a[1]), .A2(b[12]), .ZN(y[28]) );
  OR2_X1 U80bar ( .A1(abar[1]), .A2(bbar[12]), .ZN(ybar[28]) );
  AND2_X1 U81 ( .A1(a[1]), .A2(b[11]), .ZN(y[27]) );
  OR2_X1 U81bar ( .A1(abar[1]), .A2(bbar[11]), .ZN(ybar[27]) );
  AND2_X1 U82 ( .A1(a[1]), .A2(b[10]), .ZN(y[26]) );
  OR2_X1 U82bar ( .A1(abar[1]), .A2(bbar[10]), .ZN(ybar[26]) );
  AND2_X1 U83 ( .A1(a[1]), .A2(b[9]), .ZN(y[25]) );
  OR2_X1 U83bar ( .A1(abar[1]), .A2(bbar[9]), .ZN(ybar[25]) );
  AND2_X1 U84 ( .A1(a[15]), .A2(b[15]), .ZN(y[255]) );
  OR2_X1 U84bar ( .A1(abar[15]), .A2(bbar[15]), .ZN(ybar[255]) );
  AND2_X1 U85 ( .A1(a[15]), .A2(b[14]), .ZN(y[254]) );
  OR2_X1 U85bar ( .A1(abar[15]), .A2(bbar[14]), .ZN(ybar[254]) );
  AND2_X1 U86 ( .A1(a[15]), .A2(b[13]), .ZN(y[253]) );
  OR2_X1 U86bar ( .A1(abar[15]), .A2(bbar[13]), .ZN(ybar[253]) );
  AND2_X1 U87 ( .A1(a[15]), .A2(b[12]), .ZN(y[252]) );
  OR2_X1 U87bar ( .A1(abar[15]), .A2(bbar[12]), .ZN(ybar[252]) );
  AND2_X1 U88 ( .A1(a[15]), .A2(b[11]), .ZN(y[251]) );
  OR2_X1 U88bar ( .A1(abar[15]), .A2(bbar[11]), .ZN(ybar[251]) );
  AND2_X1 U89 ( .A1(a[15]), .A2(b[10]), .ZN(y[250]) );
  OR2_X1 U89bar ( .A1(abar[15]), .A2(bbar[10]), .ZN(ybar[250]) );
  AND2_X1 U90 ( .A1(a[1]), .A2(b[8]), .ZN(y[24]) );
  OR2_X1 U90bar ( .A1(abar[1]), .A2(bbar[8]), .ZN(ybar[24]) );
  AND2_X1 U91 ( .A1(a[15]), .A2(b[9]), .ZN(y[249]) );
  OR2_X1 U91bar ( .A1(abar[15]), .A2(bbar[9]), .ZN(ybar[249]) );
  AND2_X1 U92 ( .A1(a[15]), .A2(b[8]), .ZN(y[248]) );
  OR2_X1 U92bar ( .A1(abar[15]), .A2(bbar[8]), .ZN(ybar[248]) );
  AND2_X1 U93 ( .A1(a[15]), .A2(b[7]), .ZN(y[247]) );
  OR2_X1 U93bar ( .A1(abar[15]), .A2(bbar[7]), .ZN(ybar[247]) );
  AND2_X1 U94 ( .A1(a[15]), .A2(b[6]), .ZN(y[246]) );
  OR2_X1 U94bar ( .A1(abar[15]), .A2(bbar[6]), .ZN(ybar[246]) );
  AND2_X1 U95 ( .A1(a[15]), .A2(b[5]), .ZN(y[245]) );
  OR2_X1 U95bar ( .A1(abar[15]), .A2(bbar[5]), .ZN(ybar[245]) );
  AND2_X1 U96 ( .A1(a[15]), .A2(b[4]), .ZN(y[244]) );
  OR2_X1 U96bar ( .A1(abar[15]), .A2(bbar[4]), .ZN(ybar[244]) );
  AND2_X1 U97 ( .A1(a[15]), .A2(b[3]), .ZN(y[243]) );
  OR2_X1 U97bar ( .A1(abar[15]), .A2(bbar[3]), .ZN(ybar[243]) );
  AND2_X1 U98 ( .A1(a[15]), .A2(b[2]), .ZN(y[242]) );
  OR2_X1 U98bar ( .A1(abar[15]), .A2(bbar[2]), .ZN(ybar[242]) );
  AND2_X1 U99 ( .A1(a[15]), .A2(b[1]), .ZN(y[241]) );
  OR2_X1 U99bar ( .A1(abar[15]), .A2(bbar[1]), .ZN(ybar[241]) );
  AND2_X1 U100 ( .A1(a[15]), .A2(b[0]), .ZN(y[240]) );
  OR2_X1 U100bar ( .A1(abar[15]), .A2(bbar[0]), .ZN(ybar[240]) );
  AND2_X1 U101 ( .A1(a[1]), .A2(b[7]), .ZN(y[23]) );
  OR2_X1 U101bar ( .A1(abar[1]), .A2(bbar[7]), .ZN(ybar[23]) );
  AND2_X1 U102 ( .A1(a[14]), .A2(b[15]), .ZN(y[239]) );
  OR2_X1 U102bar ( .A1(abar[14]), .A2(bbar[15]), .ZN(ybar[239]) );
  AND2_X1 U103 ( .A1(a[14]), .A2(b[14]), .ZN(y[238]) );
  OR2_X1 U103bar ( .A1(abar[14]), .A2(bbar[14]), .ZN(ybar[238]) );
  AND2_X1 U104 ( .A1(a[14]), .A2(b[13]), .ZN(y[237]) );
  OR2_X1 U104bar ( .A1(abar[14]), .A2(bbar[13]), .ZN(ybar[237]) );
  AND2_X1 U105 ( .A1(a[14]), .A2(b[12]), .ZN(y[236]) );
  OR2_X1 U105bar ( .A1(abar[14]), .A2(bbar[12]), .ZN(ybar[236]) );
  AND2_X1 U106 ( .A1(a[14]), .A2(b[11]), .ZN(y[235]) );
  OR2_X1 U106bar ( .A1(abar[14]), .A2(bbar[11]), .ZN(ybar[235]) );
  AND2_X1 U107 ( .A1(a[14]), .A2(b[10]), .ZN(y[234]) );
  OR2_X1 U107bar ( .A1(abar[14]), .A2(bbar[10]), .ZN(ybar[234]) );
  AND2_X1 U108 ( .A1(a[14]), .A2(b[9]), .ZN(y[233]) );
  OR2_X1 U108bar ( .A1(abar[14]), .A2(bbar[9]), .ZN(ybar[233]) );
  AND2_X1 U109 ( .A1(a[14]), .A2(b[8]), .ZN(y[232]) );
  OR2_X1 U109bar ( .A1(abar[14]), .A2(bbar[8]), .ZN(ybar[232]) );
  AND2_X1 U110 ( .A1(a[14]), .A2(b[7]), .ZN(y[231]) );
  OR2_X1 U110bar ( .A1(abar[14]), .A2(bbar[7]), .ZN(ybar[231]) );
  AND2_X1 U111 ( .A1(a[14]), .A2(b[6]), .ZN(y[230]) );
  OR2_X1 U111bar ( .A1(abar[14]), .A2(bbar[6]), .ZN(ybar[230]) );
  AND2_X1 U112 ( .A1(a[1]), .A2(b[6]), .ZN(y[22]) );
  OR2_X1 U112bar ( .A1(abar[1]), .A2(bbar[6]), .ZN(ybar[22]) );
  AND2_X1 U113 ( .A1(a[14]), .A2(b[5]), .ZN(y[229]) );
  OR2_X1 U113bar ( .A1(abar[14]), .A2(bbar[5]), .ZN(ybar[229]) );
  AND2_X1 U114 ( .A1(a[14]), .A2(b[4]), .ZN(y[228]) );
  OR2_X1 U114bar ( .A1(abar[14]), .A2(bbar[4]), .ZN(ybar[228]) );
  AND2_X1 U115 ( .A1(a[14]), .A2(b[3]), .ZN(y[227]) );
  OR2_X1 U115bar ( .A1(abar[14]), .A2(bbar[3]), .ZN(ybar[227]) );
  AND2_X1 U116 ( .A1(a[14]), .A2(b[2]), .ZN(y[226]) );
  OR2_X1 U116bar ( .A1(abar[14]), .A2(bbar[2]), .ZN(ybar[226]) );
  AND2_X1 U117 ( .A1(a[14]), .A2(b[1]), .ZN(y[225]) );
  OR2_X1 U117bar ( .A1(abar[14]), .A2(bbar[1]), .ZN(ybar[225]) );
  AND2_X1 U118 ( .A1(a[14]), .A2(b[0]), .ZN(y[224]) );
  OR2_X1 U118bar ( .A1(abar[14]), .A2(bbar[0]), .ZN(ybar[224]) );
  AND2_X1 U119 ( .A1(a[13]), .A2(b[15]), .ZN(y[223]) );
  OR2_X1 U119bar ( .A1(abar[13]), .A2(bbar[15]), .ZN(ybar[223]) );
  AND2_X1 U120 ( .A1(a[13]), .A2(b[14]), .ZN(y[222]) );
  OR2_X1 U120bar ( .A1(abar[13]), .A2(bbar[14]), .ZN(ybar[222]) );
  AND2_X1 U121 ( .A1(a[13]), .A2(b[13]), .ZN(y[221]) );
  OR2_X1 U121bar ( .A1(abar[13]), .A2(bbar[13]), .ZN(ybar[221]) );
  AND2_X1 U122 ( .A1(a[13]), .A2(b[12]), .ZN(y[220]) );
  OR2_X1 U122bar ( .A1(abar[13]), .A2(bbar[12]), .ZN(ybar[220]) );
  AND2_X1 U123 ( .A1(a[1]), .A2(b[5]), .ZN(y[21]) );
  OR2_X1 U123bar ( .A1(abar[1]), .A2(bbar[5]), .ZN(ybar[21]) );
  AND2_X1 U124 ( .A1(a[13]), .A2(b[11]), .ZN(y[219]) );
  OR2_X1 U124bar ( .A1(abar[13]), .A2(bbar[11]), .ZN(ybar[219]) );
  AND2_X1 U125 ( .A1(a[13]), .A2(b[10]), .ZN(y[218]) );
  OR2_X1 U125bar ( .A1(abar[13]), .A2(bbar[10]), .ZN(ybar[218]) );
  AND2_X1 U126 ( .A1(a[13]), .A2(b[9]), .ZN(y[217]) );
  OR2_X1 U126bar ( .A1(abar[13]), .A2(bbar[9]), .ZN(ybar[217]) );
  AND2_X1 U127 ( .A1(a[13]), .A2(b[8]), .ZN(y[216]) );
  OR2_X1 U127bar ( .A1(abar[13]), .A2(bbar[8]), .ZN(ybar[216]) );
  AND2_X1 U128 ( .A1(a[13]), .A2(b[7]), .ZN(y[215]) );
  OR2_X1 U128bar ( .A1(abar[13]), .A2(bbar[7]), .ZN(ybar[215]) );
  AND2_X1 U129 ( .A1(a[13]), .A2(b[6]), .ZN(y[214]) );
  OR2_X1 U129bar ( .A1(abar[13]), .A2(bbar[6]), .ZN(ybar[214]) );
  AND2_X1 U130 ( .A1(a[13]), .A2(b[5]), .ZN(y[213]) );
  OR2_X1 U130bar ( .A1(abar[13]), .A2(bbar[5]), .ZN(ybar[213]) );
  AND2_X1 U131 ( .A1(a[13]), .A2(b[4]), .ZN(y[212]) );
  OR2_X1 U131bar ( .A1(abar[13]), .A2(bbar[4]), .ZN(ybar[212]) );
  AND2_X1 U132 ( .A1(a[13]), .A2(b[3]), .ZN(y[211]) );
  OR2_X1 U132bar ( .A1(abar[13]), .A2(bbar[3]), .ZN(ybar[211]) );
  AND2_X1 U133 ( .A1(a[13]), .A2(b[2]), .ZN(y[210]) );
  OR2_X1 U133bar ( .A1(abar[13]), .A2(bbar[2]), .ZN(ybar[210]) );
  AND2_X1 U134 ( .A1(a[1]), .A2(b[4]), .ZN(y[20]) );
  OR2_X1 U134bar ( .A1(abar[1]), .A2(bbar[4]), .ZN(ybar[20]) );
  AND2_X1 U135 ( .A1(a[13]), .A2(b[1]), .ZN(y[209]) );
  OR2_X1 U135bar ( .A1(abar[13]), .A2(bbar[1]), .ZN(ybar[209]) );
  AND2_X1 U136 ( .A1(a[13]), .A2(b[0]), .ZN(y[208]) );
  OR2_X1 U136bar ( .A1(abar[13]), .A2(bbar[0]), .ZN(ybar[208]) );
  AND2_X1 U137 ( .A1(a[12]), .A2(b[15]), .ZN(y[207]) );
  OR2_X1 U137bar ( .A1(abar[12]), .A2(bbar[15]), .ZN(ybar[207]) );
  AND2_X1 U138 ( .A1(a[12]), .A2(b[14]), .ZN(y[206]) );
  OR2_X1 U138bar ( .A1(abar[12]), .A2(bbar[14]), .ZN(ybar[206]) );
  AND2_X1 U139 ( .A1(a[12]), .A2(b[13]), .ZN(y[205]) );
  OR2_X1 U139bar ( .A1(abar[12]), .A2(bbar[13]), .ZN(ybar[205]) );
  AND2_X1 U140 ( .A1(a[12]), .A2(b[12]), .ZN(y[204]) );
  OR2_X1 U140bar ( .A1(abar[12]), .A2(bbar[12]), .ZN(ybar[204]) );
  AND2_X1 U141 ( .A1(a[12]), .A2(b[11]), .ZN(y[203]) );
  OR2_X1 U141bar ( .A1(abar[12]), .A2(bbar[11]), .ZN(ybar[203]) );
  AND2_X1 U142 ( .A1(a[12]), .A2(b[10]), .ZN(y[202]) );
  OR2_X1 U142bar ( .A1(abar[12]), .A2(bbar[10]), .ZN(ybar[202]) );
  AND2_X1 U143 ( .A1(a[12]), .A2(b[9]), .ZN(y[201]) );
  OR2_X1 U143bar ( .A1(abar[12]), .A2(bbar[9]), .ZN(ybar[201]) );
  AND2_X1 U144 ( .A1(a[12]), .A2(b[8]), .ZN(y[200]) );
  OR2_X1 U144bar ( .A1(abar[12]), .A2(bbar[8]), .ZN(ybar[200]) );
  AND2_X1 U145 ( .A1(b[1]), .A2(a[0]), .ZN(y[1]) );
  OR2_X1 U145bar ( .A1(bbar[1]), .A2(abar[0]), .ZN(ybar[1]) );
  AND2_X1 U146 ( .A1(a[1]), .A2(b[3]), .ZN(y[19]) );
  OR2_X1 U146bar ( .A1(abar[1]), .A2(bbar[3]), .ZN(ybar[19]) );
  AND2_X1 U147 ( .A1(a[12]), .A2(b[7]), .ZN(y[199]) );
  OR2_X1 U147bar ( .A1(abar[12]), .A2(bbar[7]), .ZN(ybar[199]) );
  AND2_X1 U148 ( .A1(a[12]), .A2(b[6]), .ZN(y[198]) );
  OR2_X1 U148bar ( .A1(abar[12]), .A2(bbar[6]), .ZN(ybar[198]) );
  AND2_X1 U149 ( .A1(a[12]), .A2(b[5]), .ZN(y[197]) );
  OR2_X1 U149bar ( .A1(abar[12]), .A2(bbar[5]), .ZN(ybar[197]) );
  AND2_X1 U150 ( .A1(a[12]), .A2(b[4]), .ZN(y[196]) );
  OR2_X1 U150bar ( .A1(abar[12]), .A2(bbar[4]), .ZN(ybar[196]) );
  AND2_X1 U151 ( .A1(a[12]), .A2(b[3]), .ZN(y[195]) );
  OR2_X1 U151bar ( .A1(abar[12]), .A2(bbar[3]), .ZN(ybar[195]) );
  AND2_X1 U152 ( .A1(a[12]), .A2(b[2]), .ZN(y[194]) );
  OR2_X1 U152bar ( .A1(abar[12]), .A2(bbar[2]), .ZN(ybar[194]) );
  AND2_X1 U153 ( .A1(a[12]), .A2(b[1]), .ZN(y[193]) );
  OR2_X1 U153bar ( .A1(abar[12]), .A2(bbar[1]), .ZN(ybar[193]) );
  AND2_X1 U154 ( .A1(a[12]), .A2(b[0]), .ZN(y[192]) );
  OR2_X1 U154bar ( .A1(abar[12]), .A2(bbar[0]), .ZN(ybar[192]) );
  AND2_X1 U155 ( .A1(a[11]), .A2(b[15]), .ZN(y[191]) );
  OR2_X1 U155bar ( .A1(abar[11]), .A2(bbar[15]), .ZN(ybar[191]) );
  AND2_X1 U156 ( .A1(a[11]), .A2(b[14]), .ZN(y[190]) );
  OR2_X1 U156bar ( .A1(abar[11]), .A2(bbar[14]), .ZN(ybar[190]) );
  AND2_X1 U157 ( .A1(a[1]), .A2(b[2]), .ZN(y[18]) );
  OR2_X1 U157bar ( .A1(abar[1]), .A2(bbar[2]), .ZN(ybar[18]) );
  AND2_X1 U158 ( .A1(a[11]), .A2(b[13]), .ZN(y[189]) );
  OR2_X1 U158bar ( .A1(abar[11]), .A2(bbar[13]), .ZN(ybar[189]) );
  AND2_X1 U159 ( .A1(a[11]), .A2(b[12]), .ZN(y[188]) );
  OR2_X1 U159bar ( .A1(abar[11]), .A2(bbar[12]), .ZN(ybar[188]) );
  AND2_X1 U160 ( .A1(a[11]), .A2(b[11]), .ZN(y[187]) );
  OR2_X1 U160bar ( .A1(abar[11]), .A2(bbar[11]), .ZN(ybar[187]) );
  AND2_X1 U161 ( .A1(a[11]), .A2(b[10]), .ZN(y[186]) );
  OR2_X1 U161bar ( .A1(abar[11]), .A2(bbar[10]), .ZN(ybar[186]) );
  AND2_X1 U162 ( .A1(a[11]), .A2(b[9]), .ZN(y[185]) );
  OR2_X1 U162bar ( .A1(abar[11]), .A2(bbar[9]), .ZN(ybar[185]) );
  AND2_X1 U163 ( .A1(a[11]), .A2(b[8]), .ZN(y[184]) );
  OR2_X1 U163bar ( .A1(abar[11]), .A2(bbar[8]), .ZN(ybar[184]) );
  AND2_X1 U164 ( .A1(a[11]), .A2(b[7]), .ZN(y[183]) );
  OR2_X1 U164bar ( .A1(abar[11]), .A2(bbar[7]), .ZN(ybar[183]) );
  AND2_X1 U165 ( .A1(a[11]), .A2(b[6]), .ZN(y[182]) );
  OR2_X1 U165bar ( .A1(abar[11]), .A2(bbar[6]), .ZN(ybar[182]) );
  AND2_X1 U166 ( .A1(a[11]), .A2(b[5]), .ZN(y[181]) );
  OR2_X1 U166bar ( .A1(abar[11]), .A2(bbar[5]), .ZN(ybar[181]) );
  AND2_X1 U167 ( .A1(a[11]), .A2(b[4]), .ZN(y[180]) );
  OR2_X1 U167bar ( .A1(abar[11]), .A2(bbar[4]), .ZN(ybar[180]) );
  AND2_X1 U168 ( .A1(a[1]), .A2(b[1]), .ZN(y[17]) );
  OR2_X1 U168bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[17]) );
  AND2_X1 U169 ( .A1(a[11]), .A2(b[3]), .ZN(y[179]) );
  OR2_X1 U169bar ( .A1(abar[11]), .A2(bbar[3]), .ZN(ybar[179]) );
  AND2_X1 U170 ( .A1(a[11]), .A2(b[2]), .ZN(y[178]) );
  OR2_X1 U170bar ( .A1(abar[11]), .A2(bbar[2]), .ZN(ybar[178]) );
  AND2_X1 U171 ( .A1(a[11]), .A2(b[1]), .ZN(y[177]) );
  OR2_X1 U171bar ( .A1(abar[11]), .A2(bbar[1]), .ZN(ybar[177]) );
  AND2_X1 U172 ( .A1(a[11]), .A2(b[0]), .ZN(y[176]) );
  OR2_X1 U172bar ( .A1(abar[11]), .A2(bbar[0]), .ZN(ybar[176]) );
  AND2_X1 U173 ( .A1(a[10]), .A2(b[15]), .ZN(y[175]) );
  OR2_X1 U173bar ( .A1(abar[10]), .A2(bbar[15]), .ZN(ybar[175]) );
  AND2_X1 U174 ( .A1(a[10]), .A2(b[14]), .ZN(y[174]) );
  OR2_X1 U174bar ( .A1(abar[10]), .A2(bbar[14]), .ZN(ybar[174]) );
  AND2_X1 U175 ( .A1(a[10]), .A2(b[13]), .ZN(y[173]) );
  OR2_X1 U175bar ( .A1(abar[10]), .A2(bbar[13]), .ZN(ybar[173]) );
  AND2_X1 U176 ( .A1(a[10]), .A2(b[12]), .ZN(y[172]) );
  OR2_X1 U176bar ( .A1(abar[10]), .A2(bbar[12]), .ZN(ybar[172]) );
  AND2_X1 U177 ( .A1(a[10]), .A2(b[11]), .ZN(y[171]) );
  OR2_X1 U177bar ( .A1(abar[10]), .A2(bbar[11]), .ZN(ybar[171]) );
  AND2_X1 U178 ( .A1(a[10]), .A2(b[10]), .ZN(y[170]) );
  OR2_X1 U178bar ( .A1(abar[10]), .A2(bbar[10]), .ZN(ybar[170]) );
  AND2_X1 U179 ( .A1(a[1]), .A2(b[0]), .ZN(y[16]) );
  OR2_X1 U179bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[16]) );
  AND2_X1 U180 ( .A1(a[10]), .A2(b[9]), .ZN(y[169]) );
  OR2_X1 U180bar ( .A1(abar[10]), .A2(bbar[9]), .ZN(ybar[169]) );
  AND2_X1 U181 ( .A1(a[10]), .A2(b[8]), .ZN(y[168]) );
  OR2_X1 U181bar ( .A1(abar[10]), .A2(bbar[8]), .ZN(ybar[168]) );
  AND2_X1 U182 ( .A1(a[10]), .A2(b[7]), .ZN(y[167]) );
  OR2_X1 U182bar ( .A1(abar[10]), .A2(bbar[7]), .ZN(ybar[167]) );
  AND2_X1 U183 ( .A1(a[10]), .A2(b[6]), .ZN(y[166]) );
  OR2_X1 U183bar ( .A1(abar[10]), .A2(bbar[6]), .ZN(ybar[166]) );
  AND2_X1 U184 ( .A1(a[10]), .A2(b[5]), .ZN(y[165]) );
  OR2_X1 U184bar ( .A1(abar[10]), .A2(bbar[5]), .ZN(ybar[165]) );
  AND2_X1 U185 ( .A1(a[10]), .A2(b[4]), .ZN(y[164]) );
  OR2_X1 U185bar ( .A1(abar[10]), .A2(bbar[4]), .ZN(ybar[164]) );
  AND2_X1 U186 ( .A1(a[10]), .A2(b[3]), .ZN(y[163]) );
  OR2_X1 U186bar ( .A1(abar[10]), .A2(bbar[3]), .ZN(ybar[163]) );
  AND2_X1 U187 ( .A1(a[10]), .A2(b[2]), .ZN(y[162]) );
  OR2_X1 U187bar ( .A1(abar[10]), .A2(bbar[2]), .ZN(ybar[162]) );
  AND2_X1 U188 ( .A1(a[10]), .A2(b[1]), .ZN(y[161]) );
  OR2_X1 U188bar ( .A1(abar[10]), .A2(bbar[1]), .ZN(ybar[161]) );
  AND2_X1 U189 ( .A1(a[10]), .A2(b[0]), .ZN(y[160]) );
  OR2_X1 U189bar ( .A1(abar[10]), .A2(bbar[0]), .ZN(ybar[160]) );
  AND2_X1 U190 ( .A1(b[15]), .A2(a[0]), .ZN(y[15]) );
  OR2_X1 U190bar ( .A1(bbar[15]), .A2(abar[0]), .ZN(ybar[15]) );
  AND2_X1 U191 ( .A1(a[9]), .A2(b[15]), .ZN(y[159]) );
  OR2_X1 U191bar ( .A1(abar[9]), .A2(bbar[15]), .ZN(ybar[159]) );
  AND2_X1 U192 ( .A1(a[9]), .A2(b[14]), .ZN(y[158]) );
  OR2_X1 U192bar ( .A1(abar[9]), .A2(bbar[14]), .ZN(ybar[158]) );
  AND2_X1 U193 ( .A1(a[9]), .A2(b[13]), .ZN(y[157]) );
  OR2_X1 U193bar ( .A1(abar[9]), .A2(bbar[13]), .ZN(ybar[157]) );
  AND2_X1 U194 ( .A1(a[9]), .A2(b[12]), .ZN(y[156]) );
  OR2_X1 U194bar ( .A1(abar[9]), .A2(bbar[12]), .ZN(ybar[156]) );
  AND2_X1 U195 ( .A1(a[9]), .A2(b[11]), .ZN(y[155]) );
  OR2_X1 U195bar ( .A1(abar[9]), .A2(bbar[11]), .ZN(ybar[155]) );
  AND2_X1 U196 ( .A1(a[9]), .A2(b[10]), .ZN(y[154]) );
  OR2_X1 U196bar ( .A1(abar[9]), .A2(bbar[10]), .ZN(ybar[154]) );
  AND2_X1 U197 ( .A1(a[9]), .A2(b[9]), .ZN(y[153]) );
  OR2_X1 U197bar ( .A1(abar[9]), .A2(bbar[9]), .ZN(ybar[153]) );
  AND2_X1 U198 ( .A1(a[9]), .A2(b[8]), .ZN(y[152]) );
  OR2_X1 U198bar ( .A1(abar[9]), .A2(bbar[8]), .ZN(ybar[152]) );
  AND2_X1 U199 ( .A1(a[9]), .A2(b[7]), .ZN(y[151]) );
  OR2_X1 U199bar ( .A1(abar[9]), .A2(bbar[7]), .ZN(ybar[151]) );
  AND2_X1 U200 ( .A1(a[9]), .A2(b[6]), .ZN(y[150]) );
  OR2_X1 U200bar ( .A1(abar[9]), .A2(bbar[6]), .ZN(ybar[150]) );
  AND2_X1 U201 ( .A1(b[14]), .A2(a[0]), .ZN(y[14]) );
  OR2_X1 U201bar ( .A1(bbar[14]), .A2(abar[0]), .ZN(ybar[14]) );
  AND2_X1 U202 ( .A1(a[9]), .A2(b[5]), .ZN(y[149]) );
  OR2_X1 U202bar ( .A1(abar[9]), .A2(bbar[5]), .ZN(ybar[149]) );
  AND2_X1 U203 ( .A1(a[9]), .A2(b[4]), .ZN(y[148]) );
  OR2_X1 U203bar ( .A1(abar[9]), .A2(bbar[4]), .ZN(ybar[148]) );
  AND2_X1 U204 ( .A1(a[9]), .A2(b[3]), .ZN(y[147]) );
  OR2_X1 U204bar ( .A1(abar[9]), .A2(bbar[3]), .ZN(ybar[147]) );
  AND2_X1 U205 ( .A1(a[9]), .A2(b[2]), .ZN(y[146]) );
  OR2_X1 U205bar ( .A1(abar[9]), .A2(bbar[2]), .ZN(ybar[146]) );
  AND2_X1 U206 ( .A1(a[9]), .A2(b[1]), .ZN(y[145]) );
  OR2_X1 U206bar ( .A1(abar[9]), .A2(bbar[1]), .ZN(ybar[145]) );
  AND2_X1 U207 ( .A1(a[9]), .A2(b[0]), .ZN(y[144]) );
  OR2_X1 U207bar ( .A1(abar[9]), .A2(bbar[0]), .ZN(ybar[144]) );
  AND2_X1 U208 ( .A1(a[8]), .A2(b[15]), .ZN(y[143]) );
  OR2_X1 U208bar ( .A1(abar[8]), .A2(bbar[15]), .ZN(ybar[143]) );
  AND2_X1 U209 ( .A1(a[8]), .A2(b[14]), .ZN(y[142]) );
  OR2_X1 U209bar ( .A1(abar[8]), .A2(bbar[14]), .ZN(ybar[142]) );
  AND2_X1 U210 ( .A1(a[8]), .A2(b[13]), .ZN(y[141]) );
  OR2_X1 U210bar ( .A1(abar[8]), .A2(bbar[13]), .ZN(ybar[141]) );
  AND2_X1 U211 ( .A1(a[8]), .A2(b[12]), .ZN(y[140]) );
  OR2_X1 U211bar ( .A1(abar[8]), .A2(bbar[12]), .ZN(ybar[140]) );
  AND2_X1 U212 ( .A1(b[13]), .A2(a[0]), .ZN(y[13]) );
  OR2_X1 U212bar ( .A1(bbar[13]), .A2(abar[0]), .ZN(ybar[13]) );
  AND2_X1 U213 ( .A1(a[8]), .A2(b[11]), .ZN(y[139]) );
  OR2_X1 U213bar ( .A1(abar[8]), .A2(bbar[11]), .ZN(ybar[139]) );
  AND2_X1 U214 ( .A1(a[8]), .A2(b[10]), .ZN(y[138]) );
  OR2_X1 U214bar ( .A1(abar[8]), .A2(bbar[10]), .ZN(ybar[138]) );
  AND2_X1 U215 ( .A1(a[8]), .A2(b[9]), .ZN(y[137]) );
  OR2_X1 U215bar ( .A1(abar[8]), .A2(bbar[9]), .ZN(ybar[137]) );
  AND2_X1 U216 ( .A1(a[8]), .A2(b[8]), .ZN(y[136]) );
  OR2_X1 U216bar ( .A1(abar[8]), .A2(bbar[8]), .ZN(ybar[136]) );
  AND2_X1 U217 ( .A1(a[8]), .A2(b[7]), .ZN(y[135]) );
  OR2_X1 U217bar ( .A1(abar[8]), .A2(bbar[7]), .ZN(ybar[135]) );
  AND2_X1 U218 ( .A1(a[8]), .A2(b[6]), .ZN(y[134]) );
  OR2_X1 U218bar ( .A1(abar[8]), .A2(bbar[6]), .ZN(ybar[134]) );
  AND2_X1 U219 ( .A1(a[8]), .A2(b[5]), .ZN(y[133]) );
  OR2_X1 U219bar ( .A1(abar[8]), .A2(bbar[5]), .ZN(ybar[133]) );
  AND2_X1 U220 ( .A1(a[8]), .A2(b[4]), .ZN(y[132]) );
  OR2_X1 U220bar ( .A1(abar[8]), .A2(bbar[4]), .ZN(ybar[132]) );
  AND2_X1 U221 ( .A1(a[8]), .A2(b[3]), .ZN(y[131]) );
  OR2_X1 U221bar ( .A1(abar[8]), .A2(bbar[3]), .ZN(ybar[131]) );
  AND2_X1 U222 ( .A1(a[8]), .A2(b[2]), .ZN(y[130]) );
  OR2_X1 U222bar ( .A1(abar[8]), .A2(bbar[2]), .ZN(ybar[130]) );
  AND2_X1 U223 ( .A1(b[12]), .A2(a[0]), .ZN(y[12]) );
  OR2_X1 U223bar ( .A1(bbar[12]), .A2(abar[0]), .ZN(ybar[12]) );
  AND2_X1 U224 ( .A1(a[8]), .A2(b[1]), .ZN(y[129]) );
  OR2_X1 U224bar ( .A1(abar[8]), .A2(bbar[1]), .ZN(ybar[129]) );
  AND2_X1 U225 ( .A1(a[8]), .A2(b[0]), .ZN(y[128]) );
  OR2_X1 U225bar ( .A1(abar[8]), .A2(bbar[0]), .ZN(ybar[128]) );
  AND2_X1 U226 ( .A1(a[7]), .A2(b[15]), .ZN(y[127]) );
  OR2_X1 U226bar ( .A1(abar[7]), .A2(bbar[15]), .ZN(ybar[127]) );
  AND2_X1 U227 ( .A1(a[7]), .A2(b[14]), .ZN(y[126]) );
  OR2_X1 U227bar ( .A1(abar[7]), .A2(bbar[14]), .ZN(ybar[126]) );
  AND2_X1 U228 ( .A1(a[7]), .A2(b[13]), .ZN(y[125]) );
  OR2_X1 U228bar ( .A1(abar[7]), .A2(bbar[13]), .ZN(ybar[125]) );
  AND2_X1 U229 ( .A1(a[7]), .A2(b[12]), .ZN(y[124]) );
  OR2_X1 U229bar ( .A1(abar[7]), .A2(bbar[12]), .ZN(ybar[124]) );
  AND2_X1 U230 ( .A1(a[7]), .A2(b[11]), .ZN(y[123]) );
  OR2_X1 U230bar ( .A1(abar[7]), .A2(bbar[11]), .ZN(ybar[123]) );
  AND2_X1 U231 ( .A1(a[7]), .A2(b[10]), .ZN(y[122]) );
  OR2_X1 U231bar ( .A1(abar[7]), .A2(bbar[10]), .ZN(ybar[122]) );
  AND2_X1 U232 ( .A1(a[7]), .A2(b[9]), .ZN(y[121]) );
  OR2_X1 U232bar ( .A1(abar[7]), .A2(bbar[9]), .ZN(ybar[121]) );
  AND2_X1 U233 ( .A1(a[7]), .A2(b[8]), .ZN(y[120]) );
  OR2_X1 U233bar ( .A1(abar[7]), .A2(bbar[8]), .ZN(ybar[120]) );
  AND2_X1 U234 ( .A1(b[11]), .A2(a[0]), .ZN(y[11]) );
  OR2_X1 U234bar ( .A1(bbar[11]), .A2(abar[0]), .ZN(ybar[11]) );
  AND2_X1 U235 ( .A1(a[7]), .A2(b[7]), .ZN(y[119]) );
  OR2_X1 U235bar ( .A1(abar[7]), .A2(bbar[7]), .ZN(ybar[119]) );
  AND2_X1 U236 ( .A1(a[7]), .A2(b[6]), .ZN(y[118]) );
  OR2_X1 U236bar ( .A1(abar[7]), .A2(bbar[6]), .ZN(ybar[118]) );
  AND2_X1 U237 ( .A1(a[7]), .A2(b[5]), .ZN(y[117]) );
  OR2_X1 U237bar ( .A1(abar[7]), .A2(bbar[5]), .ZN(ybar[117]) );
  AND2_X1 U238 ( .A1(a[7]), .A2(b[4]), .ZN(y[116]) );
  OR2_X1 U238bar ( .A1(abar[7]), .A2(bbar[4]), .ZN(ybar[116]) );
  AND2_X1 U239 ( .A1(a[7]), .A2(b[3]), .ZN(y[115]) );
  OR2_X1 U239bar ( .A1(abar[7]), .A2(bbar[3]), .ZN(ybar[115]) );
  AND2_X1 U240 ( .A1(a[7]), .A2(b[2]), .ZN(y[114]) );
  OR2_X1 U240bar ( .A1(abar[7]), .A2(bbar[2]), .ZN(ybar[114]) );
  AND2_X1 U241 ( .A1(a[7]), .A2(b[1]), .ZN(y[113]) );
  OR2_X1 U241bar ( .A1(abar[7]), .A2(bbar[1]), .ZN(ybar[113]) );
  AND2_X1 U242 ( .A1(a[7]), .A2(b[0]), .ZN(y[112]) );
  OR2_X1 U242bar ( .A1(abar[7]), .A2(bbar[0]), .ZN(ybar[112]) );
  AND2_X1 U243 ( .A1(b[15]), .A2(a[6]), .ZN(y[111]) );
  OR2_X1 U243bar ( .A1(bbar[15]), .A2(abar[6]), .ZN(ybar[111]) );
  AND2_X1 U244 ( .A1(b[14]), .A2(a[6]), .ZN(y[110]) );
  OR2_X1 U244bar ( .A1(bbar[14]), .A2(abar[6]), .ZN(ybar[110]) );
  AND2_X1 U245 ( .A1(b[10]), .A2(a[0]), .ZN(y[10]) );
  OR2_X1 U245bar ( .A1(bbar[10]), .A2(abar[0]), .ZN(ybar[10]) );
  AND2_X1 U246 ( .A1(b[13]), .A2(a[6]), .ZN(y[109]) );
  OR2_X1 U246bar ( .A1(bbar[13]), .A2(abar[6]), .ZN(ybar[109]) );
  AND2_X1 U247 ( .A1(b[12]), .A2(a[6]), .ZN(y[108]) );
  OR2_X1 U247bar ( .A1(bbar[12]), .A2(abar[6]), .ZN(ybar[108]) );
  AND2_X1 U248 ( .A1(b[11]), .A2(a[6]), .ZN(y[107]) );
  OR2_X1 U248bar ( .A1(bbar[11]), .A2(abar[6]), .ZN(ybar[107]) );
  AND2_X1 U249 ( .A1(b[10]), .A2(a[6]), .ZN(y[106]) );
  OR2_X1 U249bar ( .A1(bbar[10]), .A2(abar[6]), .ZN(ybar[106]) );
  AND2_X1 U250 ( .A1(a[6]), .A2(b[9]), .ZN(y[105]) );
  OR2_X1 U250bar ( .A1(abar[6]), .A2(bbar[9]), .ZN(ybar[105]) );
  AND2_X1 U251 ( .A1(b[8]), .A2(a[6]), .ZN(y[104]) );
  OR2_X1 U251bar ( .A1(bbar[8]), .A2(abar[6]), .ZN(ybar[104]) );
  AND2_X1 U252 ( .A1(b[7]), .A2(a[6]), .ZN(y[103]) );
  OR2_X1 U252bar ( .A1(bbar[7]), .A2(abar[6]), .ZN(ybar[103]) );
  AND2_X1 U253 ( .A1(b[6]), .A2(a[6]), .ZN(y[102]) );
  OR2_X1 U253bar ( .A1(bbar[6]), .A2(abar[6]), .ZN(ybar[102]) );
  AND2_X1 U254 ( .A1(b[5]), .A2(a[6]), .ZN(y[101]) );
  OR2_X1 U254bar ( .A1(bbar[5]), .A2(abar[6]), .ZN(ybar[101]) );
  AND2_X1 U255 ( .A1(b[4]), .A2(a[6]), .ZN(y[100]) );
  OR2_X1 U255bar ( .A1(bbar[4]), .A2(abar[6]), .ZN(ybar[100]) );
  AND2_X1 U256 ( .A1(b[0]), .A2(a[0]), .ZN(y[0]) );
  OR2_X1 U256bar ( .A1(bbar[0]), .A2(abar[0]), .ZN(ybar[0]) );
endmodule

module decode_3 ( in, inbar, out, outbar );

  input wire [7:0] in;
  input wire [7:0] inbar;
//input_done

  output wire [255:0] out;
  output wire [255:0] outbar;
//output_done

  wire [15:0] level1;
  wire [31:0] level2;
  wire [15:0] level1bar;
  wire [31:0] level2bar;
//wire_done

  CD2_12 cd_l1_1 ( .a(in[1]), .abar(inbar[1]), .b(in[0]), .bbar(inbar[0]), .y(level1[3:0]), .ybar(level1bar[3:0]) );
  CD2_11 cd_l1_2 ( .a(in[3]), .abar(inbar[3]), .b(in[2]), .bbar(inbar[2]), .y(level1[7:4]), .ybar(level1bar[7:4]) );
  CD2_10 cd_l1_3 ( .a(in[5]), .abar(inbar[5]), .b(in[4]), .bbar(inbar[4]), .y(level1[11:8]), .ybar(level1bar[11:8]) );
  CD2_9 cd_l1_4 ( .a(in[7]), .abar(inbar[7]), .b(in[6]), .bbar(inbar[6]), .y(level1[15:12]), .ybar(level1bar[15:12]) );

  CD4_6 cd_l2_1 ( .a(level1[7:4]), .abar(level1bar[7:4]), .b(level1[3:0]), .bbar(level1bar[3:0]), 
        .y(level2[15:0]), .ybar(level2bar[15:0]) );
  CD4_5 cd_l2_2 ( .a(level1[15:12]), .abar(level1bar[15:12]), .b(level1[11:8]), .bbar(level1bar[11:8]), 
        .y(level2[31:16]), .ybar(level2bar[31:16]) );
  CD16_3 cd_l3 ( .a(level2[31:16]), .abar(level2bar[31:16]), .b(level2[15:0]), .bbar(level2bar[15:0]), 
        .y(out), .ybar(outbar) );
endmodule

module encode_3 ( in, inbar, out, outbar );

  input wire [255:0] in;
  input wire [255:0] inbar;
//input_done

  output wire [7:0] out;
  output wire [7:0] outbar;
//output_done

  wire in_81;
  wire in_80;
  wire in_79;
  wire in_78;
  wire in_77;
  wire in_76;
  wire in_75;
  wire in_74;
  wire in_73;
  wire in_72;
  wire in_71;
  wire in_70;
  wire in_69;
  wire in_68;
  wire in_67;
  wire in_66;
  wire in_65;
  wire in_64;
  wire in_63;
  wire in_62;
  wire in_61;
  wire in_60;
  wire in_59;
  wire in_58;
  wire in_57;
  wire in_56;
  wire in_55;
  wire in_54;
  wire in_53;
  wire in_52;
  wire in_51;
  wire in_50;
  wire in_49;
  wire in_48;
  wire in_47;
  wire in_46;
  wire in_45;
  wire in_44;
  wire in_43;
  wire in_42;
  wire in_41;
  wire in_40;
  wire in_39;
  wire in_38;
  wire in_37;
  wire in_36;
  wire in_35;
  wire in_34;
  wire in_33;
  wire in_32;
  wire in_31;
  wire in_30;
  wire in_29;
  wire in_28;
  wire in_27;
  wire in_26;
  wire in_25;
  wire in_24;
  wire in_23;
  wire in_22;
  wire in_21;
  wire in_20;
  wire in_19;
  wire in_18;
  wire in_17;
  wire in_16;
  wire in_15;
  wire in_14;
  wire in_13;
  wire in_12;
  wire in_11;
  wire in_10;
  wire in_9;
  wire in_8;
  wire in_7;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_3;
  wire in_2;
  wire in_1;
  wire in_0;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire in_81bar;
  wire in_80bar;
  wire in_79bar;
  wire in_78bar;
  wire in_77bar;
  wire in_76bar;
  wire in_75bar;
  wire in_74bar;
  wire in_73bar;
  wire in_72bar;
  wire in_71bar;
  wire in_70bar;
  wire in_69bar;
  wire in_68bar;
  wire in_67bar;
  wire in_66bar;
  wire in_65bar;
  wire in_64bar;
  wire in_63bar;
  wire in_62bar;
  wire in_61bar;
  wire in_60bar;
  wire in_59bar;
  wire in_58bar;
  wire in_57bar;
  wire in_56bar;
  wire in_55bar;
  wire in_54bar;
  wire in_53bar;
  wire in_52bar;
  wire in_51bar;
  wire in_50bar;
  wire in_49bar;
  wire in_48bar;
  wire in_47bar;
  wire in_46bar;
  wire in_45bar;
  wire in_44bar;
  wire in_43bar;
  wire in_42bar;
  wire in_41bar;
  wire in_40bar;
  wire in_39bar;
  wire in_38bar;
  wire in_37bar;
  wire in_36bar;
  wire in_35bar;
  wire in_34bar;
  wire in_33bar;
  wire in_32bar;
  wire in_31bar;
  wire in_30bar;
  wire in_29bar;
  wire in_28bar;
  wire in_27bar;
  wire in_26bar;
  wire in_25bar;
  wire in_24bar;
  wire in_23bar;
  wire in_22bar;
  wire in_21bar;
  wire in_20bar;
  wire in_19bar;
  wire in_18bar;
  wire in_17bar;
  wire in_16bar;
  wire in_15bar;
  wire in_14bar;
  wire in_13bar;
  wire in_12bar;
  wire in_11bar;
  wire in_10bar;
  wire in_9bar;
  wire in_8bar;
  wire in_7bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_3bar;
  wire in_2bar;
  wire in_1bar;
  wire in_0bar;
  wire n487bar;
  wire n488bar;
  wire n489bar;
  wire n490bar;
  wire n491bar;
  wire n492bar;
  wire n493bar;
  wire n494bar;
  wire n495bar;
  wire n496bar;
  wire n497bar;
  wire n498bar;
  wire n499bar;
  wire n500bar;
  wire n501bar;
  wire n502bar;
  wire n503bar;
  wire n504bar;
  wire n505bar;
  wire n506bar;
  wire n507bar;
  wire n508bar;
  wire n509bar;
  wire n510bar;
  wire n511bar;
  wire n512bar;
  wire n513bar;
  wire n514bar;
  wire n515bar;
  wire n516bar;
  wire n517bar;
  wire n518bar;
  wire n519bar;
  wire n520bar;
  wire n521bar;
  wire n522bar;
  wire n523bar;
  wire n524bar;
  wire n525bar;
  wire n526bar;
  wire n527bar;
  wire n528bar;
  wire n529bar;
  wire n530bar;
  wire n531bar;
  wire n532bar;
  wire n533bar;
  wire n534bar;
  wire n535bar;
  wire n536bar;
  wire n537bar;
  wire n538bar;
  wire n539bar;
  wire n540bar;
  wire n541bar;
  wire n542bar;
  wire n543bar;
  wire n544bar;
  wire n545bar;
  wire n546bar;
  wire n547bar;
  wire n548bar;
  wire n549bar;
  wire n550bar;
  wire n551bar;
  wire n552bar;
  wire n553bar;
  wire n554bar;
  wire n555bar;
  wire n556bar;
  wire n557bar;
  wire n558bar;
  wire n559bar;
  wire n560bar;
  wire n561bar;
  wire n562bar;
  wire n563bar;
  wire n564bar;
  wire n565bar;
  wire n566bar;
  wire n567bar;
  wire n568bar;
  wire n569bar;
  wire n570bar;
  wire n571bar;
  wire n572bar;
  wire n573bar;
  wire n574bar;
  wire n575bar;
  wire n576bar;
  wire n577bar;
  wire n578bar;
  wire n579bar;
  wire n580bar;
  wire n581bar;
  wire n582bar;
  wire n583bar;
  wire n584bar;
  wire n585bar;
  wire n586bar;
  wire n587bar;
  wire n588bar;
  wire n589bar;
  wire n590bar;
  wire n591bar;
  wire n592bar;
  wire n593bar;
  wire n594bar;
  wire n595bar;
  wire n596bar;
  wire n597bar;
  wire n598bar;
  wire n599bar;
  wire n600bar;
  wire n601bar;
  wire n602bar;
  wire n603bar;
  wire n604bar;
  wire n605bar;
  wire n606bar;
  wire n607bar;
  wire n608bar;
  wire n609bar;
  wire n610bar;
  wire n611bar;
  wire n612bar;
  wire n613bar;
  wire n614bar;
  wire n615bar;
  wire n616bar;
  wire n617bar;
  wire n618bar;
  wire n619bar;
  wire n620bar;
  wire n621bar;
  wire n622bar;
  wire n623bar;
  wire n624bar;
  wire n625bar;
  wire n626bar;
  wire n627bar;
  wire n628bar;
  wire n629bar;
  wire n630bar;
  wire n631bar;
  wire n632bar;
  wire n633bar;
  wire n634bar;
  wire n635bar;
  wire n636bar;
  wire n637bar;
  wire n638bar;
  wire n639bar;
  wire n640bar;
  wire n641bar;
  wire n642bar;
  wire n643bar;
  wire n644bar;
  wire n645bar;
  wire n646bar;
  wire n647bar;
  wire n648bar;
  wire n649bar;
  wire n650bar;
  wire n651bar;
  wire n652bar;
  wire n653bar;
  wire n654bar;
  wire n655bar;
  wire n656bar;
  wire n657bar;
  wire n658bar;
  wire n659bar;
  wire n660bar;
  wire n661bar;
  wire n662bar;
  wire n663bar;
  wire n664bar;
  wire n665bar;
  wire n666bar;
  wire n667bar;
  wire n668bar;
  wire n669bar;
  wire n670bar;
  wire n671bar;
  wire n672bar;
  wire n673bar;
  wire n674bar;
  wire n675bar;
  wire n676bar;
  wire n677bar;
  wire n678bar;
  wire n679bar;
  wire n680bar;
  wire n681bar;
  wire n682bar;
  wire n683bar;
  wire n684bar;
  wire n685bar;
  wire n686bar;
  wire n687bar;
  wire n688bar;
  wire n689bar;
  wire n690bar;
  wire n691bar;
  wire n692bar;
  wire n693bar;
  wire n694bar;
  wire n695bar;
  wire n696bar;
  wire n697bar;
  wire n698bar;
  wire n699bar;
  wire n700bar;
  wire n701bar;
  wire n702bar;
  wire n703bar;
  wire n704bar;
  wire n705bar;
  wire n706bar;
  wire n707bar;
  wire n708bar;
  wire n709bar;
  wire n710bar;
  wire n711bar;
  wire n712bar;
  wire n713bar;
  wire n714bar;
  wire n715bar;
  wire n716bar;
  wire n717bar;
  wire n718bar;
  wire n719bar;
  wire n720bar;
  wire n721bar;
  wire n722bar;
  wire n723bar;
  wire n724bar;
  wire n725bar;
  wire n726bar;
  wire n727bar;
  wire n728bar;
  wire n729bar;
  wire n730bar;
  wire n731bar;
  wire n732bar;
  wire n733bar;
  wire n734bar;
  wire n735bar;
  wire n736bar;
  wire n737bar;
  wire n738bar;
  wire n739bar;
  wire n740bar;
  wire n741bar;
  wire n742bar;
  wire n743bar;
  wire n744bar;
  wire n745bar;
  wire n746bar;
  wire n747bar;
  wire n748bar;
  wire n749bar;
  wire n750bar;
  wire n751bar;
  wire n752bar;
  wire n753bar;
  wire n754bar;
  wire n755bar;
  wire n756bar;
  wire n757bar;
  wire n758bar;
  wire n759bar;
  wire n760bar;
  wire n761bar;
  wire n762bar;
  wire n763bar;
  wire n764bar;
  wire n765bar;
  wire n766bar;
  wire n767bar;
  wire n768bar;
  wire n769bar;
  wire n770bar;
  wire n771bar;
  wire n772bar;
  wire n773bar;
  wire n774bar;
  wire n775bar;
  wire n776bar;
  wire n777bar;
  wire n778bar;
  wire n779bar;
  wire n780bar;
  wire n781bar;
  wire n782bar;
  wire n783bar;
  wire n784bar;
  wire n785bar;
  wire n786bar;
  wire n787bar;
  wire n788bar;
  wire n789bar;
  wire n790bar;
  wire n791bar;
  wire n792bar;
  wire n793bar;
  wire n794bar;
  wire n795bar;
  wire n796bar;
  wire n797bar;
  wire n798bar;
  wire n799bar;
  wire n800bar;
  wire n801bar;
  wire n802bar;
  wire n803bar;
  wire n804bar;
  wire n805bar;
  wire n806bar;
  wire n807bar;
  wire n808bar;
  wire n809bar;
  wire n810bar;
  wire n811bar;
  wire n812bar;
  wire n813bar;
  wire n814bar;
  wire n815bar;
  wire n816bar;
  wire n817bar;
  wire n818bar;
  wire n819bar;
  wire n820bar;
  wire n821bar;
  wire n822bar;
  wire n823bar;
  wire n824bar;
  wire n825bar;
  wire n826bar;
  wire n827bar;
  wire n828bar;
  wire n829bar;
  wire n830bar;
  wire n831bar;
  wire n832bar;
  wire n833bar;
  wire n834bar;
  wire n835bar;
  wire n836bar;
  wire n837bar;
  wire n838bar;
  wire n839bar;
  wire n840bar;
  wire n841bar;
  wire n842bar;
  wire n843bar;
  wire n844bar;
  wire n845bar;
  wire n846bar;
  wire n847bar;
  wire n848bar;
  wire n849bar;
  wire n850bar;
  wire n851bar;
  wire n852bar;
  wire n853bar;
  wire n854bar;
  wire n855bar;
  wire n856bar;
  wire n857bar;
  wire n858bar;
  wire n859bar;
  wire n860bar;
  wire n861bar;
  wire n862bar;
  wire n863bar;
  wire n864bar;
  wire n865bar;
  wire n866bar;
  wire n867bar;
  wire n868bar;
  wire n869bar;
  wire n870bar;
  wire n871bar;
  wire n872bar;
  wire n873bar;
  wire n874bar;
  wire n875bar;
  wire n876bar;
  wire n877bar;
  wire n878bar;
  wire n879bar;
  wire n880bar;
  wire n881bar;
  wire n882bar;
  wire n883bar;
  wire n884bar;
  wire n885bar;
  wire n886bar;
  wire n887bar;
  wire n888bar;
  wire n889bar;
  wire n890bar;
  wire n891bar;
  wire n892bar;
  wire n893bar;
  wire n894bar;
  wire n895bar;
  wire n896bar;
  wire n897bar;
  wire n898bar;
  wire n899bar;
  wire n900bar;
  wire n901bar;
  wire n902bar;
  wire n903bar;
  wire n904bar;
  wire n905bar;
  wire n906bar;
  wire n907bar;
  wire n908bar;
  wire n909bar;
  wire n910bar;
  wire n911bar;
  wire n912bar;
  wire n913bar;
  wire n914bar;
  wire n915bar;
  wire n916bar;
  wire n917bar;
  wire n918bar;
  wire n919bar;
  wire n920bar;
  wire n921bar;
  wire n922bar;
  wire n923bar;
  wire n924bar;
  wire n925bar;
  wire n926bar;
  wire n927bar;
  wire n928bar;
  wire n929bar;
  wire n930bar;
  wire n931bar;
  wire n932bar;
  wire n933bar;
  wire n934bar;
  wire n935bar;
  wire n936bar;
  wire n937bar;
  wire n938bar;
  wire n939bar;
  wire n940bar;
  wire n941bar;
  wire n942bar;
  wire n943bar;
  wire n944bar;
  wire n945bar;
  wire n946bar;
  wire n947bar;
  wire n948bar;
  wire n949bar;
  wire n950bar;
  wire n951bar;
  wire n952bar;
  wire n953bar;
  wire n954bar;
  wire n955bar;
  wire n956bar;
  wire n957bar;
  wire n958bar;
  wire n959bar;
  wire n960bar;
  wire n961bar;
  wire n962bar;
  wire n963bar;
  wire n964bar;
  wire n965bar;
  wire n966bar;
  wire n967bar;
  wire n968bar;
  wire n969bar;
  wire n970bar;
  wire n971bar;
  wire n972bar;
//wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];
  assign in_81bar = inbar[81];
  assign in_80bar = inbar[80];
  assign in_79bar = inbar[79];
  assign in_78bar = inbar[78];
  assign in_77bar = inbar[77];
  assign in_76bar = inbar[76];
  assign in_75bar = inbar[75];
  assign in_74bar = inbar[74];
  assign in_73bar = inbar[73];
  assign in_72bar = inbar[72];
  assign in_71bar = inbar[71];
  assign in_70bar = inbar[70];
  assign in_69bar = inbar[69];
  assign in_68bar = inbar[68];
  assign in_67bar = inbar[67];
  assign in_66bar = inbar[66];
  assign in_65bar = inbar[65];
  assign in_64bar = inbar[64];
  assign in_63bar = inbar[63];
  assign in_62bar = inbar[62];
  assign in_61bar = inbar[61];
  assign in_60bar = inbar[60];
  assign in_59bar = inbar[59];
  assign in_58bar = inbar[58];
  assign in_57bar = inbar[57];
  assign in_56bar = inbar[56];
  assign in_55bar = inbar[55];
  assign in_54bar = inbar[54];
  assign in_53bar = inbar[53];
  assign in_52bar = inbar[52];
  assign in_51bar = inbar[51];
  assign in_50bar = inbar[50];
  assign in_49bar = inbar[49];
  assign in_48bar = inbar[48];
  assign in_47bar = inbar[47];
  assign in_46bar = inbar[46];
  assign in_45bar = inbar[45];
  assign in_44bar = inbar[44];
  assign in_43bar = inbar[43];
  assign in_42bar = inbar[42];
  assign in_41bar = inbar[41];
  assign in_40bar = inbar[40];
  assign in_39bar = inbar[39];
  assign in_38bar = inbar[38];
  assign in_37bar = inbar[37];
  assign in_36bar = inbar[36];
  assign in_35bar = inbar[35];
  assign in_34bar = inbar[34];
  assign in_33bar = inbar[33];
  assign in_32bar = inbar[32];
  assign in_31bar = inbar[31];
  assign in_30bar = inbar[30];
  assign in_29bar = inbar[29];
  assign in_28bar = inbar[28];
  assign in_27bar = inbar[27];
  assign in_26bar = inbar[26];
  assign in_25bar = inbar[25];
  assign in_24bar = inbar[24];
  assign in_23bar = inbar[23];
  assign in_22bar = inbar[22];
  assign in_21bar = inbar[21];
  assign in_20bar = inbar[20];
  assign in_19bar = inbar[19];
  assign in_18bar = inbar[18];
  assign in_17bar = inbar[17];
  assign in_16bar = inbar[16];
  assign in_15bar = inbar[15];
  assign in_14bar = inbar[14];
  assign in_13bar = inbar[13];
  assign in_12bar = inbar[12];
  assign in_11bar = inbar[11];
  assign in_10bar = inbar[10];
  assign in_9bar = inbar[9];
  assign in_8bar = inbar[8];
  assign in_7bar = inbar[7];
  assign in_6bar = inbar[6];
  assign in_5bar = inbar[5];
  assign in_4bar = inbar[4];
  assign in_3bar = inbar[3];
  assign in_2bar = inbar[2];
  assign in_1bar = inbar[1];
  assign in_0bar = inbar[0];
//assign_done

  OR2_X1 U1 ( .A1(n972), .A2(n971), .ZN(out[7]) );
  AND2_X1 U1bar ( .A1(n972bar), .A2(n971bar), .ZN(outbar[7]) );
  OR2_X1 U2 ( .A1(n970), .A2(n969), .ZN(n971) );
  AND2_X1 U2bar ( .A1(n970bar), .A2(n969bar), .ZN(n971bar) );
  OR2_X1 U3 ( .A1(n968), .A2(n967), .ZN(n969) );
  AND2_X1 U3bar ( .A1(n968bar), .A2(n967bar), .ZN(n969bar) );
  OR2_X1 U4 ( .A1(n966), .A2(n965), .ZN(n967) );
  AND2_X1 U4bar ( .A1(n966bar), .A2(n965bar), .ZN(n967bar) );
  OR2_X1 U5 ( .A1(n964), .A2(n963), .ZN(n968) );
  AND2_X1 U5bar ( .A1(n964bar), .A2(n963bar), .ZN(n968bar) );
  OR2_X1 U6 ( .A1(in[116]), .A2(n962), .ZN(n963) );
  AND2_X1 U6bar ( .A1(inbar[116]), .A2(n962bar), .ZN(n963bar) );
  OR2_X1 U7 ( .A1(n961), .A2(n960), .ZN(n970) );
  AND2_X1 U7bar ( .A1(n961bar), .A2(n960bar), .ZN(n970bar) );
  OR2_X1 U8 ( .A1(in[150]), .A2(in[127]), .ZN(n960) );
  AND2_X1 U8bar ( .A1(inbar[150]), .A2(inbar[127]), .ZN(n960bar) );
  OR2_X1 U9 ( .A1(in[160]), .A2(n959), .ZN(n961) );
  AND2_X1 U9bar ( .A1(inbar[160]), .A2(n959bar), .ZN(n961bar) );
  OR2_X1 U10 ( .A1(in[252]), .A2(in[168]), .ZN(n959) );
  AND2_X1 U10bar ( .A1(inbar[252]), .A2(inbar[168]), .ZN(n959bar) );
  OR2_X1 U11 ( .A1(n958), .A2(n957), .ZN(n972) );
  AND2_X1 U11bar ( .A1(n958bar), .A2(n957bar), .ZN(n972bar) );
  OR2_X1 U12 ( .A1(n956), .A2(n955), .ZN(n957) );
  AND2_X1 U12bar ( .A1(n956bar), .A2(n955bar), .ZN(n957bar) );
  OR2_X1 U13 ( .A1(in_17), .A2(in[96]), .ZN(n955) );
  AND2_X1 U13bar ( .A1(in_17bar), .A2(inbar[96]), .ZN(n955bar) );
  OR2_X1 U14 ( .A1(in_23), .A2(n954), .ZN(n956) );
  AND2_X1 U14bar ( .A1(in_23bar), .A2(n954bar), .ZN(n956bar) );
  OR2_X1 U15 ( .A1(in_31), .A2(in_26), .ZN(n954) );
  AND2_X1 U15bar ( .A1(in_31bar), .A2(in_26bar), .ZN(n954bar) );
  OR2_X1 U16 ( .A1(n953), .A2(n952), .ZN(n958) );
  AND2_X1 U16bar ( .A1(n953bar), .A2(n952bar), .ZN(n958bar) );
  OR2_X1 U17 ( .A1(in_58), .A2(in_4), .ZN(n952) );
  AND2_X1 U17bar ( .A1(in_58bar), .A2(in_4bar), .ZN(n952bar) );
  OR2_X1 U18 ( .A1(in_59), .A2(n951), .ZN(n953) );
  AND2_X1 U18bar ( .A1(in_59bar), .A2(n951bar), .ZN(n953bar) );
  OR2_X1 U19 ( .A1(in_71), .A2(in_62), .ZN(n951) );
  AND2_X1 U19bar ( .A1(in_71bar), .A2(in_62bar), .ZN(n951bar) );
  OR2_X1 U20 ( .A1(n950), .A2(n949), .ZN(out[6]) );
  AND2_X1 U20bar ( .A1(n950bar), .A2(n949bar), .ZN(outbar[6]) );
  OR2_X1 U21 ( .A1(n948), .A2(n947), .ZN(n949) );
  AND2_X1 U21bar ( .A1(n948bar), .A2(n947bar), .ZN(n949bar) );
  OR2_X1 U22 ( .A1(n946), .A2(n945), .ZN(n947) );
  AND2_X1 U22bar ( .A1(n946bar), .A2(n945bar), .ZN(n947bar) );
  OR2_X1 U23 ( .A1(n944), .A2(n943), .ZN(n945) );
  AND2_X1 U23bar ( .A1(n944bar), .A2(n943bar), .ZN(n945bar) );
  OR2_X1 U24 ( .A1(n942), .A2(n941), .ZN(n946) );
  AND2_X1 U24bar ( .A1(n942bar), .A2(n941bar), .ZN(n946bar) );
  OR2_X1 U25 ( .A1(in[101]), .A2(n940), .ZN(n941) );
  AND2_X1 U25bar ( .A1(inbar[101]), .A2(n940bar), .ZN(n941bar) );
  OR2_X1 U26 ( .A1(n939), .A2(n938), .ZN(n948) );
  AND2_X1 U26bar ( .A1(n939bar), .A2(n938bar), .ZN(n948bar) );
  OR2_X1 U27 ( .A1(in[114]), .A2(in[104]), .ZN(n938) );
  AND2_X1 U27bar ( .A1(inbar[114]), .A2(inbar[104]), .ZN(n938bar) );
  OR2_X1 U28 ( .A1(in[128]), .A2(n937), .ZN(n939) );
  AND2_X1 U28bar ( .A1(inbar[128]), .A2(n937bar), .ZN(n939bar) );
  OR2_X1 U29 ( .A1(in[136]), .A2(in[134]), .ZN(n937) );
  AND2_X1 U29bar ( .A1(inbar[136]), .A2(inbar[134]), .ZN(n937bar) );
  OR2_X1 U30 ( .A1(n936), .A2(n935), .ZN(n950) );
  AND2_X1 U30bar ( .A1(n936bar), .A2(n935bar), .ZN(n950bar) );
  OR2_X1 U31 ( .A1(n934), .A2(n933), .ZN(n935) );
  AND2_X1 U31bar ( .A1(n934bar), .A2(n933bar), .ZN(n935bar) );
  OR2_X1 U32 ( .A1(in[177]), .A2(in[164]), .ZN(n933) );
  AND2_X1 U32bar ( .A1(inbar[177]), .A2(inbar[164]), .ZN(n933bar) );
  OR2_X1 U33 ( .A1(in[212]), .A2(n932), .ZN(n934) );
  AND2_X1 U33bar ( .A1(inbar[212]), .A2(n932bar), .ZN(n934bar) );
  OR2_X1 U34 ( .A1(in[248]), .A2(in[221]), .ZN(n932) );
  AND2_X1 U34bar ( .A1(inbar[248]), .A2(inbar[221]), .ZN(n932bar) );
  OR2_X1 U35 ( .A1(n931), .A2(n930), .ZN(n936) );
  AND2_X1 U35bar ( .A1(n931bar), .A2(n930bar), .ZN(n936bar) );
  OR2_X1 U36 ( .A1(in_18), .A2(in[93]), .ZN(n930) );
  AND2_X1 U36bar ( .A1(in_18bar), .A2(inbar[93]), .ZN(n930bar) );
  OR2_X1 U37 ( .A1(in_31), .A2(n929), .ZN(n931) );
  AND2_X1 U37bar ( .A1(in_31bar), .A2(n929bar), .ZN(n931bar) );
  OR2_X1 U38 ( .A1(in_7), .A2(in_39), .ZN(n929) );
  AND2_X1 U38bar ( .A1(in_7bar), .A2(in_39bar), .ZN(n929bar) );
  OR2_X1 U39 ( .A1(n928), .A2(n927), .ZN(out[5]) );
  AND2_X1 U39bar ( .A1(n928bar), .A2(n927bar), .ZN(outbar[5]) );
  OR2_X1 U40 ( .A1(n926), .A2(n925), .ZN(n927) );
  AND2_X1 U40bar ( .A1(n926bar), .A2(n925bar), .ZN(n927bar) );
  OR2_X1 U41 ( .A1(n924), .A2(n923), .ZN(n925) );
  AND2_X1 U41bar ( .A1(n924bar), .A2(n923bar), .ZN(n925bar) );
  OR2_X1 U42 ( .A1(n922), .A2(n921), .ZN(n923) );
  AND2_X1 U42bar ( .A1(n922bar), .A2(n921bar), .ZN(n923bar) );
  OR2_X1 U43 ( .A1(n940), .A2(n920), .ZN(n924) );
  AND2_X1 U43bar ( .A1(n940bar), .A2(n920bar), .ZN(n924bar) );
  OR2_X1 U44 ( .A1(in[111]), .A2(n919), .ZN(n920) );
  AND2_X1 U44bar ( .A1(inbar[111]), .A2(n919bar), .ZN(n920bar) );
  OR2_X1 U45 ( .A1(n918), .A2(n917), .ZN(n940) );
  AND2_X1 U45bar ( .A1(n918bar), .A2(n917bar), .ZN(n940bar) );
  OR2_X1 U46 ( .A1(n916), .A2(n915), .ZN(n917) );
  AND2_X1 U46bar ( .A1(n916bar), .A2(n915bar), .ZN(n917bar) );
  OR2_X1 U47 ( .A1(n914), .A2(n913), .ZN(n915) );
  AND2_X1 U47bar ( .A1(n914bar), .A2(n913bar), .ZN(n915bar) );
  OR2_X1 U48 ( .A1(in[140]), .A2(in[131]), .ZN(n913) );
  AND2_X1 U48bar ( .A1(inbar[140]), .A2(inbar[131]), .ZN(n913bar) );
  OR2_X1 U49 ( .A1(in[160]), .A2(in[144]), .ZN(n914) );
  AND2_X1 U49bar ( .A1(inbar[160]), .A2(inbar[144]), .ZN(n914bar) );
  OR2_X1 U50 ( .A1(n912), .A2(n911), .ZN(n916) );
  AND2_X1 U50bar ( .A1(n912bar), .A2(n911bar), .ZN(n916bar) );
  OR2_X1 U51 ( .A1(in[179]), .A2(in[174]), .ZN(n911) );
  AND2_X1 U51bar ( .A1(inbar[179]), .A2(inbar[174]), .ZN(n911bar) );
  OR2_X1 U52 ( .A1(in[188]), .A2(in[184]), .ZN(n912) );
  AND2_X1 U52bar ( .A1(inbar[188]), .A2(inbar[184]), .ZN(n912bar) );
  OR2_X1 U53 ( .A1(n910), .A2(n909), .ZN(n918) );
  AND2_X1 U53bar ( .A1(n910bar), .A2(n909bar), .ZN(n918bar) );
  OR2_X1 U54 ( .A1(n908), .A2(n907), .ZN(n909) );
  AND2_X1 U54bar ( .A1(n908bar), .A2(n907bar), .ZN(n909bar) );
  OR2_X1 U55 ( .A1(in[216]), .A2(in[200]), .ZN(n907) );
  AND2_X1 U55bar ( .A1(inbar[216]), .A2(inbar[200]), .ZN(n907bar) );
  OR2_X1 U56 ( .A1(in[228]), .A2(in[224]), .ZN(n908) );
  AND2_X1 U56bar ( .A1(inbar[228]), .A2(inbar[224]), .ZN(n908bar) );
  OR2_X1 U57 ( .A1(n906), .A2(n905), .ZN(n910) );
  AND2_X1 U57bar ( .A1(n906bar), .A2(n905bar), .ZN(n910bar) );
  OR2_X1 U58 ( .A1(in[247]), .A2(in[235]), .ZN(n905) );
  AND2_X1 U58bar ( .A1(inbar[247]), .A2(inbar[235]), .ZN(n905bar) );
  OR2_X1 U59 ( .A1(in_42), .A2(in[83]), .ZN(n906) );
  AND2_X1 U59bar ( .A1(in_42bar), .A2(inbar[83]), .ZN(n906bar) );
  OR2_X1 U60 ( .A1(n904), .A2(n903), .ZN(n926) );
  AND2_X1 U60bar ( .A1(n904bar), .A2(n903bar), .ZN(n926bar) );
  OR2_X1 U61 ( .A1(in[166]), .A2(in[123]), .ZN(n903) );
  AND2_X1 U61bar ( .A1(inbar[166]), .A2(inbar[123]), .ZN(n903bar) );
  OR2_X1 U62 ( .A1(in[170]), .A2(n902), .ZN(n904) );
  AND2_X1 U62bar ( .A1(inbar[170]), .A2(n902bar), .ZN(n904bar) );
  OR2_X1 U63 ( .A1(in[194]), .A2(in[183]), .ZN(n902) );
  AND2_X1 U63bar ( .A1(inbar[194]), .A2(inbar[183]), .ZN(n902bar) );
  OR2_X1 U64 ( .A1(n901), .A2(n900), .ZN(n928) );
  AND2_X1 U64bar ( .A1(n901bar), .A2(n900bar), .ZN(n928bar) );
  OR2_X1 U65 ( .A1(n899), .A2(n898), .ZN(n900) );
  AND2_X1 U65bar ( .A1(n899bar), .A2(n898bar), .ZN(n900bar) );
  OR2_X1 U66 ( .A1(in[241]), .A2(in[238]), .ZN(n898) );
  AND2_X1 U66bar ( .A1(inbar[241]), .A2(inbar[238]), .ZN(n898bar) );
  OR2_X1 U67 ( .A1(in[250]), .A2(n897), .ZN(n899) );
  AND2_X1 U67bar ( .A1(inbar[250]), .A2(n897bar), .ZN(n899bar) );
  OR2_X1 U68 ( .A1(in_24), .A2(in[84]), .ZN(n897) );
  AND2_X1 U68bar ( .A1(in_24bar), .A2(inbar[84]), .ZN(n897bar) );
  OR2_X1 U69 ( .A1(n896), .A2(n895), .ZN(n901) );
  AND2_X1 U69bar ( .A1(n896bar), .A2(n895bar), .ZN(n901bar) );
  OR2_X1 U70 ( .A1(in_41), .A2(in_29), .ZN(n895) );
  AND2_X1 U70bar ( .A1(in_41bar), .A2(in_29bar), .ZN(n895bar) );
  OR2_X1 U71 ( .A1(in_66), .A2(n894), .ZN(n896) );
  AND2_X1 U71bar ( .A1(in_66bar), .A2(n894bar), .ZN(n896bar) );
  OR2_X1 U72 ( .A1(in_76), .A2(in_71), .ZN(n894) );
  AND2_X1 U72bar ( .A1(in_76bar), .A2(in_71bar), .ZN(n894bar) );
  OR2_X1 U73 ( .A1(n893), .A2(n892), .ZN(out[4]) );
  AND2_X1 U73bar ( .A1(n893bar), .A2(n892bar), .ZN(outbar[4]) );
  OR2_X1 U74 ( .A1(n891), .A2(n890), .ZN(n892) );
  AND2_X1 U74bar ( .A1(n891bar), .A2(n890bar), .ZN(n892bar) );
  OR2_X1 U75 ( .A1(n889), .A2(n888), .ZN(n890) );
  AND2_X1 U75bar ( .A1(n889bar), .A2(n888bar), .ZN(n890bar) );
  OR2_X1 U76 ( .A1(n922), .A2(n887), .ZN(n888) );
  AND2_X1 U76bar ( .A1(n922bar), .A2(n887bar), .ZN(n888bar) );
  OR2_X1 U77 ( .A1(n886), .A2(n885), .ZN(n922) );
  AND2_X1 U77bar ( .A1(n886bar), .A2(n885bar), .ZN(n922bar) );
  OR2_X1 U78 ( .A1(n884), .A2(n883), .ZN(n885) );
  AND2_X1 U78bar ( .A1(n884bar), .A2(n883bar), .ZN(n885bar) );
  OR2_X1 U79 ( .A1(n882), .A2(n881), .ZN(n883) );
  AND2_X1 U79bar ( .A1(n882bar), .A2(n881bar), .ZN(n883bar) );
  OR2_X1 U80 ( .A1(in[118]), .A2(in[109]), .ZN(n881) );
  AND2_X1 U80bar ( .A1(inbar[118]), .A2(inbar[109]), .ZN(n881bar) );
  OR2_X1 U81 ( .A1(in[139]), .A2(in[120]), .ZN(n882) );
  AND2_X1 U81bar ( .A1(inbar[139]), .A2(inbar[120]), .ZN(n882bar) );
  OR2_X1 U82 ( .A1(n880), .A2(n879), .ZN(n884) );
  AND2_X1 U82bar ( .A1(n880bar), .A2(n879bar), .ZN(n884bar) );
  OR2_X1 U83 ( .A1(in[198]), .A2(in[154]), .ZN(n879) );
  AND2_X1 U83bar ( .A1(inbar[198]), .A2(inbar[154]), .ZN(n879bar) );
  OR2_X1 U84 ( .A1(in[210]), .A2(in[205]), .ZN(n880) );
  AND2_X1 U84bar ( .A1(inbar[210]), .A2(inbar[205]), .ZN(n880bar) );
  OR2_X1 U85 ( .A1(n878), .A2(n877), .ZN(n886) );
  AND2_X1 U85bar ( .A1(n878bar), .A2(n877bar), .ZN(n886bar) );
  OR2_X1 U86 ( .A1(n876), .A2(n875), .ZN(n877) );
  AND2_X1 U86bar ( .A1(n876bar), .A2(n875bar), .ZN(n877bar) );
  OR2_X1 U87 ( .A1(in[219]), .A2(in[217]), .ZN(n875) );
  AND2_X1 U87bar ( .A1(inbar[219]), .A2(inbar[217]), .ZN(n875bar) );
  OR2_X1 U88 ( .A1(in[86]), .A2(in[252]), .ZN(n876) );
  AND2_X1 U88bar ( .A1(inbar[86]), .A2(inbar[252]), .ZN(n876bar) );
  OR2_X1 U89 ( .A1(n874), .A2(n873), .ZN(n878) );
  AND2_X1 U89bar ( .A1(n874bar), .A2(n873bar), .ZN(n878bar) );
  OR2_X1 U90 ( .A1(in_40), .A2(in[91]), .ZN(n873) );
  AND2_X1 U90bar ( .A1(in_40bar), .A2(inbar[91]), .ZN(n873bar) );
  OR2_X1 U91 ( .A1(in_8), .A2(in_46), .ZN(n874) );
  AND2_X1 U91bar ( .A1(in_8bar), .A2(in_46bar), .ZN(n874bar) );
  OR2_X1 U92 ( .A1(n872), .A2(n871), .ZN(n889) );
  AND2_X1 U92bar ( .A1(n872bar), .A2(n871bar), .ZN(n889bar) );
  OR2_X1 U93 ( .A1(in[117]), .A2(n943), .ZN(n871) );
  AND2_X1 U93bar ( .A1(inbar[117]), .A2(n943bar), .ZN(n871bar) );
  OR2_X1 U94 ( .A1(n870), .A2(n869), .ZN(n943) );
  AND2_X1 U94bar ( .A1(n870bar), .A2(n869bar), .ZN(n943bar) );
  OR2_X1 U95 ( .A1(n868), .A2(n867), .ZN(n869) );
  AND2_X1 U95bar ( .A1(n868bar), .A2(n867bar), .ZN(n869bar) );
  OR2_X1 U96 ( .A1(n866), .A2(n865), .ZN(n867) );
  AND2_X1 U96bar ( .A1(n866bar), .A2(n865bar), .ZN(n867bar) );
  OR2_X1 U97 ( .A1(n864), .A2(n863), .ZN(n865) );
  AND2_X1 U97bar ( .A1(n864bar), .A2(n863bar), .ZN(n865bar) );
  OR2_X1 U98 ( .A1(in[108]), .A2(n919), .ZN(n866) );
  AND2_X1 U98bar ( .A1(inbar[108]), .A2(n919bar), .ZN(n866bar) );
  OR2_X1 U99 ( .A1(n862), .A2(n861), .ZN(n919) );
  AND2_X1 U99bar ( .A1(n862bar), .A2(n861bar), .ZN(n919bar) );
  OR2_X1 U100 ( .A1(n860), .A2(n859), .ZN(n861) );
  AND2_X1 U100bar ( .A1(n860bar), .A2(n859bar), .ZN(n861bar) );
  OR2_X1 U101 ( .A1(n858), .A2(n857), .ZN(n859) );
  AND2_X1 U101bar ( .A1(n858bar), .A2(n857bar), .ZN(n859bar) );
  OR2_X1 U102 ( .A1(in[119]), .A2(in[105]), .ZN(n857) );
  AND2_X1 U102bar ( .A1(inbar[119]), .A2(inbar[105]), .ZN(n857bar) );
  OR2_X1 U103 ( .A1(in[186]), .A2(in[175]), .ZN(n858) );
  AND2_X1 U103bar ( .A1(inbar[186]), .A2(inbar[175]), .ZN(n858bar) );
  OR2_X1 U104 ( .A1(n856), .A2(n855), .ZN(n860) );
  AND2_X1 U104bar ( .A1(n856bar), .A2(n855bar), .ZN(n860bar) );
  OR2_X1 U105 ( .A1(in[202]), .A2(in[193]), .ZN(n855) );
  AND2_X1 U105bar ( .A1(inbar[202]), .A2(inbar[193]), .ZN(n855bar) );
  OR2_X1 U106 ( .A1(in[225]), .A2(in[208]), .ZN(n856) );
  AND2_X1 U106bar ( .A1(inbar[225]), .A2(inbar[208]), .ZN(n856bar) );
  OR2_X1 U107 ( .A1(n854), .A2(n853), .ZN(n862) );
  AND2_X1 U107bar ( .A1(n854bar), .A2(n853bar), .ZN(n862bar) );
  OR2_X1 U108 ( .A1(n852), .A2(n851), .ZN(n853) );
  AND2_X1 U108bar ( .A1(n852bar), .A2(n851bar), .ZN(n853bar) );
  OR2_X1 U109 ( .A1(in_1), .A2(in[85]), .ZN(n851) );
  AND2_X1 U109bar ( .A1(in_1bar), .A2(inbar[85]), .ZN(n851bar) );
  OR2_X1 U110 ( .A1(in_23), .A2(in_19), .ZN(n852) );
  AND2_X1 U110bar ( .A1(in_23bar), .A2(in_19bar), .ZN(n852bar) );
  OR2_X1 U111 ( .A1(n850), .A2(n849), .ZN(n854) );
  AND2_X1 U111bar ( .A1(n850bar), .A2(n849bar), .ZN(n854bar) );
  OR2_X1 U112 ( .A1(in_43), .A2(in_33), .ZN(n849) );
  AND2_X1 U112bar ( .A1(in_43bar), .A2(in_33bar), .ZN(n849bar) );
  OR2_X1 U113 ( .A1(in_63), .A2(in_44), .ZN(n850) );
  AND2_X1 U113bar ( .A1(in_63bar), .A2(in_44bar), .ZN(n850bar) );
  OR2_X1 U114 ( .A1(n848), .A2(n847), .ZN(n868) );
  AND2_X1 U114bar ( .A1(n848bar), .A2(n847bar), .ZN(n868bar) );
  OR2_X1 U115 ( .A1(in[141]), .A2(in[112]), .ZN(n847) );
  AND2_X1 U115bar ( .A1(inbar[141]), .A2(inbar[112]), .ZN(n847bar) );
  OR2_X1 U116 ( .A1(in[147]), .A2(n846), .ZN(n848) );
  AND2_X1 U116bar ( .A1(inbar[147]), .A2(n846bar), .ZN(n848bar) );
  OR2_X1 U117 ( .A1(in[181]), .A2(in[167]), .ZN(n846) );
  AND2_X1 U117bar ( .A1(inbar[181]), .A2(inbar[167]), .ZN(n846bar) );
  OR2_X1 U118 ( .A1(n845), .A2(n844), .ZN(n870) );
  AND2_X1 U118bar ( .A1(n845bar), .A2(n844bar), .ZN(n870bar) );
  OR2_X1 U119 ( .A1(n843), .A2(n842), .ZN(n844) );
  AND2_X1 U119bar ( .A1(n843bar), .A2(n842bar), .ZN(n844bar) );
  OR2_X1 U120 ( .A1(in[229]), .A2(in[201]), .ZN(n842) );
  AND2_X1 U120bar ( .A1(inbar[229]), .A2(inbar[201]), .ZN(n842bar) );
  OR2_X1 U121 ( .A1(in[237]), .A2(n841), .ZN(n843) );
  AND2_X1 U121bar ( .A1(inbar[237]), .A2(n841bar), .ZN(n843bar) );
  OR2_X1 U122 ( .A1(in[94]), .A2(in[253]), .ZN(n841) );
  AND2_X1 U122bar ( .A1(inbar[94]), .A2(inbar[253]), .ZN(n841bar) );
  OR2_X1 U123 ( .A1(n840), .A2(n839), .ZN(n845) );
  AND2_X1 U123bar ( .A1(n840bar), .A2(n839bar), .ZN(n845bar) );
  OR2_X1 U124 ( .A1(in_21), .A2(in[96]), .ZN(n839) );
  AND2_X1 U124bar ( .A1(in_21bar), .A2(inbar[96]), .ZN(n839bar) );
  OR2_X1 U125 ( .A1(in_25), .A2(n838), .ZN(n840) );
  AND2_X1 U125bar ( .A1(in_25bar), .A2(n838bar), .ZN(n840bar) );
  OR2_X1 U126 ( .A1(in_81), .A2(in_45), .ZN(n838) );
  AND2_X1 U126bar ( .A1(in_81bar), .A2(in_45bar), .ZN(n838bar) );
  OR2_X1 U127 ( .A1(n837), .A2(n836), .ZN(n891) );
  AND2_X1 U127bar ( .A1(n837bar), .A2(n836bar), .ZN(n891bar) );
  OR2_X1 U128 ( .A1(in[142]), .A2(in[124]), .ZN(n836) );
  AND2_X1 U128bar ( .A1(inbar[142]), .A2(inbar[124]), .ZN(n836bar) );
  OR2_X1 U129 ( .A1(in[150]), .A2(n835), .ZN(n837) );
  AND2_X1 U129bar ( .A1(inbar[150]), .A2(n835bar), .ZN(n837bar) );
  OR2_X1 U130 ( .A1(in[172]), .A2(in[155]), .ZN(n835) );
  AND2_X1 U130bar ( .A1(inbar[172]), .A2(inbar[155]), .ZN(n835bar) );
  OR2_X1 U131 ( .A1(n834), .A2(n833), .ZN(n893) );
  AND2_X1 U131bar ( .A1(n834bar), .A2(n833bar), .ZN(n893bar) );
  OR2_X1 U132 ( .A1(n832), .A2(n831), .ZN(n833) );
  AND2_X1 U132bar ( .A1(n832bar), .A2(n831bar), .ZN(n833bar) );
  OR2_X1 U133 ( .A1(in[196]), .A2(in[173]), .ZN(n831) );
  AND2_X1 U133bar ( .A1(inbar[196]), .A2(inbar[173]), .ZN(n831bar) );
  OR2_X1 U134 ( .A1(in[222]), .A2(n830), .ZN(n832) );
  AND2_X1 U134bar ( .A1(inbar[222]), .A2(n830bar), .ZN(n832bar) );
  OR2_X1 U135 ( .A1(in[227]), .A2(in[226]), .ZN(n830) );
  AND2_X1 U135bar ( .A1(inbar[227]), .A2(inbar[226]), .ZN(n830bar) );
  OR2_X1 U136 ( .A1(n829), .A2(n828), .ZN(n834) );
  AND2_X1 U136bar ( .A1(n829bar), .A2(n828bar), .ZN(n834bar) );
  OR2_X1 U137 ( .A1(in[249]), .A2(in[231]), .ZN(n828) );
  AND2_X1 U137bar ( .A1(inbar[249]), .A2(inbar[231]), .ZN(n828bar) );
  OR2_X1 U138 ( .A1(in_28), .A2(n827), .ZN(n829) );
  AND2_X1 U138bar ( .A1(in_28bar), .A2(n827bar), .ZN(n829bar) );
  OR2_X1 U139 ( .A1(in_52), .A2(in_47), .ZN(n827) );
  AND2_X1 U139bar ( .A1(in_52bar), .A2(in_47bar), .ZN(n827bar) );
  OR2_X1 U140 ( .A1(n826), .A2(n825), .ZN(out[3]) );
  AND2_X1 U140bar ( .A1(n826bar), .A2(n825bar), .ZN(outbar[3]) );
  OR2_X1 U141 ( .A1(n824), .A2(n823), .ZN(n825) );
  AND2_X1 U141bar ( .A1(n824bar), .A2(n823bar), .ZN(n825bar) );
  OR2_X1 U142 ( .A1(n822), .A2(n821), .ZN(n823) );
  AND2_X1 U142bar ( .A1(n822bar), .A2(n821bar), .ZN(n823bar) );
  OR2_X1 U143 ( .A1(n820), .A2(n819), .ZN(n821) );
  AND2_X1 U143bar ( .A1(n820bar), .A2(n819bar), .ZN(n821bar) );
  OR2_X1 U144 ( .A1(n964), .A2(n818), .ZN(n822) );
  AND2_X1 U144bar ( .A1(n964bar), .A2(n818bar), .ZN(n822bar) );
  OR2_X1 U145 ( .A1(in[118]), .A2(n817), .ZN(n818) );
  AND2_X1 U145bar ( .A1(inbar[118]), .A2(n817bar), .ZN(n818bar) );
  OR2_X1 U146 ( .A1(n816), .A2(n815), .ZN(n964) );
  AND2_X1 U146bar ( .A1(n816bar), .A2(n815bar), .ZN(n964bar) );
  OR2_X1 U147 ( .A1(n814), .A2(n813), .ZN(n815) );
  AND2_X1 U147bar ( .A1(n814bar), .A2(n813bar), .ZN(n815bar) );
  OR2_X1 U148 ( .A1(n812), .A2(n811), .ZN(n813) );
  AND2_X1 U148bar ( .A1(n812bar), .A2(n811bar), .ZN(n813bar) );
  OR2_X1 U149 ( .A1(in[122]), .A2(in[111]), .ZN(n811) );
  AND2_X1 U149bar ( .A1(inbar[122]), .A2(inbar[111]), .ZN(n811bar) );
  OR2_X1 U150 ( .A1(in[154]), .A2(in[151]), .ZN(n812) );
  AND2_X1 U150bar ( .A1(inbar[154]), .A2(inbar[151]), .ZN(n812bar) );
  OR2_X1 U151 ( .A1(n810), .A2(n809), .ZN(n814) );
  AND2_X1 U151bar ( .A1(n810bar), .A2(n809bar), .ZN(n814bar) );
  OR2_X1 U152 ( .A1(in[187]), .A2(in[177]), .ZN(n809) );
  AND2_X1 U152bar ( .A1(inbar[187]), .A2(inbar[177]), .ZN(n809bar) );
  OR2_X1 U153 ( .A1(in[200]), .A2(in[192]), .ZN(n810) );
  AND2_X1 U153bar ( .A1(inbar[200]), .A2(inbar[192]), .ZN(n810bar) );
  OR2_X1 U154 ( .A1(n808), .A2(n807), .ZN(n816) );
  AND2_X1 U154bar ( .A1(n808bar), .A2(n807bar), .ZN(n816bar) );
  OR2_X1 U155 ( .A1(n806), .A2(n805), .ZN(n807) );
  AND2_X1 U155bar ( .A1(n806bar), .A2(n805bar), .ZN(n807bar) );
  OR2_X1 U156 ( .A1(in[225]), .A2(in[207]), .ZN(n805) );
  AND2_X1 U156bar ( .A1(inbar[225]), .A2(inbar[207]), .ZN(n805bar) );
  OR2_X1 U157 ( .A1(in[98]), .A2(in[226]), .ZN(n806) );
  AND2_X1 U157bar ( .A1(inbar[98]), .A2(inbar[226]), .ZN(n806bar) );
  OR2_X1 U158 ( .A1(n804), .A2(n803), .ZN(n808) );
  AND2_X1 U158bar ( .A1(n804bar), .A2(n803bar), .ZN(n808bar) );
  OR2_X1 U159 ( .A1(in_20), .A2(in_16), .ZN(n803) );
  AND2_X1 U159bar ( .A1(in_20bar), .A2(in_16bar), .ZN(n803bar) );
  OR2_X1 U160 ( .A1(in_55), .A2(in_45), .ZN(n804) );
  AND2_X1 U160bar ( .A1(in_55bar), .A2(in_45bar), .ZN(n804bar) );
  OR2_X1 U161 ( .A1(n802), .A2(n801), .ZN(n824) );
  AND2_X1 U161bar ( .A1(n802bar), .A2(n801bar), .ZN(n824bar) );
  OR2_X1 U162 ( .A1(in[162]), .A2(in[149]), .ZN(n801) );
  AND2_X1 U162bar ( .A1(inbar[162]), .A2(inbar[149]), .ZN(n801bar) );
  OR2_X1 U163 ( .A1(in[163]), .A2(n800), .ZN(n802) );
  AND2_X1 U163bar ( .A1(inbar[163]), .A2(n800bar), .ZN(n802bar) );
  OR2_X1 U164 ( .A1(in[191]), .A2(in[189]), .ZN(n800) );
  AND2_X1 U164bar ( .A1(inbar[191]), .A2(inbar[189]), .ZN(n800bar) );
  OR2_X1 U165 ( .A1(n799), .A2(n798), .ZN(n826) );
  AND2_X1 U165bar ( .A1(n799bar), .A2(n798bar), .ZN(n826bar) );
  OR2_X1 U166 ( .A1(n797), .A2(n796), .ZN(n798) );
  AND2_X1 U166bar ( .A1(n797bar), .A2(n796bar), .ZN(n798bar) );
  OR2_X1 U167 ( .A1(in[212]), .A2(in[193]), .ZN(n796) );
  AND2_X1 U167bar ( .A1(inbar[212]), .A2(inbar[193]), .ZN(n796bar) );
  OR2_X1 U168 ( .A1(in[238]), .A2(n795), .ZN(n797) );
  AND2_X1 U168bar ( .A1(inbar[238]), .A2(n795bar), .ZN(n797bar) );
  OR2_X1 U169 ( .A1(in[88]), .A2(in[247]), .ZN(n795) );
  AND2_X1 U169bar ( .A1(inbar[88]), .A2(inbar[247]), .ZN(n795bar) );
  OR2_X1 U170 ( .A1(n794), .A2(n793), .ZN(n799) );
  AND2_X1 U170bar ( .A1(n794bar), .A2(n793bar), .ZN(n799bar) );
  OR2_X1 U171 ( .A1(in[94]), .A2(in[92]), .ZN(n793) );
  AND2_X1 U171bar ( .A1(inbar[94]), .A2(inbar[92]), .ZN(n793bar) );
  OR2_X1 U172 ( .A1(in_52), .A2(n792), .ZN(n794) );
  AND2_X1 U172bar ( .A1(in_52bar), .A2(n792bar), .ZN(n794bar) );
  OR2_X1 U173 ( .A1(in_70), .A2(in_67), .ZN(n792) );
  AND2_X1 U173bar ( .A1(in_70bar), .A2(in_67bar), .ZN(n792bar) );
  OR2_X1 U174 ( .A1(n791), .A2(n790), .ZN(out[2]) );
  AND2_X1 U174bar ( .A1(n791bar), .A2(n790bar), .ZN(outbar[2]) );
  OR2_X1 U175 ( .A1(n789), .A2(n788), .ZN(n790) );
  AND2_X1 U175bar ( .A1(n789bar), .A2(n788bar), .ZN(n790bar) );
  OR2_X1 U176 ( .A1(n787), .A2(n786), .ZN(n788) );
  AND2_X1 U176bar ( .A1(n787bar), .A2(n786bar), .ZN(n788bar) );
  OR2_X1 U177 ( .A1(n819), .A2(n785), .ZN(n786) );
  AND2_X1 U177bar ( .A1(n819bar), .A2(n785bar), .ZN(n786bar) );
  OR2_X1 U178 ( .A1(n784), .A2(n783), .ZN(n819) );
  AND2_X1 U178bar ( .A1(n784bar), .A2(n783bar), .ZN(n819bar) );
  OR2_X1 U179 ( .A1(n782), .A2(n781), .ZN(n783) );
  AND2_X1 U179bar ( .A1(n782bar), .A2(n781bar), .ZN(n783bar) );
  OR2_X1 U180 ( .A1(n780), .A2(n779), .ZN(n781) );
  AND2_X1 U180bar ( .A1(n780bar), .A2(n779bar), .ZN(n781bar) );
  OR2_X1 U181 ( .A1(n962), .A2(n778), .ZN(n779) );
  AND2_X1 U181bar ( .A1(n962bar), .A2(n778bar), .ZN(n779bar) );
  OR2_X1 U182 ( .A1(n777), .A2(n776), .ZN(n962) );
  AND2_X1 U182bar ( .A1(n777bar), .A2(n776bar), .ZN(n962bar) );
  OR2_X1 U183 ( .A1(n775), .A2(n774), .ZN(n776) );
  AND2_X1 U183bar ( .A1(n775bar), .A2(n774bar), .ZN(n776bar) );
  OR2_X1 U184 ( .A1(n773), .A2(n772), .ZN(n774) );
  AND2_X1 U184bar ( .A1(n773bar), .A2(n772bar), .ZN(n774bar) );
  OR2_X1 U185 ( .A1(in[131]), .A2(in[120]), .ZN(n772) );
  AND2_X1 U185bar ( .A1(inbar[131]), .A2(inbar[120]), .ZN(n772bar) );
  OR2_X1 U186 ( .A1(in[153]), .A2(in[147]), .ZN(n773) );
  AND2_X1 U186bar ( .A1(inbar[153]), .A2(inbar[147]), .ZN(n773bar) );
  OR2_X1 U187 ( .A1(n771), .A2(n770), .ZN(n775) );
  AND2_X1 U187bar ( .A1(n771bar), .A2(n770bar), .ZN(n775bar) );
  OR2_X1 U188 ( .A1(in[170]), .A2(in[156]), .ZN(n770) );
  AND2_X1 U188bar ( .A1(inbar[170]), .A2(inbar[156]), .ZN(n770bar) );
  OR2_X1 U189 ( .A1(in[223]), .A2(in[190]), .ZN(n771) );
  AND2_X1 U189bar ( .A1(inbar[223]), .A2(inbar[190]), .ZN(n771bar) );
  OR2_X1 U190 ( .A1(n769), .A2(n768), .ZN(n777) );
  AND2_X1 U190bar ( .A1(n769bar), .A2(n768bar), .ZN(n777bar) );
  OR2_X1 U191 ( .A1(n767), .A2(n766), .ZN(n768) );
  AND2_X1 U191bar ( .A1(n767bar), .A2(n766bar), .ZN(n768bar) );
  OR2_X1 U192 ( .A1(in[236]), .A2(in[230]), .ZN(n766) );
  AND2_X1 U192bar ( .A1(inbar[236]), .A2(inbar[230]), .ZN(n766bar) );
  OR2_X1 U193 ( .A1(in[85]), .A2(in[240]), .ZN(n767) );
  AND2_X1 U193bar ( .A1(inbar[85]), .A2(inbar[240]), .ZN(n767bar) );
  OR2_X1 U194 ( .A1(n765), .A2(n764), .ZN(n769) );
  AND2_X1 U194bar ( .A1(n765bar), .A2(n764bar), .ZN(n769bar) );
  OR2_X1 U195 ( .A1(in_12), .A2(in[90]), .ZN(n764) );
  AND2_X1 U195bar ( .A1(in_12bar), .A2(inbar[90]), .ZN(n764bar) );
  OR2_X1 U196 ( .A1(in_39), .A2(in_28), .ZN(n765) );
  AND2_X1 U196bar ( .A1(in_39bar), .A2(in_28bar), .ZN(n765bar) );
  OR2_X1 U197 ( .A1(in[109]), .A2(n763), .ZN(n780) );
  AND2_X1 U197bar ( .A1(inbar[109]), .A2(n763bar), .ZN(n780bar) );
  OR2_X1 U198 ( .A1(n762), .A2(n761), .ZN(n782) );
  AND2_X1 U198bar ( .A1(n762bar), .A2(n761bar), .ZN(n782bar) );
  OR2_X1 U199 ( .A1(in[138]), .A2(in[129]), .ZN(n761) );
  AND2_X1 U199bar ( .A1(inbar[138]), .A2(inbar[129]), .ZN(n761bar) );
  OR2_X1 U200 ( .A1(in[157]), .A2(n760), .ZN(n762) );
  AND2_X1 U200bar ( .A1(inbar[157]), .A2(n760bar), .ZN(n762bar) );
  OR2_X1 U201 ( .A1(in[182]), .A2(in[167]), .ZN(n760) );
  AND2_X1 U201bar ( .A1(inbar[182]), .A2(inbar[167]), .ZN(n760bar) );
  OR2_X1 U202 ( .A1(n759), .A2(n758), .ZN(n784) );
  AND2_X1 U202bar ( .A1(n759bar), .A2(n758bar), .ZN(n784bar) );
  OR2_X1 U203 ( .A1(n757), .A2(n756), .ZN(n758) );
  AND2_X1 U203bar ( .A1(n757bar), .A2(n756bar), .ZN(n758bar) );
  OR2_X1 U204 ( .A1(in[195]), .A2(in[184]), .ZN(n756) );
  AND2_X1 U204bar ( .A1(inbar[195]), .A2(inbar[184]), .ZN(n756bar) );
  OR2_X1 U205 ( .A1(in[196]), .A2(n755), .ZN(n757) );
  AND2_X1 U205bar ( .A1(inbar[196]), .A2(n755bar), .ZN(n757bar) );
  OR2_X1 U206 ( .A1(in[215]), .A2(in[209]), .ZN(n755) );
  AND2_X1 U206bar ( .A1(inbar[215]), .A2(inbar[209]), .ZN(n755bar) );
  OR2_X1 U207 ( .A1(n754), .A2(n753), .ZN(n759) );
  AND2_X1 U207bar ( .A1(n754bar), .A2(n753bar), .ZN(n759bar) );
  OR2_X1 U208 ( .A1(in[93]), .A2(in[233]), .ZN(n753) );
  AND2_X1 U208bar ( .A1(inbar[93]), .A2(inbar[233]), .ZN(n753bar) );
  OR2_X1 U209 ( .A1(in_1), .A2(n752), .ZN(n754) );
  AND2_X1 U209bar ( .A1(in_1bar), .A2(n752bar), .ZN(n754bar) );
  OR2_X1 U210 ( .A1(in_69), .A2(in_66), .ZN(n752) );
  AND2_X1 U210bar ( .A1(in_69bar), .A2(in_66bar), .ZN(n752bar) );
  OR2_X1 U211 ( .A1(n966), .A2(n751), .ZN(n787) );
  AND2_X1 U211bar ( .A1(n966bar), .A2(n751bar), .ZN(n787bar) );
  OR2_X1 U212 ( .A1(in[134]), .A2(n750), .ZN(n751) );
  AND2_X1 U212bar ( .A1(inbar[134]), .A2(n750bar), .ZN(n751bar) );
  OR2_X1 U213 ( .A1(n749), .A2(n748), .ZN(n966) );
  AND2_X1 U213bar ( .A1(n749bar), .A2(n748bar), .ZN(n966bar) );
  OR2_X1 U214 ( .A1(n747), .A2(n746), .ZN(n748) );
  AND2_X1 U214bar ( .A1(n747bar), .A2(n746bar), .ZN(n748bar) );
  OR2_X1 U215 ( .A1(n745), .A2(n744), .ZN(n746) );
  AND2_X1 U215bar ( .A1(n745bar), .A2(n744bar), .ZN(n746bar) );
  OR2_X1 U216 ( .A1(in[136]), .A2(in[121]), .ZN(n744) );
  AND2_X1 U216bar ( .A1(inbar[136]), .A2(inbar[121]), .ZN(n744bar) );
  OR2_X1 U217 ( .A1(in[186]), .A2(in[174]), .ZN(n745) );
  AND2_X1 U217bar ( .A1(inbar[186]), .A2(inbar[174]), .ZN(n745bar) );
  OR2_X1 U218 ( .A1(n743), .A2(n742), .ZN(n747) );
  AND2_X1 U218bar ( .A1(n743bar), .A2(n742bar), .ZN(n747bar) );
  OR2_X1 U219 ( .A1(in[198]), .A2(in[197]), .ZN(n742) );
  AND2_X1 U219bar ( .A1(inbar[198]), .A2(inbar[197]), .ZN(n742bar) );
  OR2_X1 U220 ( .A1(in[214]), .A2(in[199]), .ZN(n743) );
  AND2_X1 U220bar ( .A1(inbar[214]), .A2(inbar[199]), .ZN(n743bar) );
  OR2_X1 U221 ( .A1(n741), .A2(n740), .ZN(n749) );
  AND2_X1 U221bar ( .A1(n741bar), .A2(n740bar), .ZN(n749bar) );
  OR2_X1 U222 ( .A1(n739), .A2(n738), .ZN(n740) );
  AND2_X1 U222bar ( .A1(n739bar), .A2(n738bar), .ZN(n740bar) );
  OR2_X1 U223 ( .A1(in[231]), .A2(in[220]), .ZN(n738) );
  AND2_X1 U223bar ( .A1(inbar[231]), .A2(inbar[220]), .ZN(n738bar) );
  OR2_X1 U224 ( .A1(in_25), .A2(in[245]), .ZN(n739) );
  AND2_X1 U224bar ( .A1(in_25bar), .A2(inbar[245]), .ZN(n739bar) );
  OR2_X1 U225 ( .A1(n737), .A2(n736), .ZN(n741) );
  AND2_X1 U225bar ( .A1(n737bar), .A2(n736bar), .ZN(n741bar) );
  OR2_X1 U226 ( .A1(in_53), .A2(in_29), .ZN(n736) );
  AND2_X1 U226bar ( .A1(in_53bar), .A2(in_29bar), .ZN(n736bar) );
  OR2_X1 U227 ( .A1(in_79), .A2(in_74), .ZN(n737) );
  AND2_X1 U227bar ( .A1(in_79bar), .A2(in_74bar), .ZN(n737bar) );
  OR2_X1 U228 ( .A1(n735), .A2(n734), .ZN(n789) );
  AND2_X1 U228bar ( .A1(n735bar), .A2(n734bar), .ZN(n789bar) );
  OR2_X1 U229 ( .A1(in[152]), .A2(in[140]), .ZN(n734) );
  AND2_X1 U229bar ( .A1(inbar[152]), .A2(inbar[140]), .ZN(n734bar) );
  OR2_X1 U230 ( .A1(in[155]), .A2(n733), .ZN(n735) );
  AND2_X1 U230bar ( .A1(inbar[155]), .A2(n733bar), .ZN(n735bar) );
  OR2_X1 U231 ( .A1(in[166]), .A2(in[165]), .ZN(n733) );
  AND2_X1 U231bar ( .A1(inbar[166]), .A2(inbar[165]), .ZN(n733bar) );
  OR2_X1 U232 ( .A1(n732), .A2(n731), .ZN(n791) );
  AND2_X1 U232bar ( .A1(n732bar), .A2(n731bar), .ZN(n791bar) );
  OR2_X1 U233 ( .A1(n730), .A2(n729), .ZN(n731) );
  AND2_X1 U233bar ( .A1(n730bar), .A2(n729bar), .ZN(n731bar) );
  OR2_X1 U234 ( .A1(in[202]), .A2(in[185]), .ZN(n729) );
  AND2_X1 U234bar ( .A1(inbar[202]), .A2(inbar[185]), .ZN(n729bar) );
  OR2_X1 U235 ( .A1(in[211]), .A2(n728), .ZN(n730) );
  AND2_X1 U235bar ( .A1(inbar[211]), .A2(n728bar), .ZN(n730bar) );
  OR2_X1 U236 ( .A1(in[255]), .A2(in[253]), .ZN(n728) );
  AND2_X1 U236bar ( .A1(inbar[255]), .A2(inbar[253]), .ZN(n728bar) );
  OR2_X1 U237 ( .A1(n727), .A2(n726), .ZN(n732) );
  AND2_X1 U237bar ( .A1(n727bar), .A2(n726bar), .ZN(n732bar) );
  OR2_X1 U238 ( .A1(in_35), .A2(in_15), .ZN(n726) );
  AND2_X1 U238bar ( .A1(in_35bar), .A2(in_15bar), .ZN(n726bar) );
  OR2_X1 U239 ( .A1(in_36), .A2(n725), .ZN(n727) );
  AND2_X1 U239bar ( .A1(in_36bar), .A2(n725bar), .ZN(n727bar) );
  OR2_X1 U240 ( .A1(in_48), .A2(in_40), .ZN(n725) );
  AND2_X1 U240bar ( .A1(in_48bar), .A2(in_40bar), .ZN(n725bar) );
  OR2_X1 U241 ( .A1(n724), .A2(n723), .ZN(out[1]) );
  AND2_X1 U241bar ( .A1(n724bar), .A2(n723bar), .ZN(outbar[1]) );
  OR2_X1 U242 ( .A1(n722), .A2(n721), .ZN(n723) );
  AND2_X1 U242bar ( .A1(n722bar), .A2(n721bar), .ZN(n723bar) );
  OR2_X1 U243 ( .A1(n720), .A2(n719), .ZN(n721) );
  AND2_X1 U243bar ( .A1(n720bar), .A2(n719bar), .ZN(n721bar) );
  OR2_X1 U244 ( .A1(n921), .A2(n887), .ZN(n719) );
  AND2_X1 U244bar ( .A1(n921bar), .A2(n887bar), .ZN(n719bar) );
  OR2_X1 U245 ( .A1(n718), .A2(n717), .ZN(n887) );
  AND2_X1 U245bar ( .A1(n718bar), .A2(n717bar), .ZN(n887bar) );
  OR2_X1 U246 ( .A1(n716), .A2(n715), .ZN(n717) );
  AND2_X1 U246bar ( .A1(n716bar), .A2(n715bar), .ZN(n717bar) );
  OR2_X1 U247 ( .A1(n714), .A2(n713), .ZN(n715) );
  AND2_X1 U247bar ( .A1(n714bar), .A2(n713bar), .ZN(n715bar) );
  OR2_X1 U248 ( .A1(in[116]), .A2(in[110]), .ZN(n713) );
  AND2_X1 U248bar ( .A1(inbar[116]), .A2(inbar[110]), .ZN(n713bar) );
  OR2_X1 U249 ( .A1(in[133]), .A2(in[130]), .ZN(n714) );
  AND2_X1 U249bar ( .A1(inbar[133]), .A2(inbar[130]), .ZN(n714bar) );
  OR2_X1 U250 ( .A1(n712), .A2(n711), .ZN(n716) );
  AND2_X1 U250bar ( .A1(n712bar), .A2(n711bar), .ZN(n716bar) );
  OR2_X1 U251 ( .A1(in[203]), .A2(in[135]), .ZN(n711) );
  AND2_X1 U251bar ( .A1(inbar[203]), .A2(inbar[135]), .ZN(n711bar) );
  OR2_X1 U252 ( .A1(in[232]), .A2(in[223]), .ZN(n712) );
  AND2_X1 U252bar ( .A1(inbar[232]), .A2(inbar[223]), .ZN(n712bar) );
  OR2_X1 U253 ( .A1(n710), .A2(n709), .ZN(n718) );
  AND2_X1 U253bar ( .A1(n710bar), .A2(n709bar), .ZN(n718bar) );
  OR2_X1 U254 ( .A1(n708), .A2(n707), .ZN(n709) );
  AND2_X1 U254bar ( .A1(n708bar), .A2(n707bar), .ZN(n709bar) );
  OR2_X1 U255 ( .A1(in[255]), .A2(in[233]), .ZN(n707) );
  AND2_X1 U255bar ( .A1(inbar[255]), .A2(inbar[233]), .ZN(n707bar) );
  OR2_X1 U256 ( .A1(in_53), .A2(in_34), .ZN(n708) );
  AND2_X1 U256bar ( .A1(in_53bar), .A2(in_34bar), .ZN(n708bar) );
  OR2_X1 U257 ( .A1(n706), .A2(n705), .ZN(n710) );
  AND2_X1 U257bar ( .A1(n706bar), .A2(n705bar), .ZN(n710bar) );
  OR2_X1 U258 ( .A1(in_57), .A2(in_55), .ZN(n705) );
  AND2_X1 U258bar ( .A1(in_57bar), .A2(in_55bar), .ZN(n705bar) );
  OR2_X1 U259 ( .A1(in_68), .A2(in_67), .ZN(n706) );
  AND2_X1 U259bar ( .A1(in_68bar), .A2(in_67bar), .ZN(n706bar) );
  OR2_X1 U260 ( .A1(n704), .A2(n703), .ZN(n921) );
  AND2_X1 U260bar ( .A1(n704bar), .A2(n703bar), .ZN(n921bar) );
  OR2_X1 U261 ( .A1(n702), .A2(n701), .ZN(n703) );
  AND2_X1 U261bar ( .A1(n702bar), .A2(n701bar), .ZN(n703bar) );
  OR2_X1 U262 ( .A1(n700), .A2(n699), .ZN(n701) );
  AND2_X1 U262bar ( .A1(n700bar), .A2(n699bar), .ZN(n701bar) );
  OR2_X1 U263 ( .A1(n944), .A2(n872), .ZN(n699) );
  AND2_X1 U263bar ( .A1(n944bar), .A2(n872bar), .ZN(n699bar) );
  OR2_X1 U264 ( .A1(n698), .A2(n697), .ZN(n872) );
  AND2_X1 U264bar ( .A1(n698bar), .A2(n697bar), .ZN(n872bar) );
  OR2_X1 U265 ( .A1(n696), .A2(n695), .ZN(n697) );
  AND2_X1 U265bar ( .A1(n696bar), .A2(n695bar), .ZN(n697bar) );
  OR2_X1 U266 ( .A1(n694), .A2(n693), .ZN(n695) );
  AND2_X1 U266bar ( .A1(n694bar), .A2(n693bar), .ZN(n695bar) );
  OR2_X1 U267 ( .A1(in[121]), .A2(in[102]), .ZN(n693) );
  AND2_X1 U267bar ( .A1(inbar[121]), .A2(inbar[102]), .ZN(n693bar) );
  OR2_X1 U268 ( .A1(in[162]), .A2(in[161]), .ZN(n694) );
  AND2_X1 U268bar ( .A1(inbar[162]), .A2(inbar[161]), .ZN(n694bar) );
  OR2_X1 U269 ( .A1(n692), .A2(n691), .ZN(n696) );
  AND2_X1 U269bar ( .A1(n692bar), .A2(n691bar), .ZN(n696bar) );
  OR2_X1 U270 ( .A1(in[192]), .A2(in[178]), .ZN(n691) );
  AND2_X1 U270bar ( .A1(inbar[192]), .A2(inbar[178]), .ZN(n691bar) );
  OR2_X1 U271 ( .A1(in[244]), .A2(in[209]), .ZN(n692) );
  AND2_X1 U271bar ( .A1(inbar[244]), .A2(inbar[209]), .ZN(n692bar) );
  OR2_X1 U272 ( .A1(n690), .A2(n689), .ZN(n698) );
  AND2_X1 U272bar ( .A1(n690bar), .A2(n689bar), .ZN(n698bar) );
  OR2_X1 U273 ( .A1(n688), .A2(n687), .ZN(n689) );
  AND2_X1 U273bar ( .A1(n688bar), .A2(n687bar), .ZN(n689bar) );
  OR2_X1 U274 ( .A1(in[90]), .A2(in[254]), .ZN(n687) );
  AND2_X1 U274bar ( .A1(inbar[90]), .A2(inbar[254]), .ZN(n687bar) );
  OR2_X1 U275 ( .A1(in_36), .A2(in_32), .ZN(n688) );
  AND2_X1 U275bar ( .A1(in_36bar), .A2(in_32bar), .ZN(n688bar) );
  OR2_X1 U276 ( .A1(n686), .A2(n685), .ZN(n690) );
  AND2_X1 U276bar ( .A1(n686bar), .A2(n685bar), .ZN(n690bar) );
  OR2_X1 U277 ( .A1(in_62), .A2(in_37), .ZN(n685) );
  AND2_X1 U277bar ( .A1(in_62bar), .A2(in_37bar), .ZN(n685bar) );
  OR2_X1 U278 ( .A1(in_75), .A2(in_73), .ZN(n686) );
  AND2_X1 U278bar ( .A1(in_75bar), .A2(in_73bar), .ZN(n686bar) );
  OR2_X1 U279 ( .A1(n684), .A2(n683), .ZN(n944) );
  AND2_X1 U279bar ( .A1(n684bar), .A2(n683bar), .ZN(n944bar) );
  OR2_X1 U280 ( .A1(n682), .A2(n681), .ZN(n683) );
  AND2_X1 U280bar ( .A1(n682bar), .A2(n681bar), .ZN(n683bar) );
  OR2_X1 U281 ( .A1(n680), .A2(n679), .ZN(n681) );
  AND2_X1 U281bar ( .A1(n680bar), .A2(n679bar), .ZN(n681bar) );
  OR2_X1 U282 ( .A1(in[171]), .A2(in[153]), .ZN(n679) );
  AND2_X1 U282bar ( .A1(inbar[171]), .A2(inbar[153]), .ZN(n679bar) );
  OR2_X1 U283 ( .A1(in[187]), .A2(in[176]), .ZN(n680) );
  AND2_X1 U283bar ( .A1(inbar[187]), .A2(inbar[176]), .ZN(n680bar) );
  OR2_X1 U284 ( .A1(n678), .A2(n677), .ZN(n682) );
  AND2_X1 U284bar ( .A1(n678bar), .A2(n677bar), .ZN(n682bar) );
  OR2_X1 U285 ( .A1(in[245]), .A2(in[211]), .ZN(n677) );
  AND2_X1 U285bar ( .A1(inbar[245]), .A2(inbar[211]), .ZN(n677bar) );
  OR2_X1 U286 ( .A1(in[97]), .A2(in[88]), .ZN(n678) );
  AND2_X1 U286bar ( .A1(inbar[97]), .A2(inbar[88]), .ZN(n678bar) );
  OR2_X1 U287 ( .A1(n676), .A2(n675), .ZN(n684) );
  AND2_X1 U287bar ( .A1(n676bar), .A2(n675bar), .ZN(n684bar) );
  OR2_X1 U288 ( .A1(n674), .A2(n673), .ZN(n675) );
  AND2_X1 U288bar ( .A1(n674bar), .A2(n673bar), .ZN(n675bar) );
  OR2_X1 U289 ( .A1(in_10), .A2(in_0), .ZN(n673) );
  AND2_X1 U289bar ( .A1(in_10bar), .A2(in_0bar), .ZN(n673bar) );
  OR2_X1 U290 ( .A1(in_59), .A2(in_5), .ZN(n674) );
  AND2_X1 U290bar ( .A1(in_59bar), .A2(in_5bar), .ZN(n674bar) );
  OR2_X1 U291 ( .A1(n672), .A2(n671), .ZN(n676) );
  AND2_X1 U291bar ( .A1(n672bar), .A2(n671bar), .ZN(n676bar) );
  OR2_X1 U292 ( .A1(in_60), .A2(in_6), .ZN(n671) );
  AND2_X1 U292bar ( .A1(in_60bar), .A2(in_6bar), .ZN(n671bar) );
  OR2_X1 U293 ( .A1(in_77), .A2(in_69), .ZN(n672) );
  AND2_X1 U293bar ( .A1(in_77bar), .A2(in_69bar), .ZN(n672bar) );
  OR2_X1 U294 ( .A1(in[113]), .A2(n864), .ZN(n700) );
  AND2_X1 U294bar ( .A1(inbar[113]), .A2(n864bar), .ZN(n700bar) );
  OR2_X1 U295 ( .A1(n670), .A2(n669), .ZN(n864) );
  AND2_X1 U295bar ( .A1(n670bar), .A2(n669bar), .ZN(n864bar) );
  OR2_X1 U296 ( .A1(n668), .A2(n667), .ZN(n669) );
  AND2_X1 U296bar ( .A1(n668bar), .A2(n667bar), .ZN(n669bar) );
  OR2_X1 U297 ( .A1(n666), .A2(n665), .ZN(n667) );
  AND2_X1 U297bar ( .A1(n666bar), .A2(n665bar), .ZN(n667bar) );
  OR2_X1 U298 ( .A1(in[125]), .A2(in[107]), .ZN(n665) );
  AND2_X1 U298bar ( .A1(inbar[125]), .A2(inbar[107]), .ZN(n665bar) );
  OR2_X1 U299 ( .A1(in[138]), .A2(in[126]), .ZN(n666) );
  AND2_X1 U299bar ( .A1(inbar[138]), .A2(inbar[126]), .ZN(n666bar) );
  OR2_X1 U300 ( .A1(n664), .A2(n663), .ZN(n668) );
  AND2_X1 U300bar ( .A1(n664bar), .A2(n663bar), .ZN(n668bar) );
  OR2_X1 U301 ( .A1(in[189]), .A2(in[143]), .ZN(n663) );
  AND2_X1 U301bar ( .A1(inbar[189]), .A2(inbar[143]), .ZN(n663bar) );
  OR2_X1 U302 ( .A1(in[99]), .A2(in[214]), .ZN(n664) );
  AND2_X1 U302bar ( .A1(inbar[99]), .A2(inbar[214]), .ZN(n664bar) );
  OR2_X1 U303 ( .A1(n662), .A2(n661), .ZN(n670) );
  AND2_X1 U303bar ( .A1(n662bar), .A2(n661bar), .ZN(n670bar) );
  OR2_X1 U304 ( .A1(n660), .A2(n659), .ZN(n661) );
  AND2_X1 U304bar ( .A1(n660bar), .A2(n659bar), .ZN(n661bar) );
  OR2_X1 U305 ( .A1(in_15), .A2(in_12), .ZN(n659) );
  AND2_X1 U305bar ( .A1(in_15bar), .A2(in_12bar), .ZN(n659bar) );
  OR2_X1 U306 ( .A1(in_20), .A2(in_2), .ZN(n660) );
  AND2_X1 U306bar ( .A1(in_20bar), .A2(in_2bar), .ZN(n660bar) );
  OR2_X1 U307 ( .A1(n658), .A2(n657), .ZN(n662) );
  AND2_X1 U307bar ( .A1(n658bar), .A2(n657bar), .ZN(n662bar) );
  OR2_X1 U308 ( .A1(in_30), .A2(in_3), .ZN(n657) );
  AND2_X1 U308bar ( .A1(in_30bar), .A2(in_3bar), .ZN(n657bar) );
  OR2_X1 U309 ( .A1(in_4), .A2(in_38), .ZN(n658) );
  AND2_X1 U309bar ( .A1(in_4bar), .A2(in_38bar), .ZN(n658bar) );
  OR2_X1 U310 ( .A1(n656), .A2(n655), .ZN(n702) );
  AND2_X1 U310bar ( .A1(n656bar), .A2(n655bar), .ZN(n702bar) );
  OR2_X1 U311 ( .A1(in[148]), .A2(in[137]), .ZN(n655) );
  AND2_X1 U311bar ( .A1(inbar[148]), .A2(inbar[137]), .ZN(n655bar) );
  OR2_X1 U312 ( .A1(in[149]), .A2(n654), .ZN(n656) );
  AND2_X1 U312bar ( .A1(inbar[149]), .A2(n654bar), .ZN(n656bar) );
  OR2_X1 U313 ( .A1(in[195]), .A2(in[190]), .ZN(n654) );
  AND2_X1 U313bar ( .A1(inbar[195]), .A2(inbar[190]), .ZN(n654bar) );
  OR2_X1 U314 ( .A1(n653), .A2(n652), .ZN(n704) );
  AND2_X1 U314bar ( .A1(n653bar), .A2(n652bar), .ZN(n704bar) );
  OR2_X1 U315 ( .A1(n651), .A2(n650), .ZN(n652) );
  AND2_X1 U315bar ( .A1(n651bar), .A2(n650bar), .ZN(n652bar) );
  OR2_X1 U316 ( .A1(in[98]), .A2(in[197]), .ZN(n650) );
  AND2_X1 U316bar ( .A1(inbar[98]), .A2(inbar[197]), .ZN(n650bar) );
  OR2_X1 U317 ( .A1(in_11), .A2(n649), .ZN(n651) );
  AND2_X1 U317bar ( .A1(in_11bar), .A2(n649bar), .ZN(n651bar) );
  OR2_X1 U318 ( .A1(in_26), .A2(in_14), .ZN(n649) );
  AND2_X1 U318bar ( .A1(in_26bar), .A2(in_14bar), .ZN(n649bar) );
  OR2_X1 U319 ( .A1(n648), .A2(n647), .ZN(n653) );
  AND2_X1 U319bar ( .A1(n648bar), .A2(n647bar), .ZN(n653bar) );
  OR2_X1 U320 ( .A1(in_35), .A2(in_27), .ZN(n647) );
  AND2_X1 U320bar ( .A1(in_35bar), .A2(in_27bar), .ZN(n647bar) );
  OR2_X1 U321 ( .A1(in_50), .A2(n646), .ZN(n648) );
  AND2_X1 U321bar ( .A1(in_50bar), .A2(n646bar), .ZN(n648bar) );
  OR2_X1 U322 ( .A1(in_78), .A2(in_61), .ZN(n646) );
  AND2_X1 U322bar ( .A1(in_78bar), .A2(in_61bar), .ZN(n646bar) );
  OR2_X1 U323 ( .A1(n942), .A2(n645), .ZN(n720) );
  AND2_X1 U323bar ( .A1(n942bar), .A2(n645bar), .ZN(n720bar) );
  OR2_X1 U324 ( .A1(in[106]), .A2(n863), .ZN(n645) );
  AND2_X1 U324bar ( .A1(inbar[106]), .A2(n863bar), .ZN(n645bar) );
  OR2_X1 U325 ( .A1(n644), .A2(n643), .ZN(n863) );
  AND2_X1 U325bar ( .A1(n644bar), .A2(n643bar), .ZN(n863bar) );
  OR2_X1 U326 ( .A1(n642), .A2(n641), .ZN(n643) );
  AND2_X1 U326bar ( .A1(n642bar), .A2(n641bar), .ZN(n643bar) );
  OR2_X1 U327 ( .A1(n640), .A2(n639), .ZN(n641) );
  AND2_X1 U327bar ( .A1(n640bar), .A2(n639bar), .ZN(n641bar) );
  OR2_X1 U328 ( .A1(in[127]), .A2(in[122]), .ZN(n639) );
  AND2_X1 U328bar ( .A1(inbar[127]), .A2(inbar[122]), .ZN(n639bar) );
  OR2_X1 U329 ( .A1(in[156]), .A2(in[132]), .ZN(n640) );
  AND2_X1 U329bar ( .A1(inbar[156]), .A2(inbar[132]), .ZN(n640bar) );
  OR2_X1 U330 ( .A1(n638), .A2(n637), .ZN(n642) );
  AND2_X1 U330bar ( .A1(n638bar), .A2(n637bar), .ZN(n642bar) );
  OR2_X1 U331 ( .A1(in[159]), .A2(in[157]), .ZN(n637) );
  AND2_X1 U331bar ( .A1(inbar[159]), .A2(inbar[157]), .ZN(n637bar) );
  OR2_X1 U332 ( .A1(in[185]), .A2(in[169]), .ZN(n638) );
  AND2_X1 U332bar ( .A1(inbar[185]), .A2(inbar[169]), .ZN(n638bar) );
  OR2_X1 U333 ( .A1(n636), .A2(n635), .ZN(n644) );
  AND2_X1 U333bar ( .A1(n636bar), .A2(n635bar), .ZN(n644bar) );
  OR2_X1 U334 ( .A1(n634), .A2(n633), .ZN(n635) );
  AND2_X1 U334bar ( .A1(n634bar), .A2(n633bar), .ZN(n635bar) );
  OR2_X1 U335 ( .A1(in[239]), .A2(in[218]), .ZN(n633) );
  AND2_X1 U335bar ( .A1(inbar[239]), .A2(inbar[218]), .ZN(n633bar) );
  OR2_X1 U336 ( .A1(in_13), .A2(in[87]), .ZN(n634) );
  AND2_X1 U336bar ( .A1(in_13bar), .A2(inbar[87]), .ZN(n634bar) );
  OR2_X1 U337 ( .A1(n632), .A2(n631), .ZN(n636) );
  AND2_X1 U337bar ( .A1(n632bar), .A2(n631bar), .ZN(n636bar) );
  OR2_X1 U338 ( .A1(in_72), .A2(in_70), .ZN(n631) );
  AND2_X1 U338bar ( .A1(in_72bar), .A2(in_70bar), .ZN(n631bar) );
  OR2_X1 U339 ( .A1(in_80), .A2(in_74), .ZN(n632) );
  AND2_X1 U339bar ( .A1(in_80bar), .A2(in_74bar), .ZN(n632bar) );
  OR2_X1 U340 ( .A1(n630), .A2(n629), .ZN(n942) );
  AND2_X1 U340bar ( .A1(n630bar), .A2(n629bar), .ZN(n942bar) );
  OR2_X1 U341 ( .A1(n628), .A2(n627), .ZN(n629) );
  AND2_X1 U341bar ( .A1(n628bar), .A2(n627bar), .ZN(n629bar) );
  OR2_X1 U342 ( .A1(n626), .A2(n625), .ZN(n627) );
  AND2_X1 U342bar ( .A1(n626bar), .A2(n625bar), .ZN(n627bar) );
  OR2_X1 U343 ( .A1(in[146]), .A2(in[100]), .ZN(n625) );
  AND2_X1 U343bar ( .A1(inbar[146]), .A2(inbar[100]), .ZN(n625bar) );
  OR2_X1 U344 ( .A1(in[168]), .A2(in[152]), .ZN(n626) );
  AND2_X1 U344bar ( .A1(inbar[168]), .A2(inbar[152]), .ZN(n626bar) );
  OR2_X1 U345 ( .A1(n624), .A2(n623), .ZN(n628) );
  AND2_X1 U345bar ( .A1(n624bar), .A2(n623bar), .ZN(n628bar) );
  OR2_X1 U346 ( .A1(in[199]), .A2(in[182]), .ZN(n623) );
  AND2_X1 U346bar ( .A1(inbar[199]), .A2(inbar[182]), .ZN(n623bar) );
  OR2_X1 U347 ( .A1(in[236]), .A2(in[204]), .ZN(n624) );
  AND2_X1 U347bar ( .A1(inbar[236]), .A2(inbar[204]), .ZN(n624bar) );
  OR2_X1 U348 ( .A1(n622), .A2(n621), .ZN(n630) );
  AND2_X1 U348bar ( .A1(n622bar), .A2(n621bar), .ZN(n630bar) );
  OR2_X1 U349 ( .A1(n620), .A2(n619), .ZN(n621) );
  AND2_X1 U349bar ( .A1(n620bar), .A2(n619bar), .ZN(n621bar) );
  OR2_X1 U350 ( .A1(in[89]), .A2(in[246]), .ZN(n619) );
  AND2_X1 U350bar ( .A1(inbar[89]), .A2(inbar[246]), .ZN(n619bar) );
  OR2_X1 U351 ( .A1(in[95]), .A2(in[92]), .ZN(n620) );
  AND2_X1 U351bar ( .A1(inbar[95]), .A2(inbar[92]), .ZN(n620bar) );
  OR2_X1 U352 ( .A1(n618), .A2(n617), .ZN(n622) );
  AND2_X1 U352bar ( .A1(n618bar), .A2(n617bar), .ZN(n622bar) );
  OR2_X1 U353 ( .A1(in_22), .A2(in_16), .ZN(n617) );
  AND2_X1 U353bar ( .A1(in_22bar), .A2(in_16bar), .ZN(n617bar) );
  OR2_X1 U354 ( .A1(in_51), .A2(in_49), .ZN(n618) );
  AND2_X1 U354bar ( .A1(in_51bar), .A2(in_49bar), .ZN(n618bar) );
  OR2_X1 U355 ( .A1(n616), .A2(n615), .ZN(n722) );
  AND2_X1 U355bar ( .A1(n616bar), .A2(n615bar), .ZN(n722bar) );
  OR2_X1 U356 ( .A1(in[158]), .A2(in[115]), .ZN(n615) );
  AND2_X1 U356bar ( .A1(inbar[158]), .A2(inbar[115]), .ZN(n615bar) );
  OR2_X1 U357 ( .A1(in[163]), .A2(n614), .ZN(n616) );
  AND2_X1 U357bar ( .A1(inbar[163]), .A2(n614bar), .ZN(n616bar) );
  OR2_X1 U358 ( .A1(in[206]), .A2(in[165]), .ZN(n614) );
  AND2_X1 U358bar ( .A1(inbar[206]), .A2(inbar[165]), .ZN(n614bar) );
  OR2_X1 U359 ( .A1(n613), .A2(n612), .ZN(n724) );
  AND2_X1 U359bar ( .A1(n613bar), .A2(n612bar), .ZN(n724bar) );
  OR2_X1 U360 ( .A1(n611), .A2(n610), .ZN(n612) );
  AND2_X1 U360bar ( .A1(n611bar), .A2(n610bar), .ZN(n612bar) );
  OR2_X1 U361 ( .A1(in[213]), .A2(in[207]), .ZN(n610) );
  AND2_X1 U361bar ( .A1(inbar[213]), .A2(inbar[207]), .ZN(n610bar) );
  OR2_X1 U362 ( .A1(in[215]), .A2(n609), .ZN(n611) );
  AND2_X1 U362bar ( .A1(inbar[215]), .A2(n609bar), .ZN(n611bar) );
  OR2_X1 U363 ( .A1(in[230]), .A2(in[220]), .ZN(n609) );
  AND2_X1 U363bar ( .A1(inbar[230]), .A2(inbar[220]), .ZN(n609bar) );
  OR2_X1 U364 ( .A1(n608), .A2(n607), .ZN(n613) );
  AND2_X1 U364bar ( .A1(n608bar), .A2(n607bar), .ZN(n613bar) );
  OR2_X1 U365 ( .A1(in[251]), .A2(in[234]), .ZN(n607) );
  AND2_X1 U365bar ( .A1(inbar[251]), .A2(inbar[234]), .ZN(n607bar) );
  OR2_X1 U366 ( .A1(in_17), .A2(n606), .ZN(n608) );
  AND2_X1 U366bar ( .A1(in_17bar), .A2(n606bar), .ZN(n608bar) );
  OR2_X1 U367 ( .A1(in_65), .A2(in_56), .ZN(n606) );
  AND2_X1 U367bar ( .A1(in_65bar), .A2(in_56bar), .ZN(n606bar) );
  OR2_X1 U368 ( .A1(n605), .A2(n604), .ZN(out[0]) );
  AND2_X1 U368bar ( .A1(n605bar), .A2(n604bar), .ZN(outbar[0]) );
  OR2_X1 U369 ( .A1(n603), .A2(n602), .ZN(n604) );
  AND2_X1 U369bar ( .A1(n603bar), .A2(n602bar), .ZN(n604bar) );
  OR2_X1 U370 ( .A1(n601), .A2(n600), .ZN(n602) );
  AND2_X1 U370bar ( .A1(n601bar), .A2(n600bar), .ZN(n602bar) );
  OR2_X1 U371 ( .A1(n820), .A2(n785), .ZN(n600) );
  AND2_X1 U371bar ( .A1(n820bar), .A2(n785bar), .ZN(n600bar) );
  OR2_X1 U372 ( .A1(n599), .A2(n598), .ZN(n785) );
  AND2_X1 U372bar ( .A1(n599bar), .A2(n598bar), .ZN(n785bar) );
  OR2_X1 U373 ( .A1(n597), .A2(n596), .ZN(n598) );
  AND2_X1 U373bar ( .A1(n597bar), .A2(n596bar), .ZN(n598bar) );
  OR2_X1 U374 ( .A1(n595), .A2(n594), .ZN(n596) );
  AND2_X1 U374bar ( .A1(n595bar), .A2(n594bar), .ZN(n596bar) );
  OR2_X1 U375 ( .A1(in[135]), .A2(in[104]), .ZN(n594) );
  AND2_X1 U375bar ( .A1(inbar[135]), .A2(inbar[104]), .ZN(n594bar) );
  OR2_X1 U376 ( .A1(in[188]), .A2(in[178]), .ZN(n595) );
  AND2_X1 U376bar ( .A1(inbar[188]), .A2(inbar[178]), .ZN(n595bar) );
  OR2_X1 U377 ( .A1(n593), .A2(n592), .ZN(n597) );
  AND2_X1 U377bar ( .A1(n593bar), .A2(n592bar), .ZN(n597bar) );
  OR2_X1 U378 ( .A1(in[217]), .A2(in[194]), .ZN(n592) );
  AND2_X1 U378bar ( .A1(inbar[217]), .A2(inbar[194]), .ZN(n592bar) );
  OR2_X1 U379 ( .A1(in[237]), .A2(in[218]), .ZN(n593) );
  AND2_X1 U379bar ( .A1(inbar[237]), .A2(inbar[218]), .ZN(n593bar) );
  OR2_X1 U380 ( .A1(n591), .A2(n590), .ZN(n599) );
  AND2_X1 U380bar ( .A1(n591bar), .A2(n590bar), .ZN(n599bar) );
  OR2_X1 U381 ( .A1(n589), .A2(n588), .ZN(n590) );
  AND2_X1 U381bar ( .A1(n589bar), .A2(n588bar), .ZN(n590bar) );
  OR2_X1 U382 ( .A1(in_2), .A2(in_10), .ZN(n588) );
  AND2_X1 U382bar ( .A1(in_2bar), .A2(in_10bar), .ZN(n588bar) );
  OR2_X1 U383 ( .A1(in_47), .A2(in_22), .ZN(n589) );
  AND2_X1 U383bar ( .A1(in_47bar), .A2(in_22bar), .ZN(n589bar) );
  OR2_X1 U384 ( .A1(n587), .A2(n586), .ZN(n591) );
  AND2_X1 U384bar ( .A1(n587bar), .A2(n586bar), .ZN(n591bar) );
  OR2_X1 U385 ( .A1(in_56), .A2(in_54), .ZN(n586) );
  AND2_X1 U385bar ( .A1(in_56bar), .A2(in_54bar), .ZN(n586bar) );
  OR2_X1 U386 ( .A1(in_63), .A2(in_61), .ZN(n587) );
  AND2_X1 U386bar ( .A1(in_63bar), .A2(in_61bar), .ZN(n587bar) );
  OR2_X1 U387 ( .A1(n585), .A2(n584), .ZN(n820) );
  AND2_X1 U387bar ( .A1(n585bar), .A2(n584bar), .ZN(n820bar) );
  OR2_X1 U388 ( .A1(n583), .A2(n582), .ZN(n584) );
  AND2_X1 U388bar ( .A1(n583bar), .A2(n582bar), .ZN(n584bar) );
  OR2_X1 U389 ( .A1(n581), .A2(n580), .ZN(n582) );
  AND2_X1 U389bar ( .A1(n581bar), .A2(n580bar), .ZN(n582bar) );
  OR2_X1 U390 ( .A1(in[158]), .A2(in[142]), .ZN(n580) );
  AND2_X1 U390bar ( .A1(inbar[158]), .A2(inbar[142]), .ZN(n580bar) );
  OR2_X1 U391 ( .A1(in[175]), .A2(in[164]), .ZN(n581) );
  AND2_X1 U391bar ( .A1(inbar[175]), .A2(inbar[164]), .ZN(n581bar) );
  OR2_X1 U392 ( .A1(n579), .A2(n578), .ZN(n583) );
  AND2_X1 U392bar ( .A1(n579bar), .A2(n578bar), .ZN(n583bar) );
  OR2_X1 U393 ( .A1(in[228]), .A2(in[204]), .ZN(n578) );
  AND2_X1 U393bar ( .A1(inbar[228]), .A2(inbar[204]), .ZN(n578bar) );
  OR2_X1 U394 ( .A1(in[91]), .A2(in[87]), .ZN(n579) );
  AND2_X1 U394bar ( .A1(inbar[91]), .A2(inbar[87]), .ZN(n579bar) );
  OR2_X1 U395 ( .A1(n577), .A2(n576), .ZN(n585) );
  AND2_X1 U395bar ( .A1(n577bar), .A2(n576bar), .ZN(n585bar) );
  OR2_X1 U396 ( .A1(n575), .A2(n574), .ZN(n576) );
  AND2_X1 U396bar ( .A1(n575bar), .A2(n574bar), .ZN(n576bar) );
  OR2_X1 U397 ( .A1(in_21), .A2(in_11), .ZN(n574) );
  AND2_X1 U397bar ( .A1(in_21bar), .A2(in_11bar), .ZN(n574bar) );
  OR2_X1 U398 ( .A1(in_5), .A2(in_3), .ZN(n575) );
  AND2_X1 U398bar ( .A1(in_5bar), .A2(in_3bar), .ZN(n575bar) );
  OR2_X1 U399 ( .A1(n573), .A2(n572), .ZN(n577) );
  AND2_X1 U399bar ( .A1(n573bar), .A2(n572bar), .ZN(n577bar) );
  OR2_X1 U400 ( .A1(in_68), .A2(in_64), .ZN(n572) );
  AND2_X1 U400bar ( .A1(in_68bar), .A2(in_64bar), .ZN(n572bar) );
  OR2_X1 U401 ( .A1(in_76), .A2(in_73), .ZN(n573) );
  AND2_X1 U401bar ( .A1(in_76bar), .A2(in_73bar), .ZN(n573bar) );
  OR2_X1 U402 ( .A1(n778), .A2(n571), .ZN(n601) );
  AND2_X1 U402bar ( .A1(n778bar), .A2(n571bar), .ZN(n601bar) );
  OR2_X1 U403 ( .A1(in[100]), .A2(n965), .ZN(n571) );
  AND2_X1 U403bar ( .A1(inbar[100]), .A2(n965bar), .ZN(n571bar) );
  OR2_X1 U404 ( .A1(n570), .A2(n569), .ZN(n965) );
  AND2_X1 U404bar ( .A1(n570bar), .A2(n569bar), .ZN(n965bar) );
  OR2_X1 U405 ( .A1(n568), .A2(n567), .ZN(n569) );
  AND2_X1 U405bar ( .A1(n568bar), .A2(n567bar), .ZN(n569bar) );
  OR2_X1 U406 ( .A1(n566), .A2(n565), .ZN(n567) );
  AND2_X1 U406bar ( .A1(n566bar), .A2(n565bar), .ZN(n567bar) );
  OR2_X1 U407 ( .A1(n817), .A2(n750), .ZN(n565) );
  AND2_X1 U407bar ( .A1(n817bar), .A2(n750bar), .ZN(n565bar) );
  OR2_X1 U408 ( .A1(n564), .A2(n563), .ZN(n750) );
  AND2_X1 U408bar ( .A1(n564bar), .A2(n563bar), .ZN(n750bar) );
  OR2_X1 U409 ( .A1(n562), .A2(n561), .ZN(n563) );
  AND2_X1 U409bar ( .A1(n562bar), .A2(n561bar), .ZN(n563bar) );
  OR2_X1 U410 ( .A1(n560), .A2(n559), .ZN(n561) );
  AND2_X1 U410bar ( .A1(n560bar), .A2(n559bar), .ZN(n561bar) );
  OR2_X1 U411 ( .A1(in[119]), .A2(in[103]), .ZN(n559) );
  AND2_X1 U411bar ( .A1(inbar[119]), .A2(inbar[103]), .ZN(n559bar) );
  OR2_X1 U412 ( .A1(in[137]), .A2(in[133]), .ZN(n560) );
  AND2_X1 U412bar ( .A1(inbar[137]), .A2(inbar[133]), .ZN(n560bar) );
  OR2_X1 U413 ( .A1(n558), .A2(n557), .ZN(n562) );
  AND2_X1 U413bar ( .A1(n558bar), .A2(n557bar), .ZN(n562bar) );
  OR2_X1 U414 ( .A1(in[176]), .A2(in[173]), .ZN(n557) );
  AND2_X1 U414bar ( .A1(inbar[176]), .A2(inbar[173]), .ZN(n557bar) );
  OR2_X1 U415 ( .A1(in[210]), .A2(in[181]), .ZN(n558) );
  AND2_X1 U415bar ( .A1(inbar[210]), .A2(inbar[181]), .ZN(n558bar) );
  OR2_X1 U416 ( .A1(n556), .A2(n555), .ZN(n564) );
  AND2_X1 U416bar ( .A1(n556bar), .A2(n555bar), .ZN(n564bar) );
  OR2_X1 U417 ( .A1(n554), .A2(n553), .ZN(n555) );
  AND2_X1 U417bar ( .A1(n554bar), .A2(n553bar), .ZN(n555bar) );
  OR2_X1 U418 ( .A1(in_13), .A2(in[234]), .ZN(n553) );
  AND2_X1 U418bar ( .A1(in_13bar), .A2(inbar[234]), .ZN(n553bar) );
  OR2_X1 U419 ( .A1(in_38), .A2(in_32), .ZN(n554) );
  AND2_X1 U419bar ( .A1(in_38bar), .A2(in_32bar), .ZN(n554bar) );
  OR2_X1 U420 ( .A1(n552), .A2(n551), .ZN(n556) );
  AND2_X1 U420bar ( .A1(n552bar), .A2(n551bar), .ZN(n556bar) );
  OR2_X1 U421 ( .A1(in_42), .A2(in_41), .ZN(n551) );
  AND2_X1 U421bar ( .A1(in_42bar), .A2(in_41bar), .ZN(n551bar) );
  OR2_X1 U422 ( .A1(in_7), .A2(in_49), .ZN(n552) );
  AND2_X1 U422bar ( .A1(in_7bar), .A2(in_49bar), .ZN(n552bar) );
  OR2_X1 U423 ( .A1(n550), .A2(n549), .ZN(n817) );
  AND2_X1 U423bar ( .A1(n550bar), .A2(n549bar), .ZN(n817bar) );
  OR2_X1 U424 ( .A1(n548), .A2(n547), .ZN(n549) );
  AND2_X1 U424bar ( .A1(n548bar), .A2(n547bar), .ZN(n549bar) );
  OR2_X1 U425 ( .A1(n546), .A2(n545), .ZN(n547) );
  AND2_X1 U425bar ( .A1(n546bar), .A2(n545bar), .ZN(n547bar) );
  OR2_X1 U426 ( .A1(in[159]), .A2(in[105]), .ZN(n545) );
  AND2_X1 U426bar ( .A1(inbar[159]), .A2(inbar[105]), .ZN(n545bar) );
  OR2_X1 U427 ( .A1(in[206]), .A2(in[183]), .ZN(n546) );
  AND2_X1 U427bar ( .A1(inbar[206]), .A2(inbar[183]), .ZN(n546bar) );
  OR2_X1 U428 ( .A1(n544), .A2(n543), .ZN(n548) );
  AND2_X1 U428bar ( .A1(n544bar), .A2(n543bar), .ZN(n548bar) );
  OR2_X1 U429 ( .A1(in[229]), .A2(in[219]), .ZN(n543) );
  AND2_X1 U429bar ( .A1(inbar[229]), .A2(inbar[219]), .ZN(n543bar) );
  OR2_X1 U430 ( .A1(in[235]), .A2(in[232]), .ZN(n544) );
  AND2_X1 U430bar ( .A1(inbar[235]), .A2(inbar[232]), .ZN(n544bar) );
  OR2_X1 U431 ( .A1(n542), .A2(n541), .ZN(n550) );
  AND2_X1 U431bar ( .A1(n542bar), .A2(n541bar), .ZN(n550bar) );
  OR2_X1 U432 ( .A1(n540), .A2(n539), .ZN(n541) );
  AND2_X1 U432bar ( .A1(n540bar), .A2(n539bar), .ZN(n541bar) );
  OR2_X1 U433 ( .A1(in[249]), .A2(in[242]), .ZN(n539) );
  AND2_X1 U433bar ( .A1(inbar[249]), .A2(inbar[242]), .ZN(n539bar) );
  OR2_X1 U434 ( .A1(in[89]), .A2(in[254]), .ZN(n540) );
  AND2_X1 U434bar ( .A1(inbar[89]), .A2(inbar[254]), .ZN(n540bar) );
  OR2_X1 U435 ( .A1(n538), .A2(n537), .ZN(n542) );
  AND2_X1 U435bar ( .A1(n538bar), .A2(n537bar), .ZN(n542bar) );
  OR2_X1 U436 ( .A1(in_14), .A2(in[99]), .ZN(n537) );
  AND2_X1 U436bar ( .A1(in_14bar), .A2(inbar[99]), .ZN(n537bar) );
  OR2_X1 U437 ( .A1(in_60), .A2(in_18), .ZN(n538) );
  AND2_X1 U437bar ( .A1(in_60bar), .A2(in_18bar), .ZN(n538bar) );
  OR2_X1 U438 ( .A1(in[113]), .A2(n763), .ZN(n566) );
  AND2_X1 U438bar ( .A1(inbar[113]), .A2(n763bar), .ZN(n566bar) );
  OR2_X1 U439 ( .A1(n536), .A2(n535), .ZN(n763) );
  AND2_X1 U439bar ( .A1(n536bar), .A2(n535bar), .ZN(n763bar) );
  OR2_X1 U440 ( .A1(n534), .A2(n533), .ZN(n535) );
  AND2_X1 U440bar ( .A1(n534bar), .A2(n533bar), .ZN(n535bar) );
  OR2_X1 U441 ( .A1(n532), .A2(n531), .ZN(n533) );
  AND2_X1 U441bar ( .A1(n532bar), .A2(n531bar), .ZN(n533bar) );
  OR2_X1 U442 ( .A1(in[115]), .A2(in[110]), .ZN(n531) );
  AND2_X1 U442bar ( .A1(inbar[115]), .A2(inbar[110]), .ZN(n531bar) );
  OR2_X1 U443 ( .A1(in[125]), .A2(in[117]), .ZN(n532) );
  AND2_X1 U443bar ( .A1(inbar[125]), .A2(inbar[117]), .ZN(n532bar) );
  OR2_X1 U444 ( .A1(n530), .A2(n529), .ZN(n534) );
  AND2_X1 U444bar ( .A1(n530bar), .A2(n529bar), .ZN(n534bar) );
  OR2_X1 U445 ( .A1(in[180]), .A2(in[128]), .ZN(n529) );
  AND2_X1 U445bar ( .A1(inbar[180]), .A2(inbar[128]), .ZN(n529bar) );
  OR2_X1 U446 ( .A1(in[205]), .A2(in[201]), .ZN(n530) );
  AND2_X1 U446bar ( .A1(inbar[205]), .A2(inbar[201]), .ZN(n530bar) );
  OR2_X1 U447 ( .A1(n528), .A2(n527), .ZN(n536) );
  AND2_X1 U447bar ( .A1(n528bar), .A2(n527bar), .ZN(n536bar) );
  OR2_X1 U448 ( .A1(n526), .A2(n525), .ZN(n527) );
  AND2_X1 U448bar ( .A1(n526bar), .A2(n525bar), .ZN(n527bar) );
  OR2_X1 U449 ( .A1(in[244]), .A2(in[239]), .ZN(n525) );
  AND2_X1 U449bar ( .A1(inbar[244]), .A2(inbar[239]), .ZN(n525bar) );
  OR2_X1 U450 ( .A1(in[95]), .A2(in[83]), .ZN(n526) );
  AND2_X1 U450bar ( .A1(inbar[95]), .A2(inbar[83]), .ZN(n526bar) );
  OR2_X1 U451 ( .A1(n524), .A2(n523), .ZN(n528) );
  AND2_X1 U451bar ( .A1(n524bar), .A2(n523bar), .ZN(n528bar) );
  OR2_X1 U452 ( .A1(in_24), .A2(in[97]), .ZN(n523) );
  AND2_X1 U452bar ( .A1(in_24bar), .A2(inbar[97]), .ZN(n523bar) );
  OR2_X1 U453 ( .A1(in_33), .A2(in_27), .ZN(n524) );
  AND2_X1 U453bar ( .A1(in_33bar), .A2(in_27bar), .ZN(n524bar) );
  OR2_X1 U454 ( .A1(n522), .A2(n521), .ZN(n568) );
  AND2_X1 U454bar ( .A1(n522bar), .A2(n521bar), .ZN(n568bar) );
  OR2_X1 U455 ( .A1(in[145]), .A2(in[126]), .ZN(n521) );
  AND2_X1 U455bar ( .A1(inbar[145]), .A2(inbar[126]), .ZN(n521bar) );
  OR2_X1 U456 ( .A1(in[169]), .A2(n520), .ZN(n522) );
  AND2_X1 U456bar ( .A1(inbar[169]), .A2(n520bar), .ZN(n522bar) );
  OR2_X1 U457 ( .A1(in[221]), .A2(in[172]), .ZN(n520) );
  AND2_X1 U457bar ( .A1(inbar[221]), .A2(inbar[172]), .ZN(n520bar) );
  OR2_X1 U458 ( .A1(n519), .A2(n518), .ZN(n570) );
  AND2_X1 U458bar ( .A1(n519bar), .A2(n518bar), .ZN(n570bar) );
  OR2_X1 U459 ( .A1(n517), .A2(n516), .ZN(n518) );
  AND2_X1 U459bar ( .A1(n517bar), .A2(n516bar), .ZN(n518bar) );
  OR2_X1 U460 ( .A1(in[241]), .A2(in[224]), .ZN(n516) );
  AND2_X1 U460bar ( .A1(inbar[241]), .A2(inbar[224]), .ZN(n516bar) );
  OR2_X1 U461 ( .A1(in[86]), .A2(n515), .ZN(n517) );
  AND2_X1 U461bar ( .A1(inbar[86]), .A2(n515bar), .ZN(n517bar) );
  OR2_X1 U462 ( .A1(in_43), .A2(in_34), .ZN(n515) );
  AND2_X1 U462bar ( .A1(in_43bar), .A2(in_34bar), .ZN(n515bar) );
  OR2_X1 U463 ( .A1(n514), .A2(n513), .ZN(n519) );
  AND2_X1 U463bar ( .A1(n514bar), .A2(n513bar), .ZN(n519bar) );
  OR2_X1 U464 ( .A1(in_65), .A2(in_51), .ZN(n513) );
  AND2_X1 U464bar ( .A1(in_65bar), .A2(in_51bar), .ZN(n513bar) );
  OR2_X1 U465 ( .A1(in_75), .A2(n512), .ZN(n514) );
  AND2_X1 U465bar ( .A1(in_75bar), .A2(n512bar), .ZN(n514bar) );
  OR2_X1 U466 ( .A1(in_81), .A2(in_77), .ZN(n512) );
  AND2_X1 U466bar ( .A1(in_81bar), .A2(in_77bar), .ZN(n512bar) );
  OR2_X1 U467 ( .A1(n511), .A2(n510), .ZN(n778) );
  AND2_X1 U467bar ( .A1(n511bar), .A2(n510bar), .ZN(n778bar) );
  OR2_X1 U468 ( .A1(n509), .A2(n508), .ZN(n510) );
  AND2_X1 U468bar ( .A1(n509bar), .A2(n508bar), .ZN(n510bar) );
  OR2_X1 U469 ( .A1(n507), .A2(n506), .ZN(n508) );
  AND2_X1 U469bar ( .A1(n507bar), .A2(n506bar), .ZN(n508bar) );
  OR2_X1 U470 ( .A1(in[107]), .A2(in[101]), .ZN(n506) );
  AND2_X1 U470bar ( .A1(inbar[107]), .A2(inbar[101]), .ZN(n506bar) );
  OR2_X1 U471 ( .A1(in[139]), .A2(in[132]), .ZN(n507) );
  AND2_X1 U471bar ( .A1(inbar[139]), .A2(inbar[132]), .ZN(n507bar) );
  OR2_X1 U472 ( .A1(n505), .A2(n504), .ZN(n509) );
  AND2_X1 U472bar ( .A1(n505bar), .A2(n504bar), .ZN(n509bar) );
  OR2_X1 U473 ( .A1(in[146]), .A2(in[141]), .ZN(n504) );
  AND2_X1 U473bar ( .A1(inbar[146]), .A2(inbar[141]), .ZN(n504bar) );
  OR2_X1 U474 ( .A1(in[203]), .A2(in[179]), .ZN(n505) );
  AND2_X1 U474bar ( .A1(inbar[203]), .A2(inbar[179]), .ZN(n505bar) );
  OR2_X1 U475 ( .A1(n503), .A2(n502), .ZN(n511) );
  AND2_X1 U475bar ( .A1(n503bar), .A2(n502bar), .ZN(n511bar) );
  OR2_X1 U476 ( .A1(n501), .A2(n500), .ZN(n502) );
  AND2_X1 U476bar ( .A1(n501bar), .A2(n500bar), .ZN(n502bar) );
  OR2_X1 U477 ( .A1(in[243]), .A2(in[222]), .ZN(n500) );
  AND2_X1 U477bar ( .A1(inbar[243]), .A2(inbar[222]), .ZN(n500bar) );
  OR2_X1 U478 ( .A1(in[251]), .A2(in[250]), .ZN(n501) );
  AND2_X1 U478bar ( .A1(inbar[251]), .A2(inbar[250]), .ZN(n501bar) );
  OR2_X1 U479 ( .A1(n499), .A2(n498), .ZN(n503) );
  AND2_X1 U479bar ( .A1(n499bar), .A2(n498bar), .ZN(n503bar) );
  OR2_X1 U480 ( .A1(in_37), .A2(in_19), .ZN(n498) );
  AND2_X1 U480bar ( .A1(in_37bar), .A2(in_19bar), .ZN(n498bar) );
  OR2_X1 U481 ( .A1(in_78), .A2(in_6), .ZN(n499) );
  AND2_X1 U481bar ( .A1(in_78bar), .A2(in_6bar), .ZN(n499bar) );
  OR2_X1 U482 ( .A1(n497), .A2(n496), .ZN(n603) );
  AND2_X1 U482bar ( .A1(n497bar), .A2(n496bar), .ZN(n603bar) );
  OR2_X1 U483 ( .A1(in[112]), .A2(in[102]), .ZN(n496) );
  AND2_X1 U483bar ( .A1(inbar[112]), .A2(inbar[102]), .ZN(n496bar) );
  OR2_X1 U484 ( .A1(in[123]), .A2(n495), .ZN(n497) );
  AND2_X1 U484bar ( .A1(inbar[123]), .A2(n495bar), .ZN(n497bar) );
  OR2_X1 U485 ( .A1(in[143]), .A2(in[130]), .ZN(n495) );
  AND2_X1 U485bar ( .A1(inbar[143]), .A2(inbar[130]), .ZN(n495bar) );
  OR2_X1 U486 ( .A1(n494), .A2(n493), .ZN(n605) );
  AND2_X1 U486bar ( .A1(n494bar), .A2(n493bar), .ZN(n605bar) );
  OR2_X1 U487 ( .A1(n492), .A2(n491), .ZN(n493) );
  AND2_X1 U487bar ( .A1(n492bar), .A2(n491bar), .ZN(n493bar) );
  OR2_X1 U488 ( .A1(in[216]), .A2(in[213]), .ZN(n491) );
  AND2_X1 U488bar ( .A1(inbar[216]), .A2(inbar[213]), .ZN(n491bar) );
  OR2_X1 U489 ( .A1(in[227]), .A2(n490), .ZN(n492) );
  AND2_X1 U489bar ( .A1(inbar[227]), .A2(n490bar), .ZN(n492bar) );
  OR2_X1 U490 ( .A1(in_0), .A2(in[248]), .ZN(n490) );
  AND2_X1 U490bar ( .A1(in_0bar), .A2(inbar[248]), .ZN(n490bar) );
  OR2_X1 U491 ( .A1(n489), .A2(n488), .ZN(n494) );
  AND2_X1 U491bar ( .A1(n489bar), .A2(n488bar), .ZN(n494bar) );
  OR2_X1 U492 ( .A1(in_46), .A2(in_44), .ZN(n488) );
  AND2_X1 U492bar ( .A1(in_46bar), .A2(in_44bar), .ZN(n488bar) );
  OR2_X1 U493 ( .A1(in_50), .A2(n487), .ZN(n489) );
  AND2_X1 U493bar ( .A1(in_50bar), .A2(n487bar), .ZN(n489bar) );
  OR2_X1 U494 ( .A1(in_9), .A2(in_80), .ZN(n487) );
  AND2_X1 U494bar ( .A1(in_9bar), .A2(in_80bar), .ZN(n487bar) );
endmodule

module sBox_3 ( in, inbar, out, outbar );

  input wire [7:0] in;
  input wire [7:0] inbar;
//input_done

  output wire [7:0] out;
  output wire [7:0] outbar;
//output_done

  wire [255:0] decodeOut;
  wire [255:0] decodeOutbar;
//wire_done

  decode_3 dec ( .in(in), .inbar(inbar), .out(decodeOut), .outbar(decodeOutbar) );
  encode_3 enc ( .in(decodeOut), .inbar(decodeOutbar), .out(out), .outbar(outbar) );
endmodule

module CD2_13 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD2_14 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD2_15 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD2_16 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD4_7 ( a, abar, b, bbar, y, ybar );

  input wire [3:0] a;
  input wire [3:0] b;
  input wire [3:0] abar;
  input wire [3:0] bbar;
//input_done

  output wire [15:0] y;
  output wire [15:0] ybar;
//output_done

//wire_done

  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]) );
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]) );
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]) );
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]) );
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]) );
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]) );
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]) );
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]) );
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]) );
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]) );
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]) );
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]) );
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]) );
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]) );
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]) );
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]) );
endmodule

module CD4_8 ( a, abar, b, bbar, y, ybar );

  input wire [3:0] a;
  input wire [3:0] b;
  input wire [3:0] abar;
  input wire [3:0] bbar;
//input_done

  output wire [15:0] y;
  output wire [15:0] ybar;
//output_done

//wire_done

  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]) );
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]) );
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]) );
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]) );
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]) );
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]) );
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]) );
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]) );
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]) );
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]) );
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]) );
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]) );
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]) );
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]) );
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]) );
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]) );
endmodule

module CD16_4 ( a, abar, b, bbar, y, ybar );

  input wire [15:0] a;
  input wire [15:0] b;
  input wire [15:0] abar;
  input wire [15:0] bbar;
//input_done

  output wire [255:0] y;
  output wire [255:0] ybar;
//output_done

//wire_done

  AND2_X1 U1 ( .A1(b[9]), .A2(a[0]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[9]), .A2(abar[0]), .ZN(ybar[9]) );
  AND2_X1 U2 ( .A1(b[3]), .A2(a[6]), .ZN(y[99]) );
  OR2_X1 U2bar ( .A1(bbar[3]), .A2(abar[6]), .ZN(ybar[99]) );
  AND2_X1 U3 ( .A1(b[2]), .A2(a[6]), .ZN(y[98]) );
  OR2_X1 U3bar ( .A1(bbar[2]), .A2(abar[6]), .ZN(ybar[98]) );
  AND2_X1 U4 ( .A1(b[1]), .A2(a[6]), .ZN(y[97]) );
  OR2_X1 U4bar ( .A1(bbar[1]), .A2(abar[6]), .ZN(ybar[97]) );
  AND2_X1 U5 ( .A1(b[0]), .A2(a[6]), .ZN(y[96]) );
  OR2_X1 U5bar ( .A1(bbar[0]), .A2(abar[6]), .ZN(ybar[96]) );
  AND2_X1 U6 ( .A1(b[15]), .A2(a[5]), .ZN(y[95]) );
  OR2_X1 U6bar ( .A1(bbar[15]), .A2(abar[5]), .ZN(ybar[95]) );
  AND2_X1 U7 ( .A1(b[14]), .A2(a[5]), .ZN(y[94]) );
  OR2_X1 U7bar ( .A1(bbar[14]), .A2(abar[5]), .ZN(ybar[94]) );
  AND2_X1 U8 ( .A1(b[13]), .A2(a[5]), .ZN(y[93]) );
  OR2_X1 U8bar ( .A1(bbar[13]), .A2(abar[5]), .ZN(ybar[93]) );
  AND2_X1 U9 ( .A1(b[12]), .A2(a[5]), .ZN(y[92]) );
  OR2_X1 U9bar ( .A1(bbar[12]), .A2(abar[5]), .ZN(ybar[92]) );
  AND2_X1 U10 ( .A1(b[11]), .A2(a[5]), .ZN(y[91]) );
  OR2_X1 U10bar ( .A1(bbar[11]), .A2(abar[5]), .ZN(ybar[91]) );
  AND2_X1 U11 ( .A1(b[10]), .A2(a[5]), .ZN(y[90]) );
  OR2_X1 U11bar ( .A1(bbar[10]), .A2(abar[5]), .ZN(ybar[90]) );
  AND2_X1 U12 ( .A1(b[8]), .A2(a[0]), .ZN(y[8]) );
  OR2_X1 U12bar ( .A1(bbar[8]), .A2(abar[0]), .ZN(ybar[8]) );
  AND2_X1 U13 ( .A1(a[5]), .A2(b[9]), .ZN(y[89]) );
  OR2_X1 U13bar ( .A1(abar[5]), .A2(bbar[9]), .ZN(ybar[89]) );
  AND2_X1 U14 ( .A1(b[8]), .A2(a[5]), .ZN(y[88]) );
  OR2_X1 U14bar ( .A1(bbar[8]), .A2(abar[5]), .ZN(ybar[88]) );
  AND2_X1 U15 ( .A1(b[7]), .A2(a[5]), .ZN(y[87]) );
  OR2_X1 U15bar ( .A1(bbar[7]), .A2(abar[5]), .ZN(ybar[87]) );
  AND2_X1 U16 ( .A1(b[6]), .A2(a[5]), .ZN(y[86]) );
  OR2_X1 U16bar ( .A1(bbar[6]), .A2(abar[5]), .ZN(ybar[86]) );
  AND2_X1 U17 ( .A1(b[5]), .A2(a[5]), .ZN(y[85]) );
  OR2_X1 U17bar ( .A1(bbar[5]), .A2(abar[5]), .ZN(ybar[85]) );
  AND2_X1 U18 ( .A1(b[4]), .A2(a[5]), .ZN(y[84]) );
  OR2_X1 U18bar ( .A1(bbar[4]), .A2(abar[5]), .ZN(ybar[84]) );
  AND2_X1 U19 ( .A1(a[5]), .A2(b[3]), .ZN(y[83]) );
  OR2_X1 U19bar ( .A1(abar[5]), .A2(bbar[3]), .ZN(ybar[83]) );
  AND2_X1 U20 ( .A1(a[5]), .A2(b[2]), .ZN(y[82]) );
  OR2_X1 U20bar ( .A1(abar[5]), .A2(bbar[2]), .ZN(ybar[82]) );
  AND2_X1 U21 ( .A1(a[5]), .A2(b[1]), .ZN(y[81]) );
  OR2_X1 U21bar ( .A1(abar[5]), .A2(bbar[1]), .ZN(ybar[81]) );
  AND2_X1 U22 ( .A1(a[5]), .A2(b[0]), .ZN(y[80]) );
  OR2_X1 U22bar ( .A1(abar[5]), .A2(bbar[0]), .ZN(ybar[80]) );
  AND2_X1 U23 ( .A1(b[7]), .A2(a[0]), .ZN(y[7]) );
  OR2_X1 U23bar ( .A1(bbar[7]), .A2(abar[0]), .ZN(ybar[7]) );
  AND2_X1 U24 ( .A1(a[4]), .A2(b[15]), .ZN(y[79]) );
  OR2_X1 U24bar ( .A1(abar[4]), .A2(bbar[15]), .ZN(ybar[79]) );
  AND2_X1 U25 ( .A1(a[4]), .A2(b[14]), .ZN(y[78]) );
  OR2_X1 U25bar ( .A1(abar[4]), .A2(bbar[14]), .ZN(ybar[78]) );
  AND2_X1 U26 ( .A1(a[4]), .A2(b[13]), .ZN(y[77]) );
  OR2_X1 U26bar ( .A1(abar[4]), .A2(bbar[13]), .ZN(ybar[77]) );
  AND2_X1 U27 ( .A1(a[4]), .A2(b[12]), .ZN(y[76]) );
  OR2_X1 U27bar ( .A1(abar[4]), .A2(bbar[12]), .ZN(ybar[76]) );
  AND2_X1 U28 ( .A1(a[4]), .A2(b[11]), .ZN(y[75]) );
  OR2_X1 U28bar ( .A1(abar[4]), .A2(bbar[11]), .ZN(ybar[75]) );
  AND2_X1 U29 ( .A1(a[4]), .A2(b[10]), .ZN(y[74]) );
  OR2_X1 U29bar ( .A1(abar[4]), .A2(bbar[10]), .ZN(ybar[74]) );
  AND2_X1 U30 ( .A1(a[4]), .A2(b[9]), .ZN(y[73]) );
  OR2_X1 U30bar ( .A1(abar[4]), .A2(bbar[9]), .ZN(ybar[73]) );
  AND2_X1 U31 ( .A1(a[4]), .A2(b[8]), .ZN(y[72]) );
  OR2_X1 U31bar ( .A1(abar[4]), .A2(bbar[8]), .ZN(ybar[72]) );
  AND2_X1 U32 ( .A1(a[4]), .A2(b[7]), .ZN(y[71]) );
  OR2_X1 U32bar ( .A1(abar[4]), .A2(bbar[7]), .ZN(ybar[71]) );
  AND2_X1 U33 ( .A1(a[4]), .A2(b[6]), .ZN(y[70]) );
  OR2_X1 U33bar ( .A1(abar[4]), .A2(bbar[6]), .ZN(ybar[70]) );
  AND2_X1 U34 ( .A1(b[6]), .A2(a[0]), .ZN(y[6]) );
  OR2_X1 U34bar ( .A1(bbar[6]), .A2(abar[0]), .ZN(ybar[6]) );
  AND2_X1 U35 ( .A1(a[4]), .A2(b[5]), .ZN(y[69]) );
  OR2_X1 U35bar ( .A1(abar[4]), .A2(bbar[5]), .ZN(ybar[69]) );
  AND2_X1 U36 ( .A1(a[4]), .A2(b[4]), .ZN(y[68]) );
  OR2_X1 U36bar ( .A1(abar[4]), .A2(bbar[4]), .ZN(ybar[68]) );
  AND2_X1 U37 ( .A1(a[4]), .A2(b[3]), .ZN(y[67]) );
  OR2_X1 U37bar ( .A1(abar[4]), .A2(bbar[3]), .ZN(ybar[67]) );
  AND2_X1 U38 ( .A1(a[4]), .A2(b[2]), .ZN(y[66]) );
  OR2_X1 U38bar ( .A1(abar[4]), .A2(bbar[2]), .ZN(ybar[66]) );
  AND2_X1 U39 ( .A1(a[4]), .A2(b[1]), .ZN(y[65]) );
  OR2_X1 U39bar ( .A1(abar[4]), .A2(bbar[1]), .ZN(ybar[65]) );
  AND2_X1 U40 ( .A1(a[4]), .A2(b[0]), .ZN(y[64]) );
  OR2_X1 U40bar ( .A1(abar[4]), .A2(bbar[0]), .ZN(ybar[64]) );
  AND2_X1 U41 ( .A1(a[3]), .A2(b[15]), .ZN(y[63]) );
  OR2_X1 U41bar ( .A1(abar[3]), .A2(bbar[15]), .ZN(ybar[63]) );
  AND2_X1 U42 ( .A1(a[3]), .A2(b[14]), .ZN(y[62]) );
  OR2_X1 U42bar ( .A1(abar[3]), .A2(bbar[14]), .ZN(ybar[62]) );
  AND2_X1 U43 ( .A1(a[3]), .A2(b[13]), .ZN(y[61]) );
  OR2_X1 U43bar ( .A1(abar[3]), .A2(bbar[13]), .ZN(ybar[61]) );
  AND2_X1 U44 ( .A1(a[3]), .A2(b[12]), .ZN(y[60]) );
  OR2_X1 U44bar ( .A1(abar[3]), .A2(bbar[12]), .ZN(ybar[60]) );
  AND2_X1 U45 ( .A1(b[5]), .A2(a[0]), .ZN(y[5]) );
  OR2_X1 U45bar ( .A1(bbar[5]), .A2(abar[0]), .ZN(ybar[5]) );
  AND2_X1 U46 ( .A1(a[3]), .A2(b[11]), .ZN(y[59]) );
  OR2_X1 U46bar ( .A1(abar[3]), .A2(bbar[11]), .ZN(ybar[59]) );
  AND2_X1 U47 ( .A1(a[3]), .A2(b[10]), .ZN(y[58]) );
  OR2_X1 U47bar ( .A1(abar[3]), .A2(bbar[10]), .ZN(ybar[58]) );
  AND2_X1 U48 ( .A1(a[3]), .A2(b[9]), .ZN(y[57]) );
  OR2_X1 U48bar ( .A1(abar[3]), .A2(bbar[9]), .ZN(ybar[57]) );
  AND2_X1 U49 ( .A1(a[3]), .A2(b[8]), .ZN(y[56]) );
  OR2_X1 U49bar ( .A1(abar[3]), .A2(bbar[8]), .ZN(ybar[56]) );
  AND2_X1 U50 ( .A1(a[3]), .A2(b[7]), .ZN(y[55]) );
  OR2_X1 U50bar ( .A1(abar[3]), .A2(bbar[7]), .ZN(ybar[55]) );
  AND2_X1 U51 ( .A1(a[3]), .A2(b[6]), .ZN(y[54]) );
  OR2_X1 U51bar ( .A1(abar[3]), .A2(bbar[6]), .ZN(ybar[54]) );
  AND2_X1 U52 ( .A1(a[3]), .A2(b[5]), .ZN(y[53]) );
  OR2_X1 U52bar ( .A1(abar[3]), .A2(bbar[5]), .ZN(ybar[53]) );
  AND2_X1 U53 ( .A1(a[3]), .A2(b[4]), .ZN(y[52]) );
  OR2_X1 U53bar ( .A1(abar[3]), .A2(bbar[4]), .ZN(ybar[52]) );
  AND2_X1 U54 ( .A1(a[3]), .A2(b[3]), .ZN(y[51]) );
  OR2_X1 U54bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[51]) );
  AND2_X1 U55 ( .A1(a[3]), .A2(b[2]), .ZN(y[50]) );
  OR2_X1 U55bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[50]) );
  AND2_X1 U56 ( .A1(b[4]), .A2(a[0]), .ZN(y[4]) );
  OR2_X1 U56bar ( .A1(bbar[4]), .A2(abar[0]), .ZN(ybar[4]) );
  AND2_X1 U57 ( .A1(a[3]), .A2(b[1]), .ZN(y[49]) );
  OR2_X1 U57bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[49]) );
  AND2_X1 U58 ( .A1(a[3]), .A2(b[0]), .ZN(y[48]) );
  OR2_X1 U58bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[48]) );
  AND2_X1 U59 ( .A1(a[2]), .A2(b[15]), .ZN(y[47]) );
  OR2_X1 U59bar ( .A1(abar[2]), .A2(bbar[15]), .ZN(ybar[47]) );
  AND2_X1 U60 ( .A1(a[2]), .A2(b[14]), .ZN(y[46]) );
  OR2_X1 U60bar ( .A1(abar[2]), .A2(bbar[14]), .ZN(ybar[46]) );
  AND2_X1 U61 ( .A1(a[2]), .A2(b[13]), .ZN(y[45]) );
  OR2_X1 U61bar ( .A1(abar[2]), .A2(bbar[13]), .ZN(ybar[45]) );
  AND2_X1 U62 ( .A1(a[2]), .A2(b[12]), .ZN(y[44]) );
  OR2_X1 U62bar ( .A1(abar[2]), .A2(bbar[12]), .ZN(ybar[44]) );
  AND2_X1 U63 ( .A1(a[2]), .A2(b[11]), .ZN(y[43]) );
  OR2_X1 U63bar ( .A1(abar[2]), .A2(bbar[11]), .ZN(ybar[43]) );
  AND2_X1 U64 ( .A1(a[2]), .A2(b[10]), .ZN(y[42]) );
  OR2_X1 U64bar ( .A1(abar[2]), .A2(bbar[10]), .ZN(ybar[42]) );
  AND2_X1 U65 ( .A1(a[2]), .A2(b[9]), .ZN(y[41]) );
  OR2_X1 U65bar ( .A1(abar[2]), .A2(bbar[9]), .ZN(ybar[41]) );
  AND2_X1 U66 ( .A1(a[2]), .A2(b[8]), .ZN(y[40]) );
  OR2_X1 U66bar ( .A1(abar[2]), .A2(bbar[8]), .ZN(ybar[40]) );
  AND2_X1 U67 ( .A1(b[3]), .A2(a[0]), .ZN(y[3]) );
  OR2_X1 U67bar ( .A1(bbar[3]), .A2(abar[0]), .ZN(ybar[3]) );
  AND2_X1 U68 ( .A1(a[2]), .A2(b[7]), .ZN(y[39]) );
  OR2_X1 U68bar ( .A1(abar[2]), .A2(bbar[7]), .ZN(ybar[39]) );
  AND2_X1 U69 ( .A1(a[2]), .A2(b[6]), .ZN(y[38]) );
  OR2_X1 U69bar ( .A1(abar[2]), .A2(bbar[6]), .ZN(ybar[38]) );
  AND2_X1 U70 ( .A1(a[2]), .A2(b[5]), .ZN(y[37]) );
  OR2_X1 U70bar ( .A1(abar[2]), .A2(bbar[5]), .ZN(ybar[37]) );
  AND2_X1 U71 ( .A1(a[2]), .A2(b[4]), .ZN(y[36]) );
  OR2_X1 U71bar ( .A1(abar[2]), .A2(bbar[4]), .ZN(ybar[36]) );
  AND2_X1 U72 ( .A1(a[2]), .A2(b[3]), .ZN(y[35]) );
  OR2_X1 U72bar ( .A1(abar[2]), .A2(bbar[3]), .ZN(ybar[35]) );
  AND2_X1 U73 ( .A1(a[2]), .A2(b[2]), .ZN(y[34]) );
  OR2_X1 U73bar ( .A1(abar[2]), .A2(bbar[2]), .ZN(ybar[34]) );
  AND2_X1 U74 ( .A1(a[2]), .A2(b[1]), .ZN(y[33]) );
  OR2_X1 U74bar ( .A1(abar[2]), .A2(bbar[1]), .ZN(ybar[33]) );
  AND2_X1 U75 ( .A1(a[2]), .A2(b[0]), .ZN(y[32]) );
  OR2_X1 U75bar ( .A1(abar[2]), .A2(bbar[0]), .ZN(ybar[32]) );
  AND2_X1 U76 ( .A1(a[1]), .A2(b[15]), .ZN(y[31]) );
  OR2_X1 U76bar ( .A1(abar[1]), .A2(bbar[15]), .ZN(ybar[31]) );
  AND2_X1 U77 ( .A1(a[1]), .A2(b[14]), .ZN(y[30]) );
  OR2_X1 U77bar ( .A1(abar[1]), .A2(bbar[14]), .ZN(ybar[30]) );
  AND2_X1 U78 ( .A1(b[2]), .A2(a[0]), .ZN(y[2]) );
  OR2_X1 U78bar ( .A1(bbar[2]), .A2(abar[0]), .ZN(ybar[2]) );
  AND2_X1 U79 ( .A1(a[1]), .A2(b[13]), .ZN(y[29]) );
  OR2_X1 U79bar ( .A1(abar[1]), .A2(bbar[13]), .ZN(ybar[29]) );
  AND2_X1 U80 ( .A1(a[1]), .A2(b[12]), .ZN(y[28]) );
  OR2_X1 U80bar ( .A1(abar[1]), .A2(bbar[12]), .ZN(ybar[28]) );
  AND2_X1 U81 ( .A1(a[1]), .A2(b[11]), .ZN(y[27]) );
  OR2_X1 U81bar ( .A1(abar[1]), .A2(bbar[11]), .ZN(ybar[27]) );
  AND2_X1 U82 ( .A1(a[1]), .A2(b[10]), .ZN(y[26]) );
  OR2_X1 U82bar ( .A1(abar[1]), .A2(bbar[10]), .ZN(ybar[26]) );
  AND2_X1 U83 ( .A1(a[1]), .A2(b[9]), .ZN(y[25]) );
  OR2_X1 U83bar ( .A1(abar[1]), .A2(bbar[9]), .ZN(ybar[25]) );
  AND2_X1 U84 ( .A1(a[15]), .A2(b[15]), .ZN(y[255]) );
  OR2_X1 U84bar ( .A1(abar[15]), .A2(bbar[15]), .ZN(ybar[255]) );
  AND2_X1 U85 ( .A1(a[15]), .A2(b[14]), .ZN(y[254]) );
  OR2_X1 U85bar ( .A1(abar[15]), .A2(bbar[14]), .ZN(ybar[254]) );
  AND2_X1 U86 ( .A1(a[15]), .A2(b[13]), .ZN(y[253]) );
  OR2_X1 U86bar ( .A1(abar[15]), .A2(bbar[13]), .ZN(ybar[253]) );
  AND2_X1 U87 ( .A1(a[15]), .A2(b[12]), .ZN(y[252]) );
  OR2_X1 U87bar ( .A1(abar[15]), .A2(bbar[12]), .ZN(ybar[252]) );
  AND2_X1 U88 ( .A1(a[15]), .A2(b[11]), .ZN(y[251]) );
  OR2_X1 U88bar ( .A1(abar[15]), .A2(bbar[11]), .ZN(ybar[251]) );
  AND2_X1 U89 ( .A1(a[15]), .A2(b[10]), .ZN(y[250]) );
  OR2_X1 U89bar ( .A1(abar[15]), .A2(bbar[10]), .ZN(ybar[250]) );
  AND2_X1 U90 ( .A1(a[1]), .A2(b[8]), .ZN(y[24]) );
  OR2_X1 U90bar ( .A1(abar[1]), .A2(bbar[8]), .ZN(ybar[24]) );
  AND2_X1 U91 ( .A1(a[15]), .A2(b[9]), .ZN(y[249]) );
  OR2_X1 U91bar ( .A1(abar[15]), .A2(bbar[9]), .ZN(ybar[249]) );
  AND2_X1 U92 ( .A1(a[15]), .A2(b[8]), .ZN(y[248]) );
  OR2_X1 U92bar ( .A1(abar[15]), .A2(bbar[8]), .ZN(ybar[248]) );
  AND2_X1 U93 ( .A1(a[15]), .A2(b[7]), .ZN(y[247]) );
  OR2_X1 U93bar ( .A1(abar[15]), .A2(bbar[7]), .ZN(ybar[247]) );
  AND2_X1 U94 ( .A1(a[15]), .A2(b[6]), .ZN(y[246]) );
  OR2_X1 U94bar ( .A1(abar[15]), .A2(bbar[6]), .ZN(ybar[246]) );
  AND2_X1 U95 ( .A1(a[15]), .A2(b[5]), .ZN(y[245]) );
  OR2_X1 U95bar ( .A1(abar[15]), .A2(bbar[5]), .ZN(ybar[245]) );
  AND2_X1 U96 ( .A1(a[15]), .A2(b[4]), .ZN(y[244]) );
  OR2_X1 U96bar ( .A1(abar[15]), .A2(bbar[4]), .ZN(ybar[244]) );
  AND2_X1 U97 ( .A1(a[15]), .A2(b[3]), .ZN(y[243]) );
  OR2_X1 U97bar ( .A1(abar[15]), .A2(bbar[3]), .ZN(ybar[243]) );
  AND2_X1 U98 ( .A1(a[15]), .A2(b[2]), .ZN(y[242]) );
  OR2_X1 U98bar ( .A1(abar[15]), .A2(bbar[2]), .ZN(ybar[242]) );
  AND2_X1 U99 ( .A1(a[15]), .A2(b[1]), .ZN(y[241]) );
  OR2_X1 U99bar ( .A1(abar[15]), .A2(bbar[1]), .ZN(ybar[241]) );
  AND2_X1 U100 ( .A1(a[15]), .A2(b[0]), .ZN(y[240]) );
  OR2_X1 U100bar ( .A1(abar[15]), .A2(bbar[0]), .ZN(ybar[240]) );
  AND2_X1 U101 ( .A1(a[1]), .A2(b[7]), .ZN(y[23]) );
  OR2_X1 U101bar ( .A1(abar[1]), .A2(bbar[7]), .ZN(ybar[23]) );
  AND2_X1 U102 ( .A1(a[14]), .A2(b[15]), .ZN(y[239]) );
  OR2_X1 U102bar ( .A1(abar[14]), .A2(bbar[15]), .ZN(ybar[239]) );
  AND2_X1 U103 ( .A1(a[14]), .A2(b[14]), .ZN(y[238]) );
  OR2_X1 U103bar ( .A1(abar[14]), .A2(bbar[14]), .ZN(ybar[238]) );
  AND2_X1 U104 ( .A1(a[14]), .A2(b[13]), .ZN(y[237]) );
  OR2_X1 U104bar ( .A1(abar[14]), .A2(bbar[13]), .ZN(ybar[237]) );
  AND2_X1 U105 ( .A1(a[14]), .A2(b[12]), .ZN(y[236]) );
  OR2_X1 U105bar ( .A1(abar[14]), .A2(bbar[12]), .ZN(ybar[236]) );
  AND2_X1 U106 ( .A1(a[14]), .A2(b[11]), .ZN(y[235]) );
  OR2_X1 U106bar ( .A1(abar[14]), .A2(bbar[11]), .ZN(ybar[235]) );
  AND2_X1 U107 ( .A1(a[14]), .A2(b[10]), .ZN(y[234]) );
  OR2_X1 U107bar ( .A1(abar[14]), .A2(bbar[10]), .ZN(ybar[234]) );
  AND2_X1 U108 ( .A1(a[14]), .A2(b[9]), .ZN(y[233]) );
  OR2_X1 U108bar ( .A1(abar[14]), .A2(bbar[9]), .ZN(ybar[233]) );
  AND2_X1 U109 ( .A1(a[14]), .A2(b[8]), .ZN(y[232]) );
  OR2_X1 U109bar ( .A1(abar[14]), .A2(bbar[8]), .ZN(ybar[232]) );
  AND2_X1 U110 ( .A1(a[14]), .A2(b[7]), .ZN(y[231]) );
  OR2_X1 U110bar ( .A1(abar[14]), .A2(bbar[7]), .ZN(ybar[231]) );
  AND2_X1 U111 ( .A1(a[14]), .A2(b[6]), .ZN(y[230]) );
  OR2_X1 U111bar ( .A1(abar[14]), .A2(bbar[6]), .ZN(ybar[230]) );
  AND2_X1 U112 ( .A1(a[1]), .A2(b[6]), .ZN(y[22]) );
  OR2_X1 U112bar ( .A1(abar[1]), .A2(bbar[6]), .ZN(ybar[22]) );
  AND2_X1 U113 ( .A1(a[14]), .A2(b[5]), .ZN(y[229]) );
  OR2_X1 U113bar ( .A1(abar[14]), .A2(bbar[5]), .ZN(ybar[229]) );
  AND2_X1 U114 ( .A1(a[14]), .A2(b[4]), .ZN(y[228]) );
  OR2_X1 U114bar ( .A1(abar[14]), .A2(bbar[4]), .ZN(ybar[228]) );
  AND2_X1 U115 ( .A1(a[14]), .A2(b[3]), .ZN(y[227]) );
  OR2_X1 U115bar ( .A1(abar[14]), .A2(bbar[3]), .ZN(ybar[227]) );
  AND2_X1 U116 ( .A1(a[14]), .A2(b[2]), .ZN(y[226]) );
  OR2_X1 U116bar ( .A1(abar[14]), .A2(bbar[2]), .ZN(ybar[226]) );
  AND2_X1 U117 ( .A1(a[14]), .A2(b[1]), .ZN(y[225]) );
  OR2_X1 U117bar ( .A1(abar[14]), .A2(bbar[1]), .ZN(ybar[225]) );
  AND2_X1 U118 ( .A1(a[14]), .A2(b[0]), .ZN(y[224]) );
  OR2_X1 U118bar ( .A1(abar[14]), .A2(bbar[0]), .ZN(ybar[224]) );
  AND2_X1 U119 ( .A1(a[13]), .A2(b[15]), .ZN(y[223]) );
  OR2_X1 U119bar ( .A1(abar[13]), .A2(bbar[15]), .ZN(ybar[223]) );
  AND2_X1 U120 ( .A1(a[13]), .A2(b[14]), .ZN(y[222]) );
  OR2_X1 U120bar ( .A1(abar[13]), .A2(bbar[14]), .ZN(ybar[222]) );
  AND2_X1 U121 ( .A1(a[13]), .A2(b[13]), .ZN(y[221]) );
  OR2_X1 U121bar ( .A1(abar[13]), .A2(bbar[13]), .ZN(ybar[221]) );
  AND2_X1 U122 ( .A1(a[13]), .A2(b[12]), .ZN(y[220]) );
  OR2_X1 U122bar ( .A1(abar[13]), .A2(bbar[12]), .ZN(ybar[220]) );
  AND2_X1 U123 ( .A1(a[1]), .A2(b[5]), .ZN(y[21]) );
  OR2_X1 U123bar ( .A1(abar[1]), .A2(bbar[5]), .ZN(ybar[21]) );
  AND2_X1 U124 ( .A1(a[13]), .A2(b[11]), .ZN(y[219]) );
  OR2_X1 U124bar ( .A1(abar[13]), .A2(bbar[11]), .ZN(ybar[219]) );
  AND2_X1 U125 ( .A1(a[13]), .A2(b[10]), .ZN(y[218]) );
  OR2_X1 U125bar ( .A1(abar[13]), .A2(bbar[10]), .ZN(ybar[218]) );
  AND2_X1 U126 ( .A1(a[13]), .A2(b[9]), .ZN(y[217]) );
  OR2_X1 U126bar ( .A1(abar[13]), .A2(bbar[9]), .ZN(ybar[217]) );
  AND2_X1 U127 ( .A1(a[13]), .A2(b[8]), .ZN(y[216]) );
  OR2_X1 U127bar ( .A1(abar[13]), .A2(bbar[8]), .ZN(ybar[216]) );
  AND2_X1 U128 ( .A1(a[13]), .A2(b[7]), .ZN(y[215]) );
  OR2_X1 U128bar ( .A1(abar[13]), .A2(bbar[7]), .ZN(ybar[215]) );
  AND2_X1 U129 ( .A1(a[13]), .A2(b[6]), .ZN(y[214]) );
  OR2_X1 U129bar ( .A1(abar[13]), .A2(bbar[6]), .ZN(ybar[214]) );
  AND2_X1 U130 ( .A1(a[13]), .A2(b[5]), .ZN(y[213]) );
  OR2_X1 U130bar ( .A1(abar[13]), .A2(bbar[5]), .ZN(ybar[213]) );
  AND2_X1 U131 ( .A1(a[13]), .A2(b[4]), .ZN(y[212]) );
  OR2_X1 U131bar ( .A1(abar[13]), .A2(bbar[4]), .ZN(ybar[212]) );
  AND2_X1 U132 ( .A1(a[13]), .A2(b[3]), .ZN(y[211]) );
  OR2_X1 U132bar ( .A1(abar[13]), .A2(bbar[3]), .ZN(ybar[211]) );
  AND2_X1 U133 ( .A1(a[13]), .A2(b[2]), .ZN(y[210]) );
  OR2_X1 U133bar ( .A1(abar[13]), .A2(bbar[2]), .ZN(ybar[210]) );
  AND2_X1 U134 ( .A1(a[1]), .A2(b[4]), .ZN(y[20]) );
  OR2_X1 U134bar ( .A1(abar[1]), .A2(bbar[4]), .ZN(ybar[20]) );
  AND2_X1 U135 ( .A1(a[13]), .A2(b[1]), .ZN(y[209]) );
  OR2_X1 U135bar ( .A1(abar[13]), .A2(bbar[1]), .ZN(ybar[209]) );
  AND2_X1 U136 ( .A1(a[13]), .A2(b[0]), .ZN(y[208]) );
  OR2_X1 U136bar ( .A1(abar[13]), .A2(bbar[0]), .ZN(ybar[208]) );
  AND2_X1 U137 ( .A1(a[12]), .A2(b[15]), .ZN(y[207]) );
  OR2_X1 U137bar ( .A1(abar[12]), .A2(bbar[15]), .ZN(ybar[207]) );
  AND2_X1 U138 ( .A1(a[12]), .A2(b[14]), .ZN(y[206]) );
  OR2_X1 U138bar ( .A1(abar[12]), .A2(bbar[14]), .ZN(ybar[206]) );
  AND2_X1 U139 ( .A1(a[12]), .A2(b[13]), .ZN(y[205]) );
  OR2_X1 U139bar ( .A1(abar[12]), .A2(bbar[13]), .ZN(ybar[205]) );
  AND2_X1 U140 ( .A1(a[12]), .A2(b[12]), .ZN(y[204]) );
  OR2_X1 U140bar ( .A1(abar[12]), .A2(bbar[12]), .ZN(ybar[204]) );
  AND2_X1 U141 ( .A1(a[12]), .A2(b[11]), .ZN(y[203]) );
  OR2_X1 U141bar ( .A1(abar[12]), .A2(bbar[11]), .ZN(ybar[203]) );
  AND2_X1 U142 ( .A1(a[12]), .A2(b[10]), .ZN(y[202]) );
  OR2_X1 U142bar ( .A1(abar[12]), .A2(bbar[10]), .ZN(ybar[202]) );
  AND2_X1 U143 ( .A1(a[12]), .A2(b[9]), .ZN(y[201]) );
  OR2_X1 U143bar ( .A1(abar[12]), .A2(bbar[9]), .ZN(ybar[201]) );
  AND2_X1 U144 ( .A1(a[12]), .A2(b[8]), .ZN(y[200]) );
  OR2_X1 U144bar ( .A1(abar[12]), .A2(bbar[8]), .ZN(ybar[200]) );
  AND2_X1 U145 ( .A1(b[1]), .A2(a[0]), .ZN(y[1]) );
  OR2_X1 U145bar ( .A1(bbar[1]), .A2(abar[0]), .ZN(ybar[1]) );
  AND2_X1 U146 ( .A1(a[1]), .A2(b[3]), .ZN(y[19]) );
  OR2_X1 U146bar ( .A1(abar[1]), .A2(bbar[3]), .ZN(ybar[19]) );
  AND2_X1 U147 ( .A1(a[12]), .A2(b[7]), .ZN(y[199]) );
  OR2_X1 U147bar ( .A1(abar[12]), .A2(bbar[7]), .ZN(ybar[199]) );
  AND2_X1 U148 ( .A1(a[12]), .A2(b[6]), .ZN(y[198]) );
  OR2_X1 U148bar ( .A1(abar[12]), .A2(bbar[6]), .ZN(ybar[198]) );
  AND2_X1 U149 ( .A1(a[12]), .A2(b[5]), .ZN(y[197]) );
  OR2_X1 U149bar ( .A1(abar[12]), .A2(bbar[5]), .ZN(ybar[197]) );
  AND2_X1 U150 ( .A1(a[12]), .A2(b[4]), .ZN(y[196]) );
  OR2_X1 U150bar ( .A1(abar[12]), .A2(bbar[4]), .ZN(ybar[196]) );
  AND2_X1 U151 ( .A1(a[12]), .A2(b[3]), .ZN(y[195]) );
  OR2_X1 U151bar ( .A1(abar[12]), .A2(bbar[3]), .ZN(ybar[195]) );
  AND2_X1 U152 ( .A1(a[12]), .A2(b[2]), .ZN(y[194]) );
  OR2_X1 U152bar ( .A1(abar[12]), .A2(bbar[2]), .ZN(ybar[194]) );
  AND2_X1 U153 ( .A1(a[12]), .A2(b[1]), .ZN(y[193]) );
  OR2_X1 U153bar ( .A1(abar[12]), .A2(bbar[1]), .ZN(ybar[193]) );
  AND2_X1 U154 ( .A1(a[12]), .A2(b[0]), .ZN(y[192]) );
  OR2_X1 U154bar ( .A1(abar[12]), .A2(bbar[0]), .ZN(ybar[192]) );
  AND2_X1 U155 ( .A1(a[11]), .A2(b[15]), .ZN(y[191]) );
  OR2_X1 U155bar ( .A1(abar[11]), .A2(bbar[15]), .ZN(ybar[191]) );
  AND2_X1 U156 ( .A1(a[11]), .A2(b[14]), .ZN(y[190]) );
  OR2_X1 U156bar ( .A1(abar[11]), .A2(bbar[14]), .ZN(ybar[190]) );
  AND2_X1 U157 ( .A1(a[1]), .A2(b[2]), .ZN(y[18]) );
  OR2_X1 U157bar ( .A1(abar[1]), .A2(bbar[2]), .ZN(ybar[18]) );
  AND2_X1 U158 ( .A1(a[11]), .A2(b[13]), .ZN(y[189]) );
  OR2_X1 U158bar ( .A1(abar[11]), .A2(bbar[13]), .ZN(ybar[189]) );
  AND2_X1 U159 ( .A1(a[11]), .A2(b[12]), .ZN(y[188]) );
  OR2_X1 U159bar ( .A1(abar[11]), .A2(bbar[12]), .ZN(ybar[188]) );
  AND2_X1 U160 ( .A1(a[11]), .A2(b[11]), .ZN(y[187]) );
  OR2_X1 U160bar ( .A1(abar[11]), .A2(bbar[11]), .ZN(ybar[187]) );
  AND2_X1 U161 ( .A1(a[11]), .A2(b[10]), .ZN(y[186]) );
  OR2_X1 U161bar ( .A1(abar[11]), .A2(bbar[10]), .ZN(ybar[186]) );
  AND2_X1 U162 ( .A1(a[11]), .A2(b[9]), .ZN(y[185]) );
  OR2_X1 U162bar ( .A1(abar[11]), .A2(bbar[9]), .ZN(ybar[185]) );
  AND2_X1 U163 ( .A1(a[11]), .A2(b[8]), .ZN(y[184]) );
  OR2_X1 U163bar ( .A1(abar[11]), .A2(bbar[8]), .ZN(ybar[184]) );
  AND2_X1 U164 ( .A1(a[11]), .A2(b[7]), .ZN(y[183]) );
  OR2_X1 U164bar ( .A1(abar[11]), .A2(bbar[7]), .ZN(ybar[183]) );
  AND2_X1 U165 ( .A1(a[11]), .A2(b[6]), .ZN(y[182]) );
  OR2_X1 U165bar ( .A1(abar[11]), .A2(bbar[6]), .ZN(ybar[182]) );
  AND2_X1 U166 ( .A1(a[11]), .A2(b[5]), .ZN(y[181]) );
  OR2_X1 U166bar ( .A1(abar[11]), .A2(bbar[5]), .ZN(ybar[181]) );
  AND2_X1 U167 ( .A1(a[11]), .A2(b[4]), .ZN(y[180]) );
  OR2_X1 U167bar ( .A1(abar[11]), .A2(bbar[4]), .ZN(ybar[180]) );
  AND2_X1 U168 ( .A1(a[1]), .A2(b[1]), .ZN(y[17]) );
  OR2_X1 U168bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[17]) );
  AND2_X1 U169 ( .A1(a[11]), .A2(b[3]), .ZN(y[179]) );
  OR2_X1 U169bar ( .A1(abar[11]), .A2(bbar[3]), .ZN(ybar[179]) );
  AND2_X1 U170 ( .A1(a[11]), .A2(b[2]), .ZN(y[178]) );
  OR2_X1 U170bar ( .A1(abar[11]), .A2(bbar[2]), .ZN(ybar[178]) );
  AND2_X1 U171 ( .A1(a[11]), .A2(b[1]), .ZN(y[177]) );
  OR2_X1 U171bar ( .A1(abar[11]), .A2(bbar[1]), .ZN(ybar[177]) );
  AND2_X1 U172 ( .A1(a[11]), .A2(b[0]), .ZN(y[176]) );
  OR2_X1 U172bar ( .A1(abar[11]), .A2(bbar[0]), .ZN(ybar[176]) );
  AND2_X1 U173 ( .A1(a[10]), .A2(b[15]), .ZN(y[175]) );
  OR2_X1 U173bar ( .A1(abar[10]), .A2(bbar[15]), .ZN(ybar[175]) );
  AND2_X1 U174 ( .A1(a[10]), .A2(b[14]), .ZN(y[174]) );
  OR2_X1 U174bar ( .A1(abar[10]), .A2(bbar[14]), .ZN(ybar[174]) );
  AND2_X1 U175 ( .A1(a[10]), .A2(b[13]), .ZN(y[173]) );
  OR2_X1 U175bar ( .A1(abar[10]), .A2(bbar[13]), .ZN(ybar[173]) );
  AND2_X1 U176 ( .A1(a[10]), .A2(b[12]), .ZN(y[172]) );
  OR2_X1 U176bar ( .A1(abar[10]), .A2(bbar[12]), .ZN(ybar[172]) );
  AND2_X1 U177 ( .A1(a[10]), .A2(b[11]), .ZN(y[171]) );
  OR2_X1 U177bar ( .A1(abar[10]), .A2(bbar[11]), .ZN(ybar[171]) );
  AND2_X1 U178 ( .A1(a[10]), .A2(b[10]), .ZN(y[170]) );
  OR2_X1 U178bar ( .A1(abar[10]), .A2(bbar[10]), .ZN(ybar[170]) );
  AND2_X1 U179 ( .A1(a[1]), .A2(b[0]), .ZN(y[16]) );
  OR2_X1 U179bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[16]) );
  AND2_X1 U180 ( .A1(a[10]), .A2(b[9]), .ZN(y[169]) );
  OR2_X1 U180bar ( .A1(abar[10]), .A2(bbar[9]), .ZN(ybar[169]) );
  AND2_X1 U181 ( .A1(a[10]), .A2(b[8]), .ZN(y[168]) );
  OR2_X1 U181bar ( .A1(abar[10]), .A2(bbar[8]), .ZN(ybar[168]) );
  AND2_X1 U182 ( .A1(a[10]), .A2(b[7]), .ZN(y[167]) );
  OR2_X1 U182bar ( .A1(abar[10]), .A2(bbar[7]), .ZN(ybar[167]) );
  AND2_X1 U183 ( .A1(a[10]), .A2(b[6]), .ZN(y[166]) );
  OR2_X1 U183bar ( .A1(abar[10]), .A2(bbar[6]), .ZN(ybar[166]) );
  AND2_X1 U184 ( .A1(a[10]), .A2(b[5]), .ZN(y[165]) );
  OR2_X1 U184bar ( .A1(abar[10]), .A2(bbar[5]), .ZN(ybar[165]) );
  AND2_X1 U185 ( .A1(a[10]), .A2(b[4]), .ZN(y[164]) );
  OR2_X1 U185bar ( .A1(abar[10]), .A2(bbar[4]), .ZN(ybar[164]) );
  AND2_X1 U186 ( .A1(a[10]), .A2(b[3]), .ZN(y[163]) );
  OR2_X1 U186bar ( .A1(abar[10]), .A2(bbar[3]), .ZN(ybar[163]) );
  AND2_X1 U187 ( .A1(a[10]), .A2(b[2]), .ZN(y[162]) );
  OR2_X1 U187bar ( .A1(abar[10]), .A2(bbar[2]), .ZN(ybar[162]) );
  AND2_X1 U188 ( .A1(a[10]), .A2(b[1]), .ZN(y[161]) );
  OR2_X1 U188bar ( .A1(abar[10]), .A2(bbar[1]), .ZN(ybar[161]) );
  AND2_X1 U189 ( .A1(a[10]), .A2(b[0]), .ZN(y[160]) );
  OR2_X1 U189bar ( .A1(abar[10]), .A2(bbar[0]), .ZN(ybar[160]) );
  AND2_X1 U190 ( .A1(b[15]), .A2(a[0]), .ZN(y[15]) );
  OR2_X1 U190bar ( .A1(bbar[15]), .A2(abar[0]), .ZN(ybar[15]) );
  AND2_X1 U191 ( .A1(a[9]), .A2(b[15]), .ZN(y[159]) );
  OR2_X1 U191bar ( .A1(abar[9]), .A2(bbar[15]), .ZN(ybar[159]) );
  AND2_X1 U192 ( .A1(a[9]), .A2(b[14]), .ZN(y[158]) );
  OR2_X1 U192bar ( .A1(abar[9]), .A2(bbar[14]), .ZN(ybar[158]) );
  AND2_X1 U193 ( .A1(a[9]), .A2(b[13]), .ZN(y[157]) );
  OR2_X1 U193bar ( .A1(abar[9]), .A2(bbar[13]), .ZN(ybar[157]) );
  AND2_X1 U194 ( .A1(a[9]), .A2(b[12]), .ZN(y[156]) );
  OR2_X1 U194bar ( .A1(abar[9]), .A2(bbar[12]), .ZN(ybar[156]) );
  AND2_X1 U195 ( .A1(a[9]), .A2(b[11]), .ZN(y[155]) );
  OR2_X1 U195bar ( .A1(abar[9]), .A2(bbar[11]), .ZN(ybar[155]) );
  AND2_X1 U196 ( .A1(a[9]), .A2(b[10]), .ZN(y[154]) );
  OR2_X1 U196bar ( .A1(abar[9]), .A2(bbar[10]), .ZN(ybar[154]) );
  AND2_X1 U197 ( .A1(a[9]), .A2(b[9]), .ZN(y[153]) );
  OR2_X1 U197bar ( .A1(abar[9]), .A2(bbar[9]), .ZN(ybar[153]) );
  AND2_X1 U198 ( .A1(a[9]), .A2(b[8]), .ZN(y[152]) );
  OR2_X1 U198bar ( .A1(abar[9]), .A2(bbar[8]), .ZN(ybar[152]) );
  AND2_X1 U199 ( .A1(a[9]), .A2(b[7]), .ZN(y[151]) );
  OR2_X1 U199bar ( .A1(abar[9]), .A2(bbar[7]), .ZN(ybar[151]) );
  AND2_X1 U200 ( .A1(a[9]), .A2(b[6]), .ZN(y[150]) );
  OR2_X1 U200bar ( .A1(abar[9]), .A2(bbar[6]), .ZN(ybar[150]) );
  AND2_X1 U201 ( .A1(b[14]), .A2(a[0]), .ZN(y[14]) );
  OR2_X1 U201bar ( .A1(bbar[14]), .A2(abar[0]), .ZN(ybar[14]) );
  AND2_X1 U202 ( .A1(a[9]), .A2(b[5]), .ZN(y[149]) );
  OR2_X1 U202bar ( .A1(abar[9]), .A2(bbar[5]), .ZN(ybar[149]) );
  AND2_X1 U203 ( .A1(a[9]), .A2(b[4]), .ZN(y[148]) );
  OR2_X1 U203bar ( .A1(abar[9]), .A2(bbar[4]), .ZN(ybar[148]) );
  AND2_X1 U204 ( .A1(a[9]), .A2(b[3]), .ZN(y[147]) );
  OR2_X1 U204bar ( .A1(abar[9]), .A2(bbar[3]), .ZN(ybar[147]) );
  AND2_X1 U205 ( .A1(a[9]), .A2(b[2]), .ZN(y[146]) );
  OR2_X1 U205bar ( .A1(abar[9]), .A2(bbar[2]), .ZN(ybar[146]) );
  AND2_X1 U206 ( .A1(a[9]), .A2(b[1]), .ZN(y[145]) );
  OR2_X1 U206bar ( .A1(abar[9]), .A2(bbar[1]), .ZN(ybar[145]) );
  AND2_X1 U207 ( .A1(a[9]), .A2(b[0]), .ZN(y[144]) );
  OR2_X1 U207bar ( .A1(abar[9]), .A2(bbar[0]), .ZN(ybar[144]) );
  AND2_X1 U208 ( .A1(a[8]), .A2(b[15]), .ZN(y[143]) );
  OR2_X1 U208bar ( .A1(abar[8]), .A2(bbar[15]), .ZN(ybar[143]) );
  AND2_X1 U209 ( .A1(a[8]), .A2(b[14]), .ZN(y[142]) );
  OR2_X1 U209bar ( .A1(abar[8]), .A2(bbar[14]), .ZN(ybar[142]) );
  AND2_X1 U210 ( .A1(a[8]), .A2(b[13]), .ZN(y[141]) );
  OR2_X1 U210bar ( .A1(abar[8]), .A2(bbar[13]), .ZN(ybar[141]) );
  AND2_X1 U211 ( .A1(a[8]), .A2(b[12]), .ZN(y[140]) );
  OR2_X1 U211bar ( .A1(abar[8]), .A2(bbar[12]), .ZN(ybar[140]) );
  AND2_X1 U212 ( .A1(b[13]), .A2(a[0]), .ZN(y[13]) );
  OR2_X1 U212bar ( .A1(bbar[13]), .A2(abar[0]), .ZN(ybar[13]) );
  AND2_X1 U213 ( .A1(a[8]), .A2(b[11]), .ZN(y[139]) );
  OR2_X1 U213bar ( .A1(abar[8]), .A2(bbar[11]), .ZN(ybar[139]) );
  AND2_X1 U214 ( .A1(a[8]), .A2(b[10]), .ZN(y[138]) );
  OR2_X1 U214bar ( .A1(abar[8]), .A2(bbar[10]), .ZN(ybar[138]) );
  AND2_X1 U215 ( .A1(a[8]), .A2(b[9]), .ZN(y[137]) );
  OR2_X1 U215bar ( .A1(abar[8]), .A2(bbar[9]), .ZN(ybar[137]) );
  AND2_X1 U216 ( .A1(a[8]), .A2(b[8]), .ZN(y[136]) );
  OR2_X1 U216bar ( .A1(abar[8]), .A2(bbar[8]), .ZN(ybar[136]) );
  AND2_X1 U217 ( .A1(a[8]), .A2(b[7]), .ZN(y[135]) );
  OR2_X1 U217bar ( .A1(abar[8]), .A2(bbar[7]), .ZN(ybar[135]) );
  AND2_X1 U218 ( .A1(a[8]), .A2(b[6]), .ZN(y[134]) );
  OR2_X1 U218bar ( .A1(abar[8]), .A2(bbar[6]), .ZN(ybar[134]) );
  AND2_X1 U219 ( .A1(a[8]), .A2(b[5]), .ZN(y[133]) );
  OR2_X1 U219bar ( .A1(abar[8]), .A2(bbar[5]), .ZN(ybar[133]) );
  AND2_X1 U220 ( .A1(a[8]), .A2(b[4]), .ZN(y[132]) );
  OR2_X1 U220bar ( .A1(abar[8]), .A2(bbar[4]), .ZN(ybar[132]) );
  AND2_X1 U221 ( .A1(a[8]), .A2(b[3]), .ZN(y[131]) );
  OR2_X1 U221bar ( .A1(abar[8]), .A2(bbar[3]), .ZN(ybar[131]) );
  AND2_X1 U222 ( .A1(a[8]), .A2(b[2]), .ZN(y[130]) );
  OR2_X1 U222bar ( .A1(abar[8]), .A2(bbar[2]), .ZN(ybar[130]) );
  AND2_X1 U223 ( .A1(b[12]), .A2(a[0]), .ZN(y[12]) );
  OR2_X1 U223bar ( .A1(bbar[12]), .A2(abar[0]), .ZN(ybar[12]) );
  AND2_X1 U224 ( .A1(a[8]), .A2(b[1]), .ZN(y[129]) );
  OR2_X1 U224bar ( .A1(abar[8]), .A2(bbar[1]), .ZN(ybar[129]) );
  AND2_X1 U225 ( .A1(a[8]), .A2(b[0]), .ZN(y[128]) );
  OR2_X1 U225bar ( .A1(abar[8]), .A2(bbar[0]), .ZN(ybar[128]) );
  AND2_X1 U226 ( .A1(a[7]), .A2(b[15]), .ZN(y[127]) );
  OR2_X1 U226bar ( .A1(abar[7]), .A2(bbar[15]), .ZN(ybar[127]) );
  AND2_X1 U227 ( .A1(a[7]), .A2(b[14]), .ZN(y[126]) );
  OR2_X1 U227bar ( .A1(abar[7]), .A2(bbar[14]), .ZN(ybar[126]) );
  AND2_X1 U228 ( .A1(a[7]), .A2(b[13]), .ZN(y[125]) );
  OR2_X1 U228bar ( .A1(abar[7]), .A2(bbar[13]), .ZN(ybar[125]) );
  AND2_X1 U229 ( .A1(a[7]), .A2(b[12]), .ZN(y[124]) );
  OR2_X1 U229bar ( .A1(abar[7]), .A2(bbar[12]), .ZN(ybar[124]) );
  AND2_X1 U230 ( .A1(a[7]), .A2(b[11]), .ZN(y[123]) );
  OR2_X1 U230bar ( .A1(abar[7]), .A2(bbar[11]), .ZN(ybar[123]) );
  AND2_X1 U231 ( .A1(a[7]), .A2(b[10]), .ZN(y[122]) );
  OR2_X1 U231bar ( .A1(abar[7]), .A2(bbar[10]), .ZN(ybar[122]) );
  AND2_X1 U232 ( .A1(a[7]), .A2(b[9]), .ZN(y[121]) );
  OR2_X1 U232bar ( .A1(abar[7]), .A2(bbar[9]), .ZN(ybar[121]) );
  AND2_X1 U233 ( .A1(a[7]), .A2(b[8]), .ZN(y[120]) );
  OR2_X1 U233bar ( .A1(abar[7]), .A2(bbar[8]), .ZN(ybar[120]) );
  AND2_X1 U234 ( .A1(b[11]), .A2(a[0]), .ZN(y[11]) );
  OR2_X1 U234bar ( .A1(bbar[11]), .A2(abar[0]), .ZN(ybar[11]) );
  AND2_X1 U235 ( .A1(a[7]), .A2(b[7]), .ZN(y[119]) );
  OR2_X1 U235bar ( .A1(abar[7]), .A2(bbar[7]), .ZN(ybar[119]) );
  AND2_X1 U236 ( .A1(a[7]), .A2(b[6]), .ZN(y[118]) );
  OR2_X1 U236bar ( .A1(abar[7]), .A2(bbar[6]), .ZN(ybar[118]) );
  AND2_X1 U237 ( .A1(a[7]), .A2(b[5]), .ZN(y[117]) );
  OR2_X1 U237bar ( .A1(abar[7]), .A2(bbar[5]), .ZN(ybar[117]) );
  AND2_X1 U238 ( .A1(a[7]), .A2(b[4]), .ZN(y[116]) );
  OR2_X1 U238bar ( .A1(abar[7]), .A2(bbar[4]), .ZN(ybar[116]) );
  AND2_X1 U239 ( .A1(a[7]), .A2(b[3]), .ZN(y[115]) );
  OR2_X1 U239bar ( .A1(abar[7]), .A2(bbar[3]), .ZN(ybar[115]) );
  AND2_X1 U240 ( .A1(a[7]), .A2(b[2]), .ZN(y[114]) );
  OR2_X1 U240bar ( .A1(abar[7]), .A2(bbar[2]), .ZN(ybar[114]) );
  AND2_X1 U241 ( .A1(a[7]), .A2(b[1]), .ZN(y[113]) );
  OR2_X1 U241bar ( .A1(abar[7]), .A2(bbar[1]), .ZN(ybar[113]) );
  AND2_X1 U242 ( .A1(a[7]), .A2(b[0]), .ZN(y[112]) );
  OR2_X1 U242bar ( .A1(abar[7]), .A2(bbar[0]), .ZN(ybar[112]) );
  AND2_X1 U243 ( .A1(b[15]), .A2(a[6]), .ZN(y[111]) );
  OR2_X1 U243bar ( .A1(bbar[15]), .A2(abar[6]), .ZN(ybar[111]) );
  AND2_X1 U244 ( .A1(b[14]), .A2(a[6]), .ZN(y[110]) );
  OR2_X1 U244bar ( .A1(bbar[14]), .A2(abar[6]), .ZN(ybar[110]) );
  AND2_X1 U245 ( .A1(b[10]), .A2(a[0]), .ZN(y[10]) );
  OR2_X1 U245bar ( .A1(bbar[10]), .A2(abar[0]), .ZN(ybar[10]) );
  AND2_X1 U246 ( .A1(b[13]), .A2(a[6]), .ZN(y[109]) );
  OR2_X1 U246bar ( .A1(bbar[13]), .A2(abar[6]), .ZN(ybar[109]) );
  AND2_X1 U247 ( .A1(b[12]), .A2(a[6]), .ZN(y[108]) );
  OR2_X1 U247bar ( .A1(bbar[12]), .A2(abar[6]), .ZN(ybar[108]) );
  AND2_X1 U248 ( .A1(b[11]), .A2(a[6]), .ZN(y[107]) );
  OR2_X1 U248bar ( .A1(bbar[11]), .A2(abar[6]), .ZN(ybar[107]) );
  AND2_X1 U249 ( .A1(b[10]), .A2(a[6]), .ZN(y[106]) );
  OR2_X1 U249bar ( .A1(bbar[10]), .A2(abar[6]), .ZN(ybar[106]) );
  AND2_X1 U250 ( .A1(a[6]), .A2(b[9]), .ZN(y[105]) );
  OR2_X1 U250bar ( .A1(abar[6]), .A2(bbar[9]), .ZN(ybar[105]) );
  AND2_X1 U251 ( .A1(b[8]), .A2(a[6]), .ZN(y[104]) );
  OR2_X1 U251bar ( .A1(bbar[8]), .A2(abar[6]), .ZN(ybar[104]) );
  AND2_X1 U252 ( .A1(b[7]), .A2(a[6]), .ZN(y[103]) );
  OR2_X1 U252bar ( .A1(bbar[7]), .A2(abar[6]), .ZN(ybar[103]) );
  AND2_X1 U253 ( .A1(b[6]), .A2(a[6]), .ZN(y[102]) );
  OR2_X1 U253bar ( .A1(bbar[6]), .A2(abar[6]), .ZN(ybar[102]) );
  AND2_X1 U254 ( .A1(b[5]), .A2(a[6]), .ZN(y[101]) );
  OR2_X1 U254bar ( .A1(bbar[5]), .A2(abar[6]), .ZN(ybar[101]) );
  AND2_X1 U255 ( .A1(b[4]), .A2(a[6]), .ZN(y[100]) );
  OR2_X1 U255bar ( .A1(bbar[4]), .A2(abar[6]), .ZN(ybar[100]) );
  AND2_X1 U256 ( .A1(b[0]), .A2(a[0]), .ZN(y[0]) );
  OR2_X1 U256bar ( .A1(bbar[0]), .A2(abar[0]), .ZN(ybar[0]) );
endmodule

module decode_4 ( in, inbar, out, outbar );

  input wire [7:0] in;
  input wire [7:0] inbar;
//input_done

  output wire [255:0] out;
  output wire [255:0] outbar;
//output_done

  wire [15:0] level1;
  wire [31:0] level2;
  wire [15:0] level1bar;
  wire [31:0] level2bar;
//wire_done

  CD2_16 cd_l1_1 ( .a(in[1]), .abar(inbar[1]), .b(in[0]), .bbar(inbar[0]), .y(level1[3:0]), .ybar(level1bar[3:0]) );
  CD2_15 cd_l1_2 ( .a(in[3]), .abar(inbar[3]), .b(in[2]), .bbar(inbar[2]), .y(level1[7:4]), .ybar(level1bar[7:4]) );
  CD2_14 cd_l1_3 ( .a(in[5]), .abar(inbar[5]), .b(in[4]), .bbar(inbar[4]), .y(level1[11:8]), .ybar(level1bar[11:8]) );
  CD2_13 cd_l1_4 ( .a(in[7]), .abar(inbar[7]), .b(in[6]), .bbar(inbar[6]), .y(level1[15:12]), .ybar(level1bar[15:12]) );

  CD4_8 cd_l2_1 ( .a(level1[7:4]), .abar(level1bar[7:4]), .b(level1[3:0]), .bbar(level1bar[3:0]), 
        .y(level2[15:0]), .ybar(level2bar[15:0]) );
  CD4_7 cd_l2_2 ( .a(level1[15:12]), .abar(level1bar[15:12]), .b(level1[11:8]), .bbar(level1bar[11:8]), 
        .y(level2[31:16]), .ybar(level2bar[31:16]) );
  CD16_4 cd_l3 ( .a(level2[31:16]), .abar(level2bar[31:16]), .b(level2[15:0]), .bbar(level2bar[15:0]), 
        .y(out), .ybar(outbar) );
endmodule

module encode_4 ( in, inbar, out, outbar );

  input wire [255:0] in;
  input wire [255:0] inbar;
//input_done

  output wire [7:0] out;
  output wire [7:0] outbar;
//output_done

  wire in_81;
  wire in_80;
  wire in_79;
  wire in_78;
  wire in_77;
  wire in_76;
  wire in_75;
  wire in_74;
  wire in_73;
  wire in_72;
  wire in_71;
  wire in_70;
  wire in_69;
  wire in_68;
  wire in_67;
  wire in_66;
  wire in_65;
  wire in_64;
  wire in_63;
  wire in_62;
  wire in_61;
  wire in_60;
  wire in_59;
  wire in_58;
  wire in_57;
  wire in_56;
  wire in_55;
  wire in_54;
  wire in_53;
  wire in_52;
  wire in_51;
  wire in_50;
  wire in_49;
  wire in_48;
  wire in_47;
  wire in_46;
  wire in_45;
  wire in_44;
  wire in_43;
  wire in_42;
  wire in_41;
  wire in_40;
  wire in_39;
  wire in_38;
  wire in_37;
  wire in_36;
  wire in_35;
  wire in_34;
  wire in_33;
  wire in_32;
  wire in_31;
  wire in_30;
  wire in_29;
  wire in_28;
  wire in_27;
  wire in_26;
  wire in_25;
  wire in_24;
  wire in_23;
  wire in_22;
  wire in_21;
  wire in_20;
  wire in_19;
  wire in_18;
  wire in_17;
  wire in_16;
  wire in_15;
  wire in_14;
  wire in_13;
  wire in_12;
  wire in_11;
  wire in_10;
  wire in_9;
  wire in_8;
  wire in_7;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_3;
  wire in_2;
  wire in_1;
  wire in_0;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire in_81bar;
  wire in_80bar;
  wire in_79bar;
  wire in_78bar;
  wire in_77bar;
  wire in_76bar;
  wire in_75bar;
  wire in_74bar;
  wire in_73bar;
  wire in_72bar;
  wire in_71bar;
  wire in_70bar;
  wire in_69bar;
  wire in_68bar;
  wire in_67bar;
  wire in_66bar;
  wire in_65bar;
  wire in_64bar;
  wire in_63bar;
  wire in_62bar;
  wire in_61bar;
  wire in_60bar;
  wire in_59bar;
  wire in_58bar;
  wire in_57bar;
  wire in_56bar;
  wire in_55bar;
  wire in_54bar;
  wire in_53bar;
  wire in_52bar;
  wire in_51bar;
  wire in_50bar;
  wire in_49bar;
  wire in_48bar;
  wire in_47bar;
  wire in_46bar;
  wire in_45bar;
  wire in_44bar;
  wire in_43bar;
  wire in_42bar;
  wire in_41bar;
  wire in_40bar;
  wire in_39bar;
  wire in_38bar;
  wire in_37bar;
  wire in_36bar;
  wire in_35bar;
  wire in_34bar;
  wire in_33bar;
  wire in_32bar;
  wire in_31bar;
  wire in_30bar;
  wire in_29bar;
  wire in_28bar;
  wire in_27bar;
  wire in_26bar;
  wire in_25bar;
  wire in_24bar;
  wire in_23bar;
  wire in_22bar;
  wire in_21bar;
  wire in_20bar;
  wire in_19bar;
  wire in_18bar;
  wire in_17bar;
  wire in_16bar;
  wire in_15bar;
  wire in_14bar;
  wire in_13bar;
  wire in_12bar;
  wire in_11bar;
  wire in_10bar;
  wire in_9bar;
  wire in_8bar;
  wire in_7bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_3bar;
  wire in_2bar;
  wire in_1bar;
  wire in_0bar;
  wire n487bar;
  wire n488bar;
  wire n489bar;
  wire n490bar;
  wire n491bar;
  wire n492bar;
  wire n493bar;
  wire n494bar;
  wire n495bar;
  wire n496bar;
  wire n497bar;
  wire n498bar;
  wire n499bar;
  wire n500bar;
  wire n501bar;
  wire n502bar;
  wire n503bar;
  wire n504bar;
  wire n505bar;
  wire n506bar;
  wire n507bar;
  wire n508bar;
  wire n509bar;
  wire n510bar;
  wire n511bar;
  wire n512bar;
  wire n513bar;
  wire n514bar;
  wire n515bar;
  wire n516bar;
  wire n517bar;
  wire n518bar;
  wire n519bar;
  wire n520bar;
  wire n521bar;
  wire n522bar;
  wire n523bar;
  wire n524bar;
  wire n525bar;
  wire n526bar;
  wire n527bar;
  wire n528bar;
  wire n529bar;
  wire n530bar;
  wire n531bar;
  wire n532bar;
  wire n533bar;
  wire n534bar;
  wire n535bar;
  wire n536bar;
  wire n537bar;
  wire n538bar;
  wire n539bar;
  wire n540bar;
  wire n541bar;
  wire n542bar;
  wire n543bar;
  wire n544bar;
  wire n545bar;
  wire n546bar;
  wire n547bar;
  wire n548bar;
  wire n549bar;
  wire n550bar;
  wire n551bar;
  wire n552bar;
  wire n553bar;
  wire n554bar;
  wire n555bar;
  wire n556bar;
  wire n557bar;
  wire n558bar;
  wire n559bar;
  wire n560bar;
  wire n561bar;
  wire n562bar;
  wire n563bar;
  wire n564bar;
  wire n565bar;
  wire n566bar;
  wire n567bar;
  wire n568bar;
  wire n569bar;
  wire n570bar;
  wire n571bar;
  wire n572bar;
  wire n573bar;
  wire n574bar;
  wire n575bar;
  wire n576bar;
  wire n577bar;
  wire n578bar;
  wire n579bar;
  wire n580bar;
  wire n581bar;
  wire n582bar;
  wire n583bar;
  wire n584bar;
  wire n585bar;
  wire n586bar;
  wire n587bar;
  wire n588bar;
  wire n589bar;
  wire n590bar;
  wire n591bar;
  wire n592bar;
  wire n593bar;
  wire n594bar;
  wire n595bar;
  wire n596bar;
  wire n597bar;
  wire n598bar;
  wire n599bar;
  wire n600bar;
  wire n601bar;
  wire n602bar;
  wire n603bar;
  wire n604bar;
  wire n605bar;
  wire n606bar;
  wire n607bar;
  wire n608bar;
  wire n609bar;
  wire n610bar;
  wire n611bar;
  wire n612bar;
  wire n613bar;
  wire n614bar;
  wire n615bar;
  wire n616bar;
  wire n617bar;
  wire n618bar;
  wire n619bar;
  wire n620bar;
  wire n621bar;
  wire n622bar;
  wire n623bar;
  wire n624bar;
  wire n625bar;
  wire n626bar;
  wire n627bar;
  wire n628bar;
  wire n629bar;
  wire n630bar;
  wire n631bar;
  wire n632bar;
  wire n633bar;
  wire n634bar;
  wire n635bar;
  wire n636bar;
  wire n637bar;
  wire n638bar;
  wire n639bar;
  wire n640bar;
  wire n641bar;
  wire n642bar;
  wire n643bar;
  wire n644bar;
  wire n645bar;
  wire n646bar;
  wire n647bar;
  wire n648bar;
  wire n649bar;
  wire n650bar;
  wire n651bar;
  wire n652bar;
  wire n653bar;
  wire n654bar;
  wire n655bar;
  wire n656bar;
  wire n657bar;
  wire n658bar;
  wire n659bar;
  wire n660bar;
  wire n661bar;
  wire n662bar;
  wire n663bar;
  wire n664bar;
  wire n665bar;
  wire n666bar;
  wire n667bar;
  wire n668bar;
  wire n669bar;
  wire n670bar;
  wire n671bar;
  wire n672bar;
  wire n673bar;
  wire n674bar;
  wire n675bar;
  wire n676bar;
  wire n677bar;
  wire n678bar;
  wire n679bar;
  wire n680bar;
  wire n681bar;
  wire n682bar;
  wire n683bar;
  wire n684bar;
  wire n685bar;
  wire n686bar;
  wire n687bar;
  wire n688bar;
  wire n689bar;
  wire n690bar;
  wire n691bar;
  wire n692bar;
  wire n693bar;
  wire n694bar;
  wire n695bar;
  wire n696bar;
  wire n697bar;
  wire n698bar;
  wire n699bar;
  wire n700bar;
  wire n701bar;
  wire n702bar;
  wire n703bar;
  wire n704bar;
  wire n705bar;
  wire n706bar;
  wire n707bar;
  wire n708bar;
  wire n709bar;
  wire n710bar;
  wire n711bar;
  wire n712bar;
  wire n713bar;
  wire n714bar;
  wire n715bar;
  wire n716bar;
  wire n717bar;
  wire n718bar;
  wire n719bar;
  wire n720bar;
  wire n721bar;
  wire n722bar;
  wire n723bar;
  wire n724bar;
  wire n725bar;
  wire n726bar;
  wire n727bar;
  wire n728bar;
  wire n729bar;
  wire n730bar;
  wire n731bar;
  wire n732bar;
  wire n733bar;
  wire n734bar;
  wire n735bar;
  wire n736bar;
  wire n737bar;
  wire n738bar;
  wire n739bar;
  wire n740bar;
  wire n741bar;
  wire n742bar;
  wire n743bar;
  wire n744bar;
  wire n745bar;
  wire n746bar;
  wire n747bar;
  wire n748bar;
  wire n749bar;
  wire n750bar;
  wire n751bar;
  wire n752bar;
  wire n753bar;
  wire n754bar;
  wire n755bar;
  wire n756bar;
  wire n757bar;
  wire n758bar;
  wire n759bar;
  wire n760bar;
  wire n761bar;
  wire n762bar;
  wire n763bar;
  wire n764bar;
  wire n765bar;
  wire n766bar;
  wire n767bar;
  wire n768bar;
  wire n769bar;
  wire n770bar;
  wire n771bar;
  wire n772bar;
  wire n773bar;
  wire n774bar;
  wire n775bar;
  wire n776bar;
  wire n777bar;
  wire n778bar;
  wire n779bar;
  wire n780bar;
  wire n781bar;
  wire n782bar;
  wire n783bar;
  wire n784bar;
  wire n785bar;
  wire n786bar;
  wire n787bar;
  wire n788bar;
  wire n789bar;
  wire n790bar;
  wire n791bar;
  wire n792bar;
  wire n793bar;
  wire n794bar;
  wire n795bar;
  wire n796bar;
  wire n797bar;
  wire n798bar;
  wire n799bar;
  wire n800bar;
  wire n801bar;
  wire n802bar;
  wire n803bar;
  wire n804bar;
  wire n805bar;
  wire n806bar;
  wire n807bar;
  wire n808bar;
  wire n809bar;
  wire n810bar;
  wire n811bar;
  wire n812bar;
  wire n813bar;
  wire n814bar;
  wire n815bar;
  wire n816bar;
  wire n817bar;
  wire n818bar;
  wire n819bar;
  wire n820bar;
  wire n821bar;
  wire n822bar;
  wire n823bar;
  wire n824bar;
  wire n825bar;
  wire n826bar;
  wire n827bar;
  wire n828bar;
  wire n829bar;
  wire n830bar;
  wire n831bar;
  wire n832bar;
  wire n833bar;
  wire n834bar;
  wire n835bar;
  wire n836bar;
  wire n837bar;
  wire n838bar;
  wire n839bar;
  wire n840bar;
  wire n841bar;
  wire n842bar;
  wire n843bar;
  wire n844bar;
  wire n845bar;
  wire n846bar;
  wire n847bar;
  wire n848bar;
  wire n849bar;
  wire n850bar;
  wire n851bar;
  wire n852bar;
  wire n853bar;
  wire n854bar;
  wire n855bar;
  wire n856bar;
  wire n857bar;
  wire n858bar;
  wire n859bar;
  wire n860bar;
  wire n861bar;
  wire n862bar;
  wire n863bar;
  wire n864bar;
  wire n865bar;
  wire n866bar;
  wire n867bar;
  wire n868bar;
  wire n869bar;
  wire n870bar;
  wire n871bar;
  wire n872bar;
  wire n873bar;
  wire n874bar;
  wire n875bar;
  wire n876bar;
  wire n877bar;
  wire n878bar;
  wire n879bar;
  wire n880bar;
  wire n881bar;
  wire n882bar;
  wire n883bar;
  wire n884bar;
  wire n885bar;
  wire n886bar;
  wire n887bar;
  wire n888bar;
  wire n889bar;
  wire n890bar;
  wire n891bar;
  wire n892bar;
  wire n893bar;
  wire n894bar;
  wire n895bar;
  wire n896bar;
  wire n897bar;
  wire n898bar;
  wire n899bar;
  wire n900bar;
  wire n901bar;
  wire n902bar;
  wire n903bar;
  wire n904bar;
  wire n905bar;
  wire n906bar;
  wire n907bar;
  wire n908bar;
  wire n909bar;
  wire n910bar;
  wire n911bar;
  wire n912bar;
  wire n913bar;
  wire n914bar;
  wire n915bar;
  wire n916bar;
  wire n917bar;
  wire n918bar;
  wire n919bar;
  wire n920bar;
  wire n921bar;
  wire n922bar;
  wire n923bar;
  wire n924bar;
  wire n925bar;
  wire n926bar;
  wire n927bar;
  wire n928bar;
  wire n929bar;
  wire n930bar;
  wire n931bar;
  wire n932bar;
  wire n933bar;
  wire n934bar;
  wire n935bar;
  wire n936bar;
  wire n937bar;
  wire n938bar;
  wire n939bar;
  wire n940bar;
  wire n941bar;
  wire n942bar;
  wire n943bar;
  wire n944bar;
  wire n945bar;
  wire n946bar;
  wire n947bar;
  wire n948bar;
  wire n949bar;
  wire n950bar;
  wire n951bar;
  wire n952bar;
  wire n953bar;
  wire n954bar;
  wire n955bar;
  wire n956bar;
  wire n957bar;
  wire n958bar;
  wire n959bar;
  wire n960bar;
  wire n961bar;
  wire n962bar;
  wire n963bar;
  wire n964bar;
  wire n965bar;
  wire n966bar;
  wire n967bar;
  wire n968bar;
  wire n969bar;
  wire n970bar;
  wire n971bar;
  wire n972bar;
//wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];
  assign in_81bar = inbar[81];
  assign in_80bar = inbar[80];
  assign in_79bar = inbar[79];
  assign in_78bar = inbar[78];
  assign in_77bar = inbar[77];
  assign in_76bar = inbar[76];
  assign in_75bar = inbar[75];
  assign in_74bar = inbar[74];
  assign in_73bar = inbar[73];
  assign in_72bar = inbar[72];
  assign in_71bar = inbar[71];
  assign in_70bar = inbar[70];
  assign in_69bar = inbar[69];
  assign in_68bar = inbar[68];
  assign in_67bar = inbar[67];
  assign in_66bar = inbar[66];
  assign in_65bar = inbar[65];
  assign in_64bar = inbar[64];
  assign in_63bar = inbar[63];
  assign in_62bar = inbar[62];
  assign in_61bar = inbar[61];
  assign in_60bar = inbar[60];
  assign in_59bar = inbar[59];
  assign in_58bar = inbar[58];
  assign in_57bar = inbar[57];
  assign in_56bar = inbar[56];
  assign in_55bar = inbar[55];
  assign in_54bar = inbar[54];
  assign in_53bar = inbar[53];
  assign in_52bar = inbar[52];
  assign in_51bar = inbar[51];
  assign in_50bar = inbar[50];
  assign in_49bar = inbar[49];
  assign in_48bar = inbar[48];
  assign in_47bar = inbar[47];
  assign in_46bar = inbar[46];
  assign in_45bar = inbar[45];
  assign in_44bar = inbar[44];
  assign in_43bar = inbar[43];
  assign in_42bar = inbar[42];
  assign in_41bar = inbar[41];
  assign in_40bar = inbar[40];
  assign in_39bar = inbar[39];
  assign in_38bar = inbar[38];
  assign in_37bar = inbar[37];
  assign in_36bar = inbar[36];
  assign in_35bar = inbar[35];
  assign in_34bar = inbar[34];
  assign in_33bar = inbar[33];
  assign in_32bar = inbar[32];
  assign in_31bar = inbar[31];
  assign in_30bar = inbar[30];
  assign in_29bar = inbar[29];
  assign in_28bar = inbar[28];
  assign in_27bar = inbar[27];
  assign in_26bar = inbar[26];
  assign in_25bar = inbar[25];
  assign in_24bar = inbar[24];
  assign in_23bar = inbar[23];
  assign in_22bar = inbar[22];
  assign in_21bar = inbar[21];
  assign in_20bar = inbar[20];
  assign in_19bar = inbar[19];
  assign in_18bar = inbar[18];
  assign in_17bar = inbar[17];
  assign in_16bar = inbar[16];
  assign in_15bar = inbar[15];
  assign in_14bar = inbar[14];
  assign in_13bar = inbar[13];
  assign in_12bar = inbar[12];
  assign in_11bar = inbar[11];
  assign in_10bar = inbar[10];
  assign in_9bar = inbar[9];
  assign in_8bar = inbar[8];
  assign in_7bar = inbar[7];
  assign in_6bar = inbar[6];
  assign in_5bar = inbar[5];
  assign in_4bar = inbar[4];
  assign in_3bar = inbar[3];
  assign in_2bar = inbar[2];
  assign in_1bar = inbar[1];
  assign in_0bar = inbar[0];
//assign_done

  OR2_X1 U1 ( .A1(n972), .A2(n971), .ZN(out[7]) );
  AND2_X1 U1bar ( .A1(n972bar), .A2(n971bar), .ZN(outbar[7]) );
  OR2_X1 U2 ( .A1(n970), .A2(n969), .ZN(n971) );
  AND2_X1 U2bar ( .A1(n970bar), .A2(n969bar), .ZN(n971bar) );
  OR2_X1 U3 ( .A1(n968), .A2(n967), .ZN(n969) );
  AND2_X1 U3bar ( .A1(n968bar), .A2(n967bar), .ZN(n969bar) );
  OR2_X1 U4 ( .A1(n966), .A2(n965), .ZN(n967) );
  AND2_X1 U4bar ( .A1(n966bar), .A2(n965bar), .ZN(n967bar) );
  OR2_X1 U5 ( .A1(n964), .A2(n963), .ZN(n968) );
  AND2_X1 U5bar ( .A1(n964bar), .A2(n963bar), .ZN(n968bar) );
  OR2_X1 U6 ( .A1(in[116]), .A2(n962), .ZN(n963) );
  AND2_X1 U6bar ( .A1(inbar[116]), .A2(n962bar), .ZN(n963bar) );
  OR2_X1 U7 ( .A1(n961), .A2(n960), .ZN(n970) );
  AND2_X1 U7bar ( .A1(n961bar), .A2(n960bar), .ZN(n970bar) );
  OR2_X1 U8 ( .A1(in[150]), .A2(in[127]), .ZN(n960) );
  AND2_X1 U8bar ( .A1(inbar[150]), .A2(inbar[127]), .ZN(n960bar) );
  OR2_X1 U9 ( .A1(in[160]), .A2(n959), .ZN(n961) );
  AND2_X1 U9bar ( .A1(inbar[160]), .A2(n959bar), .ZN(n961bar) );
  OR2_X1 U10 ( .A1(in[252]), .A2(in[168]), .ZN(n959) );
  AND2_X1 U10bar ( .A1(inbar[252]), .A2(inbar[168]), .ZN(n959bar) );
  OR2_X1 U11 ( .A1(n958), .A2(n957), .ZN(n972) );
  AND2_X1 U11bar ( .A1(n958bar), .A2(n957bar), .ZN(n972bar) );
  OR2_X1 U12 ( .A1(n956), .A2(n955), .ZN(n957) );
  AND2_X1 U12bar ( .A1(n956bar), .A2(n955bar), .ZN(n957bar) );
  OR2_X1 U13 ( .A1(in_17), .A2(in[96]), .ZN(n955) );
  AND2_X1 U13bar ( .A1(in_17bar), .A2(inbar[96]), .ZN(n955bar) );
  OR2_X1 U14 ( .A1(in_23), .A2(n954), .ZN(n956) );
  AND2_X1 U14bar ( .A1(in_23bar), .A2(n954bar), .ZN(n956bar) );
  OR2_X1 U15 ( .A1(in_31), .A2(in_26), .ZN(n954) );
  AND2_X1 U15bar ( .A1(in_31bar), .A2(in_26bar), .ZN(n954bar) );
  OR2_X1 U16 ( .A1(n953), .A2(n952), .ZN(n958) );
  AND2_X1 U16bar ( .A1(n953bar), .A2(n952bar), .ZN(n958bar) );
  OR2_X1 U17 ( .A1(in_58), .A2(in_4), .ZN(n952) );
  AND2_X1 U17bar ( .A1(in_58bar), .A2(in_4bar), .ZN(n952bar) );
  OR2_X1 U18 ( .A1(in_59), .A2(n951), .ZN(n953) );
  AND2_X1 U18bar ( .A1(in_59bar), .A2(n951bar), .ZN(n953bar) );
  OR2_X1 U19 ( .A1(in_71), .A2(in_62), .ZN(n951) );
  AND2_X1 U19bar ( .A1(in_71bar), .A2(in_62bar), .ZN(n951bar) );
  OR2_X1 U20 ( .A1(n950), .A2(n949), .ZN(out[6]) );
  AND2_X1 U20bar ( .A1(n950bar), .A2(n949bar), .ZN(outbar[6]) );
  OR2_X1 U21 ( .A1(n948), .A2(n947), .ZN(n949) );
  AND2_X1 U21bar ( .A1(n948bar), .A2(n947bar), .ZN(n949bar) );
  OR2_X1 U22 ( .A1(n946), .A2(n945), .ZN(n947) );
  AND2_X1 U22bar ( .A1(n946bar), .A2(n945bar), .ZN(n947bar) );
  OR2_X1 U23 ( .A1(n944), .A2(n943), .ZN(n945) );
  AND2_X1 U23bar ( .A1(n944bar), .A2(n943bar), .ZN(n945bar) );
  OR2_X1 U24 ( .A1(n942), .A2(n941), .ZN(n946) );
  AND2_X1 U24bar ( .A1(n942bar), .A2(n941bar), .ZN(n946bar) );
  OR2_X1 U25 ( .A1(in[101]), .A2(n940), .ZN(n941) );
  AND2_X1 U25bar ( .A1(inbar[101]), .A2(n940bar), .ZN(n941bar) );
  OR2_X1 U26 ( .A1(n939), .A2(n938), .ZN(n948) );
  AND2_X1 U26bar ( .A1(n939bar), .A2(n938bar), .ZN(n948bar) );
  OR2_X1 U27 ( .A1(in[114]), .A2(in[104]), .ZN(n938) );
  AND2_X1 U27bar ( .A1(inbar[114]), .A2(inbar[104]), .ZN(n938bar) );
  OR2_X1 U28 ( .A1(in[128]), .A2(n937), .ZN(n939) );
  AND2_X1 U28bar ( .A1(inbar[128]), .A2(n937bar), .ZN(n939bar) );
  OR2_X1 U29 ( .A1(in[136]), .A2(in[134]), .ZN(n937) );
  AND2_X1 U29bar ( .A1(inbar[136]), .A2(inbar[134]), .ZN(n937bar) );
  OR2_X1 U30 ( .A1(n936), .A2(n935), .ZN(n950) );
  AND2_X1 U30bar ( .A1(n936bar), .A2(n935bar), .ZN(n950bar) );
  OR2_X1 U31 ( .A1(n934), .A2(n933), .ZN(n935) );
  AND2_X1 U31bar ( .A1(n934bar), .A2(n933bar), .ZN(n935bar) );
  OR2_X1 U32 ( .A1(in[177]), .A2(in[164]), .ZN(n933) );
  AND2_X1 U32bar ( .A1(inbar[177]), .A2(inbar[164]), .ZN(n933bar) );
  OR2_X1 U33 ( .A1(in[212]), .A2(n932), .ZN(n934) );
  AND2_X1 U33bar ( .A1(inbar[212]), .A2(n932bar), .ZN(n934bar) );
  OR2_X1 U34 ( .A1(in[248]), .A2(in[221]), .ZN(n932) );
  AND2_X1 U34bar ( .A1(inbar[248]), .A2(inbar[221]), .ZN(n932bar) );
  OR2_X1 U35 ( .A1(n931), .A2(n930), .ZN(n936) );
  AND2_X1 U35bar ( .A1(n931bar), .A2(n930bar), .ZN(n936bar) );
  OR2_X1 U36 ( .A1(in_18), .A2(in[93]), .ZN(n930) );
  AND2_X1 U36bar ( .A1(in_18bar), .A2(inbar[93]), .ZN(n930bar) );
  OR2_X1 U37 ( .A1(in_31), .A2(n929), .ZN(n931) );
  AND2_X1 U37bar ( .A1(in_31bar), .A2(n929bar), .ZN(n931bar) );
  OR2_X1 U38 ( .A1(in_7), .A2(in_39), .ZN(n929) );
  AND2_X1 U38bar ( .A1(in_7bar), .A2(in_39bar), .ZN(n929bar) );
  OR2_X1 U39 ( .A1(n928), .A2(n927), .ZN(out[5]) );
  AND2_X1 U39bar ( .A1(n928bar), .A2(n927bar), .ZN(outbar[5]) );
  OR2_X1 U40 ( .A1(n926), .A2(n925), .ZN(n927) );
  AND2_X1 U40bar ( .A1(n926bar), .A2(n925bar), .ZN(n927bar) );
  OR2_X1 U41 ( .A1(n924), .A2(n923), .ZN(n925) );
  AND2_X1 U41bar ( .A1(n924bar), .A2(n923bar), .ZN(n925bar) );
  OR2_X1 U42 ( .A1(n922), .A2(n921), .ZN(n923) );
  AND2_X1 U42bar ( .A1(n922bar), .A2(n921bar), .ZN(n923bar) );
  OR2_X1 U43 ( .A1(n940), .A2(n920), .ZN(n924) );
  AND2_X1 U43bar ( .A1(n940bar), .A2(n920bar), .ZN(n924bar) );
  OR2_X1 U44 ( .A1(in[111]), .A2(n919), .ZN(n920) );
  AND2_X1 U44bar ( .A1(inbar[111]), .A2(n919bar), .ZN(n920bar) );
  OR2_X1 U45 ( .A1(n918), .A2(n917), .ZN(n940) );
  AND2_X1 U45bar ( .A1(n918bar), .A2(n917bar), .ZN(n940bar) );
  OR2_X1 U46 ( .A1(n916), .A2(n915), .ZN(n917) );
  AND2_X1 U46bar ( .A1(n916bar), .A2(n915bar), .ZN(n917bar) );
  OR2_X1 U47 ( .A1(n914), .A2(n913), .ZN(n915) );
  AND2_X1 U47bar ( .A1(n914bar), .A2(n913bar), .ZN(n915bar) );
  OR2_X1 U48 ( .A1(in[140]), .A2(in[131]), .ZN(n913) );
  AND2_X1 U48bar ( .A1(inbar[140]), .A2(inbar[131]), .ZN(n913bar) );
  OR2_X1 U49 ( .A1(in[160]), .A2(in[144]), .ZN(n914) );
  AND2_X1 U49bar ( .A1(inbar[160]), .A2(inbar[144]), .ZN(n914bar) );
  OR2_X1 U50 ( .A1(n912), .A2(n911), .ZN(n916) );
  AND2_X1 U50bar ( .A1(n912bar), .A2(n911bar), .ZN(n916bar) );
  OR2_X1 U51 ( .A1(in[179]), .A2(in[174]), .ZN(n911) );
  AND2_X1 U51bar ( .A1(inbar[179]), .A2(inbar[174]), .ZN(n911bar) );
  OR2_X1 U52 ( .A1(in[188]), .A2(in[184]), .ZN(n912) );
  AND2_X1 U52bar ( .A1(inbar[188]), .A2(inbar[184]), .ZN(n912bar) );
  OR2_X1 U53 ( .A1(n910), .A2(n909), .ZN(n918) );
  AND2_X1 U53bar ( .A1(n910bar), .A2(n909bar), .ZN(n918bar) );
  OR2_X1 U54 ( .A1(n908), .A2(n907), .ZN(n909) );
  AND2_X1 U54bar ( .A1(n908bar), .A2(n907bar), .ZN(n909bar) );
  OR2_X1 U55 ( .A1(in[216]), .A2(in[200]), .ZN(n907) );
  AND2_X1 U55bar ( .A1(inbar[216]), .A2(inbar[200]), .ZN(n907bar) );
  OR2_X1 U56 ( .A1(in[228]), .A2(in[224]), .ZN(n908) );
  AND2_X1 U56bar ( .A1(inbar[228]), .A2(inbar[224]), .ZN(n908bar) );
  OR2_X1 U57 ( .A1(n906), .A2(n905), .ZN(n910) );
  AND2_X1 U57bar ( .A1(n906bar), .A2(n905bar), .ZN(n910bar) );
  OR2_X1 U58 ( .A1(in[247]), .A2(in[235]), .ZN(n905) );
  AND2_X1 U58bar ( .A1(inbar[247]), .A2(inbar[235]), .ZN(n905bar) );
  OR2_X1 U59 ( .A1(in_42), .A2(in[83]), .ZN(n906) );
  AND2_X1 U59bar ( .A1(in_42bar), .A2(inbar[83]), .ZN(n906bar) );
  OR2_X1 U60 ( .A1(n904), .A2(n903), .ZN(n926) );
  AND2_X1 U60bar ( .A1(n904bar), .A2(n903bar), .ZN(n926bar) );
  OR2_X1 U61 ( .A1(in[166]), .A2(in[123]), .ZN(n903) );
  AND2_X1 U61bar ( .A1(inbar[166]), .A2(inbar[123]), .ZN(n903bar) );
  OR2_X1 U62 ( .A1(in[170]), .A2(n902), .ZN(n904) );
  AND2_X1 U62bar ( .A1(inbar[170]), .A2(n902bar), .ZN(n904bar) );
  OR2_X1 U63 ( .A1(in[194]), .A2(in[183]), .ZN(n902) );
  AND2_X1 U63bar ( .A1(inbar[194]), .A2(inbar[183]), .ZN(n902bar) );
  OR2_X1 U64 ( .A1(n901), .A2(n900), .ZN(n928) );
  AND2_X1 U64bar ( .A1(n901bar), .A2(n900bar), .ZN(n928bar) );
  OR2_X1 U65 ( .A1(n899), .A2(n898), .ZN(n900) );
  AND2_X1 U65bar ( .A1(n899bar), .A2(n898bar), .ZN(n900bar) );
  OR2_X1 U66 ( .A1(in[241]), .A2(in[238]), .ZN(n898) );
  AND2_X1 U66bar ( .A1(inbar[241]), .A2(inbar[238]), .ZN(n898bar) );
  OR2_X1 U67 ( .A1(in[250]), .A2(n897), .ZN(n899) );
  AND2_X1 U67bar ( .A1(inbar[250]), .A2(n897bar), .ZN(n899bar) );
  OR2_X1 U68 ( .A1(in_24), .A2(in[84]), .ZN(n897) );
  AND2_X1 U68bar ( .A1(in_24bar), .A2(inbar[84]), .ZN(n897bar) );
  OR2_X1 U69 ( .A1(n896), .A2(n895), .ZN(n901) );
  AND2_X1 U69bar ( .A1(n896bar), .A2(n895bar), .ZN(n901bar) );
  OR2_X1 U70 ( .A1(in_41), .A2(in_29), .ZN(n895) );
  AND2_X1 U70bar ( .A1(in_41bar), .A2(in_29bar), .ZN(n895bar) );
  OR2_X1 U71 ( .A1(in_66), .A2(n894), .ZN(n896) );
  AND2_X1 U71bar ( .A1(in_66bar), .A2(n894bar), .ZN(n896bar) );
  OR2_X1 U72 ( .A1(in_76), .A2(in_71), .ZN(n894) );
  AND2_X1 U72bar ( .A1(in_76bar), .A2(in_71bar), .ZN(n894bar) );
  OR2_X1 U73 ( .A1(n893), .A2(n892), .ZN(out[4]) );
  AND2_X1 U73bar ( .A1(n893bar), .A2(n892bar), .ZN(outbar[4]) );
  OR2_X1 U74 ( .A1(n891), .A2(n890), .ZN(n892) );
  AND2_X1 U74bar ( .A1(n891bar), .A2(n890bar), .ZN(n892bar) );
  OR2_X1 U75 ( .A1(n889), .A2(n888), .ZN(n890) );
  AND2_X1 U75bar ( .A1(n889bar), .A2(n888bar), .ZN(n890bar) );
  OR2_X1 U76 ( .A1(n922), .A2(n887), .ZN(n888) );
  AND2_X1 U76bar ( .A1(n922bar), .A2(n887bar), .ZN(n888bar) );
  OR2_X1 U77 ( .A1(n886), .A2(n885), .ZN(n922) );
  AND2_X1 U77bar ( .A1(n886bar), .A2(n885bar), .ZN(n922bar) );
  OR2_X1 U78 ( .A1(n884), .A2(n883), .ZN(n885) );
  AND2_X1 U78bar ( .A1(n884bar), .A2(n883bar), .ZN(n885bar) );
  OR2_X1 U79 ( .A1(n882), .A2(n881), .ZN(n883) );
  AND2_X1 U79bar ( .A1(n882bar), .A2(n881bar), .ZN(n883bar) );
  OR2_X1 U80 ( .A1(in[118]), .A2(in[109]), .ZN(n881) );
  AND2_X1 U80bar ( .A1(inbar[118]), .A2(inbar[109]), .ZN(n881bar) );
  OR2_X1 U81 ( .A1(in[139]), .A2(in[120]), .ZN(n882) );
  AND2_X1 U81bar ( .A1(inbar[139]), .A2(inbar[120]), .ZN(n882bar) );
  OR2_X1 U82 ( .A1(n880), .A2(n879), .ZN(n884) );
  AND2_X1 U82bar ( .A1(n880bar), .A2(n879bar), .ZN(n884bar) );
  OR2_X1 U83 ( .A1(in[198]), .A2(in[154]), .ZN(n879) );
  AND2_X1 U83bar ( .A1(inbar[198]), .A2(inbar[154]), .ZN(n879bar) );
  OR2_X1 U84 ( .A1(in[210]), .A2(in[205]), .ZN(n880) );
  AND2_X1 U84bar ( .A1(inbar[210]), .A2(inbar[205]), .ZN(n880bar) );
  OR2_X1 U85 ( .A1(n878), .A2(n877), .ZN(n886) );
  AND2_X1 U85bar ( .A1(n878bar), .A2(n877bar), .ZN(n886bar) );
  OR2_X1 U86 ( .A1(n876), .A2(n875), .ZN(n877) );
  AND2_X1 U86bar ( .A1(n876bar), .A2(n875bar), .ZN(n877bar) );
  OR2_X1 U87 ( .A1(in[219]), .A2(in[217]), .ZN(n875) );
  AND2_X1 U87bar ( .A1(inbar[219]), .A2(inbar[217]), .ZN(n875bar) );
  OR2_X1 U88 ( .A1(in[86]), .A2(in[252]), .ZN(n876) );
  AND2_X1 U88bar ( .A1(inbar[86]), .A2(inbar[252]), .ZN(n876bar) );
  OR2_X1 U89 ( .A1(n874), .A2(n873), .ZN(n878) );
  AND2_X1 U89bar ( .A1(n874bar), .A2(n873bar), .ZN(n878bar) );
  OR2_X1 U90 ( .A1(in_40), .A2(in[91]), .ZN(n873) );
  AND2_X1 U90bar ( .A1(in_40bar), .A2(inbar[91]), .ZN(n873bar) );
  OR2_X1 U91 ( .A1(in_8), .A2(in_46), .ZN(n874) );
  AND2_X1 U91bar ( .A1(in_8bar), .A2(in_46bar), .ZN(n874bar) );
  OR2_X1 U92 ( .A1(n872), .A2(n871), .ZN(n889) );
  AND2_X1 U92bar ( .A1(n872bar), .A2(n871bar), .ZN(n889bar) );
  OR2_X1 U93 ( .A1(in[117]), .A2(n943), .ZN(n871) );
  AND2_X1 U93bar ( .A1(inbar[117]), .A2(n943bar), .ZN(n871bar) );
  OR2_X1 U94 ( .A1(n870), .A2(n869), .ZN(n943) );
  AND2_X1 U94bar ( .A1(n870bar), .A2(n869bar), .ZN(n943bar) );
  OR2_X1 U95 ( .A1(n868), .A2(n867), .ZN(n869) );
  AND2_X1 U95bar ( .A1(n868bar), .A2(n867bar), .ZN(n869bar) );
  OR2_X1 U96 ( .A1(n866), .A2(n865), .ZN(n867) );
  AND2_X1 U96bar ( .A1(n866bar), .A2(n865bar), .ZN(n867bar) );
  OR2_X1 U97 ( .A1(n864), .A2(n863), .ZN(n865) );
  AND2_X1 U97bar ( .A1(n864bar), .A2(n863bar), .ZN(n865bar) );
  OR2_X1 U98 ( .A1(in[108]), .A2(n919), .ZN(n866) );
  AND2_X1 U98bar ( .A1(inbar[108]), .A2(n919bar), .ZN(n866bar) );
  OR2_X1 U99 ( .A1(n862), .A2(n861), .ZN(n919) );
  AND2_X1 U99bar ( .A1(n862bar), .A2(n861bar), .ZN(n919bar) );
  OR2_X1 U100 ( .A1(n860), .A2(n859), .ZN(n861) );
  AND2_X1 U100bar ( .A1(n860bar), .A2(n859bar), .ZN(n861bar) );
  OR2_X1 U101 ( .A1(n858), .A2(n857), .ZN(n859) );
  AND2_X1 U101bar ( .A1(n858bar), .A2(n857bar), .ZN(n859bar) );
  OR2_X1 U102 ( .A1(in[119]), .A2(in[105]), .ZN(n857) );
  AND2_X1 U102bar ( .A1(inbar[119]), .A2(inbar[105]), .ZN(n857bar) );
  OR2_X1 U103 ( .A1(in[186]), .A2(in[175]), .ZN(n858) );
  AND2_X1 U103bar ( .A1(inbar[186]), .A2(inbar[175]), .ZN(n858bar) );
  OR2_X1 U104 ( .A1(n856), .A2(n855), .ZN(n860) );
  AND2_X1 U104bar ( .A1(n856bar), .A2(n855bar), .ZN(n860bar) );
  OR2_X1 U105 ( .A1(in[202]), .A2(in[193]), .ZN(n855) );
  AND2_X1 U105bar ( .A1(inbar[202]), .A2(inbar[193]), .ZN(n855bar) );
  OR2_X1 U106 ( .A1(in[225]), .A2(in[208]), .ZN(n856) );
  AND2_X1 U106bar ( .A1(inbar[225]), .A2(inbar[208]), .ZN(n856bar) );
  OR2_X1 U107 ( .A1(n854), .A2(n853), .ZN(n862) );
  AND2_X1 U107bar ( .A1(n854bar), .A2(n853bar), .ZN(n862bar) );
  OR2_X1 U108 ( .A1(n852), .A2(n851), .ZN(n853) );
  AND2_X1 U108bar ( .A1(n852bar), .A2(n851bar), .ZN(n853bar) );
  OR2_X1 U109 ( .A1(in_1), .A2(in[85]), .ZN(n851) );
  AND2_X1 U109bar ( .A1(in_1bar), .A2(inbar[85]), .ZN(n851bar) );
  OR2_X1 U110 ( .A1(in_23), .A2(in_19), .ZN(n852) );
  AND2_X1 U110bar ( .A1(in_23bar), .A2(in_19bar), .ZN(n852bar) );
  OR2_X1 U111 ( .A1(n850), .A2(n849), .ZN(n854) );
  AND2_X1 U111bar ( .A1(n850bar), .A2(n849bar), .ZN(n854bar) );
  OR2_X1 U112 ( .A1(in_43), .A2(in_33), .ZN(n849) );
  AND2_X1 U112bar ( .A1(in_43bar), .A2(in_33bar), .ZN(n849bar) );
  OR2_X1 U113 ( .A1(in_63), .A2(in_44), .ZN(n850) );
  AND2_X1 U113bar ( .A1(in_63bar), .A2(in_44bar), .ZN(n850bar) );
  OR2_X1 U114 ( .A1(n848), .A2(n847), .ZN(n868) );
  AND2_X1 U114bar ( .A1(n848bar), .A2(n847bar), .ZN(n868bar) );
  OR2_X1 U115 ( .A1(in[141]), .A2(in[112]), .ZN(n847) );
  AND2_X1 U115bar ( .A1(inbar[141]), .A2(inbar[112]), .ZN(n847bar) );
  OR2_X1 U116 ( .A1(in[147]), .A2(n846), .ZN(n848) );
  AND2_X1 U116bar ( .A1(inbar[147]), .A2(n846bar), .ZN(n848bar) );
  OR2_X1 U117 ( .A1(in[181]), .A2(in[167]), .ZN(n846) );
  AND2_X1 U117bar ( .A1(inbar[181]), .A2(inbar[167]), .ZN(n846bar) );
  OR2_X1 U118 ( .A1(n845), .A2(n844), .ZN(n870) );
  AND2_X1 U118bar ( .A1(n845bar), .A2(n844bar), .ZN(n870bar) );
  OR2_X1 U119 ( .A1(n843), .A2(n842), .ZN(n844) );
  AND2_X1 U119bar ( .A1(n843bar), .A2(n842bar), .ZN(n844bar) );
  OR2_X1 U120 ( .A1(in[229]), .A2(in[201]), .ZN(n842) );
  AND2_X1 U120bar ( .A1(inbar[229]), .A2(inbar[201]), .ZN(n842bar) );
  OR2_X1 U121 ( .A1(in[237]), .A2(n841), .ZN(n843) );
  AND2_X1 U121bar ( .A1(inbar[237]), .A2(n841bar), .ZN(n843bar) );
  OR2_X1 U122 ( .A1(in[94]), .A2(in[253]), .ZN(n841) );
  AND2_X1 U122bar ( .A1(inbar[94]), .A2(inbar[253]), .ZN(n841bar) );
  OR2_X1 U123 ( .A1(n840), .A2(n839), .ZN(n845) );
  AND2_X1 U123bar ( .A1(n840bar), .A2(n839bar), .ZN(n845bar) );
  OR2_X1 U124 ( .A1(in_21), .A2(in[96]), .ZN(n839) );
  AND2_X1 U124bar ( .A1(in_21bar), .A2(inbar[96]), .ZN(n839bar) );
  OR2_X1 U125 ( .A1(in_25), .A2(n838), .ZN(n840) );
  AND2_X1 U125bar ( .A1(in_25bar), .A2(n838bar), .ZN(n840bar) );
  OR2_X1 U126 ( .A1(in_81), .A2(in_45), .ZN(n838) );
  AND2_X1 U126bar ( .A1(in_81bar), .A2(in_45bar), .ZN(n838bar) );
  OR2_X1 U127 ( .A1(n837), .A2(n836), .ZN(n891) );
  AND2_X1 U127bar ( .A1(n837bar), .A2(n836bar), .ZN(n891bar) );
  OR2_X1 U128 ( .A1(in[142]), .A2(in[124]), .ZN(n836) );
  AND2_X1 U128bar ( .A1(inbar[142]), .A2(inbar[124]), .ZN(n836bar) );
  OR2_X1 U129 ( .A1(in[150]), .A2(n835), .ZN(n837) );
  AND2_X1 U129bar ( .A1(inbar[150]), .A2(n835bar), .ZN(n837bar) );
  OR2_X1 U130 ( .A1(in[172]), .A2(in[155]), .ZN(n835) );
  AND2_X1 U130bar ( .A1(inbar[172]), .A2(inbar[155]), .ZN(n835bar) );
  OR2_X1 U131 ( .A1(n834), .A2(n833), .ZN(n893) );
  AND2_X1 U131bar ( .A1(n834bar), .A2(n833bar), .ZN(n893bar) );
  OR2_X1 U132 ( .A1(n832), .A2(n831), .ZN(n833) );
  AND2_X1 U132bar ( .A1(n832bar), .A2(n831bar), .ZN(n833bar) );
  OR2_X1 U133 ( .A1(in[196]), .A2(in[173]), .ZN(n831) );
  AND2_X1 U133bar ( .A1(inbar[196]), .A2(inbar[173]), .ZN(n831bar) );
  OR2_X1 U134 ( .A1(in[222]), .A2(n830), .ZN(n832) );
  AND2_X1 U134bar ( .A1(inbar[222]), .A2(n830bar), .ZN(n832bar) );
  OR2_X1 U135 ( .A1(in[227]), .A2(in[226]), .ZN(n830) );
  AND2_X1 U135bar ( .A1(inbar[227]), .A2(inbar[226]), .ZN(n830bar) );
  OR2_X1 U136 ( .A1(n829), .A2(n828), .ZN(n834) );
  AND2_X1 U136bar ( .A1(n829bar), .A2(n828bar), .ZN(n834bar) );
  OR2_X1 U137 ( .A1(in[249]), .A2(in[231]), .ZN(n828) );
  AND2_X1 U137bar ( .A1(inbar[249]), .A2(inbar[231]), .ZN(n828bar) );
  OR2_X1 U138 ( .A1(in_28), .A2(n827), .ZN(n829) );
  AND2_X1 U138bar ( .A1(in_28bar), .A2(n827bar), .ZN(n829bar) );
  OR2_X1 U139 ( .A1(in_52), .A2(in_47), .ZN(n827) );
  AND2_X1 U139bar ( .A1(in_52bar), .A2(in_47bar), .ZN(n827bar) );
  OR2_X1 U140 ( .A1(n826), .A2(n825), .ZN(out[3]) );
  AND2_X1 U140bar ( .A1(n826bar), .A2(n825bar), .ZN(outbar[3]) );
  OR2_X1 U141 ( .A1(n824), .A2(n823), .ZN(n825) );
  AND2_X1 U141bar ( .A1(n824bar), .A2(n823bar), .ZN(n825bar) );
  OR2_X1 U142 ( .A1(n822), .A2(n821), .ZN(n823) );
  AND2_X1 U142bar ( .A1(n822bar), .A2(n821bar), .ZN(n823bar) );
  OR2_X1 U143 ( .A1(n820), .A2(n819), .ZN(n821) );
  AND2_X1 U143bar ( .A1(n820bar), .A2(n819bar), .ZN(n821bar) );
  OR2_X1 U144 ( .A1(n964), .A2(n818), .ZN(n822) );
  AND2_X1 U144bar ( .A1(n964bar), .A2(n818bar), .ZN(n822bar) );
  OR2_X1 U145 ( .A1(in[118]), .A2(n817), .ZN(n818) );
  AND2_X1 U145bar ( .A1(inbar[118]), .A2(n817bar), .ZN(n818bar) );
  OR2_X1 U146 ( .A1(n816), .A2(n815), .ZN(n964) );
  AND2_X1 U146bar ( .A1(n816bar), .A2(n815bar), .ZN(n964bar) );
  OR2_X1 U147 ( .A1(n814), .A2(n813), .ZN(n815) );
  AND2_X1 U147bar ( .A1(n814bar), .A2(n813bar), .ZN(n815bar) );
  OR2_X1 U148 ( .A1(n812), .A2(n811), .ZN(n813) );
  AND2_X1 U148bar ( .A1(n812bar), .A2(n811bar), .ZN(n813bar) );
  OR2_X1 U149 ( .A1(in[122]), .A2(in[111]), .ZN(n811) );
  AND2_X1 U149bar ( .A1(inbar[122]), .A2(inbar[111]), .ZN(n811bar) );
  OR2_X1 U150 ( .A1(in[154]), .A2(in[151]), .ZN(n812) );
  AND2_X1 U150bar ( .A1(inbar[154]), .A2(inbar[151]), .ZN(n812bar) );
  OR2_X1 U151 ( .A1(n810), .A2(n809), .ZN(n814) );
  AND2_X1 U151bar ( .A1(n810bar), .A2(n809bar), .ZN(n814bar) );
  OR2_X1 U152 ( .A1(in[187]), .A2(in[177]), .ZN(n809) );
  AND2_X1 U152bar ( .A1(inbar[187]), .A2(inbar[177]), .ZN(n809bar) );
  OR2_X1 U153 ( .A1(in[200]), .A2(in[192]), .ZN(n810) );
  AND2_X1 U153bar ( .A1(inbar[200]), .A2(inbar[192]), .ZN(n810bar) );
  OR2_X1 U154 ( .A1(n808), .A2(n807), .ZN(n816) );
  AND2_X1 U154bar ( .A1(n808bar), .A2(n807bar), .ZN(n816bar) );
  OR2_X1 U155 ( .A1(n806), .A2(n805), .ZN(n807) );
  AND2_X1 U155bar ( .A1(n806bar), .A2(n805bar), .ZN(n807bar) );
  OR2_X1 U156 ( .A1(in[225]), .A2(in[207]), .ZN(n805) );
  AND2_X1 U156bar ( .A1(inbar[225]), .A2(inbar[207]), .ZN(n805bar) );
  OR2_X1 U157 ( .A1(in[98]), .A2(in[226]), .ZN(n806) );
  AND2_X1 U157bar ( .A1(inbar[98]), .A2(inbar[226]), .ZN(n806bar) );
  OR2_X1 U158 ( .A1(n804), .A2(n803), .ZN(n808) );
  AND2_X1 U158bar ( .A1(n804bar), .A2(n803bar), .ZN(n808bar) );
  OR2_X1 U159 ( .A1(in_20), .A2(in_16), .ZN(n803) );
  AND2_X1 U159bar ( .A1(in_20bar), .A2(in_16bar), .ZN(n803bar) );
  OR2_X1 U160 ( .A1(in_55), .A2(in_45), .ZN(n804) );
  AND2_X1 U160bar ( .A1(in_55bar), .A2(in_45bar), .ZN(n804bar) );
  OR2_X1 U161 ( .A1(n802), .A2(n801), .ZN(n824) );
  AND2_X1 U161bar ( .A1(n802bar), .A2(n801bar), .ZN(n824bar) );
  OR2_X1 U162 ( .A1(in[162]), .A2(in[149]), .ZN(n801) );
  AND2_X1 U162bar ( .A1(inbar[162]), .A2(inbar[149]), .ZN(n801bar) );
  OR2_X1 U163 ( .A1(in[163]), .A2(n800), .ZN(n802) );
  AND2_X1 U163bar ( .A1(inbar[163]), .A2(n800bar), .ZN(n802bar) );
  OR2_X1 U164 ( .A1(in[191]), .A2(in[189]), .ZN(n800) );
  AND2_X1 U164bar ( .A1(inbar[191]), .A2(inbar[189]), .ZN(n800bar) );
  OR2_X1 U165 ( .A1(n799), .A2(n798), .ZN(n826) );
  AND2_X1 U165bar ( .A1(n799bar), .A2(n798bar), .ZN(n826bar) );
  OR2_X1 U166 ( .A1(n797), .A2(n796), .ZN(n798) );
  AND2_X1 U166bar ( .A1(n797bar), .A2(n796bar), .ZN(n798bar) );
  OR2_X1 U167 ( .A1(in[212]), .A2(in[193]), .ZN(n796) );
  AND2_X1 U167bar ( .A1(inbar[212]), .A2(inbar[193]), .ZN(n796bar) );
  OR2_X1 U168 ( .A1(in[238]), .A2(n795), .ZN(n797) );
  AND2_X1 U168bar ( .A1(inbar[238]), .A2(n795bar), .ZN(n797bar) );
  OR2_X1 U169 ( .A1(in[88]), .A2(in[247]), .ZN(n795) );
  AND2_X1 U169bar ( .A1(inbar[88]), .A2(inbar[247]), .ZN(n795bar) );
  OR2_X1 U170 ( .A1(n794), .A2(n793), .ZN(n799) );
  AND2_X1 U170bar ( .A1(n794bar), .A2(n793bar), .ZN(n799bar) );
  OR2_X1 U171 ( .A1(in[94]), .A2(in[92]), .ZN(n793) );
  AND2_X1 U171bar ( .A1(inbar[94]), .A2(inbar[92]), .ZN(n793bar) );
  OR2_X1 U172 ( .A1(in_52), .A2(n792), .ZN(n794) );
  AND2_X1 U172bar ( .A1(in_52bar), .A2(n792bar), .ZN(n794bar) );
  OR2_X1 U173 ( .A1(in_70), .A2(in_67), .ZN(n792) );
  AND2_X1 U173bar ( .A1(in_70bar), .A2(in_67bar), .ZN(n792bar) );
  OR2_X1 U174 ( .A1(n791), .A2(n790), .ZN(out[2]) );
  AND2_X1 U174bar ( .A1(n791bar), .A2(n790bar), .ZN(outbar[2]) );
  OR2_X1 U175 ( .A1(n789), .A2(n788), .ZN(n790) );
  AND2_X1 U175bar ( .A1(n789bar), .A2(n788bar), .ZN(n790bar) );
  OR2_X1 U176 ( .A1(n787), .A2(n786), .ZN(n788) );
  AND2_X1 U176bar ( .A1(n787bar), .A2(n786bar), .ZN(n788bar) );
  OR2_X1 U177 ( .A1(n819), .A2(n785), .ZN(n786) );
  AND2_X1 U177bar ( .A1(n819bar), .A2(n785bar), .ZN(n786bar) );
  OR2_X1 U178 ( .A1(n784), .A2(n783), .ZN(n819) );
  AND2_X1 U178bar ( .A1(n784bar), .A2(n783bar), .ZN(n819bar) );
  OR2_X1 U179 ( .A1(n782), .A2(n781), .ZN(n783) );
  AND2_X1 U179bar ( .A1(n782bar), .A2(n781bar), .ZN(n783bar) );
  OR2_X1 U180 ( .A1(n780), .A2(n779), .ZN(n781) );
  AND2_X1 U180bar ( .A1(n780bar), .A2(n779bar), .ZN(n781bar) );
  OR2_X1 U181 ( .A1(n962), .A2(n778), .ZN(n779) );
  AND2_X1 U181bar ( .A1(n962bar), .A2(n778bar), .ZN(n779bar) );
  OR2_X1 U182 ( .A1(n777), .A2(n776), .ZN(n962) );
  AND2_X1 U182bar ( .A1(n777bar), .A2(n776bar), .ZN(n962bar) );
  OR2_X1 U183 ( .A1(n775), .A2(n774), .ZN(n776) );
  AND2_X1 U183bar ( .A1(n775bar), .A2(n774bar), .ZN(n776bar) );
  OR2_X1 U184 ( .A1(n773), .A2(n772), .ZN(n774) );
  AND2_X1 U184bar ( .A1(n773bar), .A2(n772bar), .ZN(n774bar) );
  OR2_X1 U185 ( .A1(in[131]), .A2(in[120]), .ZN(n772) );
  AND2_X1 U185bar ( .A1(inbar[131]), .A2(inbar[120]), .ZN(n772bar) );
  OR2_X1 U186 ( .A1(in[153]), .A2(in[147]), .ZN(n773) );
  AND2_X1 U186bar ( .A1(inbar[153]), .A2(inbar[147]), .ZN(n773bar) );
  OR2_X1 U187 ( .A1(n771), .A2(n770), .ZN(n775) );
  AND2_X1 U187bar ( .A1(n771bar), .A2(n770bar), .ZN(n775bar) );
  OR2_X1 U188 ( .A1(in[170]), .A2(in[156]), .ZN(n770) );
  AND2_X1 U188bar ( .A1(inbar[170]), .A2(inbar[156]), .ZN(n770bar) );
  OR2_X1 U189 ( .A1(in[223]), .A2(in[190]), .ZN(n771) );
  AND2_X1 U189bar ( .A1(inbar[223]), .A2(inbar[190]), .ZN(n771bar) );
  OR2_X1 U190 ( .A1(n769), .A2(n768), .ZN(n777) );
  AND2_X1 U190bar ( .A1(n769bar), .A2(n768bar), .ZN(n777bar) );
  OR2_X1 U191 ( .A1(n767), .A2(n766), .ZN(n768) );
  AND2_X1 U191bar ( .A1(n767bar), .A2(n766bar), .ZN(n768bar) );
  OR2_X1 U192 ( .A1(in[236]), .A2(in[230]), .ZN(n766) );
  AND2_X1 U192bar ( .A1(inbar[236]), .A2(inbar[230]), .ZN(n766bar) );
  OR2_X1 U193 ( .A1(in[85]), .A2(in[240]), .ZN(n767) );
  AND2_X1 U193bar ( .A1(inbar[85]), .A2(inbar[240]), .ZN(n767bar) );
  OR2_X1 U194 ( .A1(n765), .A2(n764), .ZN(n769) );
  AND2_X1 U194bar ( .A1(n765bar), .A2(n764bar), .ZN(n769bar) );
  OR2_X1 U195 ( .A1(in_12), .A2(in[90]), .ZN(n764) );
  AND2_X1 U195bar ( .A1(in_12bar), .A2(inbar[90]), .ZN(n764bar) );
  OR2_X1 U196 ( .A1(in_39), .A2(in_28), .ZN(n765) );
  AND2_X1 U196bar ( .A1(in_39bar), .A2(in_28bar), .ZN(n765bar) );
  OR2_X1 U197 ( .A1(in[109]), .A2(n763), .ZN(n780) );
  AND2_X1 U197bar ( .A1(inbar[109]), .A2(n763bar), .ZN(n780bar) );
  OR2_X1 U198 ( .A1(n762), .A2(n761), .ZN(n782) );
  AND2_X1 U198bar ( .A1(n762bar), .A2(n761bar), .ZN(n782bar) );
  OR2_X1 U199 ( .A1(in[138]), .A2(in[129]), .ZN(n761) );
  AND2_X1 U199bar ( .A1(inbar[138]), .A2(inbar[129]), .ZN(n761bar) );
  OR2_X1 U200 ( .A1(in[157]), .A2(n760), .ZN(n762) );
  AND2_X1 U200bar ( .A1(inbar[157]), .A2(n760bar), .ZN(n762bar) );
  OR2_X1 U201 ( .A1(in[182]), .A2(in[167]), .ZN(n760) );
  AND2_X1 U201bar ( .A1(inbar[182]), .A2(inbar[167]), .ZN(n760bar) );
  OR2_X1 U202 ( .A1(n759), .A2(n758), .ZN(n784) );
  AND2_X1 U202bar ( .A1(n759bar), .A2(n758bar), .ZN(n784bar) );
  OR2_X1 U203 ( .A1(n757), .A2(n756), .ZN(n758) );
  AND2_X1 U203bar ( .A1(n757bar), .A2(n756bar), .ZN(n758bar) );
  OR2_X1 U204 ( .A1(in[195]), .A2(in[184]), .ZN(n756) );
  AND2_X1 U204bar ( .A1(inbar[195]), .A2(inbar[184]), .ZN(n756bar) );
  OR2_X1 U205 ( .A1(in[196]), .A2(n755), .ZN(n757) );
  AND2_X1 U205bar ( .A1(inbar[196]), .A2(n755bar), .ZN(n757bar) );
  OR2_X1 U206 ( .A1(in[215]), .A2(in[209]), .ZN(n755) );
  AND2_X1 U206bar ( .A1(inbar[215]), .A2(inbar[209]), .ZN(n755bar) );
  OR2_X1 U207 ( .A1(n754), .A2(n753), .ZN(n759) );
  AND2_X1 U207bar ( .A1(n754bar), .A2(n753bar), .ZN(n759bar) );
  OR2_X1 U208 ( .A1(in[93]), .A2(in[233]), .ZN(n753) );
  AND2_X1 U208bar ( .A1(inbar[93]), .A2(inbar[233]), .ZN(n753bar) );
  OR2_X1 U209 ( .A1(in_1), .A2(n752), .ZN(n754) );
  AND2_X1 U209bar ( .A1(in_1bar), .A2(n752bar), .ZN(n754bar) );
  OR2_X1 U210 ( .A1(in_69), .A2(in_66), .ZN(n752) );
  AND2_X1 U210bar ( .A1(in_69bar), .A2(in_66bar), .ZN(n752bar) );
  OR2_X1 U211 ( .A1(n966), .A2(n751), .ZN(n787) );
  AND2_X1 U211bar ( .A1(n966bar), .A2(n751bar), .ZN(n787bar) );
  OR2_X1 U212 ( .A1(in[134]), .A2(n750), .ZN(n751) );
  AND2_X1 U212bar ( .A1(inbar[134]), .A2(n750bar), .ZN(n751bar) );
  OR2_X1 U213 ( .A1(n749), .A2(n748), .ZN(n966) );
  AND2_X1 U213bar ( .A1(n749bar), .A2(n748bar), .ZN(n966bar) );
  OR2_X1 U214 ( .A1(n747), .A2(n746), .ZN(n748) );
  AND2_X1 U214bar ( .A1(n747bar), .A2(n746bar), .ZN(n748bar) );
  OR2_X1 U215 ( .A1(n745), .A2(n744), .ZN(n746) );
  AND2_X1 U215bar ( .A1(n745bar), .A2(n744bar), .ZN(n746bar) );
  OR2_X1 U216 ( .A1(in[136]), .A2(in[121]), .ZN(n744) );
  AND2_X1 U216bar ( .A1(inbar[136]), .A2(inbar[121]), .ZN(n744bar) );
  OR2_X1 U217 ( .A1(in[186]), .A2(in[174]), .ZN(n745) );
  AND2_X1 U217bar ( .A1(inbar[186]), .A2(inbar[174]), .ZN(n745bar) );
  OR2_X1 U218 ( .A1(n743), .A2(n742), .ZN(n747) );
  AND2_X1 U218bar ( .A1(n743bar), .A2(n742bar), .ZN(n747bar) );
  OR2_X1 U219 ( .A1(in[198]), .A2(in[197]), .ZN(n742) );
  AND2_X1 U219bar ( .A1(inbar[198]), .A2(inbar[197]), .ZN(n742bar) );
  OR2_X1 U220 ( .A1(in[214]), .A2(in[199]), .ZN(n743) );
  AND2_X1 U220bar ( .A1(inbar[214]), .A2(inbar[199]), .ZN(n743bar) );
  OR2_X1 U221 ( .A1(n741), .A2(n740), .ZN(n749) );
  AND2_X1 U221bar ( .A1(n741bar), .A2(n740bar), .ZN(n749bar) );
  OR2_X1 U222 ( .A1(n739), .A2(n738), .ZN(n740) );
  AND2_X1 U222bar ( .A1(n739bar), .A2(n738bar), .ZN(n740bar) );
  OR2_X1 U223 ( .A1(in[231]), .A2(in[220]), .ZN(n738) );
  AND2_X1 U223bar ( .A1(inbar[231]), .A2(inbar[220]), .ZN(n738bar) );
  OR2_X1 U224 ( .A1(in_25), .A2(in[245]), .ZN(n739) );
  AND2_X1 U224bar ( .A1(in_25bar), .A2(inbar[245]), .ZN(n739bar) );
  OR2_X1 U225 ( .A1(n737), .A2(n736), .ZN(n741) );
  AND2_X1 U225bar ( .A1(n737bar), .A2(n736bar), .ZN(n741bar) );
  OR2_X1 U226 ( .A1(in_53), .A2(in_29), .ZN(n736) );
  AND2_X1 U226bar ( .A1(in_53bar), .A2(in_29bar), .ZN(n736bar) );
  OR2_X1 U227 ( .A1(in_79), .A2(in_74), .ZN(n737) );
  AND2_X1 U227bar ( .A1(in_79bar), .A2(in_74bar), .ZN(n737bar) );
  OR2_X1 U228 ( .A1(n735), .A2(n734), .ZN(n789) );
  AND2_X1 U228bar ( .A1(n735bar), .A2(n734bar), .ZN(n789bar) );
  OR2_X1 U229 ( .A1(in[152]), .A2(in[140]), .ZN(n734) );
  AND2_X1 U229bar ( .A1(inbar[152]), .A2(inbar[140]), .ZN(n734bar) );
  OR2_X1 U230 ( .A1(in[155]), .A2(n733), .ZN(n735) );
  AND2_X1 U230bar ( .A1(inbar[155]), .A2(n733bar), .ZN(n735bar) );
  OR2_X1 U231 ( .A1(in[166]), .A2(in[165]), .ZN(n733) );
  AND2_X1 U231bar ( .A1(inbar[166]), .A2(inbar[165]), .ZN(n733bar) );
  OR2_X1 U232 ( .A1(n732), .A2(n731), .ZN(n791) );
  AND2_X1 U232bar ( .A1(n732bar), .A2(n731bar), .ZN(n791bar) );
  OR2_X1 U233 ( .A1(n730), .A2(n729), .ZN(n731) );
  AND2_X1 U233bar ( .A1(n730bar), .A2(n729bar), .ZN(n731bar) );
  OR2_X1 U234 ( .A1(in[202]), .A2(in[185]), .ZN(n729) );
  AND2_X1 U234bar ( .A1(inbar[202]), .A2(inbar[185]), .ZN(n729bar) );
  OR2_X1 U235 ( .A1(in[211]), .A2(n728), .ZN(n730) );
  AND2_X1 U235bar ( .A1(inbar[211]), .A2(n728bar), .ZN(n730bar) );
  OR2_X1 U236 ( .A1(in[255]), .A2(in[253]), .ZN(n728) );
  AND2_X1 U236bar ( .A1(inbar[255]), .A2(inbar[253]), .ZN(n728bar) );
  OR2_X1 U237 ( .A1(n727), .A2(n726), .ZN(n732) );
  AND2_X1 U237bar ( .A1(n727bar), .A2(n726bar), .ZN(n732bar) );
  OR2_X1 U238 ( .A1(in_35), .A2(in_15), .ZN(n726) );
  AND2_X1 U238bar ( .A1(in_35bar), .A2(in_15bar), .ZN(n726bar) );
  OR2_X1 U239 ( .A1(in_36), .A2(n725), .ZN(n727) );
  AND2_X1 U239bar ( .A1(in_36bar), .A2(n725bar), .ZN(n727bar) );
  OR2_X1 U240 ( .A1(in_48), .A2(in_40), .ZN(n725) );
  AND2_X1 U240bar ( .A1(in_48bar), .A2(in_40bar), .ZN(n725bar) );
  OR2_X1 U241 ( .A1(n724), .A2(n723), .ZN(out[1]) );
  AND2_X1 U241bar ( .A1(n724bar), .A2(n723bar), .ZN(outbar[1]) );
  OR2_X1 U242 ( .A1(n722), .A2(n721), .ZN(n723) );
  AND2_X1 U242bar ( .A1(n722bar), .A2(n721bar), .ZN(n723bar) );
  OR2_X1 U243 ( .A1(n720), .A2(n719), .ZN(n721) );
  AND2_X1 U243bar ( .A1(n720bar), .A2(n719bar), .ZN(n721bar) );
  OR2_X1 U244 ( .A1(n921), .A2(n887), .ZN(n719) );
  AND2_X1 U244bar ( .A1(n921bar), .A2(n887bar), .ZN(n719bar) );
  OR2_X1 U245 ( .A1(n718), .A2(n717), .ZN(n887) );
  AND2_X1 U245bar ( .A1(n718bar), .A2(n717bar), .ZN(n887bar) );
  OR2_X1 U246 ( .A1(n716), .A2(n715), .ZN(n717) );
  AND2_X1 U246bar ( .A1(n716bar), .A2(n715bar), .ZN(n717bar) );
  OR2_X1 U247 ( .A1(n714), .A2(n713), .ZN(n715) );
  AND2_X1 U247bar ( .A1(n714bar), .A2(n713bar), .ZN(n715bar) );
  OR2_X1 U248 ( .A1(in[116]), .A2(in[110]), .ZN(n713) );
  AND2_X1 U248bar ( .A1(inbar[116]), .A2(inbar[110]), .ZN(n713bar) );
  OR2_X1 U249 ( .A1(in[133]), .A2(in[130]), .ZN(n714) );
  AND2_X1 U249bar ( .A1(inbar[133]), .A2(inbar[130]), .ZN(n714bar) );
  OR2_X1 U250 ( .A1(n712), .A2(n711), .ZN(n716) );
  AND2_X1 U250bar ( .A1(n712bar), .A2(n711bar), .ZN(n716bar) );
  OR2_X1 U251 ( .A1(in[203]), .A2(in[135]), .ZN(n711) );
  AND2_X1 U251bar ( .A1(inbar[203]), .A2(inbar[135]), .ZN(n711bar) );
  OR2_X1 U252 ( .A1(in[232]), .A2(in[223]), .ZN(n712) );
  AND2_X1 U252bar ( .A1(inbar[232]), .A2(inbar[223]), .ZN(n712bar) );
  OR2_X1 U253 ( .A1(n710), .A2(n709), .ZN(n718) );
  AND2_X1 U253bar ( .A1(n710bar), .A2(n709bar), .ZN(n718bar) );
  OR2_X1 U254 ( .A1(n708), .A2(n707), .ZN(n709) );
  AND2_X1 U254bar ( .A1(n708bar), .A2(n707bar), .ZN(n709bar) );
  OR2_X1 U255 ( .A1(in[255]), .A2(in[233]), .ZN(n707) );
  AND2_X1 U255bar ( .A1(inbar[255]), .A2(inbar[233]), .ZN(n707bar) );
  OR2_X1 U256 ( .A1(in_53), .A2(in_34), .ZN(n708) );
  AND2_X1 U256bar ( .A1(in_53bar), .A2(in_34bar), .ZN(n708bar) );
  OR2_X1 U257 ( .A1(n706), .A2(n705), .ZN(n710) );
  AND2_X1 U257bar ( .A1(n706bar), .A2(n705bar), .ZN(n710bar) );
  OR2_X1 U258 ( .A1(in_57), .A2(in_55), .ZN(n705) );
  AND2_X1 U258bar ( .A1(in_57bar), .A2(in_55bar), .ZN(n705bar) );
  OR2_X1 U259 ( .A1(in_68), .A2(in_67), .ZN(n706) );
  AND2_X1 U259bar ( .A1(in_68bar), .A2(in_67bar), .ZN(n706bar) );
  OR2_X1 U260 ( .A1(n704), .A2(n703), .ZN(n921) );
  AND2_X1 U260bar ( .A1(n704bar), .A2(n703bar), .ZN(n921bar) );
  OR2_X1 U261 ( .A1(n702), .A2(n701), .ZN(n703) );
  AND2_X1 U261bar ( .A1(n702bar), .A2(n701bar), .ZN(n703bar) );
  OR2_X1 U262 ( .A1(n700), .A2(n699), .ZN(n701) );
  AND2_X1 U262bar ( .A1(n700bar), .A2(n699bar), .ZN(n701bar) );
  OR2_X1 U263 ( .A1(n944), .A2(n872), .ZN(n699) );
  AND2_X1 U263bar ( .A1(n944bar), .A2(n872bar), .ZN(n699bar) );
  OR2_X1 U264 ( .A1(n698), .A2(n697), .ZN(n872) );
  AND2_X1 U264bar ( .A1(n698bar), .A2(n697bar), .ZN(n872bar) );
  OR2_X1 U265 ( .A1(n696), .A2(n695), .ZN(n697) );
  AND2_X1 U265bar ( .A1(n696bar), .A2(n695bar), .ZN(n697bar) );
  OR2_X1 U266 ( .A1(n694), .A2(n693), .ZN(n695) );
  AND2_X1 U266bar ( .A1(n694bar), .A2(n693bar), .ZN(n695bar) );
  OR2_X1 U267 ( .A1(in[121]), .A2(in[102]), .ZN(n693) );
  AND2_X1 U267bar ( .A1(inbar[121]), .A2(inbar[102]), .ZN(n693bar) );
  OR2_X1 U268 ( .A1(in[162]), .A2(in[161]), .ZN(n694) );
  AND2_X1 U268bar ( .A1(inbar[162]), .A2(inbar[161]), .ZN(n694bar) );
  OR2_X1 U269 ( .A1(n692), .A2(n691), .ZN(n696) );
  AND2_X1 U269bar ( .A1(n692bar), .A2(n691bar), .ZN(n696bar) );
  OR2_X1 U270 ( .A1(in[192]), .A2(in[178]), .ZN(n691) );
  AND2_X1 U270bar ( .A1(inbar[192]), .A2(inbar[178]), .ZN(n691bar) );
  OR2_X1 U271 ( .A1(in[244]), .A2(in[209]), .ZN(n692) );
  AND2_X1 U271bar ( .A1(inbar[244]), .A2(inbar[209]), .ZN(n692bar) );
  OR2_X1 U272 ( .A1(n690), .A2(n689), .ZN(n698) );
  AND2_X1 U272bar ( .A1(n690bar), .A2(n689bar), .ZN(n698bar) );
  OR2_X1 U273 ( .A1(n688), .A2(n687), .ZN(n689) );
  AND2_X1 U273bar ( .A1(n688bar), .A2(n687bar), .ZN(n689bar) );
  OR2_X1 U274 ( .A1(in[90]), .A2(in[254]), .ZN(n687) );
  AND2_X1 U274bar ( .A1(inbar[90]), .A2(inbar[254]), .ZN(n687bar) );
  OR2_X1 U275 ( .A1(in_36), .A2(in_32), .ZN(n688) );
  AND2_X1 U275bar ( .A1(in_36bar), .A2(in_32bar), .ZN(n688bar) );
  OR2_X1 U276 ( .A1(n686), .A2(n685), .ZN(n690) );
  AND2_X1 U276bar ( .A1(n686bar), .A2(n685bar), .ZN(n690bar) );
  OR2_X1 U277 ( .A1(in_62), .A2(in_37), .ZN(n685) );
  AND2_X1 U277bar ( .A1(in_62bar), .A2(in_37bar), .ZN(n685bar) );
  OR2_X1 U278 ( .A1(in_75), .A2(in_73), .ZN(n686) );
  AND2_X1 U278bar ( .A1(in_75bar), .A2(in_73bar), .ZN(n686bar) );
  OR2_X1 U279 ( .A1(n684), .A2(n683), .ZN(n944) );
  AND2_X1 U279bar ( .A1(n684bar), .A2(n683bar), .ZN(n944bar) );
  OR2_X1 U280 ( .A1(n682), .A2(n681), .ZN(n683) );
  AND2_X1 U280bar ( .A1(n682bar), .A2(n681bar), .ZN(n683bar) );
  OR2_X1 U281 ( .A1(n680), .A2(n679), .ZN(n681) );
  AND2_X1 U281bar ( .A1(n680bar), .A2(n679bar), .ZN(n681bar) );
  OR2_X1 U282 ( .A1(in[171]), .A2(in[153]), .ZN(n679) );
  AND2_X1 U282bar ( .A1(inbar[171]), .A2(inbar[153]), .ZN(n679bar) );
  OR2_X1 U283 ( .A1(in[187]), .A2(in[176]), .ZN(n680) );
  AND2_X1 U283bar ( .A1(inbar[187]), .A2(inbar[176]), .ZN(n680bar) );
  OR2_X1 U284 ( .A1(n678), .A2(n677), .ZN(n682) );
  AND2_X1 U284bar ( .A1(n678bar), .A2(n677bar), .ZN(n682bar) );
  OR2_X1 U285 ( .A1(in[245]), .A2(in[211]), .ZN(n677) );
  AND2_X1 U285bar ( .A1(inbar[245]), .A2(inbar[211]), .ZN(n677bar) );
  OR2_X1 U286 ( .A1(in[97]), .A2(in[88]), .ZN(n678) );
  AND2_X1 U286bar ( .A1(inbar[97]), .A2(inbar[88]), .ZN(n678bar) );
  OR2_X1 U287 ( .A1(n676), .A2(n675), .ZN(n684) );
  AND2_X1 U287bar ( .A1(n676bar), .A2(n675bar), .ZN(n684bar) );
  OR2_X1 U288 ( .A1(n674), .A2(n673), .ZN(n675) );
  AND2_X1 U288bar ( .A1(n674bar), .A2(n673bar), .ZN(n675bar) );
  OR2_X1 U289 ( .A1(in_10), .A2(in_0), .ZN(n673) );
  AND2_X1 U289bar ( .A1(in_10bar), .A2(in_0bar), .ZN(n673bar) );
  OR2_X1 U290 ( .A1(in_59), .A2(in_5), .ZN(n674) );
  AND2_X1 U290bar ( .A1(in_59bar), .A2(in_5bar), .ZN(n674bar) );
  OR2_X1 U291 ( .A1(n672), .A2(n671), .ZN(n676) );
  AND2_X1 U291bar ( .A1(n672bar), .A2(n671bar), .ZN(n676bar) );
  OR2_X1 U292 ( .A1(in_60), .A2(in_6), .ZN(n671) );
  AND2_X1 U292bar ( .A1(in_60bar), .A2(in_6bar), .ZN(n671bar) );
  OR2_X1 U293 ( .A1(in_77), .A2(in_69), .ZN(n672) );
  AND2_X1 U293bar ( .A1(in_77bar), .A2(in_69bar), .ZN(n672bar) );
  OR2_X1 U294 ( .A1(in[113]), .A2(n864), .ZN(n700) );
  AND2_X1 U294bar ( .A1(inbar[113]), .A2(n864bar), .ZN(n700bar) );
  OR2_X1 U295 ( .A1(n670), .A2(n669), .ZN(n864) );
  AND2_X1 U295bar ( .A1(n670bar), .A2(n669bar), .ZN(n864bar) );
  OR2_X1 U296 ( .A1(n668), .A2(n667), .ZN(n669) );
  AND2_X1 U296bar ( .A1(n668bar), .A2(n667bar), .ZN(n669bar) );
  OR2_X1 U297 ( .A1(n666), .A2(n665), .ZN(n667) );
  AND2_X1 U297bar ( .A1(n666bar), .A2(n665bar), .ZN(n667bar) );
  OR2_X1 U298 ( .A1(in[125]), .A2(in[107]), .ZN(n665) );
  AND2_X1 U298bar ( .A1(inbar[125]), .A2(inbar[107]), .ZN(n665bar) );
  OR2_X1 U299 ( .A1(in[138]), .A2(in[126]), .ZN(n666) );
  AND2_X1 U299bar ( .A1(inbar[138]), .A2(inbar[126]), .ZN(n666bar) );
  OR2_X1 U300 ( .A1(n664), .A2(n663), .ZN(n668) );
  AND2_X1 U300bar ( .A1(n664bar), .A2(n663bar), .ZN(n668bar) );
  OR2_X1 U301 ( .A1(in[189]), .A2(in[143]), .ZN(n663) );
  AND2_X1 U301bar ( .A1(inbar[189]), .A2(inbar[143]), .ZN(n663bar) );
  OR2_X1 U302 ( .A1(in[99]), .A2(in[214]), .ZN(n664) );
  AND2_X1 U302bar ( .A1(inbar[99]), .A2(inbar[214]), .ZN(n664bar) );
  OR2_X1 U303 ( .A1(n662), .A2(n661), .ZN(n670) );
  AND2_X1 U303bar ( .A1(n662bar), .A2(n661bar), .ZN(n670bar) );
  OR2_X1 U304 ( .A1(n660), .A2(n659), .ZN(n661) );
  AND2_X1 U304bar ( .A1(n660bar), .A2(n659bar), .ZN(n661bar) );
  OR2_X1 U305 ( .A1(in_15), .A2(in_12), .ZN(n659) );
  AND2_X1 U305bar ( .A1(in_15bar), .A2(in_12bar), .ZN(n659bar) );
  OR2_X1 U306 ( .A1(in_20), .A2(in_2), .ZN(n660) );
  AND2_X1 U306bar ( .A1(in_20bar), .A2(in_2bar), .ZN(n660bar) );
  OR2_X1 U307 ( .A1(n658), .A2(n657), .ZN(n662) );
  AND2_X1 U307bar ( .A1(n658bar), .A2(n657bar), .ZN(n662bar) );
  OR2_X1 U308 ( .A1(in_30), .A2(in_3), .ZN(n657) );
  AND2_X1 U308bar ( .A1(in_30bar), .A2(in_3bar), .ZN(n657bar) );
  OR2_X1 U309 ( .A1(in_4), .A2(in_38), .ZN(n658) );
  AND2_X1 U309bar ( .A1(in_4bar), .A2(in_38bar), .ZN(n658bar) );
  OR2_X1 U310 ( .A1(n656), .A2(n655), .ZN(n702) );
  AND2_X1 U310bar ( .A1(n656bar), .A2(n655bar), .ZN(n702bar) );
  OR2_X1 U311 ( .A1(in[148]), .A2(in[137]), .ZN(n655) );
  AND2_X1 U311bar ( .A1(inbar[148]), .A2(inbar[137]), .ZN(n655bar) );
  OR2_X1 U312 ( .A1(in[149]), .A2(n654), .ZN(n656) );
  AND2_X1 U312bar ( .A1(inbar[149]), .A2(n654bar), .ZN(n656bar) );
  OR2_X1 U313 ( .A1(in[195]), .A2(in[190]), .ZN(n654) );
  AND2_X1 U313bar ( .A1(inbar[195]), .A2(inbar[190]), .ZN(n654bar) );
  OR2_X1 U314 ( .A1(n653), .A2(n652), .ZN(n704) );
  AND2_X1 U314bar ( .A1(n653bar), .A2(n652bar), .ZN(n704bar) );
  OR2_X1 U315 ( .A1(n651), .A2(n650), .ZN(n652) );
  AND2_X1 U315bar ( .A1(n651bar), .A2(n650bar), .ZN(n652bar) );
  OR2_X1 U316 ( .A1(in[98]), .A2(in[197]), .ZN(n650) );
  AND2_X1 U316bar ( .A1(inbar[98]), .A2(inbar[197]), .ZN(n650bar) );
  OR2_X1 U317 ( .A1(in_11), .A2(n649), .ZN(n651) );
  AND2_X1 U317bar ( .A1(in_11bar), .A2(n649bar), .ZN(n651bar) );
  OR2_X1 U318 ( .A1(in_26), .A2(in_14), .ZN(n649) );
  AND2_X1 U318bar ( .A1(in_26bar), .A2(in_14bar), .ZN(n649bar) );
  OR2_X1 U319 ( .A1(n648), .A2(n647), .ZN(n653) );
  AND2_X1 U319bar ( .A1(n648bar), .A2(n647bar), .ZN(n653bar) );
  OR2_X1 U320 ( .A1(in_35), .A2(in_27), .ZN(n647) );
  AND2_X1 U320bar ( .A1(in_35bar), .A2(in_27bar), .ZN(n647bar) );
  OR2_X1 U321 ( .A1(in_50), .A2(n646), .ZN(n648) );
  AND2_X1 U321bar ( .A1(in_50bar), .A2(n646bar), .ZN(n648bar) );
  OR2_X1 U322 ( .A1(in_78), .A2(in_61), .ZN(n646) );
  AND2_X1 U322bar ( .A1(in_78bar), .A2(in_61bar), .ZN(n646bar) );
  OR2_X1 U323 ( .A1(n942), .A2(n645), .ZN(n720) );
  AND2_X1 U323bar ( .A1(n942bar), .A2(n645bar), .ZN(n720bar) );
  OR2_X1 U324 ( .A1(in[106]), .A2(n863), .ZN(n645) );
  AND2_X1 U324bar ( .A1(inbar[106]), .A2(n863bar), .ZN(n645bar) );
  OR2_X1 U325 ( .A1(n644), .A2(n643), .ZN(n863) );
  AND2_X1 U325bar ( .A1(n644bar), .A2(n643bar), .ZN(n863bar) );
  OR2_X1 U326 ( .A1(n642), .A2(n641), .ZN(n643) );
  AND2_X1 U326bar ( .A1(n642bar), .A2(n641bar), .ZN(n643bar) );
  OR2_X1 U327 ( .A1(n640), .A2(n639), .ZN(n641) );
  AND2_X1 U327bar ( .A1(n640bar), .A2(n639bar), .ZN(n641bar) );
  OR2_X1 U328 ( .A1(in[127]), .A2(in[122]), .ZN(n639) );
  AND2_X1 U328bar ( .A1(inbar[127]), .A2(inbar[122]), .ZN(n639bar) );
  OR2_X1 U329 ( .A1(in[156]), .A2(in[132]), .ZN(n640) );
  AND2_X1 U329bar ( .A1(inbar[156]), .A2(inbar[132]), .ZN(n640bar) );
  OR2_X1 U330 ( .A1(n638), .A2(n637), .ZN(n642) );
  AND2_X1 U330bar ( .A1(n638bar), .A2(n637bar), .ZN(n642bar) );
  OR2_X1 U331 ( .A1(in[159]), .A2(in[157]), .ZN(n637) );
  AND2_X1 U331bar ( .A1(inbar[159]), .A2(inbar[157]), .ZN(n637bar) );
  OR2_X1 U332 ( .A1(in[185]), .A2(in[169]), .ZN(n638) );
  AND2_X1 U332bar ( .A1(inbar[185]), .A2(inbar[169]), .ZN(n638bar) );
  OR2_X1 U333 ( .A1(n636), .A2(n635), .ZN(n644) );
  AND2_X1 U333bar ( .A1(n636bar), .A2(n635bar), .ZN(n644bar) );
  OR2_X1 U334 ( .A1(n634), .A2(n633), .ZN(n635) );
  AND2_X1 U334bar ( .A1(n634bar), .A2(n633bar), .ZN(n635bar) );
  OR2_X1 U335 ( .A1(in[239]), .A2(in[218]), .ZN(n633) );
  AND2_X1 U335bar ( .A1(inbar[239]), .A2(inbar[218]), .ZN(n633bar) );
  OR2_X1 U336 ( .A1(in_13), .A2(in[87]), .ZN(n634) );
  AND2_X1 U336bar ( .A1(in_13bar), .A2(inbar[87]), .ZN(n634bar) );
  OR2_X1 U337 ( .A1(n632), .A2(n631), .ZN(n636) );
  AND2_X1 U337bar ( .A1(n632bar), .A2(n631bar), .ZN(n636bar) );
  OR2_X1 U338 ( .A1(in_72), .A2(in_70), .ZN(n631) );
  AND2_X1 U338bar ( .A1(in_72bar), .A2(in_70bar), .ZN(n631bar) );
  OR2_X1 U339 ( .A1(in_80), .A2(in_74), .ZN(n632) );
  AND2_X1 U339bar ( .A1(in_80bar), .A2(in_74bar), .ZN(n632bar) );
  OR2_X1 U340 ( .A1(n630), .A2(n629), .ZN(n942) );
  AND2_X1 U340bar ( .A1(n630bar), .A2(n629bar), .ZN(n942bar) );
  OR2_X1 U341 ( .A1(n628), .A2(n627), .ZN(n629) );
  AND2_X1 U341bar ( .A1(n628bar), .A2(n627bar), .ZN(n629bar) );
  OR2_X1 U342 ( .A1(n626), .A2(n625), .ZN(n627) );
  AND2_X1 U342bar ( .A1(n626bar), .A2(n625bar), .ZN(n627bar) );
  OR2_X1 U343 ( .A1(in[146]), .A2(in[100]), .ZN(n625) );
  AND2_X1 U343bar ( .A1(inbar[146]), .A2(inbar[100]), .ZN(n625bar) );
  OR2_X1 U344 ( .A1(in[168]), .A2(in[152]), .ZN(n626) );
  AND2_X1 U344bar ( .A1(inbar[168]), .A2(inbar[152]), .ZN(n626bar) );
  OR2_X1 U345 ( .A1(n624), .A2(n623), .ZN(n628) );
  AND2_X1 U345bar ( .A1(n624bar), .A2(n623bar), .ZN(n628bar) );
  OR2_X1 U346 ( .A1(in[199]), .A2(in[182]), .ZN(n623) );
  AND2_X1 U346bar ( .A1(inbar[199]), .A2(inbar[182]), .ZN(n623bar) );
  OR2_X1 U347 ( .A1(in[236]), .A2(in[204]), .ZN(n624) );
  AND2_X1 U347bar ( .A1(inbar[236]), .A2(inbar[204]), .ZN(n624bar) );
  OR2_X1 U348 ( .A1(n622), .A2(n621), .ZN(n630) );
  AND2_X1 U348bar ( .A1(n622bar), .A2(n621bar), .ZN(n630bar) );
  OR2_X1 U349 ( .A1(n620), .A2(n619), .ZN(n621) );
  AND2_X1 U349bar ( .A1(n620bar), .A2(n619bar), .ZN(n621bar) );
  OR2_X1 U350 ( .A1(in[89]), .A2(in[246]), .ZN(n619) );
  AND2_X1 U350bar ( .A1(inbar[89]), .A2(inbar[246]), .ZN(n619bar) );
  OR2_X1 U351 ( .A1(in[95]), .A2(in[92]), .ZN(n620) );
  AND2_X1 U351bar ( .A1(inbar[95]), .A2(inbar[92]), .ZN(n620bar) );
  OR2_X1 U352 ( .A1(n618), .A2(n617), .ZN(n622) );
  AND2_X1 U352bar ( .A1(n618bar), .A2(n617bar), .ZN(n622bar) );
  OR2_X1 U353 ( .A1(in_22), .A2(in_16), .ZN(n617) );
  AND2_X1 U353bar ( .A1(in_22bar), .A2(in_16bar), .ZN(n617bar) );
  OR2_X1 U354 ( .A1(in_51), .A2(in_49), .ZN(n618) );
  AND2_X1 U354bar ( .A1(in_51bar), .A2(in_49bar), .ZN(n618bar) );
  OR2_X1 U355 ( .A1(n616), .A2(n615), .ZN(n722) );
  AND2_X1 U355bar ( .A1(n616bar), .A2(n615bar), .ZN(n722bar) );
  OR2_X1 U356 ( .A1(in[158]), .A2(in[115]), .ZN(n615) );
  AND2_X1 U356bar ( .A1(inbar[158]), .A2(inbar[115]), .ZN(n615bar) );
  OR2_X1 U357 ( .A1(in[163]), .A2(n614), .ZN(n616) );
  AND2_X1 U357bar ( .A1(inbar[163]), .A2(n614bar), .ZN(n616bar) );
  OR2_X1 U358 ( .A1(in[206]), .A2(in[165]), .ZN(n614) );
  AND2_X1 U358bar ( .A1(inbar[206]), .A2(inbar[165]), .ZN(n614bar) );
  OR2_X1 U359 ( .A1(n613), .A2(n612), .ZN(n724) );
  AND2_X1 U359bar ( .A1(n613bar), .A2(n612bar), .ZN(n724bar) );
  OR2_X1 U360 ( .A1(n611), .A2(n610), .ZN(n612) );
  AND2_X1 U360bar ( .A1(n611bar), .A2(n610bar), .ZN(n612bar) );
  OR2_X1 U361 ( .A1(in[213]), .A2(in[207]), .ZN(n610) );
  AND2_X1 U361bar ( .A1(inbar[213]), .A2(inbar[207]), .ZN(n610bar) );
  OR2_X1 U362 ( .A1(in[215]), .A2(n609), .ZN(n611) );
  AND2_X1 U362bar ( .A1(inbar[215]), .A2(n609bar), .ZN(n611bar) );
  OR2_X1 U363 ( .A1(in[230]), .A2(in[220]), .ZN(n609) );
  AND2_X1 U363bar ( .A1(inbar[230]), .A2(inbar[220]), .ZN(n609bar) );
  OR2_X1 U364 ( .A1(n608), .A2(n607), .ZN(n613) );
  AND2_X1 U364bar ( .A1(n608bar), .A2(n607bar), .ZN(n613bar) );
  OR2_X1 U365 ( .A1(in[251]), .A2(in[234]), .ZN(n607) );
  AND2_X1 U365bar ( .A1(inbar[251]), .A2(inbar[234]), .ZN(n607bar) );
  OR2_X1 U366 ( .A1(in_17), .A2(n606), .ZN(n608) );
  AND2_X1 U366bar ( .A1(in_17bar), .A2(n606bar), .ZN(n608bar) );
  OR2_X1 U367 ( .A1(in_65), .A2(in_56), .ZN(n606) );
  AND2_X1 U367bar ( .A1(in_65bar), .A2(in_56bar), .ZN(n606bar) );
  OR2_X1 U368 ( .A1(n605), .A2(n604), .ZN(out[0]) );
  AND2_X1 U368bar ( .A1(n605bar), .A2(n604bar), .ZN(outbar[0]) );
  OR2_X1 U369 ( .A1(n603), .A2(n602), .ZN(n604) );
  AND2_X1 U369bar ( .A1(n603bar), .A2(n602bar), .ZN(n604bar) );
  OR2_X1 U370 ( .A1(n601), .A2(n600), .ZN(n602) );
  AND2_X1 U370bar ( .A1(n601bar), .A2(n600bar), .ZN(n602bar) );
  OR2_X1 U371 ( .A1(n820), .A2(n785), .ZN(n600) );
  AND2_X1 U371bar ( .A1(n820bar), .A2(n785bar), .ZN(n600bar) );
  OR2_X1 U372 ( .A1(n599), .A2(n598), .ZN(n785) );
  AND2_X1 U372bar ( .A1(n599bar), .A2(n598bar), .ZN(n785bar) );
  OR2_X1 U373 ( .A1(n597), .A2(n596), .ZN(n598) );
  AND2_X1 U373bar ( .A1(n597bar), .A2(n596bar), .ZN(n598bar) );
  OR2_X1 U374 ( .A1(n595), .A2(n594), .ZN(n596) );
  AND2_X1 U374bar ( .A1(n595bar), .A2(n594bar), .ZN(n596bar) );
  OR2_X1 U375 ( .A1(in[135]), .A2(in[104]), .ZN(n594) );
  AND2_X1 U375bar ( .A1(inbar[135]), .A2(inbar[104]), .ZN(n594bar) );
  OR2_X1 U376 ( .A1(in[188]), .A2(in[178]), .ZN(n595) );
  AND2_X1 U376bar ( .A1(inbar[188]), .A2(inbar[178]), .ZN(n595bar) );
  OR2_X1 U377 ( .A1(n593), .A2(n592), .ZN(n597) );
  AND2_X1 U377bar ( .A1(n593bar), .A2(n592bar), .ZN(n597bar) );
  OR2_X1 U378 ( .A1(in[217]), .A2(in[194]), .ZN(n592) );
  AND2_X1 U378bar ( .A1(inbar[217]), .A2(inbar[194]), .ZN(n592bar) );
  OR2_X1 U379 ( .A1(in[237]), .A2(in[218]), .ZN(n593) );
  AND2_X1 U379bar ( .A1(inbar[237]), .A2(inbar[218]), .ZN(n593bar) );
  OR2_X1 U380 ( .A1(n591), .A2(n590), .ZN(n599) );
  AND2_X1 U380bar ( .A1(n591bar), .A2(n590bar), .ZN(n599bar) );
  OR2_X1 U381 ( .A1(n589), .A2(n588), .ZN(n590) );
  AND2_X1 U381bar ( .A1(n589bar), .A2(n588bar), .ZN(n590bar) );
  OR2_X1 U382 ( .A1(in_2), .A2(in_10), .ZN(n588) );
  AND2_X1 U382bar ( .A1(in_2bar), .A2(in_10bar), .ZN(n588bar) );
  OR2_X1 U383 ( .A1(in_47), .A2(in_22), .ZN(n589) );
  AND2_X1 U383bar ( .A1(in_47bar), .A2(in_22bar), .ZN(n589bar) );
  OR2_X1 U384 ( .A1(n587), .A2(n586), .ZN(n591) );
  AND2_X1 U384bar ( .A1(n587bar), .A2(n586bar), .ZN(n591bar) );
  OR2_X1 U385 ( .A1(in_56), .A2(in_54), .ZN(n586) );
  AND2_X1 U385bar ( .A1(in_56bar), .A2(in_54bar), .ZN(n586bar) );
  OR2_X1 U386 ( .A1(in_63), .A2(in_61), .ZN(n587) );
  AND2_X1 U386bar ( .A1(in_63bar), .A2(in_61bar), .ZN(n587bar) );
  OR2_X1 U387 ( .A1(n585), .A2(n584), .ZN(n820) );
  AND2_X1 U387bar ( .A1(n585bar), .A2(n584bar), .ZN(n820bar) );
  OR2_X1 U388 ( .A1(n583), .A2(n582), .ZN(n584) );
  AND2_X1 U388bar ( .A1(n583bar), .A2(n582bar), .ZN(n584bar) );
  OR2_X1 U389 ( .A1(n581), .A2(n580), .ZN(n582) );
  AND2_X1 U389bar ( .A1(n581bar), .A2(n580bar), .ZN(n582bar) );
  OR2_X1 U390 ( .A1(in[158]), .A2(in[142]), .ZN(n580) );
  AND2_X1 U390bar ( .A1(inbar[158]), .A2(inbar[142]), .ZN(n580bar) );
  OR2_X1 U391 ( .A1(in[175]), .A2(in[164]), .ZN(n581) );
  AND2_X1 U391bar ( .A1(inbar[175]), .A2(inbar[164]), .ZN(n581bar) );
  OR2_X1 U392 ( .A1(n579), .A2(n578), .ZN(n583) );
  AND2_X1 U392bar ( .A1(n579bar), .A2(n578bar), .ZN(n583bar) );
  OR2_X1 U393 ( .A1(in[228]), .A2(in[204]), .ZN(n578) );
  AND2_X1 U393bar ( .A1(inbar[228]), .A2(inbar[204]), .ZN(n578bar) );
  OR2_X1 U394 ( .A1(in[91]), .A2(in[87]), .ZN(n579) );
  AND2_X1 U394bar ( .A1(inbar[91]), .A2(inbar[87]), .ZN(n579bar) );
  OR2_X1 U395 ( .A1(n577), .A2(n576), .ZN(n585) );
  AND2_X1 U395bar ( .A1(n577bar), .A2(n576bar), .ZN(n585bar) );
  OR2_X1 U396 ( .A1(n575), .A2(n574), .ZN(n576) );
  AND2_X1 U396bar ( .A1(n575bar), .A2(n574bar), .ZN(n576bar) );
  OR2_X1 U397 ( .A1(in_21), .A2(in_11), .ZN(n574) );
  AND2_X1 U397bar ( .A1(in_21bar), .A2(in_11bar), .ZN(n574bar) );
  OR2_X1 U398 ( .A1(in_5), .A2(in_3), .ZN(n575) );
  AND2_X1 U398bar ( .A1(in_5bar), .A2(in_3bar), .ZN(n575bar) );
  OR2_X1 U399 ( .A1(n573), .A2(n572), .ZN(n577) );
  AND2_X1 U399bar ( .A1(n573bar), .A2(n572bar), .ZN(n577bar) );
  OR2_X1 U400 ( .A1(in_68), .A2(in_64), .ZN(n572) );
  AND2_X1 U400bar ( .A1(in_68bar), .A2(in_64bar), .ZN(n572bar) );
  OR2_X1 U401 ( .A1(in_76), .A2(in_73), .ZN(n573) );
  AND2_X1 U401bar ( .A1(in_76bar), .A2(in_73bar), .ZN(n573bar) );
  OR2_X1 U402 ( .A1(n778), .A2(n571), .ZN(n601) );
  AND2_X1 U402bar ( .A1(n778bar), .A2(n571bar), .ZN(n601bar) );
  OR2_X1 U403 ( .A1(in[100]), .A2(n965), .ZN(n571) );
  AND2_X1 U403bar ( .A1(inbar[100]), .A2(n965bar), .ZN(n571bar) );
  OR2_X1 U404 ( .A1(n570), .A2(n569), .ZN(n965) );
  AND2_X1 U404bar ( .A1(n570bar), .A2(n569bar), .ZN(n965bar) );
  OR2_X1 U405 ( .A1(n568), .A2(n567), .ZN(n569) );
  AND2_X1 U405bar ( .A1(n568bar), .A2(n567bar), .ZN(n569bar) );
  OR2_X1 U406 ( .A1(n566), .A2(n565), .ZN(n567) );
  AND2_X1 U406bar ( .A1(n566bar), .A2(n565bar), .ZN(n567bar) );
  OR2_X1 U407 ( .A1(n817), .A2(n750), .ZN(n565) );
  AND2_X1 U407bar ( .A1(n817bar), .A2(n750bar), .ZN(n565bar) );
  OR2_X1 U408 ( .A1(n564), .A2(n563), .ZN(n750) );
  AND2_X1 U408bar ( .A1(n564bar), .A2(n563bar), .ZN(n750bar) );
  OR2_X1 U409 ( .A1(n562), .A2(n561), .ZN(n563) );
  AND2_X1 U409bar ( .A1(n562bar), .A2(n561bar), .ZN(n563bar) );
  OR2_X1 U410 ( .A1(n560), .A2(n559), .ZN(n561) );
  AND2_X1 U410bar ( .A1(n560bar), .A2(n559bar), .ZN(n561bar) );
  OR2_X1 U411 ( .A1(in[119]), .A2(in[103]), .ZN(n559) );
  AND2_X1 U411bar ( .A1(inbar[119]), .A2(inbar[103]), .ZN(n559bar) );
  OR2_X1 U412 ( .A1(in[137]), .A2(in[133]), .ZN(n560) );
  AND2_X1 U412bar ( .A1(inbar[137]), .A2(inbar[133]), .ZN(n560bar) );
  OR2_X1 U413 ( .A1(n558), .A2(n557), .ZN(n562) );
  AND2_X1 U413bar ( .A1(n558bar), .A2(n557bar), .ZN(n562bar) );
  OR2_X1 U414 ( .A1(in[176]), .A2(in[173]), .ZN(n557) );
  AND2_X1 U414bar ( .A1(inbar[176]), .A2(inbar[173]), .ZN(n557bar) );
  OR2_X1 U415 ( .A1(in[210]), .A2(in[181]), .ZN(n558) );
  AND2_X1 U415bar ( .A1(inbar[210]), .A2(inbar[181]), .ZN(n558bar) );
  OR2_X1 U416 ( .A1(n556), .A2(n555), .ZN(n564) );
  AND2_X1 U416bar ( .A1(n556bar), .A2(n555bar), .ZN(n564bar) );
  OR2_X1 U417 ( .A1(n554), .A2(n553), .ZN(n555) );
  AND2_X1 U417bar ( .A1(n554bar), .A2(n553bar), .ZN(n555bar) );
  OR2_X1 U418 ( .A1(in_13), .A2(in[234]), .ZN(n553) );
  AND2_X1 U418bar ( .A1(in_13bar), .A2(inbar[234]), .ZN(n553bar) );
  OR2_X1 U419 ( .A1(in_38), .A2(in_32), .ZN(n554) );
  AND2_X1 U419bar ( .A1(in_38bar), .A2(in_32bar), .ZN(n554bar) );
  OR2_X1 U420 ( .A1(n552), .A2(n551), .ZN(n556) );
  AND2_X1 U420bar ( .A1(n552bar), .A2(n551bar), .ZN(n556bar) );
  OR2_X1 U421 ( .A1(in_42), .A2(in_41), .ZN(n551) );
  AND2_X1 U421bar ( .A1(in_42bar), .A2(in_41bar), .ZN(n551bar) );
  OR2_X1 U422 ( .A1(in_7), .A2(in_49), .ZN(n552) );
  AND2_X1 U422bar ( .A1(in_7bar), .A2(in_49bar), .ZN(n552bar) );
  OR2_X1 U423 ( .A1(n550), .A2(n549), .ZN(n817) );
  AND2_X1 U423bar ( .A1(n550bar), .A2(n549bar), .ZN(n817bar) );
  OR2_X1 U424 ( .A1(n548), .A2(n547), .ZN(n549) );
  AND2_X1 U424bar ( .A1(n548bar), .A2(n547bar), .ZN(n549bar) );
  OR2_X1 U425 ( .A1(n546), .A2(n545), .ZN(n547) );
  AND2_X1 U425bar ( .A1(n546bar), .A2(n545bar), .ZN(n547bar) );
  OR2_X1 U426 ( .A1(in[159]), .A2(in[105]), .ZN(n545) );
  AND2_X1 U426bar ( .A1(inbar[159]), .A2(inbar[105]), .ZN(n545bar) );
  OR2_X1 U427 ( .A1(in[206]), .A2(in[183]), .ZN(n546) );
  AND2_X1 U427bar ( .A1(inbar[206]), .A2(inbar[183]), .ZN(n546bar) );
  OR2_X1 U428 ( .A1(n544), .A2(n543), .ZN(n548) );
  AND2_X1 U428bar ( .A1(n544bar), .A2(n543bar), .ZN(n548bar) );
  OR2_X1 U429 ( .A1(in[229]), .A2(in[219]), .ZN(n543) );
  AND2_X1 U429bar ( .A1(inbar[229]), .A2(inbar[219]), .ZN(n543bar) );
  OR2_X1 U430 ( .A1(in[235]), .A2(in[232]), .ZN(n544) );
  AND2_X1 U430bar ( .A1(inbar[235]), .A2(inbar[232]), .ZN(n544bar) );
  OR2_X1 U431 ( .A1(n542), .A2(n541), .ZN(n550) );
  AND2_X1 U431bar ( .A1(n542bar), .A2(n541bar), .ZN(n550bar) );
  OR2_X1 U432 ( .A1(n540), .A2(n539), .ZN(n541) );
  AND2_X1 U432bar ( .A1(n540bar), .A2(n539bar), .ZN(n541bar) );
  OR2_X1 U433 ( .A1(in[249]), .A2(in[242]), .ZN(n539) );
  AND2_X1 U433bar ( .A1(inbar[249]), .A2(inbar[242]), .ZN(n539bar) );
  OR2_X1 U434 ( .A1(in[89]), .A2(in[254]), .ZN(n540) );
  AND2_X1 U434bar ( .A1(inbar[89]), .A2(inbar[254]), .ZN(n540bar) );
  OR2_X1 U435 ( .A1(n538), .A2(n537), .ZN(n542) );
  AND2_X1 U435bar ( .A1(n538bar), .A2(n537bar), .ZN(n542bar) );
  OR2_X1 U436 ( .A1(in_14), .A2(in[99]), .ZN(n537) );
  AND2_X1 U436bar ( .A1(in_14bar), .A2(inbar[99]), .ZN(n537bar) );
  OR2_X1 U437 ( .A1(in_60), .A2(in_18), .ZN(n538) );
  AND2_X1 U437bar ( .A1(in_60bar), .A2(in_18bar), .ZN(n538bar) );
  OR2_X1 U438 ( .A1(in[113]), .A2(n763), .ZN(n566) );
  AND2_X1 U438bar ( .A1(inbar[113]), .A2(n763bar), .ZN(n566bar) );
  OR2_X1 U439 ( .A1(n536), .A2(n535), .ZN(n763) );
  AND2_X1 U439bar ( .A1(n536bar), .A2(n535bar), .ZN(n763bar) );
  OR2_X1 U440 ( .A1(n534), .A2(n533), .ZN(n535) );
  AND2_X1 U440bar ( .A1(n534bar), .A2(n533bar), .ZN(n535bar) );
  OR2_X1 U441 ( .A1(n532), .A2(n531), .ZN(n533) );
  AND2_X1 U441bar ( .A1(n532bar), .A2(n531bar), .ZN(n533bar) );
  OR2_X1 U442 ( .A1(in[115]), .A2(in[110]), .ZN(n531) );
  AND2_X1 U442bar ( .A1(inbar[115]), .A2(inbar[110]), .ZN(n531bar) );
  OR2_X1 U443 ( .A1(in[125]), .A2(in[117]), .ZN(n532) );
  AND2_X1 U443bar ( .A1(inbar[125]), .A2(inbar[117]), .ZN(n532bar) );
  OR2_X1 U444 ( .A1(n530), .A2(n529), .ZN(n534) );
  AND2_X1 U444bar ( .A1(n530bar), .A2(n529bar), .ZN(n534bar) );
  OR2_X1 U445 ( .A1(in[180]), .A2(in[128]), .ZN(n529) );
  AND2_X1 U445bar ( .A1(inbar[180]), .A2(inbar[128]), .ZN(n529bar) );
  OR2_X1 U446 ( .A1(in[205]), .A2(in[201]), .ZN(n530) );
  AND2_X1 U446bar ( .A1(inbar[205]), .A2(inbar[201]), .ZN(n530bar) );
  OR2_X1 U447 ( .A1(n528), .A2(n527), .ZN(n536) );
  AND2_X1 U447bar ( .A1(n528bar), .A2(n527bar), .ZN(n536bar) );
  OR2_X1 U448 ( .A1(n526), .A2(n525), .ZN(n527) );
  AND2_X1 U448bar ( .A1(n526bar), .A2(n525bar), .ZN(n527bar) );
  OR2_X1 U449 ( .A1(in[244]), .A2(in[239]), .ZN(n525) );
  AND2_X1 U449bar ( .A1(inbar[244]), .A2(inbar[239]), .ZN(n525bar) );
  OR2_X1 U450 ( .A1(in[95]), .A2(in[83]), .ZN(n526) );
  AND2_X1 U450bar ( .A1(inbar[95]), .A2(inbar[83]), .ZN(n526bar) );
  OR2_X1 U451 ( .A1(n524), .A2(n523), .ZN(n528) );
  AND2_X1 U451bar ( .A1(n524bar), .A2(n523bar), .ZN(n528bar) );
  OR2_X1 U452 ( .A1(in_24), .A2(in[97]), .ZN(n523) );
  AND2_X1 U452bar ( .A1(in_24bar), .A2(inbar[97]), .ZN(n523bar) );
  OR2_X1 U453 ( .A1(in_33), .A2(in_27), .ZN(n524) );
  AND2_X1 U453bar ( .A1(in_33bar), .A2(in_27bar), .ZN(n524bar) );
  OR2_X1 U454 ( .A1(n522), .A2(n521), .ZN(n568) );
  AND2_X1 U454bar ( .A1(n522bar), .A2(n521bar), .ZN(n568bar) );
  OR2_X1 U455 ( .A1(in[145]), .A2(in[126]), .ZN(n521) );
  AND2_X1 U455bar ( .A1(inbar[145]), .A2(inbar[126]), .ZN(n521bar) );
  OR2_X1 U456 ( .A1(in[169]), .A2(n520), .ZN(n522) );
  AND2_X1 U456bar ( .A1(inbar[169]), .A2(n520bar), .ZN(n522bar) );
  OR2_X1 U457 ( .A1(in[221]), .A2(in[172]), .ZN(n520) );
  AND2_X1 U457bar ( .A1(inbar[221]), .A2(inbar[172]), .ZN(n520bar) );
  OR2_X1 U458 ( .A1(n519), .A2(n518), .ZN(n570) );
  AND2_X1 U458bar ( .A1(n519bar), .A2(n518bar), .ZN(n570bar) );
  OR2_X1 U459 ( .A1(n517), .A2(n516), .ZN(n518) );
  AND2_X1 U459bar ( .A1(n517bar), .A2(n516bar), .ZN(n518bar) );
  OR2_X1 U460 ( .A1(in[241]), .A2(in[224]), .ZN(n516) );
  AND2_X1 U460bar ( .A1(inbar[241]), .A2(inbar[224]), .ZN(n516bar) );
  OR2_X1 U461 ( .A1(in[86]), .A2(n515), .ZN(n517) );
  AND2_X1 U461bar ( .A1(inbar[86]), .A2(n515bar), .ZN(n517bar) );
  OR2_X1 U462 ( .A1(in_43), .A2(in_34), .ZN(n515) );
  AND2_X1 U462bar ( .A1(in_43bar), .A2(in_34bar), .ZN(n515bar) );
  OR2_X1 U463 ( .A1(n514), .A2(n513), .ZN(n519) );
  AND2_X1 U463bar ( .A1(n514bar), .A2(n513bar), .ZN(n519bar) );
  OR2_X1 U464 ( .A1(in_65), .A2(in_51), .ZN(n513) );
  AND2_X1 U464bar ( .A1(in_65bar), .A2(in_51bar), .ZN(n513bar) );
  OR2_X1 U465 ( .A1(in_75), .A2(n512), .ZN(n514) );
  AND2_X1 U465bar ( .A1(in_75bar), .A2(n512bar), .ZN(n514bar) );
  OR2_X1 U466 ( .A1(in_81), .A2(in_77), .ZN(n512) );
  AND2_X1 U466bar ( .A1(in_81bar), .A2(in_77bar), .ZN(n512bar) );
  OR2_X1 U467 ( .A1(n511), .A2(n510), .ZN(n778) );
  AND2_X1 U467bar ( .A1(n511bar), .A2(n510bar), .ZN(n778bar) );
  OR2_X1 U468 ( .A1(n509), .A2(n508), .ZN(n510) );
  AND2_X1 U468bar ( .A1(n509bar), .A2(n508bar), .ZN(n510bar) );
  OR2_X1 U469 ( .A1(n507), .A2(n506), .ZN(n508) );
  AND2_X1 U469bar ( .A1(n507bar), .A2(n506bar), .ZN(n508bar) );
  OR2_X1 U470 ( .A1(in[107]), .A2(in[101]), .ZN(n506) );
  AND2_X1 U470bar ( .A1(inbar[107]), .A2(inbar[101]), .ZN(n506bar) );
  OR2_X1 U471 ( .A1(in[139]), .A2(in[132]), .ZN(n507) );
  AND2_X1 U471bar ( .A1(inbar[139]), .A2(inbar[132]), .ZN(n507bar) );
  OR2_X1 U472 ( .A1(n505), .A2(n504), .ZN(n509) );
  AND2_X1 U472bar ( .A1(n505bar), .A2(n504bar), .ZN(n509bar) );
  OR2_X1 U473 ( .A1(in[146]), .A2(in[141]), .ZN(n504) );
  AND2_X1 U473bar ( .A1(inbar[146]), .A2(inbar[141]), .ZN(n504bar) );
  OR2_X1 U474 ( .A1(in[203]), .A2(in[179]), .ZN(n505) );
  AND2_X1 U474bar ( .A1(inbar[203]), .A2(inbar[179]), .ZN(n505bar) );
  OR2_X1 U475 ( .A1(n503), .A2(n502), .ZN(n511) );
  AND2_X1 U475bar ( .A1(n503bar), .A2(n502bar), .ZN(n511bar) );
  OR2_X1 U476 ( .A1(n501), .A2(n500), .ZN(n502) );
  AND2_X1 U476bar ( .A1(n501bar), .A2(n500bar), .ZN(n502bar) );
  OR2_X1 U477 ( .A1(in[243]), .A2(in[222]), .ZN(n500) );
  AND2_X1 U477bar ( .A1(inbar[243]), .A2(inbar[222]), .ZN(n500bar) );
  OR2_X1 U478 ( .A1(in[251]), .A2(in[250]), .ZN(n501) );
  AND2_X1 U478bar ( .A1(inbar[251]), .A2(inbar[250]), .ZN(n501bar) );
  OR2_X1 U479 ( .A1(n499), .A2(n498), .ZN(n503) );
  AND2_X1 U479bar ( .A1(n499bar), .A2(n498bar), .ZN(n503bar) );
  OR2_X1 U480 ( .A1(in_37), .A2(in_19), .ZN(n498) );
  AND2_X1 U480bar ( .A1(in_37bar), .A2(in_19bar), .ZN(n498bar) );
  OR2_X1 U481 ( .A1(in_78), .A2(in_6), .ZN(n499) );
  AND2_X1 U481bar ( .A1(in_78bar), .A2(in_6bar), .ZN(n499bar) );
  OR2_X1 U482 ( .A1(n497), .A2(n496), .ZN(n603) );
  AND2_X1 U482bar ( .A1(n497bar), .A2(n496bar), .ZN(n603bar) );
  OR2_X1 U483 ( .A1(in[112]), .A2(in[102]), .ZN(n496) );
  AND2_X1 U483bar ( .A1(inbar[112]), .A2(inbar[102]), .ZN(n496bar) );
  OR2_X1 U484 ( .A1(in[123]), .A2(n495), .ZN(n497) );
  AND2_X1 U484bar ( .A1(inbar[123]), .A2(n495bar), .ZN(n497bar) );
  OR2_X1 U485 ( .A1(in[143]), .A2(in[130]), .ZN(n495) );
  AND2_X1 U485bar ( .A1(inbar[143]), .A2(inbar[130]), .ZN(n495bar) );
  OR2_X1 U486 ( .A1(n494), .A2(n493), .ZN(n605) );
  AND2_X1 U486bar ( .A1(n494bar), .A2(n493bar), .ZN(n605bar) );
  OR2_X1 U487 ( .A1(n492), .A2(n491), .ZN(n493) );
  AND2_X1 U487bar ( .A1(n492bar), .A2(n491bar), .ZN(n493bar) );
  OR2_X1 U488 ( .A1(in[216]), .A2(in[213]), .ZN(n491) );
  AND2_X1 U488bar ( .A1(inbar[216]), .A2(inbar[213]), .ZN(n491bar) );
  OR2_X1 U489 ( .A1(in[227]), .A2(n490), .ZN(n492) );
  AND2_X1 U489bar ( .A1(inbar[227]), .A2(n490bar), .ZN(n492bar) );
  OR2_X1 U490 ( .A1(in_0), .A2(in[248]), .ZN(n490) );
  AND2_X1 U490bar ( .A1(in_0bar), .A2(inbar[248]), .ZN(n490bar) );
  OR2_X1 U491 ( .A1(n489), .A2(n488), .ZN(n494) );
  AND2_X1 U491bar ( .A1(n489bar), .A2(n488bar), .ZN(n494bar) );
  OR2_X1 U492 ( .A1(in_46), .A2(in_44), .ZN(n488) );
  AND2_X1 U492bar ( .A1(in_46bar), .A2(in_44bar), .ZN(n488bar) );
  OR2_X1 U493 ( .A1(in_50), .A2(n487), .ZN(n489) );
  AND2_X1 U493bar ( .A1(in_50bar), .A2(n487bar), .ZN(n489bar) );
  OR2_X1 U494 ( .A1(in_9), .A2(in_80), .ZN(n487) );
  AND2_X1 U494bar ( .A1(in_9bar), .A2(in_80bar), .ZN(n487bar) );
endmodule

module sBox_4 ( in, inbar, out, outbar );

  input wire [7:0] in;
  input wire [7:0] inbar;
//input_done

  output wire [7:0] out;
  output wire [7:0] outbar;
//output_done

  wire [255:0] decodeOut;
  wire [255:0] decodeOutbar;
//wire_done

  decode_4 dec ( .in(in), .inbar(inbar), .out(decodeOut), .outbar(decodeOutbar) );
  encode_4 enc ( .in(decodeOut), .inbar(decodeOutbar), .out(out), .outbar(outbar) );
endmodule

module CD2_17 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD2_18 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD2_19 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD2_20 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD4_9 ( a, abar, b, bbar, y, ybar );

  input wire [3:0] a;
  input wire [3:0] b;
  input wire [3:0] abar;
  input wire [3:0] bbar;
//input_done

  output wire [15:0] y;
  output wire [15:0] ybar;
//output_done

//wire_done

  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]) );
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]) );
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]) );
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]) );
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]) );
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]) );
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]) );
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]) );
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]) );
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]) );
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]) );
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]) );
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]) );
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]) );
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]) );
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]) );
endmodule

module CD4_10 ( a, abar, b, bbar, y, ybar );

  input wire [3:0] a;
  input wire [3:0] b;
  input wire [3:0] abar;
  input wire [3:0] bbar;
//input_done

  output wire [15:0] y;
  output wire [15:0] ybar;
//output_done

//wire_done

  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]) );
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]) );
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]) );
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]) );
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]) );
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]) );
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]) );
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]) );
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]) );
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]) );
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]) );
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]) );
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]) );
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]) );
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]) );
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]) );
endmodule

module CD16_5 ( a, abar, b, bbar, y, ybar );

  input wire [15:0] a;
  input wire [15:0] b;
  input wire [15:0] abar;
  input wire [15:0] bbar;
//input_done

  output wire [255:0] y;
  output wire [255:0] ybar;
//output_done

//wire_done

  AND2_X1 U1 ( .A1(b[9]), .A2(a[0]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[9]), .A2(abar[0]), .ZN(ybar[9]) );
  AND2_X1 U2 ( .A1(b[3]), .A2(a[6]), .ZN(y[99]) );
  OR2_X1 U2bar ( .A1(bbar[3]), .A2(abar[6]), .ZN(ybar[99]) );
  AND2_X1 U3 ( .A1(b[2]), .A2(a[6]), .ZN(y[98]) );
  OR2_X1 U3bar ( .A1(bbar[2]), .A2(abar[6]), .ZN(ybar[98]) );
  AND2_X1 U4 ( .A1(b[1]), .A2(a[6]), .ZN(y[97]) );
  OR2_X1 U4bar ( .A1(bbar[1]), .A2(abar[6]), .ZN(ybar[97]) );
  AND2_X1 U5 ( .A1(b[0]), .A2(a[6]), .ZN(y[96]) );
  OR2_X1 U5bar ( .A1(bbar[0]), .A2(abar[6]), .ZN(ybar[96]) );
  AND2_X1 U6 ( .A1(b[15]), .A2(a[5]), .ZN(y[95]) );
  OR2_X1 U6bar ( .A1(bbar[15]), .A2(abar[5]), .ZN(ybar[95]) );
  AND2_X1 U7 ( .A1(b[14]), .A2(a[5]), .ZN(y[94]) );
  OR2_X1 U7bar ( .A1(bbar[14]), .A2(abar[5]), .ZN(ybar[94]) );
  AND2_X1 U8 ( .A1(b[13]), .A2(a[5]), .ZN(y[93]) );
  OR2_X1 U8bar ( .A1(bbar[13]), .A2(abar[5]), .ZN(ybar[93]) );
  AND2_X1 U9 ( .A1(b[12]), .A2(a[5]), .ZN(y[92]) );
  OR2_X1 U9bar ( .A1(bbar[12]), .A2(abar[5]), .ZN(ybar[92]) );
  AND2_X1 U10 ( .A1(b[11]), .A2(a[5]), .ZN(y[91]) );
  OR2_X1 U10bar ( .A1(bbar[11]), .A2(abar[5]), .ZN(ybar[91]) );
  AND2_X1 U11 ( .A1(b[10]), .A2(a[5]), .ZN(y[90]) );
  OR2_X1 U11bar ( .A1(bbar[10]), .A2(abar[5]), .ZN(ybar[90]) );
  AND2_X1 U12 ( .A1(b[8]), .A2(a[0]), .ZN(y[8]) );
  OR2_X1 U12bar ( .A1(bbar[8]), .A2(abar[0]), .ZN(ybar[8]) );
  AND2_X1 U13 ( .A1(a[5]), .A2(b[9]), .ZN(y[89]) );
  OR2_X1 U13bar ( .A1(abar[5]), .A2(bbar[9]), .ZN(ybar[89]) );
  AND2_X1 U14 ( .A1(b[8]), .A2(a[5]), .ZN(y[88]) );
  OR2_X1 U14bar ( .A1(bbar[8]), .A2(abar[5]), .ZN(ybar[88]) );
  AND2_X1 U15 ( .A1(b[7]), .A2(a[5]), .ZN(y[87]) );
  OR2_X1 U15bar ( .A1(bbar[7]), .A2(abar[5]), .ZN(ybar[87]) );
  AND2_X1 U16 ( .A1(b[6]), .A2(a[5]), .ZN(y[86]) );
  OR2_X1 U16bar ( .A1(bbar[6]), .A2(abar[5]), .ZN(ybar[86]) );
  AND2_X1 U17 ( .A1(b[5]), .A2(a[5]), .ZN(y[85]) );
  OR2_X1 U17bar ( .A1(bbar[5]), .A2(abar[5]), .ZN(ybar[85]) );
  AND2_X1 U18 ( .A1(b[4]), .A2(a[5]), .ZN(y[84]) );
  OR2_X1 U18bar ( .A1(bbar[4]), .A2(abar[5]), .ZN(ybar[84]) );
  AND2_X1 U19 ( .A1(a[5]), .A2(b[3]), .ZN(y[83]) );
  OR2_X1 U19bar ( .A1(abar[5]), .A2(bbar[3]), .ZN(ybar[83]) );
  AND2_X1 U20 ( .A1(a[5]), .A2(b[2]), .ZN(y[82]) );
  OR2_X1 U20bar ( .A1(abar[5]), .A2(bbar[2]), .ZN(ybar[82]) );
  AND2_X1 U21 ( .A1(a[5]), .A2(b[1]), .ZN(y[81]) );
  OR2_X1 U21bar ( .A1(abar[5]), .A2(bbar[1]), .ZN(ybar[81]) );
  AND2_X1 U22 ( .A1(a[5]), .A2(b[0]), .ZN(y[80]) );
  OR2_X1 U22bar ( .A1(abar[5]), .A2(bbar[0]), .ZN(ybar[80]) );
  AND2_X1 U23 ( .A1(b[7]), .A2(a[0]), .ZN(y[7]) );
  OR2_X1 U23bar ( .A1(bbar[7]), .A2(abar[0]), .ZN(ybar[7]) );
  AND2_X1 U24 ( .A1(a[4]), .A2(b[15]), .ZN(y[79]) );
  OR2_X1 U24bar ( .A1(abar[4]), .A2(bbar[15]), .ZN(ybar[79]) );
  AND2_X1 U25 ( .A1(a[4]), .A2(b[14]), .ZN(y[78]) );
  OR2_X1 U25bar ( .A1(abar[4]), .A2(bbar[14]), .ZN(ybar[78]) );
  AND2_X1 U26 ( .A1(a[4]), .A2(b[13]), .ZN(y[77]) );
  OR2_X1 U26bar ( .A1(abar[4]), .A2(bbar[13]), .ZN(ybar[77]) );
  AND2_X1 U27 ( .A1(a[4]), .A2(b[12]), .ZN(y[76]) );
  OR2_X1 U27bar ( .A1(abar[4]), .A2(bbar[12]), .ZN(ybar[76]) );
  AND2_X1 U28 ( .A1(a[4]), .A2(b[11]), .ZN(y[75]) );
  OR2_X1 U28bar ( .A1(abar[4]), .A2(bbar[11]), .ZN(ybar[75]) );
  AND2_X1 U29 ( .A1(a[4]), .A2(b[10]), .ZN(y[74]) );
  OR2_X1 U29bar ( .A1(abar[4]), .A2(bbar[10]), .ZN(ybar[74]) );
  AND2_X1 U30 ( .A1(a[4]), .A2(b[9]), .ZN(y[73]) );
  OR2_X1 U30bar ( .A1(abar[4]), .A2(bbar[9]), .ZN(ybar[73]) );
  AND2_X1 U31 ( .A1(a[4]), .A2(b[8]), .ZN(y[72]) );
  OR2_X1 U31bar ( .A1(abar[4]), .A2(bbar[8]), .ZN(ybar[72]) );
  AND2_X1 U32 ( .A1(a[4]), .A2(b[7]), .ZN(y[71]) );
  OR2_X1 U32bar ( .A1(abar[4]), .A2(bbar[7]), .ZN(ybar[71]) );
  AND2_X1 U33 ( .A1(a[4]), .A2(b[6]), .ZN(y[70]) );
  OR2_X1 U33bar ( .A1(abar[4]), .A2(bbar[6]), .ZN(ybar[70]) );
  AND2_X1 U34 ( .A1(b[6]), .A2(a[0]), .ZN(y[6]) );
  OR2_X1 U34bar ( .A1(bbar[6]), .A2(abar[0]), .ZN(ybar[6]) );
  AND2_X1 U35 ( .A1(a[4]), .A2(b[5]), .ZN(y[69]) );
  OR2_X1 U35bar ( .A1(abar[4]), .A2(bbar[5]), .ZN(ybar[69]) );
  AND2_X1 U36 ( .A1(a[4]), .A2(b[4]), .ZN(y[68]) );
  OR2_X1 U36bar ( .A1(abar[4]), .A2(bbar[4]), .ZN(ybar[68]) );
  AND2_X1 U37 ( .A1(a[4]), .A2(b[3]), .ZN(y[67]) );
  OR2_X1 U37bar ( .A1(abar[4]), .A2(bbar[3]), .ZN(ybar[67]) );
  AND2_X1 U38 ( .A1(a[4]), .A2(b[2]), .ZN(y[66]) );
  OR2_X1 U38bar ( .A1(abar[4]), .A2(bbar[2]), .ZN(ybar[66]) );
  AND2_X1 U39 ( .A1(a[4]), .A2(b[1]), .ZN(y[65]) );
  OR2_X1 U39bar ( .A1(abar[4]), .A2(bbar[1]), .ZN(ybar[65]) );
  AND2_X1 U40 ( .A1(a[4]), .A2(b[0]), .ZN(y[64]) );
  OR2_X1 U40bar ( .A1(abar[4]), .A2(bbar[0]), .ZN(ybar[64]) );
  AND2_X1 U41 ( .A1(a[3]), .A2(b[15]), .ZN(y[63]) );
  OR2_X1 U41bar ( .A1(abar[3]), .A2(bbar[15]), .ZN(ybar[63]) );
  AND2_X1 U42 ( .A1(a[3]), .A2(b[14]), .ZN(y[62]) );
  OR2_X1 U42bar ( .A1(abar[3]), .A2(bbar[14]), .ZN(ybar[62]) );
  AND2_X1 U43 ( .A1(a[3]), .A2(b[13]), .ZN(y[61]) );
  OR2_X1 U43bar ( .A1(abar[3]), .A2(bbar[13]), .ZN(ybar[61]) );
  AND2_X1 U44 ( .A1(a[3]), .A2(b[12]), .ZN(y[60]) );
  OR2_X1 U44bar ( .A1(abar[3]), .A2(bbar[12]), .ZN(ybar[60]) );
  AND2_X1 U45 ( .A1(b[5]), .A2(a[0]), .ZN(y[5]) );
  OR2_X1 U45bar ( .A1(bbar[5]), .A2(abar[0]), .ZN(ybar[5]) );
  AND2_X1 U46 ( .A1(a[3]), .A2(b[11]), .ZN(y[59]) );
  OR2_X1 U46bar ( .A1(abar[3]), .A2(bbar[11]), .ZN(ybar[59]) );
  AND2_X1 U47 ( .A1(a[3]), .A2(b[10]), .ZN(y[58]) );
  OR2_X1 U47bar ( .A1(abar[3]), .A2(bbar[10]), .ZN(ybar[58]) );
  AND2_X1 U48 ( .A1(a[3]), .A2(b[9]), .ZN(y[57]) );
  OR2_X1 U48bar ( .A1(abar[3]), .A2(bbar[9]), .ZN(ybar[57]) );
  AND2_X1 U49 ( .A1(a[3]), .A2(b[8]), .ZN(y[56]) );
  OR2_X1 U49bar ( .A1(abar[3]), .A2(bbar[8]), .ZN(ybar[56]) );
  AND2_X1 U50 ( .A1(a[3]), .A2(b[7]), .ZN(y[55]) );
  OR2_X1 U50bar ( .A1(abar[3]), .A2(bbar[7]), .ZN(ybar[55]) );
  AND2_X1 U51 ( .A1(a[3]), .A2(b[6]), .ZN(y[54]) );
  OR2_X1 U51bar ( .A1(abar[3]), .A2(bbar[6]), .ZN(ybar[54]) );
  AND2_X1 U52 ( .A1(a[3]), .A2(b[5]), .ZN(y[53]) );
  OR2_X1 U52bar ( .A1(abar[3]), .A2(bbar[5]), .ZN(ybar[53]) );
  AND2_X1 U53 ( .A1(a[3]), .A2(b[4]), .ZN(y[52]) );
  OR2_X1 U53bar ( .A1(abar[3]), .A2(bbar[4]), .ZN(ybar[52]) );
  AND2_X1 U54 ( .A1(a[3]), .A2(b[3]), .ZN(y[51]) );
  OR2_X1 U54bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[51]) );
  AND2_X1 U55 ( .A1(a[3]), .A2(b[2]), .ZN(y[50]) );
  OR2_X1 U55bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[50]) );
  AND2_X1 U56 ( .A1(b[4]), .A2(a[0]), .ZN(y[4]) );
  OR2_X1 U56bar ( .A1(bbar[4]), .A2(abar[0]), .ZN(ybar[4]) );
  AND2_X1 U57 ( .A1(a[3]), .A2(b[1]), .ZN(y[49]) );
  OR2_X1 U57bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[49]) );
  AND2_X1 U58 ( .A1(a[3]), .A2(b[0]), .ZN(y[48]) );
  OR2_X1 U58bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[48]) );
  AND2_X1 U59 ( .A1(a[2]), .A2(b[15]), .ZN(y[47]) );
  OR2_X1 U59bar ( .A1(abar[2]), .A2(bbar[15]), .ZN(ybar[47]) );
  AND2_X1 U60 ( .A1(a[2]), .A2(b[14]), .ZN(y[46]) );
  OR2_X1 U60bar ( .A1(abar[2]), .A2(bbar[14]), .ZN(ybar[46]) );
  AND2_X1 U61 ( .A1(a[2]), .A2(b[13]), .ZN(y[45]) );
  OR2_X1 U61bar ( .A1(abar[2]), .A2(bbar[13]), .ZN(ybar[45]) );
  AND2_X1 U62 ( .A1(a[2]), .A2(b[12]), .ZN(y[44]) );
  OR2_X1 U62bar ( .A1(abar[2]), .A2(bbar[12]), .ZN(ybar[44]) );
  AND2_X1 U63 ( .A1(a[2]), .A2(b[11]), .ZN(y[43]) );
  OR2_X1 U63bar ( .A1(abar[2]), .A2(bbar[11]), .ZN(ybar[43]) );
  AND2_X1 U64 ( .A1(a[2]), .A2(b[10]), .ZN(y[42]) );
  OR2_X1 U64bar ( .A1(abar[2]), .A2(bbar[10]), .ZN(ybar[42]) );
  AND2_X1 U65 ( .A1(a[2]), .A2(b[9]), .ZN(y[41]) );
  OR2_X1 U65bar ( .A1(abar[2]), .A2(bbar[9]), .ZN(ybar[41]) );
  AND2_X1 U66 ( .A1(a[2]), .A2(b[8]), .ZN(y[40]) );
  OR2_X1 U66bar ( .A1(abar[2]), .A2(bbar[8]), .ZN(ybar[40]) );
  AND2_X1 U67 ( .A1(b[3]), .A2(a[0]), .ZN(y[3]) );
  OR2_X1 U67bar ( .A1(bbar[3]), .A2(abar[0]), .ZN(ybar[3]) );
  AND2_X1 U68 ( .A1(a[2]), .A2(b[7]), .ZN(y[39]) );
  OR2_X1 U68bar ( .A1(abar[2]), .A2(bbar[7]), .ZN(ybar[39]) );
  AND2_X1 U69 ( .A1(a[2]), .A2(b[6]), .ZN(y[38]) );
  OR2_X1 U69bar ( .A1(abar[2]), .A2(bbar[6]), .ZN(ybar[38]) );
  AND2_X1 U70 ( .A1(a[2]), .A2(b[5]), .ZN(y[37]) );
  OR2_X1 U70bar ( .A1(abar[2]), .A2(bbar[5]), .ZN(ybar[37]) );
  AND2_X1 U71 ( .A1(a[2]), .A2(b[4]), .ZN(y[36]) );
  OR2_X1 U71bar ( .A1(abar[2]), .A2(bbar[4]), .ZN(ybar[36]) );
  AND2_X1 U72 ( .A1(a[2]), .A2(b[3]), .ZN(y[35]) );
  OR2_X1 U72bar ( .A1(abar[2]), .A2(bbar[3]), .ZN(ybar[35]) );
  AND2_X1 U73 ( .A1(a[2]), .A2(b[2]), .ZN(y[34]) );
  OR2_X1 U73bar ( .A1(abar[2]), .A2(bbar[2]), .ZN(ybar[34]) );
  AND2_X1 U74 ( .A1(a[2]), .A2(b[1]), .ZN(y[33]) );
  OR2_X1 U74bar ( .A1(abar[2]), .A2(bbar[1]), .ZN(ybar[33]) );
  AND2_X1 U75 ( .A1(a[2]), .A2(b[0]), .ZN(y[32]) );
  OR2_X1 U75bar ( .A1(abar[2]), .A2(bbar[0]), .ZN(ybar[32]) );
  AND2_X1 U76 ( .A1(a[1]), .A2(b[15]), .ZN(y[31]) );
  OR2_X1 U76bar ( .A1(abar[1]), .A2(bbar[15]), .ZN(ybar[31]) );
  AND2_X1 U77 ( .A1(a[1]), .A2(b[14]), .ZN(y[30]) );
  OR2_X1 U77bar ( .A1(abar[1]), .A2(bbar[14]), .ZN(ybar[30]) );
  AND2_X1 U78 ( .A1(b[2]), .A2(a[0]), .ZN(y[2]) );
  OR2_X1 U78bar ( .A1(bbar[2]), .A2(abar[0]), .ZN(ybar[2]) );
  AND2_X1 U79 ( .A1(a[1]), .A2(b[13]), .ZN(y[29]) );
  OR2_X1 U79bar ( .A1(abar[1]), .A2(bbar[13]), .ZN(ybar[29]) );
  AND2_X1 U80 ( .A1(a[1]), .A2(b[12]), .ZN(y[28]) );
  OR2_X1 U80bar ( .A1(abar[1]), .A2(bbar[12]), .ZN(ybar[28]) );
  AND2_X1 U81 ( .A1(a[1]), .A2(b[11]), .ZN(y[27]) );
  OR2_X1 U81bar ( .A1(abar[1]), .A2(bbar[11]), .ZN(ybar[27]) );
  AND2_X1 U82 ( .A1(a[1]), .A2(b[10]), .ZN(y[26]) );
  OR2_X1 U82bar ( .A1(abar[1]), .A2(bbar[10]), .ZN(ybar[26]) );
  AND2_X1 U83 ( .A1(a[1]), .A2(b[9]), .ZN(y[25]) );
  OR2_X1 U83bar ( .A1(abar[1]), .A2(bbar[9]), .ZN(ybar[25]) );
  AND2_X1 U84 ( .A1(a[15]), .A2(b[15]), .ZN(y[255]) );
  OR2_X1 U84bar ( .A1(abar[15]), .A2(bbar[15]), .ZN(ybar[255]) );
  AND2_X1 U85 ( .A1(a[15]), .A2(b[14]), .ZN(y[254]) );
  OR2_X1 U85bar ( .A1(abar[15]), .A2(bbar[14]), .ZN(ybar[254]) );
  AND2_X1 U86 ( .A1(a[15]), .A2(b[13]), .ZN(y[253]) );
  OR2_X1 U86bar ( .A1(abar[15]), .A2(bbar[13]), .ZN(ybar[253]) );
  AND2_X1 U87 ( .A1(a[15]), .A2(b[12]), .ZN(y[252]) );
  OR2_X1 U87bar ( .A1(abar[15]), .A2(bbar[12]), .ZN(ybar[252]) );
  AND2_X1 U88 ( .A1(a[15]), .A2(b[11]), .ZN(y[251]) );
  OR2_X1 U88bar ( .A1(abar[15]), .A2(bbar[11]), .ZN(ybar[251]) );
  AND2_X1 U89 ( .A1(a[15]), .A2(b[10]), .ZN(y[250]) );
  OR2_X1 U89bar ( .A1(abar[15]), .A2(bbar[10]), .ZN(ybar[250]) );
  AND2_X1 U90 ( .A1(a[1]), .A2(b[8]), .ZN(y[24]) );
  OR2_X1 U90bar ( .A1(abar[1]), .A2(bbar[8]), .ZN(ybar[24]) );
  AND2_X1 U91 ( .A1(a[15]), .A2(b[9]), .ZN(y[249]) );
  OR2_X1 U91bar ( .A1(abar[15]), .A2(bbar[9]), .ZN(ybar[249]) );
  AND2_X1 U92 ( .A1(a[15]), .A2(b[8]), .ZN(y[248]) );
  OR2_X1 U92bar ( .A1(abar[15]), .A2(bbar[8]), .ZN(ybar[248]) );
  AND2_X1 U93 ( .A1(a[15]), .A2(b[7]), .ZN(y[247]) );
  OR2_X1 U93bar ( .A1(abar[15]), .A2(bbar[7]), .ZN(ybar[247]) );
  AND2_X1 U94 ( .A1(a[15]), .A2(b[6]), .ZN(y[246]) );
  OR2_X1 U94bar ( .A1(abar[15]), .A2(bbar[6]), .ZN(ybar[246]) );
  AND2_X1 U95 ( .A1(a[15]), .A2(b[5]), .ZN(y[245]) );
  OR2_X1 U95bar ( .A1(abar[15]), .A2(bbar[5]), .ZN(ybar[245]) );
  AND2_X1 U96 ( .A1(a[15]), .A2(b[4]), .ZN(y[244]) );
  OR2_X1 U96bar ( .A1(abar[15]), .A2(bbar[4]), .ZN(ybar[244]) );
  AND2_X1 U97 ( .A1(a[15]), .A2(b[3]), .ZN(y[243]) );
  OR2_X1 U97bar ( .A1(abar[15]), .A2(bbar[3]), .ZN(ybar[243]) );
  AND2_X1 U98 ( .A1(a[15]), .A2(b[2]), .ZN(y[242]) );
  OR2_X1 U98bar ( .A1(abar[15]), .A2(bbar[2]), .ZN(ybar[242]) );
  AND2_X1 U99 ( .A1(a[15]), .A2(b[1]), .ZN(y[241]) );
  OR2_X1 U99bar ( .A1(abar[15]), .A2(bbar[1]), .ZN(ybar[241]) );
  AND2_X1 U100 ( .A1(a[15]), .A2(b[0]), .ZN(y[240]) );
  OR2_X1 U100bar ( .A1(abar[15]), .A2(bbar[0]), .ZN(ybar[240]) );
  AND2_X1 U101 ( .A1(a[1]), .A2(b[7]), .ZN(y[23]) );
  OR2_X1 U101bar ( .A1(abar[1]), .A2(bbar[7]), .ZN(ybar[23]) );
  AND2_X1 U102 ( .A1(a[14]), .A2(b[15]), .ZN(y[239]) );
  OR2_X1 U102bar ( .A1(abar[14]), .A2(bbar[15]), .ZN(ybar[239]) );
  AND2_X1 U103 ( .A1(a[14]), .A2(b[14]), .ZN(y[238]) );
  OR2_X1 U103bar ( .A1(abar[14]), .A2(bbar[14]), .ZN(ybar[238]) );
  AND2_X1 U104 ( .A1(a[14]), .A2(b[13]), .ZN(y[237]) );
  OR2_X1 U104bar ( .A1(abar[14]), .A2(bbar[13]), .ZN(ybar[237]) );
  AND2_X1 U105 ( .A1(a[14]), .A2(b[12]), .ZN(y[236]) );
  OR2_X1 U105bar ( .A1(abar[14]), .A2(bbar[12]), .ZN(ybar[236]) );
  AND2_X1 U106 ( .A1(a[14]), .A2(b[11]), .ZN(y[235]) );
  OR2_X1 U106bar ( .A1(abar[14]), .A2(bbar[11]), .ZN(ybar[235]) );
  AND2_X1 U107 ( .A1(a[14]), .A2(b[10]), .ZN(y[234]) );
  OR2_X1 U107bar ( .A1(abar[14]), .A2(bbar[10]), .ZN(ybar[234]) );
  AND2_X1 U108 ( .A1(a[14]), .A2(b[9]), .ZN(y[233]) );
  OR2_X1 U108bar ( .A1(abar[14]), .A2(bbar[9]), .ZN(ybar[233]) );
  AND2_X1 U109 ( .A1(a[14]), .A2(b[8]), .ZN(y[232]) );
  OR2_X1 U109bar ( .A1(abar[14]), .A2(bbar[8]), .ZN(ybar[232]) );
  AND2_X1 U110 ( .A1(a[14]), .A2(b[7]), .ZN(y[231]) );
  OR2_X1 U110bar ( .A1(abar[14]), .A2(bbar[7]), .ZN(ybar[231]) );
  AND2_X1 U111 ( .A1(a[14]), .A2(b[6]), .ZN(y[230]) );
  OR2_X1 U111bar ( .A1(abar[14]), .A2(bbar[6]), .ZN(ybar[230]) );
  AND2_X1 U112 ( .A1(a[1]), .A2(b[6]), .ZN(y[22]) );
  OR2_X1 U112bar ( .A1(abar[1]), .A2(bbar[6]), .ZN(ybar[22]) );
  AND2_X1 U113 ( .A1(a[14]), .A2(b[5]), .ZN(y[229]) );
  OR2_X1 U113bar ( .A1(abar[14]), .A2(bbar[5]), .ZN(ybar[229]) );
  AND2_X1 U114 ( .A1(a[14]), .A2(b[4]), .ZN(y[228]) );
  OR2_X1 U114bar ( .A1(abar[14]), .A2(bbar[4]), .ZN(ybar[228]) );
  AND2_X1 U115 ( .A1(a[14]), .A2(b[3]), .ZN(y[227]) );
  OR2_X1 U115bar ( .A1(abar[14]), .A2(bbar[3]), .ZN(ybar[227]) );
  AND2_X1 U116 ( .A1(a[14]), .A2(b[2]), .ZN(y[226]) );
  OR2_X1 U116bar ( .A1(abar[14]), .A2(bbar[2]), .ZN(ybar[226]) );
  AND2_X1 U117 ( .A1(a[14]), .A2(b[1]), .ZN(y[225]) );
  OR2_X1 U117bar ( .A1(abar[14]), .A2(bbar[1]), .ZN(ybar[225]) );
  AND2_X1 U118 ( .A1(a[14]), .A2(b[0]), .ZN(y[224]) );
  OR2_X1 U118bar ( .A1(abar[14]), .A2(bbar[0]), .ZN(ybar[224]) );
  AND2_X1 U119 ( .A1(a[13]), .A2(b[15]), .ZN(y[223]) );
  OR2_X1 U119bar ( .A1(abar[13]), .A2(bbar[15]), .ZN(ybar[223]) );
  AND2_X1 U120 ( .A1(a[13]), .A2(b[14]), .ZN(y[222]) );
  OR2_X1 U120bar ( .A1(abar[13]), .A2(bbar[14]), .ZN(ybar[222]) );
  AND2_X1 U121 ( .A1(a[13]), .A2(b[13]), .ZN(y[221]) );
  OR2_X1 U121bar ( .A1(abar[13]), .A2(bbar[13]), .ZN(ybar[221]) );
  AND2_X1 U122 ( .A1(a[13]), .A2(b[12]), .ZN(y[220]) );
  OR2_X1 U122bar ( .A1(abar[13]), .A2(bbar[12]), .ZN(ybar[220]) );
  AND2_X1 U123 ( .A1(a[1]), .A2(b[5]), .ZN(y[21]) );
  OR2_X1 U123bar ( .A1(abar[1]), .A2(bbar[5]), .ZN(ybar[21]) );
  AND2_X1 U124 ( .A1(a[13]), .A2(b[11]), .ZN(y[219]) );
  OR2_X1 U124bar ( .A1(abar[13]), .A2(bbar[11]), .ZN(ybar[219]) );
  AND2_X1 U125 ( .A1(a[13]), .A2(b[10]), .ZN(y[218]) );
  OR2_X1 U125bar ( .A1(abar[13]), .A2(bbar[10]), .ZN(ybar[218]) );
  AND2_X1 U126 ( .A1(a[13]), .A2(b[9]), .ZN(y[217]) );
  OR2_X1 U126bar ( .A1(abar[13]), .A2(bbar[9]), .ZN(ybar[217]) );
  AND2_X1 U127 ( .A1(a[13]), .A2(b[8]), .ZN(y[216]) );
  OR2_X1 U127bar ( .A1(abar[13]), .A2(bbar[8]), .ZN(ybar[216]) );
  AND2_X1 U128 ( .A1(a[13]), .A2(b[7]), .ZN(y[215]) );
  OR2_X1 U128bar ( .A1(abar[13]), .A2(bbar[7]), .ZN(ybar[215]) );
  AND2_X1 U129 ( .A1(a[13]), .A2(b[6]), .ZN(y[214]) );
  OR2_X1 U129bar ( .A1(abar[13]), .A2(bbar[6]), .ZN(ybar[214]) );
  AND2_X1 U130 ( .A1(a[13]), .A2(b[5]), .ZN(y[213]) );
  OR2_X1 U130bar ( .A1(abar[13]), .A2(bbar[5]), .ZN(ybar[213]) );
  AND2_X1 U131 ( .A1(a[13]), .A2(b[4]), .ZN(y[212]) );
  OR2_X1 U131bar ( .A1(abar[13]), .A2(bbar[4]), .ZN(ybar[212]) );
  AND2_X1 U132 ( .A1(a[13]), .A2(b[3]), .ZN(y[211]) );
  OR2_X1 U132bar ( .A1(abar[13]), .A2(bbar[3]), .ZN(ybar[211]) );
  AND2_X1 U133 ( .A1(a[13]), .A2(b[2]), .ZN(y[210]) );
  OR2_X1 U133bar ( .A1(abar[13]), .A2(bbar[2]), .ZN(ybar[210]) );
  AND2_X1 U134 ( .A1(a[1]), .A2(b[4]), .ZN(y[20]) );
  OR2_X1 U134bar ( .A1(abar[1]), .A2(bbar[4]), .ZN(ybar[20]) );
  AND2_X1 U135 ( .A1(a[13]), .A2(b[1]), .ZN(y[209]) );
  OR2_X1 U135bar ( .A1(abar[13]), .A2(bbar[1]), .ZN(ybar[209]) );
  AND2_X1 U136 ( .A1(a[13]), .A2(b[0]), .ZN(y[208]) );
  OR2_X1 U136bar ( .A1(abar[13]), .A2(bbar[0]), .ZN(ybar[208]) );
  AND2_X1 U137 ( .A1(a[12]), .A2(b[15]), .ZN(y[207]) );
  OR2_X1 U137bar ( .A1(abar[12]), .A2(bbar[15]), .ZN(ybar[207]) );
  AND2_X1 U138 ( .A1(a[12]), .A2(b[14]), .ZN(y[206]) );
  OR2_X1 U138bar ( .A1(abar[12]), .A2(bbar[14]), .ZN(ybar[206]) );
  AND2_X1 U139 ( .A1(a[12]), .A2(b[13]), .ZN(y[205]) );
  OR2_X1 U139bar ( .A1(abar[12]), .A2(bbar[13]), .ZN(ybar[205]) );
  AND2_X1 U140 ( .A1(a[12]), .A2(b[12]), .ZN(y[204]) );
  OR2_X1 U140bar ( .A1(abar[12]), .A2(bbar[12]), .ZN(ybar[204]) );
  AND2_X1 U141 ( .A1(a[12]), .A2(b[11]), .ZN(y[203]) );
  OR2_X1 U141bar ( .A1(abar[12]), .A2(bbar[11]), .ZN(ybar[203]) );
  AND2_X1 U142 ( .A1(a[12]), .A2(b[10]), .ZN(y[202]) );
  OR2_X1 U142bar ( .A1(abar[12]), .A2(bbar[10]), .ZN(ybar[202]) );
  AND2_X1 U143 ( .A1(a[12]), .A2(b[9]), .ZN(y[201]) );
  OR2_X1 U143bar ( .A1(abar[12]), .A2(bbar[9]), .ZN(ybar[201]) );
  AND2_X1 U144 ( .A1(a[12]), .A2(b[8]), .ZN(y[200]) );
  OR2_X1 U144bar ( .A1(abar[12]), .A2(bbar[8]), .ZN(ybar[200]) );
  AND2_X1 U145 ( .A1(b[1]), .A2(a[0]), .ZN(y[1]) );
  OR2_X1 U145bar ( .A1(bbar[1]), .A2(abar[0]), .ZN(ybar[1]) );
  AND2_X1 U146 ( .A1(a[1]), .A2(b[3]), .ZN(y[19]) );
  OR2_X1 U146bar ( .A1(abar[1]), .A2(bbar[3]), .ZN(ybar[19]) );
  AND2_X1 U147 ( .A1(a[12]), .A2(b[7]), .ZN(y[199]) );
  OR2_X1 U147bar ( .A1(abar[12]), .A2(bbar[7]), .ZN(ybar[199]) );
  AND2_X1 U148 ( .A1(a[12]), .A2(b[6]), .ZN(y[198]) );
  OR2_X1 U148bar ( .A1(abar[12]), .A2(bbar[6]), .ZN(ybar[198]) );
  AND2_X1 U149 ( .A1(a[12]), .A2(b[5]), .ZN(y[197]) );
  OR2_X1 U149bar ( .A1(abar[12]), .A2(bbar[5]), .ZN(ybar[197]) );
  AND2_X1 U150 ( .A1(a[12]), .A2(b[4]), .ZN(y[196]) );
  OR2_X1 U150bar ( .A1(abar[12]), .A2(bbar[4]), .ZN(ybar[196]) );
  AND2_X1 U151 ( .A1(a[12]), .A2(b[3]), .ZN(y[195]) );
  OR2_X1 U151bar ( .A1(abar[12]), .A2(bbar[3]), .ZN(ybar[195]) );
  AND2_X1 U152 ( .A1(a[12]), .A2(b[2]), .ZN(y[194]) );
  OR2_X1 U152bar ( .A1(abar[12]), .A2(bbar[2]), .ZN(ybar[194]) );
  AND2_X1 U153 ( .A1(a[12]), .A2(b[1]), .ZN(y[193]) );
  OR2_X1 U153bar ( .A1(abar[12]), .A2(bbar[1]), .ZN(ybar[193]) );
  AND2_X1 U154 ( .A1(a[12]), .A2(b[0]), .ZN(y[192]) );
  OR2_X1 U154bar ( .A1(abar[12]), .A2(bbar[0]), .ZN(ybar[192]) );
  AND2_X1 U155 ( .A1(a[11]), .A2(b[15]), .ZN(y[191]) );
  OR2_X1 U155bar ( .A1(abar[11]), .A2(bbar[15]), .ZN(ybar[191]) );
  AND2_X1 U156 ( .A1(a[11]), .A2(b[14]), .ZN(y[190]) );
  OR2_X1 U156bar ( .A1(abar[11]), .A2(bbar[14]), .ZN(ybar[190]) );
  AND2_X1 U157 ( .A1(a[1]), .A2(b[2]), .ZN(y[18]) );
  OR2_X1 U157bar ( .A1(abar[1]), .A2(bbar[2]), .ZN(ybar[18]) );
  AND2_X1 U158 ( .A1(a[11]), .A2(b[13]), .ZN(y[189]) );
  OR2_X1 U158bar ( .A1(abar[11]), .A2(bbar[13]), .ZN(ybar[189]) );
  AND2_X1 U159 ( .A1(a[11]), .A2(b[12]), .ZN(y[188]) );
  OR2_X1 U159bar ( .A1(abar[11]), .A2(bbar[12]), .ZN(ybar[188]) );
  AND2_X1 U160 ( .A1(a[11]), .A2(b[11]), .ZN(y[187]) );
  OR2_X1 U160bar ( .A1(abar[11]), .A2(bbar[11]), .ZN(ybar[187]) );
  AND2_X1 U161 ( .A1(a[11]), .A2(b[10]), .ZN(y[186]) );
  OR2_X1 U161bar ( .A1(abar[11]), .A2(bbar[10]), .ZN(ybar[186]) );
  AND2_X1 U162 ( .A1(a[11]), .A2(b[9]), .ZN(y[185]) );
  OR2_X1 U162bar ( .A1(abar[11]), .A2(bbar[9]), .ZN(ybar[185]) );
  AND2_X1 U163 ( .A1(a[11]), .A2(b[8]), .ZN(y[184]) );
  OR2_X1 U163bar ( .A1(abar[11]), .A2(bbar[8]), .ZN(ybar[184]) );
  AND2_X1 U164 ( .A1(a[11]), .A2(b[7]), .ZN(y[183]) );
  OR2_X1 U164bar ( .A1(abar[11]), .A2(bbar[7]), .ZN(ybar[183]) );
  AND2_X1 U165 ( .A1(a[11]), .A2(b[6]), .ZN(y[182]) );
  OR2_X1 U165bar ( .A1(abar[11]), .A2(bbar[6]), .ZN(ybar[182]) );
  AND2_X1 U166 ( .A1(a[11]), .A2(b[5]), .ZN(y[181]) );
  OR2_X1 U166bar ( .A1(abar[11]), .A2(bbar[5]), .ZN(ybar[181]) );
  AND2_X1 U167 ( .A1(a[11]), .A2(b[4]), .ZN(y[180]) );
  OR2_X1 U167bar ( .A1(abar[11]), .A2(bbar[4]), .ZN(ybar[180]) );
  AND2_X1 U168 ( .A1(a[1]), .A2(b[1]), .ZN(y[17]) );
  OR2_X1 U168bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[17]) );
  AND2_X1 U169 ( .A1(a[11]), .A2(b[3]), .ZN(y[179]) );
  OR2_X1 U169bar ( .A1(abar[11]), .A2(bbar[3]), .ZN(ybar[179]) );
  AND2_X1 U170 ( .A1(a[11]), .A2(b[2]), .ZN(y[178]) );
  OR2_X1 U170bar ( .A1(abar[11]), .A2(bbar[2]), .ZN(ybar[178]) );
  AND2_X1 U171 ( .A1(a[11]), .A2(b[1]), .ZN(y[177]) );
  OR2_X1 U171bar ( .A1(abar[11]), .A2(bbar[1]), .ZN(ybar[177]) );
  AND2_X1 U172 ( .A1(a[11]), .A2(b[0]), .ZN(y[176]) );
  OR2_X1 U172bar ( .A1(abar[11]), .A2(bbar[0]), .ZN(ybar[176]) );
  AND2_X1 U173 ( .A1(a[10]), .A2(b[15]), .ZN(y[175]) );
  OR2_X1 U173bar ( .A1(abar[10]), .A2(bbar[15]), .ZN(ybar[175]) );
  AND2_X1 U174 ( .A1(a[10]), .A2(b[14]), .ZN(y[174]) );
  OR2_X1 U174bar ( .A1(abar[10]), .A2(bbar[14]), .ZN(ybar[174]) );
  AND2_X1 U175 ( .A1(a[10]), .A2(b[13]), .ZN(y[173]) );
  OR2_X1 U175bar ( .A1(abar[10]), .A2(bbar[13]), .ZN(ybar[173]) );
  AND2_X1 U176 ( .A1(a[10]), .A2(b[12]), .ZN(y[172]) );
  OR2_X1 U176bar ( .A1(abar[10]), .A2(bbar[12]), .ZN(ybar[172]) );
  AND2_X1 U177 ( .A1(a[10]), .A2(b[11]), .ZN(y[171]) );
  OR2_X1 U177bar ( .A1(abar[10]), .A2(bbar[11]), .ZN(ybar[171]) );
  AND2_X1 U178 ( .A1(a[10]), .A2(b[10]), .ZN(y[170]) );
  OR2_X1 U178bar ( .A1(abar[10]), .A2(bbar[10]), .ZN(ybar[170]) );
  AND2_X1 U179 ( .A1(a[1]), .A2(b[0]), .ZN(y[16]) );
  OR2_X1 U179bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[16]) );
  AND2_X1 U180 ( .A1(a[10]), .A2(b[9]), .ZN(y[169]) );
  OR2_X1 U180bar ( .A1(abar[10]), .A2(bbar[9]), .ZN(ybar[169]) );
  AND2_X1 U181 ( .A1(a[10]), .A2(b[8]), .ZN(y[168]) );
  OR2_X1 U181bar ( .A1(abar[10]), .A2(bbar[8]), .ZN(ybar[168]) );
  AND2_X1 U182 ( .A1(a[10]), .A2(b[7]), .ZN(y[167]) );
  OR2_X1 U182bar ( .A1(abar[10]), .A2(bbar[7]), .ZN(ybar[167]) );
  AND2_X1 U183 ( .A1(a[10]), .A2(b[6]), .ZN(y[166]) );
  OR2_X1 U183bar ( .A1(abar[10]), .A2(bbar[6]), .ZN(ybar[166]) );
  AND2_X1 U184 ( .A1(a[10]), .A2(b[5]), .ZN(y[165]) );
  OR2_X1 U184bar ( .A1(abar[10]), .A2(bbar[5]), .ZN(ybar[165]) );
  AND2_X1 U185 ( .A1(a[10]), .A2(b[4]), .ZN(y[164]) );
  OR2_X1 U185bar ( .A1(abar[10]), .A2(bbar[4]), .ZN(ybar[164]) );
  AND2_X1 U186 ( .A1(a[10]), .A2(b[3]), .ZN(y[163]) );
  OR2_X1 U186bar ( .A1(abar[10]), .A2(bbar[3]), .ZN(ybar[163]) );
  AND2_X1 U187 ( .A1(a[10]), .A2(b[2]), .ZN(y[162]) );
  OR2_X1 U187bar ( .A1(abar[10]), .A2(bbar[2]), .ZN(ybar[162]) );
  AND2_X1 U188 ( .A1(a[10]), .A2(b[1]), .ZN(y[161]) );
  OR2_X1 U188bar ( .A1(abar[10]), .A2(bbar[1]), .ZN(ybar[161]) );
  AND2_X1 U189 ( .A1(a[10]), .A2(b[0]), .ZN(y[160]) );
  OR2_X1 U189bar ( .A1(abar[10]), .A2(bbar[0]), .ZN(ybar[160]) );
  AND2_X1 U190 ( .A1(b[15]), .A2(a[0]), .ZN(y[15]) );
  OR2_X1 U190bar ( .A1(bbar[15]), .A2(abar[0]), .ZN(ybar[15]) );
  AND2_X1 U191 ( .A1(a[9]), .A2(b[15]), .ZN(y[159]) );
  OR2_X1 U191bar ( .A1(abar[9]), .A2(bbar[15]), .ZN(ybar[159]) );
  AND2_X1 U192 ( .A1(a[9]), .A2(b[14]), .ZN(y[158]) );
  OR2_X1 U192bar ( .A1(abar[9]), .A2(bbar[14]), .ZN(ybar[158]) );
  AND2_X1 U193 ( .A1(a[9]), .A2(b[13]), .ZN(y[157]) );
  OR2_X1 U193bar ( .A1(abar[9]), .A2(bbar[13]), .ZN(ybar[157]) );
  AND2_X1 U194 ( .A1(a[9]), .A2(b[12]), .ZN(y[156]) );
  OR2_X1 U194bar ( .A1(abar[9]), .A2(bbar[12]), .ZN(ybar[156]) );
  AND2_X1 U195 ( .A1(a[9]), .A2(b[11]), .ZN(y[155]) );
  OR2_X1 U195bar ( .A1(abar[9]), .A2(bbar[11]), .ZN(ybar[155]) );
  AND2_X1 U196 ( .A1(a[9]), .A2(b[10]), .ZN(y[154]) );
  OR2_X1 U196bar ( .A1(abar[9]), .A2(bbar[10]), .ZN(ybar[154]) );
  AND2_X1 U197 ( .A1(a[9]), .A2(b[9]), .ZN(y[153]) );
  OR2_X1 U197bar ( .A1(abar[9]), .A2(bbar[9]), .ZN(ybar[153]) );
  AND2_X1 U198 ( .A1(a[9]), .A2(b[8]), .ZN(y[152]) );
  OR2_X1 U198bar ( .A1(abar[9]), .A2(bbar[8]), .ZN(ybar[152]) );
  AND2_X1 U199 ( .A1(a[9]), .A2(b[7]), .ZN(y[151]) );
  OR2_X1 U199bar ( .A1(abar[9]), .A2(bbar[7]), .ZN(ybar[151]) );
  AND2_X1 U200 ( .A1(a[9]), .A2(b[6]), .ZN(y[150]) );
  OR2_X1 U200bar ( .A1(abar[9]), .A2(bbar[6]), .ZN(ybar[150]) );
  AND2_X1 U201 ( .A1(b[14]), .A2(a[0]), .ZN(y[14]) );
  OR2_X1 U201bar ( .A1(bbar[14]), .A2(abar[0]), .ZN(ybar[14]) );
  AND2_X1 U202 ( .A1(a[9]), .A2(b[5]), .ZN(y[149]) );
  OR2_X1 U202bar ( .A1(abar[9]), .A2(bbar[5]), .ZN(ybar[149]) );
  AND2_X1 U203 ( .A1(a[9]), .A2(b[4]), .ZN(y[148]) );
  OR2_X1 U203bar ( .A1(abar[9]), .A2(bbar[4]), .ZN(ybar[148]) );
  AND2_X1 U204 ( .A1(a[9]), .A2(b[3]), .ZN(y[147]) );
  OR2_X1 U204bar ( .A1(abar[9]), .A2(bbar[3]), .ZN(ybar[147]) );
  AND2_X1 U205 ( .A1(a[9]), .A2(b[2]), .ZN(y[146]) );
  OR2_X1 U205bar ( .A1(abar[9]), .A2(bbar[2]), .ZN(ybar[146]) );
  AND2_X1 U206 ( .A1(a[9]), .A2(b[1]), .ZN(y[145]) );
  OR2_X1 U206bar ( .A1(abar[9]), .A2(bbar[1]), .ZN(ybar[145]) );
  AND2_X1 U207 ( .A1(a[9]), .A2(b[0]), .ZN(y[144]) );
  OR2_X1 U207bar ( .A1(abar[9]), .A2(bbar[0]), .ZN(ybar[144]) );
  AND2_X1 U208 ( .A1(a[8]), .A2(b[15]), .ZN(y[143]) );
  OR2_X1 U208bar ( .A1(abar[8]), .A2(bbar[15]), .ZN(ybar[143]) );
  AND2_X1 U209 ( .A1(a[8]), .A2(b[14]), .ZN(y[142]) );
  OR2_X1 U209bar ( .A1(abar[8]), .A2(bbar[14]), .ZN(ybar[142]) );
  AND2_X1 U210 ( .A1(a[8]), .A2(b[13]), .ZN(y[141]) );
  OR2_X1 U210bar ( .A1(abar[8]), .A2(bbar[13]), .ZN(ybar[141]) );
  AND2_X1 U211 ( .A1(a[8]), .A2(b[12]), .ZN(y[140]) );
  OR2_X1 U211bar ( .A1(abar[8]), .A2(bbar[12]), .ZN(ybar[140]) );
  AND2_X1 U212 ( .A1(b[13]), .A2(a[0]), .ZN(y[13]) );
  OR2_X1 U212bar ( .A1(bbar[13]), .A2(abar[0]), .ZN(ybar[13]) );
  AND2_X1 U213 ( .A1(a[8]), .A2(b[11]), .ZN(y[139]) );
  OR2_X1 U213bar ( .A1(abar[8]), .A2(bbar[11]), .ZN(ybar[139]) );
  AND2_X1 U214 ( .A1(a[8]), .A2(b[10]), .ZN(y[138]) );
  OR2_X1 U214bar ( .A1(abar[8]), .A2(bbar[10]), .ZN(ybar[138]) );
  AND2_X1 U215 ( .A1(a[8]), .A2(b[9]), .ZN(y[137]) );
  OR2_X1 U215bar ( .A1(abar[8]), .A2(bbar[9]), .ZN(ybar[137]) );
  AND2_X1 U216 ( .A1(a[8]), .A2(b[8]), .ZN(y[136]) );
  OR2_X1 U216bar ( .A1(abar[8]), .A2(bbar[8]), .ZN(ybar[136]) );
  AND2_X1 U217 ( .A1(a[8]), .A2(b[7]), .ZN(y[135]) );
  OR2_X1 U217bar ( .A1(abar[8]), .A2(bbar[7]), .ZN(ybar[135]) );
  AND2_X1 U218 ( .A1(a[8]), .A2(b[6]), .ZN(y[134]) );
  OR2_X1 U218bar ( .A1(abar[8]), .A2(bbar[6]), .ZN(ybar[134]) );
  AND2_X1 U219 ( .A1(a[8]), .A2(b[5]), .ZN(y[133]) );
  OR2_X1 U219bar ( .A1(abar[8]), .A2(bbar[5]), .ZN(ybar[133]) );
  AND2_X1 U220 ( .A1(a[8]), .A2(b[4]), .ZN(y[132]) );
  OR2_X1 U220bar ( .A1(abar[8]), .A2(bbar[4]), .ZN(ybar[132]) );
  AND2_X1 U221 ( .A1(a[8]), .A2(b[3]), .ZN(y[131]) );
  OR2_X1 U221bar ( .A1(abar[8]), .A2(bbar[3]), .ZN(ybar[131]) );
  AND2_X1 U222 ( .A1(a[8]), .A2(b[2]), .ZN(y[130]) );
  OR2_X1 U222bar ( .A1(abar[8]), .A2(bbar[2]), .ZN(ybar[130]) );
  AND2_X1 U223 ( .A1(b[12]), .A2(a[0]), .ZN(y[12]) );
  OR2_X1 U223bar ( .A1(bbar[12]), .A2(abar[0]), .ZN(ybar[12]) );
  AND2_X1 U224 ( .A1(a[8]), .A2(b[1]), .ZN(y[129]) );
  OR2_X1 U224bar ( .A1(abar[8]), .A2(bbar[1]), .ZN(ybar[129]) );
  AND2_X1 U225 ( .A1(a[8]), .A2(b[0]), .ZN(y[128]) );
  OR2_X1 U225bar ( .A1(abar[8]), .A2(bbar[0]), .ZN(ybar[128]) );
  AND2_X1 U226 ( .A1(a[7]), .A2(b[15]), .ZN(y[127]) );
  OR2_X1 U226bar ( .A1(abar[7]), .A2(bbar[15]), .ZN(ybar[127]) );
  AND2_X1 U227 ( .A1(a[7]), .A2(b[14]), .ZN(y[126]) );
  OR2_X1 U227bar ( .A1(abar[7]), .A2(bbar[14]), .ZN(ybar[126]) );
  AND2_X1 U228 ( .A1(a[7]), .A2(b[13]), .ZN(y[125]) );
  OR2_X1 U228bar ( .A1(abar[7]), .A2(bbar[13]), .ZN(ybar[125]) );
  AND2_X1 U229 ( .A1(a[7]), .A2(b[12]), .ZN(y[124]) );
  OR2_X1 U229bar ( .A1(abar[7]), .A2(bbar[12]), .ZN(ybar[124]) );
  AND2_X1 U230 ( .A1(a[7]), .A2(b[11]), .ZN(y[123]) );
  OR2_X1 U230bar ( .A1(abar[7]), .A2(bbar[11]), .ZN(ybar[123]) );
  AND2_X1 U231 ( .A1(a[7]), .A2(b[10]), .ZN(y[122]) );
  OR2_X1 U231bar ( .A1(abar[7]), .A2(bbar[10]), .ZN(ybar[122]) );
  AND2_X1 U232 ( .A1(a[7]), .A2(b[9]), .ZN(y[121]) );
  OR2_X1 U232bar ( .A1(abar[7]), .A2(bbar[9]), .ZN(ybar[121]) );
  AND2_X1 U233 ( .A1(a[7]), .A2(b[8]), .ZN(y[120]) );
  OR2_X1 U233bar ( .A1(abar[7]), .A2(bbar[8]), .ZN(ybar[120]) );
  AND2_X1 U234 ( .A1(b[11]), .A2(a[0]), .ZN(y[11]) );
  OR2_X1 U234bar ( .A1(bbar[11]), .A2(abar[0]), .ZN(ybar[11]) );
  AND2_X1 U235 ( .A1(a[7]), .A2(b[7]), .ZN(y[119]) );
  OR2_X1 U235bar ( .A1(abar[7]), .A2(bbar[7]), .ZN(ybar[119]) );
  AND2_X1 U236 ( .A1(a[7]), .A2(b[6]), .ZN(y[118]) );
  OR2_X1 U236bar ( .A1(abar[7]), .A2(bbar[6]), .ZN(ybar[118]) );
  AND2_X1 U237 ( .A1(a[7]), .A2(b[5]), .ZN(y[117]) );
  OR2_X1 U237bar ( .A1(abar[7]), .A2(bbar[5]), .ZN(ybar[117]) );
  AND2_X1 U238 ( .A1(a[7]), .A2(b[4]), .ZN(y[116]) );
  OR2_X1 U238bar ( .A1(abar[7]), .A2(bbar[4]), .ZN(ybar[116]) );
  AND2_X1 U239 ( .A1(a[7]), .A2(b[3]), .ZN(y[115]) );
  OR2_X1 U239bar ( .A1(abar[7]), .A2(bbar[3]), .ZN(ybar[115]) );
  AND2_X1 U240 ( .A1(a[7]), .A2(b[2]), .ZN(y[114]) );
  OR2_X1 U240bar ( .A1(abar[7]), .A2(bbar[2]), .ZN(ybar[114]) );
  AND2_X1 U241 ( .A1(a[7]), .A2(b[1]), .ZN(y[113]) );
  OR2_X1 U241bar ( .A1(abar[7]), .A2(bbar[1]), .ZN(ybar[113]) );
  AND2_X1 U242 ( .A1(a[7]), .A2(b[0]), .ZN(y[112]) );
  OR2_X1 U242bar ( .A1(abar[7]), .A2(bbar[0]), .ZN(ybar[112]) );
  AND2_X1 U243 ( .A1(b[15]), .A2(a[6]), .ZN(y[111]) );
  OR2_X1 U243bar ( .A1(bbar[15]), .A2(abar[6]), .ZN(ybar[111]) );
  AND2_X1 U244 ( .A1(b[14]), .A2(a[6]), .ZN(y[110]) );
  OR2_X1 U244bar ( .A1(bbar[14]), .A2(abar[6]), .ZN(ybar[110]) );
  AND2_X1 U245 ( .A1(b[10]), .A2(a[0]), .ZN(y[10]) );
  OR2_X1 U245bar ( .A1(bbar[10]), .A2(abar[0]), .ZN(ybar[10]) );
  AND2_X1 U246 ( .A1(b[13]), .A2(a[6]), .ZN(y[109]) );
  OR2_X1 U246bar ( .A1(bbar[13]), .A2(abar[6]), .ZN(ybar[109]) );
  AND2_X1 U247 ( .A1(b[12]), .A2(a[6]), .ZN(y[108]) );
  OR2_X1 U247bar ( .A1(bbar[12]), .A2(abar[6]), .ZN(ybar[108]) );
  AND2_X1 U248 ( .A1(b[11]), .A2(a[6]), .ZN(y[107]) );
  OR2_X1 U248bar ( .A1(bbar[11]), .A2(abar[6]), .ZN(ybar[107]) );
  AND2_X1 U249 ( .A1(b[10]), .A2(a[6]), .ZN(y[106]) );
  OR2_X1 U249bar ( .A1(bbar[10]), .A2(abar[6]), .ZN(ybar[106]) );
  AND2_X1 U250 ( .A1(a[6]), .A2(b[9]), .ZN(y[105]) );
  OR2_X1 U250bar ( .A1(abar[6]), .A2(bbar[9]), .ZN(ybar[105]) );
  AND2_X1 U251 ( .A1(b[8]), .A2(a[6]), .ZN(y[104]) );
  OR2_X1 U251bar ( .A1(bbar[8]), .A2(abar[6]), .ZN(ybar[104]) );
  AND2_X1 U252 ( .A1(b[7]), .A2(a[6]), .ZN(y[103]) );
  OR2_X1 U252bar ( .A1(bbar[7]), .A2(abar[6]), .ZN(ybar[103]) );
  AND2_X1 U253 ( .A1(b[6]), .A2(a[6]), .ZN(y[102]) );
  OR2_X1 U253bar ( .A1(bbar[6]), .A2(abar[6]), .ZN(ybar[102]) );
  AND2_X1 U254 ( .A1(b[5]), .A2(a[6]), .ZN(y[101]) );
  OR2_X1 U254bar ( .A1(bbar[5]), .A2(abar[6]), .ZN(ybar[101]) );
  AND2_X1 U255 ( .A1(b[4]), .A2(a[6]), .ZN(y[100]) );
  OR2_X1 U255bar ( .A1(bbar[4]), .A2(abar[6]), .ZN(ybar[100]) );
  AND2_X1 U256 ( .A1(b[0]), .A2(a[0]), .ZN(y[0]) );
  OR2_X1 U256bar ( .A1(bbar[0]), .A2(abar[0]), .ZN(ybar[0]) );
endmodule

module decode_5 ( in, inbar, out, outbar );

  input wire [7:0] in;
  input wire [7:0] inbar;
//input_done

  output wire [255:0] out;
  output wire [255:0] outbar;
//output_done

  wire [15:0] level1;
  wire [31:0] level2;
  wire [15:0] level1bar;
  wire [31:0] level2bar;
//wire_done

  CD2_20 cd_l1_1 ( .a(in[1]), .abar(inbar[1]), .b(in[0]), .bbar(inbar[0]), .y(level1[3:0]), .ybar(level1bar[3:0]) );
  CD2_19 cd_l1_2 ( .a(in[3]), .abar(inbar[3]), .b(in[2]), .bbar(inbar[2]), .y(level1[7:4]), .ybar(level1bar[7:4]) );
  CD2_18 cd_l1_3 ( .a(in[5]), .abar(inbar[5]), .b(in[4]), .bbar(inbar[4]), .y(level1[11:8]), .ybar(level1bar[11:8]) );
  CD2_17 cd_l1_4 ( .a(in[7]), .abar(inbar[7]), .b(in[6]), .bbar(inbar[6]), .y(level1[15:12]), .ybar(level1bar[15:12]) );

  CD4_10 cd_l2_1 ( .a(level1[7:4]), .abar(level1bar[7:4]), .b(level1[3:0]), .bbar(level1bar[3:0]), 
        .y(level2[15:0]), .ybar(level2bar[15:0]) );
  CD4_9 cd_l2_2 ( .a(level1[15:12]), .abar(level1bar[15:12]), .b(level1[11:8]), .bbar(level1bar[11:8]), 
        .y(level2[31:16]), .ybar(level2bar[31:16]) );
  CD16_5 cd_l3 ( .a(level2[31:16]), .abar(level2bar[31:16]), .b(level2[15:0]), .bbar(level2bar[15:0]), 
        .y(out), .ybar(outbar) );
endmodule

module encode_5 ( in, inbar, out, outbar );

  input wire [255:0] in;
  input wire [255:0] inbar;
//input_done

  output wire [7:0] out;
  output wire [7:0] outbar;
//output_done

  wire in_81;
  wire in_80;
  wire in_79;
  wire in_78;
  wire in_77;
  wire in_76;
  wire in_75;
  wire in_74;
  wire in_73;
  wire in_72;
  wire in_71;
  wire in_70;
  wire in_69;
  wire in_68;
  wire in_67;
  wire in_66;
  wire in_65;
  wire in_64;
  wire in_63;
  wire in_62;
  wire in_61;
  wire in_60;
  wire in_59;
  wire in_58;
  wire in_57;
  wire in_56;
  wire in_55;
  wire in_54;
  wire in_53;
  wire in_52;
  wire in_51;
  wire in_50;
  wire in_49;
  wire in_48;
  wire in_47;
  wire in_46;
  wire in_45;
  wire in_44;
  wire in_43;
  wire in_42;
  wire in_41;
  wire in_40;
  wire in_39;
  wire in_38;
  wire in_37;
  wire in_36;
  wire in_35;
  wire in_34;
  wire in_33;
  wire in_32;
  wire in_31;
  wire in_30;
  wire in_29;
  wire in_28;
  wire in_27;
  wire in_26;
  wire in_25;
  wire in_24;
  wire in_23;
  wire in_22;
  wire in_21;
  wire in_20;
  wire in_19;
  wire in_18;
  wire in_17;
  wire in_16;
  wire in_15;
  wire in_14;
  wire in_13;
  wire in_12;
  wire in_11;
  wire in_10;
  wire in_9;
  wire in_8;
  wire in_7;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_3;
  wire in_2;
  wire in_1;
  wire in_0;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire in_81bar;
  wire in_80bar;
  wire in_79bar;
  wire in_78bar;
  wire in_77bar;
  wire in_76bar;
  wire in_75bar;
  wire in_74bar;
  wire in_73bar;
  wire in_72bar;
  wire in_71bar;
  wire in_70bar;
  wire in_69bar;
  wire in_68bar;
  wire in_67bar;
  wire in_66bar;
  wire in_65bar;
  wire in_64bar;
  wire in_63bar;
  wire in_62bar;
  wire in_61bar;
  wire in_60bar;
  wire in_59bar;
  wire in_58bar;
  wire in_57bar;
  wire in_56bar;
  wire in_55bar;
  wire in_54bar;
  wire in_53bar;
  wire in_52bar;
  wire in_51bar;
  wire in_50bar;
  wire in_49bar;
  wire in_48bar;
  wire in_47bar;
  wire in_46bar;
  wire in_45bar;
  wire in_44bar;
  wire in_43bar;
  wire in_42bar;
  wire in_41bar;
  wire in_40bar;
  wire in_39bar;
  wire in_38bar;
  wire in_37bar;
  wire in_36bar;
  wire in_35bar;
  wire in_34bar;
  wire in_33bar;
  wire in_32bar;
  wire in_31bar;
  wire in_30bar;
  wire in_29bar;
  wire in_28bar;
  wire in_27bar;
  wire in_26bar;
  wire in_25bar;
  wire in_24bar;
  wire in_23bar;
  wire in_22bar;
  wire in_21bar;
  wire in_20bar;
  wire in_19bar;
  wire in_18bar;
  wire in_17bar;
  wire in_16bar;
  wire in_15bar;
  wire in_14bar;
  wire in_13bar;
  wire in_12bar;
  wire in_11bar;
  wire in_10bar;
  wire in_9bar;
  wire in_8bar;
  wire in_7bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_3bar;
  wire in_2bar;
  wire in_1bar;
  wire in_0bar;
  wire n487bar;
  wire n488bar;
  wire n489bar;
  wire n490bar;
  wire n491bar;
  wire n492bar;
  wire n493bar;
  wire n494bar;
  wire n495bar;
  wire n496bar;
  wire n497bar;
  wire n498bar;
  wire n499bar;
  wire n500bar;
  wire n501bar;
  wire n502bar;
  wire n503bar;
  wire n504bar;
  wire n505bar;
  wire n506bar;
  wire n507bar;
  wire n508bar;
  wire n509bar;
  wire n510bar;
  wire n511bar;
  wire n512bar;
  wire n513bar;
  wire n514bar;
  wire n515bar;
  wire n516bar;
  wire n517bar;
  wire n518bar;
  wire n519bar;
  wire n520bar;
  wire n521bar;
  wire n522bar;
  wire n523bar;
  wire n524bar;
  wire n525bar;
  wire n526bar;
  wire n527bar;
  wire n528bar;
  wire n529bar;
  wire n530bar;
  wire n531bar;
  wire n532bar;
  wire n533bar;
  wire n534bar;
  wire n535bar;
  wire n536bar;
  wire n537bar;
  wire n538bar;
  wire n539bar;
  wire n540bar;
  wire n541bar;
  wire n542bar;
  wire n543bar;
  wire n544bar;
  wire n545bar;
  wire n546bar;
  wire n547bar;
  wire n548bar;
  wire n549bar;
  wire n550bar;
  wire n551bar;
  wire n552bar;
  wire n553bar;
  wire n554bar;
  wire n555bar;
  wire n556bar;
  wire n557bar;
  wire n558bar;
  wire n559bar;
  wire n560bar;
  wire n561bar;
  wire n562bar;
  wire n563bar;
  wire n564bar;
  wire n565bar;
  wire n566bar;
  wire n567bar;
  wire n568bar;
  wire n569bar;
  wire n570bar;
  wire n571bar;
  wire n572bar;
  wire n573bar;
  wire n574bar;
  wire n575bar;
  wire n576bar;
  wire n577bar;
  wire n578bar;
  wire n579bar;
  wire n580bar;
  wire n581bar;
  wire n582bar;
  wire n583bar;
  wire n584bar;
  wire n585bar;
  wire n586bar;
  wire n587bar;
  wire n588bar;
  wire n589bar;
  wire n590bar;
  wire n591bar;
  wire n592bar;
  wire n593bar;
  wire n594bar;
  wire n595bar;
  wire n596bar;
  wire n597bar;
  wire n598bar;
  wire n599bar;
  wire n600bar;
  wire n601bar;
  wire n602bar;
  wire n603bar;
  wire n604bar;
  wire n605bar;
  wire n606bar;
  wire n607bar;
  wire n608bar;
  wire n609bar;
  wire n610bar;
  wire n611bar;
  wire n612bar;
  wire n613bar;
  wire n614bar;
  wire n615bar;
  wire n616bar;
  wire n617bar;
  wire n618bar;
  wire n619bar;
  wire n620bar;
  wire n621bar;
  wire n622bar;
  wire n623bar;
  wire n624bar;
  wire n625bar;
  wire n626bar;
  wire n627bar;
  wire n628bar;
  wire n629bar;
  wire n630bar;
  wire n631bar;
  wire n632bar;
  wire n633bar;
  wire n634bar;
  wire n635bar;
  wire n636bar;
  wire n637bar;
  wire n638bar;
  wire n639bar;
  wire n640bar;
  wire n641bar;
  wire n642bar;
  wire n643bar;
  wire n644bar;
  wire n645bar;
  wire n646bar;
  wire n647bar;
  wire n648bar;
  wire n649bar;
  wire n650bar;
  wire n651bar;
  wire n652bar;
  wire n653bar;
  wire n654bar;
  wire n655bar;
  wire n656bar;
  wire n657bar;
  wire n658bar;
  wire n659bar;
  wire n660bar;
  wire n661bar;
  wire n662bar;
  wire n663bar;
  wire n664bar;
  wire n665bar;
  wire n666bar;
  wire n667bar;
  wire n668bar;
  wire n669bar;
  wire n670bar;
  wire n671bar;
  wire n672bar;
  wire n673bar;
  wire n674bar;
  wire n675bar;
  wire n676bar;
  wire n677bar;
  wire n678bar;
  wire n679bar;
  wire n680bar;
  wire n681bar;
  wire n682bar;
  wire n683bar;
  wire n684bar;
  wire n685bar;
  wire n686bar;
  wire n687bar;
  wire n688bar;
  wire n689bar;
  wire n690bar;
  wire n691bar;
  wire n692bar;
  wire n693bar;
  wire n694bar;
  wire n695bar;
  wire n696bar;
  wire n697bar;
  wire n698bar;
  wire n699bar;
  wire n700bar;
  wire n701bar;
  wire n702bar;
  wire n703bar;
  wire n704bar;
  wire n705bar;
  wire n706bar;
  wire n707bar;
  wire n708bar;
  wire n709bar;
  wire n710bar;
  wire n711bar;
  wire n712bar;
  wire n713bar;
  wire n714bar;
  wire n715bar;
  wire n716bar;
  wire n717bar;
  wire n718bar;
  wire n719bar;
  wire n720bar;
  wire n721bar;
  wire n722bar;
  wire n723bar;
  wire n724bar;
  wire n725bar;
  wire n726bar;
  wire n727bar;
  wire n728bar;
  wire n729bar;
  wire n730bar;
  wire n731bar;
  wire n732bar;
  wire n733bar;
  wire n734bar;
  wire n735bar;
  wire n736bar;
  wire n737bar;
  wire n738bar;
  wire n739bar;
  wire n740bar;
  wire n741bar;
  wire n742bar;
  wire n743bar;
  wire n744bar;
  wire n745bar;
  wire n746bar;
  wire n747bar;
  wire n748bar;
  wire n749bar;
  wire n750bar;
  wire n751bar;
  wire n752bar;
  wire n753bar;
  wire n754bar;
  wire n755bar;
  wire n756bar;
  wire n757bar;
  wire n758bar;
  wire n759bar;
  wire n760bar;
  wire n761bar;
  wire n762bar;
  wire n763bar;
  wire n764bar;
  wire n765bar;
  wire n766bar;
  wire n767bar;
  wire n768bar;
  wire n769bar;
  wire n770bar;
  wire n771bar;
  wire n772bar;
  wire n773bar;
  wire n774bar;
  wire n775bar;
  wire n776bar;
  wire n777bar;
  wire n778bar;
  wire n779bar;
  wire n780bar;
  wire n781bar;
  wire n782bar;
  wire n783bar;
  wire n784bar;
  wire n785bar;
  wire n786bar;
  wire n787bar;
  wire n788bar;
  wire n789bar;
  wire n790bar;
  wire n791bar;
  wire n792bar;
  wire n793bar;
  wire n794bar;
  wire n795bar;
  wire n796bar;
  wire n797bar;
  wire n798bar;
  wire n799bar;
  wire n800bar;
  wire n801bar;
  wire n802bar;
  wire n803bar;
  wire n804bar;
  wire n805bar;
  wire n806bar;
  wire n807bar;
  wire n808bar;
  wire n809bar;
  wire n810bar;
  wire n811bar;
  wire n812bar;
  wire n813bar;
  wire n814bar;
  wire n815bar;
  wire n816bar;
  wire n817bar;
  wire n818bar;
  wire n819bar;
  wire n820bar;
  wire n821bar;
  wire n822bar;
  wire n823bar;
  wire n824bar;
  wire n825bar;
  wire n826bar;
  wire n827bar;
  wire n828bar;
  wire n829bar;
  wire n830bar;
  wire n831bar;
  wire n832bar;
  wire n833bar;
  wire n834bar;
  wire n835bar;
  wire n836bar;
  wire n837bar;
  wire n838bar;
  wire n839bar;
  wire n840bar;
  wire n841bar;
  wire n842bar;
  wire n843bar;
  wire n844bar;
  wire n845bar;
  wire n846bar;
  wire n847bar;
  wire n848bar;
  wire n849bar;
  wire n850bar;
  wire n851bar;
  wire n852bar;
  wire n853bar;
  wire n854bar;
  wire n855bar;
  wire n856bar;
  wire n857bar;
  wire n858bar;
  wire n859bar;
  wire n860bar;
  wire n861bar;
  wire n862bar;
  wire n863bar;
  wire n864bar;
  wire n865bar;
  wire n866bar;
  wire n867bar;
  wire n868bar;
  wire n869bar;
  wire n870bar;
  wire n871bar;
  wire n872bar;
  wire n873bar;
  wire n874bar;
  wire n875bar;
  wire n876bar;
  wire n877bar;
  wire n878bar;
  wire n879bar;
  wire n880bar;
  wire n881bar;
  wire n882bar;
  wire n883bar;
  wire n884bar;
  wire n885bar;
  wire n886bar;
  wire n887bar;
  wire n888bar;
  wire n889bar;
  wire n890bar;
  wire n891bar;
  wire n892bar;
  wire n893bar;
  wire n894bar;
  wire n895bar;
  wire n896bar;
  wire n897bar;
  wire n898bar;
  wire n899bar;
  wire n900bar;
  wire n901bar;
  wire n902bar;
  wire n903bar;
  wire n904bar;
  wire n905bar;
  wire n906bar;
  wire n907bar;
  wire n908bar;
  wire n909bar;
  wire n910bar;
  wire n911bar;
  wire n912bar;
  wire n913bar;
  wire n914bar;
  wire n915bar;
  wire n916bar;
  wire n917bar;
  wire n918bar;
  wire n919bar;
  wire n920bar;
  wire n921bar;
  wire n922bar;
  wire n923bar;
  wire n924bar;
  wire n925bar;
  wire n926bar;
  wire n927bar;
  wire n928bar;
  wire n929bar;
  wire n930bar;
  wire n931bar;
  wire n932bar;
  wire n933bar;
  wire n934bar;
  wire n935bar;
  wire n936bar;
  wire n937bar;
  wire n938bar;
  wire n939bar;
  wire n940bar;
  wire n941bar;
  wire n942bar;
  wire n943bar;
  wire n944bar;
  wire n945bar;
  wire n946bar;
  wire n947bar;
  wire n948bar;
  wire n949bar;
  wire n950bar;
  wire n951bar;
  wire n952bar;
  wire n953bar;
  wire n954bar;
  wire n955bar;
  wire n956bar;
  wire n957bar;
  wire n958bar;
  wire n959bar;
  wire n960bar;
  wire n961bar;
  wire n962bar;
  wire n963bar;
  wire n964bar;
  wire n965bar;
  wire n966bar;
  wire n967bar;
  wire n968bar;
  wire n969bar;
  wire n970bar;
  wire n971bar;
  wire n972bar;
//wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];
  assign in_81bar = inbar[81];
  assign in_80bar = inbar[80];
  assign in_79bar = inbar[79];
  assign in_78bar = inbar[78];
  assign in_77bar = inbar[77];
  assign in_76bar = inbar[76];
  assign in_75bar = inbar[75];
  assign in_74bar = inbar[74];
  assign in_73bar = inbar[73];
  assign in_72bar = inbar[72];
  assign in_71bar = inbar[71];
  assign in_70bar = inbar[70];
  assign in_69bar = inbar[69];
  assign in_68bar = inbar[68];
  assign in_67bar = inbar[67];
  assign in_66bar = inbar[66];
  assign in_65bar = inbar[65];
  assign in_64bar = inbar[64];
  assign in_63bar = inbar[63];
  assign in_62bar = inbar[62];
  assign in_61bar = inbar[61];
  assign in_60bar = inbar[60];
  assign in_59bar = inbar[59];
  assign in_58bar = inbar[58];
  assign in_57bar = inbar[57];
  assign in_56bar = inbar[56];
  assign in_55bar = inbar[55];
  assign in_54bar = inbar[54];
  assign in_53bar = inbar[53];
  assign in_52bar = inbar[52];
  assign in_51bar = inbar[51];
  assign in_50bar = inbar[50];
  assign in_49bar = inbar[49];
  assign in_48bar = inbar[48];
  assign in_47bar = inbar[47];
  assign in_46bar = inbar[46];
  assign in_45bar = inbar[45];
  assign in_44bar = inbar[44];
  assign in_43bar = inbar[43];
  assign in_42bar = inbar[42];
  assign in_41bar = inbar[41];
  assign in_40bar = inbar[40];
  assign in_39bar = inbar[39];
  assign in_38bar = inbar[38];
  assign in_37bar = inbar[37];
  assign in_36bar = inbar[36];
  assign in_35bar = inbar[35];
  assign in_34bar = inbar[34];
  assign in_33bar = inbar[33];
  assign in_32bar = inbar[32];
  assign in_31bar = inbar[31];
  assign in_30bar = inbar[30];
  assign in_29bar = inbar[29];
  assign in_28bar = inbar[28];
  assign in_27bar = inbar[27];
  assign in_26bar = inbar[26];
  assign in_25bar = inbar[25];
  assign in_24bar = inbar[24];
  assign in_23bar = inbar[23];
  assign in_22bar = inbar[22];
  assign in_21bar = inbar[21];
  assign in_20bar = inbar[20];
  assign in_19bar = inbar[19];
  assign in_18bar = inbar[18];
  assign in_17bar = inbar[17];
  assign in_16bar = inbar[16];
  assign in_15bar = inbar[15];
  assign in_14bar = inbar[14];
  assign in_13bar = inbar[13];
  assign in_12bar = inbar[12];
  assign in_11bar = inbar[11];
  assign in_10bar = inbar[10];
  assign in_9bar = inbar[9];
  assign in_8bar = inbar[8];
  assign in_7bar = inbar[7];
  assign in_6bar = inbar[6];
  assign in_5bar = inbar[5];
  assign in_4bar = inbar[4];
  assign in_3bar = inbar[3];
  assign in_2bar = inbar[2];
  assign in_1bar = inbar[1];
  assign in_0bar = inbar[0];
//assign_done

  OR2_X1 U1 ( .A1(n972), .A2(n971), .ZN(out[7]) );
  AND2_X1 U1bar ( .A1(n972bar), .A2(n971bar), .ZN(outbar[7]) );
  OR2_X1 U2 ( .A1(n970), .A2(n969), .ZN(n971) );
  AND2_X1 U2bar ( .A1(n970bar), .A2(n969bar), .ZN(n971bar) );
  OR2_X1 U3 ( .A1(n968), .A2(n967), .ZN(n969) );
  AND2_X1 U3bar ( .A1(n968bar), .A2(n967bar), .ZN(n969bar) );
  OR2_X1 U4 ( .A1(n966), .A2(n965), .ZN(n967) );
  AND2_X1 U4bar ( .A1(n966bar), .A2(n965bar), .ZN(n967bar) );
  OR2_X1 U5 ( .A1(n964), .A2(n963), .ZN(n968) );
  AND2_X1 U5bar ( .A1(n964bar), .A2(n963bar), .ZN(n968bar) );
  OR2_X1 U6 ( .A1(in[116]), .A2(n962), .ZN(n963) );
  AND2_X1 U6bar ( .A1(inbar[116]), .A2(n962bar), .ZN(n963bar) );
  OR2_X1 U7 ( .A1(n961), .A2(n960), .ZN(n970) );
  AND2_X1 U7bar ( .A1(n961bar), .A2(n960bar), .ZN(n970bar) );
  OR2_X1 U8 ( .A1(in[150]), .A2(in[127]), .ZN(n960) );
  AND2_X1 U8bar ( .A1(inbar[150]), .A2(inbar[127]), .ZN(n960bar) );
  OR2_X1 U9 ( .A1(in[160]), .A2(n959), .ZN(n961) );
  AND2_X1 U9bar ( .A1(inbar[160]), .A2(n959bar), .ZN(n961bar) );
  OR2_X1 U10 ( .A1(in[252]), .A2(in[168]), .ZN(n959) );
  AND2_X1 U10bar ( .A1(inbar[252]), .A2(inbar[168]), .ZN(n959bar) );
  OR2_X1 U11 ( .A1(n958), .A2(n957), .ZN(n972) );
  AND2_X1 U11bar ( .A1(n958bar), .A2(n957bar), .ZN(n972bar) );
  OR2_X1 U12 ( .A1(n956), .A2(n955), .ZN(n957) );
  AND2_X1 U12bar ( .A1(n956bar), .A2(n955bar), .ZN(n957bar) );
  OR2_X1 U13 ( .A1(in_17), .A2(in[96]), .ZN(n955) );
  AND2_X1 U13bar ( .A1(in_17bar), .A2(inbar[96]), .ZN(n955bar) );
  OR2_X1 U14 ( .A1(in_23), .A2(n954), .ZN(n956) );
  AND2_X1 U14bar ( .A1(in_23bar), .A2(n954bar), .ZN(n956bar) );
  OR2_X1 U15 ( .A1(in_31), .A2(in_26), .ZN(n954) );
  AND2_X1 U15bar ( .A1(in_31bar), .A2(in_26bar), .ZN(n954bar) );
  OR2_X1 U16 ( .A1(n953), .A2(n952), .ZN(n958) );
  AND2_X1 U16bar ( .A1(n953bar), .A2(n952bar), .ZN(n958bar) );
  OR2_X1 U17 ( .A1(in_58), .A2(in_4), .ZN(n952) );
  AND2_X1 U17bar ( .A1(in_58bar), .A2(in_4bar), .ZN(n952bar) );
  OR2_X1 U18 ( .A1(in_59), .A2(n951), .ZN(n953) );
  AND2_X1 U18bar ( .A1(in_59bar), .A2(n951bar), .ZN(n953bar) );
  OR2_X1 U19 ( .A1(in_71), .A2(in_62), .ZN(n951) );
  AND2_X1 U19bar ( .A1(in_71bar), .A2(in_62bar), .ZN(n951bar) );
  OR2_X1 U20 ( .A1(n950), .A2(n949), .ZN(out[6]) );
  AND2_X1 U20bar ( .A1(n950bar), .A2(n949bar), .ZN(outbar[6]) );
  OR2_X1 U21 ( .A1(n948), .A2(n947), .ZN(n949) );
  AND2_X1 U21bar ( .A1(n948bar), .A2(n947bar), .ZN(n949bar) );
  OR2_X1 U22 ( .A1(n946), .A2(n945), .ZN(n947) );
  AND2_X1 U22bar ( .A1(n946bar), .A2(n945bar), .ZN(n947bar) );
  OR2_X1 U23 ( .A1(n944), .A2(n943), .ZN(n945) );
  AND2_X1 U23bar ( .A1(n944bar), .A2(n943bar), .ZN(n945bar) );
  OR2_X1 U24 ( .A1(n942), .A2(n941), .ZN(n946) );
  AND2_X1 U24bar ( .A1(n942bar), .A2(n941bar), .ZN(n946bar) );
  OR2_X1 U25 ( .A1(in[101]), .A2(n940), .ZN(n941) );
  AND2_X1 U25bar ( .A1(inbar[101]), .A2(n940bar), .ZN(n941bar) );
  OR2_X1 U26 ( .A1(n939), .A2(n938), .ZN(n948) );
  AND2_X1 U26bar ( .A1(n939bar), .A2(n938bar), .ZN(n948bar) );
  OR2_X1 U27 ( .A1(in[114]), .A2(in[104]), .ZN(n938) );
  AND2_X1 U27bar ( .A1(inbar[114]), .A2(inbar[104]), .ZN(n938bar) );
  OR2_X1 U28 ( .A1(in[128]), .A2(n937), .ZN(n939) );
  AND2_X1 U28bar ( .A1(inbar[128]), .A2(n937bar), .ZN(n939bar) );
  OR2_X1 U29 ( .A1(in[136]), .A2(in[134]), .ZN(n937) );
  AND2_X1 U29bar ( .A1(inbar[136]), .A2(inbar[134]), .ZN(n937bar) );
  OR2_X1 U30 ( .A1(n936), .A2(n935), .ZN(n950) );
  AND2_X1 U30bar ( .A1(n936bar), .A2(n935bar), .ZN(n950bar) );
  OR2_X1 U31 ( .A1(n934), .A2(n933), .ZN(n935) );
  AND2_X1 U31bar ( .A1(n934bar), .A2(n933bar), .ZN(n935bar) );
  OR2_X1 U32 ( .A1(in[177]), .A2(in[164]), .ZN(n933) );
  AND2_X1 U32bar ( .A1(inbar[177]), .A2(inbar[164]), .ZN(n933bar) );
  OR2_X1 U33 ( .A1(in[212]), .A2(n932), .ZN(n934) );
  AND2_X1 U33bar ( .A1(inbar[212]), .A2(n932bar), .ZN(n934bar) );
  OR2_X1 U34 ( .A1(in[248]), .A2(in[221]), .ZN(n932) );
  AND2_X1 U34bar ( .A1(inbar[248]), .A2(inbar[221]), .ZN(n932bar) );
  OR2_X1 U35 ( .A1(n931), .A2(n930), .ZN(n936) );
  AND2_X1 U35bar ( .A1(n931bar), .A2(n930bar), .ZN(n936bar) );
  OR2_X1 U36 ( .A1(in_18), .A2(in[93]), .ZN(n930) );
  AND2_X1 U36bar ( .A1(in_18bar), .A2(inbar[93]), .ZN(n930bar) );
  OR2_X1 U37 ( .A1(in_31), .A2(n929), .ZN(n931) );
  AND2_X1 U37bar ( .A1(in_31bar), .A2(n929bar), .ZN(n931bar) );
  OR2_X1 U38 ( .A1(in_7), .A2(in_39), .ZN(n929) );
  AND2_X1 U38bar ( .A1(in_7bar), .A2(in_39bar), .ZN(n929bar) );
  OR2_X1 U39 ( .A1(n928), .A2(n927), .ZN(out[5]) );
  AND2_X1 U39bar ( .A1(n928bar), .A2(n927bar), .ZN(outbar[5]) );
  OR2_X1 U40 ( .A1(n926), .A2(n925), .ZN(n927) );
  AND2_X1 U40bar ( .A1(n926bar), .A2(n925bar), .ZN(n927bar) );
  OR2_X1 U41 ( .A1(n924), .A2(n923), .ZN(n925) );
  AND2_X1 U41bar ( .A1(n924bar), .A2(n923bar), .ZN(n925bar) );
  OR2_X1 U42 ( .A1(n922), .A2(n921), .ZN(n923) );
  AND2_X1 U42bar ( .A1(n922bar), .A2(n921bar), .ZN(n923bar) );
  OR2_X1 U43 ( .A1(n940), .A2(n920), .ZN(n924) );
  AND2_X1 U43bar ( .A1(n940bar), .A2(n920bar), .ZN(n924bar) );
  OR2_X1 U44 ( .A1(in[111]), .A2(n919), .ZN(n920) );
  AND2_X1 U44bar ( .A1(inbar[111]), .A2(n919bar), .ZN(n920bar) );
  OR2_X1 U45 ( .A1(n918), .A2(n917), .ZN(n940) );
  AND2_X1 U45bar ( .A1(n918bar), .A2(n917bar), .ZN(n940bar) );
  OR2_X1 U46 ( .A1(n916), .A2(n915), .ZN(n917) );
  AND2_X1 U46bar ( .A1(n916bar), .A2(n915bar), .ZN(n917bar) );
  OR2_X1 U47 ( .A1(n914), .A2(n913), .ZN(n915) );
  AND2_X1 U47bar ( .A1(n914bar), .A2(n913bar), .ZN(n915bar) );
  OR2_X1 U48 ( .A1(in[140]), .A2(in[131]), .ZN(n913) );
  AND2_X1 U48bar ( .A1(inbar[140]), .A2(inbar[131]), .ZN(n913bar) );
  OR2_X1 U49 ( .A1(in[160]), .A2(in[144]), .ZN(n914) );
  AND2_X1 U49bar ( .A1(inbar[160]), .A2(inbar[144]), .ZN(n914bar) );
  OR2_X1 U50 ( .A1(n912), .A2(n911), .ZN(n916) );
  AND2_X1 U50bar ( .A1(n912bar), .A2(n911bar), .ZN(n916bar) );
  OR2_X1 U51 ( .A1(in[179]), .A2(in[174]), .ZN(n911) );
  AND2_X1 U51bar ( .A1(inbar[179]), .A2(inbar[174]), .ZN(n911bar) );
  OR2_X1 U52 ( .A1(in[188]), .A2(in[184]), .ZN(n912) );
  AND2_X1 U52bar ( .A1(inbar[188]), .A2(inbar[184]), .ZN(n912bar) );
  OR2_X1 U53 ( .A1(n910), .A2(n909), .ZN(n918) );
  AND2_X1 U53bar ( .A1(n910bar), .A2(n909bar), .ZN(n918bar) );
  OR2_X1 U54 ( .A1(n908), .A2(n907), .ZN(n909) );
  AND2_X1 U54bar ( .A1(n908bar), .A2(n907bar), .ZN(n909bar) );
  OR2_X1 U55 ( .A1(in[216]), .A2(in[200]), .ZN(n907) );
  AND2_X1 U55bar ( .A1(inbar[216]), .A2(inbar[200]), .ZN(n907bar) );
  OR2_X1 U56 ( .A1(in[228]), .A2(in[224]), .ZN(n908) );
  AND2_X1 U56bar ( .A1(inbar[228]), .A2(inbar[224]), .ZN(n908bar) );
  OR2_X1 U57 ( .A1(n906), .A2(n905), .ZN(n910) );
  AND2_X1 U57bar ( .A1(n906bar), .A2(n905bar), .ZN(n910bar) );
  OR2_X1 U58 ( .A1(in[247]), .A2(in[235]), .ZN(n905) );
  AND2_X1 U58bar ( .A1(inbar[247]), .A2(inbar[235]), .ZN(n905bar) );
  OR2_X1 U59 ( .A1(in_42), .A2(in[83]), .ZN(n906) );
  AND2_X1 U59bar ( .A1(in_42bar), .A2(inbar[83]), .ZN(n906bar) );
  OR2_X1 U60 ( .A1(n904), .A2(n903), .ZN(n926) );
  AND2_X1 U60bar ( .A1(n904bar), .A2(n903bar), .ZN(n926bar) );
  OR2_X1 U61 ( .A1(in[166]), .A2(in[123]), .ZN(n903) );
  AND2_X1 U61bar ( .A1(inbar[166]), .A2(inbar[123]), .ZN(n903bar) );
  OR2_X1 U62 ( .A1(in[170]), .A2(n902), .ZN(n904) );
  AND2_X1 U62bar ( .A1(inbar[170]), .A2(n902bar), .ZN(n904bar) );
  OR2_X1 U63 ( .A1(in[194]), .A2(in[183]), .ZN(n902) );
  AND2_X1 U63bar ( .A1(inbar[194]), .A2(inbar[183]), .ZN(n902bar) );
  OR2_X1 U64 ( .A1(n901), .A2(n900), .ZN(n928) );
  AND2_X1 U64bar ( .A1(n901bar), .A2(n900bar), .ZN(n928bar) );
  OR2_X1 U65 ( .A1(n899), .A2(n898), .ZN(n900) );
  AND2_X1 U65bar ( .A1(n899bar), .A2(n898bar), .ZN(n900bar) );
  OR2_X1 U66 ( .A1(in[241]), .A2(in[238]), .ZN(n898) );
  AND2_X1 U66bar ( .A1(inbar[241]), .A2(inbar[238]), .ZN(n898bar) );
  OR2_X1 U67 ( .A1(in[250]), .A2(n897), .ZN(n899) );
  AND2_X1 U67bar ( .A1(inbar[250]), .A2(n897bar), .ZN(n899bar) );
  OR2_X1 U68 ( .A1(in_24), .A2(in[84]), .ZN(n897) );
  AND2_X1 U68bar ( .A1(in_24bar), .A2(inbar[84]), .ZN(n897bar) );
  OR2_X1 U69 ( .A1(n896), .A2(n895), .ZN(n901) );
  AND2_X1 U69bar ( .A1(n896bar), .A2(n895bar), .ZN(n901bar) );
  OR2_X1 U70 ( .A1(in_41), .A2(in_29), .ZN(n895) );
  AND2_X1 U70bar ( .A1(in_41bar), .A2(in_29bar), .ZN(n895bar) );
  OR2_X1 U71 ( .A1(in_66), .A2(n894), .ZN(n896) );
  AND2_X1 U71bar ( .A1(in_66bar), .A2(n894bar), .ZN(n896bar) );
  OR2_X1 U72 ( .A1(in_76), .A2(in_71), .ZN(n894) );
  AND2_X1 U72bar ( .A1(in_76bar), .A2(in_71bar), .ZN(n894bar) );
  OR2_X1 U73 ( .A1(n893), .A2(n892), .ZN(out[4]) );
  AND2_X1 U73bar ( .A1(n893bar), .A2(n892bar), .ZN(outbar[4]) );
  OR2_X1 U74 ( .A1(n891), .A2(n890), .ZN(n892) );
  AND2_X1 U74bar ( .A1(n891bar), .A2(n890bar), .ZN(n892bar) );
  OR2_X1 U75 ( .A1(n889), .A2(n888), .ZN(n890) );
  AND2_X1 U75bar ( .A1(n889bar), .A2(n888bar), .ZN(n890bar) );
  OR2_X1 U76 ( .A1(n922), .A2(n887), .ZN(n888) );
  AND2_X1 U76bar ( .A1(n922bar), .A2(n887bar), .ZN(n888bar) );
  OR2_X1 U77 ( .A1(n886), .A2(n885), .ZN(n922) );
  AND2_X1 U77bar ( .A1(n886bar), .A2(n885bar), .ZN(n922bar) );
  OR2_X1 U78 ( .A1(n884), .A2(n883), .ZN(n885) );
  AND2_X1 U78bar ( .A1(n884bar), .A2(n883bar), .ZN(n885bar) );
  OR2_X1 U79 ( .A1(n882), .A2(n881), .ZN(n883) );
  AND2_X1 U79bar ( .A1(n882bar), .A2(n881bar), .ZN(n883bar) );
  OR2_X1 U80 ( .A1(in[118]), .A2(in[109]), .ZN(n881) );
  AND2_X1 U80bar ( .A1(inbar[118]), .A2(inbar[109]), .ZN(n881bar) );
  OR2_X1 U81 ( .A1(in[139]), .A2(in[120]), .ZN(n882) );
  AND2_X1 U81bar ( .A1(inbar[139]), .A2(inbar[120]), .ZN(n882bar) );
  OR2_X1 U82 ( .A1(n880), .A2(n879), .ZN(n884) );
  AND2_X1 U82bar ( .A1(n880bar), .A2(n879bar), .ZN(n884bar) );
  OR2_X1 U83 ( .A1(in[198]), .A2(in[154]), .ZN(n879) );
  AND2_X1 U83bar ( .A1(inbar[198]), .A2(inbar[154]), .ZN(n879bar) );
  OR2_X1 U84 ( .A1(in[210]), .A2(in[205]), .ZN(n880) );
  AND2_X1 U84bar ( .A1(inbar[210]), .A2(inbar[205]), .ZN(n880bar) );
  OR2_X1 U85 ( .A1(n878), .A2(n877), .ZN(n886) );
  AND2_X1 U85bar ( .A1(n878bar), .A2(n877bar), .ZN(n886bar) );
  OR2_X1 U86 ( .A1(n876), .A2(n875), .ZN(n877) );
  AND2_X1 U86bar ( .A1(n876bar), .A2(n875bar), .ZN(n877bar) );
  OR2_X1 U87 ( .A1(in[219]), .A2(in[217]), .ZN(n875) );
  AND2_X1 U87bar ( .A1(inbar[219]), .A2(inbar[217]), .ZN(n875bar) );
  OR2_X1 U88 ( .A1(in[86]), .A2(in[252]), .ZN(n876) );
  AND2_X1 U88bar ( .A1(inbar[86]), .A2(inbar[252]), .ZN(n876bar) );
  OR2_X1 U89 ( .A1(n874), .A2(n873), .ZN(n878) );
  AND2_X1 U89bar ( .A1(n874bar), .A2(n873bar), .ZN(n878bar) );
  OR2_X1 U90 ( .A1(in_40), .A2(in[91]), .ZN(n873) );
  AND2_X1 U90bar ( .A1(in_40bar), .A2(inbar[91]), .ZN(n873bar) );
  OR2_X1 U91 ( .A1(in_8), .A2(in_46), .ZN(n874) );
  AND2_X1 U91bar ( .A1(in_8bar), .A2(in_46bar), .ZN(n874bar) );
  OR2_X1 U92 ( .A1(n872), .A2(n871), .ZN(n889) );
  AND2_X1 U92bar ( .A1(n872bar), .A2(n871bar), .ZN(n889bar) );
  OR2_X1 U93 ( .A1(in[117]), .A2(n943), .ZN(n871) );
  AND2_X1 U93bar ( .A1(inbar[117]), .A2(n943bar), .ZN(n871bar) );
  OR2_X1 U94 ( .A1(n870), .A2(n869), .ZN(n943) );
  AND2_X1 U94bar ( .A1(n870bar), .A2(n869bar), .ZN(n943bar) );
  OR2_X1 U95 ( .A1(n868), .A2(n867), .ZN(n869) );
  AND2_X1 U95bar ( .A1(n868bar), .A2(n867bar), .ZN(n869bar) );
  OR2_X1 U96 ( .A1(n866), .A2(n865), .ZN(n867) );
  AND2_X1 U96bar ( .A1(n866bar), .A2(n865bar), .ZN(n867bar) );
  OR2_X1 U97 ( .A1(n864), .A2(n863), .ZN(n865) );
  AND2_X1 U97bar ( .A1(n864bar), .A2(n863bar), .ZN(n865bar) );
  OR2_X1 U98 ( .A1(in[108]), .A2(n919), .ZN(n866) );
  AND2_X1 U98bar ( .A1(inbar[108]), .A2(n919bar), .ZN(n866bar) );
  OR2_X1 U99 ( .A1(n862), .A2(n861), .ZN(n919) );
  AND2_X1 U99bar ( .A1(n862bar), .A2(n861bar), .ZN(n919bar) );
  OR2_X1 U100 ( .A1(n860), .A2(n859), .ZN(n861) );
  AND2_X1 U100bar ( .A1(n860bar), .A2(n859bar), .ZN(n861bar) );
  OR2_X1 U101 ( .A1(n858), .A2(n857), .ZN(n859) );
  AND2_X1 U101bar ( .A1(n858bar), .A2(n857bar), .ZN(n859bar) );
  OR2_X1 U102 ( .A1(in[119]), .A2(in[105]), .ZN(n857) );
  AND2_X1 U102bar ( .A1(inbar[119]), .A2(inbar[105]), .ZN(n857bar) );
  OR2_X1 U103 ( .A1(in[186]), .A2(in[175]), .ZN(n858) );
  AND2_X1 U103bar ( .A1(inbar[186]), .A2(inbar[175]), .ZN(n858bar) );
  OR2_X1 U104 ( .A1(n856), .A2(n855), .ZN(n860) );
  AND2_X1 U104bar ( .A1(n856bar), .A2(n855bar), .ZN(n860bar) );
  OR2_X1 U105 ( .A1(in[202]), .A2(in[193]), .ZN(n855) );
  AND2_X1 U105bar ( .A1(inbar[202]), .A2(inbar[193]), .ZN(n855bar) );
  OR2_X1 U106 ( .A1(in[225]), .A2(in[208]), .ZN(n856) );
  AND2_X1 U106bar ( .A1(inbar[225]), .A2(inbar[208]), .ZN(n856bar) );
  OR2_X1 U107 ( .A1(n854), .A2(n853), .ZN(n862) );
  AND2_X1 U107bar ( .A1(n854bar), .A2(n853bar), .ZN(n862bar) );
  OR2_X1 U108 ( .A1(n852), .A2(n851), .ZN(n853) );
  AND2_X1 U108bar ( .A1(n852bar), .A2(n851bar), .ZN(n853bar) );
  OR2_X1 U109 ( .A1(in_1), .A2(in[85]), .ZN(n851) );
  AND2_X1 U109bar ( .A1(in_1bar), .A2(inbar[85]), .ZN(n851bar) );
  OR2_X1 U110 ( .A1(in_23), .A2(in_19), .ZN(n852) );
  AND2_X1 U110bar ( .A1(in_23bar), .A2(in_19bar), .ZN(n852bar) );
  OR2_X1 U111 ( .A1(n850), .A2(n849), .ZN(n854) );
  AND2_X1 U111bar ( .A1(n850bar), .A2(n849bar), .ZN(n854bar) );
  OR2_X1 U112 ( .A1(in_43), .A2(in_33), .ZN(n849) );
  AND2_X1 U112bar ( .A1(in_43bar), .A2(in_33bar), .ZN(n849bar) );
  OR2_X1 U113 ( .A1(in_63), .A2(in_44), .ZN(n850) );
  AND2_X1 U113bar ( .A1(in_63bar), .A2(in_44bar), .ZN(n850bar) );
  OR2_X1 U114 ( .A1(n848), .A2(n847), .ZN(n868) );
  AND2_X1 U114bar ( .A1(n848bar), .A2(n847bar), .ZN(n868bar) );
  OR2_X1 U115 ( .A1(in[141]), .A2(in[112]), .ZN(n847) );
  AND2_X1 U115bar ( .A1(inbar[141]), .A2(inbar[112]), .ZN(n847bar) );
  OR2_X1 U116 ( .A1(in[147]), .A2(n846), .ZN(n848) );
  AND2_X1 U116bar ( .A1(inbar[147]), .A2(n846bar), .ZN(n848bar) );
  OR2_X1 U117 ( .A1(in[181]), .A2(in[167]), .ZN(n846) );
  AND2_X1 U117bar ( .A1(inbar[181]), .A2(inbar[167]), .ZN(n846bar) );
  OR2_X1 U118 ( .A1(n845), .A2(n844), .ZN(n870) );
  AND2_X1 U118bar ( .A1(n845bar), .A2(n844bar), .ZN(n870bar) );
  OR2_X1 U119 ( .A1(n843), .A2(n842), .ZN(n844) );
  AND2_X1 U119bar ( .A1(n843bar), .A2(n842bar), .ZN(n844bar) );
  OR2_X1 U120 ( .A1(in[229]), .A2(in[201]), .ZN(n842) );
  AND2_X1 U120bar ( .A1(inbar[229]), .A2(inbar[201]), .ZN(n842bar) );
  OR2_X1 U121 ( .A1(in[237]), .A2(n841), .ZN(n843) );
  AND2_X1 U121bar ( .A1(inbar[237]), .A2(n841bar), .ZN(n843bar) );
  OR2_X1 U122 ( .A1(in[94]), .A2(in[253]), .ZN(n841) );
  AND2_X1 U122bar ( .A1(inbar[94]), .A2(inbar[253]), .ZN(n841bar) );
  OR2_X1 U123 ( .A1(n840), .A2(n839), .ZN(n845) );
  AND2_X1 U123bar ( .A1(n840bar), .A2(n839bar), .ZN(n845bar) );
  OR2_X1 U124 ( .A1(in_21), .A2(in[96]), .ZN(n839) );
  AND2_X1 U124bar ( .A1(in_21bar), .A2(inbar[96]), .ZN(n839bar) );
  OR2_X1 U125 ( .A1(in_25), .A2(n838), .ZN(n840) );
  AND2_X1 U125bar ( .A1(in_25bar), .A2(n838bar), .ZN(n840bar) );
  OR2_X1 U126 ( .A1(in_81), .A2(in_45), .ZN(n838) );
  AND2_X1 U126bar ( .A1(in_81bar), .A2(in_45bar), .ZN(n838bar) );
  OR2_X1 U127 ( .A1(n837), .A2(n836), .ZN(n891) );
  AND2_X1 U127bar ( .A1(n837bar), .A2(n836bar), .ZN(n891bar) );
  OR2_X1 U128 ( .A1(in[142]), .A2(in[124]), .ZN(n836) );
  AND2_X1 U128bar ( .A1(inbar[142]), .A2(inbar[124]), .ZN(n836bar) );
  OR2_X1 U129 ( .A1(in[150]), .A2(n835), .ZN(n837) );
  AND2_X1 U129bar ( .A1(inbar[150]), .A2(n835bar), .ZN(n837bar) );
  OR2_X1 U130 ( .A1(in[172]), .A2(in[155]), .ZN(n835) );
  AND2_X1 U130bar ( .A1(inbar[172]), .A2(inbar[155]), .ZN(n835bar) );
  OR2_X1 U131 ( .A1(n834), .A2(n833), .ZN(n893) );
  AND2_X1 U131bar ( .A1(n834bar), .A2(n833bar), .ZN(n893bar) );
  OR2_X1 U132 ( .A1(n832), .A2(n831), .ZN(n833) );
  AND2_X1 U132bar ( .A1(n832bar), .A2(n831bar), .ZN(n833bar) );
  OR2_X1 U133 ( .A1(in[196]), .A2(in[173]), .ZN(n831) );
  AND2_X1 U133bar ( .A1(inbar[196]), .A2(inbar[173]), .ZN(n831bar) );
  OR2_X1 U134 ( .A1(in[222]), .A2(n830), .ZN(n832) );
  AND2_X1 U134bar ( .A1(inbar[222]), .A2(n830bar), .ZN(n832bar) );
  OR2_X1 U135 ( .A1(in[227]), .A2(in[226]), .ZN(n830) );
  AND2_X1 U135bar ( .A1(inbar[227]), .A2(inbar[226]), .ZN(n830bar) );
  OR2_X1 U136 ( .A1(n829), .A2(n828), .ZN(n834) );
  AND2_X1 U136bar ( .A1(n829bar), .A2(n828bar), .ZN(n834bar) );
  OR2_X1 U137 ( .A1(in[249]), .A2(in[231]), .ZN(n828) );
  AND2_X1 U137bar ( .A1(inbar[249]), .A2(inbar[231]), .ZN(n828bar) );
  OR2_X1 U138 ( .A1(in_28), .A2(n827), .ZN(n829) );
  AND2_X1 U138bar ( .A1(in_28bar), .A2(n827bar), .ZN(n829bar) );
  OR2_X1 U139 ( .A1(in_52), .A2(in_47), .ZN(n827) );
  AND2_X1 U139bar ( .A1(in_52bar), .A2(in_47bar), .ZN(n827bar) );
  OR2_X1 U140 ( .A1(n826), .A2(n825), .ZN(out[3]) );
  AND2_X1 U140bar ( .A1(n826bar), .A2(n825bar), .ZN(outbar[3]) );
  OR2_X1 U141 ( .A1(n824), .A2(n823), .ZN(n825) );
  AND2_X1 U141bar ( .A1(n824bar), .A2(n823bar), .ZN(n825bar) );
  OR2_X1 U142 ( .A1(n822), .A2(n821), .ZN(n823) );
  AND2_X1 U142bar ( .A1(n822bar), .A2(n821bar), .ZN(n823bar) );
  OR2_X1 U143 ( .A1(n820), .A2(n819), .ZN(n821) );
  AND2_X1 U143bar ( .A1(n820bar), .A2(n819bar), .ZN(n821bar) );
  OR2_X1 U144 ( .A1(n964), .A2(n818), .ZN(n822) );
  AND2_X1 U144bar ( .A1(n964bar), .A2(n818bar), .ZN(n822bar) );
  OR2_X1 U145 ( .A1(in[118]), .A2(n817), .ZN(n818) );
  AND2_X1 U145bar ( .A1(inbar[118]), .A2(n817bar), .ZN(n818bar) );
  OR2_X1 U146 ( .A1(n816), .A2(n815), .ZN(n964) );
  AND2_X1 U146bar ( .A1(n816bar), .A2(n815bar), .ZN(n964bar) );
  OR2_X1 U147 ( .A1(n814), .A2(n813), .ZN(n815) );
  AND2_X1 U147bar ( .A1(n814bar), .A2(n813bar), .ZN(n815bar) );
  OR2_X1 U148 ( .A1(n812), .A2(n811), .ZN(n813) );
  AND2_X1 U148bar ( .A1(n812bar), .A2(n811bar), .ZN(n813bar) );
  OR2_X1 U149 ( .A1(in[122]), .A2(in[111]), .ZN(n811) );
  AND2_X1 U149bar ( .A1(inbar[122]), .A2(inbar[111]), .ZN(n811bar) );
  OR2_X1 U150 ( .A1(in[154]), .A2(in[151]), .ZN(n812) );
  AND2_X1 U150bar ( .A1(inbar[154]), .A2(inbar[151]), .ZN(n812bar) );
  OR2_X1 U151 ( .A1(n810), .A2(n809), .ZN(n814) );
  AND2_X1 U151bar ( .A1(n810bar), .A2(n809bar), .ZN(n814bar) );
  OR2_X1 U152 ( .A1(in[187]), .A2(in[177]), .ZN(n809) );
  AND2_X1 U152bar ( .A1(inbar[187]), .A2(inbar[177]), .ZN(n809bar) );
  OR2_X1 U153 ( .A1(in[200]), .A2(in[192]), .ZN(n810) );
  AND2_X1 U153bar ( .A1(inbar[200]), .A2(inbar[192]), .ZN(n810bar) );
  OR2_X1 U154 ( .A1(n808), .A2(n807), .ZN(n816) );
  AND2_X1 U154bar ( .A1(n808bar), .A2(n807bar), .ZN(n816bar) );
  OR2_X1 U155 ( .A1(n806), .A2(n805), .ZN(n807) );
  AND2_X1 U155bar ( .A1(n806bar), .A2(n805bar), .ZN(n807bar) );
  OR2_X1 U156 ( .A1(in[225]), .A2(in[207]), .ZN(n805) );
  AND2_X1 U156bar ( .A1(inbar[225]), .A2(inbar[207]), .ZN(n805bar) );
  OR2_X1 U157 ( .A1(in[98]), .A2(in[226]), .ZN(n806) );
  AND2_X1 U157bar ( .A1(inbar[98]), .A2(inbar[226]), .ZN(n806bar) );
  OR2_X1 U158 ( .A1(n804), .A2(n803), .ZN(n808) );
  AND2_X1 U158bar ( .A1(n804bar), .A2(n803bar), .ZN(n808bar) );
  OR2_X1 U159 ( .A1(in_20), .A2(in_16), .ZN(n803) );
  AND2_X1 U159bar ( .A1(in_20bar), .A2(in_16bar), .ZN(n803bar) );
  OR2_X1 U160 ( .A1(in_55), .A2(in_45), .ZN(n804) );
  AND2_X1 U160bar ( .A1(in_55bar), .A2(in_45bar), .ZN(n804bar) );
  OR2_X1 U161 ( .A1(n802), .A2(n801), .ZN(n824) );
  AND2_X1 U161bar ( .A1(n802bar), .A2(n801bar), .ZN(n824bar) );
  OR2_X1 U162 ( .A1(in[162]), .A2(in[149]), .ZN(n801) );
  AND2_X1 U162bar ( .A1(inbar[162]), .A2(inbar[149]), .ZN(n801bar) );
  OR2_X1 U163 ( .A1(in[163]), .A2(n800), .ZN(n802) );
  AND2_X1 U163bar ( .A1(inbar[163]), .A2(n800bar), .ZN(n802bar) );
  OR2_X1 U164 ( .A1(in[191]), .A2(in[189]), .ZN(n800) );
  AND2_X1 U164bar ( .A1(inbar[191]), .A2(inbar[189]), .ZN(n800bar) );
  OR2_X1 U165 ( .A1(n799), .A2(n798), .ZN(n826) );
  AND2_X1 U165bar ( .A1(n799bar), .A2(n798bar), .ZN(n826bar) );
  OR2_X1 U166 ( .A1(n797), .A2(n796), .ZN(n798) );
  AND2_X1 U166bar ( .A1(n797bar), .A2(n796bar), .ZN(n798bar) );
  OR2_X1 U167 ( .A1(in[212]), .A2(in[193]), .ZN(n796) );
  AND2_X1 U167bar ( .A1(inbar[212]), .A2(inbar[193]), .ZN(n796bar) );
  OR2_X1 U168 ( .A1(in[238]), .A2(n795), .ZN(n797) );
  AND2_X1 U168bar ( .A1(inbar[238]), .A2(n795bar), .ZN(n797bar) );
  OR2_X1 U169 ( .A1(in[88]), .A2(in[247]), .ZN(n795) );
  AND2_X1 U169bar ( .A1(inbar[88]), .A2(inbar[247]), .ZN(n795bar) );
  OR2_X1 U170 ( .A1(n794), .A2(n793), .ZN(n799) );
  AND2_X1 U170bar ( .A1(n794bar), .A2(n793bar), .ZN(n799bar) );
  OR2_X1 U171 ( .A1(in[94]), .A2(in[92]), .ZN(n793) );
  AND2_X1 U171bar ( .A1(inbar[94]), .A2(inbar[92]), .ZN(n793bar) );
  OR2_X1 U172 ( .A1(in_52), .A2(n792), .ZN(n794) );
  AND2_X1 U172bar ( .A1(in_52bar), .A2(n792bar), .ZN(n794bar) );
  OR2_X1 U173 ( .A1(in_70), .A2(in_67), .ZN(n792) );
  AND2_X1 U173bar ( .A1(in_70bar), .A2(in_67bar), .ZN(n792bar) );
  OR2_X1 U174 ( .A1(n791), .A2(n790), .ZN(out[2]) );
  AND2_X1 U174bar ( .A1(n791bar), .A2(n790bar), .ZN(outbar[2]) );
  OR2_X1 U175 ( .A1(n789), .A2(n788), .ZN(n790) );
  AND2_X1 U175bar ( .A1(n789bar), .A2(n788bar), .ZN(n790bar) );
  OR2_X1 U176 ( .A1(n787), .A2(n786), .ZN(n788) );
  AND2_X1 U176bar ( .A1(n787bar), .A2(n786bar), .ZN(n788bar) );
  OR2_X1 U177 ( .A1(n819), .A2(n785), .ZN(n786) );
  AND2_X1 U177bar ( .A1(n819bar), .A2(n785bar), .ZN(n786bar) );
  OR2_X1 U178 ( .A1(n784), .A2(n783), .ZN(n819) );
  AND2_X1 U178bar ( .A1(n784bar), .A2(n783bar), .ZN(n819bar) );
  OR2_X1 U179 ( .A1(n782), .A2(n781), .ZN(n783) );
  AND2_X1 U179bar ( .A1(n782bar), .A2(n781bar), .ZN(n783bar) );
  OR2_X1 U180 ( .A1(n780), .A2(n779), .ZN(n781) );
  AND2_X1 U180bar ( .A1(n780bar), .A2(n779bar), .ZN(n781bar) );
  OR2_X1 U181 ( .A1(n962), .A2(n778), .ZN(n779) );
  AND2_X1 U181bar ( .A1(n962bar), .A2(n778bar), .ZN(n779bar) );
  OR2_X1 U182 ( .A1(n777), .A2(n776), .ZN(n962) );
  AND2_X1 U182bar ( .A1(n777bar), .A2(n776bar), .ZN(n962bar) );
  OR2_X1 U183 ( .A1(n775), .A2(n774), .ZN(n776) );
  AND2_X1 U183bar ( .A1(n775bar), .A2(n774bar), .ZN(n776bar) );
  OR2_X1 U184 ( .A1(n773), .A2(n772), .ZN(n774) );
  AND2_X1 U184bar ( .A1(n773bar), .A2(n772bar), .ZN(n774bar) );
  OR2_X1 U185 ( .A1(in[131]), .A2(in[120]), .ZN(n772) );
  AND2_X1 U185bar ( .A1(inbar[131]), .A2(inbar[120]), .ZN(n772bar) );
  OR2_X1 U186 ( .A1(in[153]), .A2(in[147]), .ZN(n773) );
  AND2_X1 U186bar ( .A1(inbar[153]), .A2(inbar[147]), .ZN(n773bar) );
  OR2_X1 U187 ( .A1(n771), .A2(n770), .ZN(n775) );
  AND2_X1 U187bar ( .A1(n771bar), .A2(n770bar), .ZN(n775bar) );
  OR2_X1 U188 ( .A1(in[170]), .A2(in[156]), .ZN(n770) );
  AND2_X1 U188bar ( .A1(inbar[170]), .A2(inbar[156]), .ZN(n770bar) );
  OR2_X1 U189 ( .A1(in[223]), .A2(in[190]), .ZN(n771) );
  AND2_X1 U189bar ( .A1(inbar[223]), .A2(inbar[190]), .ZN(n771bar) );
  OR2_X1 U190 ( .A1(n769), .A2(n768), .ZN(n777) );
  AND2_X1 U190bar ( .A1(n769bar), .A2(n768bar), .ZN(n777bar) );
  OR2_X1 U191 ( .A1(n767), .A2(n766), .ZN(n768) );
  AND2_X1 U191bar ( .A1(n767bar), .A2(n766bar), .ZN(n768bar) );
  OR2_X1 U192 ( .A1(in[236]), .A2(in[230]), .ZN(n766) );
  AND2_X1 U192bar ( .A1(inbar[236]), .A2(inbar[230]), .ZN(n766bar) );
  OR2_X1 U193 ( .A1(in[85]), .A2(in[240]), .ZN(n767) );
  AND2_X1 U193bar ( .A1(inbar[85]), .A2(inbar[240]), .ZN(n767bar) );
  OR2_X1 U194 ( .A1(n765), .A2(n764), .ZN(n769) );
  AND2_X1 U194bar ( .A1(n765bar), .A2(n764bar), .ZN(n769bar) );
  OR2_X1 U195 ( .A1(in_12), .A2(in[90]), .ZN(n764) );
  AND2_X1 U195bar ( .A1(in_12bar), .A2(inbar[90]), .ZN(n764bar) );
  OR2_X1 U196 ( .A1(in_39), .A2(in_28), .ZN(n765) );
  AND2_X1 U196bar ( .A1(in_39bar), .A2(in_28bar), .ZN(n765bar) );
  OR2_X1 U197 ( .A1(in[109]), .A2(n763), .ZN(n780) );
  AND2_X1 U197bar ( .A1(inbar[109]), .A2(n763bar), .ZN(n780bar) );
  OR2_X1 U198 ( .A1(n762), .A2(n761), .ZN(n782) );
  AND2_X1 U198bar ( .A1(n762bar), .A2(n761bar), .ZN(n782bar) );
  OR2_X1 U199 ( .A1(in[138]), .A2(in[129]), .ZN(n761) );
  AND2_X1 U199bar ( .A1(inbar[138]), .A2(inbar[129]), .ZN(n761bar) );
  OR2_X1 U200 ( .A1(in[157]), .A2(n760), .ZN(n762) );
  AND2_X1 U200bar ( .A1(inbar[157]), .A2(n760bar), .ZN(n762bar) );
  OR2_X1 U201 ( .A1(in[182]), .A2(in[167]), .ZN(n760) );
  AND2_X1 U201bar ( .A1(inbar[182]), .A2(inbar[167]), .ZN(n760bar) );
  OR2_X1 U202 ( .A1(n759), .A2(n758), .ZN(n784) );
  AND2_X1 U202bar ( .A1(n759bar), .A2(n758bar), .ZN(n784bar) );
  OR2_X1 U203 ( .A1(n757), .A2(n756), .ZN(n758) );
  AND2_X1 U203bar ( .A1(n757bar), .A2(n756bar), .ZN(n758bar) );
  OR2_X1 U204 ( .A1(in[195]), .A2(in[184]), .ZN(n756) );
  AND2_X1 U204bar ( .A1(inbar[195]), .A2(inbar[184]), .ZN(n756bar) );
  OR2_X1 U205 ( .A1(in[196]), .A2(n755), .ZN(n757) );
  AND2_X1 U205bar ( .A1(inbar[196]), .A2(n755bar), .ZN(n757bar) );
  OR2_X1 U206 ( .A1(in[215]), .A2(in[209]), .ZN(n755) );
  AND2_X1 U206bar ( .A1(inbar[215]), .A2(inbar[209]), .ZN(n755bar) );
  OR2_X1 U207 ( .A1(n754), .A2(n753), .ZN(n759) );
  AND2_X1 U207bar ( .A1(n754bar), .A2(n753bar), .ZN(n759bar) );
  OR2_X1 U208 ( .A1(in[93]), .A2(in[233]), .ZN(n753) );
  AND2_X1 U208bar ( .A1(inbar[93]), .A2(inbar[233]), .ZN(n753bar) );
  OR2_X1 U209 ( .A1(in_1), .A2(n752), .ZN(n754) );
  AND2_X1 U209bar ( .A1(in_1bar), .A2(n752bar), .ZN(n754bar) );
  OR2_X1 U210 ( .A1(in_69), .A2(in_66), .ZN(n752) );
  AND2_X1 U210bar ( .A1(in_69bar), .A2(in_66bar), .ZN(n752bar) );
  OR2_X1 U211 ( .A1(n966), .A2(n751), .ZN(n787) );
  AND2_X1 U211bar ( .A1(n966bar), .A2(n751bar), .ZN(n787bar) );
  OR2_X1 U212 ( .A1(in[134]), .A2(n750), .ZN(n751) );
  AND2_X1 U212bar ( .A1(inbar[134]), .A2(n750bar), .ZN(n751bar) );
  OR2_X1 U213 ( .A1(n749), .A2(n748), .ZN(n966) );
  AND2_X1 U213bar ( .A1(n749bar), .A2(n748bar), .ZN(n966bar) );
  OR2_X1 U214 ( .A1(n747), .A2(n746), .ZN(n748) );
  AND2_X1 U214bar ( .A1(n747bar), .A2(n746bar), .ZN(n748bar) );
  OR2_X1 U215 ( .A1(n745), .A2(n744), .ZN(n746) );
  AND2_X1 U215bar ( .A1(n745bar), .A2(n744bar), .ZN(n746bar) );
  OR2_X1 U216 ( .A1(in[136]), .A2(in[121]), .ZN(n744) );
  AND2_X1 U216bar ( .A1(inbar[136]), .A2(inbar[121]), .ZN(n744bar) );
  OR2_X1 U217 ( .A1(in[186]), .A2(in[174]), .ZN(n745) );
  AND2_X1 U217bar ( .A1(inbar[186]), .A2(inbar[174]), .ZN(n745bar) );
  OR2_X1 U218 ( .A1(n743), .A2(n742), .ZN(n747) );
  AND2_X1 U218bar ( .A1(n743bar), .A2(n742bar), .ZN(n747bar) );
  OR2_X1 U219 ( .A1(in[198]), .A2(in[197]), .ZN(n742) );
  AND2_X1 U219bar ( .A1(inbar[198]), .A2(inbar[197]), .ZN(n742bar) );
  OR2_X1 U220 ( .A1(in[214]), .A2(in[199]), .ZN(n743) );
  AND2_X1 U220bar ( .A1(inbar[214]), .A2(inbar[199]), .ZN(n743bar) );
  OR2_X1 U221 ( .A1(n741), .A2(n740), .ZN(n749) );
  AND2_X1 U221bar ( .A1(n741bar), .A2(n740bar), .ZN(n749bar) );
  OR2_X1 U222 ( .A1(n739), .A2(n738), .ZN(n740) );
  AND2_X1 U222bar ( .A1(n739bar), .A2(n738bar), .ZN(n740bar) );
  OR2_X1 U223 ( .A1(in[231]), .A2(in[220]), .ZN(n738) );
  AND2_X1 U223bar ( .A1(inbar[231]), .A2(inbar[220]), .ZN(n738bar) );
  OR2_X1 U224 ( .A1(in_25), .A2(in[245]), .ZN(n739) );
  AND2_X1 U224bar ( .A1(in_25bar), .A2(inbar[245]), .ZN(n739bar) );
  OR2_X1 U225 ( .A1(n737), .A2(n736), .ZN(n741) );
  AND2_X1 U225bar ( .A1(n737bar), .A2(n736bar), .ZN(n741bar) );
  OR2_X1 U226 ( .A1(in_53), .A2(in_29), .ZN(n736) );
  AND2_X1 U226bar ( .A1(in_53bar), .A2(in_29bar), .ZN(n736bar) );
  OR2_X1 U227 ( .A1(in_79), .A2(in_74), .ZN(n737) );
  AND2_X1 U227bar ( .A1(in_79bar), .A2(in_74bar), .ZN(n737bar) );
  OR2_X1 U228 ( .A1(n735), .A2(n734), .ZN(n789) );
  AND2_X1 U228bar ( .A1(n735bar), .A2(n734bar), .ZN(n789bar) );
  OR2_X1 U229 ( .A1(in[152]), .A2(in[140]), .ZN(n734) );
  AND2_X1 U229bar ( .A1(inbar[152]), .A2(inbar[140]), .ZN(n734bar) );
  OR2_X1 U230 ( .A1(in[155]), .A2(n733), .ZN(n735) );
  AND2_X1 U230bar ( .A1(inbar[155]), .A2(n733bar), .ZN(n735bar) );
  OR2_X1 U231 ( .A1(in[166]), .A2(in[165]), .ZN(n733) );
  AND2_X1 U231bar ( .A1(inbar[166]), .A2(inbar[165]), .ZN(n733bar) );
  OR2_X1 U232 ( .A1(n732), .A2(n731), .ZN(n791) );
  AND2_X1 U232bar ( .A1(n732bar), .A2(n731bar), .ZN(n791bar) );
  OR2_X1 U233 ( .A1(n730), .A2(n729), .ZN(n731) );
  AND2_X1 U233bar ( .A1(n730bar), .A2(n729bar), .ZN(n731bar) );
  OR2_X1 U234 ( .A1(in[202]), .A2(in[185]), .ZN(n729) );
  AND2_X1 U234bar ( .A1(inbar[202]), .A2(inbar[185]), .ZN(n729bar) );
  OR2_X1 U235 ( .A1(in[211]), .A2(n728), .ZN(n730) );
  AND2_X1 U235bar ( .A1(inbar[211]), .A2(n728bar), .ZN(n730bar) );
  OR2_X1 U236 ( .A1(in[255]), .A2(in[253]), .ZN(n728) );
  AND2_X1 U236bar ( .A1(inbar[255]), .A2(inbar[253]), .ZN(n728bar) );
  OR2_X1 U237 ( .A1(n727), .A2(n726), .ZN(n732) );
  AND2_X1 U237bar ( .A1(n727bar), .A2(n726bar), .ZN(n732bar) );
  OR2_X1 U238 ( .A1(in_35), .A2(in_15), .ZN(n726) );
  AND2_X1 U238bar ( .A1(in_35bar), .A2(in_15bar), .ZN(n726bar) );
  OR2_X1 U239 ( .A1(in_36), .A2(n725), .ZN(n727) );
  AND2_X1 U239bar ( .A1(in_36bar), .A2(n725bar), .ZN(n727bar) );
  OR2_X1 U240 ( .A1(in_48), .A2(in_40), .ZN(n725) );
  AND2_X1 U240bar ( .A1(in_48bar), .A2(in_40bar), .ZN(n725bar) );
  OR2_X1 U241 ( .A1(n724), .A2(n723), .ZN(out[1]) );
  AND2_X1 U241bar ( .A1(n724bar), .A2(n723bar), .ZN(outbar[1]) );
  OR2_X1 U242 ( .A1(n722), .A2(n721), .ZN(n723) );
  AND2_X1 U242bar ( .A1(n722bar), .A2(n721bar), .ZN(n723bar) );
  OR2_X1 U243 ( .A1(n720), .A2(n719), .ZN(n721) );
  AND2_X1 U243bar ( .A1(n720bar), .A2(n719bar), .ZN(n721bar) );
  OR2_X1 U244 ( .A1(n921), .A2(n887), .ZN(n719) );
  AND2_X1 U244bar ( .A1(n921bar), .A2(n887bar), .ZN(n719bar) );
  OR2_X1 U245 ( .A1(n718), .A2(n717), .ZN(n887) );
  AND2_X1 U245bar ( .A1(n718bar), .A2(n717bar), .ZN(n887bar) );
  OR2_X1 U246 ( .A1(n716), .A2(n715), .ZN(n717) );
  AND2_X1 U246bar ( .A1(n716bar), .A2(n715bar), .ZN(n717bar) );
  OR2_X1 U247 ( .A1(n714), .A2(n713), .ZN(n715) );
  AND2_X1 U247bar ( .A1(n714bar), .A2(n713bar), .ZN(n715bar) );
  OR2_X1 U248 ( .A1(in[116]), .A2(in[110]), .ZN(n713) );
  AND2_X1 U248bar ( .A1(inbar[116]), .A2(inbar[110]), .ZN(n713bar) );
  OR2_X1 U249 ( .A1(in[133]), .A2(in[130]), .ZN(n714) );
  AND2_X1 U249bar ( .A1(inbar[133]), .A2(inbar[130]), .ZN(n714bar) );
  OR2_X1 U250 ( .A1(n712), .A2(n711), .ZN(n716) );
  AND2_X1 U250bar ( .A1(n712bar), .A2(n711bar), .ZN(n716bar) );
  OR2_X1 U251 ( .A1(in[203]), .A2(in[135]), .ZN(n711) );
  AND2_X1 U251bar ( .A1(inbar[203]), .A2(inbar[135]), .ZN(n711bar) );
  OR2_X1 U252 ( .A1(in[232]), .A2(in[223]), .ZN(n712) );
  AND2_X1 U252bar ( .A1(inbar[232]), .A2(inbar[223]), .ZN(n712bar) );
  OR2_X1 U253 ( .A1(n710), .A2(n709), .ZN(n718) );
  AND2_X1 U253bar ( .A1(n710bar), .A2(n709bar), .ZN(n718bar) );
  OR2_X1 U254 ( .A1(n708), .A2(n707), .ZN(n709) );
  AND2_X1 U254bar ( .A1(n708bar), .A2(n707bar), .ZN(n709bar) );
  OR2_X1 U255 ( .A1(in[255]), .A2(in[233]), .ZN(n707) );
  AND2_X1 U255bar ( .A1(inbar[255]), .A2(inbar[233]), .ZN(n707bar) );
  OR2_X1 U256 ( .A1(in_53), .A2(in_34), .ZN(n708) );
  AND2_X1 U256bar ( .A1(in_53bar), .A2(in_34bar), .ZN(n708bar) );
  OR2_X1 U257 ( .A1(n706), .A2(n705), .ZN(n710) );
  AND2_X1 U257bar ( .A1(n706bar), .A2(n705bar), .ZN(n710bar) );
  OR2_X1 U258 ( .A1(in_57), .A2(in_55), .ZN(n705) );
  AND2_X1 U258bar ( .A1(in_57bar), .A2(in_55bar), .ZN(n705bar) );
  OR2_X1 U259 ( .A1(in_68), .A2(in_67), .ZN(n706) );
  AND2_X1 U259bar ( .A1(in_68bar), .A2(in_67bar), .ZN(n706bar) );
  OR2_X1 U260 ( .A1(n704), .A2(n703), .ZN(n921) );
  AND2_X1 U260bar ( .A1(n704bar), .A2(n703bar), .ZN(n921bar) );
  OR2_X1 U261 ( .A1(n702), .A2(n701), .ZN(n703) );
  AND2_X1 U261bar ( .A1(n702bar), .A2(n701bar), .ZN(n703bar) );
  OR2_X1 U262 ( .A1(n700), .A2(n699), .ZN(n701) );
  AND2_X1 U262bar ( .A1(n700bar), .A2(n699bar), .ZN(n701bar) );
  OR2_X1 U263 ( .A1(n944), .A2(n872), .ZN(n699) );
  AND2_X1 U263bar ( .A1(n944bar), .A2(n872bar), .ZN(n699bar) );
  OR2_X1 U264 ( .A1(n698), .A2(n697), .ZN(n872) );
  AND2_X1 U264bar ( .A1(n698bar), .A2(n697bar), .ZN(n872bar) );
  OR2_X1 U265 ( .A1(n696), .A2(n695), .ZN(n697) );
  AND2_X1 U265bar ( .A1(n696bar), .A2(n695bar), .ZN(n697bar) );
  OR2_X1 U266 ( .A1(n694), .A2(n693), .ZN(n695) );
  AND2_X1 U266bar ( .A1(n694bar), .A2(n693bar), .ZN(n695bar) );
  OR2_X1 U267 ( .A1(in[121]), .A2(in[102]), .ZN(n693) );
  AND2_X1 U267bar ( .A1(inbar[121]), .A2(inbar[102]), .ZN(n693bar) );
  OR2_X1 U268 ( .A1(in[162]), .A2(in[161]), .ZN(n694) );
  AND2_X1 U268bar ( .A1(inbar[162]), .A2(inbar[161]), .ZN(n694bar) );
  OR2_X1 U269 ( .A1(n692), .A2(n691), .ZN(n696) );
  AND2_X1 U269bar ( .A1(n692bar), .A2(n691bar), .ZN(n696bar) );
  OR2_X1 U270 ( .A1(in[192]), .A2(in[178]), .ZN(n691) );
  AND2_X1 U270bar ( .A1(inbar[192]), .A2(inbar[178]), .ZN(n691bar) );
  OR2_X1 U271 ( .A1(in[244]), .A2(in[209]), .ZN(n692) );
  AND2_X1 U271bar ( .A1(inbar[244]), .A2(inbar[209]), .ZN(n692bar) );
  OR2_X1 U272 ( .A1(n690), .A2(n689), .ZN(n698) );
  AND2_X1 U272bar ( .A1(n690bar), .A2(n689bar), .ZN(n698bar) );
  OR2_X1 U273 ( .A1(n688), .A2(n687), .ZN(n689) );
  AND2_X1 U273bar ( .A1(n688bar), .A2(n687bar), .ZN(n689bar) );
  OR2_X1 U274 ( .A1(in[90]), .A2(in[254]), .ZN(n687) );
  AND2_X1 U274bar ( .A1(inbar[90]), .A2(inbar[254]), .ZN(n687bar) );
  OR2_X1 U275 ( .A1(in_36), .A2(in_32), .ZN(n688) );
  AND2_X1 U275bar ( .A1(in_36bar), .A2(in_32bar), .ZN(n688bar) );
  OR2_X1 U276 ( .A1(n686), .A2(n685), .ZN(n690) );
  AND2_X1 U276bar ( .A1(n686bar), .A2(n685bar), .ZN(n690bar) );
  OR2_X1 U277 ( .A1(in_62), .A2(in_37), .ZN(n685) );
  AND2_X1 U277bar ( .A1(in_62bar), .A2(in_37bar), .ZN(n685bar) );
  OR2_X1 U278 ( .A1(in_75), .A2(in_73), .ZN(n686) );
  AND2_X1 U278bar ( .A1(in_75bar), .A2(in_73bar), .ZN(n686bar) );
  OR2_X1 U279 ( .A1(n684), .A2(n683), .ZN(n944) );
  AND2_X1 U279bar ( .A1(n684bar), .A2(n683bar), .ZN(n944bar) );
  OR2_X1 U280 ( .A1(n682), .A2(n681), .ZN(n683) );
  AND2_X1 U280bar ( .A1(n682bar), .A2(n681bar), .ZN(n683bar) );
  OR2_X1 U281 ( .A1(n680), .A2(n679), .ZN(n681) );
  AND2_X1 U281bar ( .A1(n680bar), .A2(n679bar), .ZN(n681bar) );
  OR2_X1 U282 ( .A1(in[171]), .A2(in[153]), .ZN(n679) );
  AND2_X1 U282bar ( .A1(inbar[171]), .A2(inbar[153]), .ZN(n679bar) );
  OR2_X1 U283 ( .A1(in[187]), .A2(in[176]), .ZN(n680) );
  AND2_X1 U283bar ( .A1(inbar[187]), .A2(inbar[176]), .ZN(n680bar) );
  OR2_X1 U284 ( .A1(n678), .A2(n677), .ZN(n682) );
  AND2_X1 U284bar ( .A1(n678bar), .A2(n677bar), .ZN(n682bar) );
  OR2_X1 U285 ( .A1(in[245]), .A2(in[211]), .ZN(n677) );
  AND2_X1 U285bar ( .A1(inbar[245]), .A2(inbar[211]), .ZN(n677bar) );
  OR2_X1 U286 ( .A1(in[97]), .A2(in[88]), .ZN(n678) );
  AND2_X1 U286bar ( .A1(inbar[97]), .A2(inbar[88]), .ZN(n678bar) );
  OR2_X1 U287 ( .A1(n676), .A2(n675), .ZN(n684) );
  AND2_X1 U287bar ( .A1(n676bar), .A2(n675bar), .ZN(n684bar) );
  OR2_X1 U288 ( .A1(n674), .A2(n673), .ZN(n675) );
  AND2_X1 U288bar ( .A1(n674bar), .A2(n673bar), .ZN(n675bar) );
  OR2_X1 U289 ( .A1(in_10), .A2(in_0), .ZN(n673) );
  AND2_X1 U289bar ( .A1(in_10bar), .A2(in_0bar), .ZN(n673bar) );
  OR2_X1 U290 ( .A1(in_59), .A2(in_5), .ZN(n674) );
  AND2_X1 U290bar ( .A1(in_59bar), .A2(in_5bar), .ZN(n674bar) );
  OR2_X1 U291 ( .A1(n672), .A2(n671), .ZN(n676) );
  AND2_X1 U291bar ( .A1(n672bar), .A2(n671bar), .ZN(n676bar) );
  OR2_X1 U292 ( .A1(in_60), .A2(in_6), .ZN(n671) );
  AND2_X1 U292bar ( .A1(in_60bar), .A2(in_6bar), .ZN(n671bar) );
  OR2_X1 U293 ( .A1(in_77), .A2(in_69), .ZN(n672) );
  AND2_X1 U293bar ( .A1(in_77bar), .A2(in_69bar), .ZN(n672bar) );
  OR2_X1 U294 ( .A1(in[113]), .A2(n864), .ZN(n700) );
  AND2_X1 U294bar ( .A1(inbar[113]), .A2(n864bar), .ZN(n700bar) );
  OR2_X1 U295 ( .A1(n670), .A2(n669), .ZN(n864) );
  AND2_X1 U295bar ( .A1(n670bar), .A2(n669bar), .ZN(n864bar) );
  OR2_X1 U296 ( .A1(n668), .A2(n667), .ZN(n669) );
  AND2_X1 U296bar ( .A1(n668bar), .A2(n667bar), .ZN(n669bar) );
  OR2_X1 U297 ( .A1(n666), .A2(n665), .ZN(n667) );
  AND2_X1 U297bar ( .A1(n666bar), .A2(n665bar), .ZN(n667bar) );
  OR2_X1 U298 ( .A1(in[125]), .A2(in[107]), .ZN(n665) );
  AND2_X1 U298bar ( .A1(inbar[125]), .A2(inbar[107]), .ZN(n665bar) );
  OR2_X1 U299 ( .A1(in[138]), .A2(in[126]), .ZN(n666) );
  AND2_X1 U299bar ( .A1(inbar[138]), .A2(inbar[126]), .ZN(n666bar) );
  OR2_X1 U300 ( .A1(n664), .A2(n663), .ZN(n668) );
  AND2_X1 U300bar ( .A1(n664bar), .A2(n663bar), .ZN(n668bar) );
  OR2_X1 U301 ( .A1(in[189]), .A2(in[143]), .ZN(n663) );
  AND2_X1 U301bar ( .A1(inbar[189]), .A2(inbar[143]), .ZN(n663bar) );
  OR2_X1 U302 ( .A1(in[99]), .A2(in[214]), .ZN(n664) );
  AND2_X1 U302bar ( .A1(inbar[99]), .A2(inbar[214]), .ZN(n664bar) );
  OR2_X1 U303 ( .A1(n662), .A2(n661), .ZN(n670) );
  AND2_X1 U303bar ( .A1(n662bar), .A2(n661bar), .ZN(n670bar) );
  OR2_X1 U304 ( .A1(n660), .A2(n659), .ZN(n661) );
  AND2_X1 U304bar ( .A1(n660bar), .A2(n659bar), .ZN(n661bar) );
  OR2_X1 U305 ( .A1(in_15), .A2(in_12), .ZN(n659) );
  AND2_X1 U305bar ( .A1(in_15bar), .A2(in_12bar), .ZN(n659bar) );
  OR2_X1 U306 ( .A1(in_20), .A2(in_2), .ZN(n660) );
  AND2_X1 U306bar ( .A1(in_20bar), .A2(in_2bar), .ZN(n660bar) );
  OR2_X1 U307 ( .A1(n658), .A2(n657), .ZN(n662) );
  AND2_X1 U307bar ( .A1(n658bar), .A2(n657bar), .ZN(n662bar) );
  OR2_X1 U308 ( .A1(in_30), .A2(in_3), .ZN(n657) );
  AND2_X1 U308bar ( .A1(in_30bar), .A2(in_3bar), .ZN(n657bar) );
  OR2_X1 U309 ( .A1(in_4), .A2(in_38), .ZN(n658) );
  AND2_X1 U309bar ( .A1(in_4bar), .A2(in_38bar), .ZN(n658bar) );
  OR2_X1 U310 ( .A1(n656), .A2(n655), .ZN(n702) );
  AND2_X1 U310bar ( .A1(n656bar), .A2(n655bar), .ZN(n702bar) );
  OR2_X1 U311 ( .A1(in[148]), .A2(in[137]), .ZN(n655) );
  AND2_X1 U311bar ( .A1(inbar[148]), .A2(inbar[137]), .ZN(n655bar) );
  OR2_X1 U312 ( .A1(in[149]), .A2(n654), .ZN(n656) );
  AND2_X1 U312bar ( .A1(inbar[149]), .A2(n654bar), .ZN(n656bar) );
  OR2_X1 U313 ( .A1(in[195]), .A2(in[190]), .ZN(n654) );
  AND2_X1 U313bar ( .A1(inbar[195]), .A2(inbar[190]), .ZN(n654bar) );
  OR2_X1 U314 ( .A1(n653), .A2(n652), .ZN(n704) );
  AND2_X1 U314bar ( .A1(n653bar), .A2(n652bar), .ZN(n704bar) );
  OR2_X1 U315 ( .A1(n651), .A2(n650), .ZN(n652) );
  AND2_X1 U315bar ( .A1(n651bar), .A2(n650bar), .ZN(n652bar) );
  OR2_X1 U316 ( .A1(in[98]), .A2(in[197]), .ZN(n650) );
  AND2_X1 U316bar ( .A1(inbar[98]), .A2(inbar[197]), .ZN(n650bar) );
  OR2_X1 U317 ( .A1(in_11), .A2(n649), .ZN(n651) );
  AND2_X1 U317bar ( .A1(in_11bar), .A2(n649bar), .ZN(n651bar) );
  OR2_X1 U318 ( .A1(in_26), .A2(in_14), .ZN(n649) );
  AND2_X1 U318bar ( .A1(in_26bar), .A2(in_14bar), .ZN(n649bar) );
  OR2_X1 U319 ( .A1(n648), .A2(n647), .ZN(n653) );
  AND2_X1 U319bar ( .A1(n648bar), .A2(n647bar), .ZN(n653bar) );
  OR2_X1 U320 ( .A1(in_35), .A2(in_27), .ZN(n647) );
  AND2_X1 U320bar ( .A1(in_35bar), .A2(in_27bar), .ZN(n647bar) );
  OR2_X1 U321 ( .A1(in_50), .A2(n646), .ZN(n648) );
  AND2_X1 U321bar ( .A1(in_50bar), .A2(n646bar), .ZN(n648bar) );
  OR2_X1 U322 ( .A1(in_78), .A2(in_61), .ZN(n646) );
  AND2_X1 U322bar ( .A1(in_78bar), .A2(in_61bar), .ZN(n646bar) );
  OR2_X1 U323 ( .A1(n942), .A2(n645), .ZN(n720) );
  AND2_X1 U323bar ( .A1(n942bar), .A2(n645bar), .ZN(n720bar) );
  OR2_X1 U324 ( .A1(in[106]), .A2(n863), .ZN(n645) );
  AND2_X1 U324bar ( .A1(inbar[106]), .A2(n863bar), .ZN(n645bar) );
  OR2_X1 U325 ( .A1(n644), .A2(n643), .ZN(n863) );
  AND2_X1 U325bar ( .A1(n644bar), .A2(n643bar), .ZN(n863bar) );
  OR2_X1 U326 ( .A1(n642), .A2(n641), .ZN(n643) );
  AND2_X1 U326bar ( .A1(n642bar), .A2(n641bar), .ZN(n643bar) );
  OR2_X1 U327 ( .A1(n640), .A2(n639), .ZN(n641) );
  AND2_X1 U327bar ( .A1(n640bar), .A2(n639bar), .ZN(n641bar) );
  OR2_X1 U328 ( .A1(in[127]), .A2(in[122]), .ZN(n639) );
  AND2_X1 U328bar ( .A1(inbar[127]), .A2(inbar[122]), .ZN(n639bar) );
  OR2_X1 U329 ( .A1(in[156]), .A2(in[132]), .ZN(n640) );
  AND2_X1 U329bar ( .A1(inbar[156]), .A2(inbar[132]), .ZN(n640bar) );
  OR2_X1 U330 ( .A1(n638), .A2(n637), .ZN(n642) );
  AND2_X1 U330bar ( .A1(n638bar), .A2(n637bar), .ZN(n642bar) );
  OR2_X1 U331 ( .A1(in[159]), .A2(in[157]), .ZN(n637) );
  AND2_X1 U331bar ( .A1(inbar[159]), .A2(inbar[157]), .ZN(n637bar) );
  OR2_X1 U332 ( .A1(in[185]), .A2(in[169]), .ZN(n638) );
  AND2_X1 U332bar ( .A1(inbar[185]), .A2(inbar[169]), .ZN(n638bar) );
  OR2_X1 U333 ( .A1(n636), .A2(n635), .ZN(n644) );
  AND2_X1 U333bar ( .A1(n636bar), .A2(n635bar), .ZN(n644bar) );
  OR2_X1 U334 ( .A1(n634), .A2(n633), .ZN(n635) );
  AND2_X1 U334bar ( .A1(n634bar), .A2(n633bar), .ZN(n635bar) );
  OR2_X1 U335 ( .A1(in[239]), .A2(in[218]), .ZN(n633) );
  AND2_X1 U335bar ( .A1(inbar[239]), .A2(inbar[218]), .ZN(n633bar) );
  OR2_X1 U336 ( .A1(in_13), .A2(in[87]), .ZN(n634) );
  AND2_X1 U336bar ( .A1(in_13bar), .A2(inbar[87]), .ZN(n634bar) );
  OR2_X1 U337 ( .A1(n632), .A2(n631), .ZN(n636) );
  AND2_X1 U337bar ( .A1(n632bar), .A2(n631bar), .ZN(n636bar) );
  OR2_X1 U338 ( .A1(in_72), .A2(in_70), .ZN(n631) );
  AND2_X1 U338bar ( .A1(in_72bar), .A2(in_70bar), .ZN(n631bar) );
  OR2_X1 U339 ( .A1(in_80), .A2(in_74), .ZN(n632) );
  AND2_X1 U339bar ( .A1(in_80bar), .A2(in_74bar), .ZN(n632bar) );
  OR2_X1 U340 ( .A1(n630), .A2(n629), .ZN(n942) );
  AND2_X1 U340bar ( .A1(n630bar), .A2(n629bar), .ZN(n942bar) );
  OR2_X1 U341 ( .A1(n628), .A2(n627), .ZN(n629) );
  AND2_X1 U341bar ( .A1(n628bar), .A2(n627bar), .ZN(n629bar) );
  OR2_X1 U342 ( .A1(n626), .A2(n625), .ZN(n627) );
  AND2_X1 U342bar ( .A1(n626bar), .A2(n625bar), .ZN(n627bar) );
  OR2_X1 U343 ( .A1(in[146]), .A2(in[100]), .ZN(n625) );
  AND2_X1 U343bar ( .A1(inbar[146]), .A2(inbar[100]), .ZN(n625bar) );
  OR2_X1 U344 ( .A1(in[168]), .A2(in[152]), .ZN(n626) );
  AND2_X1 U344bar ( .A1(inbar[168]), .A2(inbar[152]), .ZN(n626bar) );
  OR2_X1 U345 ( .A1(n624), .A2(n623), .ZN(n628) );
  AND2_X1 U345bar ( .A1(n624bar), .A2(n623bar), .ZN(n628bar) );
  OR2_X1 U346 ( .A1(in[199]), .A2(in[182]), .ZN(n623) );
  AND2_X1 U346bar ( .A1(inbar[199]), .A2(inbar[182]), .ZN(n623bar) );
  OR2_X1 U347 ( .A1(in[236]), .A2(in[204]), .ZN(n624) );
  AND2_X1 U347bar ( .A1(inbar[236]), .A2(inbar[204]), .ZN(n624bar) );
  OR2_X1 U348 ( .A1(n622), .A2(n621), .ZN(n630) );
  AND2_X1 U348bar ( .A1(n622bar), .A2(n621bar), .ZN(n630bar) );
  OR2_X1 U349 ( .A1(n620), .A2(n619), .ZN(n621) );
  AND2_X1 U349bar ( .A1(n620bar), .A2(n619bar), .ZN(n621bar) );
  OR2_X1 U350 ( .A1(in[89]), .A2(in[246]), .ZN(n619) );
  AND2_X1 U350bar ( .A1(inbar[89]), .A2(inbar[246]), .ZN(n619bar) );
  OR2_X1 U351 ( .A1(in[95]), .A2(in[92]), .ZN(n620) );
  AND2_X1 U351bar ( .A1(inbar[95]), .A2(inbar[92]), .ZN(n620bar) );
  OR2_X1 U352 ( .A1(n618), .A2(n617), .ZN(n622) );
  AND2_X1 U352bar ( .A1(n618bar), .A2(n617bar), .ZN(n622bar) );
  OR2_X1 U353 ( .A1(in_22), .A2(in_16), .ZN(n617) );
  AND2_X1 U353bar ( .A1(in_22bar), .A2(in_16bar), .ZN(n617bar) );
  OR2_X1 U354 ( .A1(in_51), .A2(in_49), .ZN(n618) );
  AND2_X1 U354bar ( .A1(in_51bar), .A2(in_49bar), .ZN(n618bar) );
  OR2_X1 U355 ( .A1(n616), .A2(n615), .ZN(n722) );
  AND2_X1 U355bar ( .A1(n616bar), .A2(n615bar), .ZN(n722bar) );
  OR2_X1 U356 ( .A1(in[158]), .A2(in[115]), .ZN(n615) );
  AND2_X1 U356bar ( .A1(inbar[158]), .A2(inbar[115]), .ZN(n615bar) );
  OR2_X1 U357 ( .A1(in[163]), .A2(n614), .ZN(n616) );
  AND2_X1 U357bar ( .A1(inbar[163]), .A2(n614bar), .ZN(n616bar) );
  OR2_X1 U358 ( .A1(in[206]), .A2(in[165]), .ZN(n614) );
  AND2_X1 U358bar ( .A1(inbar[206]), .A2(inbar[165]), .ZN(n614bar) );
  OR2_X1 U359 ( .A1(n613), .A2(n612), .ZN(n724) );
  AND2_X1 U359bar ( .A1(n613bar), .A2(n612bar), .ZN(n724bar) );
  OR2_X1 U360 ( .A1(n611), .A2(n610), .ZN(n612) );
  AND2_X1 U360bar ( .A1(n611bar), .A2(n610bar), .ZN(n612bar) );
  OR2_X1 U361 ( .A1(in[213]), .A2(in[207]), .ZN(n610) );
  AND2_X1 U361bar ( .A1(inbar[213]), .A2(inbar[207]), .ZN(n610bar) );
  OR2_X1 U362 ( .A1(in[215]), .A2(n609), .ZN(n611) );
  AND2_X1 U362bar ( .A1(inbar[215]), .A2(n609bar), .ZN(n611bar) );
  OR2_X1 U363 ( .A1(in[230]), .A2(in[220]), .ZN(n609) );
  AND2_X1 U363bar ( .A1(inbar[230]), .A2(inbar[220]), .ZN(n609bar) );
  OR2_X1 U364 ( .A1(n608), .A2(n607), .ZN(n613) );
  AND2_X1 U364bar ( .A1(n608bar), .A2(n607bar), .ZN(n613bar) );
  OR2_X1 U365 ( .A1(in[251]), .A2(in[234]), .ZN(n607) );
  AND2_X1 U365bar ( .A1(inbar[251]), .A2(inbar[234]), .ZN(n607bar) );
  OR2_X1 U366 ( .A1(in_17), .A2(n606), .ZN(n608) );
  AND2_X1 U366bar ( .A1(in_17bar), .A2(n606bar), .ZN(n608bar) );
  OR2_X1 U367 ( .A1(in_65), .A2(in_56), .ZN(n606) );
  AND2_X1 U367bar ( .A1(in_65bar), .A2(in_56bar), .ZN(n606bar) );
  OR2_X1 U368 ( .A1(n605), .A2(n604), .ZN(out[0]) );
  AND2_X1 U368bar ( .A1(n605bar), .A2(n604bar), .ZN(outbar[0]) );
  OR2_X1 U369 ( .A1(n603), .A2(n602), .ZN(n604) );
  AND2_X1 U369bar ( .A1(n603bar), .A2(n602bar), .ZN(n604bar) );
  OR2_X1 U370 ( .A1(n601), .A2(n600), .ZN(n602) );
  AND2_X1 U370bar ( .A1(n601bar), .A2(n600bar), .ZN(n602bar) );
  OR2_X1 U371 ( .A1(n820), .A2(n785), .ZN(n600) );
  AND2_X1 U371bar ( .A1(n820bar), .A2(n785bar), .ZN(n600bar) );
  OR2_X1 U372 ( .A1(n599), .A2(n598), .ZN(n785) );
  AND2_X1 U372bar ( .A1(n599bar), .A2(n598bar), .ZN(n785bar) );
  OR2_X1 U373 ( .A1(n597), .A2(n596), .ZN(n598) );
  AND2_X1 U373bar ( .A1(n597bar), .A2(n596bar), .ZN(n598bar) );
  OR2_X1 U374 ( .A1(n595), .A2(n594), .ZN(n596) );
  AND2_X1 U374bar ( .A1(n595bar), .A2(n594bar), .ZN(n596bar) );
  OR2_X1 U375 ( .A1(in[135]), .A2(in[104]), .ZN(n594) );
  AND2_X1 U375bar ( .A1(inbar[135]), .A2(inbar[104]), .ZN(n594bar) );
  OR2_X1 U376 ( .A1(in[188]), .A2(in[178]), .ZN(n595) );
  AND2_X1 U376bar ( .A1(inbar[188]), .A2(inbar[178]), .ZN(n595bar) );
  OR2_X1 U377 ( .A1(n593), .A2(n592), .ZN(n597) );
  AND2_X1 U377bar ( .A1(n593bar), .A2(n592bar), .ZN(n597bar) );
  OR2_X1 U378 ( .A1(in[217]), .A2(in[194]), .ZN(n592) );
  AND2_X1 U378bar ( .A1(inbar[217]), .A2(inbar[194]), .ZN(n592bar) );
  OR2_X1 U379 ( .A1(in[237]), .A2(in[218]), .ZN(n593) );
  AND2_X1 U379bar ( .A1(inbar[237]), .A2(inbar[218]), .ZN(n593bar) );
  OR2_X1 U380 ( .A1(n591), .A2(n590), .ZN(n599) );
  AND2_X1 U380bar ( .A1(n591bar), .A2(n590bar), .ZN(n599bar) );
  OR2_X1 U381 ( .A1(n589), .A2(n588), .ZN(n590) );
  AND2_X1 U381bar ( .A1(n589bar), .A2(n588bar), .ZN(n590bar) );
  OR2_X1 U382 ( .A1(in_2), .A2(in_10), .ZN(n588) );
  AND2_X1 U382bar ( .A1(in_2bar), .A2(in_10bar), .ZN(n588bar) );
  OR2_X1 U383 ( .A1(in_47), .A2(in_22), .ZN(n589) );
  AND2_X1 U383bar ( .A1(in_47bar), .A2(in_22bar), .ZN(n589bar) );
  OR2_X1 U384 ( .A1(n587), .A2(n586), .ZN(n591) );
  AND2_X1 U384bar ( .A1(n587bar), .A2(n586bar), .ZN(n591bar) );
  OR2_X1 U385 ( .A1(in_56), .A2(in_54), .ZN(n586) );
  AND2_X1 U385bar ( .A1(in_56bar), .A2(in_54bar), .ZN(n586bar) );
  OR2_X1 U386 ( .A1(in_63), .A2(in_61), .ZN(n587) );
  AND2_X1 U386bar ( .A1(in_63bar), .A2(in_61bar), .ZN(n587bar) );
  OR2_X1 U387 ( .A1(n585), .A2(n584), .ZN(n820) );
  AND2_X1 U387bar ( .A1(n585bar), .A2(n584bar), .ZN(n820bar) );
  OR2_X1 U388 ( .A1(n583), .A2(n582), .ZN(n584) );
  AND2_X1 U388bar ( .A1(n583bar), .A2(n582bar), .ZN(n584bar) );
  OR2_X1 U389 ( .A1(n581), .A2(n580), .ZN(n582) );
  AND2_X1 U389bar ( .A1(n581bar), .A2(n580bar), .ZN(n582bar) );
  OR2_X1 U390 ( .A1(in[158]), .A2(in[142]), .ZN(n580) );
  AND2_X1 U390bar ( .A1(inbar[158]), .A2(inbar[142]), .ZN(n580bar) );
  OR2_X1 U391 ( .A1(in[175]), .A2(in[164]), .ZN(n581) );
  AND2_X1 U391bar ( .A1(inbar[175]), .A2(inbar[164]), .ZN(n581bar) );
  OR2_X1 U392 ( .A1(n579), .A2(n578), .ZN(n583) );
  AND2_X1 U392bar ( .A1(n579bar), .A2(n578bar), .ZN(n583bar) );
  OR2_X1 U393 ( .A1(in[228]), .A2(in[204]), .ZN(n578) );
  AND2_X1 U393bar ( .A1(inbar[228]), .A2(inbar[204]), .ZN(n578bar) );
  OR2_X1 U394 ( .A1(in[91]), .A2(in[87]), .ZN(n579) );
  AND2_X1 U394bar ( .A1(inbar[91]), .A2(inbar[87]), .ZN(n579bar) );
  OR2_X1 U395 ( .A1(n577), .A2(n576), .ZN(n585) );
  AND2_X1 U395bar ( .A1(n577bar), .A2(n576bar), .ZN(n585bar) );
  OR2_X1 U396 ( .A1(n575), .A2(n574), .ZN(n576) );
  AND2_X1 U396bar ( .A1(n575bar), .A2(n574bar), .ZN(n576bar) );
  OR2_X1 U397 ( .A1(in_21), .A2(in_11), .ZN(n574) );
  AND2_X1 U397bar ( .A1(in_21bar), .A2(in_11bar), .ZN(n574bar) );
  OR2_X1 U398 ( .A1(in_5), .A2(in_3), .ZN(n575) );
  AND2_X1 U398bar ( .A1(in_5bar), .A2(in_3bar), .ZN(n575bar) );
  OR2_X1 U399 ( .A1(n573), .A2(n572), .ZN(n577) );
  AND2_X1 U399bar ( .A1(n573bar), .A2(n572bar), .ZN(n577bar) );
  OR2_X1 U400 ( .A1(in_68), .A2(in_64), .ZN(n572) );
  AND2_X1 U400bar ( .A1(in_68bar), .A2(in_64bar), .ZN(n572bar) );
  OR2_X1 U401 ( .A1(in_76), .A2(in_73), .ZN(n573) );
  AND2_X1 U401bar ( .A1(in_76bar), .A2(in_73bar), .ZN(n573bar) );
  OR2_X1 U402 ( .A1(n778), .A2(n571), .ZN(n601) );
  AND2_X1 U402bar ( .A1(n778bar), .A2(n571bar), .ZN(n601bar) );
  OR2_X1 U403 ( .A1(in[100]), .A2(n965), .ZN(n571) );
  AND2_X1 U403bar ( .A1(inbar[100]), .A2(n965bar), .ZN(n571bar) );
  OR2_X1 U404 ( .A1(n570), .A2(n569), .ZN(n965) );
  AND2_X1 U404bar ( .A1(n570bar), .A2(n569bar), .ZN(n965bar) );
  OR2_X1 U405 ( .A1(n568), .A2(n567), .ZN(n569) );
  AND2_X1 U405bar ( .A1(n568bar), .A2(n567bar), .ZN(n569bar) );
  OR2_X1 U406 ( .A1(n566), .A2(n565), .ZN(n567) );
  AND2_X1 U406bar ( .A1(n566bar), .A2(n565bar), .ZN(n567bar) );
  OR2_X1 U407 ( .A1(n817), .A2(n750), .ZN(n565) );
  AND2_X1 U407bar ( .A1(n817bar), .A2(n750bar), .ZN(n565bar) );
  OR2_X1 U408 ( .A1(n564), .A2(n563), .ZN(n750) );
  AND2_X1 U408bar ( .A1(n564bar), .A2(n563bar), .ZN(n750bar) );
  OR2_X1 U409 ( .A1(n562), .A2(n561), .ZN(n563) );
  AND2_X1 U409bar ( .A1(n562bar), .A2(n561bar), .ZN(n563bar) );
  OR2_X1 U410 ( .A1(n560), .A2(n559), .ZN(n561) );
  AND2_X1 U410bar ( .A1(n560bar), .A2(n559bar), .ZN(n561bar) );
  OR2_X1 U411 ( .A1(in[119]), .A2(in[103]), .ZN(n559) );
  AND2_X1 U411bar ( .A1(inbar[119]), .A2(inbar[103]), .ZN(n559bar) );
  OR2_X1 U412 ( .A1(in[137]), .A2(in[133]), .ZN(n560) );
  AND2_X1 U412bar ( .A1(inbar[137]), .A2(inbar[133]), .ZN(n560bar) );
  OR2_X1 U413 ( .A1(n558), .A2(n557), .ZN(n562) );
  AND2_X1 U413bar ( .A1(n558bar), .A2(n557bar), .ZN(n562bar) );
  OR2_X1 U414 ( .A1(in[176]), .A2(in[173]), .ZN(n557) );
  AND2_X1 U414bar ( .A1(inbar[176]), .A2(inbar[173]), .ZN(n557bar) );
  OR2_X1 U415 ( .A1(in[210]), .A2(in[181]), .ZN(n558) );
  AND2_X1 U415bar ( .A1(inbar[210]), .A2(inbar[181]), .ZN(n558bar) );
  OR2_X1 U416 ( .A1(n556), .A2(n555), .ZN(n564) );
  AND2_X1 U416bar ( .A1(n556bar), .A2(n555bar), .ZN(n564bar) );
  OR2_X1 U417 ( .A1(n554), .A2(n553), .ZN(n555) );
  AND2_X1 U417bar ( .A1(n554bar), .A2(n553bar), .ZN(n555bar) );
  OR2_X1 U418 ( .A1(in_13), .A2(in[234]), .ZN(n553) );
  AND2_X1 U418bar ( .A1(in_13bar), .A2(inbar[234]), .ZN(n553bar) );
  OR2_X1 U419 ( .A1(in_38), .A2(in_32), .ZN(n554) );
  AND2_X1 U419bar ( .A1(in_38bar), .A2(in_32bar), .ZN(n554bar) );
  OR2_X1 U420 ( .A1(n552), .A2(n551), .ZN(n556) );
  AND2_X1 U420bar ( .A1(n552bar), .A2(n551bar), .ZN(n556bar) );
  OR2_X1 U421 ( .A1(in_42), .A2(in_41), .ZN(n551) );
  AND2_X1 U421bar ( .A1(in_42bar), .A2(in_41bar), .ZN(n551bar) );
  OR2_X1 U422 ( .A1(in_7), .A2(in_49), .ZN(n552) );
  AND2_X1 U422bar ( .A1(in_7bar), .A2(in_49bar), .ZN(n552bar) );
  OR2_X1 U423 ( .A1(n550), .A2(n549), .ZN(n817) );
  AND2_X1 U423bar ( .A1(n550bar), .A2(n549bar), .ZN(n817bar) );
  OR2_X1 U424 ( .A1(n548), .A2(n547), .ZN(n549) );
  AND2_X1 U424bar ( .A1(n548bar), .A2(n547bar), .ZN(n549bar) );
  OR2_X1 U425 ( .A1(n546), .A2(n545), .ZN(n547) );
  AND2_X1 U425bar ( .A1(n546bar), .A2(n545bar), .ZN(n547bar) );
  OR2_X1 U426 ( .A1(in[159]), .A2(in[105]), .ZN(n545) );
  AND2_X1 U426bar ( .A1(inbar[159]), .A2(inbar[105]), .ZN(n545bar) );
  OR2_X1 U427 ( .A1(in[206]), .A2(in[183]), .ZN(n546) );
  AND2_X1 U427bar ( .A1(inbar[206]), .A2(inbar[183]), .ZN(n546bar) );
  OR2_X1 U428 ( .A1(n544), .A2(n543), .ZN(n548) );
  AND2_X1 U428bar ( .A1(n544bar), .A2(n543bar), .ZN(n548bar) );
  OR2_X1 U429 ( .A1(in[229]), .A2(in[219]), .ZN(n543) );
  AND2_X1 U429bar ( .A1(inbar[229]), .A2(inbar[219]), .ZN(n543bar) );
  OR2_X1 U430 ( .A1(in[235]), .A2(in[232]), .ZN(n544) );
  AND2_X1 U430bar ( .A1(inbar[235]), .A2(inbar[232]), .ZN(n544bar) );
  OR2_X1 U431 ( .A1(n542), .A2(n541), .ZN(n550) );
  AND2_X1 U431bar ( .A1(n542bar), .A2(n541bar), .ZN(n550bar) );
  OR2_X1 U432 ( .A1(n540), .A2(n539), .ZN(n541) );
  AND2_X1 U432bar ( .A1(n540bar), .A2(n539bar), .ZN(n541bar) );
  OR2_X1 U433 ( .A1(in[249]), .A2(in[242]), .ZN(n539) );
  AND2_X1 U433bar ( .A1(inbar[249]), .A2(inbar[242]), .ZN(n539bar) );
  OR2_X1 U434 ( .A1(in[89]), .A2(in[254]), .ZN(n540) );
  AND2_X1 U434bar ( .A1(inbar[89]), .A2(inbar[254]), .ZN(n540bar) );
  OR2_X1 U435 ( .A1(n538), .A2(n537), .ZN(n542) );
  AND2_X1 U435bar ( .A1(n538bar), .A2(n537bar), .ZN(n542bar) );
  OR2_X1 U436 ( .A1(in_14), .A2(in[99]), .ZN(n537) );
  AND2_X1 U436bar ( .A1(in_14bar), .A2(inbar[99]), .ZN(n537bar) );
  OR2_X1 U437 ( .A1(in_60), .A2(in_18), .ZN(n538) );
  AND2_X1 U437bar ( .A1(in_60bar), .A2(in_18bar), .ZN(n538bar) );
  OR2_X1 U438 ( .A1(in[113]), .A2(n763), .ZN(n566) );
  AND2_X1 U438bar ( .A1(inbar[113]), .A2(n763bar), .ZN(n566bar) );
  OR2_X1 U439 ( .A1(n536), .A2(n535), .ZN(n763) );
  AND2_X1 U439bar ( .A1(n536bar), .A2(n535bar), .ZN(n763bar) );
  OR2_X1 U440 ( .A1(n534), .A2(n533), .ZN(n535) );
  AND2_X1 U440bar ( .A1(n534bar), .A2(n533bar), .ZN(n535bar) );
  OR2_X1 U441 ( .A1(n532), .A2(n531), .ZN(n533) );
  AND2_X1 U441bar ( .A1(n532bar), .A2(n531bar), .ZN(n533bar) );
  OR2_X1 U442 ( .A1(in[115]), .A2(in[110]), .ZN(n531) );
  AND2_X1 U442bar ( .A1(inbar[115]), .A2(inbar[110]), .ZN(n531bar) );
  OR2_X1 U443 ( .A1(in[125]), .A2(in[117]), .ZN(n532) );
  AND2_X1 U443bar ( .A1(inbar[125]), .A2(inbar[117]), .ZN(n532bar) );
  OR2_X1 U444 ( .A1(n530), .A2(n529), .ZN(n534) );
  AND2_X1 U444bar ( .A1(n530bar), .A2(n529bar), .ZN(n534bar) );
  OR2_X1 U445 ( .A1(in[180]), .A2(in[128]), .ZN(n529) );
  AND2_X1 U445bar ( .A1(inbar[180]), .A2(inbar[128]), .ZN(n529bar) );
  OR2_X1 U446 ( .A1(in[205]), .A2(in[201]), .ZN(n530) );
  AND2_X1 U446bar ( .A1(inbar[205]), .A2(inbar[201]), .ZN(n530bar) );
  OR2_X1 U447 ( .A1(n528), .A2(n527), .ZN(n536) );
  AND2_X1 U447bar ( .A1(n528bar), .A2(n527bar), .ZN(n536bar) );
  OR2_X1 U448 ( .A1(n526), .A2(n525), .ZN(n527) );
  AND2_X1 U448bar ( .A1(n526bar), .A2(n525bar), .ZN(n527bar) );
  OR2_X1 U449 ( .A1(in[244]), .A2(in[239]), .ZN(n525) );
  AND2_X1 U449bar ( .A1(inbar[244]), .A2(inbar[239]), .ZN(n525bar) );
  OR2_X1 U450 ( .A1(in[95]), .A2(in[83]), .ZN(n526) );
  AND2_X1 U450bar ( .A1(inbar[95]), .A2(inbar[83]), .ZN(n526bar) );
  OR2_X1 U451 ( .A1(n524), .A2(n523), .ZN(n528) );
  AND2_X1 U451bar ( .A1(n524bar), .A2(n523bar), .ZN(n528bar) );
  OR2_X1 U452 ( .A1(in_24), .A2(in[97]), .ZN(n523) );
  AND2_X1 U452bar ( .A1(in_24bar), .A2(inbar[97]), .ZN(n523bar) );
  OR2_X1 U453 ( .A1(in_33), .A2(in_27), .ZN(n524) );
  AND2_X1 U453bar ( .A1(in_33bar), .A2(in_27bar), .ZN(n524bar) );
  OR2_X1 U454 ( .A1(n522), .A2(n521), .ZN(n568) );
  AND2_X1 U454bar ( .A1(n522bar), .A2(n521bar), .ZN(n568bar) );
  OR2_X1 U455 ( .A1(in[145]), .A2(in[126]), .ZN(n521) );
  AND2_X1 U455bar ( .A1(inbar[145]), .A2(inbar[126]), .ZN(n521bar) );
  OR2_X1 U456 ( .A1(in[169]), .A2(n520), .ZN(n522) );
  AND2_X1 U456bar ( .A1(inbar[169]), .A2(n520bar), .ZN(n522bar) );
  OR2_X1 U457 ( .A1(in[221]), .A2(in[172]), .ZN(n520) );
  AND2_X1 U457bar ( .A1(inbar[221]), .A2(inbar[172]), .ZN(n520bar) );
  OR2_X1 U458 ( .A1(n519), .A2(n518), .ZN(n570) );
  AND2_X1 U458bar ( .A1(n519bar), .A2(n518bar), .ZN(n570bar) );
  OR2_X1 U459 ( .A1(n517), .A2(n516), .ZN(n518) );
  AND2_X1 U459bar ( .A1(n517bar), .A2(n516bar), .ZN(n518bar) );
  OR2_X1 U460 ( .A1(in[241]), .A2(in[224]), .ZN(n516) );
  AND2_X1 U460bar ( .A1(inbar[241]), .A2(inbar[224]), .ZN(n516bar) );
  OR2_X1 U461 ( .A1(in[86]), .A2(n515), .ZN(n517) );
  AND2_X1 U461bar ( .A1(inbar[86]), .A2(n515bar), .ZN(n517bar) );
  OR2_X1 U462 ( .A1(in_43), .A2(in_34), .ZN(n515) );
  AND2_X1 U462bar ( .A1(in_43bar), .A2(in_34bar), .ZN(n515bar) );
  OR2_X1 U463 ( .A1(n514), .A2(n513), .ZN(n519) );
  AND2_X1 U463bar ( .A1(n514bar), .A2(n513bar), .ZN(n519bar) );
  OR2_X1 U464 ( .A1(in_65), .A2(in_51), .ZN(n513) );
  AND2_X1 U464bar ( .A1(in_65bar), .A2(in_51bar), .ZN(n513bar) );
  OR2_X1 U465 ( .A1(in_75), .A2(n512), .ZN(n514) );
  AND2_X1 U465bar ( .A1(in_75bar), .A2(n512bar), .ZN(n514bar) );
  OR2_X1 U466 ( .A1(in_81), .A2(in_77), .ZN(n512) );
  AND2_X1 U466bar ( .A1(in_81bar), .A2(in_77bar), .ZN(n512bar) );
  OR2_X1 U467 ( .A1(n511), .A2(n510), .ZN(n778) );
  AND2_X1 U467bar ( .A1(n511bar), .A2(n510bar), .ZN(n778bar) );
  OR2_X1 U468 ( .A1(n509), .A2(n508), .ZN(n510) );
  AND2_X1 U468bar ( .A1(n509bar), .A2(n508bar), .ZN(n510bar) );
  OR2_X1 U469 ( .A1(n507), .A2(n506), .ZN(n508) );
  AND2_X1 U469bar ( .A1(n507bar), .A2(n506bar), .ZN(n508bar) );
  OR2_X1 U470 ( .A1(in[107]), .A2(in[101]), .ZN(n506) );
  AND2_X1 U470bar ( .A1(inbar[107]), .A2(inbar[101]), .ZN(n506bar) );
  OR2_X1 U471 ( .A1(in[139]), .A2(in[132]), .ZN(n507) );
  AND2_X1 U471bar ( .A1(inbar[139]), .A2(inbar[132]), .ZN(n507bar) );
  OR2_X1 U472 ( .A1(n505), .A2(n504), .ZN(n509) );
  AND2_X1 U472bar ( .A1(n505bar), .A2(n504bar), .ZN(n509bar) );
  OR2_X1 U473 ( .A1(in[146]), .A2(in[141]), .ZN(n504) );
  AND2_X1 U473bar ( .A1(inbar[146]), .A2(inbar[141]), .ZN(n504bar) );
  OR2_X1 U474 ( .A1(in[203]), .A2(in[179]), .ZN(n505) );
  AND2_X1 U474bar ( .A1(inbar[203]), .A2(inbar[179]), .ZN(n505bar) );
  OR2_X1 U475 ( .A1(n503), .A2(n502), .ZN(n511) );
  AND2_X1 U475bar ( .A1(n503bar), .A2(n502bar), .ZN(n511bar) );
  OR2_X1 U476 ( .A1(n501), .A2(n500), .ZN(n502) );
  AND2_X1 U476bar ( .A1(n501bar), .A2(n500bar), .ZN(n502bar) );
  OR2_X1 U477 ( .A1(in[243]), .A2(in[222]), .ZN(n500) );
  AND2_X1 U477bar ( .A1(inbar[243]), .A2(inbar[222]), .ZN(n500bar) );
  OR2_X1 U478 ( .A1(in[251]), .A2(in[250]), .ZN(n501) );
  AND2_X1 U478bar ( .A1(inbar[251]), .A2(inbar[250]), .ZN(n501bar) );
  OR2_X1 U479 ( .A1(n499), .A2(n498), .ZN(n503) );
  AND2_X1 U479bar ( .A1(n499bar), .A2(n498bar), .ZN(n503bar) );
  OR2_X1 U480 ( .A1(in_37), .A2(in_19), .ZN(n498) );
  AND2_X1 U480bar ( .A1(in_37bar), .A2(in_19bar), .ZN(n498bar) );
  OR2_X1 U481 ( .A1(in_78), .A2(in_6), .ZN(n499) );
  AND2_X1 U481bar ( .A1(in_78bar), .A2(in_6bar), .ZN(n499bar) );
  OR2_X1 U482 ( .A1(n497), .A2(n496), .ZN(n603) );
  AND2_X1 U482bar ( .A1(n497bar), .A2(n496bar), .ZN(n603bar) );
  OR2_X1 U483 ( .A1(in[112]), .A2(in[102]), .ZN(n496) );
  AND2_X1 U483bar ( .A1(inbar[112]), .A2(inbar[102]), .ZN(n496bar) );
  OR2_X1 U484 ( .A1(in[123]), .A2(n495), .ZN(n497) );
  AND2_X1 U484bar ( .A1(inbar[123]), .A2(n495bar), .ZN(n497bar) );
  OR2_X1 U485 ( .A1(in[143]), .A2(in[130]), .ZN(n495) );
  AND2_X1 U485bar ( .A1(inbar[143]), .A2(inbar[130]), .ZN(n495bar) );
  OR2_X1 U486 ( .A1(n494), .A2(n493), .ZN(n605) );
  AND2_X1 U486bar ( .A1(n494bar), .A2(n493bar), .ZN(n605bar) );
  OR2_X1 U487 ( .A1(n492), .A2(n491), .ZN(n493) );
  AND2_X1 U487bar ( .A1(n492bar), .A2(n491bar), .ZN(n493bar) );
  OR2_X1 U488 ( .A1(in[216]), .A2(in[213]), .ZN(n491) );
  AND2_X1 U488bar ( .A1(inbar[216]), .A2(inbar[213]), .ZN(n491bar) );
  OR2_X1 U489 ( .A1(in[227]), .A2(n490), .ZN(n492) );
  AND2_X1 U489bar ( .A1(inbar[227]), .A2(n490bar), .ZN(n492bar) );
  OR2_X1 U490 ( .A1(in_0), .A2(in[248]), .ZN(n490) );
  AND2_X1 U490bar ( .A1(in_0bar), .A2(inbar[248]), .ZN(n490bar) );
  OR2_X1 U491 ( .A1(n489), .A2(n488), .ZN(n494) );
  AND2_X1 U491bar ( .A1(n489bar), .A2(n488bar), .ZN(n494bar) );
  OR2_X1 U492 ( .A1(in_46), .A2(in_44), .ZN(n488) );
  AND2_X1 U492bar ( .A1(in_46bar), .A2(in_44bar), .ZN(n488bar) );
  OR2_X1 U493 ( .A1(in_50), .A2(n487), .ZN(n489) );
  AND2_X1 U493bar ( .A1(in_50bar), .A2(n487bar), .ZN(n489bar) );
  OR2_X1 U494 ( .A1(in_9), .A2(in_80), .ZN(n487) );
  AND2_X1 U494bar ( .A1(in_9bar), .A2(in_80bar), .ZN(n487bar) );
endmodule

module sBox_5 ( in, inbar, out, outbar );

  input wire [7:0] in;
  input wire [7:0] inbar;
//input_done

  output wire [7:0] out;
  output wire [7:0] outbar;
//output_done

  wire [255:0] decodeOut;
  wire [255:0] decodeOutbar;
//wire_done

  decode_5 dec ( .in(in), .inbar(inbar), .out(decodeOut), .outbar(decodeOutbar) );
  encode_5 enc ( .in(decodeOut), .inbar(decodeOutbar), .out(out), .outbar(outbar) );
endmodule

module CD2_21 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD2_22 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD2_23 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD2_24 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD4_11 ( a, abar, b, bbar, y, ybar );

  input wire [3:0] a;
  input wire [3:0] b;
  input wire [3:0] abar;
  input wire [3:0] bbar;
//input_done

  output wire [15:0] y;
  output wire [15:0] ybar;
//output_done

//wire_done

  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]) );
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]) );
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]) );
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]) );
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]) );
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]) );
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]) );
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]) );
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]) );
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]) );
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]) );
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]) );
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]) );
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]) );
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]) );
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]) );
endmodule

module CD4_12( a, abar, b, bbar, y, ybar );

  input wire [3:0] a;
  input wire [3:0] b;
  input wire [3:0] abar;
  input wire [3:0] bbar;
//input_done

  output wire [15:0] y;
  output wire [15:0] ybar;
//output_done

//wire_done

  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]) );
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]) );
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]) );
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]) );
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]) );
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]) );
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]) );
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]) );
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]) );
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]) );
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]) );
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]) );
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]) );
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]) );
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]) );
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]) );
endmodule

module CD16_6 ( a, abar, b, bbar, y, ybar );

  input wire [15:0] a;
  input wire [15:0] b;
  input wire [15:0] abar;
  input wire [15:0] bbar;
//input_done

  output wire [255:0] y;
  output wire [255:0] ybar;
//output_done

//wire_done

  AND2_X1 U1 ( .A1(b[9]), .A2(a[0]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[9]), .A2(abar[0]), .ZN(ybar[9]) );
  AND2_X1 U2 ( .A1(b[3]), .A2(a[6]), .ZN(y[99]) );
  OR2_X1 U2bar ( .A1(bbar[3]), .A2(abar[6]), .ZN(ybar[99]) );
  AND2_X1 U3 ( .A1(b[2]), .A2(a[6]), .ZN(y[98]) );
  OR2_X1 U3bar ( .A1(bbar[2]), .A2(abar[6]), .ZN(ybar[98]) );
  AND2_X1 U4 ( .A1(b[1]), .A2(a[6]), .ZN(y[97]) );
  OR2_X1 U4bar ( .A1(bbar[1]), .A2(abar[6]), .ZN(ybar[97]) );
  AND2_X1 U5 ( .A1(b[0]), .A2(a[6]), .ZN(y[96]) );
  OR2_X1 U5bar ( .A1(bbar[0]), .A2(abar[6]), .ZN(ybar[96]) );
  AND2_X1 U6 ( .A1(b[15]), .A2(a[5]), .ZN(y[95]) );
  OR2_X1 U6bar ( .A1(bbar[15]), .A2(abar[5]), .ZN(ybar[95]) );
  AND2_X1 U7 ( .A1(b[14]), .A2(a[5]), .ZN(y[94]) );
  OR2_X1 U7bar ( .A1(bbar[14]), .A2(abar[5]), .ZN(ybar[94]) );
  AND2_X1 U8 ( .A1(b[13]), .A2(a[5]), .ZN(y[93]) );
  OR2_X1 U8bar ( .A1(bbar[13]), .A2(abar[5]), .ZN(ybar[93]) );
  AND2_X1 U9 ( .A1(b[12]), .A2(a[5]), .ZN(y[92]) );
  OR2_X1 U9bar ( .A1(bbar[12]), .A2(abar[5]), .ZN(ybar[92]) );
  AND2_X1 U10 ( .A1(b[11]), .A2(a[5]), .ZN(y[91]) );
  OR2_X1 U10bar ( .A1(bbar[11]), .A2(abar[5]), .ZN(ybar[91]) );
  AND2_X1 U11 ( .A1(b[10]), .A2(a[5]), .ZN(y[90]) );
  OR2_X1 U11bar ( .A1(bbar[10]), .A2(abar[5]), .ZN(ybar[90]) );
  AND2_X1 U12 ( .A1(b[8]), .A2(a[0]), .ZN(y[8]) );
  OR2_X1 U12bar ( .A1(bbar[8]), .A2(abar[0]), .ZN(ybar[8]) );
  AND2_X1 U13 ( .A1(a[5]), .A2(b[9]), .ZN(y[89]) );
  OR2_X1 U13bar ( .A1(abar[5]), .A2(bbar[9]), .ZN(ybar[89]) );
  AND2_X1 U14 ( .A1(b[8]), .A2(a[5]), .ZN(y[88]) );
  OR2_X1 U14bar ( .A1(bbar[8]), .A2(abar[5]), .ZN(ybar[88]) );
  AND2_X1 U15 ( .A1(b[7]), .A2(a[5]), .ZN(y[87]) );
  OR2_X1 U15bar ( .A1(bbar[7]), .A2(abar[5]), .ZN(ybar[87]) );
  AND2_X1 U16 ( .A1(b[6]), .A2(a[5]), .ZN(y[86]) );
  OR2_X1 U16bar ( .A1(bbar[6]), .A2(abar[5]), .ZN(ybar[86]) );
  AND2_X1 U17 ( .A1(b[5]), .A2(a[5]), .ZN(y[85]) );
  OR2_X1 U17bar ( .A1(bbar[5]), .A2(abar[5]), .ZN(ybar[85]) );
  AND2_X1 U18 ( .A1(b[4]), .A2(a[5]), .ZN(y[84]) );
  OR2_X1 U18bar ( .A1(bbar[4]), .A2(abar[5]), .ZN(ybar[84]) );
  AND2_X1 U19 ( .A1(a[5]), .A2(b[3]), .ZN(y[83]) );
  OR2_X1 U19bar ( .A1(abar[5]), .A2(bbar[3]), .ZN(ybar[83]) );
  AND2_X1 U20 ( .A1(a[5]), .A2(b[2]), .ZN(y[82]) );
  OR2_X1 U20bar ( .A1(abar[5]), .A2(bbar[2]), .ZN(ybar[82]) );
  AND2_X1 U21 ( .A1(a[5]), .A2(b[1]), .ZN(y[81]) );
  OR2_X1 U21bar ( .A1(abar[5]), .A2(bbar[1]), .ZN(ybar[81]) );
  AND2_X1 U22 ( .A1(a[5]), .A2(b[0]), .ZN(y[80]) );
  OR2_X1 U22bar ( .A1(abar[5]), .A2(bbar[0]), .ZN(ybar[80]) );
  AND2_X1 U23 ( .A1(b[7]), .A2(a[0]), .ZN(y[7]) );
  OR2_X1 U23bar ( .A1(bbar[7]), .A2(abar[0]), .ZN(ybar[7]) );
  AND2_X1 U24 ( .A1(a[4]), .A2(b[15]), .ZN(y[79]) );
  OR2_X1 U24bar ( .A1(abar[4]), .A2(bbar[15]), .ZN(ybar[79]) );
  AND2_X1 U25 ( .A1(a[4]), .A2(b[14]), .ZN(y[78]) );
  OR2_X1 U25bar ( .A1(abar[4]), .A2(bbar[14]), .ZN(ybar[78]) );
  AND2_X1 U26 ( .A1(a[4]), .A2(b[13]), .ZN(y[77]) );
  OR2_X1 U26bar ( .A1(abar[4]), .A2(bbar[13]), .ZN(ybar[77]) );
  AND2_X1 U27 ( .A1(a[4]), .A2(b[12]), .ZN(y[76]) );
  OR2_X1 U27bar ( .A1(abar[4]), .A2(bbar[12]), .ZN(ybar[76]) );
  AND2_X1 U28 ( .A1(a[4]), .A2(b[11]), .ZN(y[75]) );
  OR2_X1 U28bar ( .A1(abar[4]), .A2(bbar[11]), .ZN(ybar[75]) );
  AND2_X1 U29 ( .A1(a[4]), .A2(b[10]), .ZN(y[74]) );
  OR2_X1 U29bar ( .A1(abar[4]), .A2(bbar[10]), .ZN(ybar[74]) );
  AND2_X1 U30 ( .A1(a[4]), .A2(b[9]), .ZN(y[73]) );
  OR2_X1 U30bar ( .A1(abar[4]), .A2(bbar[9]), .ZN(ybar[73]) );
  AND2_X1 U31 ( .A1(a[4]), .A2(b[8]), .ZN(y[72]) );
  OR2_X1 U31bar ( .A1(abar[4]), .A2(bbar[8]), .ZN(ybar[72]) );
  AND2_X1 U32 ( .A1(a[4]), .A2(b[7]), .ZN(y[71]) );
  OR2_X1 U32bar ( .A1(abar[4]), .A2(bbar[7]), .ZN(ybar[71]) );
  AND2_X1 U33 ( .A1(a[4]), .A2(b[6]), .ZN(y[70]) );
  OR2_X1 U33bar ( .A1(abar[4]), .A2(bbar[6]), .ZN(ybar[70]) );
  AND2_X1 U34 ( .A1(b[6]), .A2(a[0]), .ZN(y[6]) );
  OR2_X1 U34bar ( .A1(bbar[6]), .A2(abar[0]), .ZN(ybar[6]) );
  AND2_X1 U35 ( .A1(a[4]), .A2(b[5]), .ZN(y[69]) );
  OR2_X1 U35bar ( .A1(abar[4]), .A2(bbar[5]), .ZN(ybar[69]) );
  AND2_X1 U36 ( .A1(a[4]), .A2(b[4]), .ZN(y[68]) );
  OR2_X1 U36bar ( .A1(abar[4]), .A2(bbar[4]), .ZN(ybar[68]) );
  AND2_X1 U37 ( .A1(a[4]), .A2(b[3]), .ZN(y[67]) );
  OR2_X1 U37bar ( .A1(abar[4]), .A2(bbar[3]), .ZN(ybar[67]) );
  AND2_X1 U38 ( .A1(a[4]), .A2(b[2]), .ZN(y[66]) );
  OR2_X1 U38bar ( .A1(abar[4]), .A2(bbar[2]), .ZN(ybar[66]) );
  AND2_X1 U39 ( .A1(a[4]), .A2(b[1]), .ZN(y[65]) );
  OR2_X1 U39bar ( .A1(abar[4]), .A2(bbar[1]), .ZN(ybar[65]) );
  AND2_X1 U40 ( .A1(a[4]), .A2(b[0]), .ZN(y[64]) );
  OR2_X1 U40bar ( .A1(abar[4]), .A2(bbar[0]), .ZN(ybar[64]) );
  AND2_X1 U41 ( .A1(a[3]), .A2(b[15]), .ZN(y[63]) );
  OR2_X1 U41bar ( .A1(abar[3]), .A2(bbar[15]), .ZN(ybar[63]) );
  AND2_X1 U42 ( .A1(a[3]), .A2(b[14]), .ZN(y[62]) );
  OR2_X1 U42bar ( .A1(abar[3]), .A2(bbar[14]), .ZN(ybar[62]) );
  AND2_X1 U43 ( .A1(a[3]), .A2(b[13]), .ZN(y[61]) );
  OR2_X1 U43bar ( .A1(abar[3]), .A2(bbar[13]), .ZN(ybar[61]) );
  AND2_X1 U44 ( .A1(a[3]), .A2(b[12]), .ZN(y[60]) );
  OR2_X1 U44bar ( .A1(abar[3]), .A2(bbar[12]), .ZN(ybar[60]) );
  AND2_X1 U45 ( .A1(b[5]), .A2(a[0]), .ZN(y[5]) );
  OR2_X1 U45bar ( .A1(bbar[5]), .A2(abar[0]), .ZN(ybar[5]) );
  AND2_X1 U46 ( .A1(a[3]), .A2(b[11]), .ZN(y[59]) );
  OR2_X1 U46bar ( .A1(abar[3]), .A2(bbar[11]), .ZN(ybar[59]) );
  AND2_X1 U47 ( .A1(a[3]), .A2(b[10]), .ZN(y[58]) );
  OR2_X1 U47bar ( .A1(abar[3]), .A2(bbar[10]), .ZN(ybar[58]) );
  AND2_X1 U48 ( .A1(a[3]), .A2(b[9]), .ZN(y[57]) );
  OR2_X1 U48bar ( .A1(abar[3]), .A2(bbar[9]), .ZN(ybar[57]) );
  AND2_X1 U49 ( .A1(a[3]), .A2(b[8]), .ZN(y[56]) );
  OR2_X1 U49bar ( .A1(abar[3]), .A2(bbar[8]), .ZN(ybar[56]) );
  AND2_X1 U50 ( .A1(a[3]), .A2(b[7]), .ZN(y[55]) );
  OR2_X1 U50bar ( .A1(abar[3]), .A2(bbar[7]), .ZN(ybar[55]) );
  AND2_X1 U51 ( .A1(a[3]), .A2(b[6]), .ZN(y[54]) );
  OR2_X1 U51bar ( .A1(abar[3]), .A2(bbar[6]), .ZN(ybar[54]) );
  AND2_X1 U52 ( .A1(a[3]), .A2(b[5]), .ZN(y[53]) );
  OR2_X1 U52bar ( .A1(abar[3]), .A2(bbar[5]), .ZN(ybar[53]) );
  AND2_X1 U53 ( .A1(a[3]), .A2(b[4]), .ZN(y[52]) );
  OR2_X1 U53bar ( .A1(abar[3]), .A2(bbar[4]), .ZN(ybar[52]) );
  AND2_X1 U54 ( .A1(a[3]), .A2(b[3]), .ZN(y[51]) );
  OR2_X1 U54bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[51]) );
  AND2_X1 U55 ( .A1(a[3]), .A2(b[2]), .ZN(y[50]) );
  OR2_X1 U55bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[50]) );
  AND2_X1 U56 ( .A1(b[4]), .A2(a[0]), .ZN(y[4]) );
  OR2_X1 U56bar ( .A1(bbar[4]), .A2(abar[0]), .ZN(ybar[4]) );
  AND2_X1 U57 ( .A1(a[3]), .A2(b[1]), .ZN(y[49]) );
  OR2_X1 U57bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[49]) );
  AND2_X1 U58 ( .A1(a[3]), .A2(b[0]), .ZN(y[48]) );
  OR2_X1 U58bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[48]) );
  AND2_X1 U59 ( .A1(a[2]), .A2(b[15]), .ZN(y[47]) );
  OR2_X1 U59bar ( .A1(abar[2]), .A2(bbar[15]), .ZN(ybar[47]) );
  AND2_X1 U60 ( .A1(a[2]), .A2(b[14]), .ZN(y[46]) );
  OR2_X1 U60bar ( .A1(abar[2]), .A2(bbar[14]), .ZN(ybar[46]) );
  AND2_X1 U61 ( .A1(a[2]), .A2(b[13]), .ZN(y[45]) );
  OR2_X1 U61bar ( .A1(abar[2]), .A2(bbar[13]), .ZN(ybar[45]) );
  AND2_X1 U62 ( .A1(a[2]), .A2(b[12]), .ZN(y[44]) );
  OR2_X1 U62bar ( .A1(abar[2]), .A2(bbar[12]), .ZN(ybar[44]) );
  AND2_X1 U63 ( .A1(a[2]), .A2(b[11]), .ZN(y[43]) );
  OR2_X1 U63bar ( .A1(abar[2]), .A2(bbar[11]), .ZN(ybar[43]) );
  AND2_X1 U64 ( .A1(a[2]), .A2(b[10]), .ZN(y[42]) );
  OR2_X1 U64bar ( .A1(abar[2]), .A2(bbar[10]), .ZN(ybar[42]) );
  AND2_X1 U65 ( .A1(a[2]), .A2(b[9]), .ZN(y[41]) );
  OR2_X1 U65bar ( .A1(abar[2]), .A2(bbar[9]), .ZN(ybar[41]) );
  AND2_X1 U66 ( .A1(a[2]), .A2(b[8]), .ZN(y[40]) );
  OR2_X1 U66bar ( .A1(abar[2]), .A2(bbar[8]), .ZN(ybar[40]) );
  AND2_X1 U67 ( .A1(b[3]), .A2(a[0]), .ZN(y[3]) );
  OR2_X1 U67bar ( .A1(bbar[3]), .A2(abar[0]), .ZN(ybar[3]) );
  AND2_X1 U68 ( .A1(a[2]), .A2(b[7]), .ZN(y[39]) );
  OR2_X1 U68bar ( .A1(abar[2]), .A2(bbar[7]), .ZN(ybar[39]) );
  AND2_X1 U69 ( .A1(a[2]), .A2(b[6]), .ZN(y[38]) );
  OR2_X1 U69bar ( .A1(abar[2]), .A2(bbar[6]), .ZN(ybar[38]) );
  AND2_X1 U70 ( .A1(a[2]), .A2(b[5]), .ZN(y[37]) );
  OR2_X1 U70bar ( .A1(abar[2]), .A2(bbar[5]), .ZN(ybar[37]) );
  AND2_X1 U71 ( .A1(a[2]), .A2(b[4]), .ZN(y[36]) );
  OR2_X1 U71bar ( .A1(abar[2]), .A2(bbar[4]), .ZN(ybar[36]) );
  AND2_X1 U72 ( .A1(a[2]), .A2(b[3]), .ZN(y[35]) );
  OR2_X1 U72bar ( .A1(abar[2]), .A2(bbar[3]), .ZN(ybar[35]) );
  AND2_X1 U73 ( .A1(a[2]), .A2(b[2]), .ZN(y[34]) );
  OR2_X1 U73bar ( .A1(abar[2]), .A2(bbar[2]), .ZN(ybar[34]) );
  AND2_X1 U74 ( .A1(a[2]), .A2(b[1]), .ZN(y[33]) );
  OR2_X1 U74bar ( .A1(abar[2]), .A2(bbar[1]), .ZN(ybar[33]) );
  AND2_X1 U75 ( .A1(a[2]), .A2(b[0]), .ZN(y[32]) );
  OR2_X1 U75bar ( .A1(abar[2]), .A2(bbar[0]), .ZN(ybar[32]) );
  AND2_X1 U76 ( .A1(a[1]), .A2(b[15]), .ZN(y[31]) );
  OR2_X1 U76bar ( .A1(abar[1]), .A2(bbar[15]), .ZN(ybar[31]) );
  AND2_X1 U77 ( .A1(a[1]), .A2(b[14]), .ZN(y[30]) );
  OR2_X1 U77bar ( .A1(abar[1]), .A2(bbar[14]), .ZN(ybar[30]) );
  AND2_X1 U78 ( .A1(b[2]), .A2(a[0]), .ZN(y[2]) );
  OR2_X1 U78bar ( .A1(bbar[2]), .A2(abar[0]), .ZN(ybar[2]) );
  AND2_X1 U79 ( .A1(a[1]), .A2(b[13]), .ZN(y[29]) );
  OR2_X1 U79bar ( .A1(abar[1]), .A2(bbar[13]), .ZN(ybar[29]) );
  AND2_X1 U80 ( .A1(a[1]), .A2(b[12]), .ZN(y[28]) );
  OR2_X1 U80bar ( .A1(abar[1]), .A2(bbar[12]), .ZN(ybar[28]) );
  AND2_X1 U81 ( .A1(a[1]), .A2(b[11]), .ZN(y[27]) );
  OR2_X1 U81bar ( .A1(abar[1]), .A2(bbar[11]), .ZN(ybar[27]) );
  AND2_X1 U82 ( .A1(a[1]), .A2(b[10]), .ZN(y[26]) );
  OR2_X1 U82bar ( .A1(abar[1]), .A2(bbar[10]), .ZN(ybar[26]) );
  AND2_X1 U83 ( .A1(a[1]), .A2(b[9]), .ZN(y[25]) );
  OR2_X1 U83bar ( .A1(abar[1]), .A2(bbar[9]), .ZN(ybar[25]) );
  AND2_X1 U84 ( .A1(a[15]), .A2(b[15]), .ZN(y[255]) );
  OR2_X1 U84bar ( .A1(abar[15]), .A2(bbar[15]), .ZN(ybar[255]) );
  AND2_X1 U85 ( .A1(a[15]), .A2(b[14]), .ZN(y[254]) );
  OR2_X1 U85bar ( .A1(abar[15]), .A2(bbar[14]), .ZN(ybar[254]) );
  AND2_X1 U86 ( .A1(a[15]), .A2(b[13]), .ZN(y[253]) );
  OR2_X1 U86bar ( .A1(abar[15]), .A2(bbar[13]), .ZN(ybar[253]) );
  AND2_X1 U87 ( .A1(a[15]), .A2(b[12]), .ZN(y[252]) );
  OR2_X1 U87bar ( .A1(abar[15]), .A2(bbar[12]), .ZN(ybar[252]) );
  AND2_X1 U88 ( .A1(a[15]), .A2(b[11]), .ZN(y[251]) );
  OR2_X1 U88bar ( .A1(abar[15]), .A2(bbar[11]), .ZN(ybar[251]) );
  AND2_X1 U89 ( .A1(a[15]), .A2(b[10]), .ZN(y[250]) );
  OR2_X1 U89bar ( .A1(abar[15]), .A2(bbar[10]), .ZN(ybar[250]) );
  AND2_X1 U90 ( .A1(a[1]), .A2(b[8]), .ZN(y[24]) );
  OR2_X1 U90bar ( .A1(abar[1]), .A2(bbar[8]), .ZN(ybar[24]) );
  AND2_X1 U91 ( .A1(a[15]), .A2(b[9]), .ZN(y[249]) );
  OR2_X1 U91bar ( .A1(abar[15]), .A2(bbar[9]), .ZN(ybar[249]) );
  AND2_X1 U92 ( .A1(a[15]), .A2(b[8]), .ZN(y[248]) );
  OR2_X1 U92bar ( .A1(abar[15]), .A2(bbar[8]), .ZN(ybar[248]) );
  AND2_X1 U93 ( .A1(a[15]), .A2(b[7]), .ZN(y[247]) );
  OR2_X1 U93bar ( .A1(abar[15]), .A2(bbar[7]), .ZN(ybar[247]) );
  AND2_X1 U94 ( .A1(a[15]), .A2(b[6]), .ZN(y[246]) );
  OR2_X1 U94bar ( .A1(abar[15]), .A2(bbar[6]), .ZN(ybar[246]) );
  AND2_X1 U95 ( .A1(a[15]), .A2(b[5]), .ZN(y[245]) );
  OR2_X1 U95bar ( .A1(abar[15]), .A2(bbar[5]), .ZN(ybar[245]) );
  AND2_X1 U96 ( .A1(a[15]), .A2(b[4]), .ZN(y[244]) );
  OR2_X1 U96bar ( .A1(abar[15]), .A2(bbar[4]), .ZN(ybar[244]) );
  AND2_X1 U97 ( .A1(a[15]), .A2(b[3]), .ZN(y[243]) );
  OR2_X1 U97bar ( .A1(abar[15]), .A2(bbar[3]), .ZN(ybar[243]) );
  AND2_X1 U98 ( .A1(a[15]), .A2(b[2]), .ZN(y[242]) );
  OR2_X1 U98bar ( .A1(abar[15]), .A2(bbar[2]), .ZN(ybar[242]) );
  AND2_X1 U99 ( .A1(a[15]), .A2(b[1]), .ZN(y[241]) );
  OR2_X1 U99bar ( .A1(abar[15]), .A2(bbar[1]), .ZN(ybar[241]) );
  AND2_X1 U100 ( .A1(a[15]), .A2(b[0]), .ZN(y[240]) );
  OR2_X1 U100bar ( .A1(abar[15]), .A2(bbar[0]), .ZN(ybar[240]) );
  AND2_X1 U101 ( .A1(a[1]), .A2(b[7]), .ZN(y[23]) );
  OR2_X1 U101bar ( .A1(abar[1]), .A2(bbar[7]), .ZN(ybar[23]) );
  AND2_X1 U102 ( .A1(a[14]), .A2(b[15]), .ZN(y[239]) );
  OR2_X1 U102bar ( .A1(abar[14]), .A2(bbar[15]), .ZN(ybar[239]) );
  AND2_X1 U103 ( .A1(a[14]), .A2(b[14]), .ZN(y[238]) );
  OR2_X1 U103bar ( .A1(abar[14]), .A2(bbar[14]), .ZN(ybar[238]) );
  AND2_X1 U104 ( .A1(a[14]), .A2(b[13]), .ZN(y[237]) );
  OR2_X1 U104bar ( .A1(abar[14]), .A2(bbar[13]), .ZN(ybar[237]) );
  AND2_X1 U105 ( .A1(a[14]), .A2(b[12]), .ZN(y[236]) );
  OR2_X1 U105bar ( .A1(abar[14]), .A2(bbar[12]), .ZN(ybar[236]) );
  AND2_X1 U106 ( .A1(a[14]), .A2(b[11]), .ZN(y[235]) );
  OR2_X1 U106bar ( .A1(abar[14]), .A2(bbar[11]), .ZN(ybar[235]) );
  AND2_X1 U107 ( .A1(a[14]), .A2(b[10]), .ZN(y[234]) );
  OR2_X1 U107bar ( .A1(abar[14]), .A2(bbar[10]), .ZN(ybar[234]) );
  AND2_X1 U108 ( .A1(a[14]), .A2(b[9]), .ZN(y[233]) );
  OR2_X1 U108bar ( .A1(abar[14]), .A2(bbar[9]), .ZN(ybar[233]) );
  AND2_X1 U109 ( .A1(a[14]), .A2(b[8]), .ZN(y[232]) );
  OR2_X1 U109bar ( .A1(abar[14]), .A2(bbar[8]), .ZN(ybar[232]) );
  AND2_X1 U110 ( .A1(a[14]), .A2(b[7]), .ZN(y[231]) );
  OR2_X1 U110bar ( .A1(abar[14]), .A2(bbar[7]), .ZN(ybar[231]) );
  AND2_X1 U111 ( .A1(a[14]), .A2(b[6]), .ZN(y[230]) );
  OR2_X1 U111bar ( .A1(abar[14]), .A2(bbar[6]), .ZN(ybar[230]) );
  AND2_X1 U112 ( .A1(a[1]), .A2(b[6]), .ZN(y[22]) );
  OR2_X1 U112bar ( .A1(abar[1]), .A2(bbar[6]), .ZN(ybar[22]) );
  AND2_X1 U113 ( .A1(a[14]), .A2(b[5]), .ZN(y[229]) );
  OR2_X1 U113bar ( .A1(abar[14]), .A2(bbar[5]), .ZN(ybar[229]) );
  AND2_X1 U114 ( .A1(a[14]), .A2(b[4]), .ZN(y[228]) );
  OR2_X1 U114bar ( .A1(abar[14]), .A2(bbar[4]), .ZN(ybar[228]) );
  AND2_X1 U115 ( .A1(a[14]), .A2(b[3]), .ZN(y[227]) );
  OR2_X1 U115bar ( .A1(abar[14]), .A2(bbar[3]), .ZN(ybar[227]) );
  AND2_X1 U116 ( .A1(a[14]), .A2(b[2]), .ZN(y[226]) );
  OR2_X1 U116bar ( .A1(abar[14]), .A2(bbar[2]), .ZN(ybar[226]) );
  AND2_X1 U117 ( .A1(a[14]), .A2(b[1]), .ZN(y[225]) );
  OR2_X1 U117bar ( .A1(abar[14]), .A2(bbar[1]), .ZN(ybar[225]) );
  AND2_X1 U118 ( .A1(a[14]), .A2(b[0]), .ZN(y[224]) );
  OR2_X1 U118bar ( .A1(abar[14]), .A2(bbar[0]), .ZN(ybar[224]) );
  AND2_X1 U119 ( .A1(a[13]), .A2(b[15]), .ZN(y[223]) );
  OR2_X1 U119bar ( .A1(abar[13]), .A2(bbar[15]), .ZN(ybar[223]) );
  AND2_X1 U120 ( .A1(a[13]), .A2(b[14]), .ZN(y[222]) );
  OR2_X1 U120bar ( .A1(abar[13]), .A2(bbar[14]), .ZN(ybar[222]) );
  AND2_X1 U121 ( .A1(a[13]), .A2(b[13]), .ZN(y[221]) );
  OR2_X1 U121bar ( .A1(abar[13]), .A2(bbar[13]), .ZN(ybar[221]) );
  AND2_X1 U122 ( .A1(a[13]), .A2(b[12]), .ZN(y[220]) );
  OR2_X1 U122bar ( .A1(abar[13]), .A2(bbar[12]), .ZN(ybar[220]) );
  AND2_X1 U123 ( .A1(a[1]), .A2(b[5]), .ZN(y[21]) );
  OR2_X1 U123bar ( .A1(abar[1]), .A2(bbar[5]), .ZN(ybar[21]) );
  AND2_X1 U124 ( .A1(a[13]), .A2(b[11]), .ZN(y[219]) );
  OR2_X1 U124bar ( .A1(abar[13]), .A2(bbar[11]), .ZN(ybar[219]) );
  AND2_X1 U125 ( .A1(a[13]), .A2(b[10]), .ZN(y[218]) );
  OR2_X1 U125bar ( .A1(abar[13]), .A2(bbar[10]), .ZN(ybar[218]) );
  AND2_X1 U126 ( .A1(a[13]), .A2(b[9]), .ZN(y[217]) );
  OR2_X1 U126bar ( .A1(abar[13]), .A2(bbar[9]), .ZN(ybar[217]) );
  AND2_X1 U127 ( .A1(a[13]), .A2(b[8]), .ZN(y[216]) );
  OR2_X1 U127bar ( .A1(abar[13]), .A2(bbar[8]), .ZN(ybar[216]) );
  AND2_X1 U128 ( .A1(a[13]), .A2(b[7]), .ZN(y[215]) );
  OR2_X1 U128bar ( .A1(abar[13]), .A2(bbar[7]), .ZN(ybar[215]) );
  AND2_X1 U129 ( .A1(a[13]), .A2(b[6]), .ZN(y[214]) );
  OR2_X1 U129bar ( .A1(abar[13]), .A2(bbar[6]), .ZN(ybar[214]) );
  AND2_X1 U130 ( .A1(a[13]), .A2(b[5]), .ZN(y[213]) );
  OR2_X1 U130bar ( .A1(abar[13]), .A2(bbar[5]), .ZN(ybar[213]) );
  AND2_X1 U131 ( .A1(a[13]), .A2(b[4]), .ZN(y[212]) );
  OR2_X1 U131bar ( .A1(abar[13]), .A2(bbar[4]), .ZN(ybar[212]) );
  AND2_X1 U132 ( .A1(a[13]), .A2(b[3]), .ZN(y[211]) );
  OR2_X1 U132bar ( .A1(abar[13]), .A2(bbar[3]), .ZN(ybar[211]) );
  AND2_X1 U133 ( .A1(a[13]), .A2(b[2]), .ZN(y[210]) );
  OR2_X1 U133bar ( .A1(abar[13]), .A2(bbar[2]), .ZN(ybar[210]) );
  AND2_X1 U134 ( .A1(a[1]), .A2(b[4]), .ZN(y[20]) );
  OR2_X1 U134bar ( .A1(abar[1]), .A2(bbar[4]), .ZN(ybar[20]) );
  AND2_X1 U135 ( .A1(a[13]), .A2(b[1]), .ZN(y[209]) );
  OR2_X1 U135bar ( .A1(abar[13]), .A2(bbar[1]), .ZN(ybar[209]) );
  AND2_X1 U136 ( .A1(a[13]), .A2(b[0]), .ZN(y[208]) );
  OR2_X1 U136bar ( .A1(abar[13]), .A2(bbar[0]), .ZN(ybar[208]) );
  AND2_X1 U137 ( .A1(a[12]), .A2(b[15]), .ZN(y[207]) );
  OR2_X1 U137bar ( .A1(abar[12]), .A2(bbar[15]), .ZN(ybar[207]) );
  AND2_X1 U138 ( .A1(a[12]), .A2(b[14]), .ZN(y[206]) );
  OR2_X1 U138bar ( .A1(abar[12]), .A2(bbar[14]), .ZN(ybar[206]) );
  AND2_X1 U139 ( .A1(a[12]), .A2(b[13]), .ZN(y[205]) );
  OR2_X1 U139bar ( .A1(abar[12]), .A2(bbar[13]), .ZN(ybar[205]) );
  AND2_X1 U140 ( .A1(a[12]), .A2(b[12]), .ZN(y[204]) );
  OR2_X1 U140bar ( .A1(abar[12]), .A2(bbar[12]), .ZN(ybar[204]) );
  AND2_X1 U141 ( .A1(a[12]), .A2(b[11]), .ZN(y[203]) );
  OR2_X1 U141bar ( .A1(abar[12]), .A2(bbar[11]), .ZN(ybar[203]) );
  AND2_X1 U142 ( .A1(a[12]), .A2(b[10]), .ZN(y[202]) );
  OR2_X1 U142bar ( .A1(abar[12]), .A2(bbar[10]), .ZN(ybar[202]) );
  AND2_X1 U143 ( .A1(a[12]), .A2(b[9]), .ZN(y[201]) );
  OR2_X1 U143bar ( .A1(abar[12]), .A2(bbar[9]), .ZN(ybar[201]) );
  AND2_X1 U144 ( .A1(a[12]), .A2(b[8]), .ZN(y[200]) );
  OR2_X1 U144bar ( .A1(abar[12]), .A2(bbar[8]), .ZN(ybar[200]) );
  AND2_X1 U145 ( .A1(b[1]), .A2(a[0]), .ZN(y[1]) );
  OR2_X1 U145bar ( .A1(bbar[1]), .A2(abar[0]), .ZN(ybar[1]) );
  AND2_X1 U146 ( .A1(a[1]), .A2(b[3]), .ZN(y[19]) );
  OR2_X1 U146bar ( .A1(abar[1]), .A2(bbar[3]), .ZN(ybar[19]) );
  AND2_X1 U147 ( .A1(a[12]), .A2(b[7]), .ZN(y[199]) );
  OR2_X1 U147bar ( .A1(abar[12]), .A2(bbar[7]), .ZN(ybar[199]) );
  AND2_X1 U148 ( .A1(a[12]), .A2(b[6]), .ZN(y[198]) );
  OR2_X1 U148bar ( .A1(abar[12]), .A2(bbar[6]), .ZN(ybar[198]) );
  AND2_X1 U149 ( .A1(a[12]), .A2(b[5]), .ZN(y[197]) );
  OR2_X1 U149bar ( .A1(abar[12]), .A2(bbar[5]), .ZN(ybar[197]) );
  AND2_X1 U150 ( .A1(a[12]), .A2(b[4]), .ZN(y[196]) );
  OR2_X1 U150bar ( .A1(abar[12]), .A2(bbar[4]), .ZN(ybar[196]) );
  AND2_X1 U151 ( .A1(a[12]), .A2(b[3]), .ZN(y[195]) );
  OR2_X1 U151bar ( .A1(abar[12]), .A2(bbar[3]), .ZN(ybar[195]) );
  AND2_X1 U152 ( .A1(a[12]), .A2(b[2]), .ZN(y[194]) );
  OR2_X1 U152bar ( .A1(abar[12]), .A2(bbar[2]), .ZN(ybar[194]) );
  AND2_X1 U153 ( .A1(a[12]), .A2(b[1]), .ZN(y[193]) );
  OR2_X1 U153bar ( .A1(abar[12]), .A2(bbar[1]), .ZN(ybar[193]) );
  AND2_X1 U154 ( .A1(a[12]), .A2(b[0]), .ZN(y[192]) );
  OR2_X1 U154bar ( .A1(abar[12]), .A2(bbar[0]), .ZN(ybar[192]) );
  AND2_X1 U155 ( .A1(a[11]), .A2(b[15]), .ZN(y[191]) );
  OR2_X1 U155bar ( .A1(abar[11]), .A2(bbar[15]), .ZN(ybar[191]) );
  AND2_X1 U156 ( .A1(a[11]), .A2(b[14]), .ZN(y[190]) );
  OR2_X1 U156bar ( .A1(abar[11]), .A2(bbar[14]), .ZN(ybar[190]) );
  AND2_X1 U157 ( .A1(a[1]), .A2(b[2]), .ZN(y[18]) );
  OR2_X1 U157bar ( .A1(abar[1]), .A2(bbar[2]), .ZN(ybar[18]) );
  AND2_X1 U158 ( .A1(a[11]), .A2(b[13]), .ZN(y[189]) );
  OR2_X1 U158bar ( .A1(abar[11]), .A2(bbar[13]), .ZN(ybar[189]) );
  AND2_X1 U159 ( .A1(a[11]), .A2(b[12]), .ZN(y[188]) );
  OR2_X1 U159bar ( .A1(abar[11]), .A2(bbar[12]), .ZN(ybar[188]) );
  AND2_X1 U160 ( .A1(a[11]), .A2(b[11]), .ZN(y[187]) );
  OR2_X1 U160bar ( .A1(abar[11]), .A2(bbar[11]), .ZN(ybar[187]) );
  AND2_X1 U161 ( .A1(a[11]), .A2(b[10]), .ZN(y[186]) );
  OR2_X1 U161bar ( .A1(abar[11]), .A2(bbar[10]), .ZN(ybar[186]) );
  AND2_X1 U162 ( .A1(a[11]), .A2(b[9]), .ZN(y[185]) );
  OR2_X1 U162bar ( .A1(abar[11]), .A2(bbar[9]), .ZN(ybar[185]) );
  AND2_X1 U163 ( .A1(a[11]), .A2(b[8]), .ZN(y[184]) );
  OR2_X1 U163bar ( .A1(abar[11]), .A2(bbar[8]), .ZN(ybar[184]) );
  AND2_X1 U164 ( .A1(a[11]), .A2(b[7]), .ZN(y[183]) );
  OR2_X1 U164bar ( .A1(abar[11]), .A2(bbar[7]), .ZN(ybar[183]) );
  AND2_X1 U165 ( .A1(a[11]), .A2(b[6]), .ZN(y[182]) );
  OR2_X1 U165bar ( .A1(abar[11]), .A2(bbar[6]), .ZN(ybar[182]) );
  AND2_X1 U166 ( .A1(a[11]), .A2(b[5]), .ZN(y[181]) );
  OR2_X1 U166bar ( .A1(abar[11]), .A2(bbar[5]), .ZN(ybar[181]) );
  AND2_X1 U167 ( .A1(a[11]), .A2(b[4]), .ZN(y[180]) );
  OR2_X1 U167bar ( .A1(abar[11]), .A2(bbar[4]), .ZN(ybar[180]) );
  AND2_X1 U168 ( .A1(a[1]), .A2(b[1]), .ZN(y[17]) );
  OR2_X1 U168bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[17]) );
  AND2_X1 U169 ( .A1(a[11]), .A2(b[3]), .ZN(y[179]) );
  OR2_X1 U169bar ( .A1(abar[11]), .A2(bbar[3]), .ZN(ybar[179]) );
  AND2_X1 U170 ( .A1(a[11]), .A2(b[2]), .ZN(y[178]) );
  OR2_X1 U170bar ( .A1(abar[11]), .A2(bbar[2]), .ZN(ybar[178]) );
  AND2_X1 U171 ( .A1(a[11]), .A2(b[1]), .ZN(y[177]) );
  OR2_X1 U171bar ( .A1(abar[11]), .A2(bbar[1]), .ZN(ybar[177]) );
  AND2_X1 U172 ( .A1(a[11]), .A2(b[0]), .ZN(y[176]) );
  OR2_X1 U172bar ( .A1(abar[11]), .A2(bbar[0]), .ZN(ybar[176]) );
  AND2_X1 U173 ( .A1(a[10]), .A2(b[15]), .ZN(y[175]) );
  OR2_X1 U173bar ( .A1(abar[10]), .A2(bbar[15]), .ZN(ybar[175]) );
  AND2_X1 U174 ( .A1(a[10]), .A2(b[14]), .ZN(y[174]) );
  OR2_X1 U174bar ( .A1(abar[10]), .A2(bbar[14]), .ZN(ybar[174]) );
  AND2_X1 U175 ( .A1(a[10]), .A2(b[13]), .ZN(y[173]) );
  OR2_X1 U175bar ( .A1(abar[10]), .A2(bbar[13]), .ZN(ybar[173]) );
  AND2_X1 U176 ( .A1(a[10]), .A2(b[12]), .ZN(y[172]) );
  OR2_X1 U176bar ( .A1(abar[10]), .A2(bbar[12]), .ZN(ybar[172]) );
  AND2_X1 U177 ( .A1(a[10]), .A2(b[11]), .ZN(y[171]) );
  OR2_X1 U177bar ( .A1(abar[10]), .A2(bbar[11]), .ZN(ybar[171]) );
  AND2_X1 U178 ( .A1(a[10]), .A2(b[10]), .ZN(y[170]) );
  OR2_X1 U178bar ( .A1(abar[10]), .A2(bbar[10]), .ZN(ybar[170]) );
  AND2_X1 U179 ( .A1(a[1]), .A2(b[0]), .ZN(y[16]) );
  OR2_X1 U179bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[16]) );
  AND2_X1 U180 ( .A1(a[10]), .A2(b[9]), .ZN(y[169]) );
  OR2_X1 U180bar ( .A1(abar[10]), .A2(bbar[9]), .ZN(ybar[169]) );
  AND2_X1 U181 ( .A1(a[10]), .A2(b[8]), .ZN(y[168]) );
  OR2_X1 U181bar ( .A1(abar[10]), .A2(bbar[8]), .ZN(ybar[168]) );
  AND2_X1 U182 ( .A1(a[10]), .A2(b[7]), .ZN(y[167]) );
  OR2_X1 U182bar ( .A1(abar[10]), .A2(bbar[7]), .ZN(ybar[167]) );
  AND2_X1 U183 ( .A1(a[10]), .A2(b[6]), .ZN(y[166]) );
  OR2_X1 U183bar ( .A1(abar[10]), .A2(bbar[6]), .ZN(ybar[166]) );
  AND2_X1 U184 ( .A1(a[10]), .A2(b[5]), .ZN(y[165]) );
  OR2_X1 U184bar ( .A1(abar[10]), .A2(bbar[5]), .ZN(ybar[165]) );
  AND2_X1 U185 ( .A1(a[10]), .A2(b[4]), .ZN(y[164]) );
  OR2_X1 U185bar ( .A1(abar[10]), .A2(bbar[4]), .ZN(ybar[164]) );
  AND2_X1 U186 ( .A1(a[10]), .A2(b[3]), .ZN(y[163]) );
  OR2_X1 U186bar ( .A1(abar[10]), .A2(bbar[3]), .ZN(ybar[163]) );
  AND2_X1 U187 ( .A1(a[10]), .A2(b[2]), .ZN(y[162]) );
  OR2_X1 U187bar ( .A1(abar[10]), .A2(bbar[2]), .ZN(ybar[162]) );
  AND2_X1 U188 ( .A1(a[10]), .A2(b[1]), .ZN(y[161]) );
  OR2_X1 U188bar ( .A1(abar[10]), .A2(bbar[1]), .ZN(ybar[161]) );
  AND2_X1 U189 ( .A1(a[10]), .A2(b[0]), .ZN(y[160]) );
  OR2_X1 U189bar ( .A1(abar[10]), .A2(bbar[0]), .ZN(ybar[160]) );
  AND2_X1 U190 ( .A1(b[15]), .A2(a[0]), .ZN(y[15]) );
  OR2_X1 U190bar ( .A1(bbar[15]), .A2(abar[0]), .ZN(ybar[15]) );
  AND2_X1 U191 ( .A1(a[9]), .A2(b[15]), .ZN(y[159]) );
  OR2_X1 U191bar ( .A1(abar[9]), .A2(bbar[15]), .ZN(ybar[159]) );
  AND2_X1 U192 ( .A1(a[9]), .A2(b[14]), .ZN(y[158]) );
  OR2_X1 U192bar ( .A1(abar[9]), .A2(bbar[14]), .ZN(ybar[158]) );
  AND2_X1 U193 ( .A1(a[9]), .A2(b[13]), .ZN(y[157]) );
  OR2_X1 U193bar ( .A1(abar[9]), .A2(bbar[13]), .ZN(ybar[157]) );
  AND2_X1 U194 ( .A1(a[9]), .A2(b[12]), .ZN(y[156]) );
  OR2_X1 U194bar ( .A1(abar[9]), .A2(bbar[12]), .ZN(ybar[156]) );
  AND2_X1 U195 ( .A1(a[9]), .A2(b[11]), .ZN(y[155]) );
  OR2_X1 U195bar ( .A1(abar[9]), .A2(bbar[11]), .ZN(ybar[155]) );
  AND2_X1 U196 ( .A1(a[9]), .A2(b[10]), .ZN(y[154]) );
  OR2_X1 U196bar ( .A1(abar[9]), .A2(bbar[10]), .ZN(ybar[154]) );
  AND2_X1 U197 ( .A1(a[9]), .A2(b[9]), .ZN(y[153]) );
  OR2_X1 U197bar ( .A1(abar[9]), .A2(bbar[9]), .ZN(ybar[153]) );
  AND2_X1 U198 ( .A1(a[9]), .A2(b[8]), .ZN(y[152]) );
  OR2_X1 U198bar ( .A1(abar[9]), .A2(bbar[8]), .ZN(ybar[152]) );
  AND2_X1 U199 ( .A1(a[9]), .A2(b[7]), .ZN(y[151]) );
  OR2_X1 U199bar ( .A1(abar[9]), .A2(bbar[7]), .ZN(ybar[151]) );
  AND2_X1 U200 ( .A1(a[9]), .A2(b[6]), .ZN(y[150]) );
  OR2_X1 U200bar ( .A1(abar[9]), .A2(bbar[6]), .ZN(ybar[150]) );
  AND2_X1 U201 ( .A1(b[14]), .A2(a[0]), .ZN(y[14]) );
  OR2_X1 U201bar ( .A1(bbar[14]), .A2(abar[0]), .ZN(ybar[14]) );
  AND2_X1 U202 ( .A1(a[9]), .A2(b[5]), .ZN(y[149]) );
  OR2_X1 U202bar ( .A1(abar[9]), .A2(bbar[5]), .ZN(ybar[149]) );
  AND2_X1 U203 ( .A1(a[9]), .A2(b[4]), .ZN(y[148]) );
  OR2_X1 U203bar ( .A1(abar[9]), .A2(bbar[4]), .ZN(ybar[148]) );
  AND2_X1 U204 ( .A1(a[9]), .A2(b[3]), .ZN(y[147]) );
  OR2_X1 U204bar ( .A1(abar[9]), .A2(bbar[3]), .ZN(ybar[147]) );
  AND2_X1 U205 ( .A1(a[9]), .A2(b[2]), .ZN(y[146]) );
  OR2_X1 U205bar ( .A1(abar[9]), .A2(bbar[2]), .ZN(ybar[146]) );
  AND2_X1 U206 ( .A1(a[9]), .A2(b[1]), .ZN(y[145]) );
  OR2_X1 U206bar ( .A1(abar[9]), .A2(bbar[1]), .ZN(ybar[145]) );
  AND2_X1 U207 ( .A1(a[9]), .A2(b[0]), .ZN(y[144]) );
  OR2_X1 U207bar ( .A1(abar[9]), .A2(bbar[0]), .ZN(ybar[144]) );
  AND2_X1 U208 ( .A1(a[8]), .A2(b[15]), .ZN(y[143]) );
  OR2_X1 U208bar ( .A1(abar[8]), .A2(bbar[15]), .ZN(ybar[143]) );
  AND2_X1 U209 ( .A1(a[8]), .A2(b[14]), .ZN(y[142]) );
  OR2_X1 U209bar ( .A1(abar[8]), .A2(bbar[14]), .ZN(ybar[142]) );
  AND2_X1 U210 ( .A1(a[8]), .A2(b[13]), .ZN(y[141]) );
  OR2_X1 U210bar ( .A1(abar[8]), .A2(bbar[13]), .ZN(ybar[141]) );
  AND2_X1 U211 ( .A1(a[8]), .A2(b[12]), .ZN(y[140]) );
  OR2_X1 U211bar ( .A1(abar[8]), .A2(bbar[12]), .ZN(ybar[140]) );
  AND2_X1 U212 ( .A1(b[13]), .A2(a[0]), .ZN(y[13]) );
  OR2_X1 U212bar ( .A1(bbar[13]), .A2(abar[0]), .ZN(ybar[13]) );
  AND2_X1 U213 ( .A1(a[8]), .A2(b[11]), .ZN(y[139]) );
  OR2_X1 U213bar ( .A1(abar[8]), .A2(bbar[11]), .ZN(ybar[139]) );
  AND2_X1 U214 ( .A1(a[8]), .A2(b[10]), .ZN(y[138]) );
  OR2_X1 U214bar ( .A1(abar[8]), .A2(bbar[10]), .ZN(ybar[138]) );
  AND2_X1 U215 ( .A1(a[8]), .A2(b[9]), .ZN(y[137]) );
  OR2_X1 U215bar ( .A1(abar[8]), .A2(bbar[9]), .ZN(ybar[137]) );
  AND2_X1 U216 ( .A1(a[8]), .A2(b[8]), .ZN(y[136]) );
  OR2_X1 U216bar ( .A1(abar[8]), .A2(bbar[8]), .ZN(ybar[136]) );
  AND2_X1 U217 ( .A1(a[8]), .A2(b[7]), .ZN(y[135]) );
  OR2_X1 U217bar ( .A1(abar[8]), .A2(bbar[7]), .ZN(ybar[135]) );
  AND2_X1 U218 ( .A1(a[8]), .A2(b[6]), .ZN(y[134]) );
  OR2_X1 U218bar ( .A1(abar[8]), .A2(bbar[6]), .ZN(ybar[134]) );
  AND2_X1 U219 ( .A1(a[8]), .A2(b[5]), .ZN(y[133]) );
  OR2_X1 U219bar ( .A1(abar[8]), .A2(bbar[5]), .ZN(ybar[133]) );
  AND2_X1 U220 ( .A1(a[8]), .A2(b[4]), .ZN(y[132]) );
  OR2_X1 U220bar ( .A1(abar[8]), .A2(bbar[4]), .ZN(ybar[132]) );
  AND2_X1 U221 ( .A1(a[8]), .A2(b[3]), .ZN(y[131]) );
  OR2_X1 U221bar ( .A1(abar[8]), .A2(bbar[3]), .ZN(ybar[131]) );
  AND2_X1 U222 ( .A1(a[8]), .A2(b[2]), .ZN(y[130]) );
  OR2_X1 U222bar ( .A1(abar[8]), .A2(bbar[2]), .ZN(ybar[130]) );
  AND2_X1 U223 ( .A1(b[12]), .A2(a[0]), .ZN(y[12]) );
  OR2_X1 U223bar ( .A1(bbar[12]), .A2(abar[0]), .ZN(ybar[12]) );
  AND2_X1 U224 ( .A1(a[8]), .A2(b[1]), .ZN(y[129]) );
  OR2_X1 U224bar ( .A1(abar[8]), .A2(bbar[1]), .ZN(ybar[129]) );
  AND2_X1 U225 ( .A1(a[8]), .A2(b[0]), .ZN(y[128]) );
  OR2_X1 U225bar ( .A1(abar[8]), .A2(bbar[0]), .ZN(ybar[128]) );
  AND2_X1 U226 ( .A1(a[7]), .A2(b[15]), .ZN(y[127]) );
  OR2_X1 U226bar ( .A1(abar[7]), .A2(bbar[15]), .ZN(ybar[127]) );
  AND2_X1 U227 ( .A1(a[7]), .A2(b[14]), .ZN(y[126]) );
  OR2_X1 U227bar ( .A1(abar[7]), .A2(bbar[14]), .ZN(ybar[126]) );
  AND2_X1 U228 ( .A1(a[7]), .A2(b[13]), .ZN(y[125]) );
  OR2_X1 U228bar ( .A1(abar[7]), .A2(bbar[13]), .ZN(ybar[125]) );
  AND2_X1 U229 ( .A1(a[7]), .A2(b[12]), .ZN(y[124]) );
  OR2_X1 U229bar ( .A1(abar[7]), .A2(bbar[12]), .ZN(ybar[124]) );
  AND2_X1 U230 ( .A1(a[7]), .A2(b[11]), .ZN(y[123]) );
  OR2_X1 U230bar ( .A1(abar[7]), .A2(bbar[11]), .ZN(ybar[123]) );
  AND2_X1 U231 ( .A1(a[7]), .A2(b[10]), .ZN(y[122]) );
  OR2_X1 U231bar ( .A1(abar[7]), .A2(bbar[10]), .ZN(ybar[122]) );
  AND2_X1 U232 ( .A1(a[7]), .A2(b[9]), .ZN(y[121]) );
  OR2_X1 U232bar ( .A1(abar[7]), .A2(bbar[9]), .ZN(ybar[121]) );
  AND2_X1 U233 ( .A1(a[7]), .A2(b[8]), .ZN(y[120]) );
  OR2_X1 U233bar ( .A1(abar[7]), .A2(bbar[8]), .ZN(ybar[120]) );
  AND2_X1 U234 ( .A1(b[11]), .A2(a[0]), .ZN(y[11]) );
  OR2_X1 U234bar ( .A1(bbar[11]), .A2(abar[0]), .ZN(ybar[11]) );
  AND2_X1 U235 ( .A1(a[7]), .A2(b[7]), .ZN(y[119]) );
  OR2_X1 U235bar ( .A1(abar[7]), .A2(bbar[7]), .ZN(ybar[119]) );
  AND2_X1 U236 ( .A1(a[7]), .A2(b[6]), .ZN(y[118]) );
  OR2_X1 U236bar ( .A1(abar[7]), .A2(bbar[6]), .ZN(ybar[118]) );
  AND2_X1 U237 ( .A1(a[7]), .A2(b[5]), .ZN(y[117]) );
  OR2_X1 U237bar ( .A1(abar[7]), .A2(bbar[5]), .ZN(ybar[117]) );
  AND2_X1 U238 ( .A1(a[7]), .A2(b[4]), .ZN(y[116]) );
  OR2_X1 U238bar ( .A1(abar[7]), .A2(bbar[4]), .ZN(ybar[116]) );
  AND2_X1 U239 ( .A1(a[7]), .A2(b[3]), .ZN(y[115]) );
  OR2_X1 U239bar ( .A1(abar[7]), .A2(bbar[3]), .ZN(ybar[115]) );
  AND2_X1 U240 ( .A1(a[7]), .A2(b[2]), .ZN(y[114]) );
  OR2_X1 U240bar ( .A1(abar[7]), .A2(bbar[2]), .ZN(ybar[114]) );
  AND2_X1 U241 ( .A1(a[7]), .A2(b[1]), .ZN(y[113]) );
  OR2_X1 U241bar ( .A1(abar[7]), .A2(bbar[1]), .ZN(ybar[113]) );
  AND2_X1 U242 ( .A1(a[7]), .A2(b[0]), .ZN(y[112]) );
  OR2_X1 U242bar ( .A1(abar[7]), .A2(bbar[0]), .ZN(ybar[112]) );
  AND2_X1 U243 ( .A1(b[15]), .A2(a[6]), .ZN(y[111]) );
  OR2_X1 U243bar ( .A1(bbar[15]), .A2(abar[6]), .ZN(ybar[111]) );
  AND2_X1 U244 ( .A1(b[14]), .A2(a[6]), .ZN(y[110]) );
  OR2_X1 U244bar ( .A1(bbar[14]), .A2(abar[6]), .ZN(ybar[110]) );
  AND2_X1 U245 ( .A1(b[10]), .A2(a[0]), .ZN(y[10]) );
  OR2_X1 U245bar ( .A1(bbar[10]), .A2(abar[0]), .ZN(ybar[10]) );
  AND2_X1 U246 ( .A1(b[13]), .A2(a[6]), .ZN(y[109]) );
  OR2_X1 U246bar ( .A1(bbar[13]), .A2(abar[6]), .ZN(ybar[109]) );
  AND2_X1 U247 ( .A1(b[12]), .A2(a[6]), .ZN(y[108]) );
  OR2_X1 U247bar ( .A1(bbar[12]), .A2(abar[6]), .ZN(ybar[108]) );
  AND2_X1 U248 ( .A1(b[11]), .A2(a[6]), .ZN(y[107]) );
  OR2_X1 U248bar ( .A1(bbar[11]), .A2(abar[6]), .ZN(ybar[107]) );
  AND2_X1 U249 ( .A1(b[10]), .A2(a[6]), .ZN(y[106]) );
  OR2_X1 U249bar ( .A1(bbar[10]), .A2(abar[6]), .ZN(ybar[106]) );
  AND2_X1 U250 ( .A1(a[6]), .A2(b[9]), .ZN(y[105]) );
  OR2_X1 U250bar ( .A1(abar[6]), .A2(bbar[9]), .ZN(ybar[105]) );
  AND2_X1 U251 ( .A1(b[8]), .A2(a[6]), .ZN(y[104]) );
  OR2_X1 U251bar ( .A1(bbar[8]), .A2(abar[6]), .ZN(ybar[104]) );
  AND2_X1 U252 ( .A1(b[7]), .A2(a[6]), .ZN(y[103]) );
  OR2_X1 U252bar ( .A1(bbar[7]), .A2(abar[6]), .ZN(ybar[103]) );
  AND2_X1 U253 ( .A1(b[6]), .A2(a[6]), .ZN(y[102]) );
  OR2_X1 U253bar ( .A1(bbar[6]), .A2(abar[6]), .ZN(ybar[102]) );
  AND2_X1 U254 ( .A1(b[5]), .A2(a[6]), .ZN(y[101]) );
  OR2_X1 U254bar ( .A1(bbar[5]), .A2(abar[6]), .ZN(ybar[101]) );
  AND2_X1 U255 ( .A1(b[4]), .A2(a[6]), .ZN(y[100]) );
  OR2_X1 U255bar ( .A1(bbar[4]), .A2(abar[6]), .ZN(ybar[100]) );
  AND2_X1 U256 ( .A1(b[0]), .A2(a[0]), .ZN(y[0]) );
  OR2_X1 U256bar ( .A1(bbar[0]), .A2(abar[0]), .ZN(ybar[0]) );
endmodule

module decode_6 ( in, inbar, out, outbar );

  input wire [7:0] in;
  input wire [7:0] inbar;
//input_done

  output wire [255:0] out;
  output wire [255:0] outbar;
//output_done

  wire [15:0] level1;
  wire [31:0] level2;
  wire [15:0] level1bar;
  wire [31:0] level2bar;
//wire_done

  CD2_24 cd_l1_1 ( .a(in[1]), .abar(inbar[1]), .b(in[0]), .bbar(inbar[0]), .y(level1[3:0]), .ybar(level1bar[3:0]) );
  CD2_23 cd_l1_2 ( .a(in[3]), .abar(inbar[3]), .b(in[2]), .bbar(inbar[2]), .y(level1[7:4]), .ybar(level1bar[7:4]) );
  CD2_22 cd_l1_3 ( .a(in[5]), .abar(inbar[5]), .b(in[4]), .bbar(inbar[4]), .y(level1[11:8]), .ybar(level1bar[11:8]) );
  CD2_21 cd_l1_4 ( .a(in[7]), .abar(inbar[7]), .b(in[6]), .bbar(inbar[6]), .y(level1[15:12]), .ybar(level1bar[15:12]) );

  CD4_12 cd_l2_1 ( .a(level1[7:4]), .abar(level1bar[7:4]), .b(level1[3:0]), .bbar(level1bar[3:0]), 
        .y(level2[15:0]), .ybar(level2bar[15:0]) );
  CD4_11 cd_l2_2 ( .a(level1[15:12]), .abar(level1bar[15:12]), .b(level1[11:8]), .bbar(level1bar[11:8]), 
        .y(level2[31:16]), .ybar(level2bar[31:16]) );
  CD16_6 cd_l3 ( .a(level2[31:16]), .abar(level2bar[31:16]), .b(level2[15:0]), .bbar(level2bar[15:0]), 
        .y(out), .ybar(outbar) );
endmodule

module encode_6 ( in, inbar, out, outbar );

  input wire [255:0] in;
  input wire [255:0] inbar;
//input_done

  output wire [7:0] out;
  output wire [7:0] outbar;
//output_done

  wire in_81;
  wire in_80;
  wire in_79;
  wire in_78;
  wire in_77;
  wire in_76;
  wire in_75;
  wire in_74;
  wire in_73;
  wire in_72;
  wire in_71;
  wire in_70;
  wire in_69;
  wire in_68;
  wire in_67;
  wire in_66;
  wire in_65;
  wire in_64;
  wire in_63;
  wire in_62;
  wire in_61;
  wire in_60;
  wire in_59;
  wire in_58;
  wire in_57;
  wire in_56;
  wire in_55;
  wire in_54;
  wire in_53;
  wire in_52;
  wire in_51;
  wire in_50;
  wire in_49;
  wire in_48;
  wire in_47;
  wire in_46;
  wire in_45;
  wire in_44;
  wire in_43;
  wire in_42;
  wire in_41;
  wire in_40;
  wire in_39;
  wire in_38;
  wire in_37;
  wire in_36;
  wire in_35;
  wire in_34;
  wire in_33;
  wire in_32;
  wire in_31;
  wire in_30;
  wire in_29;
  wire in_28;
  wire in_27;
  wire in_26;
  wire in_25;
  wire in_24;
  wire in_23;
  wire in_22;
  wire in_21;
  wire in_20;
  wire in_19;
  wire in_18;
  wire in_17;
  wire in_16;
  wire in_15;
  wire in_14;
  wire in_13;
  wire in_12;
  wire in_11;
  wire in_10;
  wire in_9;
  wire in_8;
  wire in_7;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_3;
  wire in_2;
  wire in_1;
  wire in_0;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire in_81bar;
  wire in_80bar;
  wire in_79bar;
  wire in_78bar;
  wire in_77bar;
  wire in_76bar;
  wire in_75bar;
  wire in_74bar;
  wire in_73bar;
  wire in_72bar;
  wire in_71bar;
  wire in_70bar;
  wire in_69bar;
  wire in_68bar;
  wire in_67bar;
  wire in_66bar;
  wire in_65bar;
  wire in_64bar;
  wire in_63bar;
  wire in_62bar;
  wire in_61bar;
  wire in_60bar;
  wire in_59bar;
  wire in_58bar;
  wire in_57bar;
  wire in_56bar;
  wire in_55bar;
  wire in_54bar;
  wire in_53bar;
  wire in_52bar;
  wire in_51bar;
  wire in_50bar;
  wire in_49bar;
  wire in_48bar;
  wire in_47bar;
  wire in_46bar;
  wire in_45bar;
  wire in_44bar;
  wire in_43bar;
  wire in_42bar;
  wire in_41bar;
  wire in_40bar;
  wire in_39bar;
  wire in_38bar;
  wire in_37bar;
  wire in_36bar;
  wire in_35bar;
  wire in_34bar;
  wire in_33bar;
  wire in_32bar;
  wire in_31bar;
  wire in_30bar;
  wire in_29bar;
  wire in_28bar;
  wire in_27bar;
  wire in_26bar;
  wire in_25bar;
  wire in_24bar;
  wire in_23bar;
  wire in_22bar;
  wire in_21bar;
  wire in_20bar;
  wire in_19bar;
  wire in_18bar;
  wire in_17bar;
  wire in_16bar;
  wire in_15bar;
  wire in_14bar;
  wire in_13bar;
  wire in_12bar;
  wire in_11bar;
  wire in_10bar;
  wire in_9bar;
  wire in_8bar;
  wire in_7bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_3bar;
  wire in_2bar;
  wire in_1bar;
  wire in_0bar;
  wire n487bar;
  wire n488bar;
  wire n489bar;
  wire n490bar;
  wire n491bar;
  wire n492bar;
  wire n493bar;
  wire n494bar;
  wire n495bar;
  wire n496bar;
  wire n497bar;
  wire n498bar;
  wire n499bar;
  wire n500bar;
  wire n501bar;
  wire n502bar;
  wire n503bar;
  wire n504bar;
  wire n505bar;
  wire n506bar;
  wire n507bar;
  wire n508bar;
  wire n509bar;
  wire n510bar;
  wire n511bar;
  wire n512bar;
  wire n513bar;
  wire n514bar;
  wire n515bar;
  wire n516bar;
  wire n517bar;
  wire n518bar;
  wire n519bar;
  wire n520bar;
  wire n521bar;
  wire n522bar;
  wire n523bar;
  wire n524bar;
  wire n525bar;
  wire n526bar;
  wire n527bar;
  wire n528bar;
  wire n529bar;
  wire n530bar;
  wire n531bar;
  wire n532bar;
  wire n533bar;
  wire n534bar;
  wire n535bar;
  wire n536bar;
  wire n537bar;
  wire n538bar;
  wire n539bar;
  wire n540bar;
  wire n541bar;
  wire n542bar;
  wire n543bar;
  wire n544bar;
  wire n545bar;
  wire n546bar;
  wire n547bar;
  wire n548bar;
  wire n549bar;
  wire n550bar;
  wire n551bar;
  wire n552bar;
  wire n553bar;
  wire n554bar;
  wire n555bar;
  wire n556bar;
  wire n557bar;
  wire n558bar;
  wire n559bar;
  wire n560bar;
  wire n561bar;
  wire n562bar;
  wire n563bar;
  wire n564bar;
  wire n565bar;
  wire n566bar;
  wire n567bar;
  wire n568bar;
  wire n569bar;
  wire n570bar;
  wire n571bar;
  wire n572bar;
  wire n573bar;
  wire n574bar;
  wire n575bar;
  wire n576bar;
  wire n577bar;
  wire n578bar;
  wire n579bar;
  wire n580bar;
  wire n581bar;
  wire n582bar;
  wire n583bar;
  wire n584bar;
  wire n585bar;
  wire n586bar;
  wire n587bar;
  wire n588bar;
  wire n589bar;
  wire n590bar;
  wire n591bar;
  wire n592bar;
  wire n593bar;
  wire n594bar;
  wire n595bar;
  wire n596bar;
  wire n597bar;
  wire n598bar;
  wire n599bar;
  wire n600bar;
  wire n601bar;
  wire n602bar;
  wire n603bar;
  wire n604bar;
  wire n605bar;
  wire n606bar;
  wire n607bar;
  wire n608bar;
  wire n609bar;
  wire n610bar;
  wire n611bar;
  wire n612bar;
  wire n613bar;
  wire n614bar;
  wire n615bar;
  wire n616bar;
  wire n617bar;
  wire n618bar;
  wire n619bar;
  wire n620bar;
  wire n621bar;
  wire n622bar;
  wire n623bar;
  wire n624bar;
  wire n625bar;
  wire n626bar;
  wire n627bar;
  wire n628bar;
  wire n629bar;
  wire n630bar;
  wire n631bar;
  wire n632bar;
  wire n633bar;
  wire n634bar;
  wire n635bar;
  wire n636bar;
  wire n637bar;
  wire n638bar;
  wire n639bar;
  wire n640bar;
  wire n641bar;
  wire n642bar;
  wire n643bar;
  wire n644bar;
  wire n645bar;
  wire n646bar;
  wire n647bar;
  wire n648bar;
  wire n649bar;
  wire n650bar;
  wire n651bar;
  wire n652bar;
  wire n653bar;
  wire n654bar;
  wire n655bar;
  wire n656bar;
  wire n657bar;
  wire n658bar;
  wire n659bar;
  wire n660bar;
  wire n661bar;
  wire n662bar;
  wire n663bar;
  wire n664bar;
  wire n665bar;
  wire n666bar;
  wire n667bar;
  wire n668bar;
  wire n669bar;
  wire n670bar;
  wire n671bar;
  wire n672bar;
  wire n673bar;
  wire n674bar;
  wire n675bar;
  wire n676bar;
  wire n677bar;
  wire n678bar;
  wire n679bar;
  wire n680bar;
  wire n681bar;
  wire n682bar;
  wire n683bar;
  wire n684bar;
  wire n685bar;
  wire n686bar;
  wire n687bar;
  wire n688bar;
  wire n689bar;
  wire n690bar;
  wire n691bar;
  wire n692bar;
  wire n693bar;
  wire n694bar;
  wire n695bar;
  wire n696bar;
  wire n697bar;
  wire n698bar;
  wire n699bar;
  wire n700bar;
  wire n701bar;
  wire n702bar;
  wire n703bar;
  wire n704bar;
  wire n705bar;
  wire n706bar;
  wire n707bar;
  wire n708bar;
  wire n709bar;
  wire n710bar;
  wire n711bar;
  wire n712bar;
  wire n713bar;
  wire n714bar;
  wire n715bar;
  wire n716bar;
  wire n717bar;
  wire n718bar;
  wire n719bar;
  wire n720bar;
  wire n721bar;
  wire n722bar;
  wire n723bar;
  wire n724bar;
  wire n725bar;
  wire n726bar;
  wire n727bar;
  wire n728bar;
  wire n729bar;
  wire n730bar;
  wire n731bar;
  wire n732bar;
  wire n733bar;
  wire n734bar;
  wire n735bar;
  wire n736bar;
  wire n737bar;
  wire n738bar;
  wire n739bar;
  wire n740bar;
  wire n741bar;
  wire n742bar;
  wire n743bar;
  wire n744bar;
  wire n745bar;
  wire n746bar;
  wire n747bar;
  wire n748bar;
  wire n749bar;
  wire n750bar;
  wire n751bar;
  wire n752bar;
  wire n753bar;
  wire n754bar;
  wire n755bar;
  wire n756bar;
  wire n757bar;
  wire n758bar;
  wire n759bar;
  wire n760bar;
  wire n761bar;
  wire n762bar;
  wire n763bar;
  wire n764bar;
  wire n765bar;
  wire n766bar;
  wire n767bar;
  wire n768bar;
  wire n769bar;
  wire n770bar;
  wire n771bar;
  wire n772bar;
  wire n773bar;
  wire n774bar;
  wire n775bar;
  wire n776bar;
  wire n777bar;
  wire n778bar;
  wire n779bar;
  wire n780bar;
  wire n781bar;
  wire n782bar;
  wire n783bar;
  wire n784bar;
  wire n785bar;
  wire n786bar;
  wire n787bar;
  wire n788bar;
  wire n789bar;
  wire n790bar;
  wire n791bar;
  wire n792bar;
  wire n793bar;
  wire n794bar;
  wire n795bar;
  wire n796bar;
  wire n797bar;
  wire n798bar;
  wire n799bar;
  wire n800bar;
  wire n801bar;
  wire n802bar;
  wire n803bar;
  wire n804bar;
  wire n805bar;
  wire n806bar;
  wire n807bar;
  wire n808bar;
  wire n809bar;
  wire n810bar;
  wire n811bar;
  wire n812bar;
  wire n813bar;
  wire n814bar;
  wire n815bar;
  wire n816bar;
  wire n817bar;
  wire n818bar;
  wire n819bar;
  wire n820bar;
  wire n821bar;
  wire n822bar;
  wire n823bar;
  wire n824bar;
  wire n825bar;
  wire n826bar;
  wire n827bar;
  wire n828bar;
  wire n829bar;
  wire n830bar;
  wire n831bar;
  wire n832bar;
  wire n833bar;
  wire n834bar;
  wire n835bar;
  wire n836bar;
  wire n837bar;
  wire n838bar;
  wire n839bar;
  wire n840bar;
  wire n841bar;
  wire n842bar;
  wire n843bar;
  wire n844bar;
  wire n845bar;
  wire n846bar;
  wire n847bar;
  wire n848bar;
  wire n849bar;
  wire n850bar;
  wire n851bar;
  wire n852bar;
  wire n853bar;
  wire n854bar;
  wire n855bar;
  wire n856bar;
  wire n857bar;
  wire n858bar;
  wire n859bar;
  wire n860bar;
  wire n861bar;
  wire n862bar;
  wire n863bar;
  wire n864bar;
  wire n865bar;
  wire n866bar;
  wire n867bar;
  wire n868bar;
  wire n869bar;
  wire n870bar;
  wire n871bar;
  wire n872bar;
  wire n873bar;
  wire n874bar;
  wire n875bar;
  wire n876bar;
  wire n877bar;
  wire n878bar;
  wire n879bar;
  wire n880bar;
  wire n881bar;
  wire n882bar;
  wire n883bar;
  wire n884bar;
  wire n885bar;
  wire n886bar;
  wire n887bar;
  wire n888bar;
  wire n889bar;
  wire n890bar;
  wire n891bar;
  wire n892bar;
  wire n893bar;
  wire n894bar;
  wire n895bar;
  wire n896bar;
  wire n897bar;
  wire n898bar;
  wire n899bar;
  wire n900bar;
  wire n901bar;
  wire n902bar;
  wire n903bar;
  wire n904bar;
  wire n905bar;
  wire n906bar;
  wire n907bar;
  wire n908bar;
  wire n909bar;
  wire n910bar;
  wire n911bar;
  wire n912bar;
  wire n913bar;
  wire n914bar;
  wire n915bar;
  wire n916bar;
  wire n917bar;
  wire n918bar;
  wire n919bar;
  wire n920bar;
  wire n921bar;
  wire n922bar;
  wire n923bar;
  wire n924bar;
  wire n925bar;
  wire n926bar;
  wire n927bar;
  wire n928bar;
  wire n929bar;
  wire n930bar;
  wire n931bar;
  wire n932bar;
  wire n933bar;
  wire n934bar;
  wire n935bar;
  wire n936bar;
  wire n937bar;
  wire n938bar;
  wire n939bar;
  wire n940bar;
  wire n941bar;
  wire n942bar;
  wire n943bar;
  wire n944bar;
  wire n945bar;
  wire n946bar;
  wire n947bar;
  wire n948bar;
  wire n949bar;
  wire n950bar;
  wire n951bar;
  wire n952bar;
  wire n953bar;
  wire n954bar;
  wire n955bar;
  wire n956bar;
  wire n957bar;
  wire n958bar;
  wire n959bar;
  wire n960bar;
  wire n961bar;
  wire n962bar;
  wire n963bar;
  wire n964bar;
  wire n965bar;
  wire n966bar;
  wire n967bar;
  wire n968bar;
  wire n969bar;
  wire n970bar;
  wire n971bar;
  wire n972bar;
//wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];
  assign in_81bar = inbar[81];
  assign in_80bar = inbar[80];
  assign in_79bar = inbar[79];
  assign in_78bar = inbar[78];
  assign in_77bar = inbar[77];
  assign in_76bar = inbar[76];
  assign in_75bar = inbar[75];
  assign in_74bar = inbar[74];
  assign in_73bar = inbar[73];
  assign in_72bar = inbar[72];
  assign in_71bar = inbar[71];
  assign in_70bar = inbar[70];
  assign in_69bar = inbar[69];
  assign in_68bar = inbar[68];
  assign in_67bar = inbar[67];
  assign in_66bar = inbar[66];
  assign in_65bar = inbar[65];
  assign in_64bar = inbar[64];
  assign in_63bar = inbar[63];
  assign in_62bar = inbar[62];
  assign in_61bar = inbar[61];
  assign in_60bar = inbar[60];
  assign in_59bar = inbar[59];
  assign in_58bar = inbar[58];
  assign in_57bar = inbar[57];
  assign in_56bar = inbar[56];
  assign in_55bar = inbar[55];
  assign in_54bar = inbar[54];
  assign in_53bar = inbar[53];
  assign in_52bar = inbar[52];
  assign in_51bar = inbar[51];
  assign in_50bar = inbar[50];
  assign in_49bar = inbar[49];
  assign in_48bar = inbar[48];
  assign in_47bar = inbar[47];
  assign in_46bar = inbar[46];
  assign in_45bar = inbar[45];
  assign in_44bar = inbar[44];
  assign in_43bar = inbar[43];
  assign in_42bar = inbar[42];
  assign in_41bar = inbar[41];
  assign in_40bar = inbar[40];
  assign in_39bar = inbar[39];
  assign in_38bar = inbar[38];
  assign in_37bar = inbar[37];
  assign in_36bar = inbar[36];
  assign in_35bar = inbar[35];
  assign in_34bar = inbar[34];
  assign in_33bar = inbar[33];
  assign in_32bar = inbar[32];
  assign in_31bar = inbar[31];
  assign in_30bar = inbar[30];
  assign in_29bar = inbar[29];
  assign in_28bar = inbar[28];
  assign in_27bar = inbar[27];
  assign in_26bar = inbar[26];
  assign in_25bar = inbar[25];
  assign in_24bar = inbar[24];
  assign in_23bar = inbar[23];
  assign in_22bar = inbar[22];
  assign in_21bar = inbar[21];
  assign in_20bar = inbar[20];
  assign in_19bar = inbar[19];
  assign in_18bar = inbar[18];
  assign in_17bar = inbar[17];
  assign in_16bar = inbar[16];
  assign in_15bar = inbar[15];
  assign in_14bar = inbar[14];
  assign in_13bar = inbar[13];
  assign in_12bar = inbar[12];
  assign in_11bar = inbar[11];
  assign in_10bar = inbar[10];
  assign in_9bar = inbar[9];
  assign in_8bar = inbar[8];
  assign in_7bar = inbar[7];
  assign in_6bar = inbar[6];
  assign in_5bar = inbar[5];
  assign in_4bar = inbar[4];
  assign in_3bar = inbar[3];
  assign in_2bar = inbar[2];
  assign in_1bar = inbar[1];
  assign in_0bar = inbar[0];
//assign_done

  OR2_X1 U1 ( .A1(n972), .A2(n971), .ZN(out[7]) );
  AND2_X1 U1bar ( .A1(n972bar), .A2(n971bar), .ZN(outbar[7]) );
  OR2_X1 U2 ( .A1(n970), .A2(n969), .ZN(n971) );
  AND2_X1 U2bar ( .A1(n970bar), .A2(n969bar), .ZN(n971bar) );
  OR2_X1 U3 ( .A1(n968), .A2(n967), .ZN(n969) );
  AND2_X1 U3bar ( .A1(n968bar), .A2(n967bar), .ZN(n969bar) );
  OR2_X1 U4 ( .A1(n966), .A2(n965), .ZN(n967) );
  AND2_X1 U4bar ( .A1(n966bar), .A2(n965bar), .ZN(n967bar) );
  OR2_X1 U5 ( .A1(n964), .A2(n963), .ZN(n968) );
  AND2_X1 U5bar ( .A1(n964bar), .A2(n963bar), .ZN(n968bar) );
  OR2_X1 U6 ( .A1(in[116]), .A2(n962), .ZN(n963) );
  AND2_X1 U6bar ( .A1(inbar[116]), .A2(n962bar), .ZN(n963bar) );
  OR2_X1 U7 ( .A1(n961), .A2(n960), .ZN(n970) );
  AND2_X1 U7bar ( .A1(n961bar), .A2(n960bar), .ZN(n970bar) );
  OR2_X1 U8 ( .A1(in[150]), .A2(in[127]), .ZN(n960) );
  AND2_X1 U8bar ( .A1(inbar[150]), .A2(inbar[127]), .ZN(n960bar) );
  OR2_X1 U9 ( .A1(in[160]), .A2(n959), .ZN(n961) );
  AND2_X1 U9bar ( .A1(inbar[160]), .A2(n959bar), .ZN(n961bar) );
  OR2_X1 U10 ( .A1(in[252]), .A2(in[168]), .ZN(n959) );
  AND2_X1 U10bar ( .A1(inbar[252]), .A2(inbar[168]), .ZN(n959bar) );
  OR2_X1 U11 ( .A1(n958), .A2(n957), .ZN(n972) );
  AND2_X1 U11bar ( .A1(n958bar), .A2(n957bar), .ZN(n972bar) );
  OR2_X1 U12 ( .A1(n956), .A2(n955), .ZN(n957) );
  AND2_X1 U12bar ( .A1(n956bar), .A2(n955bar), .ZN(n957bar) );
  OR2_X1 U13 ( .A1(in_17), .A2(in[96]), .ZN(n955) );
  AND2_X1 U13bar ( .A1(in_17bar), .A2(inbar[96]), .ZN(n955bar) );
  OR2_X1 U14 ( .A1(in_23), .A2(n954), .ZN(n956) );
  AND2_X1 U14bar ( .A1(in_23bar), .A2(n954bar), .ZN(n956bar) );
  OR2_X1 U15 ( .A1(in_31), .A2(in_26), .ZN(n954) );
  AND2_X1 U15bar ( .A1(in_31bar), .A2(in_26bar), .ZN(n954bar) );
  OR2_X1 U16 ( .A1(n953), .A2(n952), .ZN(n958) );
  AND2_X1 U16bar ( .A1(n953bar), .A2(n952bar), .ZN(n958bar) );
  OR2_X1 U17 ( .A1(in_58), .A2(in_4), .ZN(n952) );
  AND2_X1 U17bar ( .A1(in_58bar), .A2(in_4bar), .ZN(n952bar) );
  OR2_X1 U18 ( .A1(in_59), .A2(n951), .ZN(n953) );
  AND2_X1 U18bar ( .A1(in_59bar), .A2(n951bar), .ZN(n953bar) );
  OR2_X1 U19 ( .A1(in_71), .A2(in_62), .ZN(n951) );
  AND2_X1 U19bar ( .A1(in_71bar), .A2(in_62bar), .ZN(n951bar) );
  OR2_X1 U20 ( .A1(n950), .A2(n949), .ZN(out[6]) );
  AND2_X1 U20bar ( .A1(n950bar), .A2(n949bar), .ZN(outbar[6]) );
  OR2_X1 U21 ( .A1(n948), .A2(n947), .ZN(n949) );
  AND2_X1 U21bar ( .A1(n948bar), .A2(n947bar), .ZN(n949bar) );
  OR2_X1 U22 ( .A1(n946), .A2(n945), .ZN(n947) );
  AND2_X1 U22bar ( .A1(n946bar), .A2(n945bar), .ZN(n947bar) );
  OR2_X1 U23 ( .A1(n944), .A2(n943), .ZN(n945) );
  AND2_X1 U23bar ( .A1(n944bar), .A2(n943bar), .ZN(n945bar) );
  OR2_X1 U24 ( .A1(n942), .A2(n941), .ZN(n946) );
  AND2_X1 U24bar ( .A1(n942bar), .A2(n941bar), .ZN(n946bar) );
  OR2_X1 U25 ( .A1(in[101]), .A2(n940), .ZN(n941) );
  AND2_X1 U25bar ( .A1(inbar[101]), .A2(n940bar), .ZN(n941bar) );
  OR2_X1 U26 ( .A1(n939), .A2(n938), .ZN(n948) );
  AND2_X1 U26bar ( .A1(n939bar), .A2(n938bar), .ZN(n948bar) );
  OR2_X1 U27 ( .A1(in[114]), .A2(in[104]), .ZN(n938) );
  AND2_X1 U27bar ( .A1(inbar[114]), .A2(inbar[104]), .ZN(n938bar) );
  OR2_X1 U28 ( .A1(in[128]), .A2(n937), .ZN(n939) );
  AND2_X1 U28bar ( .A1(inbar[128]), .A2(n937bar), .ZN(n939bar) );
  OR2_X1 U29 ( .A1(in[136]), .A2(in[134]), .ZN(n937) );
  AND2_X1 U29bar ( .A1(inbar[136]), .A2(inbar[134]), .ZN(n937bar) );
  OR2_X1 U30 ( .A1(n936), .A2(n935), .ZN(n950) );
  AND2_X1 U30bar ( .A1(n936bar), .A2(n935bar), .ZN(n950bar) );
  OR2_X1 U31 ( .A1(n934), .A2(n933), .ZN(n935) );
  AND2_X1 U31bar ( .A1(n934bar), .A2(n933bar), .ZN(n935bar) );
  OR2_X1 U32 ( .A1(in[177]), .A2(in[164]), .ZN(n933) );
  AND2_X1 U32bar ( .A1(inbar[177]), .A2(inbar[164]), .ZN(n933bar) );
  OR2_X1 U33 ( .A1(in[212]), .A2(n932), .ZN(n934) );
  AND2_X1 U33bar ( .A1(inbar[212]), .A2(n932bar), .ZN(n934bar) );
  OR2_X1 U34 ( .A1(in[248]), .A2(in[221]), .ZN(n932) );
  AND2_X1 U34bar ( .A1(inbar[248]), .A2(inbar[221]), .ZN(n932bar) );
  OR2_X1 U35 ( .A1(n931), .A2(n930), .ZN(n936) );
  AND2_X1 U35bar ( .A1(n931bar), .A2(n930bar), .ZN(n936bar) );
  OR2_X1 U36 ( .A1(in_18), .A2(in[93]), .ZN(n930) );
  AND2_X1 U36bar ( .A1(in_18bar), .A2(inbar[93]), .ZN(n930bar) );
  OR2_X1 U37 ( .A1(in_31), .A2(n929), .ZN(n931) );
  AND2_X1 U37bar ( .A1(in_31bar), .A2(n929bar), .ZN(n931bar) );
  OR2_X1 U38 ( .A1(in_7), .A2(in_39), .ZN(n929) );
  AND2_X1 U38bar ( .A1(in_7bar), .A2(in_39bar), .ZN(n929bar) );
  OR2_X1 U39 ( .A1(n928), .A2(n927), .ZN(out[5]) );
  AND2_X1 U39bar ( .A1(n928bar), .A2(n927bar), .ZN(outbar[5]) );
  OR2_X1 U40 ( .A1(n926), .A2(n925), .ZN(n927) );
  AND2_X1 U40bar ( .A1(n926bar), .A2(n925bar), .ZN(n927bar) );
  OR2_X1 U41 ( .A1(n924), .A2(n923), .ZN(n925) );
  AND2_X1 U41bar ( .A1(n924bar), .A2(n923bar), .ZN(n925bar) );
  OR2_X1 U42 ( .A1(n922), .A2(n921), .ZN(n923) );
  AND2_X1 U42bar ( .A1(n922bar), .A2(n921bar), .ZN(n923bar) );
  OR2_X1 U43 ( .A1(n940), .A2(n920), .ZN(n924) );
  AND2_X1 U43bar ( .A1(n940bar), .A2(n920bar), .ZN(n924bar) );
  OR2_X1 U44 ( .A1(in[111]), .A2(n919), .ZN(n920) );
  AND2_X1 U44bar ( .A1(inbar[111]), .A2(n919bar), .ZN(n920bar) );
  OR2_X1 U45 ( .A1(n918), .A2(n917), .ZN(n940) );
  AND2_X1 U45bar ( .A1(n918bar), .A2(n917bar), .ZN(n940bar) );
  OR2_X1 U46 ( .A1(n916), .A2(n915), .ZN(n917) );
  AND2_X1 U46bar ( .A1(n916bar), .A2(n915bar), .ZN(n917bar) );
  OR2_X1 U47 ( .A1(n914), .A2(n913), .ZN(n915) );
  AND2_X1 U47bar ( .A1(n914bar), .A2(n913bar), .ZN(n915bar) );
  OR2_X1 U48 ( .A1(in[140]), .A2(in[131]), .ZN(n913) );
  AND2_X1 U48bar ( .A1(inbar[140]), .A2(inbar[131]), .ZN(n913bar) );
  OR2_X1 U49 ( .A1(in[160]), .A2(in[144]), .ZN(n914) );
  AND2_X1 U49bar ( .A1(inbar[160]), .A2(inbar[144]), .ZN(n914bar) );
  OR2_X1 U50 ( .A1(n912), .A2(n911), .ZN(n916) );
  AND2_X1 U50bar ( .A1(n912bar), .A2(n911bar), .ZN(n916bar) );
  OR2_X1 U51 ( .A1(in[179]), .A2(in[174]), .ZN(n911) );
  AND2_X1 U51bar ( .A1(inbar[179]), .A2(inbar[174]), .ZN(n911bar) );
  OR2_X1 U52 ( .A1(in[188]), .A2(in[184]), .ZN(n912) );
  AND2_X1 U52bar ( .A1(inbar[188]), .A2(inbar[184]), .ZN(n912bar) );
  OR2_X1 U53 ( .A1(n910), .A2(n909), .ZN(n918) );
  AND2_X1 U53bar ( .A1(n910bar), .A2(n909bar), .ZN(n918bar) );
  OR2_X1 U54 ( .A1(n908), .A2(n907), .ZN(n909) );
  AND2_X1 U54bar ( .A1(n908bar), .A2(n907bar), .ZN(n909bar) );
  OR2_X1 U55 ( .A1(in[216]), .A2(in[200]), .ZN(n907) );
  AND2_X1 U55bar ( .A1(inbar[216]), .A2(inbar[200]), .ZN(n907bar) );
  OR2_X1 U56 ( .A1(in[228]), .A2(in[224]), .ZN(n908) );
  AND2_X1 U56bar ( .A1(inbar[228]), .A2(inbar[224]), .ZN(n908bar) );
  OR2_X1 U57 ( .A1(n906), .A2(n905), .ZN(n910) );
  AND2_X1 U57bar ( .A1(n906bar), .A2(n905bar), .ZN(n910bar) );
  OR2_X1 U58 ( .A1(in[247]), .A2(in[235]), .ZN(n905) );
  AND2_X1 U58bar ( .A1(inbar[247]), .A2(inbar[235]), .ZN(n905bar) );
  OR2_X1 U59 ( .A1(in_42), .A2(in[83]), .ZN(n906) );
  AND2_X1 U59bar ( .A1(in_42bar), .A2(inbar[83]), .ZN(n906bar) );
  OR2_X1 U60 ( .A1(n904), .A2(n903), .ZN(n926) );
  AND2_X1 U60bar ( .A1(n904bar), .A2(n903bar), .ZN(n926bar) );
  OR2_X1 U61 ( .A1(in[166]), .A2(in[123]), .ZN(n903) );
  AND2_X1 U61bar ( .A1(inbar[166]), .A2(inbar[123]), .ZN(n903bar) );
  OR2_X1 U62 ( .A1(in[170]), .A2(n902), .ZN(n904) );
  AND2_X1 U62bar ( .A1(inbar[170]), .A2(n902bar), .ZN(n904bar) );
  OR2_X1 U63 ( .A1(in[194]), .A2(in[183]), .ZN(n902) );
  AND2_X1 U63bar ( .A1(inbar[194]), .A2(inbar[183]), .ZN(n902bar) );
  OR2_X1 U64 ( .A1(n901), .A2(n900), .ZN(n928) );
  AND2_X1 U64bar ( .A1(n901bar), .A2(n900bar), .ZN(n928bar) );
  OR2_X1 U65 ( .A1(n899), .A2(n898), .ZN(n900) );
  AND2_X1 U65bar ( .A1(n899bar), .A2(n898bar), .ZN(n900bar) );
  OR2_X1 U66 ( .A1(in[241]), .A2(in[238]), .ZN(n898) );
  AND2_X1 U66bar ( .A1(inbar[241]), .A2(inbar[238]), .ZN(n898bar) );
  OR2_X1 U67 ( .A1(in[250]), .A2(n897), .ZN(n899) );
  AND2_X1 U67bar ( .A1(inbar[250]), .A2(n897bar), .ZN(n899bar) );
  OR2_X1 U68 ( .A1(in_24), .A2(in[84]), .ZN(n897) );
  AND2_X1 U68bar ( .A1(in_24bar), .A2(inbar[84]), .ZN(n897bar) );
  OR2_X1 U69 ( .A1(n896), .A2(n895), .ZN(n901) );
  AND2_X1 U69bar ( .A1(n896bar), .A2(n895bar), .ZN(n901bar) );
  OR2_X1 U70 ( .A1(in_41), .A2(in_29), .ZN(n895) );
  AND2_X1 U70bar ( .A1(in_41bar), .A2(in_29bar), .ZN(n895bar) );
  OR2_X1 U71 ( .A1(in_66), .A2(n894), .ZN(n896) );
  AND2_X1 U71bar ( .A1(in_66bar), .A2(n894bar), .ZN(n896bar) );
  OR2_X1 U72 ( .A1(in_76), .A2(in_71), .ZN(n894) );
  AND2_X1 U72bar ( .A1(in_76bar), .A2(in_71bar), .ZN(n894bar) );
  OR2_X1 U73 ( .A1(n893), .A2(n892), .ZN(out[4]) );
  AND2_X1 U73bar ( .A1(n893bar), .A2(n892bar), .ZN(outbar[4]) );
  OR2_X1 U74 ( .A1(n891), .A2(n890), .ZN(n892) );
  AND2_X1 U74bar ( .A1(n891bar), .A2(n890bar), .ZN(n892bar) );
  OR2_X1 U75 ( .A1(n889), .A2(n888), .ZN(n890) );
  AND2_X1 U75bar ( .A1(n889bar), .A2(n888bar), .ZN(n890bar) );
  OR2_X1 U76 ( .A1(n922), .A2(n887), .ZN(n888) );
  AND2_X1 U76bar ( .A1(n922bar), .A2(n887bar), .ZN(n888bar) );
  OR2_X1 U77 ( .A1(n886), .A2(n885), .ZN(n922) );
  AND2_X1 U77bar ( .A1(n886bar), .A2(n885bar), .ZN(n922bar) );
  OR2_X1 U78 ( .A1(n884), .A2(n883), .ZN(n885) );
  AND2_X1 U78bar ( .A1(n884bar), .A2(n883bar), .ZN(n885bar) );
  OR2_X1 U79 ( .A1(n882), .A2(n881), .ZN(n883) );
  AND2_X1 U79bar ( .A1(n882bar), .A2(n881bar), .ZN(n883bar) );
  OR2_X1 U80 ( .A1(in[118]), .A2(in[109]), .ZN(n881) );
  AND2_X1 U80bar ( .A1(inbar[118]), .A2(inbar[109]), .ZN(n881bar) );
  OR2_X1 U81 ( .A1(in[139]), .A2(in[120]), .ZN(n882) );
  AND2_X1 U81bar ( .A1(inbar[139]), .A2(inbar[120]), .ZN(n882bar) );
  OR2_X1 U82 ( .A1(n880), .A2(n879), .ZN(n884) );
  AND2_X1 U82bar ( .A1(n880bar), .A2(n879bar), .ZN(n884bar) );
  OR2_X1 U83 ( .A1(in[198]), .A2(in[154]), .ZN(n879) );
  AND2_X1 U83bar ( .A1(inbar[198]), .A2(inbar[154]), .ZN(n879bar) );
  OR2_X1 U84 ( .A1(in[210]), .A2(in[205]), .ZN(n880) );
  AND2_X1 U84bar ( .A1(inbar[210]), .A2(inbar[205]), .ZN(n880bar) );
  OR2_X1 U85 ( .A1(n878), .A2(n877), .ZN(n886) );
  AND2_X1 U85bar ( .A1(n878bar), .A2(n877bar), .ZN(n886bar) );
  OR2_X1 U86 ( .A1(n876), .A2(n875), .ZN(n877) );
  AND2_X1 U86bar ( .A1(n876bar), .A2(n875bar), .ZN(n877bar) );
  OR2_X1 U87 ( .A1(in[219]), .A2(in[217]), .ZN(n875) );
  AND2_X1 U87bar ( .A1(inbar[219]), .A2(inbar[217]), .ZN(n875bar) );
  OR2_X1 U88 ( .A1(in[86]), .A2(in[252]), .ZN(n876) );
  AND2_X1 U88bar ( .A1(inbar[86]), .A2(inbar[252]), .ZN(n876bar) );
  OR2_X1 U89 ( .A1(n874), .A2(n873), .ZN(n878) );
  AND2_X1 U89bar ( .A1(n874bar), .A2(n873bar), .ZN(n878bar) );
  OR2_X1 U90 ( .A1(in_40), .A2(in[91]), .ZN(n873) );
  AND2_X1 U90bar ( .A1(in_40bar), .A2(inbar[91]), .ZN(n873bar) );
  OR2_X1 U91 ( .A1(in_8), .A2(in_46), .ZN(n874) );
  AND2_X1 U91bar ( .A1(in_8bar), .A2(in_46bar), .ZN(n874bar) );
  OR2_X1 U92 ( .A1(n872), .A2(n871), .ZN(n889) );
  AND2_X1 U92bar ( .A1(n872bar), .A2(n871bar), .ZN(n889bar) );
  OR2_X1 U93 ( .A1(in[117]), .A2(n943), .ZN(n871) );
  AND2_X1 U93bar ( .A1(inbar[117]), .A2(n943bar), .ZN(n871bar) );
  OR2_X1 U94 ( .A1(n870), .A2(n869), .ZN(n943) );
  AND2_X1 U94bar ( .A1(n870bar), .A2(n869bar), .ZN(n943bar) );
  OR2_X1 U95 ( .A1(n868), .A2(n867), .ZN(n869) );
  AND2_X1 U95bar ( .A1(n868bar), .A2(n867bar), .ZN(n869bar) );
  OR2_X1 U96 ( .A1(n866), .A2(n865), .ZN(n867) );
  AND2_X1 U96bar ( .A1(n866bar), .A2(n865bar), .ZN(n867bar) );
  OR2_X1 U97 ( .A1(n864), .A2(n863), .ZN(n865) );
  AND2_X1 U97bar ( .A1(n864bar), .A2(n863bar), .ZN(n865bar) );
  OR2_X1 U98 ( .A1(in[108]), .A2(n919), .ZN(n866) );
  AND2_X1 U98bar ( .A1(inbar[108]), .A2(n919bar), .ZN(n866bar) );
  OR2_X1 U99 ( .A1(n862), .A2(n861), .ZN(n919) );
  AND2_X1 U99bar ( .A1(n862bar), .A2(n861bar), .ZN(n919bar) );
  OR2_X1 U100 ( .A1(n860), .A2(n859), .ZN(n861) );
  AND2_X1 U100bar ( .A1(n860bar), .A2(n859bar), .ZN(n861bar) );
  OR2_X1 U101 ( .A1(n858), .A2(n857), .ZN(n859) );
  AND2_X1 U101bar ( .A1(n858bar), .A2(n857bar), .ZN(n859bar) );
  OR2_X1 U102 ( .A1(in[119]), .A2(in[105]), .ZN(n857) );
  AND2_X1 U102bar ( .A1(inbar[119]), .A2(inbar[105]), .ZN(n857bar) );
  OR2_X1 U103 ( .A1(in[186]), .A2(in[175]), .ZN(n858) );
  AND2_X1 U103bar ( .A1(inbar[186]), .A2(inbar[175]), .ZN(n858bar) );
  OR2_X1 U104 ( .A1(n856), .A2(n855), .ZN(n860) );
  AND2_X1 U104bar ( .A1(n856bar), .A2(n855bar), .ZN(n860bar) );
  OR2_X1 U105 ( .A1(in[202]), .A2(in[193]), .ZN(n855) );
  AND2_X1 U105bar ( .A1(inbar[202]), .A2(inbar[193]), .ZN(n855bar) );
  OR2_X1 U106 ( .A1(in[225]), .A2(in[208]), .ZN(n856) );
  AND2_X1 U106bar ( .A1(inbar[225]), .A2(inbar[208]), .ZN(n856bar) );
  OR2_X1 U107 ( .A1(n854), .A2(n853), .ZN(n862) );
  AND2_X1 U107bar ( .A1(n854bar), .A2(n853bar), .ZN(n862bar) );
  OR2_X1 U108 ( .A1(n852), .A2(n851), .ZN(n853) );
  AND2_X1 U108bar ( .A1(n852bar), .A2(n851bar), .ZN(n853bar) );
  OR2_X1 U109 ( .A1(in_1), .A2(in[85]), .ZN(n851) );
  AND2_X1 U109bar ( .A1(in_1bar), .A2(inbar[85]), .ZN(n851bar) );
  OR2_X1 U110 ( .A1(in_23), .A2(in_19), .ZN(n852) );
  AND2_X1 U110bar ( .A1(in_23bar), .A2(in_19bar), .ZN(n852bar) );
  OR2_X1 U111 ( .A1(n850), .A2(n849), .ZN(n854) );
  AND2_X1 U111bar ( .A1(n850bar), .A2(n849bar), .ZN(n854bar) );
  OR2_X1 U112 ( .A1(in_43), .A2(in_33), .ZN(n849) );
  AND2_X1 U112bar ( .A1(in_43bar), .A2(in_33bar), .ZN(n849bar) );
  OR2_X1 U113 ( .A1(in_63), .A2(in_44), .ZN(n850) );
  AND2_X1 U113bar ( .A1(in_63bar), .A2(in_44bar), .ZN(n850bar) );
  OR2_X1 U114 ( .A1(n848), .A2(n847), .ZN(n868) );
  AND2_X1 U114bar ( .A1(n848bar), .A2(n847bar), .ZN(n868bar) );
  OR2_X1 U115 ( .A1(in[141]), .A2(in[112]), .ZN(n847) );
  AND2_X1 U115bar ( .A1(inbar[141]), .A2(inbar[112]), .ZN(n847bar) );
  OR2_X1 U116 ( .A1(in[147]), .A2(n846), .ZN(n848) );
  AND2_X1 U116bar ( .A1(inbar[147]), .A2(n846bar), .ZN(n848bar) );
  OR2_X1 U117 ( .A1(in[181]), .A2(in[167]), .ZN(n846) );
  AND2_X1 U117bar ( .A1(inbar[181]), .A2(inbar[167]), .ZN(n846bar) );
  OR2_X1 U118 ( .A1(n845), .A2(n844), .ZN(n870) );
  AND2_X1 U118bar ( .A1(n845bar), .A2(n844bar), .ZN(n870bar) );
  OR2_X1 U119 ( .A1(n843), .A2(n842), .ZN(n844) );
  AND2_X1 U119bar ( .A1(n843bar), .A2(n842bar), .ZN(n844bar) );
  OR2_X1 U120 ( .A1(in[229]), .A2(in[201]), .ZN(n842) );
  AND2_X1 U120bar ( .A1(inbar[229]), .A2(inbar[201]), .ZN(n842bar) );
  OR2_X1 U121 ( .A1(in[237]), .A2(n841), .ZN(n843) );
  AND2_X1 U121bar ( .A1(inbar[237]), .A2(n841bar), .ZN(n843bar) );
  OR2_X1 U122 ( .A1(in[94]), .A2(in[253]), .ZN(n841) );
  AND2_X1 U122bar ( .A1(inbar[94]), .A2(inbar[253]), .ZN(n841bar) );
  OR2_X1 U123 ( .A1(n840), .A2(n839), .ZN(n845) );
  AND2_X1 U123bar ( .A1(n840bar), .A2(n839bar), .ZN(n845bar) );
  OR2_X1 U124 ( .A1(in_21), .A2(in[96]), .ZN(n839) );
  AND2_X1 U124bar ( .A1(in_21bar), .A2(inbar[96]), .ZN(n839bar) );
  OR2_X1 U125 ( .A1(in_25), .A2(n838), .ZN(n840) );
  AND2_X1 U125bar ( .A1(in_25bar), .A2(n838bar), .ZN(n840bar) );
  OR2_X1 U126 ( .A1(in_81), .A2(in_45), .ZN(n838) );
  AND2_X1 U126bar ( .A1(in_81bar), .A2(in_45bar), .ZN(n838bar) );
  OR2_X1 U127 ( .A1(n837), .A2(n836), .ZN(n891) );
  AND2_X1 U127bar ( .A1(n837bar), .A2(n836bar), .ZN(n891bar) );
  OR2_X1 U128 ( .A1(in[142]), .A2(in[124]), .ZN(n836) );
  AND2_X1 U128bar ( .A1(inbar[142]), .A2(inbar[124]), .ZN(n836bar) );
  OR2_X1 U129 ( .A1(in[150]), .A2(n835), .ZN(n837) );
  AND2_X1 U129bar ( .A1(inbar[150]), .A2(n835bar), .ZN(n837bar) );
  OR2_X1 U130 ( .A1(in[172]), .A2(in[155]), .ZN(n835) );
  AND2_X1 U130bar ( .A1(inbar[172]), .A2(inbar[155]), .ZN(n835bar) );
  OR2_X1 U131 ( .A1(n834), .A2(n833), .ZN(n893) );
  AND2_X1 U131bar ( .A1(n834bar), .A2(n833bar), .ZN(n893bar) );
  OR2_X1 U132 ( .A1(n832), .A2(n831), .ZN(n833) );
  AND2_X1 U132bar ( .A1(n832bar), .A2(n831bar), .ZN(n833bar) );
  OR2_X1 U133 ( .A1(in[196]), .A2(in[173]), .ZN(n831) );
  AND2_X1 U133bar ( .A1(inbar[196]), .A2(inbar[173]), .ZN(n831bar) );
  OR2_X1 U134 ( .A1(in[222]), .A2(n830), .ZN(n832) );
  AND2_X1 U134bar ( .A1(inbar[222]), .A2(n830bar), .ZN(n832bar) );
  OR2_X1 U135 ( .A1(in[227]), .A2(in[226]), .ZN(n830) );
  AND2_X1 U135bar ( .A1(inbar[227]), .A2(inbar[226]), .ZN(n830bar) );
  OR2_X1 U136 ( .A1(n829), .A2(n828), .ZN(n834) );
  AND2_X1 U136bar ( .A1(n829bar), .A2(n828bar), .ZN(n834bar) );
  OR2_X1 U137 ( .A1(in[249]), .A2(in[231]), .ZN(n828) );
  AND2_X1 U137bar ( .A1(inbar[249]), .A2(inbar[231]), .ZN(n828bar) );
  OR2_X1 U138 ( .A1(in_28), .A2(n827), .ZN(n829) );
  AND2_X1 U138bar ( .A1(in_28bar), .A2(n827bar), .ZN(n829bar) );
  OR2_X1 U139 ( .A1(in_52), .A2(in_47), .ZN(n827) );
  AND2_X1 U139bar ( .A1(in_52bar), .A2(in_47bar), .ZN(n827bar) );
  OR2_X1 U140 ( .A1(n826), .A2(n825), .ZN(out[3]) );
  AND2_X1 U140bar ( .A1(n826bar), .A2(n825bar), .ZN(outbar[3]) );
  OR2_X1 U141 ( .A1(n824), .A2(n823), .ZN(n825) );
  AND2_X1 U141bar ( .A1(n824bar), .A2(n823bar), .ZN(n825bar) );
  OR2_X1 U142 ( .A1(n822), .A2(n821), .ZN(n823) );
  AND2_X1 U142bar ( .A1(n822bar), .A2(n821bar), .ZN(n823bar) );
  OR2_X1 U143 ( .A1(n820), .A2(n819), .ZN(n821) );
  AND2_X1 U143bar ( .A1(n820bar), .A2(n819bar), .ZN(n821bar) );
  OR2_X1 U144 ( .A1(n964), .A2(n818), .ZN(n822) );
  AND2_X1 U144bar ( .A1(n964bar), .A2(n818bar), .ZN(n822bar) );
  OR2_X1 U145 ( .A1(in[118]), .A2(n817), .ZN(n818) );
  AND2_X1 U145bar ( .A1(inbar[118]), .A2(n817bar), .ZN(n818bar) );
  OR2_X1 U146 ( .A1(n816), .A2(n815), .ZN(n964) );
  AND2_X1 U146bar ( .A1(n816bar), .A2(n815bar), .ZN(n964bar) );
  OR2_X1 U147 ( .A1(n814), .A2(n813), .ZN(n815) );
  AND2_X1 U147bar ( .A1(n814bar), .A2(n813bar), .ZN(n815bar) );
  OR2_X1 U148 ( .A1(n812), .A2(n811), .ZN(n813) );
  AND2_X1 U148bar ( .A1(n812bar), .A2(n811bar), .ZN(n813bar) );
  OR2_X1 U149 ( .A1(in[122]), .A2(in[111]), .ZN(n811) );
  AND2_X1 U149bar ( .A1(inbar[122]), .A2(inbar[111]), .ZN(n811bar) );
  OR2_X1 U150 ( .A1(in[154]), .A2(in[151]), .ZN(n812) );
  AND2_X1 U150bar ( .A1(inbar[154]), .A2(inbar[151]), .ZN(n812bar) );
  OR2_X1 U151 ( .A1(n810), .A2(n809), .ZN(n814) );
  AND2_X1 U151bar ( .A1(n810bar), .A2(n809bar), .ZN(n814bar) );
  OR2_X1 U152 ( .A1(in[187]), .A2(in[177]), .ZN(n809) );
  AND2_X1 U152bar ( .A1(inbar[187]), .A2(inbar[177]), .ZN(n809bar) );
  OR2_X1 U153 ( .A1(in[200]), .A2(in[192]), .ZN(n810) );
  AND2_X1 U153bar ( .A1(inbar[200]), .A2(inbar[192]), .ZN(n810bar) );
  OR2_X1 U154 ( .A1(n808), .A2(n807), .ZN(n816) );
  AND2_X1 U154bar ( .A1(n808bar), .A2(n807bar), .ZN(n816bar) );
  OR2_X1 U155 ( .A1(n806), .A2(n805), .ZN(n807) );
  AND2_X1 U155bar ( .A1(n806bar), .A2(n805bar), .ZN(n807bar) );
  OR2_X1 U156 ( .A1(in[225]), .A2(in[207]), .ZN(n805) );
  AND2_X1 U156bar ( .A1(inbar[225]), .A2(inbar[207]), .ZN(n805bar) );
  OR2_X1 U157 ( .A1(in[98]), .A2(in[226]), .ZN(n806) );
  AND2_X1 U157bar ( .A1(inbar[98]), .A2(inbar[226]), .ZN(n806bar) );
  OR2_X1 U158 ( .A1(n804), .A2(n803), .ZN(n808) );
  AND2_X1 U158bar ( .A1(n804bar), .A2(n803bar), .ZN(n808bar) );
  OR2_X1 U159 ( .A1(in_20), .A2(in_16), .ZN(n803) );
  AND2_X1 U159bar ( .A1(in_20bar), .A2(in_16bar), .ZN(n803bar) );
  OR2_X1 U160 ( .A1(in_55), .A2(in_45), .ZN(n804) );
  AND2_X1 U160bar ( .A1(in_55bar), .A2(in_45bar), .ZN(n804bar) );
  OR2_X1 U161 ( .A1(n802), .A2(n801), .ZN(n824) );
  AND2_X1 U161bar ( .A1(n802bar), .A2(n801bar), .ZN(n824bar) );
  OR2_X1 U162 ( .A1(in[162]), .A2(in[149]), .ZN(n801) );
  AND2_X1 U162bar ( .A1(inbar[162]), .A2(inbar[149]), .ZN(n801bar) );
  OR2_X1 U163 ( .A1(in[163]), .A2(n800), .ZN(n802) );
  AND2_X1 U163bar ( .A1(inbar[163]), .A2(n800bar), .ZN(n802bar) );
  OR2_X1 U164 ( .A1(in[191]), .A2(in[189]), .ZN(n800) );
  AND2_X1 U164bar ( .A1(inbar[191]), .A2(inbar[189]), .ZN(n800bar) );
  OR2_X1 U165 ( .A1(n799), .A2(n798), .ZN(n826) );
  AND2_X1 U165bar ( .A1(n799bar), .A2(n798bar), .ZN(n826bar) );
  OR2_X1 U166 ( .A1(n797), .A2(n796), .ZN(n798) );
  AND2_X1 U166bar ( .A1(n797bar), .A2(n796bar), .ZN(n798bar) );
  OR2_X1 U167 ( .A1(in[212]), .A2(in[193]), .ZN(n796) );
  AND2_X1 U167bar ( .A1(inbar[212]), .A2(inbar[193]), .ZN(n796bar) );
  OR2_X1 U168 ( .A1(in[238]), .A2(n795), .ZN(n797) );
  AND2_X1 U168bar ( .A1(inbar[238]), .A2(n795bar), .ZN(n797bar) );
  OR2_X1 U169 ( .A1(in[88]), .A2(in[247]), .ZN(n795) );
  AND2_X1 U169bar ( .A1(inbar[88]), .A2(inbar[247]), .ZN(n795bar) );
  OR2_X1 U170 ( .A1(n794), .A2(n793), .ZN(n799) );
  AND2_X1 U170bar ( .A1(n794bar), .A2(n793bar), .ZN(n799bar) );
  OR2_X1 U171 ( .A1(in[94]), .A2(in[92]), .ZN(n793) );
  AND2_X1 U171bar ( .A1(inbar[94]), .A2(inbar[92]), .ZN(n793bar) );
  OR2_X1 U172 ( .A1(in_52), .A2(n792), .ZN(n794) );
  AND2_X1 U172bar ( .A1(in_52bar), .A2(n792bar), .ZN(n794bar) );
  OR2_X1 U173 ( .A1(in_70), .A2(in_67), .ZN(n792) );
  AND2_X1 U173bar ( .A1(in_70bar), .A2(in_67bar), .ZN(n792bar) );
  OR2_X1 U174 ( .A1(n791), .A2(n790), .ZN(out[2]) );
  AND2_X1 U174bar ( .A1(n791bar), .A2(n790bar), .ZN(outbar[2]) );
  OR2_X1 U175 ( .A1(n789), .A2(n788), .ZN(n790) );
  AND2_X1 U175bar ( .A1(n789bar), .A2(n788bar), .ZN(n790bar) );
  OR2_X1 U176 ( .A1(n787), .A2(n786), .ZN(n788) );
  AND2_X1 U176bar ( .A1(n787bar), .A2(n786bar), .ZN(n788bar) );
  OR2_X1 U177 ( .A1(n819), .A2(n785), .ZN(n786) );
  AND2_X1 U177bar ( .A1(n819bar), .A2(n785bar), .ZN(n786bar) );
  OR2_X1 U178 ( .A1(n784), .A2(n783), .ZN(n819) );
  AND2_X1 U178bar ( .A1(n784bar), .A2(n783bar), .ZN(n819bar) );
  OR2_X1 U179 ( .A1(n782), .A2(n781), .ZN(n783) );
  AND2_X1 U179bar ( .A1(n782bar), .A2(n781bar), .ZN(n783bar) );
  OR2_X1 U180 ( .A1(n780), .A2(n779), .ZN(n781) );
  AND2_X1 U180bar ( .A1(n780bar), .A2(n779bar), .ZN(n781bar) );
  OR2_X1 U181 ( .A1(n962), .A2(n778), .ZN(n779) );
  AND2_X1 U181bar ( .A1(n962bar), .A2(n778bar), .ZN(n779bar) );
  OR2_X1 U182 ( .A1(n777), .A2(n776), .ZN(n962) );
  AND2_X1 U182bar ( .A1(n777bar), .A2(n776bar), .ZN(n962bar) );
  OR2_X1 U183 ( .A1(n775), .A2(n774), .ZN(n776) );
  AND2_X1 U183bar ( .A1(n775bar), .A2(n774bar), .ZN(n776bar) );
  OR2_X1 U184 ( .A1(n773), .A2(n772), .ZN(n774) );
  AND2_X1 U184bar ( .A1(n773bar), .A2(n772bar), .ZN(n774bar) );
  OR2_X1 U185 ( .A1(in[131]), .A2(in[120]), .ZN(n772) );
  AND2_X1 U185bar ( .A1(inbar[131]), .A2(inbar[120]), .ZN(n772bar) );
  OR2_X1 U186 ( .A1(in[153]), .A2(in[147]), .ZN(n773) );
  AND2_X1 U186bar ( .A1(inbar[153]), .A2(inbar[147]), .ZN(n773bar) );
  OR2_X1 U187 ( .A1(n771), .A2(n770), .ZN(n775) );
  AND2_X1 U187bar ( .A1(n771bar), .A2(n770bar), .ZN(n775bar) );
  OR2_X1 U188 ( .A1(in[170]), .A2(in[156]), .ZN(n770) );
  AND2_X1 U188bar ( .A1(inbar[170]), .A2(inbar[156]), .ZN(n770bar) );
  OR2_X1 U189 ( .A1(in[223]), .A2(in[190]), .ZN(n771) );
  AND2_X1 U189bar ( .A1(inbar[223]), .A2(inbar[190]), .ZN(n771bar) );
  OR2_X1 U190 ( .A1(n769), .A2(n768), .ZN(n777) );
  AND2_X1 U190bar ( .A1(n769bar), .A2(n768bar), .ZN(n777bar) );
  OR2_X1 U191 ( .A1(n767), .A2(n766), .ZN(n768) );
  AND2_X1 U191bar ( .A1(n767bar), .A2(n766bar), .ZN(n768bar) );
  OR2_X1 U192 ( .A1(in[236]), .A2(in[230]), .ZN(n766) );
  AND2_X1 U192bar ( .A1(inbar[236]), .A2(inbar[230]), .ZN(n766bar) );
  OR2_X1 U193 ( .A1(in[85]), .A2(in[240]), .ZN(n767) );
  AND2_X1 U193bar ( .A1(inbar[85]), .A2(inbar[240]), .ZN(n767bar) );
  OR2_X1 U194 ( .A1(n765), .A2(n764), .ZN(n769) );
  AND2_X1 U194bar ( .A1(n765bar), .A2(n764bar), .ZN(n769bar) );
  OR2_X1 U195 ( .A1(in_12), .A2(in[90]), .ZN(n764) );
  AND2_X1 U195bar ( .A1(in_12bar), .A2(inbar[90]), .ZN(n764bar) );
  OR2_X1 U196 ( .A1(in_39), .A2(in_28), .ZN(n765) );
  AND2_X1 U196bar ( .A1(in_39bar), .A2(in_28bar), .ZN(n765bar) );
  OR2_X1 U197 ( .A1(in[109]), .A2(n763), .ZN(n780) );
  AND2_X1 U197bar ( .A1(inbar[109]), .A2(n763bar), .ZN(n780bar) );
  OR2_X1 U198 ( .A1(n762), .A2(n761), .ZN(n782) );
  AND2_X1 U198bar ( .A1(n762bar), .A2(n761bar), .ZN(n782bar) );
  OR2_X1 U199 ( .A1(in[138]), .A2(in[129]), .ZN(n761) );
  AND2_X1 U199bar ( .A1(inbar[138]), .A2(inbar[129]), .ZN(n761bar) );
  OR2_X1 U200 ( .A1(in[157]), .A2(n760), .ZN(n762) );
  AND2_X1 U200bar ( .A1(inbar[157]), .A2(n760bar), .ZN(n762bar) );
  OR2_X1 U201 ( .A1(in[182]), .A2(in[167]), .ZN(n760) );
  AND2_X1 U201bar ( .A1(inbar[182]), .A2(inbar[167]), .ZN(n760bar) );
  OR2_X1 U202 ( .A1(n759), .A2(n758), .ZN(n784) );
  AND2_X1 U202bar ( .A1(n759bar), .A2(n758bar), .ZN(n784bar) );
  OR2_X1 U203 ( .A1(n757), .A2(n756), .ZN(n758) );
  AND2_X1 U203bar ( .A1(n757bar), .A2(n756bar), .ZN(n758bar) );
  OR2_X1 U204 ( .A1(in[195]), .A2(in[184]), .ZN(n756) );
  AND2_X1 U204bar ( .A1(inbar[195]), .A2(inbar[184]), .ZN(n756bar) );
  OR2_X1 U205 ( .A1(in[196]), .A2(n755), .ZN(n757) );
  AND2_X1 U205bar ( .A1(inbar[196]), .A2(n755bar), .ZN(n757bar) );
  OR2_X1 U206 ( .A1(in[215]), .A2(in[209]), .ZN(n755) );
  AND2_X1 U206bar ( .A1(inbar[215]), .A2(inbar[209]), .ZN(n755bar) );
  OR2_X1 U207 ( .A1(n754), .A2(n753), .ZN(n759) );
  AND2_X1 U207bar ( .A1(n754bar), .A2(n753bar), .ZN(n759bar) );
  OR2_X1 U208 ( .A1(in[93]), .A2(in[233]), .ZN(n753) );
  AND2_X1 U208bar ( .A1(inbar[93]), .A2(inbar[233]), .ZN(n753bar) );
  OR2_X1 U209 ( .A1(in_1), .A2(n752), .ZN(n754) );
  AND2_X1 U209bar ( .A1(in_1bar), .A2(n752bar), .ZN(n754bar) );
  OR2_X1 U210 ( .A1(in_69), .A2(in_66), .ZN(n752) );
  AND2_X1 U210bar ( .A1(in_69bar), .A2(in_66bar), .ZN(n752bar) );
  OR2_X1 U211 ( .A1(n966), .A2(n751), .ZN(n787) );
  AND2_X1 U211bar ( .A1(n966bar), .A2(n751bar), .ZN(n787bar) );
  OR2_X1 U212 ( .A1(in[134]), .A2(n750), .ZN(n751) );
  AND2_X1 U212bar ( .A1(inbar[134]), .A2(n750bar), .ZN(n751bar) );
  OR2_X1 U213 ( .A1(n749), .A2(n748), .ZN(n966) );
  AND2_X1 U213bar ( .A1(n749bar), .A2(n748bar), .ZN(n966bar) );
  OR2_X1 U214 ( .A1(n747), .A2(n746), .ZN(n748) );
  AND2_X1 U214bar ( .A1(n747bar), .A2(n746bar), .ZN(n748bar) );
  OR2_X1 U215 ( .A1(n745), .A2(n744), .ZN(n746) );
  AND2_X1 U215bar ( .A1(n745bar), .A2(n744bar), .ZN(n746bar) );
  OR2_X1 U216 ( .A1(in[136]), .A2(in[121]), .ZN(n744) );
  AND2_X1 U216bar ( .A1(inbar[136]), .A2(inbar[121]), .ZN(n744bar) );
  OR2_X1 U217 ( .A1(in[186]), .A2(in[174]), .ZN(n745) );
  AND2_X1 U217bar ( .A1(inbar[186]), .A2(inbar[174]), .ZN(n745bar) );
  OR2_X1 U218 ( .A1(n743), .A2(n742), .ZN(n747) );
  AND2_X1 U218bar ( .A1(n743bar), .A2(n742bar), .ZN(n747bar) );
  OR2_X1 U219 ( .A1(in[198]), .A2(in[197]), .ZN(n742) );
  AND2_X1 U219bar ( .A1(inbar[198]), .A2(inbar[197]), .ZN(n742bar) );
  OR2_X1 U220 ( .A1(in[214]), .A2(in[199]), .ZN(n743) );
  AND2_X1 U220bar ( .A1(inbar[214]), .A2(inbar[199]), .ZN(n743bar) );
  OR2_X1 U221 ( .A1(n741), .A2(n740), .ZN(n749) );
  AND2_X1 U221bar ( .A1(n741bar), .A2(n740bar), .ZN(n749bar) );
  OR2_X1 U222 ( .A1(n739), .A2(n738), .ZN(n740) );
  AND2_X1 U222bar ( .A1(n739bar), .A2(n738bar), .ZN(n740bar) );
  OR2_X1 U223 ( .A1(in[231]), .A2(in[220]), .ZN(n738) );
  AND2_X1 U223bar ( .A1(inbar[231]), .A2(inbar[220]), .ZN(n738bar) );
  OR2_X1 U224 ( .A1(in_25), .A2(in[245]), .ZN(n739) );
  AND2_X1 U224bar ( .A1(in_25bar), .A2(inbar[245]), .ZN(n739bar) );
  OR2_X1 U225 ( .A1(n737), .A2(n736), .ZN(n741) );
  AND2_X1 U225bar ( .A1(n737bar), .A2(n736bar), .ZN(n741bar) );
  OR2_X1 U226 ( .A1(in_53), .A2(in_29), .ZN(n736) );
  AND2_X1 U226bar ( .A1(in_53bar), .A2(in_29bar), .ZN(n736bar) );
  OR2_X1 U227 ( .A1(in_79), .A2(in_74), .ZN(n737) );
  AND2_X1 U227bar ( .A1(in_79bar), .A2(in_74bar), .ZN(n737bar) );
  OR2_X1 U228 ( .A1(n735), .A2(n734), .ZN(n789) );
  AND2_X1 U228bar ( .A1(n735bar), .A2(n734bar), .ZN(n789bar) );
  OR2_X1 U229 ( .A1(in[152]), .A2(in[140]), .ZN(n734) );
  AND2_X1 U229bar ( .A1(inbar[152]), .A2(inbar[140]), .ZN(n734bar) );
  OR2_X1 U230 ( .A1(in[155]), .A2(n733), .ZN(n735) );
  AND2_X1 U230bar ( .A1(inbar[155]), .A2(n733bar), .ZN(n735bar) );
  OR2_X1 U231 ( .A1(in[166]), .A2(in[165]), .ZN(n733) );
  AND2_X1 U231bar ( .A1(inbar[166]), .A2(inbar[165]), .ZN(n733bar) );
  OR2_X1 U232 ( .A1(n732), .A2(n731), .ZN(n791) );
  AND2_X1 U232bar ( .A1(n732bar), .A2(n731bar), .ZN(n791bar) );
  OR2_X1 U233 ( .A1(n730), .A2(n729), .ZN(n731) );
  AND2_X1 U233bar ( .A1(n730bar), .A2(n729bar), .ZN(n731bar) );
  OR2_X1 U234 ( .A1(in[202]), .A2(in[185]), .ZN(n729) );
  AND2_X1 U234bar ( .A1(inbar[202]), .A2(inbar[185]), .ZN(n729bar) );
  OR2_X1 U235 ( .A1(in[211]), .A2(n728), .ZN(n730) );
  AND2_X1 U235bar ( .A1(inbar[211]), .A2(n728bar), .ZN(n730bar) );
  OR2_X1 U236 ( .A1(in[255]), .A2(in[253]), .ZN(n728) );
  AND2_X1 U236bar ( .A1(inbar[255]), .A2(inbar[253]), .ZN(n728bar) );
  OR2_X1 U237 ( .A1(n727), .A2(n726), .ZN(n732) );
  AND2_X1 U237bar ( .A1(n727bar), .A2(n726bar), .ZN(n732bar) );
  OR2_X1 U238 ( .A1(in_35), .A2(in_15), .ZN(n726) );
  AND2_X1 U238bar ( .A1(in_35bar), .A2(in_15bar), .ZN(n726bar) );
  OR2_X1 U239 ( .A1(in_36), .A2(n725), .ZN(n727) );
  AND2_X1 U239bar ( .A1(in_36bar), .A2(n725bar), .ZN(n727bar) );
  OR2_X1 U240 ( .A1(in_48), .A2(in_40), .ZN(n725) );
  AND2_X1 U240bar ( .A1(in_48bar), .A2(in_40bar), .ZN(n725bar) );
  OR2_X1 U241 ( .A1(n724), .A2(n723), .ZN(out[1]) );
  AND2_X1 U241bar ( .A1(n724bar), .A2(n723bar), .ZN(outbar[1]) );
  OR2_X1 U242 ( .A1(n722), .A2(n721), .ZN(n723) );
  AND2_X1 U242bar ( .A1(n722bar), .A2(n721bar), .ZN(n723bar) );
  OR2_X1 U243 ( .A1(n720), .A2(n719), .ZN(n721) );
  AND2_X1 U243bar ( .A1(n720bar), .A2(n719bar), .ZN(n721bar) );
  OR2_X1 U244 ( .A1(n921), .A2(n887), .ZN(n719) );
  AND2_X1 U244bar ( .A1(n921bar), .A2(n887bar), .ZN(n719bar) );
  OR2_X1 U245 ( .A1(n718), .A2(n717), .ZN(n887) );
  AND2_X1 U245bar ( .A1(n718bar), .A2(n717bar), .ZN(n887bar) );
  OR2_X1 U246 ( .A1(n716), .A2(n715), .ZN(n717) );
  AND2_X1 U246bar ( .A1(n716bar), .A2(n715bar), .ZN(n717bar) );
  OR2_X1 U247 ( .A1(n714), .A2(n713), .ZN(n715) );
  AND2_X1 U247bar ( .A1(n714bar), .A2(n713bar), .ZN(n715bar) );
  OR2_X1 U248 ( .A1(in[116]), .A2(in[110]), .ZN(n713) );
  AND2_X1 U248bar ( .A1(inbar[116]), .A2(inbar[110]), .ZN(n713bar) );
  OR2_X1 U249 ( .A1(in[133]), .A2(in[130]), .ZN(n714) );
  AND2_X1 U249bar ( .A1(inbar[133]), .A2(inbar[130]), .ZN(n714bar) );
  OR2_X1 U250 ( .A1(n712), .A2(n711), .ZN(n716) );
  AND2_X1 U250bar ( .A1(n712bar), .A2(n711bar), .ZN(n716bar) );
  OR2_X1 U251 ( .A1(in[203]), .A2(in[135]), .ZN(n711) );
  AND2_X1 U251bar ( .A1(inbar[203]), .A2(inbar[135]), .ZN(n711bar) );
  OR2_X1 U252 ( .A1(in[232]), .A2(in[223]), .ZN(n712) );
  AND2_X1 U252bar ( .A1(inbar[232]), .A2(inbar[223]), .ZN(n712bar) );
  OR2_X1 U253 ( .A1(n710), .A2(n709), .ZN(n718) );
  AND2_X1 U253bar ( .A1(n710bar), .A2(n709bar), .ZN(n718bar) );
  OR2_X1 U254 ( .A1(n708), .A2(n707), .ZN(n709) );
  AND2_X1 U254bar ( .A1(n708bar), .A2(n707bar), .ZN(n709bar) );
  OR2_X1 U255 ( .A1(in[255]), .A2(in[233]), .ZN(n707) );
  AND2_X1 U255bar ( .A1(inbar[255]), .A2(inbar[233]), .ZN(n707bar) );
  OR2_X1 U256 ( .A1(in_53), .A2(in_34), .ZN(n708) );
  AND2_X1 U256bar ( .A1(in_53bar), .A2(in_34bar), .ZN(n708bar) );
  OR2_X1 U257 ( .A1(n706), .A2(n705), .ZN(n710) );
  AND2_X1 U257bar ( .A1(n706bar), .A2(n705bar), .ZN(n710bar) );
  OR2_X1 U258 ( .A1(in_57), .A2(in_55), .ZN(n705) );
  AND2_X1 U258bar ( .A1(in_57bar), .A2(in_55bar), .ZN(n705bar) );
  OR2_X1 U259 ( .A1(in_68), .A2(in_67), .ZN(n706) );
  AND2_X1 U259bar ( .A1(in_68bar), .A2(in_67bar), .ZN(n706bar) );
  OR2_X1 U260 ( .A1(n704), .A2(n703), .ZN(n921) );
  AND2_X1 U260bar ( .A1(n704bar), .A2(n703bar), .ZN(n921bar) );
  OR2_X1 U261 ( .A1(n702), .A2(n701), .ZN(n703) );
  AND2_X1 U261bar ( .A1(n702bar), .A2(n701bar), .ZN(n703bar) );
  OR2_X1 U262 ( .A1(n700), .A2(n699), .ZN(n701) );
  AND2_X1 U262bar ( .A1(n700bar), .A2(n699bar), .ZN(n701bar) );
  OR2_X1 U263 ( .A1(n944), .A2(n872), .ZN(n699) );
  AND2_X1 U263bar ( .A1(n944bar), .A2(n872bar), .ZN(n699bar) );
  OR2_X1 U264 ( .A1(n698), .A2(n697), .ZN(n872) );
  AND2_X1 U264bar ( .A1(n698bar), .A2(n697bar), .ZN(n872bar) );
  OR2_X1 U265 ( .A1(n696), .A2(n695), .ZN(n697) );
  AND2_X1 U265bar ( .A1(n696bar), .A2(n695bar), .ZN(n697bar) );
  OR2_X1 U266 ( .A1(n694), .A2(n693), .ZN(n695) );
  AND2_X1 U266bar ( .A1(n694bar), .A2(n693bar), .ZN(n695bar) );
  OR2_X1 U267 ( .A1(in[121]), .A2(in[102]), .ZN(n693) );
  AND2_X1 U267bar ( .A1(inbar[121]), .A2(inbar[102]), .ZN(n693bar) );
  OR2_X1 U268 ( .A1(in[162]), .A2(in[161]), .ZN(n694) );
  AND2_X1 U268bar ( .A1(inbar[162]), .A2(inbar[161]), .ZN(n694bar) );
  OR2_X1 U269 ( .A1(n692), .A2(n691), .ZN(n696) );
  AND2_X1 U269bar ( .A1(n692bar), .A2(n691bar), .ZN(n696bar) );
  OR2_X1 U270 ( .A1(in[192]), .A2(in[178]), .ZN(n691) );
  AND2_X1 U270bar ( .A1(inbar[192]), .A2(inbar[178]), .ZN(n691bar) );
  OR2_X1 U271 ( .A1(in[244]), .A2(in[209]), .ZN(n692) );
  AND2_X1 U271bar ( .A1(inbar[244]), .A2(inbar[209]), .ZN(n692bar) );
  OR2_X1 U272 ( .A1(n690), .A2(n689), .ZN(n698) );
  AND2_X1 U272bar ( .A1(n690bar), .A2(n689bar), .ZN(n698bar) );
  OR2_X1 U273 ( .A1(n688), .A2(n687), .ZN(n689) );
  AND2_X1 U273bar ( .A1(n688bar), .A2(n687bar), .ZN(n689bar) );
  OR2_X1 U274 ( .A1(in[90]), .A2(in[254]), .ZN(n687) );
  AND2_X1 U274bar ( .A1(inbar[90]), .A2(inbar[254]), .ZN(n687bar) );
  OR2_X1 U275 ( .A1(in_36), .A2(in_32), .ZN(n688) );
  AND2_X1 U275bar ( .A1(in_36bar), .A2(in_32bar), .ZN(n688bar) );
  OR2_X1 U276 ( .A1(n686), .A2(n685), .ZN(n690) );
  AND2_X1 U276bar ( .A1(n686bar), .A2(n685bar), .ZN(n690bar) );
  OR2_X1 U277 ( .A1(in_62), .A2(in_37), .ZN(n685) );
  AND2_X1 U277bar ( .A1(in_62bar), .A2(in_37bar), .ZN(n685bar) );
  OR2_X1 U278 ( .A1(in_75), .A2(in_73), .ZN(n686) );
  AND2_X1 U278bar ( .A1(in_75bar), .A2(in_73bar), .ZN(n686bar) );
  OR2_X1 U279 ( .A1(n684), .A2(n683), .ZN(n944) );
  AND2_X1 U279bar ( .A1(n684bar), .A2(n683bar), .ZN(n944bar) );
  OR2_X1 U280 ( .A1(n682), .A2(n681), .ZN(n683) );
  AND2_X1 U280bar ( .A1(n682bar), .A2(n681bar), .ZN(n683bar) );
  OR2_X1 U281 ( .A1(n680), .A2(n679), .ZN(n681) );
  AND2_X1 U281bar ( .A1(n680bar), .A2(n679bar), .ZN(n681bar) );
  OR2_X1 U282 ( .A1(in[171]), .A2(in[153]), .ZN(n679) );
  AND2_X1 U282bar ( .A1(inbar[171]), .A2(inbar[153]), .ZN(n679bar) );
  OR2_X1 U283 ( .A1(in[187]), .A2(in[176]), .ZN(n680) );
  AND2_X1 U283bar ( .A1(inbar[187]), .A2(inbar[176]), .ZN(n680bar) );
  OR2_X1 U284 ( .A1(n678), .A2(n677), .ZN(n682) );
  AND2_X1 U284bar ( .A1(n678bar), .A2(n677bar), .ZN(n682bar) );
  OR2_X1 U285 ( .A1(in[245]), .A2(in[211]), .ZN(n677) );
  AND2_X1 U285bar ( .A1(inbar[245]), .A2(inbar[211]), .ZN(n677bar) );
  OR2_X1 U286 ( .A1(in[97]), .A2(in[88]), .ZN(n678) );
  AND2_X1 U286bar ( .A1(inbar[97]), .A2(inbar[88]), .ZN(n678bar) );
  OR2_X1 U287 ( .A1(n676), .A2(n675), .ZN(n684) );
  AND2_X1 U287bar ( .A1(n676bar), .A2(n675bar), .ZN(n684bar) );
  OR2_X1 U288 ( .A1(n674), .A2(n673), .ZN(n675) );
  AND2_X1 U288bar ( .A1(n674bar), .A2(n673bar), .ZN(n675bar) );
  OR2_X1 U289 ( .A1(in_10), .A2(in_0), .ZN(n673) );
  AND2_X1 U289bar ( .A1(in_10bar), .A2(in_0bar), .ZN(n673bar) );
  OR2_X1 U290 ( .A1(in_59), .A2(in_5), .ZN(n674) );
  AND2_X1 U290bar ( .A1(in_59bar), .A2(in_5bar), .ZN(n674bar) );
  OR2_X1 U291 ( .A1(n672), .A2(n671), .ZN(n676) );
  AND2_X1 U291bar ( .A1(n672bar), .A2(n671bar), .ZN(n676bar) );
  OR2_X1 U292 ( .A1(in_60), .A2(in_6), .ZN(n671) );
  AND2_X1 U292bar ( .A1(in_60bar), .A2(in_6bar), .ZN(n671bar) );
  OR2_X1 U293 ( .A1(in_77), .A2(in_69), .ZN(n672) );
  AND2_X1 U293bar ( .A1(in_77bar), .A2(in_69bar), .ZN(n672bar) );
  OR2_X1 U294 ( .A1(in[113]), .A2(n864), .ZN(n700) );
  AND2_X1 U294bar ( .A1(inbar[113]), .A2(n864bar), .ZN(n700bar) );
  OR2_X1 U295 ( .A1(n670), .A2(n669), .ZN(n864) );
  AND2_X1 U295bar ( .A1(n670bar), .A2(n669bar), .ZN(n864bar) );
  OR2_X1 U296 ( .A1(n668), .A2(n667), .ZN(n669) );
  AND2_X1 U296bar ( .A1(n668bar), .A2(n667bar), .ZN(n669bar) );
  OR2_X1 U297 ( .A1(n666), .A2(n665), .ZN(n667) );
  AND2_X1 U297bar ( .A1(n666bar), .A2(n665bar), .ZN(n667bar) );
  OR2_X1 U298 ( .A1(in[125]), .A2(in[107]), .ZN(n665) );
  AND2_X1 U298bar ( .A1(inbar[125]), .A2(inbar[107]), .ZN(n665bar) );
  OR2_X1 U299 ( .A1(in[138]), .A2(in[126]), .ZN(n666) );
  AND2_X1 U299bar ( .A1(inbar[138]), .A2(inbar[126]), .ZN(n666bar) );
  OR2_X1 U300 ( .A1(n664), .A2(n663), .ZN(n668) );
  AND2_X1 U300bar ( .A1(n664bar), .A2(n663bar), .ZN(n668bar) );
  OR2_X1 U301 ( .A1(in[189]), .A2(in[143]), .ZN(n663) );
  AND2_X1 U301bar ( .A1(inbar[189]), .A2(inbar[143]), .ZN(n663bar) );
  OR2_X1 U302 ( .A1(in[99]), .A2(in[214]), .ZN(n664) );
  AND2_X1 U302bar ( .A1(inbar[99]), .A2(inbar[214]), .ZN(n664bar) );
  OR2_X1 U303 ( .A1(n662), .A2(n661), .ZN(n670) );
  AND2_X1 U303bar ( .A1(n662bar), .A2(n661bar), .ZN(n670bar) );
  OR2_X1 U304 ( .A1(n660), .A2(n659), .ZN(n661) );
  AND2_X1 U304bar ( .A1(n660bar), .A2(n659bar), .ZN(n661bar) );
  OR2_X1 U305 ( .A1(in_15), .A2(in_12), .ZN(n659) );
  AND2_X1 U305bar ( .A1(in_15bar), .A2(in_12bar), .ZN(n659bar) );
  OR2_X1 U306 ( .A1(in_20), .A2(in_2), .ZN(n660) );
  AND2_X1 U306bar ( .A1(in_20bar), .A2(in_2bar), .ZN(n660bar) );
  OR2_X1 U307 ( .A1(n658), .A2(n657), .ZN(n662) );
  AND2_X1 U307bar ( .A1(n658bar), .A2(n657bar), .ZN(n662bar) );
  OR2_X1 U308 ( .A1(in_30), .A2(in_3), .ZN(n657) );
  AND2_X1 U308bar ( .A1(in_30bar), .A2(in_3bar), .ZN(n657bar) );
  OR2_X1 U309 ( .A1(in_4), .A2(in_38), .ZN(n658) );
  AND2_X1 U309bar ( .A1(in_4bar), .A2(in_38bar), .ZN(n658bar) );
  OR2_X1 U310 ( .A1(n656), .A2(n655), .ZN(n702) );
  AND2_X1 U310bar ( .A1(n656bar), .A2(n655bar), .ZN(n702bar) );
  OR2_X1 U311 ( .A1(in[148]), .A2(in[137]), .ZN(n655) );
  AND2_X1 U311bar ( .A1(inbar[148]), .A2(inbar[137]), .ZN(n655bar) );
  OR2_X1 U312 ( .A1(in[149]), .A2(n654), .ZN(n656) );
  AND2_X1 U312bar ( .A1(inbar[149]), .A2(n654bar), .ZN(n656bar) );
  OR2_X1 U313 ( .A1(in[195]), .A2(in[190]), .ZN(n654) );
  AND2_X1 U313bar ( .A1(inbar[195]), .A2(inbar[190]), .ZN(n654bar) );
  OR2_X1 U314 ( .A1(n653), .A2(n652), .ZN(n704) );
  AND2_X1 U314bar ( .A1(n653bar), .A2(n652bar), .ZN(n704bar) );
  OR2_X1 U315 ( .A1(n651), .A2(n650), .ZN(n652) );
  AND2_X1 U315bar ( .A1(n651bar), .A2(n650bar), .ZN(n652bar) );
  OR2_X1 U316 ( .A1(in[98]), .A2(in[197]), .ZN(n650) );
  AND2_X1 U316bar ( .A1(inbar[98]), .A2(inbar[197]), .ZN(n650bar) );
  OR2_X1 U317 ( .A1(in_11), .A2(n649), .ZN(n651) );
  AND2_X1 U317bar ( .A1(in_11bar), .A2(n649bar), .ZN(n651bar) );
  OR2_X1 U318 ( .A1(in_26), .A2(in_14), .ZN(n649) );
  AND2_X1 U318bar ( .A1(in_26bar), .A2(in_14bar), .ZN(n649bar) );
  OR2_X1 U319 ( .A1(n648), .A2(n647), .ZN(n653) );
  AND2_X1 U319bar ( .A1(n648bar), .A2(n647bar), .ZN(n653bar) );
  OR2_X1 U320 ( .A1(in_35), .A2(in_27), .ZN(n647) );
  AND2_X1 U320bar ( .A1(in_35bar), .A2(in_27bar), .ZN(n647bar) );
  OR2_X1 U321 ( .A1(in_50), .A2(n646), .ZN(n648) );
  AND2_X1 U321bar ( .A1(in_50bar), .A2(n646bar), .ZN(n648bar) );
  OR2_X1 U322 ( .A1(in_78), .A2(in_61), .ZN(n646) );
  AND2_X1 U322bar ( .A1(in_78bar), .A2(in_61bar), .ZN(n646bar) );
  OR2_X1 U323 ( .A1(n942), .A2(n645), .ZN(n720) );
  AND2_X1 U323bar ( .A1(n942bar), .A2(n645bar), .ZN(n720bar) );
  OR2_X1 U324 ( .A1(in[106]), .A2(n863), .ZN(n645) );
  AND2_X1 U324bar ( .A1(inbar[106]), .A2(n863bar), .ZN(n645bar) );
  OR2_X1 U325 ( .A1(n644), .A2(n643), .ZN(n863) );
  AND2_X1 U325bar ( .A1(n644bar), .A2(n643bar), .ZN(n863bar) );
  OR2_X1 U326 ( .A1(n642), .A2(n641), .ZN(n643) );
  AND2_X1 U326bar ( .A1(n642bar), .A2(n641bar), .ZN(n643bar) );
  OR2_X1 U327 ( .A1(n640), .A2(n639), .ZN(n641) );
  AND2_X1 U327bar ( .A1(n640bar), .A2(n639bar), .ZN(n641bar) );
  OR2_X1 U328 ( .A1(in[127]), .A2(in[122]), .ZN(n639) );
  AND2_X1 U328bar ( .A1(inbar[127]), .A2(inbar[122]), .ZN(n639bar) );
  OR2_X1 U329 ( .A1(in[156]), .A2(in[132]), .ZN(n640) );
  AND2_X1 U329bar ( .A1(inbar[156]), .A2(inbar[132]), .ZN(n640bar) );
  OR2_X1 U330 ( .A1(n638), .A2(n637), .ZN(n642) );
  AND2_X1 U330bar ( .A1(n638bar), .A2(n637bar), .ZN(n642bar) );
  OR2_X1 U331 ( .A1(in[159]), .A2(in[157]), .ZN(n637) );
  AND2_X1 U331bar ( .A1(inbar[159]), .A2(inbar[157]), .ZN(n637bar) );
  OR2_X1 U332 ( .A1(in[185]), .A2(in[169]), .ZN(n638) );
  AND2_X1 U332bar ( .A1(inbar[185]), .A2(inbar[169]), .ZN(n638bar) );
  OR2_X1 U333 ( .A1(n636), .A2(n635), .ZN(n644) );
  AND2_X1 U333bar ( .A1(n636bar), .A2(n635bar), .ZN(n644bar) );
  OR2_X1 U334 ( .A1(n634), .A2(n633), .ZN(n635) );
  AND2_X1 U334bar ( .A1(n634bar), .A2(n633bar), .ZN(n635bar) );
  OR2_X1 U335 ( .A1(in[239]), .A2(in[218]), .ZN(n633) );
  AND2_X1 U335bar ( .A1(inbar[239]), .A2(inbar[218]), .ZN(n633bar) );
  OR2_X1 U336 ( .A1(in_13), .A2(in[87]), .ZN(n634) );
  AND2_X1 U336bar ( .A1(in_13bar), .A2(inbar[87]), .ZN(n634bar) );
  OR2_X1 U337 ( .A1(n632), .A2(n631), .ZN(n636) );
  AND2_X1 U337bar ( .A1(n632bar), .A2(n631bar), .ZN(n636bar) );
  OR2_X1 U338 ( .A1(in_72), .A2(in_70), .ZN(n631) );
  AND2_X1 U338bar ( .A1(in_72bar), .A2(in_70bar), .ZN(n631bar) );
  OR2_X1 U339 ( .A1(in_80), .A2(in_74), .ZN(n632) );
  AND2_X1 U339bar ( .A1(in_80bar), .A2(in_74bar), .ZN(n632bar) );
  OR2_X1 U340 ( .A1(n630), .A2(n629), .ZN(n942) );
  AND2_X1 U340bar ( .A1(n630bar), .A2(n629bar), .ZN(n942bar) );
  OR2_X1 U341 ( .A1(n628), .A2(n627), .ZN(n629) );
  AND2_X1 U341bar ( .A1(n628bar), .A2(n627bar), .ZN(n629bar) );
  OR2_X1 U342 ( .A1(n626), .A2(n625), .ZN(n627) );
  AND2_X1 U342bar ( .A1(n626bar), .A2(n625bar), .ZN(n627bar) );
  OR2_X1 U343 ( .A1(in[146]), .A2(in[100]), .ZN(n625) );
  AND2_X1 U343bar ( .A1(inbar[146]), .A2(inbar[100]), .ZN(n625bar) );
  OR2_X1 U344 ( .A1(in[168]), .A2(in[152]), .ZN(n626) );
  AND2_X1 U344bar ( .A1(inbar[168]), .A2(inbar[152]), .ZN(n626bar) );
  OR2_X1 U345 ( .A1(n624), .A2(n623), .ZN(n628) );
  AND2_X1 U345bar ( .A1(n624bar), .A2(n623bar), .ZN(n628bar) );
  OR2_X1 U346 ( .A1(in[199]), .A2(in[182]), .ZN(n623) );
  AND2_X1 U346bar ( .A1(inbar[199]), .A2(inbar[182]), .ZN(n623bar) );
  OR2_X1 U347 ( .A1(in[236]), .A2(in[204]), .ZN(n624) );
  AND2_X1 U347bar ( .A1(inbar[236]), .A2(inbar[204]), .ZN(n624bar) );
  OR2_X1 U348 ( .A1(n622), .A2(n621), .ZN(n630) );
  AND2_X1 U348bar ( .A1(n622bar), .A2(n621bar), .ZN(n630bar) );
  OR2_X1 U349 ( .A1(n620), .A2(n619), .ZN(n621) );
  AND2_X1 U349bar ( .A1(n620bar), .A2(n619bar), .ZN(n621bar) );
  OR2_X1 U350 ( .A1(in[89]), .A2(in[246]), .ZN(n619) );
  AND2_X1 U350bar ( .A1(inbar[89]), .A2(inbar[246]), .ZN(n619bar) );
  OR2_X1 U351 ( .A1(in[95]), .A2(in[92]), .ZN(n620) );
  AND2_X1 U351bar ( .A1(inbar[95]), .A2(inbar[92]), .ZN(n620bar) );
  OR2_X1 U352 ( .A1(n618), .A2(n617), .ZN(n622) );
  AND2_X1 U352bar ( .A1(n618bar), .A2(n617bar), .ZN(n622bar) );
  OR2_X1 U353 ( .A1(in_22), .A2(in_16), .ZN(n617) );
  AND2_X1 U353bar ( .A1(in_22bar), .A2(in_16bar), .ZN(n617bar) );
  OR2_X1 U354 ( .A1(in_51), .A2(in_49), .ZN(n618) );
  AND2_X1 U354bar ( .A1(in_51bar), .A2(in_49bar), .ZN(n618bar) );
  OR2_X1 U355 ( .A1(n616), .A2(n615), .ZN(n722) );
  AND2_X1 U355bar ( .A1(n616bar), .A2(n615bar), .ZN(n722bar) );
  OR2_X1 U356 ( .A1(in[158]), .A2(in[115]), .ZN(n615) );
  AND2_X1 U356bar ( .A1(inbar[158]), .A2(inbar[115]), .ZN(n615bar) );
  OR2_X1 U357 ( .A1(in[163]), .A2(n614), .ZN(n616) );
  AND2_X1 U357bar ( .A1(inbar[163]), .A2(n614bar), .ZN(n616bar) );
  OR2_X1 U358 ( .A1(in[206]), .A2(in[165]), .ZN(n614) );
  AND2_X1 U358bar ( .A1(inbar[206]), .A2(inbar[165]), .ZN(n614bar) );
  OR2_X1 U359 ( .A1(n613), .A2(n612), .ZN(n724) );
  AND2_X1 U359bar ( .A1(n613bar), .A2(n612bar), .ZN(n724bar) );
  OR2_X1 U360 ( .A1(n611), .A2(n610), .ZN(n612) );
  AND2_X1 U360bar ( .A1(n611bar), .A2(n610bar), .ZN(n612bar) );
  OR2_X1 U361 ( .A1(in[213]), .A2(in[207]), .ZN(n610) );
  AND2_X1 U361bar ( .A1(inbar[213]), .A2(inbar[207]), .ZN(n610bar) );
  OR2_X1 U362 ( .A1(in[215]), .A2(n609), .ZN(n611) );
  AND2_X1 U362bar ( .A1(inbar[215]), .A2(n609bar), .ZN(n611bar) );
  OR2_X1 U363 ( .A1(in[230]), .A2(in[220]), .ZN(n609) );
  AND2_X1 U363bar ( .A1(inbar[230]), .A2(inbar[220]), .ZN(n609bar) );
  OR2_X1 U364 ( .A1(n608), .A2(n607), .ZN(n613) );
  AND2_X1 U364bar ( .A1(n608bar), .A2(n607bar), .ZN(n613bar) );
  OR2_X1 U365 ( .A1(in[251]), .A2(in[234]), .ZN(n607) );
  AND2_X1 U365bar ( .A1(inbar[251]), .A2(inbar[234]), .ZN(n607bar) );
  OR2_X1 U366 ( .A1(in_17), .A2(n606), .ZN(n608) );
  AND2_X1 U366bar ( .A1(in_17bar), .A2(n606bar), .ZN(n608bar) );
  OR2_X1 U367 ( .A1(in_65), .A2(in_56), .ZN(n606) );
  AND2_X1 U367bar ( .A1(in_65bar), .A2(in_56bar), .ZN(n606bar) );
  OR2_X1 U368 ( .A1(n605), .A2(n604), .ZN(out[0]) );
  AND2_X1 U368bar ( .A1(n605bar), .A2(n604bar), .ZN(outbar[0]) );
  OR2_X1 U369 ( .A1(n603), .A2(n602), .ZN(n604) );
  AND2_X1 U369bar ( .A1(n603bar), .A2(n602bar), .ZN(n604bar) );
  OR2_X1 U370 ( .A1(n601), .A2(n600), .ZN(n602) );
  AND2_X1 U370bar ( .A1(n601bar), .A2(n600bar), .ZN(n602bar) );
  OR2_X1 U371 ( .A1(n820), .A2(n785), .ZN(n600) );
  AND2_X1 U371bar ( .A1(n820bar), .A2(n785bar), .ZN(n600bar) );
  OR2_X1 U372 ( .A1(n599), .A2(n598), .ZN(n785) );
  AND2_X1 U372bar ( .A1(n599bar), .A2(n598bar), .ZN(n785bar) );
  OR2_X1 U373 ( .A1(n597), .A2(n596), .ZN(n598) );
  AND2_X1 U373bar ( .A1(n597bar), .A2(n596bar), .ZN(n598bar) );
  OR2_X1 U374 ( .A1(n595), .A2(n594), .ZN(n596) );
  AND2_X1 U374bar ( .A1(n595bar), .A2(n594bar), .ZN(n596bar) );
  OR2_X1 U375 ( .A1(in[135]), .A2(in[104]), .ZN(n594) );
  AND2_X1 U375bar ( .A1(inbar[135]), .A2(inbar[104]), .ZN(n594bar) );
  OR2_X1 U376 ( .A1(in[188]), .A2(in[178]), .ZN(n595) );
  AND2_X1 U376bar ( .A1(inbar[188]), .A2(inbar[178]), .ZN(n595bar) );
  OR2_X1 U377 ( .A1(n593), .A2(n592), .ZN(n597) );
  AND2_X1 U377bar ( .A1(n593bar), .A2(n592bar), .ZN(n597bar) );
  OR2_X1 U378 ( .A1(in[217]), .A2(in[194]), .ZN(n592) );
  AND2_X1 U378bar ( .A1(inbar[217]), .A2(inbar[194]), .ZN(n592bar) );
  OR2_X1 U379 ( .A1(in[237]), .A2(in[218]), .ZN(n593) );
  AND2_X1 U379bar ( .A1(inbar[237]), .A2(inbar[218]), .ZN(n593bar) );
  OR2_X1 U380 ( .A1(n591), .A2(n590), .ZN(n599) );
  AND2_X1 U380bar ( .A1(n591bar), .A2(n590bar), .ZN(n599bar) );
  OR2_X1 U381 ( .A1(n589), .A2(n588), .ZN(n590) );
  AND2_X1 U381bar ( .A1(n589bar), .A2(n588bar), .ZN(n590bar) );
  OR2_X1 U382 ( .A1(in_2), .A2(in_10), .ZN(n588) );
  AND2_X1 U382bar ( .A1(in_2bar), .A2(in_10bar), .ZN(n588bar) );
  OR2_X1 U383 ( .A1(in_47), .A2(in_22), .ZN(n589) );
  AND2_X1 U383bar ( .A1(in_47bar), .A2(in_22bar), .ZN(n589bar) );
  OR2_X1 U384 ( .A1(n587), .A2(n586), .ZN(n591) );
  AND2_X1 U384bar ( .A1(n587bar), .A2(n586bar), .ZN(n591bar) );
  OR2_X1 U385 ( .A1(in_56), .A2(in_54), .ZN(n586) );
  AND2_X1 U385bar ( .A1(in_56bar), .A2(in_54bar), .ZN(n586bar) );
  OR2_X1 U386 ( .A1(in_63), .A2(in_61), .ZN(n587) );
  AND2_X1 U386bar ( .A1(in_63bar), .A2(in_61bar), .ZN(n587bar) );
  OR2_X1 U387 ( .A1(n585), .A2(n584), .ZN(n820) );
  AND2_X1 U387bar ( .A1(n585bar), .A2(n584bar), .ZN(n820bar) );
  OR2_X1 U388 ( .A1(n583), .A2(n582), .ZN(n584) );
  AND2_X1 U388bar ( .A1(n583bar), .A2(n582bar), .ZN(n584bar) );
  OR2_X1 U389 ( .A1(n581), .A2(n580), .ZN(n582) );
  AND2_X1 U389bar ( .A1(n581bar), .A2(n580bar), .ZN(n582bar) );
  OR2_X1 U390 ( .A1(in[158]), .A2(in[142]), .ZN(n580) );
  AND2_X1 U390bar ( .A1(inbar[158]), .A2(inbar[142]), .ZN(n580bar) );
  OR2_X1 U391 ( .A1(in[175]), .A2(in[164]), .ZN(n581) );
  AND2_X1 U391bar ( .A1(inbar[175]), .A2(inbar[164]), .ZN(n581bar) );
  OR2_X1 U392 ( .A1(n579), .A2(n578), .ZN(n583) );
  AND2_X1 U392bar ( .A1(n579bar), .A2(n578bar), .ZN(n583bar) );
  OR2_X1 U393 ( .A1(in[228]), .A2(in[204]), .ZN(n578) );
  AND2_X1 U393bar ( .A1(inbar[228]), .A2(inbar[204]), .ZN(n578bar) );
  OR2_X1 U394 ( .A1(in[91]), .A2(in[87]), .ZN(n579) );
  AND2_X1 U394bar ( .A1(inbar[91]), .A2(inbar[87]), .ZN(n579bar) );
  OR2_X1 U395 ( .A1(n577), .A2(n576), .ZN(n585) );
  AND2_X1 U395bar ( .A1(n577bar), .A2(n576bar), .ZN(n585bar) );
  OR2_X1 U396 ( .A1(n575), .A2(n574), .ZN(n576) );
  AND2_X1 U396bar ( .A1(n575bar), .A2(n574bar), .ZN(n576bar) );
  OR2_X1 U397 ( .A1(in_21), .A2(in_11), .ZN(n574) );
  AND2_X1 U397bar ( .A1(in_21bar), .A2(in_11bar), .ZN(n574bar) );
  OR2_X1 U398 ( .A1(in_5), .A2(in_3), .ZN(n575) );
  AND2_X1 U398bar ( .A1(in_5bar), .A2(in_3bar), .ZN(n575bar) );
  OR2_X1 U399 ( .A1(n573), .A2(n572), .ZN(n577) );
  AND2_X1 U399bar ( .A1(n573bar), .A2(n572bar), .ZN(n577bar) );
  OR2_X1 U400 ( .A1(in_68), .A2(in_64), .ZN(n572) );
  AND2_X1 U400bar ( .A1(in_68bar), .A2(in_64bar), .ZN(n572bar) );
  OR2_X1 U401 ( .A1(in_76), .A2(in_73), .ZN(n573) );
  AND2_X1 U401bar ( .A1(in_76bar), .A2(in_73bar), .ZN(n573bar) );
  OR2_X1 U402 ( .A1(n778), .A2(n571), .ZN(n601) );
  AND2_X1 U402bar ( .A1(n778bar), .A2(n571bar), .ZN(n601bar) );
  OR2_X1 U403 ( .A1(in[100]), .A2(n965), .ZN(n571) );
  AND2_X1 U403bar ( .A1(inbar[100]), .A2(n965bar), .ZN(n571bar) );
  OR2_X1 U404 ( .A1(n570), .A2(n569), .ZN(n965) );
  AND2_X1 U404bar ( .A1(n570bar), .A2(n569bar), .ZN(n965bar) );
  OR2_X1 U405 ( .A1(n568), .A2(n567), .ZN(n569) );
  AND2_X1 U405bar ( .A1(n568bar), .A2(n567bar), .ZN(n569bar) );
  OR2_X1 U406 ( .A1(n566), .A2(n565), .ZN(n567) );
  AND2_X1 U406bar ( .A1(n566bar), .A2(n565bar), .ZN(n567bar) );
  OR2_X1 U407 ( .A1(n817), .A2(n750), .ZN(n565) );
  AND2_X1 U407bar ( .A1(n817bar), .A2(n750bar), .ZN(n565bar) );
  OR2_X1 U408 ( .A1(n564), .A2(n563), .ZN(n750) );
  AND2_X1 U408bar ( .A1(n564bar), .A2(n563bar), .ZN(n750bar) );
  OR2_X1 U409 ( .A1(n562), .A2(n561), .ZN(n563) );
  AND2_X1 U409bar ( .A1(n562bar), .A2(n561bar), .ZN(n563bar) );
  OR2_X1 U410 ( .A1(n560), .A2(n559), .ZN(n561) );
  AND2_X1 U410bar ( .A1(n560bar), .A2(n559bar), .ZN(n561bar) );
  OR2_X1 U411 ( .A1(in[119]), .A2(in[103]), .ZN(n559) );
  AND2_X1 U411bar ( .A1(inbar[119]), .A2(inbar[103]), .ZN(n559bar) );
  OR2_X1 U412 ( .A1(in[137]), .A2(in[133]), .ZN(n560) );
  AND2_X1 U412bar ( .A1(inbar[137]), .A2(inbar[133]), .ZN(n560bar) );
  OR2_X1 U413 ( .A1(n558), .A2(n557), .ZN(n562) );
  AND2_X1 U413bar ( .A1(n558bar), .A2(n557bar), .ZN(n562bar) );
  OR2_X1 U414 ( .A1(in[176]), .A2(in[173]), .ZN(n557) );
  AND2_X1 U414bar ( .A1(inbar[176]), .A2(inbar[173]), .ZN(n557bar) );
  OR2_X1 U415 ( .A1(in[210]), .A2(in[181]), .ZN(n558) );
  AND2_X1 U415bar ( .A1(inbar[210]), .A2(inbar[181]), .ZN(n558bar) );
  OR2_X1 U416 ( .A1(n556), .A2(n555), .ZN(n564) );
  AND2_X1 U416bar ( .A1(n556bar), .A2(n555bar), .ZN(n564bar) );
  OR2_X1 U417 ( .A1(n554), .A2(n553), .ZN(n555) );
  AND2_X1 U417bar ( .A1(n554bar), .A2(n553bar), .ZN(n555bar) );
  OR2_X1 U418 ( .A1(in_13), .A2(in[234]), .ZN(n553) );
  AND2_X1 U418bar ( .A1(in_13bar), .A2(inbar[234]), .ZN(n553bar) );
  OR2_X1 U419 ( .A1(in_38), .A2(in_32), .ZN(n554) );
  AND2_X1 U419bar ( .A1(in_38bar), .A2(in_32bar), .ZN(n554bar) );
  OR2_X1 U420 ( .A1(n552), .A2(n551), .ZN(n556) );
  AND2_X1 U420bar ( .A1(n552bar), .A2(n551bar), .ZN(n556bar) );
  OR2_X1 U421 ( .A1(in_42), .A2(in_41), .ZN(n551) );
  AND2_X1 U421bar ( .A1(in_42bar), .A2(in_41bar), .ZN(n551bar) );
  OR2_X1 U422 ( .A1(in_7), .A2(in_49), .ZN(n552) );
  AND2_X1 U422bar ( .A1(in_7bar), .A2(in_49bar), .ZN(n552bar) );
  OR2_X1 U423 ( .A1(n550), .A2(n549), .ZN(n817) );
  AND2_X1 U423bar ( .A1(n550bar), .A2(n549bar), .ZN(n817bar) );
  OR2_X1 U424 ( .A1(n548), .A2(n547), .ZN(n549) );
  AND2_X1 U424bar ( .A1(n548bar), .A2(n547bar), .ZN(n549bar) );
  OR2_X1 U425 ( .A1(n546), .A2(n545), .ZN(n547) );
  AND2_X1 U425bar ( .A1(n546bar), .A2(n545bar), .ZN(n547bar) );
  OR2_X1 U426 ( .A1(in[159]), .A2(in[105]), .ZN(n545) );
  AND2_X1 U426bar ( .A1(inbar[159]), .A2(inbar[105]), .ZN(n545bar) );
  OR2_X1 U427 ( .A1(in[206]), .A2(in[183]), .ZN(n546) );
  AND2_X1 U427bar ( .A1(inbar[206]), .A2(inbar[183]), .ZN(n546bar) );
  OR2_X1 U428 ( .A1(n544), .A2(n543), .ZN(n548) );
  AND2_X1 U428bar ( .A1(n544bar), .A2(n543bar), .ZN(n548bar) );
  OR2_X1 U429 ( .A1(in[229]), .A2(in[219]), .ZN(n543) );
  AND2_X1 U429bar ( .A1(inbar[229]), .A2(inbar[219]), .ZN(n543bar) );
  OR2_X1 U430 ( .A1(in[235]), .A2(in[232]), .ZN(n544) );
  AND2_X1 U430bar ( .A1(inbar[235]), .A2(inbar[232]), .ZN(n544bar) );
  OR2_X1 U431 ( .A1(n542), .A2(n541), .ZN(n550) );
  AND2_X1 U431bar ( .A1(n542bar), .A2(n541bar), .ZN(n550bar) );
  OR2_X1 U432 ( .A1(n540), .A2(n539), .ZN(n541) );
  AND2_X1 U432bar ( .A1(n540bar), .A2(n539bar), .ZN(n541bar) );
  OR2_X1 U433 ( .A1(in[249]), .A2(in[242]), .ZN(n539) );
  AND2_X1 U433bar ( .A1(inbar[249]), .A2(inbar[242]), .ZN(n539bar) );
  OR2_X1 U434 ( .A1(in[89]), .A2(in[254]), .ZN(n540) );
  AND2_X1 U434bar ( .A1(inbar[89]), .A2(inbar[254]), .ZN(n540bar) );
  OR2_X1 U435 ( .A1(n538), .A2(n537), .ZN(n542) );
  AND2_X1 U435bar ( .A1(n538bar), .A2(n537bar), .ZN(n542bar) );
  OR2_X1 U436 ( .A1(in_14), .A2(in[99]), .ZN(n537) );
  AND2_X1 U436bar ( .A1(in_14bar), .A2(inbar[99]), .ZN(n537bar) );
  OR2_X1 U437 ( .A1(in_60), .A2(in_18), .ZN(n538) );
  AND2_X1 U437bar ( .A1(in_60bar), .A2(in_18bar), .ZN(n538bar) );
  OR2_X1 U438 ( .A1(in[113]), .A2(n763), .ZN(n566) );
  AND2_X1 U438bar ( .A1(inbar[113]), .A2(n763bar), .ZN(n566bar) );
  OR2_X1 U439 ( .A1(n536), .A2(n535), .ZN(n763) );
  AND2_X1 U439bar ( .A1(n536bar), .A2(n535bar), .ZN(n763bar) );
  OR2_X1 U440 ( .A1(n534), .A2(n533), .ZN(n535) );
  AND2_X1 U440bar ( .A1(n534bar), .A2(n533bar), .ZN(n535bar) );
  OR2_X1 U441 ( .A1(n532), .A2(n531), .ZN(n533) );
  AND2_X1 U441bar ( .A1(n532bar), .A2(n531bar), .ZN(n533bar) );
  OR2_X1 U442 ( .A1(in[115]), .A2(in[110]), .ZN(n531) );
  AND2_X1 U442bar ( .A1(inbar[115]), .A2(inbar[110]), .ZN(n531bar) );
  OR2_X1 U443 ( .A1(in[125]), .A2(in[117]), .ZN(n532) );
  AND2_X1 U443bar ( .A1(inbar[125]), .A2(inbar[117]), .ZN(n532bar) );
  OR2_X1 U444 ( .A1(n530), .A2(n529), .ZN(n534) );
  AND2_X1 U444bar ( .A1(n530bar), .A2(n529bar), .ZN(n534bar) );
  OR2_X1 U445 ( .A1(in[180]), .A2(in[128]), .ZN(n529) );
  AND2_X1 U445bar ( .A1(inbar[180]), .A2(inbar[128]), .ZN(n529bar) );
  OR2_X1 U446 ( .A1(in[205]), .A2(in[201]), .ZN(n530) );
  AND2_X1 U446bar ( .A1(inbar[205]), .A2(inbar[201]), .ZN(n530bar) );
  OR2_X1 U447 ( .A1(n528), .A2(n527), .ZN(n536) );
  AND2_X1 U447bar ( .A1(n528bar), .A2(n527bar), .ZN(n536bar) );
  OR2_X1 U448 ( .A1(n526), .A2(n525), .ZN(n527) );
  AND2_X1 U448bar ( .A1(n526bar), .A2(n525bar), .ZN(n527bar) );
  OR2_X1 U449 ( .A1(in[244]), .A2(in[239]), .ZN(n525) );
  AND2_X1 U449bar ( .A1(inbar[244]), .A2(inbar[239]), .ZN(n525bar) );
  OR2_X1 U450 ( .A1(in[95]), .A2(in[83]), .ZN(n526) );
  AND2_X1 U450bar ( .A1(inbar[95]), .A2(inbar[83]), .ZN(n526bar) );
  OR2_X1 U451 ( .A1(n524), .A2(n523), .ZN(n528) );
  AND2_X1 U451bar ( .A1(n524bar), .A2(n523bar), .ZN(n528bar) );
  OR2_X1 U452 ( .A1(in_24), .A2(in[97]), .ZN(n523) );
  AND2_X1 U452bar ( .A1(in_24bar), .A2(inbar[97]), .ZN(n523bar) );
  OR2_X1 U453 ( .A1(in_33), .A2(in_27), .ZN(n524) );
  AND2_X1 U453bar ( .A1(in_33bar), .A2(in_27bar), .ZN(n524bar) );
  OR2_X1 U454 ( .A1(n522), .A2(n521), .ZN(n568) );
  AND2_X1 U454bar ( .A1(n522bar), .A2(n521bar), .ZN(n568bar) );
  OR2_X1 U455 ( .A1(in[145]), .A2(in[126]), .ZN(n521) );
  AND2_X1 U455bar ( .A1(inbar[145]), .A2(inbar[126]), .ZN(n521bar) );
  OR2_X1 U456 ( .A1(in[169]), .A2(n520), .ZN(n522) );
  AND2_X1 U456bar ( .A1(inbar[169]), .A2(n520bar), .ZN(n522bar) );
  OR2_X1 U457 ( .A1(in[221]), .A2(in[172]), .ZN(n520) );
  AND2_X1 U457bar ( .A1(inbar[221]), .A2(inbar[172]), .ZN(n520bar) );
  OR2_X1 U458 ( .A1(n519), .A2(n518), .ZN(n570) );
  AND2_X1 U458bar ( .A1(n519bar), .A2(n518bar), .ZN(n570bar) );
  OR2_X1 U459 ( .A1(n517), .A2(n516), .ZN(n518) );
  AND2_X1 U459bar ( .A1(n517bar), .A2(n516bar), .ZN(n518bar) );
  OR2_X1 U460 ( .A1(in[241]), .A2(in[224]), .ZN(n516) );
  AND2_X1 U460bar ( .A1(inbar[241]), .A2(inbar[224]), .ZN(n516bar) );
  OR2_X1 U461 ( .A1(in[86]), .A2(n515), .ZN(n517) );
  AND2_X1 U461bar ( .A1(inbar[86]), .A2(n515bar), .ZN(n517bar) );
  OR2_X1 U462 ( .A1(in_43), .A2(in_34), .ZN(n515) );
  AND2_X1 U462bar ( .A1(in_43bar), .A2(in_34bar), .ZN(n515bar) );
  OR2_X1 U463 ( .A1(n514), .A2(n513), .ZN(n519) );
  AND2_X1 U463bar ( .A1(n514bar), .A2(n513bar), .ZN(n519bar) );
  OR2_X1 U464 ( .A1(in_65), .A2(in_51), .ZN(n513) );
  AND2_X1 U464bar ( .A1(in_65bar), .A2(in_51bar), .ZN(n513bar) );
  OR2_X1 U465 ( .A1(in_75), .A2(n512), .ZN(n514) );
  AND2_X1 U465bar ( .A1(in_75bar), .A2(n512bar), .ZN(n514bar) );
  OR2_X1 U466 ( .A1(in_81), .A2(in_77), .ZN(n512) );
  AND2_X1 U466bar ( .A1(in_81bar), .A2(in_77bar), .ZN(n512bar) );
  OR2_X1 U467 ( .A1(n511), .A2(n510), .ZN(n778) );
  AND2_X1 U467bar ( .A1(n511bar), .A2(n510bar), .ZN(n778bar) );
  OR2_X1 U468 ( .A1(n509), .A2(n508), .ZN(n510) );
  AND2_X1 U468bar ( .A1(n509bar), .A2(n508bar), .ZN(n510bar) );
  OR2_X1 U469 ( .A1(n507), .A2(n506), .ZN(n508) );
  AND2_X1 U469bar ( .A1(n507bar), .A2(n506bar), .ZN(n508bar) );
  OR2_X1 U470 ( .A1(in[107]), .A2(in[101]), .ZN(n506) );
  AND2_X1 U470bar ( .A1(inbar[107]), .A2(inbar[101]), .ZN(n506bar) );
  OR2_X1 U471 ( .A1(in[139]), .A2(in[132]), .ZN(n507) );
  AND2_X1 U471bar ( .A1(inbar[139]), .A2(inbar[132]), .ZN(n507bar) );
  OR2_X1 U472 ( .A1(n505), .A2(n504), .ZN(n509) );
  AND2_X1 U472bar ( .A1(n505bar), .A2(n504bar), .ZN(n509bar) );
  OR2_X1 U473 ( .A1(in[146]), .A2(in[141]), .ZN(n504) );
  AND2_X1 U473bar ( .A1(inbar[146]), .A2(inbar[141]), .ZN(n504bar) );
  OR2_X1 U474 ( .A1(in[203]), .A2(in[179]), .ZN(n505) );
  AND2_X1 U474bar ( .A1(inbar[203]), .A2(inbar[179]), .ZN(n505bar) );
  OR2_X1 U475 ( .A1(n503), .A2(n502), .ZN(n511) );
  AND2_X1 U475bar ( .A1(n503bar), .A2(n502bar), .ZN(n511bar) );
  OR2_X1 U476 ( .A1(n501), .A2(n500), .ZN(n502) );
  AND2_X1 U476bar ( .A1(n501bar), .A2(n500bar), .ZN(n502bar) );
  OR2_X1 U477 ( .A1(in[243]), .A2(in[222]), .ZN(n500) );
  AND2_X1 U477bar ( .A1(inbar[243]), .A2(inbar[222]), .ZN(n500bar) );
  OR2_X1 U478 ( .A1(in[251]), .A2(in[250]), .ZN(n501) );
  AND2_X1 U478bar ( .A1(inbar[251]), .A2(inbar[250]), .ZN(n501bar) );
  OR2_X1 U479 ( .A1(n499), .A2(n498), .ZN(n503) );
  AND2_X1 U479bar ( .A1(n499bar), .A2(n498bar), .ZN(n503bar) );
  OR2_X1 U480 ( .A1(in_37), .A2(in_19), .ZN(n498) );
  AND2_X1 U480bar ( .A1(in_37bar), .A2(in_19bar), .ZN(n498bar) );
  OR2_X1 U481 ( .A1(in_78), .A2(in_6), .ZN(n499) );
  AND2_X1 U481bar ( .A1(in_78bar), .A2(in_6bar), .ZN(n499bar) );
  OR2_X1 U482 ( .A1(n497), .A2(n496), .ZN(n603) );
  AND2_X1 U482bar ( .A1(n497bar), .A2(n496bar), .ZN(n603bar) );
  OR2_X1 U483 ( .A1(in[112]), .A2(in[102]), .ZN(n496) );
  AND2_X1 U483bar ( .A1(inbar[112]), .A2(inbar[102]), .ZN(n496bar) );
  OR2_X1 U484 ( .A1(in[123]), .A2(n495), .ZN(n497) );
  AND2_X1 U484bar ( .A1(inbar[123]), .A2(n495bar), .ZN(n497bar) );
  OR2_X1 U485 ( .A1(in[143]), .A2(in[130]), .ZN(n495) );
  AND2_X1 U485bar ( .A1(inbar[143]), .A2(inbar[130]), .ZN(n495bar) );
  OR2_X1 U486 ( .A1(n494), .A2(n493), .ZN(n605) );
  AND2_X1 U486bar ( .A1(n494bar), .A2(n493bar), .ZN(n605bar) );
  OR2_X1 U487 ( .A1(n492), .A2(n491), .ZN(n493) );
  AND2_X1 U487bar ( .A1(n492bar), .A2(n491bar), .ZN(n493bar) );
  OR2_X1 U488 ( .A1(in[216]), .A2(in[213]), .ZN(n491) );
  AND2_X1 U488bar ( .A1(inbar[216]), .A2(inbar[213]), .ZN(n491bar) );
  OR2_X1 U489 ( .A1(in[227]), .A2(n490), .ZN(n492) );
  AND2_X1 U489bar ( .A1(inbar[227]), .A2(n490bar), .ZN(n492bar) );
  OR2_X1 U490 ( .A1(in_0), .A2(in[248]), .ZN(n490) );
  AND2_X1 U490bar ( .A1(in_0bar), .A2(inbar[248]), .ZN(n490bar) );
  OR2_X1 U491 ( .A1(n489), .A2(n488), .ZN(n494) );
  AND2_X1 U491bar ( .A1(n489bar), .A2(n488bar), .ZN(n494bar) );
  OR2_X1 U492 ( .A1(in_46), .A2(in_44), .ZN(n488) );
  AND2_X1 U492bar ( .A1(in_46bar), .A2(in_44bar), .ZN(n488bar) );
  OR2_X1 U493 ( .A1(in_50), .A2(n487), .ZN(n489) );
  AND2_X1 U493bar ( .A1(in_50bar), .A2(n487bar), .ZN(n489bar) );
  OR2_X1 U494 ( .A1(in_9), .A2(in_80), .ZN(n487) );
  AND2_X1 U494bar ( .A1(in_9bar), .A2(in_80bar), .ZN(n487bar) );
endmodule

module sBox_6 ( in, inbar, out, outbar );

  input wire [7:0] in;
  input wire [7:0] inbar;
//input_done

  output wire [7:0] out;
  output wire [7:0] outbar;
//output_done

  wire [255:0] decodeOut;
  wire [255:0] decodeOutbar;
//wire_done

  decode_6 dec ( .in(in), .inbar(inbar), .out(decodeOut), .outbar(decodeOutbar) );
  encode_6 enc ( .in(decodeOut), .inbar(decodeOutbar), .out(out), .outbar(outbar) );
endmodule

module CD2_25 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD2_26 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD2_27 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD2_28 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD4_13 ( a, abar, b, bbar, y, ybar );

  input wire [3:0] a;
  input wire [3:0] b;
  input wire [3:0] abar;
  input wire [3:0] bbar;
//input_done

  output wire [15:0] y;
  output wire [15:0] ybar;
//output_done

//wire_done

  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]) );
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]) );
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]) );
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]) );
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]) );
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]) );
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]) );
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]) );
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]) );
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]) );
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]) );
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]) );
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]) );
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]) );
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]) );
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]) );
endmodule

module CD4_14 ( a, abar, b, bbar, y, ybar );

  input wire [3:0] a;
  input wire [3:0] b;
  input wire [3:0] abar;
  input wire [3:0] bbar;
//input_done

  output wire [15:0] y;
  output wire [15:0] ybar;
//output_done

//wire_done

  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]) );
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]) );
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]) );
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]) );
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]) );
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]) );
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]) );
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]) );
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]) );
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]) );
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]) );
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]) );
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]) );
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]) );
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]) );
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]) );
endmodule

module CD16_7 ( a, abar, b, bbar, y, ybar );

  input wire [15:0] a;
  input wire [15:0] b;
  input wire [15:0] abar;
  input wire [15:0] bbar;
//input_done

  output wire [255:0] y;
  output wire [255:0] ybar;
//output_done

//wire_done

  AND2_X1 U1 ( .A1(b[9]), .A2(a[0]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[9]), .A2(abar[0]), .ZN(ybar[9]) );
  AND2_X1 U2 ( .A1(b[3]), .A2(a[6]), .ZN(y[99]) );
  OR2_X1 U2bar ( .A1(bbar[3]), .A2(abar[6]), .ZN(ybar[99]) );
  AND2_X1 U3 ( .A1(b[2]), .A2(a[6]), .ZN(y[98]) );
  OR2_X1 U3bar ( .A1(bbar[2]), .A2(abar[6]), .ZN(ybar[98]) );
  AND2_X1 U4 ( .A1(b[1]), .A2(a[6]), .ZN(y[97]) );
  OR2_X1 U4bar ( .A1(bbar[1]), .A2(abar[6]), .ZN(ybar[97]) );
  AND2_X1 U5 ( .A1(b[0]), .A2(a[6]), .ZN(y[96]) );
  OR2_X1 U5bar ( .A1(bbar[0]), .A2(abar[6]), .ZN(ybar[96]) );
  AND2_X1 U6 ( .A1(b[15]), .A2(a[5]), .ZN(y[95]) );
  OR2_X1 U6bar ( .A1(bbar[15]), .A2(abar[5]), .ZN(ybar[95]) );
  AND2_X1 U7 ( .A1(b[14]), .A2(a[5]), .ZN(y[94]) );
  OR2_X1 U7bar ( .A1(bbar[14]), .A2(abar[5]), .ZN(ybar[94]) );
  AND2_X1 U8 ( .A1(b[13]), .A2(a[5]), .ZN(y[93]) );
  OR2_X1 U8bar ( .A1(bbar[13]), .A2(abar[5]), .ZN(ybar[93]) );
  AND2_X1 U9 ( .A1(b[12]), .A2(a[5]), .ZN(y[92]) );
  OR2_X1 U9bar ( .A1(bbar[12]), .A2(abar[5]), .ZN(ybar[92]) );
  AND2_X1 U10 ( .A1(b[11]), .A2(a[5]), .ZN(y[91]) );
  OR2_X1 U10bar ( .A1(bbar[11]), .A2(abar[5]), .ZN(ybar[91]) );
  AND2_X1 U11 ( .A1(b[10]), .A2(a[5]), .ZN(y[90]) );
  OR2_X1 U11bar ( .A1(bbar[10]), .A2(abar[5]), .ZN(ybar[90]) );
  AND2_X1 U12 ( .A1(b[8]), .A2(a[0]), .ZN(y[8]) );
  OR2_X1 U12bar ( .A1(bbar[8]), .A2(abar[0]), .ZN(ybar[8]) );
  AND2_X1 U13 ( .A1(a[5]), .A2(b[9]), .ZN(y[89]) );
  OR2_X1 U13bar ( .A1(abar[5]), .A2(bbar[9]), .ZN(ybar[89]) );
  AND2_X1 U14 ( .A1(b[8]), .A2(a[5]), .ZN(y[88]) );
  OR2_X1 U14bar ( .A1(bbar[8]), .A2(abar[5]), .ZN(ybar[88]) );
  AND2_X1 U15 ( .A1(b[7]), .A2(a[5]), .ZN(y[87]) );
  OR2_X1 U15bar ( .A1(bbar[7]), .A2(abar[5]), .ZN(ybar[87]) );
  AND2_X1 U16 ( .A1(b[6]), .A2(a[5]), .ZN(y[86]) );
  OR2_X1 U16bar ( .A1(bbar[6]), .A2(abar[5]), .ZN(ybar[86]) );
  AND2_X1 U17 ( .A1(b[5]), .A2(a[5]), .ZN(y[85]) );
  OR2_X1 U17bar ( .A1(bbar[5]), .A2(abar[5]), .ZN(ybar[85]) );
  AND2_X1 U18 ( .A1(b[4]), .A2(a[5]), .ZN(y[84]) );
  OR2_X1 U18bar ( .A1(bbar[4]), .A2(abar[5]), .ZN(ybar[84]) );
  AND2_X1 U19 ( .A1(a[5]), .A2(b[3]), .ZN(y[83]) );
  OR2_X1 U19bar ( .A1(abar[5]), .A2(bbar[3]), .ZN(ybar[83]) );
  AND2_X1 U20 ( .A1(a[5]), .A2(b[2]), .ZN(y[82]) );
  OR2_X1 U20bar ( .A1(abar[5]), .A2(bbar[2]), .ZN(ybar[82]) );
  AND2_X1 U21 ( .A1(a[5]), .A2(b[1]), .ZN(y[81]) );
  OR2_X1 U21bar ( .A1(abar[5]), .A2(bbar[1]), .ZN(ybar[81]) );
  AND2_X1 U22 ( .A1(a[5]), .A2(b[0]), .ZN(y[80]) );
  OR2_X1 U22bar ( .A1(abar[5]), .A2(bbar[0]), .ZN(ybar[80]) );
  AND2_X1 U23 ( .A1(b[7]), .A2(a[0]), .ZN(y[7]) );
  OR2_X1 U23bar ( .A1(bbar[7]), .A2(abar[0]), .ZN(ybar[7]) );
  AND2_X1 U24 ( .A1(a[4]), .A2(b[15]), .ZN(y[79]) );
  OR2_X1 U24bar ( .A1(abar[4]), .A2(bbar[15]), .ZN(ybar[79]) );
  AND2_X1 U25 ( .A1(a[4]), .A2(b[14]), .ZN(y[78]) );
  OR2_X1 U25bar ( .A1(abar[4]), .A2(bbar[14]), .ZN(ybar[78]) );
  AND2_X1 U26 ( .A1(a[4]), .A2(b[13]), .ZN(y[77]) );
  OR2_X1 U26bar ( .A1(abar[4]), .A2(bbar[13]), .ZN(ybar[77]) );
  AND2_X1 U27 ( .A1(a[4]), .A2(b[12]), .ZN(y[76]) );
  OR2_X1 U27bar ( .A1(abar[4]), .A2(bbar[12]), .ZN(ybar[76]) );
  AND2_X1 U28 ( .A1(a[4]), .A2(b[11]), .ZN(y[75]) );
  OR2_X1 U28bar ( .A1(abar[4]), .A2(bbar[11]), .ZN(ybar[75]) );
  AND2_X1 U29 ( .A1(a[4]), .A2(b[10]), .ZN(y[74]) );
  OR2_X1 U29bar ( .A1(abar[4]), .A2(bbar[10]), .ZN(ybar[74]) );
  AND2_X1 U30 ( .A1(a[4]), .A2(b[9]), .ZN(y[73]) );
  OR2_X1 U30bar ( .A1(abar[4]), .A2(bbar[9]), .ZN(ybar[73]) );
  AND2_X1 U31 ( .A1(a[4]), .A2(b[8]), .ZN(y[72]) );
  OR2_X1 U31bar ( .A1(abar[4]), .A2(bbar[8]), .ZN(ybar[72]) );
  AND2_X1 U32 ( .A1(a[4]), .A2(b[7]), .ZN(y[71]) );
  OR2_X1 U32bar ( .A1(abar[4]), .A2(bbar[7]), .ZN(ybar[71]) );
  AND2_X1 U33 ( .A1(a[4]), .A2(b[6]), .ZN(y[70]) );
  OR2_X1 U33bar ( .A1(abar[4]), .A2(bbar[6]), .ZN(ybar[70]) );
  AND2_X1 U34 ( .A1(b[6]), .A2(a[0]), .ZN(y[6]) );
  OR2_X1 U34bar ( .A1(bbar[6]), .A2(abar[0]), .ZN(ybar[6]) );
  AND2_X1 U35 ( .A1(a[4]), .A2(b[5]), .ZN(y[69]) );
  OR2_X1 U35bar ( .A1(abar[4]), .A2(bbar[5]), .ZN(ybar[69]) );
  AND2_X1 U36 ( .A1(a[4]), .A2(b[4]), .ZN(y[68]) );
  OR2_X1 U36bar ( .A1(abar[4]), .A2(bbar[4]), .ZN(ybar[68]) );
  AND2_X1 U37 ( .A1(a[4]), .A2(b[3]), .ZN(y[67]) );
  OR2_X1 U37bar ( .A1(abar[4]), .A2(bbar[3]), .ZN(ybar[67]) );
  AND2_X1 U38 ( .A1(a[4]), .A2(b[2]), .ZN(y[66]) );
  OR2_X1 U38bar ( .A1(abar[4]), .A2(bbar[2]), .ZN(ybar[66]) );
  AND2_X1 U39 ( .A1(a[4]), .A2(b[1]), .ZN(y[65]) );
  OR2_X1 U39bar ( .A1(abar[4]), .A2(bbar[1]), .ZN(ybar[65]) );
  AND2_X1 U40 ( .A1(a[4]), .A2(b[0]), .ZN(y[64]) );
  OR2_X1 U40bar ( .A1(abar[4]), .A2(bbar[0]), .ZN(ybar[64]) );
  AND2_X1 U41 ( .A1(a[3]), .A2(b[15]), .ZN(y[63]) );
  OR2_X1 U41bar ( .A1(abar[3]), .A2(bbar[15]), .ZN(ybar[63]) );
  AND2_X1 U42 ( .A1(a[3]), .A2(b[14]), .ZN(y[62]) );
  OR2_X1 U42bar ( .A1(abar[3]), .A2(bbar[14]), .ZN(ybar[62]) );
  AND2_X1 U43 ( .A1(a[3]), .A2(b[13]), .ZN(y[61]) );
  OR2_X1 U43bar ( .A1(abar[3]), .A2(bbar[13]), .ZN(ybar[61]) );
  AND2_X1 U44 ( .A1(a[3]), .A2(b[12]), .ZN(y[60]) );
  OR2_X1 U44bar ( .A1(abar[3]), .A2(bbar[12]), .ZN(ybar[60]) );
  AND2_X1 U45 ( .A1(b[5]), .A2(a[0]), .ZN(y[5]) );
  OR2_X1 U45bar ( .A1(bbar[5]), .A2(abar[0]), .ZN(ybar[5]) );
  AND2_X1 U46 ( .A1(a[3]), .A2(b[11]), .ZN(y[59]) );
  OR2_X1 U46bar ( .A1(abar[3]), .A2(bbar[11]), .ZN(ybar[59]) );
  AND2_X1 U47 ( .A1(a[3]), .A2(b[10]), .ZN(y[58]) );
  OR2_X1 U47bar ( .A1(abar[3]), .A2(bbar[10]), .ZN(ybar[58]) );
  AND2_X1 U48 ( .A1(a[3]), .A2(b[9]), .ZN(y[57]) );
  OR2_X1 U48bar ( .A1(abar[3]), .A2(bbar[9]), .ZN(ybar[57]) );
  AND2_X1 U49 ( .A1(a[3]), .A2(b[8]), .ZN(y[56]) );
  OR2_X1 U49bar ( .A1(abar[3]), .A2(bbar[8]), .ZN(ybar[56]) );
  AND2_X1 U50 ( .A1(a[3]), .A2(b[7]), .ZN(y[55]) );
  OR2_X1 U50bar ( .A1(abar[3]), .A2(bbar[7]), .ZN(ybar[55]) );
  AND2_X1 U51 ( .A1(a[3]), .A2(b[6]), .ZN(y[54]) );
  OR2_X1 U51bar ( .A1(abar[3]), .A2(bbar[6]), .ZN(ybar[54]) );
  AND2_X1 U52 ( .A1(a[3]), .A2(b[5]), .ZN(y[53]) );
  OR2_X1 U52bar ( .A1(abar[3]), .A2(bbar[5]), .ZN(ybar[53]) );
  AND2_X1 U53 ( .A1(a[3]), .A2(b[4]), .ZN(y[52]) );
  OR2_X1 U53bar ( .A1(abar[3]), .A2(bbar[4]), .ZN(ybar[52]) );
  AND2_X1 U54 ( .A1(a[3]), .A2(b[3]), .ZN(y[51]) );
  OR2_X1 U54bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[51]) );
  AND2_X1 U55 ( .A1(a[3]), .A2(b[2]), .ZN(y[50]) );
  OR2_X1 U55bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[50]) );
  AND2_X1 U56 ( .A1(b[4]), .A2(a[0]), .ZN(y[4]) );
  OR2_X1 U56bar ( .A1(bbar[4]), .A2(abar[0]), .ZN(ybar[4]) );
  AND2_X1 U57 ( .A1(a[3]), .A2(b[1]), .ZN(y[49]) );
  OR2_X1 U57bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[49]) );
  AND2_X1 U58 ( .A1(a[3]), .A2(b[0]), .ZN(y[48]) );
  OR2_X1 U58bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[48]) );
  AND2_X1 U59 ( .A1(a[2]), .A2(b[15]), .ZN(y[47]) );
  OR2_X1 U59bar ( .A1(abar[2]), .A2(bbar[15]), .ZN(ybar[47]) );
  AND2_X1 U60 ( .A1(a[2]), .A2(b[14]), .ZN(y[46]) );
  OR2_X1 U60bar ( .A1(abar[2]), .A2(bbar[14]), .ZN(ybar[46]) );
  AND2_X1 U61 ( .A1(a[2]), .A2(b[13]), .ZN(y[45]) );
  OR2_X1 U61bar ( .A1(abar[2]), .A2(bbar[13]), .ZN(ybar[45]) );
  AND2_X1 U62 ( .A1(a[2]), .A2(b[12]), .ZN(y[44]) );
  OR2_X1 U62bar ( .A1(abar[2]), .A2(bbar[12]), .ZN(ybar[44]) );
  AND2_X1 U63 ( .A1(a[2]), .A2(b[11]), .ZN(y[43]) );
  OR2_X1 U63bar ( .A1(abar[2]), .A2(bbar[11]), .ZN(ybar[43]) );
  AND2_X1 U64 ( .A1(a[2]), .A2(b[10]), .ZN(y[42]) );
  OR2_X1 U64bar ( .A1(abar[2]), .A2(bbar[10]), .ZN(ybar[42]) );
  AND2_X1 U65 ( .A1(a[2]), .A2(b[9]), .ZN(y[41]) );
  OR2_X1 U65bar ( .A1(abar[2]), .A2(bbar[9]), .ZN(ybar[41]) );
  AND2_X1 U66 ( .A1(a[2]), .A2(b[8]), .ZN(y[40]) );
  OR2_X1 U66bar ( .A1(abar[2]), .A2(bbar[8]), .ZN(ybar[40]) );
  AND2_X1 U67 ( .A1(b[3]), .A2(a[0]), .ZN(y[3]) );
  OR2_X1 U67bar ( .A1(bbar[3]), .A2(abar[0]), .ZN(ybar[3]) );
  AND2_X1 U68 ( .A1(a[2]), .A2(b[7]), .ZN(y[39]) );
  OR2_X1 U68bar ( .A1(abar[2]), .A2(bbar[7]), .ZN(ybar[39]) );
  AND2_X1 U69 ( .A1(a[2]), .A2(b[6]), .ZN(y[38]) );
  OR2_X1 U69bar ( .A1(abar[2]), .A2(bbar[6]), .ZN(ybar[38]) );
  AND2_X1 U70 ( .A1(a[2]), .A2(b[5]), .ZN(y[37]) );
  OR2_X1 U70bar ( .A1(abar[2]), .A2(bbar[5]), .ZN(ybar[37]) );
  AND2_X1 U71 ( .A1(a[2]), .A2(b[4]), .ZN(y[36]) );
  OR2_X1 U71bar ( .A1(abar[2]), .A2(bbar[4]), .ZN(ybar[36]) );
  AND2_X1 U72 ( .A1(a[2]), .A2(b[3]), .ZN(y[35]) );
  OR2_X1 U72bar ( .A1(abar[2]), .A2(bbar[3]), .ZN(ybar[35]) );
  AND2_X1 U73 ( .A1(a[2]), .A2(b[2]), .ZN(y[34]) );
  OR2_X1 U73bar ( .A1(abar[2]), .A2(bbar[2]), .ZN(ybar[34]) );
  AND2_X1 U74 ( .A1(a[2]), .A2(b[1]), .ZN(y[33]) );
  OR2_X1 U74bar ( .A1(abar[2]), .A2(bbar[1]), .ZN(ybar[33]) );
  AND2_X1 U75 ( .A1(a[2]), .A2(b[0]), .ZN(y[32]) );
  OR2_X1 U75bar ( .A1(abar[2]), .A2(bbar[0]), .ZN(ybar[32]) );
  AND2_X1 U76 ( .A1(a[1]), .A2(b[15]), .ZN(y[31]) );
  OR2_X1 U76bar ( .A1(abar[1]), .A2(bbar[15]), .ZN(ybar[31]) );
  AND2_X1 U77 ( .A1(a[1]), .A2(b[14]), .ZN(y[30]) );
  OR2_X1 U77bar ( .A1(abar[1]), .A2(bbar[14]), .ZN(ybar[30]) );
  AND2_X1 U78 ( .A1(b[2]), .A2(a[0]), .ZN(y[2]) );
  OR2_X1 U78bar ( .A1(bbar[2]), .A2(abar[0]), .ZN(ybar[2]) );
  AND2_X1 U79 ( .A1(a[1]), .A2(b[13]), .ZN(y[29]) );
  OR2_X1 U79bar ( .A1(abar[1]), .A2(bbar[13]), .ZN(ybar[29]) );
  AND2_X1 U80 ( .A1(a[1]), .A2(b[12]), .ZN(y[28]) );
  OR2_X1 U80bar ( .A1(abar[1]), .A2(bbar[12]), .ZN(ybar[28]) );
  AND2_X1 U81 ( .A1(a[1]), .A2(b[11]), .ZN(y[27]) );
  OR2_X1 U81bar ( .A1(abar[1]), .A2(bbar[11]), .ZN(ybar[27]) );
  AND2_X1 U82 ( .A1(a[1]), .A2(b[10]), .ZN(y[26]) );
  OR2_X1 U82bar ( .A1(abar[1]), .A2(bbar[10]), .ZN(ybar[26]) );
  AND2_X1 U83 ( .A1(a[1]), .A2(b[9]), .ZN(y[25]) );
  OR2_X1 U83bar ( .A1(abar[1]), .A2(bbar[9]), .ZN(ybar[25]) );
  AND2_X1 U84 ( .A1(a[15]), .A2(b[15]), .ZN(y[255]) );
  OR2_X1 U84bar ( .A1(abar[15]), .A2(bbar[15]), .ZN(ybar[255]) );
  AND2_X1 U85 ( .A1(a[15]), .A2(b[14]), .ZN(y[254]) );
  OR2_X1 U85bar ( .A1(abar[15]), .A2(bbar[14]), .ZN(ybar[254]) );
  AND2_X1 U86 ( .A1(a[15]), .A2(b[13]), .ZN(y[253]) );
  OR2_X1 U86bar ( .A1(abar[15]), .A2(bbar[13]), .ZN(ybar[253]) );
  AND2_X1 U87 ( .A1(a[15]), .A2(b[12]), .ZN(y[252]) );
  OR2_X1 U87bar ( .A1(abar[15]), .A2(bbar[12]), .ZN(ybar[252]) );
  AND2_X1 U88 ( .A1(a[15]), .A2(b[11]), .ZN(y[251]) );
  OR2_X1 U88bar ( .A1(abar[15]), .A2(bbar[11]), .ZN(ybar[251]) );
  AND2_X1 U89 ( .A1(a[15]), .A2(b[10]), .ZN(y[250]) );
  OR2_X1 U89bar ( .A1(abar[15]), .A2(bbar[10]), .ZN(ybar[250]) );
  AND2_X1 U90 ( .A1(a[1]), .A2(b[8]), .ZN(y[24]) );
  OR2_X1 U90bar ( .A1(abar[1]), .A2(bbar[8]), .ZN(ybar[24]) );
  AND2_X1 U91 ( .A1(a[15]), .A2(b[9]), .ZN(y[249]) );
  OR2_X1 U91bar ( .A1(abar[15]), .A2(bbar[9]), .ZN(ybar[249]) );
  AND2_X1 U92 ( .A1(a[15]), .A2(b[8]), .ZN(y[248]) );
  OR2_X1 U92bar ( .A1(abar[15]), .A2(bbar[8]), .ZN(ybar[248]) );
  AND2_X1 U93 ( .A1(a[15]), .A2(b[7]), .ZN(y[247]) );
  OR2_X1 U93bar ( .A1(abar[15]), .A2(bbar[7]), .ZN(ybar[247]) );
  AND2_X1 U94 ( .A1(a[15]), .A2(b[6]), .ZN(y[246]) );
  OR2_X1 U94bar ( .A1(abar[15]), .A2(bbar[6]), .ZN(ybar[246]) );
  AND2_X1 U95 ( .A1(a[15]), .A2(b[5]), .ZN(y[245]) );
  OR2_X1 U95bar ( .A1(abar[15]), .A2(bbar[5]), .ZN(ybar[245]) );
  AND2_X1 U96 ( .A1(a[15]), .A2(b[4]), .ZN(y[244]) );
  OR2_X1 U96bar ( .A1(abar[15]), .A2(bbar[4]), .ZN(ybar[244]) );
  AND2_X1 U97 ( .A1(a[15]), .A2(b[3]), .ZN(y[243]) );
  OR2_X1 U97bar ( .A1(abar[15]), .A2(bbar[3]), .ZN(ybar[243]) );
  AND2_X1 U98 ( .A1(a[15]), .A2(b[2]), .ZN(y[242]) );
  OR2_X1 U98bar ( .A1(abar[15]), .A2(bbar[2]), .ZN(ybar[242]) );
  AND2_X1 U99 ( .A1(a[15]), .A2(b[1]), .ZN(y[241]) );
  OR2_X1 U99bar ( .A1(abar[15]), .A2(bbar[1]), .ZN(ybar[241]) );
  AND2_X1 U100 ( .A1(a[15]), .A2(b[0]), .ZN(y[240]) );
  OR2_X1 U100bar ( .A1(abar[15]), .A2(bbar[0]), .ZN(ybar[240]) );
  AND2_X1 U101 ( .A1(a[1]), .A2(b[7]), .ZN(y[23]) );
  OR2_X1 U101bar ( .A1(abar[1]), .A2(bbar[7]), .ZN(ybar[23]) );
  AND2_X1 U102 ( .A1(a[14]), .A2(b[15]), .ZN(y[239]) );
  OR2_X1 U102bar ( .A1(abar[14]), .A2(bbar[15]), .ZN(ybar[239]) );
  AND2_X1 U103 ( .A1(a[14]), .A2(b[14]), .ZN(y[238]) );
  OR2_X1 U103bar ( .A1(abar[14]), .A2(bbar[14]), .ZN(ybar[238]) );
  AND2_X1 U104 ( .A1(a[14]), .A2(b[13]), .ZN(y[237]) );
  OR2_X1 U104bar ( .A1(abar[14]), .A2(bbar[13]), .ZN(ybar[237]) );
  AND2_X1 U105 ( .A1(a[14]), .A2(b[12]), .ZN(y[236]) );
  OR2_X1 U105bar ( .A1(abar[14]), .A2(bbar[12]), .ZN(ybar[236]) );
  AND2_X1 U106 ( .A1(a[14]), .A2(b[11]), .ZN(y[235]) );
  OR2_X1 U106bar ( .A1(abar[14]), .A2(bbar[11]), .ZN(ybar[235]) );
  AND2_X1 U107 ( .A1(a[14]), .A2(b[10]), .ZN(y[234]) );
  OR2_X1 U107bar ( .A1(abar[14]), .A2(bbar[10]), .ZN(ybar[234]) );
  AND2_X1 U108 ( .A1(a[14]), .A2(b[9]), .ZN(y[233]) );
  OR2_X1 U108bar ( .A1(abar[14]), .A2(bbar[9]), .ZN(ybar[233]) );
  AND2_X1 U109 ( .A1(a[14]), .A2(b[8]), .ZN(y[232]) );
  OR2_X1 U109bar ( .A1(abar[14]), .A2(bbar[8]), .ZN(ybar[232]) );
  AND2_X1 U110 ( .A1(a[14]), .A2(b[7]), .ZN(y[231]) );
  OR2_X1 U110bar ( .A1(abar[14]), .A2(bbar[7]), .ZN(ybar[231]) );
  AND2_X1 U111 ( .A1(a[14]), .A2(b[6]), .ZN(y[230]) );
  OR2_X1 U111bar ( .A1(abar[14]), .A2(bbar[6]), .ZN(ybar[230]) );
  AND2_X1 U112 ( .A1(a[1]), .A2(b[6]), .ZN(y[22]) );
  OR2_X1 U112bar ( .A1(abar[1]), .A2(bbar[6]), .ZN(ybar[22]) );
  AND2_X1 U113 ( .A1(a[14]), .A2(b[5]), .ZN(y[229]) );
  OR2_X1 U113bar ( .A1(abar[14]), .A2(bbar[5]), .ZN(ybar[229]) );
  AND2_X1 U114 ( .A1(a[14]), .A2(b[4]), .ZN(y[228]) );
  OR2_X1 U114bar ( .A1(abar[14]), .A2(bbar[4]), .ZN(ybar[228]) );
  AND2_X1 U115 ( .A1(a[14]), .A2(b[3]), .ZN(y[227]) );
  OR2_X1 U115bar ( .A1(abar[14]), .A2(bbar[3]), .ZN(ybar[227]) );
  AND2_X1 U116 ( .A1(a[14]), .A2(b[2]), .ZN(y[226]) );
  OR2_X1 U116bar ( .A1(abar[14]), .A2(bbar[2]), .ZN(ybar[226]) );
  AND2_X1 U117 ( .A1(a[14]), .A2(b[1]), .ZN(y[225]) );
  OR2_X1 U117bar ( .A1(abar[14]), .A2(bbar[1]), .ZN(ybar[225]) );
  AND2_X1 U118 ( .A1(a[14]), .A2(b[0]), .ZN(y[224]) );
  OR2_X1 U118bar ( .A1(abar[14]), .A2(bbar[0]), .ZN(ybar[224]) );
  AND2_X1 U119 ( .A1(a[13]), .A2(b[15]), .ZN(y[223]) );
  OR2_X1 U119bar ( .A1(abar[13]), .A2(bbar[15]), .ZN(ybar[223]) );
  AND2_X1 U120 ( .A1(a[13]), .A2(b[14]), .ZN(y[222]) );
  OR2_X1 U120bar ( .A1(abar[13]), .A2(bbar[14]), .ZN(ybar[222]) );
  AND2_X1 U121 ( .A1(a[13]), .A2(b[13]), .ZN(y[221]) );
  OR2_X1 U121bar ( .A1(abar[13]), .A2(bbar[13]), .ZN(ybar[221]) );
  AND2_X1 U122 ( .A1(a[13]), .A2(b[12]), .ZN(y[220]) );
  OR2_X1 U122bar ( .A1(abar[13]), .A2(bbar[12]), .ZN(ybar[220]) );
  AND2_X1 U123 ( .A1(a[1]), .A2(b[5]), .ZN(y[21]) );
  OR2_X1 U123bar ( .A1(abar[1]), .A2(bbar[5]), .ZN(ybar[21]) );
  AND2_X1 U124 ( .A1(a[13]), .A2(b[11]), .ZN(y[219]) );
  OR2_X1 U124bar ( .A1(abar[13]), .A2(bbar[11]), .ZN(ybar[219]) );
  AND2_X1 U125 ( .A1(a[13]), .A2(b[10]), .ZN(y[218]) );
  OR2_X1 U125bar ( .A1(abar[13]), .A2(bbar[10]), .ZN(ybar[218]) );
  AND2_X1 U126 ( .A1(a[13]), .A2(b[9]), .ZN(y[217]) );
  OR2_X1 U126bar ( .A1(abar[13]), .A2(bbar[9]), .ZN(ybar[217]) );
  AND2_X1 U127 ( .A1(a[13]), .A2(b[8]), .ZN(y[216]) );
  OR2_X1 U127bar ( .A1(abar[13]), .A2(bbar[8]), .ZN(ybar[216]) );
  AND2_X1 U128 ( .A1(a[13]), .A2(b[7]), .ZN(y[215]) );
  OR2_X1 U128bar ( .A1(abar[13]), .A2(bbar[7]), .ZN(ybar[215]) );
  AND2_X1 U129 ( .A1(a[13]), .A2(b[6]), .ZN(y[214]) );
  OR2_X1 U129bar ( .A1(abar[13]), .A2(bbar[6]), .ZN(ybar[214]) );
  AND2_X1 U130 ( .A1(a[13]), .A2(b[5]), .ZN(y[213]) );
  OR2_X1 U130bar ( .A1(abar[13]), .A2(bbar[5]), .ZN(ybar[213]) );
  AND2_X1 U131 ( .A1(a[13]), .A2(b[4]), .ZN(y[212]) );
  OR2_X1 U131bar ( .A1(abar[13]), .A2(bbar[4]), .ZN(ybar[212]) );
  AND2_X1 U132 ( .A1(a[13]), .A2(b[3]), .ZN(y[211]) );
  OR2_X1 U132bar ( .A1(abar[13]), .A2(bbar[3]), .ZN(ybar[211]) );
  AND2_X1 U133 ( .A1(a[13]), .A2(b[2]), .ZN(y[210]) );
  OR2_X1 U133bar ( .A1(abar[13]), .A2(bbar[2]), .ZN(ybar[210]) );
  AND2_X1 U134 ( .A1(a[1]), .A2(b[4]), .ZN(y[20]) );
  OR2_X1 U134bar ( .A1(abar[1]), .A2(bbar[4]), .ZN(ybar[20]) );
  AND2_X1 U135 ( .A1(a[13]), .A2(b[1]), .ZN(y[209]) );
  OR2_X1 U135bar ( .A1(abar[13]), .A2(bbar[1]), .ZN(ybar[209]) );
  AND2_X1 U136 ( .A1(a[13]), .A2(b[0]), .ZN(y[208]) );
  OR2_X1 U136bar ( .A1(abar[13]), .A2(bbar[0]), .ZN(ybar[208]) );
  AND2_X1 U137 ( .A1(a[12]), .A2(b[15]), .ZN(y[207]) );
  OR2_X1 U137bar ( .A1(abar[12]), .A2(bbar[15]), .ZN(ybar[207]) );
  AND2_X1 U138 ( .A1(a[12]), .A2(b[14]), .ZN(y[206]) );
  OR2_X1 U138bar ( .A1(abar[12]), .A2(bbar[14]), .ZN(ybar[206]) );
  AND2_X1 U139 ( .A1(a[12]), .A2(b[13]), .ZN(y[205]) );
  OR2_X1 U139bar ( .A1(abar[12]), .A2(bbar[13]), .ZN(ybar[205]) );
  AND2_X1 U140 ( .A1(a[12]), .A2(b[12]), .ZN(y[204]) );
  OR2_X1 U140bar ( .A1(abar[12]), .A2(bbar[12]), .ZN(ybar[204]) );
  AND2_X1 U141 ( .A1(a[12]), .A2(b[11]), .ZN(y[203]) );
  OR2_X1 U141bar ( .A1(abar[12]), .A2(bbar[11]), .ZN(ybar[203]) );
  AND2_X1 U142 ( .A1(a[12]), .A2(b[10]), .ZN(y[202]) );
  OR2_X1 U142bar ( .A1(abar[12]), .A2(bbar[10]), .ZN(ybar[202]) );
  AND2_X1 U143 ( .A1(a[12]), .A2(b[9]), .ZN(y[201]) );
  OR2_X1 U143bar ( .A1(abar[12]), .A2(bbar[9]), .ZN(ybar[201]) );
  AND2_X1 U144 ( .A1(a[12]), .A2(b[8]), .ZN(y[200]) );
  OR2_X1 U144bar ( .A1(abar[12]), .A2(bbar[8]), .ZN(ybar[200]) );
  AND2_X1 U145 ( .A1(b[1]), .A2(a[0]), .ZN(y[1]) );
  OR2_X1 U145bar ( .A1(bbar[1]), .A2(abar[0]), .ZN(ybar[1]) );
  AND2_X1 U146 ( .A1(a[1]), .A2(b[3]), .ZN(y[19]) );
  OR2_X1 U146bar ( .A1(abar[1]), .A2(bbar[3]), .ZN(ybar[19]) );
  AND2_X1 U147 ( .A1(a[12]), .A2(b[7]), .ZN(y[199]) );
  OR2_X1 U147bar ( .A1(abar[12]), .A2(bbar[7]), .ZN(ybar[199]) );
  AND2_X1 U148 ( .A1(a[12]), .A2(b[6]), .ZN(y[198]) );
  OR2_X1 U148bar ( .A1(abar[12]), .A2(bbar[6]), .ZN(ybar[198]) );
  AND2_X1 U149 ( .A1(a[12]), .A2(b[5]), .ZN(y[197]) );
  OR2_X1 U149bar ( .A1(abar[12]), .A2(bbar[5]), .ZN(ybar[197]) );
  AND2_X1 U150 ( .A1(a[12]), .A2(b[4]), .ZN(y[196]) );
  OR2_X1 U150bar ( .A1(abar[12]), .A2(bbar[4]), .ZN(ybar[196]) );
  AND2_X1 U151 ( .A1(a[12]), .A2(b[3]), .ZN(y[195]) );
  OR2_X1 U151bar ( .A1(abar[12]), .A2(bbar[3]), .ZN(ybar[195]) );
  AND2_X1 U152 ( .A1(a[12]), .A2(b[2]), .ZN(y[194]) );
  OR2_X1 U152bar ( .A1(abar[12]), .A2(bbar[2]), .ZN(ybar[194]) );
  AND2_X1 U153 ( .A1(a[12]), .A2(b[1]), .ZN(y[193]) );
  OR2_X1 U153bar ( .A1(abar[12]), .A2(bbar[1]), .ZN(ybar[193]) );
  AND2_X1 U154 ( .A1(a[12]), .A2(b[0]), .ZN(y[192]) );
  OR2_X1 U154bar ( .A1(abar[12]), .A2(bbar[0]), .ZN(ybar[192]) );
  AND2_X1 U155 ( .A1(a[11]), .A2(b[15]), .ZN(y[191]) );
  OR2_X1 U155bar ( .A1(abar[11]), .A2(bbar[15]), .ZN(ybar[191]) );
  AND2_X1 U156 ( .A1(a[11]), .A2(b[14]), .ZN(y[190]) );
  OR2_X1 U156bar ( .A1(abar[11]), .A2(bbar[14]), .ZN(ybar[190]) );
  AND2_X1 U157 ( .A1(a[1]), .A2(b[2]), .ZN(y[18]) );
  OR2_X1 U157bar ( .A1(abar[1]), .A2(bbar[2]), .ZN(ybar[18]) );
  AND2_X1 U158 ( .A1(a[11]), .A2(b[13]), .ZN(y[189]) );
  OR2_X1 U158bar ( .A1(abar[11]), .A2(bbar[13]), .ZN(ybar[189]) );
  AND2_X1 U159 ( .A1(a[11]), .A2(b[12]), .ZN(y[188]) );
  OR2_X1 U159bar ( .A1(abar[11]), .A2(bbar[12]), .ZN(ybar[188]) );
  AND2_X1 U160 ( .A1(a[11]), .A2(b[11]), .ZN(y[187]) );
  OR2_X1 U160bar ( .A1(abar[11]), .A2(bbar[11]), .ZN(ybar[187]) );
  AND2_X1 U161 ( .A1(a[11]), .A2(b[10]), .ZN(y[186]) );
  OR2_X1 U161bar ( .A1(abar[11]), .A2(bbar[10]), .ZN(ybar[186]) );
  AND2_X1 U162 ( .A1(a[11]), .A2(b[9]), .ZN(y[185]) );
  OR2_X1 U162bar ( .A1(abar[11]), .A2(bbar[9]), .ZN(ybar[185]) );
  AND2_X1 U163 ( .A1(a[11]), .A2(b[8]), .ZN(y[184]) );
  OR2_X1 U163bar ( .A1(abar[11]), .A2(bbar[8]), .ZN(ybar[184]) );
  AND2_X1 U164 ( .A1(a[11]), .A2(b[7]), .ZN(y[183]) );
  OR2_X1 U164bar ( .A1(abar[11]), .A2(bbar[7]), .ZN(ybar[183]) );
  AND2_X1 U165 ( .A1(a[11]), .A2(b[6]), .ZN(y[182]) );
  OR2_X1 U165bar ( .A1(abar[11]), .A2(bbar[6]), .ZN(ybar[182]) );
  AND2_X1 U166 ( .A1(a[11]), .A2(b[5]), .ZN(y[181]) );
  OR2_X1 U166bar ( .A1(abar[11]), .A2(bbar[5]), .ZN(ybar[181]) );
  AND2_X1 U167 ( .A1(a[11]), .A2(b[4]), .ZN(y[180]) );
  OR2_X1 U167bar ( .A1(abar[11]), .A2(bbar[4]), .ZN(ybar[180]) );
  AND2_X1 U168 ( .A1(a[1]), .A2(b[1]), .ZN(y[17]) );
  OR2_X1 U168bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[17]) );
  AND2_X1 U169 ( .A1(a[11]), .A2(b[3]), .ZN(y[179]) );
  OR2_X1 U169bar ( .A1(abar[11]), .A2(bbar[3]), .ZN(ybar[179]) );
  AND2_X1 U170 ( .A1(a[11]), .A2(b[2]), .ZN(y[178]) );
  OR2_X1 U170bar ( .A1(abar[11]), .A2(bbar[2]), .ZN(ybar[178]) );
  AND2_X1 U171 ( .A1(a[11]), .A2(b[1]), .ZN(y[177]) );
  OR2_X1 U171bar ( .A1(abar[11]), .A2(bbar[1]), .ZN(ybar[177]) );
  AND2_X1 U172 ( .A1(a[11]), .A2(b[0]), .ZN(y[176]) );
  OR2_X1 U172bar ( .A1(abar[11]), .A2(bbar[0]), .ZN(ybar[176]) );
  AND2_X1 U173 ( .A1(a[10]), .A2(b[15]), .ZN(y[175]) );
  OR2_X1 U173bar ( .A1(abar[10]), .A2(bbar[15]), .ZN(ybar[175]) );
  AND2_X1 U174 ( .A1(a[10]), .A2(b[14]), .ZN(y[174]) );
  OR2_X1 U174bar ( .A1(abar[10]), .A2(bbar[14]), .ZN(ybar[174]) );
  AND2_X1 U175 ( .A1(a[10]), .A2(b[13]), .ZN(y[173]) );
  OR2_X1 U175bar ( .A1(abar[10]), .A2(bbar[13]), .ZN(ybar[173]) );
  AND2_X1 U176 ( .A1(a[10]), .A2(b[12]), .ZN(y[172]) );
  OR2_X1 U176bar ( .A1(abar[10]), .A2(bbar[12]), .ZN(ybar[172]) );
  AND2_X1 U177 ( .A1(a[10]), .A2(b[11]), .ZN(y[171]) );
  OR2_X1 U177bar ( .A1(abar[10]), .A2(bbar[11]), .ZN(ybar[171]) );
  AND2_X1 U178 ( .A1(a[10]), .A2(b[10]), .ZN(y[170]) );
  OR2_X1 U178bar ( .A1(abar[10]), .A2(bbar[10]), .ZN(ybar[170]) );
  AND2_X1 U179 ( .A1(a[1]), .A2(b[0]), .ZN(y[16]) );
  OR2_X1 U179bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[16]) );
  AND2_X1 U180 ( .A1(a[10]), .A2(b[9]), .ZN(y[169]) );
  OR2_X1 U180bar ( .A1(abar[10]), .A2(bbar[9]), .ZN(ybar[169]) );
  AND2_X1 U181 ( .A1(a[10]), .A2(b[8]), .ZN(y[168]) );
  OR2_X1 U181bar ( .A1(abar[10]), .A2(bbar[8]), .ZN(ybar[168]) );
  AND2_X1 U182 ( .A1(a[10]), .A2(b[7]), .ZN(y[167]) );
  OR2_X1 U182bar ( .A1(abar[10]), .A2(bbar[7]), .ZN(ybar[167]) );
  AND2_X1 U183 ( .A1(a[10]), .A2(b[6]), .ZN(y[166]) );
  OR2_X1 U183bar ( .A1(abar[10]), .A2(bbar[6]), .ZN(ybar[166]) );
  AND2_X1 U184 ( .A1(a[10]), .A2(b[5]), .ZN(y[165]) );
  OR2_X1 U184bar ( .A1(abar[10]), .A2(bbar[5]), .ZN(ybar[165]) );
  AND2_X1 U185 ( .A1(a[10]), .A2(b[4]), .ZN(y[164]) );
  OR2_X1 U185bar ( .A1(abar[10]), .A2(bbar[4]), .ZN(ybar[164]) );
  AND2_X1 U186 ( .A1(a[10]), .A2(b[3]), .ZN(y[163]) );
  OR2_X1 U186bar ( .A1(abar[10]), .A2(bbar[3]), .ZN(ybar[163]) );
  AND2_X1 U187 ( .A1(a[10]), .A2(b[2]), .ZN(y[162]) );
  OR2_X1 U187bar ( .A1(abar[10]), .A2(bbar[2]), .ZN(ybar[162]) );
  AND2_X1 U188 ( .A1(a[10]), .A2(b[1]), .ZN(y[161]) );
  OR2_X1 U188bar ( .A1(abar[10]), .A2(bbar[1]), .ZN(ybar[161]) );
  AND2_X1 U189 ( .A1(a[10]), .A2(b[0]), .ZN(y[160]) );
  OR2_X1 U189bar ( .A1(abar[10]), .A2(bbar[0]), .ZN(ybar[160]) );
  AND2_X1 U190 ( .A1(b[15]), .A2(a[0]), .ZN(y[15]) );
  OR2_X1 U190bar ( .A1(bbar[15]), .A2(abar[0]), .ZN(ybar[15]) );
  AND2_X1 U191 ( .A1(a[9]), .A2(b[15]), .ZN(y[159]) );
  OR2_X1 U191bar ( .A1(abar[9]), .A2(bbar[15]), .ZN(ybar[159]) );
  AND2_X1 U192 ( .A1(a[9]), .A2(b[14]), .ZN(y[158]) );
  OR2_X1 U192bar ( .A1(abar[9]), .A2(bbar[14]), .ZN(ybar[158]) );
  AND2_X1 U193 ( .A1(a[9]), .A2(b[13]), .ZN(y[157]) );
  OR2_X1 U193bar ( .A1(abar[9]), .A2(bbar[13]), .ZN(ybar[157]) );
  AND2_X1 U194 ( .A1(a[9]), .A2(b[12]), .ZN(y[156]) );
  OR2_X1 U194bar ( .A1(abar[9]), .A2(bbar[12]), .ZN(ybar[156]) );
  AND2_X1 U195 ( .A1(a[9]), .A2(b[11]), .ZN(y[155]) );
  OR2_X1 U195bar ( .A1(abar[9]), .A2(bbar[11]), .ZN(ybar[155]) );
  AND2_X1 U196 ( .A1(a[9]), .A2(b[10]), .ZN(y[154]) );
  OR2_X1 U196bar ( .A1(abar[9]), .A2(bbar[10]), .ZN(ybar[154]) );
  AND2_X1 U197 ( .A1(a[9]), .A2(b[9]), .ZN(y[153]) );
  OR2_X1 U197bar ( .A1(abar[9]), .A2(bbar[9]), .ZN(ybar[153]) );
  AND2_X1 U198 ( .A1(a[9]), .A2(b[8]), .ZN(y[152]) );
  OR2_X1 U198bar ( .A1(abar[9]), .A2(bbar[8]), .ZN(ybar[152]) );
  AND2_X1 U199 ( .A1(a[9]), .A2(b[7]), .ZN(y[151]) );
  OR2_X1 U199bar ( .A1(abar[9]), .A2(bbar[7]), .ZN(ybar[151]) );
  AND2_X1 U200 ( .A1(a[9]), .A2(b[6]), .ZN(y[150]) );
  OR2_X1 U200bar ( .A1(abar[9]), .A2(bbar[6]), .ZN(ybar[150]) );
  AND2_X1 U201 ( .A1(b[14]), .A2(a[0]), .ZN(y[14]) );
  OR2_X1 U201bar ( .A1(bbar[14]), .A2(abar[0]), .ZN(ybar[14]) );
  AND2_X1 U202 ( .A1(a[9]), .A2(b[5]), .ZN(y[149]) );
  OR2_X1 U202bar ( .A1(abar[9]), .A2(bbar[5]), .ZN(ybar[149]) );
  AND2_X1 U203 ( .A1(a[9]), .A2(b[4]), .ZN(y[148]) );
  OR2_X1 U203bar ( .A1(abar[9]), .A2(bbar[4]), .ZN(ybar[148]) );
  AND2_X1 U204 ( .A1(a[9]), .A2(b[3]), .ZN(y[147]) );
  OR2_X1 U204bar ( .A1(abar[9]), .A2(bbar[3]), .ZN(ybar[147]) );
  AND2_X1 U205 ( .A1(a[9]), .A2(b[2]), .ZN(y[146]) );
  OR2_X1 U205bar ( .A1(abar[9]), .A2(bbar[2]), .ZN(ybar[146]) );
  AND2_X1 U206 ( .A1(a[9]), .A2(b[1]), .ZN(y[145]) );
  OR2_X1 U206bar ( .A1(abar[9]), .A2(bbar[1]), .ZN(ybar[145]) );
  AND2_X1 U207 ( .A1(a[9]), .A2(b[0]), .ZN(y[144]) );
  OR2_X1 U207bar ( .A1(abar[9]), .A2(bbar[0]), .ZN(ybar[144]) );
  AND2_X1 U208 ( .A1(a[8]), .A2(b[15]), .ZN(y[143]) );
  OR2_X1 U208bar ( .A1(abar[8]), .A2(bbar[15]), .ZN(ybar[143]) );
  AND2_X1 U209 ( .A1(a[8]), .A2(b[14]), .ZN(y[142]) );
  OR2_X1 U209bar ( .A1(abar[8]), .A2(bbar[14]), .ZN(ybar[142]) );
  AND2_X1 U210 ( .A1(a[8]), .A2(b[13]), .ZN(y[141]) );
  OR2_X1 U210bar ( .A1(abar[8]), .A2(bbar[13]), .ZN(ybar[141]) );
  AND2_X1 U211 ( .A1(a[8]), .A2(b[12]), .ZN(y[140]) );
  OR2_X1 U211bar ( .A1(abar[8]), .A2(bbar[12]), .ZN(ybar[140]) );
  AND2_X1 U212 ( .A1(b[13]), .A2(a[0]), .ZN(y[13]) );
  OR2_X1 U212bar ( .A1(bbar[13]), .A2(abar[0]), .ZN(ybar[13]) );
  AND2_X1 U213 ( .A1(a[8]), .A2(b[11]), .ZN(y[139]) );
  OR2_X1 U213bar ( .A1(abar[8]), .A2(bbar[11]), .ZN(ybar[139]) );
  AND2_X1 U214 ( .A1(a[8]), .A2(b[10]), .ZN(y[138]) );
  OR2_X1 U214bar ( .A1(abar[8]), .A2(bbar[10]), .ZN(ybar[138]) );
  AND2_X1 U215 ( .A1(a[8]), .A2(b[9]), .ZN(y[137]) );
  OR2_X1 U215bar ( .A1(abar[8]), .A2(bbar[9]), .ZN(ybar[137]) );
  AND2_X1 U216 ( .A1(a[8]), .A2(b[8]), .ZN(y[136]) );
  OR2_X1 U216bar ( .A1(abar[8]), .A2(bbar[8]), .ZN(ybar[136]) );
  AND2_X1 U217 ( .A1(a[8]), .A2(b[7]), .ZN(y[135]) );
  OR2_X1 U217bar ( .A1(abar[8]), .A2(bbar[7]), .ZN(ybar[135]) );
  AND2_X1 U218 ( .A1(a[8]), .A2(b[6]), .ZN(y[134]) );
  OR2_X1 U218bar ( .A1(abar[8]), .A2(bbar[6]), .ZN(ybar[134]) );
  AND2_X1 U219 ( .A1(a[8]), .A2(b[5]), .ZN(y[133]) );
  OR2_X1 U219bar ( .A1(abar[8]), .A2(bbar[5]), .ZN(ybar[133]) );
  AND2_X1 U220 ( .A1(a[8]), .A2(b[4]), .ZN(y[132]) );
  OR2_X1 U220bar ( .A1(abar[8]), .A2(bbar[4]), .ZN(ybar[132]) );
  AND2_X1 U221 ( .A1(a[8]), .A2(b[3]), .ZN(y[131]) );
  OR2_X1 U221bar ( .A1(abar[8]), .A2(bbar[3]), .ZN(ybar[131]) );
  AND2_X1 U222 ( .A1(a[8]), .A2(b[2]), .ZN(y[130]) );
  OR2_X1 U222bar ( .A1(abar[8]), .A2(bbar[2]), .ZN(ybar[130]) );
  AND2_X1 U223 ( .A1(b[12]), .A2(a[0]), .ZN(y[12]) );
  OR2_X1 U223bar ( .A1(bbar[12]), .A2(abar[0]), .ZN(ybar[12]) );
  AND2_X1 U224 ( .A1(a[8]), .A2(b[1]), .ZN(y[129]) );
  OR2_X1 U224bar ( .A1(abar[8]), .A2(bbar[1]), .ZN(ybar[129]) );
  AND2_X1 U225 ( .A1(a[8]), .A2(b[0]), .ZN(y[128]) );
  OR2_X1 U225bar ( .A1(abar[8]), .A2(bbar[0]), .ZN(ybar[128]) );
  AND2_X1 U226 ( .A1(a[7]), .A2(b[15]), .ZN(y[127]) );
  OR2_X1 U226bar ( .A1(abar[7]), .A2(bbar[15]), .ZN(ybar[127]) );
  AND2_X1 U227 ( .A1(a[7]), .A2(b[14]), .ZN(y[126]) );
  OR2_X1 U227bar ( .A1(abar[7]), .A2(bbar[14]), .ZN(ybar[126]) );
  AND2_X1 U228 ( .A1(a[7]), .A2(b[13]), .ZN(y[125]) );
  OR2_X1 U228bar ( .A1(abar[7]), .A2(bbar[13]), .ZN(ybar[125]) );
  AND2_X1 U229 ( .A1(a[7]), .A2(b[12]), .ZN(y[124]) );
  OR2_X1 U229bar ( .A1(abar[7]), .A2(bbar[12]), .ZN(ybar[124]) );
  AND2_X1 U230 ( .A1(a[7]), .A2(b[11]), .ZN(y[123]) );
  OR2_X1 U230bar ( .A1(abar[7]), .A2(bbar[11]), .ZN(ybar[123]) );
  AND2_X1 U231 ( .A1(a[7]), .A2(b[10]), .ZN(y[122]) );
  OR2_X1 U231bar ( .A1(abar[7]), .A2(bbar[10]), .ZN(ybar[122]) );
  AND2_X1 U232 ( .A1(a[7]), .A2(b[9]), .ZN(y[121]) );
  OR2_X1 U232bar ( .A1(abar[7]), .A2(bbar[9]), .ZN(ybar[121]) );
  AND2_X1 U233 ( .A1(a[7]), .A2(b[8]), .ZN(y[120]) );
  OR2_X1 U233bar ( .A1(abar[7]), .A2(bbar[8]), .ZN(ybar[120]) );
  AND2_X1 U234 ( .A1(b[11]), .A2(a[0]), .ZN(y[11]) );
  OR2_X1 U234bar ( .A1(bbar[11]), .A2(abar[0]), .ZN(ybar[11]) );
  AND2_X1 U235 ( .A1(a[7]), .A2(b[7]), .ZN(y[119]) );
  OR2_X1 U235bar ( .A1(abar[7]), .A2(bbar[7]), .ZN(ybar[119]) );
  AND2_X1 U236 ( .A1(a[7]), .A2(b[6]), .ZN(y[118]) );
  OR2_X1 U236bar ( .A1(abar[7]), .A2(bbar[6]), .ZN(ybar[118]) );
  AND2_X1 U237 ( .A1(a[7]), .A2(b[5]), .ZN(y[117]) );
  OR2_X1 U237bar ( .A1(abar[7]), .A2(bbar[5]), .ZN(ybar[117]) );
  AND2_X1 U238 ( .A1(a[7]), .A2(b[4]), .ZN(y[116]) );
  OR2_X1 U238bar ( .A1(abar[7]), .A2(bbar[4]), .ZN(ybar[116]) );
  AND2_X1 U239 ( .A1(a[7]), .A2(b[3]), .ZN(y[115]) );
  OR2_X1 U239bar ( .A1(abar[7]), .A2(bbar[3]), .ZN(ybar[115]) );
  AND2_X1 U240 ( .A1(a[7]), .A2(b[2]), .ZN(y[114]) );
  OR2_X1 U240bar ( .A1(abar[7]), .A2(bbar[2]), .ZN(ybar[114]) );
  AND2_X1 U241 ( .A1(a[7]), .A2(b[1]), .ZN(y[113]) );
  OR2_X1 U241bar ( .A1(abar[7]), .A2(bbar[1]), .ZN(ybar[113]) );
  AND2_X1 U242 ( .A1(a[7]), .A2(b[0]), .ZN(y[112]) );
  OR2_X1 U242bar ( .A1(abar[7]), .A2(bbar[0]), .ZN(ybar[112]) );
  AND2_X1 U243 ( .A1(b[15]), .A2(a[6]), .ZN(y[111]) );
  OR2_X1 U243bar ( .A1(bbar[15]), .A2(abar[6]), .ZN(ybar[111]) );
  AND2_X1 U244 ( .A1(b[14]), .A2(a[6]), .ZN(y[110]) );
  OR2_X1 U244bar ( .A1(bbar[14]), .A2(abar[6]), .ZN(ybar[110]) );
  AND2_X1 U245 ( .A1(b[10]), .A2(a[0]), .ZN(y[10]) );
  OR2_X1 U245bar ( .A1(bbar[10]), .A2(abar[0]), .ZN(ybar[10]) );
  AND2_X1 U246 ( .A1(b[13]), .A2(a[6]), .ZN(y[109]) );
  OR2_X1 U246bar ( .A1(bbar[13]), .A2(abar[6]), .ZN(ybar[109]) );
  AND2_X1 U247 ( .A1(b[12]), .A2(a[6]), .ZN(y[108]) );
  OR2_X1 U247bar ( .A1(bbar[12]), .A2(abar[6]), .ZN(ybar[108]) );
  AND2_X1 U248 ( .A1(b[11]), .A2(a[6]), .ZN(y[107]) );
  OR2_X1 U248bar ( .A1(bbar[11]), .A2(abar[6]), .ZN(ybar[107]) );
  AND2_X1 U249 ( .A1(b[10]), .A2(a[6]), .ZN(y[106]) );
  OR2_X1 U249bar ( .A1(bbar[10]), .A2(abar[6]), .ZN(ybar[106]) );
  AND2_X1 U250 ( .A1(a[6]), .A2(b[9]), .ZN(y[105]) );
  OR2_X1 U250bar ( .A1(abar[6]), .A2(bbar[9]), .ZN(ybar[105]) );
  AND2_X1 U251 ( .A1(b[8]), .A2(a[6]), .ZN(y[104]) );
  OR2_X1 U251bar ( .A1(bbar[8]), .A2(abar[6]), .ZN(ybar[104]) );
  AND2_X1 U252 ( .A1(b[7]), .A2(a[6]), .ZN(y[103]) );
  OR2_X1 U252bar ( .A1(bbar[7]), .A2(abar[6]), .ZN(ybar[103]) );
  AND2_X1 U253 ( .A1(b[6]), .A2(a[6]), .ZN(y[102]) );
  OR2_X1 U253bar ( .A1(bbar[6]), .A2(abar[6]), .ZN(ybar[102]) );
  AND2_X1 U254 ( .A1(b[5]), .A2(a[6]), .ZN(y[101]) );
  OR2_X1 U254bar ( .A1(bbar[5]), .A2(abar[6]), .ZN(ybar[101]) );
  AND2_X1 U255 ( .A1(b[4]), .A2(a[6]), .ZN(y[100]) );
  OR2_X1 U255bar ( .A1(bbar[4]), .A2(abar[6]), .ZN(ybar[100]) );
  AND2_X1 U256 ( .A1(b[0]), .A2(a[0]), .ZN(y[0]) );
  OR2_X1 U256bar ( .A1(bbar[0]), .A2(abar[0]), .ZN(ybar[0]) );
endmodule

module decode_7 ( in, inbar, out, outbar );

  input wire [7:0] in;
  input wire [7:0] inbar;
//input_done

  output wire [255:0] out;
  output wire [255:0] outbar;
//output_done

  wire [15:0] level1;
  wire [31:0] level2;
  wire [15:0] level1bar;
  wire [31:0] level2bar;
//wire_done

  CD2_28 cd_l1_1 ( .a(in[1]), .abar(inbar[1]), .b(in[0]), .bbar(inbar[0]), .y(level1[3:0]), .ybar(level1bar[3:0]) );
  CD2_27 cd_l1_2 ( .a(in[3]), .abar(inbar[3]), .b(in[2]), .bbar(inbar[2]), .y(level1[7:4]), .ybar(level1bar[7:4]) );
  CD2_26 cd_l1_3 ( .a(in[5]), .abar(inbar[5]), .b(in[4]), .bbar(inbar[4]), .y(level1[11:8]), .ybar(level1bar[11:8]) );
  CD2_25 cd_l1_4 ( .a(in[7]), .abar(inbar[7]), .b(in[6]), .bbar(inbar[6]), .y(level1[15:12]), .ybar(level1bar[15:12]) );

  CD4_14 cd_l2_1 ( .a(level1[7:4]), .abar(level1bar[7:4]), .b(level1[3:0]), .bbar(level1bar[3:0]), 
        .y(level2[15:0]), .ybar(level2bar[15:0]) );
  CD4_13 cd_l2_2 ( .a(level1[15:12]), .abar(level1bar[15:12]), .b(level1[11:8]), .bbar(level1bar[11:8]), 
        .y(level2[31:16]), .ybar(level2bar[31:16]) );
  CD16_7 cd_l3 ( .a(level2[31:16]), .abar(level2bar[31:16]), .b(level2[15:0]), .bbar(level2bar[15:0]), 
        .y(out), .ybar(outbar) );
endmodule

module encode_7 ( in, inbar, out, outbar );

  input wire [255:0] in;
  input wire [255:0] inbar;
//input_done

  output wire [7:0] out;
  output wire [7:0] outbar;
//output_done

  wire in_81;
  wire in_80;
  wire in_79;
  wire in_78;
  wire in_77;
  wire in_76;
  wire in_75;
  wire in_74;
  wire in_73;
  wire in_72;
  wire in_71;
  wire in_70;
  wire in_69;
  wire in_68;
  wire in_67;
  wire in_66;
  wire in_65;
  wire in_64;
  wire in_63;
  wire in_62;
  wire in_61;
  wire in_60;
  wire in_59;
  wire in_58;
  wire in_57;
  wire in_56;
  wire in_55;
  wire in_54;
  wire in_53;
  wire in_52;
  wire in_51;
  wire in_50;
  wire in_49;
  wire in_48;
  wire in_47;
  wire in_46;
  wire in_45;
  wire in_44;
  wire in_43;
  wire in_42;
  wire in_41;
  wire in_40;
  wire in_39;
  wire in_38;
  wire in_37;
  wire in_36;
  wire in_35;
  wire in_34;
  wire in_33;
  wire in_32;
  wire in_31;
  wire in_30;
  wire in_29;
  wire in_28;
  wire in_27;
  wire in_26;
  wire in_25;
  wire in_24;
  wire in_23;
  wire in_22;
  wire in_21;
  wire in_20;
  wire in_19;
  wire in_18;
  wire in_17;
  wire in_16;
  wire in_15;
  wire in_14;
  wire in_13;
  wire in_12;
  wire in_11;
  wire in_10;
  wire in_9;
  wire in_8;
  wire in_7;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_3;
  wire in_2;
  wire in_1;
  wire in_0;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire in_81bar;
  wire in_80bar;
  wire in_79bar;
  wire in_78bar;
  wire in_77bar;
  wire in_76bar;
  wire in_75bar;
  wire in_74bar;
  wire in_73bar;
  wire in_72bar;
  wire in_71bar;
  wire in_70bar;
  wire in_69bar;
  wire in_68bar;
  wire in_67bar;
  wire in_66bar;
  wire in_65bar;
  wire in_64bar;
  wire in_63bar;
  wire in_62bar;
  wire in_61bar;
  wire in_60bar;
  wire in_59bar;
  wire in_58bar;
  wire in_57bar;
  wire in_56bar;
  wire in_55bar;
  wire in_54bar;
  wire in_53bar;
  wire in_52bar;
  wire in_51bar;
  wire in_50bar;
  wire in_49bar;
  wire in_48bar;
  wire in_47bar;
  wire in_46bar;
  wire in_45bar;
  wire in_44bar;
  wire in_43bar;
  wire in_42bar;
  wire in_41bar;
  wire in_40bar;
  wire in_39bar;
  wire in_38bar;
  wire in_37bar;
  wire in_36bar;
  wire in_35bar;
  wire in_34bar;
  wire in_33bar;
  wire in_32bar;
  wire in_31bar;
  wire in_30bar;
  wire in_29bar;
  wire in_28bar;
  wire in_27bar;
  wire in_26bar;
  wire in_25bar;
  wire in_24bar;
  wire in_23bar;
  wire in_22bar;
  wire in_21bar;
  wire in_20bar;
  wire in_19bar;
  wire in_18bar;
  wire in_17bar;
  wire in_16bar;
  wire in_15bar;
  wire in_14bar;
  wire in_13bar;
  wire in_12bar;
  wire in_11bar;
  wire in_10bar;
  wire in_9bar;
  wire in_8bar;
  wire in_7bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_3bar;
  wire in_2bar;
  wire in_1bar;
  wire in_0bar;
  wire n487bar;
  wire n488bar;
  wire n489bar;
  wire n490bar;
  wire n491bar;
  wire n492bar;
  wire n493bar;
  wire n494bar;
  wire n495bar;
  wire n496bar;
  wire n497bar;
  wire n498bar;
  wire n499bar;
  wire n500bar;
  wire n501bar;
  wire n502bar;
  wire n503bar;
  wire n504bar;
  wire n505bar;
  wire n506bar;
  wire n507bar;
  wire n508bar;
  wire n509bar;
  wire n510bar;
  wire n511bar;
  wire n512bar;
  wire n513bar;
  wire n514bar;
  wire n515bar;
  wire n516bar;
  wire n517bar;
  wire n518bar;
  wire n519bar;
  wire n520bar;
  wire n521bar;
  wire n522bar;
  wire n523bar;
  wire n524bar;
  wire n525bar;
  wire n526bar;
  wire n527bar;
  wire n528bar;
  wire n529bar;
  wire n530bar;
  wire n531bar;
  wire n532bar;
  wire n533bar;
  wire n534bar;
  wire n535bar;
  wire n536bar;
  wire n537bar;
  wire n538bar;
  wire n539bar;
  wire n540bar;
  wire n541bar;
  wire n542bar;
  wire n543bar;
  wire n544bar;
  wire n545bar;
  wire n546bar;
  wire n547bar;
  wire n548bar;
  wire n549bar;
  wire n550bar;
  wire n551bar;
  wire n552bar;
  wire n553bar;
  wire n554bar;
  wire n555bar;
  wire n556bar;
  wire n557bar;
  wire n558bar;
  wire n559bar;
  wire n560bar;
  wire n561bar;
  wire n562bar;
  wire n563bar;
  wire n564bar;
  wire n565bar;
  wire n566bar;
  wire n567bar;
  wire n568bar;
  wire n569bar;
  wire n570bar;
  wire n571bar;
  wire n572bar;
  wire n573bar;
  wire n574bar;
  wire n575bar;
  wire n576bar;
  wire n577bar;
  wire n578bar;
  wire n579bar;
  wire n580bar;
  wire n581bar;
  wire n582bar;
  wire n583bar;
  wire n584bar;
  wire n585bar;
  wire n586bar;
  wire n587bar;
  wire n588bar;
  wire n589bar;
  wire n590bar;
  wire n591bar;
  wire n592bar;
  wire n593bar;
  wire n594bar;
  wire n595bar;
  wire n596bar;
  wire n597bar;
  wire n598bar;
  wire n599bar;
  wire n600bar;
  wire n601bar;
  wire n602bar;
  wire n603bar;
  wire n604bar;
  wire n605bar;
  wire n606bar;
  wire n607bar;
  wire n608bar;
  wire n609bar;
  wire n610bar;
  wire n611bar;
  wire n612bar;
  wire n613bar;
  wire n614bar;
  wire n615bar;
  wire n616bar;
  wire n617bar;
  wire n618bar;
  wire n619bar;
  wire n620bar;
  wire n621bar;
  wire n622bar;
  wire n623bar;
  wire n624bar;
  wire n625bar;
  wire n626bar;
  wire n627bar;
  wire n628bar;
  wire n629bar;
  wire n630bar;
  wire n631bar;
  wire n632bar;
  wire n633bar;
  wire n634bar;
  wire n635bar;
  wire n636bar;
  wire n637bar;
  wire n638bar;
  wire n639bar;
  wire n640bar;
  wire n641bar;
  wire n642bar;
  wire n643bar;
  wire n644bar;
  wire n645bar;
  wire n646bar;
  wire n647bar;
  wire n648bar;
  wire n649bar;
  wire n650bar;
  wire n651bar;
  wire n652bar;
  wire n653bar;
  wire n654bar;
  wire n655bar;
  wire n656bar;
  wire n657bar;
  wire n658bar;
  wire n659bar;
  wire n660bar;
  wire n661bar;
  wire n662bar;
  wire n663bar;
  wire n664bar;
  wire n665bar;
  wire n666bar;
  wire n667bar;
  wire n668bar;
  wire n669bar;
  wire n670bar;
  wire n671bar;
  wire n672bar;
  wire n673bar;
  wire n674bar;
  wire n675bar;
  wire n676bar;
  wire n677bar;
  wire n678bar;
  wire n679bar;
  wire n680bar;
  wire n681bar;
  wire n682bar;
  wire n683bar;
  wire n684bar;
  wire n685bar;
  wire n686bar;
  wire n687bar;
  wire n688bar;
  wire n689bar;
  wire n690bar;
  wire n691bar;
  wire n692bar;
  wire n693bar;
  wire n694bar;
  wire n695bar;
  wire n696bar;
  wire n697bar;
  wire n698bar;
  wire n699bar;
  wire n700bar;
  wire n701bar;
  wire n702bar;
  wire n703bar;
  wire n704bar;
  wire n705bar;
  wire n706bar;
  wire n707bar;
  wire n708bar;
  wire n709bar;
  wire n710bar;
  wire n711bar;
  wire n712bar;
  wire n713bar;
  wire n714bar;
  wire n715bar;
  wire n716bar;
  wire n717bar;
  wire n718bar;
  wire n719bar;
  wire n720bar;
  wire n721bar;
  wire n722bar;
  wire n723bar;
  wire n724bar;
  wire n725bar;
  wire n726bar;
  wire n727bar;
  wire n728bar;
  wire n729bar;
  wire n730bar;
  wire n731bar;
  wire n732bar;
  wire n733bar;
  wire n734bar;
  wire n735bar;
  wire n736bar;
  wire n737bar;
  wire n738bar;
  wire n739bar;
  wire n740bar;
  wire n741bar;
  wire n742bar;
  wire n743bar;
  wire n744bar;
  wire n745bar;
  wire n746bar;
  wire n747bar;
  wire n748bar;
  wire n749bar;
  wire n750bar;
  wire n751bar;
  wire n752bar;
  wire n753bar;
  wire n754bar;
  wire n755bar;
  wire n756bar;
  wire n757bar;
  wire n758bar;
  wire n759bar;
  wire n760bar;
  wire n761bar;
  wire n762bar;
  wire n763bar;
  wire n764bar;
  wire n765bar;
  wire n766bar;
  wire n767bar;
  wire n768bar;
  wire n769bar;
  wire n770bar;
  wire n771bar;
  wire n772bar;
  wire n773bar;
  wire n774bar;
  wire n775bar;
  wire n776bar;
  wire n777bar;
  wire n778bar;
  wire n779bar;
  wire n780bar;
  wire n781bar;
  wire n782bar;
  wire n783bar;
  wire n784bar;
  wire n785bar;
  wire n786bar;
  wire n787bar;
  wire n788bar;
  wire n789bar;
  wire n790bar;
  wire n791bar;
  wire n792bar;
  wire n793bar;
  wire n794bar;
  wire n795bar;
  wire n796bar;
  wire n797bar;
  wire n798bar;
  wire n799bar;
  wire n800bar;
  wire n801bar;
  wire n802bar;
  wire n803bar;
  wire n804bar;
  wire n805bar;
  wire n806bar;
  wire n807bar;
  wire n808bar;
  wire n809bar;
  wire n810bar;
  wire n811bar;
  wire n812bar;
  wire n813bar;
  wire n814bar;
  wire n815bar;
  wire n816bar;
  wire n817bar;
  wire n818bar;
  wire n819bar;
  wire n820bar;
  wire n821bar;
  wire n822bar;
  wire n823bar;
  wire n824bar;
  wire n825bar;
  wire n826bar;
  wire n827bar;
  wire n828bar;
  wire n829bar;
  wire n830bar;
  wire n831bar;
  wire n832bar;
  wire n833bar;
  wire n834bar;
  wire n835bar;
  wire n836bar;
  wire n837bar;
  wire n838bar;
  wire n839bar;
  wire n840bar;
  wire n841bar;
  wire n842bar;
  wire n843bar;
  wire n844bar;
  wire n845bar;
  wire n846bar;
  wire n847bar;
  wire n848bar;
  wire n849bar;
  wire n850bar;
  wire n851bar;
  wire n852bar;
  wire n853bar;
  wire n854bar;
  wire n855bar;
  wire n856bar;
  wire n857bar;
  wire n858bar;
  wire n859bar;
  wire n860bar;
  wire n861bar;
  wire n862bar;
  wire n863bar;
  wire n864bar;
  wire n865bar;
  wire n866bar;
  wire n867bar;
  wire n868bar;
  wire n869bar;
  wire n870bar;
  wire n871bar;
  wire n872bar;
  wire n873bar;
  wire n874bar;
  wire n875bar;
  wire n876bar;
  wire n877bar;
  wire n878bar;
  wire n879bar;
  wire n880bar;
  wire n881bar;
  wire n882bar;
  wire n883bar;
  wire n884bar;
  wire n885bar;
  wire n886bar;
  wire n887bar;
  wire n888bar;
  wire n889bar;
  wire n890bar;
  wire n891bar;
  wire n892bar;
  wire n893bar;
  wire n894bar;
  wire n895bar;
  wire n896bar;
  wire n897bar;
  wire n898bar;
  wire n899bar;
  wire n900bar;
  wire n901bar;
  wire n902bar;
  wire n903bar;
  wire n904bar;
  wire n905bar;
  wire n906bar;
  wire n907bar;
  wire n908bar;
  wire n909bar;
  wire n910bar;
  wire n911bar;
  wire n912bar;
  wire n913bar;
  wire n914bar;
  wire n915bar;
  wire n916bar;
  wire n917bar;
  wire n918bar;
  wire n919bar;
  wire n920bar;
  wire n921bar;
  wire n922bar;
  wire n923bar;
  wire n924bar;
  wire n925bar;
  wire n926bar;
  wire n927bar;
  wire n928bar;
  wire n929bar;
  wire n930bar;
  wire n931bar;
  wire n932bar;
  wire n933bar;
  wire n934bar;
  wire n935bar;
  wire n936bar;
  wire n937bar;
  wire n938bar;
  wire n939bar;
  wire n940bar;
  wire n941bar;
  wire n942bar;
  wire n943bar;
  wire n944bar;
  wire n945bar;
  wire n946bar;
  wire n947bar;
  wire n948bar;
  wire n949bar;
  wire n950bar;
  wire n951bar;
  wire n952bar;
  wire n953bar;
  wire n954bar;
  wire n955bar;
  wire n956bar;
  wire n957bar;
  wire n958bar;
  wire n959bar;
  wire n960bar;
  wire n961bar;
  wire n962bar;
  wire n963bar;
  wire n964bar;
  wire n965bar;
  wire n966bar;
  wire n967bar;
  wire n968bar;
  wire n969bar;
  wire n970bar;
  wire n971bar;
  wire n972bar;
//wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];
  assign in_81bar = inbar[81];
  assign in_80bar = inbar[80];
  assign in_79bar = inbar[79];
  assign in_78bar = inbar[78];
  assign in_77bar = inbar[77];
  assign in_76bar = inbar[76];
  assign in_75bar = inbar[75];
  assign in_74bar = inbar[74];
  assign in_73bar = inbar[73];
  assign in_72bar = inbar[72];
  assign in_71bar = inbar[71];
  assign in_70bar = inbar[70];
  assign in_69bar = inbar[69];
  assign in_68bar = inbar[68];
  assign in_67bar = inbar[67];
  assign in_66bar = inbar[66];
  assign in_65bar = inbar[65];
  assign in_64bar = inbar[64];
  assign in_63bar = inbar[63];
  assign in_62bar = inbar[62];
  assign in_61bar = inbar[61];
  assign in_60bar = inbar[60];
  assign in_59bar = inbar[59];
  assign in_58bar = inbar[58];
  assign in_57bar = inbar[57];
  assign in_56bar = inbar[56];
  assign in_55bar = inbar[55];
  assign in_54bar = inbar[54];
  assign in_53bar = inbar[53];
  assign in_52bar = inbar[52];
  assign in_51bar = inbar[51];
  assign in_50bar = inbar[50];
  assign in_49bar = inbar[49];
  assign in_48bar = inbar[48];
  assign in_47bar = inbar[47];
  assign in_46bar = inbar[46];
  assign in_45bar = inbar[45];
  assign in_44bar = inbar[44];
  assign in_43bar = inbar[43];
  assign in_42bar = inbar[42];
  assign in_41bar = inbar[41];
  assign in_40bar = inbar[40];
  assign in_39bar = inbar[39];
  assign in_38bar = inbar[38];
  assign in_37bar = inbar[37];
  assign in_36bar = inbar[36];
  assign in_35bar = inbar[35];
  assign in_34bar = inbar[34];
  assign in_33bar = inbar[33];
  assign in_32bar = inbar[32];
  assign in_31bar = inbar[31];
  assign in_30bar = inbar[30];
  assign in_29bar = inbar[29];
  assign in_28bar = inbar[28];
  assign in_27bar = inbar[27];
  assign in_26bar = inbar[26];
  assign in_25bar = inbar[25];
  assign in_24bar = inbar[24];
  assign in_23bar = inbar[23];
  assign in_22bar = inbar[22];
  assign in_21bar = inbar[21];
  assign in_20bar = inbar[20];
  assign in_19bar = inbar[19];
  assign in_18bar = inbar[18];
  assign in_17bar = inbar[17];
  assign in_16bar = inbar[16];
  assign in_15bar = inbar[15];
  assign in_14bar = inbar[14];
  assign in_13bar = inbar[13];
  assign in_12bar = inbar[12];
  assign in_11bar = inbar[11];
  assign in_10bar = inbar[10];
  assign in_9bar = inbar[9];
  assign in_8bar = inbar[8];
  assign in_7bar = inbar[7];
  assign in_6bar = inbar[6];
  assign in_5bar = inbar[5];
  assign in_4bar = inbar[4];
  assign in_3bar = inbar[3];
  assign in_2bar = inbar[2];
  assign in_1bar = inbar[1];
  assign in_0bar = inbar[0];
//assign_done

  OR2_X1 U1 ( .A1(n972), .A2(n971), .ZN(out[7]) );
  AND2_X1 U1bar ( .A1(n972bar), .A2(n971bar), .ZN(outbar[7]) );
  OR2_X1 U2 ( .A1(n970), .A2(n969), .ZN(n971) );
  AND2_X1 U2bar ( .A1(n970bar), .A2(n969bar), .ZN(n971bar) );
  OR2_X1 U3 ( .A1(n968), .A2(n967), .ZN(n969) );
  AND2_X1 U3bar ( .A1(n968bar), .A2(n967bar), .ZN(n969bar) );
  OR2_X1 U4 ( .A1(n966), .A2(n965), .ZN(n967) );
  AND2_X1 U4bar ( .A1(n966bar), .A2(n965bar), .ZN(n967bar) );
  OR2_X1 U5 ( .A1(n964), .A2(n963), .ZN(n968) );
  AND2_X1 U5bar ( .A1(n964bar), .A2(n963bar), .ZN(n968bar) );
  OR2_X1 U6 ( .A1(in[116]), .A2(n962), .ZN(n963) );
  AND2_X1 U6bar ( .A1(inbar[116]), .A2(n962bar), .ZN(n963bar) );
  OR2_X1 U7 ( .A1(n961), .A2(n960), .ZN(n970) );
  AND2_X1 U7bar ( .A1(n961bar), .A2(n960bar), .ZN(n970bar) );
  OR2_X1 U8 ( .A1(in[150]), .A2(in[127]), .ZN(n960) );
  AND2_X1 U8bar ( .A1(inbar[150]), .A2(inbar[127]), .ZN(n960bar) );
  OR2_X1 U9 ( .A1(in[160]), .A2(n959), .ZN(n961) );
  AND2_X1 U9bar ( .A1(inbar[160]), .A2(n959bar), .ZN(n961bar) );
  OR2_X1 U10 ( .A1(in[252]), .A2(in[168]), .ZN(n959) );
  AND2_X1 U10bar ( .A1(inbar[252]), .A2(inbar[168]), .ZN(n959bar) );
  OR2_X1 U11 ( .A1(n958), .A2(n957), .ZN(n972) );
  AND2_X1 U11bar ( .A1(n958bar), .A2(n957bar), .ZN(n972bar) );
  OR2_X1 U12 ( .A1(n956), .A2(n955), .ZN(n957) );
  AND2_X1 U12bar ( .A1(n956bar), .A2(n955bar), .ZN(n957bar) );
  OR2_X1 U13 ( .A1(in_17), .A2(in[96]), .ZN(n955) );
  AND2_X1 U13bar ( .A1(in_17bar), .A2(inbar[96]), .ZN(n955bar) );
  OR2_X1 U14 ( .A1(in_23), .A2(n954), .ZN(n956) );
  AND2_X1 U14bar ( .A1(in_23bar), .A2(n954bar), .ZN(n956bar) );
  OR2_X1 U15 ( .A1(in_31), .A2(in_26), .ZN(n954) );
  AND2_X1 U15bar ( .A1(in_31bar), .A2(in_26bar), .ZN(n954bar) );
  OR2_X1 U16 ( .A1(n953), .A2(n952), .ZN(n958) );
  AND2_X1 U16bar ( .A1(n953bar), .A2(n952bar), .ZN(n958bar) );
  OR2_X1 U17 ( .A1(in_58), .A2(in_4), .ZN(n952) );
  AND2_X1 U17bar ( .A1(in_58bar), .A2(in_4bar), .ZN(n952bar) );
  OR2_X1 U18 ( .A1(in_59), .A2(n951), .ZN(n953) );
  AND2_X1 U18bar ( .A1(in_59bar), .A2(n951bar), .ZN(n953bar) );
  OR2_X1 U19 ( .A1(in_71), .A2(in_62), .ZN(n951) );
  AND2_X1 U19bar ( .A1(in_71bar), .A2(in_62bar), .ZN(n951bar) );
  OR2_X1 U20 ( .A1(n950), .A2(n949), .ZN(out[6]) );
  AND2_X1 U20bar ( .A1(n950bar), .A2(n949bar), .ZN(outbar[6]) );
  OR2_X1 U21 ( .A1(n948), .A2(n947), .ZN(n949) );
  AND2_X1 U21bar ( .A1(n948bar), .A2(n947bar), .ZN(n949bar) );
  OR2_X1 U22 ( .A1(n946), .A2(n945), .ZN(n947) );
  AND2_X1 U22bar ( .A1(n946bar), .A2(n945bar), .ZN(n947bar) );
  OR2_X1 U23 ( .A1(n944), .A2(n943), .ZN(n945) );
  AND2_X1 U23bar ( .A1(n944bar), .A2(n943bar), .ZN(n945bar) );
  OR2_X1 U24 ( .A1(n942), .A2(n941), .ZN(n946) );
  AND2_X1 U24bar ( .A1(n942bar), .A2(n941bar), .ZN(n946bar) );
  OR2_X1 U25 ( .A1(in[101]), .A2(n940), .ZN(n941) );
  AND2_X1 U25bar ( .A1(inbar[101]), .A2(n940bar), .ZN(n941bar) );
  OR2_X1 U26 ( .A1(n939), .A2(n938), .ZN(n948) );
  AND2_X1 U26bar ( .A1(n939bar), .A2(n938bar), .ZN(n948bar) );
  OR2_X1 U27 ( .A1(in[114]), .A2(in[104]), .ZN(n938) );
  AND2_X1 U27bar ( .A1(inbar[114]), .A2(inbar[104]), .ZN(n938bar) );
  OR2_X1 U28 ( .A1(in[128]), .A2(n937), .ZN(n939) );
  AND2_X1 U28bar ( .A1(inbar[128]), .A2(n937bar), .ZN(n939bar) );
  OR2_X1 U29 ( .A1(in[136]), .A2(in[134]), .ZN(n937) );
  AND2_X1 U29bar ( .A1(inbar[136]), .A2(inbar[134]), .ZN(n937bar) );
  OR2_X1 U30 ( .A1(n936), .A2(n935), .ZN(n950) );
  AND2_X1 U30bar ( .A1(n936bar), .A2(n935bar), .ZN(n950bar) );
  OR2_X1 U31 ( .A1(n934), .A2(n933), .ZN(n935) );
  AND2_X1 U31bar ( .A1(n934bar), .A2(n933bar), .ZN(n935bar) );
  OR2_X1 U32 ( .A1(in[177]), .A2(in[164]), .ZN(n933) );
  AND2_X1 U32bar ( .A1(inbar[177]), .A2(inbar[164]), .ZN(n933bar) );
  OR2_X1 U33 ( .A1(in[212]), .A2(n932), .ZN(n934) );
  AND2_X1 U33bar ( .A1(inbar[212]), .A2(n932bar), .ZN(n934bar) );
  OR2_X1 U34 ( .A1(in[248]), .A2(in[221]), .ZN(n932) );
  AND2_X1 U34bar ( .A1(inbar[248]), .A2(inbar[221]), .ZN(n932bar) );
  OR2_X1 U35 ( .A1(n931), .A2(n930), .ZN(n936) );
  AND2_X1 U35bar ( .A1(n931bar), .A2(n930bar), .ZN(n936bar) );
  OR2_X1 U36 ( .A1(in_18), .A2(in[93]), .ZN(n930) );
  AND2_X1 U36bar ( .A1(in_18bar), .A2(inbar[93]), .ZN(n930bar) );
  OR2_X1 U37 ( .A1(in_31), .A2(n929), .ZN(n931) );
  AND2_X1 U37bar ( .A1(in_31bar), .A2(n929bar), .ZN(n931bar) );
  OR2_X1 U38 ( .A1(in_7), .A2(in_39), .ZN(n929) );
  AND2_X1 U38bar ( .A1(in_7bar), .A2(in_39bar), .ZN(n929bar) );
  OR2_X1 U39 ( .A1(n928), .A2(n927), .ZN(out[5]) );
  AND2_X1 U39bar ( .A1(n928bar), .A2(n927bar), .ZN(outbar[5]) );
  OR2_X1 U40 ( .A1(n926), .A2(n925), .ZN(n927) );
  AND2_X1 U40bar ( .A1(n926bar), .A2(n925bar), .ZN(n927bar) );
  OR2_X1 U41 ( .A1(n924), .A2(n923), .ZN(n925) );
  AND2_X1 U41bar ( .A1(n924bar), .A2(n923bar), .ZN(n925bar) );
  OR2_X1 U42 ( .A1(n922), .A2(n921), .ZN(n923) );
  AND2_X1 U42bar ( .A1(n922bar), .A2(n921bar), .ZN(n923bar) );
  OR2_X1 U43 ( .A1(n940), .A2(n920), .ZN(n924) );
  AND2_X1 U43bar ( .A1(n940bar), .A2(n920bar), .ZN(n924bar) );
  OR2_X1 U44 ( .A1(in[111]), .A2(n919), .ZN(n920) );
  AND2_X1 U44bar ( .A1(inbar[111]), .A2(n919bar), .ZN(n920bar) );
  OR2_X1 U45 ( .A1(n918), .A2(n917), .ZN(n940) );
  AND2_X1 U45bar ( .A1(n918bar), .A2(n917bar), .ZN(n940bar) );
  OR2_X1 U46 ( .A1(n916), .A2(n915), .ZN(n917) );
  AND2_X1 U46bar ( .A1(n916bar), .A2(n915bar), .ZN(n917bar) );
  OR2_X1 U47 ( .A1(n914), .A2(n913), .ZN(n915) );
  AND2_X1 U47bar ( .A1(n914bar), .A2(n913bar), .ZN(n915bar) );
  OR2_X1 U48 ( .A1(in[140]), .A2(in[131]), .ZN(n913) );
  AND2_X1 U48bar ( .A1(inbar[140]), .A2(inbar[131]), .ZN(n913bar) );
  OR2_X1 U49 ( .A1(in[160]), .A2(in[144]), .ZN(n914) );
  AND2_X1 U49bar ( .A1(inbar[160]), .A2(inbar[144]), .ZN(n914bar) );
  OR2_X1 U50 ( .A1(n912), .A2(n911), .ZN(n916) );
  AND2_X1 U50bar ( .A1(n912bar), .A2(n911bar), .ZN(n916bar) );
  OR2_X1 U51 ( .A1(in[179]), .A2(in[174]), .ZN(n911) );
  AND2_X1 U51bar ( .A1(inbar[179]), .A2(inbar[174]), .ZN(n911bar) );
  OR2_X1 U52 ( .A1(in[188]), .A2(in[184]), .ZN(n912) );
  AND2_X1 U52bar ( .A1(inbar[188]), .A2(inbar[184]), .ZN(n912bar) );
  OR2_X1 U53 ( .A1(n910), .A2(n909), .ZN(n918) );
  AND2_X1 U53bar ( .A1(n910bar), .A2(n909bar), .ZN(n918bar) );
  OR2_X1 U54 ( .A1(n908), .A2(n907), .ZN(n909) );
  AND2_X1 U54bar ( .A1(n908bar), .A2(n907bar), .ZN(n909bar) );
  OR2_X1 U55 ( .A1(in[216]), .A2(in[200]), .ZN(n907) );
  AND2_X1 U55bar ( .A1(inbar[216]), .A2(inbar[200]), .ZN(n907bar) );
  OR2_X1 U56 ( .A1(in[228]), .A2(in[224]), .ZN(n908) );
  AND2_X1 U56bar ( .A1(inbar[228]), .A2(inbar[224]), .ZN(n908bar) );
  OR2_X1 U57 ( .A1(n906), .A2(n905), .ZN(n910) );
  AND2_X1 U57bar ( .A1(n906bar), .A2(n905bar), .ZN(n910bar) );
  OR2_X1 U58 ( .A1(in[247]), .A2(in[235]), .ZN(n905) );
  AND2_X1 U58bar ( .A1(inbar[247]), .A2(inbar[235]), .ZN(n905bar) );
  OR2_X1 U59 ( .A1(in_42), .A2(in[83]), .ZN(n906) );
  AND2_X1 U59bar ( .A1(in_42bar), .A2(inbar[83]), .ZN(n906bar) );
  OR2_X1 U60 ( .A1(n904), .A2(n903), .ZN(n926) );
  AND2_X1 U60bar ( .A1(n904bar), .A2(n903bar), .ZN(n926bar) );
  OR2_X1 U61 ( .A1(in[166]), .A2(in[123]), .ZN(n903) );
  AND2_X1 U61bar ( .A1(inbar[166]), .A2(inbar[123]), .ZN(n903bar) );
  OR2_X1 U62 ( .A1(in[170]), .A2(n902), .ZN(n904) );
  AND2_X1 U62bar ( .A1(inbar[170]), .A2(n902bar), .ZN(n904bar) );
  OR2_X1 U63 ( .A1(in[194]), .A2(in[183]), .ZN(n902) );
  AND2_X1 U63bar ( .A1(inbar[194]), .A2(inbar[183]), .ZN(n902bar) );
  OR2_X1 U64 ( .A1(n901), .A2(n900), .ZN(n928) );
  AND2_X1 U64bar ( .A1(n901bar), .A2(n900bar), .ZN(n928bar) );
  OR2_X1 U65 ( .A1(n899), .A2(n898), .ZN(n900) );
  AND2_X1 U65bar ( .A1(n899bar), .A2(n898bar), .ZN(n900bar) );
  OR2_X1 U66 ( .A1(in[241]), .A2(in[238]), .ZN(n898) );
  AND2_X1 U66bar ( .A1(inbar[241]), .A2(inbar[238]), .ZN(n898bar) );
  OR2_X1 U67 ( .A1(in[250]), .A2(n897), .ZN(n899) );
  AND2_X1 U67bar ( .A1(inbar[250]), .A2(n897bar), .ZN(n899bar) );
  OR2_X1 U68 ( .A1(in_24), .A2(in[84]), .ZN(n897) );
  AND2_X1 U68bar ( .A1(in_24bar), .A2(inbar[84]), .ZN(n897bar) );
  OR2_X1 U69 ( .A1(n896), .A2(n895), .ZN(n901) );
  AND2_X1 U69bar ( .A1(n896bar), .A2(n895bar), .ZN(n901bar) );
  OR2_X1 U70 ( .A1(in_41), .A2(in_29), .ZN(n895) );
  AND2_X1 U70bar ( .A1(in_41bar), .A2(in_29bar), .ZN(n895bar) );
  OR2_X1 U71 ( .A1(in_66), .A2(n894), .ZN(n896) );
  AND2_X1 U71bar ( .A1(in_66bar), .A2(n894bar), .ZN(n896bar) );
  OR2_X1 U72 ( .A1(in_76), .A2(in_71), .ZN(n894) );
  AND2_X1 U72bar ( .A1(in_76bar), .A2(in_71bar), .ZN(n894bar) );
  OR2_X1 U73 ( .A1(n893), .A2(n892), .ZN(out[4]) );
  AND2_X1 U73bar ( .A1(n893bar), .A2(n892bar), .ZN(outbar[4]) );
  OR2_X1 U74 ( .A1(n891), .A2(n890), .ZN(n892) );
  AND2_X1 U74bar ( .A1(n891bar), .A2(n890bar), .ZN(n892bar) );
  OR2_X1 U75 ( .A1(n889), .A2(n888), .ZN(n890) );
  AND2_X1 U75bar ( .A1(n889bar), .A2(n888bar), .ZN(n890bar) );
  OR2_X1 U76 ( .A1(n922), .A2(n887), .ZN(n888) );
  AND2_X1 U76bar ( .A1(n922bar), .A2(n887bar), .ZN(n888bar) );
  OR2_X1 U77 ( .A1(n886), .A2(n885), .ZN(n922) );
  AND2_X1 U77bar ( .A1(n886bar), .A2(n885bar), .ZN(n922bar) );
  OR2_X1 U78 ( .A1(n884), .A2(n883), .ZN(n885) );
  AND2_X1 U78bar ( .A1(n884bar), .A2(n883bar), .ZN(n885bar) );
  OR2_X1 U79 ( .A1(n882), .A2(n881), .ZN(n883) );
  AND2_X1 U79bar ( .A1(n882bar), .A2(n881bar), .ZN(n883bar) );
  OR2_X1 U80 ( .A1(in[118]), .A2(in[109]), .ZN(n881) );
  AND2_X1 U80bar ( .A1(inbar[118]), .A2(inbar[109]), .ZN(n881bar) );
  OR2_X1 U81 ( .A1(in[139]), .A2(in[120]), .ZN(n882) );
  AND2_X1 U81bar ( .A1(inbar[139]), .A2(inbar[120]), .ZN(n882bar) );
  OR2_X1 U82 ( .A1(n880), .A2(n879), .ZN(n884) );
  AND2_X1 U82bar ( .A1(n880bar), .A2(n879bar), .ZN(n884bar) );
  OR2_X1 U83 ( .A1(in[198]), .A2(in[154]), .ZN(n879) );
  AND2_X1 U83bar ( .A1(inbar[198]), .A2(inbar[154]), .ZN(n879bar) );
  OR2_X1 U84 ( .A1(in[210]), .A2(in[205]), .ZN(n880) );
  AND2_X1 U84bar ( .A1(inbar[210]), .A2(inbar[205]), .ZN(n880bar) );
  OR2_X1 U85 ( .A1(n878), .A2(n877), .ZN(n886) );
  AND2_X1 U85bar ( .A1(n878bar), .A2(n877bar), .ZN(n886bar) );
  OR2_X1 U86 ( .A1(n876), .A2(n875), .ZN(n877) );
  AND2_X1 U86bar ( .A1(n876bar), .A2(n875bar), .ZN(n877bar) );
  OR2_X1 U87 ( .A1(in[219]), .A2(in[217]), .ZN(n875) );
  AND2_X1 U87bar ( .A1(inbar[219]), .A2(inbar[217]), .ZN(n875bar) );
  OR2_X1 U88 ( .A1(in[86]), .A2(in[252]), .ZN(n876) );
  AND2_X1 U88bar ( .A1(inbar[86]), .A2(inbar[252]), .ZN(n876bar) );
  OR2_X1 U89 ( .A1(n874), .A2(n873), .ZN(n878) );
  AND2_X1 U89bar ( .A1(n874bar), .A2(n873bar), .ZN(n878bar) );
  OR2_X1 U90 ( .A1(in_40), .A2(in[91]), .ZN(n873) );
  AND2_X1 U90bar ( .A1(in_40bar), .A2(inbar[91]), .ZN(n873bar) );
  OR2_X1 U91 ( .A1(in_8), .A2(in_46), .ZN(n874) );
  AND2_X1 U91bar ( .A1(in_8bar), .A2(in_46bar), .ZN(n874bar) );
  OR2_X1 U92 ( .A1(n872), .A2(n871), .ZN(n889) );
  AND2_X1 U92bar ( .A1(n872bar), .A2(n871bar), .ZN(n889bar) );
  OR2_X1 U93 ( .A1(in[117]), .A2(n943), .ZN(n871) );
  AND2_X1 U93bar ( .A1(inbar[117]), .A2(n943bar), .ZN(n871bar) );
  OR2_X1 U94 ( .A1(n870), .A2(n869), .ZN(n943) );
  AND2_X1 U94bar ( .A1(n870bar), .A2(n869bar), .ZN(n943bar) );
  OR2_X1 U95 ( .A1(n868), .A2(n867), .ZN(n869) );
  AND2_X1 U95bar ( .A1(n868bar), .A2(n867bar), .ZN(n869bar) );
  OR2_X1 U96 ( .A1(n866), .A2(n865), .ZN(n867) );
  AND2_X1 U96bar ( .A1(n866bar), .A2(n865bar), .ZN(n867bar) );
  OR2_X1 U97 ( .A1(n864), .A2(n863), .ZN(n865) );
  AND2_X1 U97bar ( .A1(n864bar), .A2(n863bar), .ZN(n865bar) );
  OR2_X1 U98 ( .A1(in[108]), .A2(n919), .ZN(n866) );
  AND2_X1 U98bar ( .A1(inbar[108]), .A2(n919bar), .ZN(n866bar) );
  OR2_X1 U99 ( .A1(n862), .A2(n861), .ZN(n919) );
  AND2_X1 U99bar ( .A1(n862bar), .A2(n861bar), .ZN(n919bar) );
  OR2_X1 U100 ( .A1(n860), .A2(n859), .ZN(n861) );
  AND2_X1 U100bar ( .A1(n860bar), .A2(n859bar), .ZN(n861bar) );
  OR2_X1 U101 ( .A1(n858), .A2(n857), .ZN(n859) );
  AND2_X1 U101bar ( .A1(n858bar), .A2(n857bar), .ZN(n859bar) );
  OR2_X1 U102 ( .A1(in[119]), .A2(in[105]), .ZN(n857) );
  AND2_X1 U102bar ( .A1(inbar[119]), .A2(inbar[105]), .ZN(n857bar) );
  OR2_X1 U103 ( .A1(in[186]), .A2(in[175]), .ZN(n858) );
  AND2_X1 U103bar ( .A1(inbar[186]), .A2(inbar[175]), .ZN(n858bar) );
  OR2_X1 U104 ( .A1(n856), .A2(n855), .ZN(n860) );
  AND2_X1 U104bar ( .A1(n856bar), .A2(n855bar), .ZN(n860bar) );
  OR2_X1 U105 ( .A1(in[202]), .A2(in[193]), .ZN(n855) );
  AND2_X1 U105bar ( .A1(inbar[202]), .A2(inbar[193]), .ZN(n855bar) );
  OR2_X1 U106 ( .A1(in[225]), .A2(in[208]), .ZN(n856) );
  AND2_X1 U106bar ( .A1(inbar[225]), .A2(inbar[208]), .ZN(n856bar) );
  OR2_X1 U107 ( .A1(n854), .A2(n853), .ZN(n862) );
  AND2_X1 U107bar ( .A1(n854bar), .A2(n853bar), .ZN(n862bar) );
  OR2_X1 U108 ( .A1(n852), .A2(n851), .ZN(n853) );
  AND2_X1 U108bar ( .A1(n852bar), .A2(n851bar), .ZN(n853bar) );
  OR2_X1 U109 ( .A1(in_1), .A2(in[85]), .ZN(n851) );
  AND2_X1 U109bar ( .A1(in_1bar), .A2(inbar[85]), .ZN(n851bar) );
  OR2_X1 U110 ( .A1(in_23), .A2(in_19), .ZN(n852) );
  AND2_X1 U110bar ( .A1(in_23bar), .A2(in_19bar), .ZN(n852bar) );
  OR2_X1 U111 ( .A1(n850), .A2(n849), .ZN(n854) );
  AND2_X1 U111bar ( .A1(n850bar), .A2(n849bar), .ZN(n854bar) );
  OR2_X1 U112 ( .A1(in_43), .A2(in_33), .ZN(n849) );
  AND2_X1 U112bar ( .A1(in_43bar), .A2(in_33bar), .ZN(n849bar) );
  OR2_X1 U113 ( .A1(in_63), .A2(in_44), .ZN(n850) );
  AND2_X1 U113bar ( .A1(in_63bar), .A2(in_44bar), .ZN(n850bar) );
  OR2_X1 U114 ( .A1(n848), .A2(n847), .ZN(n868) );
  AND2_X1 U114bar ( .A1(n848bar), .A2(n847bar), .ZN(n868bar) );
  OR2_X1 U115 ( .A1(in[141]), .A2(in[112]), .ZN(n847) );
  AND2_X1 U115bar ( .A1(inbar[141]), .A2(inbar[112]), .ZN(n847bar) );
  OR2_X1 U116 ( .A1(in[147]), .A2(n846), .ZN(n848) );
  AND2_X1 U116bar ( .A1(inbar[147]), .A2(n846bar), .ZN(n848bar) );
  OR2_X1 U117 ( .A1(in[181]), .A2(in[167]), .ZN(n846) );
  AND2_X1 U117bar ( .A1(inbar[181]), .A2(inbar[167]), .ZN(n846bar) );
  OR2_X1 U118 ( .A1(n845), .A2(n844), .ZN(n870) );
  AND2_X1 U118bar ( .A1(n845bar), .A2(n844bar), .ZN(n870bar) );
  OR2_X1 U119 ( .A1(n843), .A2(n842), .ZN(n844) );
  AND2_X1 U119bar ( .A1(n843bar), .A2(n842bar), .ZN(n844bar) );
  OR2_X1 U120 ( .A1(in[229]), .A2(in[201]), .ZN(n842) );
  AND2_X1 U120bar ( .A1(inbar[229]), .A2(inbar[201]), .ZN(n842bar) );
  OR2_X1 U121 ( .A1(in[237]), .A2(n841), .ZN(n843) );
  AND2_X1 U121bar ( .A1(inbar[237]), .A2(n841bar), .ZN(n843bar) );
  OR2_X1 U122 ( .A1(in[94]), .A2(in[253]), .ZN(n841) );
  AND2_X1 U122bar ( .A1(inbar[94]), .A2(inbar[253]), .ZN(n841bar) );
  OR2_X1 U123 ( .A1(n840), .A2(n839), .ZN(n845) );
  AND2_X1 U123bar ( .A1(n840bar), .A2(n839bar), .ZN(n845bar) );
  OR2_X1 U124 ( .A1(in_21), .A2(in[96]), .ZN(n839) );
  AND2_X1 U124bar ( .A1(in_21bar), .A2(inbar[96]), .ZN(n839bar) );
  OR2_X1 U125 ( .A1(in_25), .A2(n838), .ZN(n840) );
  AND2_X1 U125bar ( .A1(in_25bar), .A2(n838bar), .ZN(n840bar) );
  OR2_X1 U126 ( .A1(in_81), .A2(in_45), .ZN(n838) );
  AND2_X1 U126bar ( .A1(in_81bar), .A2(in_45bar), .ZN(n838bar) );
  OR2_X1 U127 ( .A1(n837), .A2(n836), .ZN(n891) );
  AND2_X1 U127bar ( .A1(n837bar), .A2(n836bar), .ZN(n891bar) );
  OR2_X1 U128 ( .A1(in[142]), .A2(in[124]), .ZN(n836) );
  AND2_X1 U128bar ( .A1(inbar[142]), .A2(inbar[124]), .ZN(n836bar) );
  OR2_X1 U129 ( .A1(in[150]), .A2(n835), .ZN(n837) );
  AND2_X1 U129bar ( .A1(inbar[150]), .A2(n835bar), .ZN(n837bar) );
  OR2_X1 U130 ( .A1(in[172]), .A2(in[155]), .ZN(n835) );
  AND2_X1 U130bar ( .A1(inbar[172]), .A2(inbar[155]), .ZN(n835bar) );
  OR2_X1 U131 ( .A1(n834), .A2(n833), .ZN(n893) );
  AND2_X1 U131bar ( .A1(n834bar), .A2(n833bar), .ZN(n893bar) );
  OR2_X1 U132 ( .A1(n832), .A2(n831), .ZN(n833) );
  AND2_X1 U132bar ( .A1(n832bar), .A2(n831bar), .ZN(n833bar) );
  OR2_X1 U133 ( .A1(in[196]), .A2(in[173]), .ZN(n831) );
  AND2_X1 U133bar ( .A1(inbar[196]), .A2(inbar[173]), .ZN(n831bar) );
  OR2_X1 U134 ( .A1(in[222]), .A2(n830), .ZN(n832) );
  AND2_X1 U134bar ( .A1(inbar[222]), .A2(n830bar), .ZN(n832bar) );
  OR2_X1 U135 ( .A1(in[227]), .A2(in[226]), .ZN(n830) );
  AND2_X1 U135bar ( .A1(inbar[227]), .A2(inbar[226]), .ZN(n830bar) );
  OR2_X1 U136 ( .A1(n829), .A2(n828), .ZN(n834) );
  AND2_X1 U136bar ( .A1(n829bar), .A2(n828bar), .ZN(n834bar) );
  OR2_X1 U137 ( .A1(in[249]), .A2(in[231]), .ZN(n828) );
  AND2_X1 U137bar ( .A1(inbar[249]), .A2(inbar[231]), .ZN(n828bar) );
  OR2_X1 U138 ( .A1(in_28), .A2(n827), .ZN(n829) );
  AND2_X1 U138bar ( .A1(in_28bar), .A2(n827bar), .ZN(n829bar) );
  OR2_X1 U139 ( .A1(in_52), .A2(in_47), .ZN(n827) );
  AND2_X1 U139bar ( .A1(in_52bar), .A2(in_47bar), .ZN(n827bar) );
  OR2_X1 U140 ( .A1(n826), .A2(n825), .ZN(out[3]) );
  AND2_X1 U140bar ( .A1(n826bar), .A2(n825bar), .ZN(outbar[3]) );
  OR2_X1 U141 ( .A1(n824), .A2(n823), .ZN(n825) );
  AND2_X1 U141bar ( .A1(n824bar), .A2(n823bar), .ZN(n825bar) );
  OR2_X1 U142 ( .A1(n822), .A2(n821), .ZN(n823) );
  AND2_X1 U142bar ( .A1(n822bar), .A2(n821bar), .ZN(n823bar) );
  OR2_X1 U143 ( .A1(n820), .A2(n819), .ZN(n821) );
  AND2_X1 U143bar ( .A1(n820bar), .A2(n819bar), .ZN(n821bar) );
  OR2_X1 U144 ( .A1(n964), .A2(n818), .ZN(n822) );
  AND2_X1 U144bar ( .A1(n964bar), .A2(n818bar), .ZN(n822bar) );
  OR2_X1 U145 ( .A1(in[118]), .A2(n817), .ZN(n818) );
  AND2_X1 U145bar ( .A1(inbar[118]), .A2(n817bar), .ZN(n818bar) );
  OR2_X1 U146 ( .A1(n816), .A2(n815), .ZN(n964) );
  AND2_X1 U146bar ( .A1(n816bar), .A2(n815bar), .ZN(n964bar) );
  OR2_X1 U147 ( .A1(n814), .A2(n813), .ZN(n815) );
  AND2_X1 U147bar ( .A1(n814bar), .A2(n813bar), .ZN(n815bar) );
  OR2_X1 U148 ( .A1(n812), .A2(n811), .ZN(n813) );
  AND2_X1 U148bar ( .A1(n812bar), .A2(n811bar), .ZN(n813bar) );
  OR2_X1 U149 ( .A1(in[122]), .A2(in[111]), .ZN(n811) );
  AND2_X1 U149bar ( .A1(inbar[122]), .A2(inbar[111]), .ZN(n811bar) );
  OR2_X1 U150 ( .A1(in[154]), .A2(in[151]), .ZN(n812) );
  AND2_X1 U150bar ( .A1(inbar[154]), .A2(inbar[151]), .ZN(n812bar) );
  OR2_X1 U151 ( .A1(n810), .A2(n809), .ZN(n814) );
  AND2_X1 U151bar ( .A1(n810bar), .A2(n809bar), .ZN(n814bar) );
  OR2_X1 U152 ( .A1(in[187]), .A2(in[177]), .ZN(n809) );
  AND2_X1 U152bar ( .A1(inbar[187]), .A2(inbar[177]), .ZN(n809bar) );
  OR2_X1 U153 ( .A1(in[200]), .A2(in[192]), .ZN(n810) );
  AND2_X1 U153bar ( .A1(inbar[200]), .A2(inbar[192]), .ZN(n810bar) );
  OR2_X1 U154 ( .A1(n808), .A2(n807), .ZN(n816) );
  AND2_X1 U154bar ( .A1(n808bar), .A2(n807bar), .ZN(n816bar) );
  OR2_X1 U155 ( .A1(n806), .A2(n805), .ZN(n807) );
  AND2_X1 U155bar ( .A1(n806bar), .A2(n805bar), .ZN(n807bar) );
  OR2_X1 U156 ( .A1(in[225]), .A2(in[207]), .ZN(n805) );
  AND2_X1 U156bar ( .A1(inbar[225]), .A2(inbar[207]), .ZN(n805bar) );
  OR2_X1 U157 ( .A1(in[98]), .A2(in[226]), .ZN(n806) );
  AND2_X1 U157bar ( .A1(inbar[98]), .A2(inbar[226]), .ZN(n806bar) );
  OR2_X1 U158 ( .A1(n804), .A2(n803), .ZN(n808) );
  AND2_X1 U158bar ( .A1(n804bar), .A2(n803bar), .ZN(n808bar) );
  OR2_X1 U159 ( .A1(in_20), .A2(in_16), .ZN(n803) );
  AND2_X1 U159bar ( .A1(in_20bar), .A2(in_16bar), .ZN(n803bar) );
  OR2_X1 U160 ( .A1(in_55), .A2(in_45), .ZN(n804) );
  AND2_X1 U160bar ( .A1(in_55bar), .A2(in_45bar), .ZN(n804bar) );
  OR2_X1 U161 ( .A1(n802), .A2(n801), .ZN(n824) );
  AND2_X1 U161bar ( .A1(n802bar), .A2(n801bar), .ZN(n824bar) );
  OR2_X1 U162 ( .A1(in[162]), .A2(in[149]), .ZN(n801) );
  AND2_X1 U162bar ( .A1(inbar[162]), .A2(inbar[149]), .ZN(n801bar) );
  OR2_X1 U163 ( .A1(in[163]), .A2(n800), .ZN(n802) );
  AND2_X1 U163bar ( .A1(inbar[163]), .A2(n800bar), .ZN(n802bar) );
  OR2_X1 U164 ( .A1(in[191]), .A2(in[189]), .ZN(n800) );
  AND2_X1 U164bar ( .A1(inbar[191]), .A2(inbar[189]), .ZN(n800bar) );
  OR2_X1 U165 ( .A1(n799), .A2(n798), .ZN(n826) );
  AND2_X1 U165bar ( .A1(n799bar), .A2(n798bar), .ZN(n826bar) );
  OR2_X1 U166 ( .A1(n797), .A2(n796), .ZN(n798) );
  AND2_X1 U166bar ( .A1(n797bar), .A2(n796bar), .ZN(n798bar) );
  OR2_X1 U167 ( .A1(in[212]), .A2(in[193]), .ZN(n796) );
  AND2_X1 U167bar ( .A1(inbar[212]), .A2(inbar[193]), .ZN(n796bar) );
  OR2_X1 U168 ( .A1(in[238]), .A2(n795), .ZN(n797) );
  AND2_X1 U168bar ( .A1(inbar[238]), .A2(n795bar), .ZN(n797bar) );
  OR2_X1 U169 ( .A1(in[88]), .A2(in[247]), .ZN(n795) );
  AND2_X1 U169bar ( .A1(inbar[88]), .A2(inbar[247]), .ZN(n795bar) );
  OR2_X1 U170 ( .A1(n794), .A2(n793), .ZN(n799) );
  AND2_X1 U170bar ( .A1(n794bar), .A2(n793bar), .ZN(n799bar) );
  OR2_X1 U171 ( .A1(in[94]), .A2(in[92]), .ZN(n793) );
  AND2_X1 U171bar ( .A1(inbar[94]), .A2(inbar[92]), .ZN(n793bar) );
  OR2_X1 U172 ( .A1(in_52), .A2(n792), .ZN(n794) );
  AND2_X1 U172bar ( .A1(in_52bar), .A2(n792bar), .ZN(n794bar) );
  OR2_X1 U173 ( .A1(in_70), .A2(in_67), .ZN(n792) );
  AND2_X1 U173bar ( .A1(in_70bar), .A2(in_67bar), .ZN(n792bar) );
  OR2_X1 U174 ( .A1(n791), .A2(n790), .ZN(out[2]) );
  AND2_X1 U174bar ( .A1(n791bar), .A2(n790bar), .ZN(outbar[2]) );
  OR2_X1 U175 ( .A1(n789), .A2(n788), .ZN(n790) );
  AND2_X1 U175bar ( .A1(n789bar), .A2(n788bar), .ZN(n790bar) );
  OR2_X1 U176 ( .A1(n787), .A2(n786), .ZN(n788) );
  AND2_X1 U176bar ( .A1(n787bar), .A2(n786bar), .ZN(n788bar) );
  OR2_X1 U177 ( .A1(n819), .A2(n785), .ZN(n786) );
  AND2_X1 U177bar ( .A1(n819bar), .A2(n785bar), .ZN(n786bar) );
  OR2_X1 U178 ( .A1(n784), .A2(n783), .ZN(n819) );
  AND2_X1 U178bar ( .A1(n784bar), .A2(n783bar), .ZN(n819bar) );
  OR2_X1 U179 ( .A1(n782), .A2(n781), .ZN(n783) );
  AND2_X1 U179bar ( .A1(n782bar), .A2(n781bar), .ZN(n783bar) );
  OR2_X1 U180 ( .A1(n780), .A2(n779), .ZN(n781) );
  AND2_X1 U180bar ( .A1(n780bar), .A2(n779bar), .ZN(n781bar) );
  OR2_X1 U181 ( .A1(n962), .A2(n778), .ZN(n779) );
  AND2_X1 U181bar ( .A1(n962bar), .A2(n778bar), .ZN(n779bar) );
  OR2_X1 U182 ( .A1(n777), .A2(n776), .ZN(n962) );
  AND2_X1 U182bar ( .A1(n777bar), .A2(n776bar), .ZN(n962bar) );
  OR2_X1 U183 ( .A1(n775), .A2(n774), .ZN(n776) );
  AND2_X1 U183bar ( .A1(n775bar), .A2(n774bar), .ZN(n776bar) );
  OR2_X1 U184 ( .A1(n773), .A2(n772), .ZN(n774) );
  AND2_X1 U184bar ( .A1(n773bar), .A2(n772bar), .ZN(n774bar) );
  OR2_X1 U185 ( .A1(in[131]), .A2(in[120]), .ZN(n772) );
  AND2_X1 U185bar ( .A1(inbar[131]), .A2(inbar[120]), .ZN(n772bar) );
  OR2_X1 U186 ( .A1(in[153]), .A2(in[147]), .ZN(n773) );
  AND2_X1 U186bar ( .A1(inbar[153]), .A2(inbar[147]), .ZN(n773bar) );
  OR2_X1 U187 ( .A1(n771), .A2(n770), .ZN(n775) );
  AND2_X1 U187bar ( .A1(n771bar), .A2(n770bar), .ZN(n775bar) );
  OR2_X1 U188 ( .A1(in[170]), .A2(in[156]), .ZN(n770) );
  AND2_X1 U188bar ( .A1(inbar[170]), .A2(inbar[156]), .ZN(n770bar) );
  OR2_X1 U189 ( .A1(in[223]), .A2(in[190]), .ZN(n771) );
  AND2_X1 U189bar ( .A1(inbar[223]), .A2(inbar[190]), .ZN(n771bar) );
  OR2_X1 U190 ( .A1(n769), .A2(n768), .ZN(n777) );
  AND2_X1 U190bar ( .A1(n769bar), .A2(n768bar), .ZN(n777bar) );
  OR2_X1 U191 ( .A1(n767), .A2(n766), .ZN(n768) );
  AND2_X1 U191bar ( .A1(n767bar), .A2(n766bar), .ZN(n768bar) );
  OR2_X1 U192 ( .A1(in[236]), .A2(in[230]), .ZN(n766) );
  AND2_X1 U192bar ( .A1(inbar[236]), .A2(inbar[230]), .ZN(n766bar) );
  OR2_X1 U193 ( .A1(in[85]), .A2(in[240]), .ZN(n767) );
  AND2_X1 U193bar ( .A1(inbar[85]), .A2(inbar[240]), .ZN(n767bar) );
  OR2_X1 U194 ( .A1(n765), .A2(n764), .ZN(n769) );
  AND2_X1 U194bar ( .A1(n765bar), .A2(n764bar), .ZN(n769bar) );
  OR2_X1 U195 ( .A1(in_12), .A2(in[90]), .ZN(n764) );
  AND2_X1 U195bar ( .A1(in_12bar), .A2(inbar[90]), .ZN(n764bar) );
  OR2_X1 U196 ( .A1(in_39), .A2(in_28), .ZN(n765) );
  AND2_X1 U196bar ( .A1(in_39bar), .A2(in_28bar), .ZN(n765bar) );
  OR2_X1 U197 ( .A1(in[109]), .A2(n763), .ZN(n780) );
  AND2_X1 U197bar ( .A1(inbar[109]), .A2(n763bar), .ZN(n780bar) );
  OR2_X1 U198 ( .A1(n762), .A2(n761), .ZN(n782) );
  AND2_X1 U198bar ( .A1(n762bar), .A2(n761bar), .ZN(n782bar) );
  OR2_X1 U199 ( .A1(in[138]), .A2(in[129]), .ZN(n761) );
  AND2_X1 U199bar ( .A1(inbar[138]), .A2(inbar[129]), .ZN(n761bar) );
  OR2_X1 U200 ( .A1(in[157]), .A2(n760), .ZN(n762) );
  AND2_X1 U200bar ( .A1(inbar[157]), .A2(n760bar), .ZN(n762bar) );
  OR2_X1 U201 ( .A1(in[182]), .A2(in[167]), .ZN(n760) );
  AND2_X1 U201bar ( .A1(inbar[182]), .A2(inbar[167]), .ZN(n760bar) );
  OR2_X1 U202 ( .A1(n759), .A2(n758), .ZN(n784) );
  AND2_X1 U202bar ( .A1(n759bar), .A2(n758bar), .ZN(n784bar) );
  OR2_X1 U203 ( .A1(n757), .A2(n756), .ZN(n758) );
  AND2_X1 U203bar ( .A1(n757bar), .A2(n756bar), .ZN(n758bar) );
  OR2_X1 U204 ( .A1(in[195]), .A2(in[184]), .ZN(n756) );
  AND2_X1 U204bar ( .A1(inbar[195]), .A2(inbar[184]), .ZN(n756bar) );
  OR2_X1 U205 ( .A1(in[196]), .A2(n755), .ZN(n757) );
  AND2_X1 U205bar ( .A1(inbar[196]), .A2(n755bar), .ZN(n757bar) );
  OR2_X1 U206 ( .A1(in[215]), .A2(in[209]), .ZN(n755) );
  AND2_X1 U206bar ( .A1(inbar[215]), .A2(inbar[209]), .ZN(n755bar) );
  OR2_X1 U207 ( .A1(n754), .A2(n753), .ZN(n759) );
  AND2_X1 U207bar ( .A1(n754bar), .A2(n753bar), .ZN(n759bar) );
  OR2_X1 U208 ( .A1(in[93]), .A2(in[233]), .ZN(n753) );
  AND2_X1 U208bar ( .A1(inbar[93]), .A2(inbar[233]), .ZN(n753bar) );
  OR2_X1 U209 ( .A1(in_1), .A2(n752), .ZN(n754) );
  AND2_X1 U209bar ( .A1(in_1bar), .A2(n752bar), .ZN(n754bar) );
  OR2_X1 U210 ( .A1(in_69), .A2(in_66), .ZN(n752) );
  AND2_X1 U210bar ( .A1(in_69bar), .A2(in_66bar), .ZN(n752bar) );
  OR2_X1 U211 ( .A1(n966), .A2(n751), .ZN(n787) );
  AND2_X1 U211bar ( .A1(n966bar), .A2(n751bar), .ZN(n787bar) );
  OR2_X1 U212 ( .A1(in[134]), .A2(n750), .ZN(n751) );
  AND2_X1 U212bar ( .A1(inbar[134]), .A2(n750bar), .ZN(n751bar) );
  OR2_X1 U213 ( .A1(n749), .A2(n748), .ZN(n966) );
  AND2_X1 U213bar ( .A1(n749bar), .A2(n748bar), .ZN(n966bar) );
  OR2_X1 U214 ( .A1(n747), .A2(n746), .ZN(n748) );
  AND2_X1 U214bar ( .A1(n747bar), .A2(n746bar), .ZN(n748bar) );
  OR2_X1 U215 ( .A1(n745), .A2(n744), .ZN(n746) );
  AND2_X1 U215bar ( .A1(n745bar), .A2(n744bar), .ZN(n746bar) );
  OR2_X1 U216 ( .A1(in[136]), .A2(in[121]), .ZN(n744) );
  AND2_X1 U216bar ( .A1(inbar[136]), .A2(inbar[121]), .ZN(n744bar) );
  OR2_X1 U217 ( .A1(in[186]), .A2(in[174]), .ZN(n745) );
  AND2_X1 U217bar ( .A1(inbar[186]), .A2(inbar[174]), .ZN(n745bar) );
  OR2_X1 U218 ( .A1(n743), .A2(n742), .ZN(n747) );
  AND2_X1 U218bar ( .A1(n743bar), .A2(n742bar), .ZN(n747bar) );
  OR2_X1 U219 ( .A1(in[198]), .A2(in[197]), .ZN(n742) );
  AND2_X1 U219bar ( .A1(inbar[198]), .A2(inbar[197]), .ZN(n742bar) );
  OR2_X1 U220 ( .A1(in[214]), .A2(in[199]), .ZN(n743) );
  AND2_X1 U220bar ( .A1(inbar[214]), .A2(inbar[199]), .ZN(n743bar) );
  OR2_X1 U221 ( .A1(n741), .A2(n740), .ZN(n749) );
  AND2_X1 U221bar ( .A1(n741bar), .A2(n740bar), .ZN(n749bar) );
  OR2_X1 U222 ( .A1(n739), .A2(n738), .ZN(n740) );
  AND2_X1 U222bar ( .A1(n739bar), .A2(n738bar), .ZN(n740bar) );
  OR2_X1 U223 ( .A1(in[231]), .A2(in[220]), .ZN(n738) );
  AND2_X1 U223bar ( .A1(inbar[231]), .A2(inbar[220]), .ZN(n738bar) );
  OR2_X1 U224 ( .A1(in_25), .A2(in[245]), .ZN(n739) );
  AND2_X1 U224bar ( .A1(in_25bar), .A2(inbar[245]), .ZN(n739bar) );
  OR2_X1 U225 ( .A1(n737), .A2(n736), .ZN(n741) );
  AND2_X1 U225bar ( .A1(n737bar), .A2(n736bar), .ZN(n741bar) );
  OR2_X1 U226 ( .A1(in_53), .A2(in_29), .ZN(n736) );
  AND2_X1 U226bar ( .A1(in_53bar), .A2(in_29bar), .ZN(n736bar) );
  OR2_X1 U227 ( .A1(in_79), .A2(in_74), .ZN(n737) );
  AND2_X1 U227bar ( .A1(in_79bar), .A2(in_74bar), .ZN(n737bar) );
  OR2_X1 U228 ( .A1(n735), .A2(n734), .ZN(n789) );
  AND2_X1 U228bar ( .A1(n735bar), .A2(n734bar), .ZN(n789bar) );
  OR2_X1 U229 ( .A1(in[152]), .A2(in[140]), .ZN(n734) );
  AND2_X1 U229bar ( .A1(inbar[152]), .A2(inbar[140]), .ZN(n734bar) );
  OR2_X1 U230 ( .A1(in[155]), .A2(n733), .ZN(n735) );
  AND2_X1 U230bar ( .A1(inbar[155]), .A2(n733bar), .ZN(n735bar) );
  OR2_X1 U231 ( .A1(in[166]), .A2(in[165]), .ZN(n733) );
  AND2_X1 U231bar ( .A1(inbar[166]), .A2(inbar[165]), .ZN(n733bar) );
  OR2_X1 U232 ( .A1(n732), .A2(n731), .ZN(n791) );
  AND2_X1 U232bar ( .A1(n732bar), .A2(n731bar), .ZN(n791bar) );
  OR2_X1 U233 ( .A1(n730), .A2(n729), .ZN(n731) );
  AND2_X1 U233bar ( .A1(n730bar), .A2(n729bar), .ZN(n731bar) );
  OR2_X1 U234 ( .A1(in[202]), .A2(in[185]), .ZN(n729) );
  AND2_X1 U234bar ( .A1(inbar[202]), .A2(inbar[185]), .ZN(n729bar) );
  OR2_X1 U235 ( .A1(in[211]), .A2(n728), .ZN(n730) );
  AND2_X1 U235bar ( .A1(inbar[211]), .A2(n728bar), .ZN(n730bar) );
  OR2_X1 U236 ( .A1(in[255]), .A2(in[253]), .ZN(n728) );
  AND2_X1 U236bar ( .A1(inbar[255]), .A2(inbar[253]), .ZN(n728bar) );
  OR2_X1 U237 ( .A1(n727), .A2(n726), .ZN(n732) );
  AND2_X1 U237bar ( .A1(n727bar), .A2(n726bar), .ZN(n732bar) );
  OR2_X1 U238 ( .A1(in_35), .A2(in_15), .ZN(n726) );
  AND2_X1 U238bar ( .A1(in_35bar), .A2(in_15bar), .ZN(n726bar) );
  OR2_X1 U239 ( .A1(in_36), .A2(n725), .ZN(n727) );
  AND2_X1 U239bar ( .A1(in_36bar), .A2(n725bar), .ZN(n727bar) );
  OR2_X1 U240 ( .A1(in_48), .A2(in_40), .ZN(n725) );
  AND2_X1 U240bar ( .A1(in_48bar), .A2(in_40bar), .ZN(n725bar) );
  OR2_X1 U241 ( .A1(n724), .A2(n723), .ZN(out[1]) );
  AND2_X1 U241bar ( .A1(n724bar), .A2(n723bar), .ZN(outbar[1]) );
  OR2_X1 U242 ( .A1(n722), .A2(n721), .ZN(n723) );
  AND2_X1 U242bar ( .A1(n722bar), .A2(n721bar), .ZN(n723bar) );
  OR2_X1 U243 ( .A1(n720), .A2(n719), .ZN(n721) );
  AND2_X1 U243bar ( .A1(n720bar), .A2(n719bar), .ZN(n721bar) );
  OR2_X1 U244 ( .A1(n921), .A2(n887), .ZN(n719) );
  AND2_X1 U244bar ( .A1(n921bar), .A2(n887bar), .ZN(n719bar) );
  OR2_X1 U245 ( .A1(n718), .A2(n717), .ZN(n887) );
  AND2_X1 U245bar ( .A1(n718bar), .A2(n717bar), .ZN(n887bar) );
  OR2_X1 U246 ( .A1(n716), .A2(n715), .ZN(n717) );
  AND2_X1 U246bar ( .A1(n716bar), .A2(n715bar), .ZN(n717bar) );
  OR2_X1 U247 ( .A1(n714), .A2(n713), .ZN(n715) );
  AND2_X1 U247bar ( .A1(n714bar), .A2(n713bar), .ZN(n715bar) );
  OR2_X1 U248 ( .A1(in[116]), .A2(in[110]), .ZN(n713) );
  AND2_X1 U248bar ( .A1(inbar[116]), .A2(inbar[110]), .ZN(n713bar) );
  OR2_X1 U249 ( .A1(in[133]), .A2(in[130]), .ZN(n714) );
  AND2_X1 U249bar ( .A1(inbar[133]), .A2(inbar[130]), .ZN(n714bar) );
  OR2_X1 U250 ( .A1(n712), .A2(n711), .ZN(n716) );
  AND2_X1 U250bar ( .A1(n712bar), .A2(n711bar), .ZN(n716bar) );
  OR2_X1 U251 ( .A1(in[203]), .A2(in[135]), .ZN(n711) );
  AND2_X1 U251bar ( .A1(inbar[203]), .A2(inbar[135]), .ZN(n711bar) );
  OR2_X1 U252 ( .A1(in[232]), .A2(in[223]), .ZN(n712) );
  AND2_X1 U252bar ( .A1(inbar[232]), .A2(inbar[223]), .ZN(n712bar) );
  OR2_X1 U253 ( .A1(n710), .A2(n709), .ZN(n718) );
  AND2_X1 U253bar ( .A1(n710bar), .A2(n709bar), .ZN(n718bar) );
  OR2_X1 U254 ( .A1(n708), .A2(n707), .ZN(n709) );
  AND2_X1 U254bar ( .A1(n708bar), .A2(n707bar), .ZN(n709bar) );
  OR2_X1 U255 ( .A1(in[255]), .A2(in[233]), .ZN(n707) );
  AND2_X1 U255bar ( .A1(inbar[255]), .A2(inbar[233]), .ZN(n707bar) );
  OR2_X1 U256 ( .A1(in_53), .A2(in_34), .ZN(n708) );
  AND2_X1 U256bar ( .A1(in_53bar), .A2(in_34bar), .ZN(n708bar) );
  OR2_X1 U257 ( .A1(n706), .A2(n705), .ZN(n710) );
  AND2_X1 U257bar ( .A1(n706bar), .A2(n705bar), .ZN(n710bar) );
  OR2_X1 U258 ( .A1(in_57), .A2(in_55), .ZN(n705) );
  AND2_X1 U258bar ( .A1(in_57bar), .A2(in_55bar), .ZN(n705bar) );
  OR2_X1 U259 ( .A1(in_68), .A2(in_67), .ZN(n706) );
  AND2_X1 U259bar ( .A1(in_68bar), .A2(in_67bar), .ZN(n706bar) );
  OR2_X1 U260 ( .A1(n704), .A2(n703), .ZN(n921) );
  AND2_X1 U260bar ( .A1(n704bar), .A2(n703bar), .ZN(n921bar) );
  OR2_X1 U261 ( .A1(n702), .A2(n701), .ZN(n703) );
  AND2_X1 U261bar ( .A1(n702bar), .A2(n701bar), .ZN(n703bar) );
  OR2_X1 U262 ( .A1(n700), .A2(n699), .ZN(n701) );
  AND2_X1 U262bar ( .A1(n700bar), .A2(n699bar), .ZN(n701bar) );
  OR2_X1 U263 ( .A1(n944), .A2(n872), .ZN(n699) );
  AND2_X1 U263bar ( .A1(n944bar), .A2(n872bar), .ZN(n699bar) );
  OR2_X1 U264 ( .A1(n698), .A2(n697), .ZN(n872) );
  AND2_X1 U264bar ( .A1(n698bar), .A2(n697bar), .ZN(n872bar) );
  OR2_X1 U265 ( .A1(n696), .A2(n695), .ZN(n697) );
  AND2_X1 U265bar ( .A1(n696bar), .A2(n695bar), .ZN(n697bar) );
  OR2_X1 U266 ( .A1(n694), .A2(n693), .ZN(n695) );
  AND2_X1 U266bar ( .A1(n694bar), .A2(n693bar), .ZN(n695bar) );
  OR2_X1 U267 ( .A1(in[121]), .A2(in[102]), .ZN(n693) );
  AND2_X1 U267bar ( .A1(inbar[121]), .A2(inbar[102]), .ZN(n693bar) );
  OR2_X1 U268 ( .A1(in[162]), .A2(in[161]), .ZN(n694) );
  AND2_X1 U268bar ( .A1(inbar[162]), .A2(inbar[161]), .ZN(n694bar) );
  OR2_X1 U269 ( .A1(n692), .A2(n691), .ZN(n696) );
  AND2_X1 U269bar ( .A1(n692bar), .A2(n691bar), .ZN(n696bar) );
  OR2_X1 U270 ( .A1(in[192]), .A2(in[178]), .ZN(n691) );
  AND2_X1 U270bar ( .A1(inbar[192]), .A2(inbar[178]), .ZN(n691bar) );
  OR2_X1 U271 ( .A1(in[244]), .A2(in[209]), .ZN(n692) );
  AND2_X1 U271bar ( .A1(inbar[244]), .A2(inbar[209]), .ZN(n692bar) );
  OR2_X1 U272 ( .A1(n690), .A2(n689), .ZN(n698) );
  AND2_X1 U272bar ( .A1(n690bar), .A2(n689bar), .ZN(n698bar) );
  OR2_X1 U273 ( .A1(n688), .A2(n687), .ZN(n689) );
  AND2_X1 U273bar ( .A1(n688bar), .A2(n687bar), .ZN(n689bar) );
  OR2_X1 U274 ( .A1(in[90]), .A2(in[254]), .ZN(n687) );
  AND2_X1 U274bar ( .A1(inbar[90]), .A2(inbar[254]), .ZN(n687bar) );
  OR2_X1 U275 ( .A1(in_36), .A2(in_32), .ZN(n688) );
  AND2_X1 U275bar ( .A1(in_36bar), .A2(in_32bar), .ZN(n688bar) );
  OR2_X1 U276 ( .A1(n686), .A2(n685), .ZN(n690) );
  AND2_X1 U276bar ( .A1(n686bar), .A2(n685bar), .ZN(n690bar) );
  OR2_X1 U277 ( .A1(in_62), .A2(in_37), .ZN(n685) );
  AND2_X1 U277bar ( .A1(in_62bar), .A2(in_37bar), .ZN(n685bar) );
  OR2_X1 U278 ( .A1(in_75), .A2(in_73), .ZN(n686) );
  AND2_X1 U278bar ( .A1(in_75bar), .A2(in_73bar), .ZN(n686bar) );
  OR2_X1 U279 ( .A1(n684), .A2(n683), .ZN(n944) );
  AND2_X1 U279bar ( .A1(n684bar), .A2(n683bar), .ZN(n944bar) );
  OR2_X1 U280 ( .A1(n682), .A2(n681), .ZN(n683) );
  AND2_X1 U280bar ( .A1(n682bar), .A2(n681bar), .ZN(n683bar) );
  OR2_X1 U281 ( .A1(n680), .A2(n679), .ZN(n681) );
  AND2_X1 U281bar ( .A1(n680bar), .A2(n679bar), .ZN(n681bar) );
  OR2_X1 U282 ( .A1(in[171]), .A2(in[153]), .ZN(n679) );
  AND2_X1 U282bar ( .A1(inbar[171]), .A2(inbar[153]), .ZN(n679bar) );
  OR2_X1 U283 ( .A1(in[187]), .A2(in[176]), .ZN(n680) );
  AND2_X1 U283bar ( .A1(inbar[187]), .A2(inbar[176]), .ZN(n680bar) );
  OR2_X1 U284 ( .A1(n678), .A2(n677), .ZN(n682) );
  AND2_X1 U284bar ( .A1(n678bar), .A2(n677bar), .ZN(n682bar) );
  OR2_X1 U285 ( .A1(in[245]), .A2(in[211]), .ZN(n677) );
  AND2_X1 U285bar ( .A1(inbar[245]), .A2(inbar[211]), .ZN(n677bar) );
  OR2_X1 U286 ( .A1(in[97]), .A2(in[88]), .ZN(n678) );
  AND2_X1 U286bar ( .A1(inbar[97]), .A2(inbar[88]), .ZN(n678bar) );
  OR2_X1 U287 ( .A1(n676), .A2(n675), .ZN(n684) );
  AND2_X1 U287bar ( .A1(n676bar), .A2(n675bar), .ZN(n684bar) );
  OR2_X1 U288 ( .A1(n674), .A2(n673), .ZN(n675) );
  AND2_X1 U288bar ( .A1(n674bar), .A2(n673bar), .ZN(n675bar) );
  OR2_X1 U289 ( .A1(in_10), .A2(in_0), .ZN(n673) );
  AND2_X1 U289bar ( .A1(in_10bar), .A2(in_0bar), .ZN(n673bar) );
  OR2_X1 U290 ( .A1(in_59), .A2(in_5), .ZN(n674) );
  AND2_X1 U290bar ( .A1(in_59bar), .A2(in_5bar), .ZN(n674bar) );
  OR2_X1 U291 ( .A1(n672), .A2(n671), .ZN(n676) );
  AND2_X1 U291bar ( .A1(n672bar), .A2(n671bar), .ZN(n676bar) );
  OR2_X1 U292 ( .A1(in_60), .A2(in_6), .ZN(n671) );
  AND2_X1 U292bar ( .A1(in_60bar), .A2(in_6bar), .ZN(n671bar) );
  OR2_X1 U293 ( .A1(in_77), .A2(in_69), .ZN(n672) );
  AND2_X1 U293bar ( .A1(in_77bar), .A2(in_69bar), .ZN(n672bar) );
  OR2_X1 U294 ( .A1(in[113]), .A2(n864), .ZN(n700) );
  AND2_X1 U294bar ( .A1(inbar[113]), .A2(n864bar), .ZN(n700bar) );
  OR2_X1 U295 ( .A1(n670), .A2(n669), .ZN(n864) );
  AND2_X1 U295bar ( .A1(n670bar), .A2(n669bar), .ZN(n864bar) );
  OR2_X1 U296 ( .A1(n668), .A2(n667), .ZN(n669) );
  AND2_X1 U296bar ( .A1(n668bar), .A2(n667bar), .ZN(n669bar) );
  OR2_X1 U297 ( .A1(n666), .A2(n665), .ZN(n667) );
  AND2_X1 U297bar ( .A1(n666bar), .A2(n665bar), .ZN(n667bar) );
  OR2_X1 U298 ( .A1(in[125]), .A2(in[107]), .ZN(n665) );
  AND2_X1 U298bar ( .A1(inbar[125]), .A2(inbar[107]), .ZN(n665bar) );
  OR2_X1 U299 ( .A1(in[138]), .A2(in[126]), .ZN(n666) );
  AND2_X1 U299bar ( .A1(inbar[138]), .A2(inbar[126]), .ZN(n666bar) );
  OR2_X1 U300 ( .A1(n664), .A2(n663), .ZN(n668) );
  AND2_X1 U300bar ( .A1(n664bar), .A2(n663bar), .ZN(n668bar) );
  OR2_X1 U301 ( .A1(in[189]), .A2(in[143]), .ZN(n663) );
  AND2_X1 U301bar ( .A1(inbar[189]), .A2(inbar[143]), .ZN(n663bar) );
  OR2_X1 U302 ( .A1(in[99]), .A2(in[214]), .ZN(n664) );
  AND2_X1 U302bar ( .A1(inbar[99]), .A2(inbar[214]), .ZN(n664bar) );
  OR2_X1 U303 ( .A1(n662), .A2(n661), .ZN(n670) );
  AND2_X1 U303bar ( .A1(n662bar), .A2(n661bar), .ZN(n670bar) );
  OR2_X1 U304 ( .A1(n660), .A2(n659), .ZN(n661) );
  AND2_X1 U304bar ( .A1(n660bar), .A2(n659bar), .ZN(n661bar) );
  OR2_X1 U305 ( .A1(in_15), .A2(in_12), .ZN(n659) );
  AND2_X1 U305bar ( .A1(in_15bar), .A2(in_12bar), .ZN(n659bar) );
  OR2_X1 U306 ( .A1(in_20), .A2(in_2), .ZN(n660) );
  AND2_X1 U306bar ( .A1(in_20bar), .A2(in_2bar), .ZN(n660bar) );
  OR2_X1 U307 ( .A1(n658), .A2(n657), .ZN(n662) );
  AND2_X1 U307bar ( .A1(n658bar), .A2(n657bar), .ZN(n662bar) );
  OR2_X1 U308 ( .A1(in_30), .A2(in_3), .ZN(n657) );
  AND2_X1 U308bar ( .A1(in_30bar), .A2(in_3bar), .ZN(n657bar) );
  OR2_X1 U309 ( .A1(in_4), .A2(in_38), .ZN(n658) );
  AND2_X1 U309bar ( .A1(in_4bar), .A2(in_38bar), .ZN(n658bar) );
  OR2_X1 U310 ( .A1(n656), .A2(n655), .ZN(n702) );
  AND2_X1 U310bar ( .A1(n656bar), .A2(n655bar), .ZN(n702bar) );
  OR2_X1 U311 ( .A1(in[148]), .A2(in[137]), .ZN(n655) );
  AND2_X1 U311bar ( .A1(inbar[148]), .A2(inbar[137]), .ZN(n655bar) );
  OR2_X1 U312 ( .A1(in[149]), .A2(n654), .ZN(n656) );
  AND2_X1 U312bar ( .A1(inbar[149]), .A2(n654bar), .ZN(n656bar) );
  OR2_X1 U313 ( .A1(in[195]), .A2(in[190]), .ZN(n654) );
  AND2_X1 U313bar ( .A1(inbar[195]), .A2(inbar[190]), .ZN(n654bar) );
  OR2_X1 U314 ( .A1(n653), .A2(n652), .ZN(n704) );
  AND2_X1 U314bar ( .A1(n653bar), .A2(n652bar), .ZN(n704bar) );
  OR2_X1 U315 ( .A1(n651), .A2(n650), .ZN(n652) );
  AND2_X1 U315bar ( .A1(n651bar), .A2(n650bar), .ZN(n652bar) );
  OR2_X1 U316 ( .A1(in[98]), .A2(in[197]), .ZN(n650) );
  AND2_X1 U316bar ( .A1(inbar[98]), .A2(inbar[197]), .ZN(n650bar) );
  OR2_X1 U317 ( .A1(in_11), .A2(n649), .ZN(n651) );
  AND2_X1 U317bar ( .A1(in_11bar), .A2(n649bar), .ZN(n651bar) );
  OR2_X1 U318 ( .A1(in_26), .A2(in_14), .ZN(n649) );
  AND2_X1 U318bar ( .A1(in_26bar), .A2(in_14bar), .ZN(n649bar) );
  OR2_X1 U319 ( .A1(n648), .A2(n647), .ZN(n653) );
  AND2_X1 U319bar ( .A1(n648bar), .A2(n647bar), .ZN(n653bar) );
  OR2_X1 U320 ( .A1(in_35), .A2(in_27), .ZN(n647) );
  AND2_X1 U320bar ( .A1(in_35bar), .A2(in_27bar), .ZN(n647bar) );
  OR2_X1 U321 ( .A1(in_50), .A2(n646), .ZN(n648) );
  AND2_X1 U321bar ( .A1(in_50bar), .A2(n646bar), .ZN(n648bar) );
  OR2_X1 U322 ( .A1(in_78), .A2(in_61), .ZN(n646) );
  AND2_X1 U322bar ( .A1(in_78bar), .A2(in_61bar), .ZN(n646bar) );
  OR2_X1 U323 ( .A1(n942), .A2(n645), .ZN(n720) );
  AND2_X1 U323bar ( .A1(n942bar), .A2(n645bar), .ZN(n720bar) );
  OR2_X1 U324 ( .A1(in[106]), .A2(n863), .ZN(n645) );
  AND2_X1 U324bar ( .A1(inbar[106]), .A2(n863bar), .ZN(n645bar) );
  OR2_X1 U325 ( .A1(n644), .A2(n643), .ZN(n863) );
  AND2_X1 U325bar ( .A1(n644bar), .A2(n643bar), .ZN(n863bar) );
  OR2_X1 U326 ( .A1(n642), .A2(n641), .ZN(n643) );
  AND2_X1 U326bar ( .A1(n642bar), .A2(n641bar), .ZN(n643bar) );
  OR2_X1 U327 ( .A1(n640), .A2(n639), .ZN(n641) );
  AND2_X1 U327bar ( .A1(n640bar), .A2(n639bar), .ZN(n641bar) );
  OR2_X1 U328 ( .A1(in[127]), .A2(in[122]), .ZN(n639) );
  AND2_X1 U328bar ( .A1(inbar[127]), .A2(inbar[122]), .ZN(n639bar) );
  OR2_X1 U329 ( .A1(in[156]), .A2(in[132]), .ZN(n640) );
  AND2_X1 U329bar ( .A1(inbar[156]), .A2(inbar[132]), .ZN(n640bar) );
  OR2_X1 U330 ( .A1(n638), .A2(n637), .ZN(n642) );
  AND2_X1 U330bar ( .A1(n638bar), .A2(n637bar), .ZN(n642bar) );
  OR2_X1 U331 ( .A1(in[159]), .A2(in[157]), .ZN(n637) );
  AND2_X1 U331bar ( .A1(inbar[159]), .A2(inbar[157]), .ZN(n637bar) );
  OR2_X1 U332 ( .A1(in[185]), .A2(in[169]), .ZN(n638) );
  AND2_X1 U332bar ( .A1(inbar[185]), .A2(inbar[169]), .ZN(n638bar) );
  OR2_X1 U333 ( .A1(n636), .A2(n635), .ZN(n644) );
  AND2_X1 U333bar ( .A1(n636bar), .A2(n635bar), .ZN(n644bar) );
  OR2_X1 U334 ( .A1(n634), .A2(n633), .ZN(n635) );
  AND2_X1 U334bar ( .A1(n634bar), .A2(n633bar), .ZN(n635bar) );
  OR2_X1 U335 ( .A1(in[239]), .A2(in[218]), .ZN(n633) );
  AND2_X1 U335bar ( .A1(inbar[239]), .A2(inbar[218]), .ZN(n633bar) );
  OR2_X1 U336 ( .A1(in_13), .A2(in[87]), .ZN(n634) );
  AND2_X1 U336bar ( .A1(in_13bar), .A2(inbar[87]), .ZN(n634bar) );
  OR2_X1 U337 ( .A1(n632), .A2(n631), .ZN(n636) );
  AND2_X1 U337bar ( .A1(n632bar), .A2(n631bar), .ZN(n636bar) );
  OR2_X1 U338 ( .A1(in_72), .A2(in_70), .ZN(n631) );
  AND2_X1 U338bar ( .A1(in_72bar), .A2(in_70bar), .ZN(n631bar) );
  OR2_X1 U339 ( .A1(in_80), .A2(in_74), .ZN(n632) );
  AND2_X1 U339bar ( .A1(in_80bar), .A2(in_74bar), .ZN(n632bar) );
  OR2_X1 U340 ( .A1(n630), .A2(n629), .ZN(n942) );
  AND2_X1 U340bar ( .A1(n630bar), .A2(n629bar), .ZN(n942bar) );
  OR2_X1 U341 ( .A1(n628), .A2(n627), .ZN(n629) );
  AND2_X1 U341bar ( .A1(n628bar), .A2(n627bar), .ZN(n629bar) );
  OR2_X1 U342 ( .A1(n626), .A2(n625), .ZN(n627) );
  AND2_X1 U342bar ( .A1(n626bar), .A2(n625bar), .ZN(n627bar) );
  OR2_X1 U343 ( .A1(in[146]), .A2(in[100]), .ZN(n625) );
  AND2_X1 U343bar ( .A1(inbar[146]), .A2(inbar[100]), .ZN(n625bar) );
  OR2_X1 U344 ( .A1(in[168]), .A2(in[152]), .ZN(n626) );
  AND2_X1 U344bar ( .A1(inbar[168]), .A2(inbar[152]), .ZN(n626bar) );
  OR2_X1 U345 ( .A1(n624), .A2(n623), .ZN(n628) );
  AND2_X1 U345bar ( .A1(n624bar), .A2(n623bar), .ZN(n628bar) );
  OR2_X1 U346 ( .A1(in[199]), .A2(in[182]), .ZN(n623) );
  AND2_X1 U346bar ( .A1(inbar[199]), .A2(inbar[182]), .ZN(n623bar) );
  OR2_X1 U347 ( .A1(in[236]), .A2(in[204]), .ZN(n624) );
  AND2_X1 U347bar ( .A1(inbar[236]), .A2(inbar[204]), .ZN(n624bar) );
  OR2_X1 U348 ( .A1(n622), .A2(n621), .ZN(n630) );
  AND2_X1 U348bar ( .A1(n622bar), .A2(n621bar), .ZN(n630bar) );
  OR2_X1 U349 ( .A1(n620), .A2(n619), .ZN(n621) );
  AND2_X1 U349bar ( .A1(n620bar), .A2(n619bar), .ZN(n621bar) );
  OR2_X1 U350 ( .A1(in[89]), .A2(in[246]), .ZN(n619) );
  AND2_X1 U350bar ( .A1(inbar[89]), .A2(inbar[246]), .ZN(n619bar) );
  OR2_X1 U351 ( .A1(in[95]), .A2(in[92]), .ZN(n620) );
  AND2_X1 U351bar ( .A1(inbar[95]), .A2(inbar[92]), .ZN(n620bar) );
  OR2_X1 U352 ( .A1(n618), .A2(n617), .ZN(n622) );
  AND2_X1 U352bar ( .A1(n618bar), .A2(n617bar), .ZN(n622bar) );
  OR2_X1 U353 ( .A1(in_22), .A2(in_16), .ZN(n617) );
  AND2_X1 U353bar ( .A1(in_22bar), .A2(in_16bar), .ZN(n617bar) );
  OR2_X1 U354 ( .A1(in_51), .A2(in_49), .ZN(n618) );
  AND2_X1 U354bar ( .A1(in_51bar), .A2(in_49bar), .ZN(n618bar) );
  OR2_X1 U355 ( .A1(n616), .A2(n615), .ZN(n722) );
  AND2_X1 U355bar ( .A1(n616bar), .A2(n615bar), .ZN(n722bar) );
  OR2_X1 U356 ( .A1(in[158]), .A2(in[115]), .ZN(n615) );
  AND2_X1 U356bar ( .A1(inbar[158]), .A2(inbar[115]), .ZN(n615bar) );
  OR2_X1 U357 ( .A1(in[163]), .A2(n614), .ZN(n616) );
  AND2_X1 U357bar ( .A1(inbar[163]), .A2(n614bar), .ZN(n616bar) );
  OR2_X1 U358 ( .A1(in[206]), .A2(in[165]), .ZN(n614) );
  AND2_X1 U358bar ( .A1(inbar[206]), .A2(inbar[165]), .ZN(n614bar) );
  OR2_X1 U359 ( .A1(n613), .A2(n612), .ZN(n724) );
  AND2_X1 U359bar ( .A1(n613bar), .A2(n612bar), .ZN(n724bar) );
  OR2_X1 U360 ( .A1(n611), .A2(n610), .ZN(n612) );
  AND2_X1 U360bar ( .A1(n611bar), .A2(n610bar), .ZN(n612bar) );
  OR2_X1 U361 ( .A1(in[213]), .A2(in[207]), .ZN(n610) );
  AND2_X1 U361bar ( .A1(inbar[213]), .A2(inbar[207]), .ZN(n610bar) );
  OR2_X1 U362 ( .A1(in[215]), .A2(n609), .ZN(n611) );
  AND2_X1 U362bar ( .A1(inbar[215]), .A2(n609bar), .ZN(n611bar) );
  OR2_X1 U363 ( .A1(in[230]), .A2(in[220]), .ZN(n609) );
  AND2_X1 U363bar ( .A1(inbar[230]), .A2(inbar[220]), .ZN(n609bar) );
  OR2_X1 U364 ( .A1(n608), .A2(n607), .ZN(n613) );
  AND2_X1 U364bar ( .A1(n608bar), .A2(n607bar), .ZN(n613bar) );
  OR2_X1 U365 ( .A1(in[251]), .A2(in[234]), .ZN(n607) );
  AND2_X1 U365bar ( .A1(inbar[251]), .A2(inbar[234]), .ZN(n607bar) );
  OR2_X1 U366 ( .A1(in_17), .A2(n606), .ZN(n608) );
  AND2_X1 U366bar ( .A1(in_17bar), .A2(n606bar), .ZN(n608bar) );
  OR2_X1 U367 ( .A1(in_65), .A2(in_56), .ZN(n606) );
  AND2_X1 U367bar ( .A1(in_65bar), .A2(in_56bar), .ZN(n606bar) );
  OR2_X1 U368 ( .A1(n605), .A2(n604), .ZN(out[0]) );
  AND2_X1 U368bar ( .A1(n605bar), .A2(n604bar), .ZN(outbar[0]) );
  OR2_X1 U369 ( .A1(n603), .A2(n602), .ZN(n604) );
  AND2_X1 U369bar ( .A1(n603bar), .A2(n602bar), .ZN(n604bar) );
  OR2_X1 U370 ( .A1(n601), .A2(n600), .ZN(n602) );
  AND2_X1 U370bar ( .A1(n601bar), .A2(n600bar), .ZN(n602bar) );
  OR2_X1 U371 ( .A1(n820), .A2(n785), .ZN(n600) );
  AND2_X1 U371bar ( .A1(n820bar), .A2(n785bar), .ZN(n600bar) );
  OR2_X1 U372 ( .A1(n599), .A2(n598), .ZN(n785) );
  AND2_X1 U372bar ( .A1(n599bar), .A2(n598bar), .ZN(n785bar) );
  OR2_X1 U373 ( .A1(n597), .A2(n596), .ZN(n598) );
  AND2_X1 U373bar ( .A1(n597bar), .A2(n596bar), .ZN(n598bar) );
  OR2_X1 U374 ( .A1(n595), .A2(n594), .ZN(n596) );
  AND2_X1 U374bar ( .A1(n595bar), .A2(n594bar), .ZN(n596bar) );
  OR2_X1 U375 ( .A1(in[135]), .A2(in[104]), .ZN(n594) );
  AND2_X1 U375bar ( .A1(inbar[135]), .A2(inbar[104]), .ZN(n594bar) );
  OR2_X1 U376 ( .A1(in[188]), .A2(in[178]), .ZN(n595) );
  AND2_X1 U376bar ( .A1(inbar[188]), .A2(inbar[178]), .ZN(n595bar) );
  OR2_X1 U377 ( .A1(n593), .A2(n592), .ZN(n597) );
  AND2_X1 U377bar ( .A1(n593bar), .A2(n592bar), .ZN(n597bar) );
  OR2_X1 U378 ( .A1(in[217]), .A2(in[194]), .ZN(n592) );
  AND2_X1 U378bar ( .A1(inbar[217]), .A2(inbar[194]), .ZN(n592bar) );
  OR2_X1 U379 ( .A1(in[237]), .A2(in[218]), .ZN(n593) );
  AND2_X1 U379bar ( .A1(inbar[237]), .A2(inbar[218]), .ZN(n593bar) );
  OR2_X1 U380 ( .A1(n591), .A2(n590), .ZN(n599) );
  AND2_X1 U380bar ( .A1(n591bar), .A2(n590bar), .ZN(n599bar) );
  OR2_X1 U381 ( .A1(n589), .A2(n588), .ZN(n590) );
  AND2_X1 U381bar ( .A1(n589bar), .A2(n588bar), .ZN(n590bar) );
  OR2_X1 U382 ( .A1(in_2), .A2(in_10), .ZN(n588) );
  AND2_X1 U382bar ( .A1(in_2bar), .A2(in_10bar), .ZN(n588bar) );
  OR2_X1 U383 ( .A1(in_47), .A2(in_22), .ZN(n589) );
  AND2_X1 U383bar ( .A1(in_47bar), .A2(in_22bar), .ZN(n589bar) );
  OR2_X1 U384 ( .A1(n587), .A2(n586), .ZN(n591) );
  AND2_X1 U384bar ( .A1(n587bar), .A2(n586bar), .ZN(n591bar) );
  OR2_X1 U385 ( .A1(in_56), .A2(in_54), .ZN(n586) );
  AND2_X1 U385bar ( .A1(in_56bar), .A2(in_54bar), .ZN(n586bar) );
  OR2_X1 U386 ( .A1(in_63), .A2(in_61), .ZN(n587) );
  AND2_X1 U386bar ( .A1(in_63bar), .A2(in_61bar), .ZN(n587bar) );
  OR2_X1 U387 ( .A1(n585), .A2(n584), .ZN(n820) );
  AND2_X1 U387bar ( .A1(n585bar), .A2(n584bar), .ZN(n820bar) );
  OR2_X1 U388 ( .A1(n583), .A2(n582), .ZN(n584) );
  AND2_X1 U388bar ( .A1(n583bar), .A2(n582bar), .ZN(n584bar) );
  OR2_X1 U389 ( .A1(n581), .A2(n580), .ZN(n582) );
  AND2_X1 U389bar ( .A1(n581bar), .A2(n580bar), .ZN(n582bar) );
  OR2_X1 U390 ( .A1(in[158]), .A2(in[142]), .ZN(n580) );
  AND2_X1 U390bar ( .A1(inbar[158]), .A2(inbar[142]), .ZN(n580bar) );
  OR2_X1 U391 ( .A1(in[175]), .A2(in[164]), .ZN(n581) );
  AND2_X1 U391bar ( .A1(inbar[175]), .A2(inbar[164]), .ZN(n581bar) );
  OR2_X1 U392 ( .A1(n579), .A2(n578), .ZN(n583) );
  AND2_X1 U392bar ( .A1(n579bar), .A2(n578bar), .ZN(n583bar) );
  OR2_X1 U393 ( .A1(in[228]), .A2(in[204]), .ZN(n578) );
  AND2_X1 U393bar ( .A1(inbar[228]), .A2(inbar[204]), .ZN(n578bar) );
  OR2_X1 U394 ( .A1(in[91]), .A2(in[87]), .ZN(n579) );
  AND2_X1 U394bar ( .A1(inbar[91]), .A2(inbar[87]), .ZN(n579bar) );
  OR2_X1 U395 ( .A1(n577), .A2(n576), .ZN(n585) );
  AND2_X1 U395bar ( .A1(n577bar), .A2(n576bar), .ZN(n585bar) );
  OR2_X1 U396 ( .A1(n575), .A2(n574), .ZN(n576) );
  AND2_X1 U396bar ( .A1(n575bar), .A2(n574bar), .ZN(n576bar) );
  OR2_X1 U397 ( .A1(in_21), .A2(in_11), .ZN(n574) );
  AND2_X1 U397bar ( .A1(in_21bar), .A2(in_11bar), .ZN(n574bar) );
  OR2_X1 U398 ( .A1(in_5), .A2(in_3), .ZN(n575) );
  AND2_X1 U398bar ( .A1(in_5bar), .A2(in_3bar), .ZN(n575bar) );
  OR2_X1 U399 ( .A1(n573), .A2(n572), .ZN(n577) );
  AND2_X1 U399bar ( .A1(n573bar), .A2(n572bar), .ZN(n577bar) );
  OR2_X1 U400 ( .A1(in_68), .A2(in_64), .ZN(n572) );
  AND2_X1 U400bar ( .A1(in_68bar), .A2(in_64bar), .ZN(n572bar) );
  OR2_X1 U401 ( .A1(in_76), .A2(in_73), .ZN(n573) );
  AND2_X1 U401bar ( .A1(in_76bar), .A2(in_73bar), .ZN(n573bar) );
  OR2_X1 U402 ( .A1(n778), .A2(n571), .ZN(n601) );
  AND2_X1 U402bar ( .A1(n778bar), .A2(n571bar), .ZN(n601bar) );
  OR2_X1 U403 ( .A1(in[100]), .A2(n965), .ZN(n571) );
  AND2_X1 U403bar ( .A1(inbar[100]), .A2(n965bar), .ZN(n571bar) );
  OR2_X1 U404 ( .A1(n570), .A2(n569), .ZN(n965) );
  AND2_X1 U404bar ( .A1(n570bar), .A2(n569bar), .ZN(n965bar) );
  OR2_X1 U405 ( .A1(n568), .A2(n567), .ZN(n569) );
  AND2_X1 U405bar ( .A1(n568bar), .A2(n567bar), .ZN(n569bar) );
  OR2_X1 U406 ( .A1(n566), .A2(n565), .ZN(n567) );
  AND2_X1 U406bar ( .A1(n566bar), .A2(n565bar), .ZN(n567bar) );
  OR2_X1 U407 ( .A1(n817), .A2(n750), .ZN(n565) );
  AND2_X1 U407bar ( .A1(n817bar), .A2(n750bar), .ZN(n565bar) );
  OR2_X1 U408 ( .A1(n564), .A2(n563), .ZN(n750) );
  AND2_X1 U408bar ( .A1(n564bar), .A2(n563bar), .ZN(n750bar) );
  OR2_X1 U409 ( .A1(n562), .A2(n561), .ZN(n563) );
  AND2_X1 U409bar ( .A1(n562bar), .A2(n561bar), .ZN(n563bar) );
  OR2_X1 U410 ( .A1(n560), .A2(n559), .ZN(n561) );
  AND2_X1 U410bar ( .A1(n560bar), .A2(n559bar), .ZN(n561bar) );
  OR2_X1 U411 ( .A1(in[119]), .A2(in[103]), .ZN(n559) );
  AND2_X1 U411bar ( .A1(inbar[119]), .A2(inbar[103]), .ZN(n559bar) );
  OR2_X1 U412 ( .A1(in[137]), .A2(in[133]), .ZN(n560) );
  AND2_X1 U412bar ( .A1(inbar[137]), .A2(inbar[133]), .ZN(n560bar) );
  OR2_X1 U413 ( .A1(n558), .A2(n557), .ZN(n562) );
  AND2_X1 U413bar ( .A1(n558bar), .A2(n557bar), .ZN(n562bar) );
  OR2_X1 U414 ( .A1(in[176]), .A2(in[173]), .ZN(n557) );
  AND2_X1 U414bar ( .A1(inbar[176]), .A2(inbar[173]), .ZN(n557bar) );
  OR2_X1 U415 ( .A1(in[210]), .A2(in[181]), .ZN(n558) );
  AND2_X1 U415bar ( .A1(inbar[210]), .A2(inbar[181]), .ZN(n558bar) );
  OR2_X1 U416 ( .A1(n556), .A2(n555), .ZN(n564) );
  AND2_X1 U416bar ( .A1(n556bar), .A2(n555bar), .ZN(n564bar) );
  OR2_X1 U417 ( .A1(n554), .A2(n553), .ZN(n555) );
  AND2_X1 U417bar ( .A1(n554bar), .A2(n553bar), .ZN(n555bar) );
  OR2_X1 U418 ( .A1(in_13), .A2(in[234]), .ZN(n553) );
  AND2_X1 U418bar ( .A1(in_13bar), .A2(inbar[234]), .ZN(n553bar) );
  OR2_X1 U419 ( .A1(in_38), .A2(in_32), .ZN(n554) );
  AND2_X1 U419bar ( .A1(in_38bar), .A2(in_32bar), .ZN(n554bar) );
  OR2_X1 U420 ( .A1(n552), .A2(n551), .ZN(n556) );
  AND2_X1 U420bar ( .A1(n552bar), .A2(n551bar), .ZN(n556bar) );
  OR2_X1 U421 ( .A1(in_42), .A2(in_41), .ZN(n551) );
  AND2_X1 U421bar ( .A1(in_42bar), .A2(in_41bar), .ZN(n551bar) );
  OR2_X1 U422 ( .A1(in_7), .A2(in_49), .ZN(n552) );
  AND2_X1 U422bar ( .A1(in_7bar), .A2(in_49bar), .ZN(n552bar) );
  OR2_X1 U423 ( .A1(n550), .A2(n549), .ZN(n817) );
  AND2_X1 U423bar ( .A1(n550bar), .A2(n549bar), .ZN(n817bar) );
  OR2_X1 U424 ( .A1(n548), .A2(n547), .ZN(n549) );
  AND2_X1 U424bar ( .A1(n548bar), .A2(n547bar), .ZN(n549bar) );
  OR2_X1 U425 ( .A1(n546), .A2(n545), .ZN(n547) );
  AND2_X1 U425bar ( .A1(n546bar), .A2(n545bar), .ZN(n547bar) );
  OR2_X1 U426 ( .A1(in[159]), .A2(in[105]), .ZN(n545) );
  AND2_X1 U426bar ( .A1(inbar[159]), .A2(inbar[105]), .ZN(n545bar) );
  OR2_X1 U427 ( .A1(in[206]), .A2(in[183]), .ZN(n546) );
  AND2_X1 U427bar ( .A1(inbar[206]), .A2(inbar[183]), .ZN(n546bar) );
  OR2_X1 U428 ( .A1(n544), .A2(n543), .ZN(n548) );
  AND2_X1 U428bar ( .A1(n544bar), .A2(n543bar), .ZN(n548bar) );
  OR2_X1 U429 ( .A1(in[229]), .A2(in[219]), .ZN(n543) );
  AND2_X1 U429bar ( .A1(inbar[229]), .A2(inbar[219]), .ZN(n543bar) );
  OR2_X1 U430 ( .A1(in[235]), .A2(in[232]), .ZN(n544) );
  AND2_X1 U430bar ( .A1(inbar[235]), .A2(inbar[232]), .ZN(n544bar) );
  OR2_X1 U431 ( .A1(n542), .A2(n541), .ZN(n550) );
  AND2_X1 U431bar ( .A1(n542bar), .A2(n541bar), .ZN(n550bar) );
  OR2_X1 U432 ( .A1(n540), .A2(n539), .ZN(n541) );
  AND2_X1 U432bar ( .A1(n540bar), .A2(n539bar), .ZN(n541bar) );
  OR2_X1 U433 ( .A1(in[249]), .A2(in[242]), .ZN(n539) );
  AND2_X1 U433bar ( .A1(inbar[249]), .A2(inbar[242]), .ZN(n539bar) );
  OR2_X1 U434 ( .A1(in[89]), .A2(in[254]), .ZN(n540) );
  AND2_X1 U434bar ( .A1(inbar[89]), .A2(inbar[254]), .ZN(n540bar) );
  OR2_X1 U435 ( .A1(n538), .A2(n537), .ZN(n542) );
  AND2_X1 U435bar ( .A1(n538bar), .A2(n537bar), .ZN(n542bar) );
  OR2_X1 U436 ( .A1(in_14), .A2(in[99]), .ZN(n537) );
  AND2_X1 U436bar ( .A1(in_14bar), .A2(inbar[99]), .ZN(n537bar) );
  OR2_X1 U437 ( .A1(in_60), .A2(in_18), .ZN(n538) );
  AND2_X1 U437bar ( .A1(in_60bar), .A2(in_18bar), .ZN(n538bar) );
  OR2_X1 U438 ( .A1(in[113]), .A2(n763), .ZN(n566) );
  AND2_X1 U438bar ( .A1(inbar[113]), .A2(n763bar), .ZN(n566bar) );
  OR2_X1 U439 ( .A1(n536), .A2(n535), .ZN(n763) );
  AND2_X1 U439bar ( .A1(n536bar), .A2(n535bar), .ZN(n763bar) );
  OR2_X1 U440 ( .A1(n534), .A2(n533), .ZN(n535) );
  AND2_X1 U440bar ( .A1(n534bar), .A2(n533bar), .ZN(n535bar) );
  OR2_X1 U441 ( .A1(n532), .A2(n531), .ZN(n533) );
  AND2_X1 U441bar ( .A1(n532bar), .A2(n531bar), .ZN(n533bar) );
  OR2_X1 U442 ( .A1(in[115]), .A2(in[110]), .ZN(n531) );
  AND2_X1 U442bar ( .A1(inbar[115]), .A2(inbar[110]), .ZN(n531bar) );
  OR2_X1 U443 ( .A1(in[125]), .A2(in[117]), .ZN(n532) );
  AND2_X1 U443bar ( .A1(inbar[125]), .A2(inbar[117]), .ZN(n532bar) );
  OR2_X1 U444 ( .A1(n530), .A2(n529), .ZN(n534) );
  AND2_X1 U444bar ( .A1(n530bar), .A2(n529bar), .ZN(n534bar) );
  OR2_X1 U445 ( .A1(in[180]), .A2(in[128]), .ZN(n529) );
  AND2_X1 U445bar ( .A1(inbar[180]), .A2(inbar[128]), .ZN(n529bar) );
  OR2_X1 U446 ( .A1(in[205]), .A2(in[201]), .ZN(n530) );
  AND2_X1 U446bar ( .A1(inbar[205]), .A2(inbar[201]), .ZN(n530bar) );
  OR2_X1 U447 ( .A1(n528), .A2(n527), .ZN(n536) );
  AND2_X1 U447bar ( .A1(n528bar), .A2(n527bar), .ZN(n536bar) );
  OR2_X1 U448 ( .A1(n526), .A2(n525), .ZN(n527) );
  AND2_X1 U448bar ( .A1(n526bar), .A2(n525bar), .ZN(n527bar) );
  OR2_X1 U449 ( .A1(in[244]), .A2(in[239]), .ZN(n525) );
  AND2_X1 U449bar ( .A1(inbar[244]), .A2(inbar[239]), .ZN(n525bar) );
  OR2_X1 U450 ( .A1(in[95]), .A2(in[83]), .ZN(n526) );
  AND2_X1 U450bar ( .A1(inbar[95]), .A2(inbar[83]), .ZN(n526bar) );
  OR2_X1 U451 ( .A1(n524), .A2(n523), .ZN(n528) );
  AND2_X1 U451bar ( .A1(n524bar), .A2(n523bar), .ZN(n528bar) );
  OR2_X1 U452 ( .A1(in_24), .A2(in[97]), .ZN(n523) );
  AND2_X1 U452bar ( .A1(in_24bar), .A2(inbar[97]), .ZN(n523bar) );
  OR2_X1 U453 ( .A1(in_33), .A2(in_27), .ZN(n524) );
  AND2_X1 U453bar ( .A1(in_33bar), .A2(in_27bar), .ZN(n524bar) );
  OR2_X1 U454 ( .A1(n522), .A2(n521), .ZN(n568) );
  AND2_X1 U454bar ( .A1(n522bar), .A2(n521bar), .ZN(n568bar) );
  OR2_X1 U455 ( .A1(in[145]), .A2(in[126]), .ZN(n521) );
  AND2_X1 U455bar ( .A1(inbar[145]), .A2(inbar[126]), .ZN(n521bar) );
  OR2_X1 U456 ( .A1(in[169]), .A2(n520), .ZN(n522) );
  AND2_X1 U456bar ( .A1(inbar[169]), .A2(n520bar), .ZN(n522bar) );
  OR2_X1 U457 ( .A1(in[221]), .A2(in[172]), .ZN(n520) );
  AND2_X1 U457bar ( .A1(inbar[221]), .A2(inbar[172]), .ZN(n520bar) );
  OR2_X1 U458 ( .A1(n519), .A2(n518), .ZN(n570) );
  AND2_X1 U458bar ( .A1(n519bar), .A2(n518bar), .ZN(n570bar) );
  OR2_X1 U459 ( .A1(n517), .A2(n516), .ZN(n518) );
  AND2_X1 U459bar ( .A1(n517bar), .A2(n516bar), .ZN(n518bar) );
  OR2_X1 U460 ( .A1(in[241]), .A2(in[224]), .ZN(n516) );
  AND2_X1 U460bar ( .A1(inbar[241]), .A2(inbar[224]), .ZN(n516bar) );
  OR2_X1 U461 ( .A1(in[86]), .A2(n515), .ZN(n517) );
  AND2_X1 U461bar ( .A1(inbar[86]), .A2(n515bar), .ZN(n517bar) );
  OR2_X1 U462 ( .A1(in_43), .A2(in_34), .ZN(n515) );
  AND2_X1 U462bar ( .A1(in_43bar), .A2(in_34bar), .ZN(n515bar) );
  OR2_X1 U463 ( .A1(n514), .A2(n513), .ZN(n519) );
  AND2_X1 U463bar ( .A1(n514bar), .A2(n513bar), .ZN(n519bar) );
  OR2_X1 U464 ( .A1(in_65), .A2(in_51), .ZN(n513) );
  AND2_X1 U464bar ( .A1(in_65bar), .A2(in_51bar), .ZN(n513bar) );
  OR2_X1 U465 ( .A1(in_75), .A2(n512), .ZN(n514) );
  AND2_X1 U465bar ( .A1(in_75bar), .A2(n512bar), .ZN(n514bar) );
  OR2_X1 U466 ( .A1(in_81), .A2(in_77), .ZN(n512) );
  AND2_X1 U466bar ( .A1(in_81bar), .A2(in_77bar), .ZN(n512bar) );
  OR2_X1 U467 ( .A1(n511), .A2(n510), .ZN(n778) );
  AND2_X1 U467bar ( .A1(n511bar), .A2(n510bar), .ZN(n778bar) );
  OR2_X1 U468 ( .A1(n509), .A2(n508), .ZN(n510) );
  AND2_X1 U468bar ( .A1(n509bar), .A2(n508bar), .ZN(n510bar) );
  OR2_X1 U469 ( .A1(n507), .A2(n506), .ZN(n508) );
  AND2_X1 U469bar ( .A1(n507bar), .A2(n506bar), .ZN(n508bar) );
  OR2_X1 U470 ( .A1(in[107]), .A2(in[101]), .ZN(n506) );
  AND2_X1 U470bar ( .A1(inbar[107]), .A2(inbar[101]), .ZN(n506bar) );
  OR2_X1 U471 ( .A1(in[139]), .A2(in[132]), .ZN(n507) );
  AND2_X1 U471bar ( .A1(inbar[139]), .A2(inbar[132]), .ZN(n507bar) );
  OR2_X1 U472 ( .A1(n505), .A2(n504), .ZN(n509) );
  AND2_X1 U472bar ( .A1(n505bar), .A2(n504bar), .ZN(n509bar) );
  OR2_X1 U473 ( .A1(in[146]), .A2(in[141]), .ZN(n504) );
  AND2_X1 U473bar ( .A1(inbar[146]), .A2(inbar[141]), .ZN(n504bar) );
  OR2_X1 U474 ( .A1(in[203]), .A2(in[179]), .ZN(n505) );
  AND2_X1 U474bar ( .A1(inbar[203]), .A2(inbar[179]), .ZN(n505bar) );
  OR2_X1 U475 ( .A1(n503), .A2(n502), .ZN(n511) );
  AND2_X1 U475bar ( .A1(n503bar), .A2(n502bar), .ZN(n511bar) );
  OR2_X1 U476 ( .A1(n501), .A2(n500), .ZN(n502) );
  AND2_X1 U476bar ( .A1(n501bar), .A2(n500bar), .ZN(n502bar) );
  OR2_X1 U477 ( .A1(in[243]), .A2(in[222]), .ZN(n500) );
  AND2_X1 U477bar ( .A1(inbar[243]), .A2(inbar[222]), .ZN(n500bar) );
  OR2_X1 U478 ( .A1(in[251]), .A2(in[250]), .ZN(n501) );
  AND2_X1 U478bar ( .A1(inbar[251]), .A2(inbar[250]), .ZN(n501bar) );
  OR2_X1 U479 ( .A1(n499), .A2(n498), .ZN(n503) );
  AND2_X1 U479bar ( .A1(n499bar), .A2(n498bar), .ZN(n503bar) );
  OR2_X1 U480 ( .A1(in_37), .A2(in_19), .ZN(n498) );
  AND2_X1 U480bar ( .A1(in_37bar), .A2(in_19bar), .ZN(n498bar) );
  OR2_X1 U481 ( .A1(in_78), .A2(in_6), .ZN(n499) );
  AND2_X1 U481bar ( .A1(in_78bar), .A2(in_6bar), .ZN(n499bar) );
  OR2_X1 U482 ( .A1(n497), .A2(n496), .ZN(n603) );
  AND2_X1 U482bar ( .A1(n497bar), .A2(n496bar), .ZN(n603bar) );
  OR2_X1 U483 ( .A1(in[112]), .A2(in[102]), .ZN(n496) );
  AND2_X1 U483bar ( .A1(inbar[112]), .A2(inbar[102]), .ZN(n496bar) );
  OR2_X1 U484 ( .A1(in[123]), .A2(n495), .ZN(n497) );
  AND2_X1 U484bar ( .A1(inbar[123]), .A2(n495bar), .ZN(n497bar) );
  OR2_X1 U485 ( .A1(in[143]), .A2(in[130]), .ZN(n495) );
  AND2_X1 U485bar ( .A1(inbar[143]), .A2(inbar[130]), .ZN(n495bar) );
  OR2_X1 U486 ( .A1(n494), .A2(n493), .ZN(n605) );
  AND2_X1 U486bar ( .A1(n494bar), .A2(n493bar), .ZN(n605bar) );
  OR2_X1 U487 ( .A1(n492), .A2(n491), .ZN(n493) );
  AND2_X1 U487bar ( .A1(n492bar), .A2(n491bar), .ZN(n493bar) );
  OR2_X1 U488 ( .A1(in[216]), .A2(in[213]), .ZN(n491) );
  AND2_X1 U488bar ( .A1(inbar[216]), .A2(inbar[213]), .ZN(n491bar) );
  OR2_X1 U489 ( .A1(in[227]), .A2(n490), .ZN(n492) );
  AND2_X1 U489bar ( .A1(inbar[227]), .A2(n490bar), .ZN(n492bar) );
  OR2_X1 U490 ( .A1(in_0), .A2(in[248]), .ZN(n490) );
  AND2_X1 U490bar ( .A1(in_0bar), .A2(inbar[248]), .ZN(n490bar) );
  OR2_X1 U491 ( .A1(n489), .A2(n488), .ZN(n494) );
  AND2_X1 U491bar ( .A1(n489bar), .A2(n488bar), .ZN(n494bar) );
  OR2_X1 U492 ( .A1(in_46), .A2(in_44), .ZN(n488) );
  AND2_X1 U492bar ( .A1(in_46bar), .A2(in_44bar), .ZN(n488bar) );
  OR2_X1 U493 ( .A1(in_50), .A2(n487), .ZN(n489) );
  AND2_X1 U493bar ( .A1(in_50bar), .A2(n487bar), .ZN(n489bar) );
  OR2_X1 U494 ( .A1(in_9), .A2(in_80), .ZN(n487) );
  AND2_X1 U494bar ( .A1(in_9bar), .A2(in_80bar), .ZN(n487bar) );
endmodule

module sBox_7 ( in, inbar, out, outbar );

  input wire [7:0] in;
  input wire [7:0] inbar;
//input_done

  output wire [7:0] out;
  output wire [7:0] outbar;
//output_done

  wire [255:0] decodeOut;
  wire [255:0] decodeOutbar;
//wire_done

  decode_7 dec ( .in(in), .inbar(inbar), .out(decodeOut), .outbar(decodeOutbar) );
  encode_7 enc ( .in(decodeOut), .inbar(decodeOutbar), .out(out), .outbar(outbar) );
endmodule

module CD2_29 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD2_30 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD2_31 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD2_32 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD4_15 ( a, abar, b, bbar, y, ybar );

  input wire [3:0] a;
  input wire [3:0] b;
  input wire [3:0] abar;
  input wire [3:0] bbar;
//input_done

  output wire [15:0] y;
  output wire [15:0] ybar;
//output_done

//wire_done

  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]) );
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]) );
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]) );
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]) );
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]) );
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]) );
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]) );
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]) );
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]) );
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]) );
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]) );
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]) );
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]) );
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]) );
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]) );
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]) );
endmodule

module CD4_16 ( a, abar, b, bbar, y, ybar );

  input wire [3:0] a;
  input wire [3:0] b;
  input wire [3:0] abar;
  input wire [3:0] bbar;
//input_done

  output wire [15:0] y;
  output wire [15:0] ybar;
//output_done

//wire_done

  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]) );
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]) );
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]) );
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]) );
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]) );
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]) );
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]) );
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]) );
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]) );
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]) );
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]) );
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]) );
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]) );
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]) );
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]) );
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]) );
endmodule

module CD16_8 ( a, abar, b, bbar, y, ybar );

  input wire [15:0] a;
  input wire [15:0] b;
  input wire [15:0] abar;
  input wire [15:0] bbar;
//input_done

  output wire [255:0] y;
  output wire [255:0] ybar;
//output_done

//wire_done

  AND2_X1 U1 ( .A1(b[9]), .A2(a[0]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[9]), .A2(abar[0]), .ZN(ybar[9]) );
  AND2_X1 U2 ( .A1(b[3]), .A2(a[6]), .ZN(y[99]) );
  OR2_X1 U2bar ( .A1(bbar[3]), .A2(abar[6]), .ZN(ybar[99]) );
  AND2_X1 U3 ( .A1(b[2]), .A2(a[6]), .ZN(y[98]) );
  OR2_X1 U3bar ( .A1(bbar[2]), .A2(abar[6]), .ZN(ybar[98]) );
  AND2_X1 U4 ( .A1(b[1]), .A2(a[6]), .ZN(y[97]) );
  OR2_X1 U4bar ( .A1(bbar[1]), .A2(abar[6]), .ZN(ybar[97]) );
  AND2_X1 U5 ( .A1(b[0]), .A2(a[6]), .ZN(y[96]) );
  OR2_X1 U5bar ( .A1(bbar[0]), .A2(abar[6]), .ZN(ybar[96]) );
  AND2_X1 U6 ( .A1(b[15]), .A2(a[5]), .ZN(y[95]) );
  OR2_X1 U6bar ( .A1(bbar[15]), .A2(abar[5]), .ZN(ybar[95]) );
  AND2_X1 U7 ( .A1(b[14]), .A2(a[5]), .ZN(y[94]) );
  OR2_X1 U7bar ( .A1(bbar[14]), .A2(abar[5]), .ZN(ybar[94]) );
  AND2_X1 U8 ( .A1(b[13]), .A2(a[5]), .ZN(y[93]) );
  OR2_X1 U8bar ( .A1(bbar[13]), .A2(abar[5]), .ZN(ybar[93]) );
  AND2_X1 U9 ( .A1(b[12]), .A2(a[5]), .ZN(y[92]) );
  OR2_X1 U9bar ( .A1(bbar[12]), .A2(abar[5]), .ZN(ybar[92]) );
  AND2_X1 U10 ( .A1(b[11]), .A2(a[5]), .ZN(y[91]) );
  OR2_X1 U10bar ( .A1(bbar[11]), .A2(abar[5]), .ZN(ybar[91]) );
  AND2_X1 U11 ( .A1(b[10]), .A2(a[5]), .ZN(y[90]) );
  OR2_X1 U11bar ( .A1(bbar[10]), .A2(abar[5]), .ZN(ybar[90]) );
  AND2_X1 U12 ( .A1(b[8]), .A2(a[0]), .ZN(y[8]) );
  OR2_X1 U12bar ( .A1(bbar[8]), .A2(abar[0]), .ZN(ybar[8]) );
  AND2_X1 U13 ( .A1(a[5]), .A2(b[9]), .ZN(y[89]) );
  OR2_X1 U13bar ( .A1(abar[5]), .A2(bbar[9]), .ZN(ybar[89]) );
  AND2_X1 U14 ( .A1(b[8]), .A2(a[5]), .ZN(y[88]) );
  OR2_X1 U14bar ( .A1(bbar[8]), .A2(abar[5]), .ZN(ybar[88]) );
  AND2_X1 U15 ( .A1(b[7]), .A2(a[5]), .ZN(y[87]) );
  OR2_X1 U15bar ( .A1(bbar[7]), .A2(abar[5]), .ZN(ybar[87]) );
  AND2_X1 U16 ( .A1(b[6]), .A2(a[5]), .ZN(y[86]) );
  OR2_X1 U16bar ( .A1(bbar[6]), .A2(abar[5]), .ZN(ybar[86]) );
  AND2_X1 U17 ( .A1(b[5]), .A2(a[5]), .ZN(y[85]) );
  OR2_X1 U17bar ( .A1(bbar[5]), .A2(abar[5]), .ZN(ybar[85]) );
  AND2_X1 U18 ( .A1(b[4]), .A2(a[5]), .ZN(y[84]) );
  OR2_X1 U18bar ( .A1(bbar[4]), .A2(abar[5]), .ZN(ybar[84]) );
  AND2_X1 U19 ( .A1(a[5]), .A2(b[3]), .ZN(y[83]) );
  OR2_X1 U19bar ( .A1(abar[5]), .A2(bbar[3]), .ZN(ybar[83]) );
  AND2_X1 U20 ( .A1(a[5]), .A2(b[2]), .ZN(y[82]) );
  OR2_X1 U20bar ( .A1(abar[5]), .A2(bbar[2]), .ZN(ybar[82]) );
  AND2_X1 U21 ( .A1(a[5]), .A2(b[1]), .ZN(y[81]) );
  OR2_X1 U21bar ( .A1(abar[5]), .A2(bbar[1]), .ZN(ybar[81]) );
  AND2_X1 U22 ( .A1(a[5]), .A2(b[0]), .ZN(y[80]) );
  OR2_X1 U22bar ( .A1(abar[5]), .A2(bbar[0]), .ZN(ybar[80]) );
  AND2_X1 U23 ( .A1(b[7]), .A2(a[0]), .ZN(y[7]) );
  OR2_X1 U23bar ( .A1(bbar[7]), .A2(abar[0]), .ZN(ybar[7]) );
  AND2_X1 U24 ( .A1(a[4]), .A2(b[15]), .ZN(y[79]) );
  OR2_X1 U24bar ( .A1(abar[4]), .A2(bbar[15]), .ZN(ybar[79]) );
  AND2_X1 U25 ( .A1(a[4]), .A2(b[14]), .ZN(y[78]) );
  OR2_X1 U25bar ( .A1(abar[4]), .A2(bbar[14]), .ZN(ybar[78]) );
  AND2_X1 U26 ( .A1(a[4]), .A2(b[13]), .ZN(y[77]) );
  OR2_X1 U26bar ( .A1(abar[4]), .A2(bbar[13]), .ZN(ybar[77]) );
  AND2_X1 U27 ( .A1(a[4]), .A2(b[12]), .ZN(y[76]) );
  OR2_X1 U27bar ( .A1(abar[4]), .A2(bbar[12]), .ZN(ybar[76]) );
  AND2_X1 U28 ( .A1(a[4]), .A2(b[11]), .ZN(y[75]) );
  OR2_X1 U28bar ( .A1(abar[4]), .A2(bbar[11]), .ZN(ybar[75]) );
  AND2_X1 U29 ( .A1(a[4]), .A2(b[10]), .ZN(y[74]) );
  OR2_X1 U29bar ( .A1(abar[4]), .A2(bbar[10]), .ZN(ybar[74]) );
  AND2_X1 U30 ( .A1(a[4]), .A2(b[9]), .ZN(y[73]) );
  OR2_X1 U30bar ( .A1(abar[4]), .A2(bbar[9]), .ZN(ybar[73]) );
  AND2_X1 U31 ( .A1(a[4]), .A2(b[8]), .ZN(y[72]) );
  OR2_X1 U31bar ( .A1(abar[4]), .A2(bbar[8]), .ZN(ybar[72]) );
  AND2_X1 U32 ( .A1(a[4]), .A2(b[7]), .ZN(y[71]) );
  OR2_X1 U32bar ( .A1(abar[4]), .A2(bbar[7]), .ZN(ybar[71]) );
  AND2_X1 U33 ( .A1(a[4]), .A2(b[6]), .ZN(y[70]) );
  OR2_X1 U33bar ( .A1(abar[4]), .A2(bbar[6]), .ZN(ybar[70]) );
  AND2_X1 U34 ( .A1(b[6]), .A2(a[0]), .ZN(y[6]) );
  OR2_X1 U34bar ( .A1(bbar[6]), .A2(abar[0]), .ZN(ybar[6]) );
  AND2_X1 U35 ( .A1(a[4]), .A2(b[5]), .ZN(y[69]) );
  OR2_X1 U35bar ( .A1(abar[4]), .A2(bbar[5]), .ZN(ybar[69]) );
  AND2_X1 U36 ( .A1(a[4]), .A2(b[4]), .ZN(y[68]) );
  OR2_X1 U36bar ( .A1(abar[4]), .A2(bbar[4]), .ZN(ybar[68]) );
  AND2_X1 U37 ( .A1(a[4]), .A2(b[3]), .ZN(y[67]) );
  OR2_X1 U37bar ( .A1(abar[4]), .A2(bbar[3]), .ZN(ybar[67]) );
  AND2_X1 U38 ( .A1(a[4]), .A2(b[2]), .ZN(y[66]) );
  OR2_X1 U38bar ( .A1(abar[4]), .A2(bbar[2]), .ZN(ybar[66]) );
  AND2_X1 U39 ( .A1(a[4]), .A2(b[1]), .ZN(y[65]) );
  OR2_X1 U39bar ( .A1(abar[4]), .A2(bbar[1]), .ZN(ybar[65]) );
  AND2_X1 U40 ( .A1(a[4]), .A2(b[0]), .ZN(y[64]) );
  OR2_X1 U40bar ( .A1(abar[4]), .A2(bbar[0]), .ZN(ybar[64]) );
  AND2_X1 U41 ( .A1(a[3]), .A2(b[15]), .ZN(y[63]) );
  OR2_X1 U41bar ( .A1(abar[3]), .A2(bbar[15]), .ZN(ybar[63]) );
  AND2_X1 U42 ( .A1(a[3]), .A2(b[14]), .ZN(y[62]) );
  OR2_X1 U42bar ( .A1(abar[3]), .A2(bbar[14]), .ZN(ybar[62]) );
  AND2_X1 U43 ( .A1(a[3]), .A2(b[13]), .ZN(y[61]) );
  OR2_X1 U43bar ( .A1(abar[3]), .A2(bbar[13]), .ZN(ybar[61]) );
  AND2_X1 U44 ( .A1(a[3]), .A2(b[12]), .ZN(y[60]) );
  OR2_X1 U44bar ( .A1(abar[3]), .A2(bbar[12]), .ZN(ybar[60]) );
  AND2_X1 U45 ( .A1(b[5]), .A2(a[0]), .ZN(y[5]) );
  OR2_X1 U45bar ( .A1(bbar[5]), .A2(abar[0]), .ZN(ybar[5]) );
  AND2_X1 U46 ( .A1(a[3]), .A2(b[11]), .ZN(y[59]) );
  OR2_X1 U46bar ( .A1(abar[3]), .A2(bbar[11]), .ZN(ybar[59]) );
  AND2_X1 U47 ( .A1(a[3]), .A2(b[10]), .ZN(y[58]) );
  OR2_X1 U47bar ( .A1(abar[3]), .A2(bbar[10]), .ZN(ybar[58]) );
  AND2_X1 U48 ( .A1(a[3]), .A2(b[9]), .ZN(y[57]) );
  OR2_X1 U48bar ( .A1(abar[3]), .A2(bbar[9]), .ZN(ybar[57]) );
  AND2_X1 U49 ( .A1(a[3]), .A2(b[8]), .ZN(y[56]) );
  OR2_X1 U49bar ( .A1(abar[3]), .A2(bbar[8]), .ZN(ybar[56]) );
  AND2_X1 U50 ( .A1(a[3]), .A2(b[7]), .ZN(y[55]) );
  OR2_X1 U50bar ( .A1(abar[3]), .A2(bbar[7]), .ZN(ybar[55]) );
  AND2_X1 U51 ( .A1(a[3]), .A2(b[6]), .ZN(y[54]) );
  OR2_X1 U51bar ( .A1(abar[3]), .A2(bbar[6]), .ZN(ybar[54]) );
  AND2_X1 U52 ( .A1(a[3]), .A2(b[5]), .ZN(y[53]) );
  OR2_X1 U52bar ( .A1(abar[3]), .A2(bbar[5]), .ZN(ybar[53]) );
  AND2_X1 U53 ( .A1(a[3]), .A2(b[4]), .ZN(y[52]) );
  OR2_X1 U53bar ( .A1(abar[3]), .A2(bbar[4]), .ZN(ybar[52]) );
  AND2_X1 U54 ( .A1(a[3]), .A2(b[3]), .ZN(y[51]) );
  OR2_X1 U54bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[51]) );
  AND2_X1 U55 ( .A1(a[3]), .A2(b[2]), .ZN(y[50]) );
  OR2_X1 U55bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[50]) );
  AND2_X1 U56 ( .A1(b[4]), .A2(a[0]), .ZN(y[4]) );
  OR2_X1 U56bar ( .A1(bbar[4]), .A2(abar[0]), .ZN(ybar[4]) );
  AND2_X1 U57 ( .A1(a[3]), .A2(b[1]), .ZN(y[49]) );
  OR2_X1 U57bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[49]) );
  AND2_X1 U58 ( .A1(a[3]), .A2(b[0]), .ZN(y[48]) );
  OR2_X1 U58bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[48]) );
  AND2_X1 U59 ( .A1(a[2]), .A2(b[15]), .ZN(y[47]) );
  OR2_X1 U59bar ( .A1(abar[2]), .A2(bbar[15]), .ZN(ybar[47]) );
  AND2_X1 U60 ( .A1(a[2]), .A2(b[14]), .ZN(y[46]) );
  OR2_X1 U60bar ( .A1(abar[2]), .A2(bbar[14]), .ZN(ybar[46]) );
  AND2_X1 U61 ( .A1(a[2]), .A2(b[13]), .ZN(y[45]) );
  OR2_X1 U61bar ( .A1(abar[2]), .A2(bbar[13]), .ZN(ybar[45]) );
  AND2_X1 U62 ( .A1(a[2]), .A2(b[12]), .ZN(y[44]) );
  OR2_X1 U62bar ( .A1(abar[2]), .A2(bbar[12]), .ZN(ybar[44]) );
  AND2_X1 U63 ( .A1(a[2]), .A2(b[11]), .ZN(y[43]) );
  OR2_X1 U63bar ( .A1(abar[2]), .A2(bbar[11]), .ZN(ybar[43]) );
  AND2_X1 U64 ( .A1(a[2]), .A2(b[10]), .ZN(y[42]) );
  OR2_X1 U64bar ( .A1(abar[2]), .A2(bbar[10]), .ZN(ybar[42]) );
  AND2_X1 U65 ( .A1(a[2]), .A2(b[9]), .ZN(y[41]) );
  OR2_X1 U65bar ( .A1(abar[2]), .A2(bbar[9]), .ZN(ybar[41]) );
  AND2_X1 U66 ( .A1(a[2]), .A2(b[8]), .ZN(y[40]) );
  OR2_X1 U66bar ( .A1(abar[2]), .A2(bbar[8]), .ZN(ybar[40]) );
  AND2_X1 U67 ( .A1(b[3]), .A2(a[0]), .ZN(y[3]) );
  OR2_X1 U67bar ( .A1(bbar[3]), .A2(abar[0]), .ZN(ybar[3]) );
  AND2_X1 U68 ( .A1(a[2]), .A2(b[7]), .ZN(y[39]) );
  OR2_X1 U68bar ( .A1(abar[2]), .A2(bbar[7]), .ZN(ybar[39]) );
  AND2_X1 U69 ( .A1(a[2]), .A2(b[6]), .ZN(y[38]) );
  OR2_X1 U69bar ( .A1(abar[2]), .A2(bbar[6]), .ZN(ybar[38]) );
  AND2_X1 U70 ( .A1(a[2]), .A2(b[5]), .ZN(y[37]) );
  OR2_X1 U70bar ( .A1(abar[2]), .A2(bbar[5]), .ZN(ybar[37]) );
  AND2_X1 U71 ( .A1(a[2]), .A2(b[4]), .ZN(y[36]) );
  OR2_X1 U71bar ( .A1(abar[2]), .A2(bbar[4]), .ZN(ybar[36]) );
  AND2_X1 U72 ( .A1(a[2]), .A2(b[3]), .ZN(y[35]) );
  OR2_X1 U72bar ( .A1(abar[2]), .A2(bbar[3]), .ZN(ybar[35]) );
  AND2_X1 U73 ( .A1(a[2]), .A2(b[2]), .ZN(y[34]) );
  OR2_X1 U73bar ( .A1(abar[2]), .A2(bbar[2]), .ZN(ybar[34]) );
  AND2_X1 U74 ( .A1(a[2]), .A2(b[1]), .ZN(y[33]) );
  OR2_X1 U74bar ( .A1(abar[2]), .A2(bbar[1]), .ZN(ybar[33]) );
  AND2_X1 U75 ( .A1(a[2]), .A2(b[0]), .ZN(y[32]) );
  OR2_X1 U75bar ( .A1(abar[2]), .A2(bbar[0]), .ZN(ybar[32]) );
  AND2_X1 U76 ( .A1(a[1]), .A2(b[15]), .ZN(y[31]) );
  OR2_X1 U76bar ( .A1(abar[1]), .A2(bbar[15]), .ZN(ybar[31]) );
  AND2_X1 U77 ( .A1(a[1]), .A2(b[14]), .ZN(y[30]) );
  OR2_X1 U77bar ( .A1(abar[1]), .A2(bbar[14]), .ZN(ybar[30]) );
  AND2_X1 U78 ( .A1(b[2]), .A2(a[0]), .ZN(y[2]) );
  OR2_X1 U78bar ( .A1(bbar[2]), .A2(abar[0]), .ZN(ybar[2]) );
  AND2_X1 U79 ( .A1(a[1]), .A2(b[13]), .ZN(y[29]) );
  OR2_X1 U79bar ( .A1(abar[1]), .A2(bbar[13]), .ZN(ybar[29]) );
  AND2_X1 U80 ( .A1(a[1]), .A2(b[12]), .ZN(y[28]) );
  OR2_X1 U80bar ( .A1(abar[1]), .A2(bbar[12]), .ZN(ybar[28]) );
  AND2_X1 U81 ( .A1(a[1]), .A2(b[11]), .ZN(y[27]) );
  OR2_X1 U81bar ( .A1(abar[1]), .A2(bbar[11]), .ZN(ybar[27]) );
  AND2_X1 U82 ( .A1(a[1]), .A2(b[10]), .ZN(y[26]) );
  OR2_X1 U82bar ( .A1(abar[1]), .A2(bbar[10]), .ZN(ybar[26]) );
  AND2_X1 U83 ( .A1(a[1]), .A2(b[9]), .ZN(y[25]) );
  OR2_X1 U83bar ( .A1(abar[1]), .A2(bbar[9]), .ZN(ybar[25]) );
  AND2_X1 U84 ( .A1(a[15]), .A2(b[15]), .ZN(y[255]) );
  OR2_X1 U84bar ( .A1(abar[15]), .A2(bbar[15]), .ZN(ybar[255]) );
  AND2_X1 U85 ( .A1(a[15]), .A2(b[14]), .ZN(y[254]) );
  OR2_X1 U85bar ( .A1(abar[15]), .A2(bbar[14]), .ZN(ybar[254]) );
  AND2_X1 U86 ( .A1(a[15]), .A2(b[13]), .ZN(y[253]) );
  OR2_X1 U86bar ( .A1(abar[15]), .A2(bbar[13]), .ZN(ybar[253]) );
  AND2_X1 U87 ( .A1(a[15]), .A2(b[12]), .ZN(y[252]) );
  OR2_X1 U87bar ( .A1(abar[15]), .A2(bbar[12]), .ZN(ybar[252]) );
  AND2_X1 U88 ( .A1(a[15]), .A2(b[11]), .ZN(y[251]) );
  OR2_X1 U88bar ( .A1(abar[15]), .A2(bbar[11]), .ZN(ybar[251]) );
  AND2_X1 U89 ( .A1(a[15]), .A2(b[10]), .ZN(y[250]) );
  OR2_X1 U89bar ( .A1(abar[15]), .A2(bbar[10]), .ZN(ybar[250]) );
  AND2_X1 U90 ( .A1(a[1]), .A2(b[8]), .ZN(y[24]) );
  OR2_X1 U90bar ( .A1(abar[1]), .A2(bbar[8]), .ZN(ybar[24]) );
  AND2_X1 U91 ( .A1(a[15]), .A2(b[9]), .ZN(y[249]) );
  OR2_X1 U91bar ( .A1(abar[15]), .A2(bbar[9]), .ZN(ybar[249]) );
  AND2_X1 U92 ( .A1(a[15]), .A2(b[8]), .ZN(y[248]) );
  OR2_X1 U92bar ( .A1(abar[15]), .A2(bbar[8]), .ZN(ybar[248]) );
  AND2_X1 U93 ( .A1(a[15]), .A2(b[7]), .ZN(y[247]) );
  OR2_X1 U93bar ( .A1(abar[15]), .A2(bbar[7]), .ZN(ybar[247]) );
  AND2_X1 U94 ( .A1(a[15]), .A2(b[6]), .ZN(y[246]) );
  OR2_X1 U94bar ( .A1(abar[15]), .A2(bbar[6]), .ZN(ybar[246]) );
  AND2_X1 U95 ( .A1(a[15]), .A2(b[5]), .ZN(y[245]) );
  OR2_X1 U95bar ( .A1(abar[15]), .A2(bbar[5]), .ZN(ybar[245]) );
  AND2_X1 U96 ( .A1(a[15]), .A2(b[4]), .ZN(y[244]) );
  OR2_X1 U96bar ( .A1(abar[15]), .A2(bbar[4]), .ZN(ybar[244]) );
  AND2_X1 U97 ( .A1(a[15]), .A2(b[3]), .ZN(y[243]) );
  OR2_X1 U97bar ( .A1(abar[15]), .A2(bbar[3]), .ZN(ybar[243]) );
  AND2_X1 U98 ( .A1(a[15]), .A2(b[2]), .ZN(y[242]) );
  OR2_X1 U98bar ( .A1(abar[15]), .A2(bbar[2]), .ZN(ybar[242]) );
  AND2_X1 U99 ( .A1(a[15]), .A2(b[1]), .ZN(y[241]) );
  OR2_X1 U99bar ( .A1(abar[15]), .A2(bbar[1]), .ZN(ybar[241]) );
  AND2_X1 U100 ( .A1(a[15]), .A2(b[0]), .ZN(y[240]) );
  OR2_X1 U100bar ( .A1(abar[15]), .A2(bbar[0]), .ZN(ybar[240]) );
  AND2_X1 U101 ( .A1(a[1]), .A2(b[7]), .ZN(y[23]) );
  OR2_X1 U101bar ( .A1(abar[1]), .A2(bbar[7]), .ZN(ybar[23]) );
  AND2_X1 U102 ( .A1(a[14]), .A2(b[15]), .ZN(y[239]) );
  OR2_X1 U102bar ( .A1(abar[14]), .A2(bbar[15]), .ZN(ybar[239]) );
  AND2_X1 U103 ( .A1(a[14]), .A2(b[14]), .ZN(y[238]) );
  OR2_X1 U103bar ( .A1(abar[14]), .A2(bbar[14]), .ZN(ybar[238]) );
  AND2_X1 U104 ( .A1(a[14]), .A2(b[13]), .ZN(y[237]) );
  OR2_X1 U104bar ( .A1(abar[14]), .A2(bbar[13]), .ZN(ybar[237]) );
  AND2_X1 U105 ( .A1(a[14]), .A2(b[12]), .ZN(y[236]) );
  OR2_X1 U105bar ( .A1(abar[14]), .A2(bbar[12]), .ZN(ybar[236]) );
  AND2_X1 U106 ( .A1(a[14]), .A2(b[11]), .ZN(y[235]) );
  OR2_X1 U106bar ( .A1(abar[14]), .A2(bbar[11]), .ZN(ybar[235]) );
  AND2_X1 U107 ( .A1(a[14]), .A2(b[10]), .ZN(y[234]) );
  OR2_X1 U107bar ( .A1(abar[14]), .A2(bbar[10]), .ZN(ybar[234]) );
  AND2_X1 U108 ( .A1(a[14]), .A2(b[9]), .ZN(y[233]) );
  OR2_X1 U108bar ( .A1(abar[14]), .A2(bbar[9]), .ZN(ybar[233]) );
  AND2_X1 U109 ( .A1(a[14]), .A2(b[8]), .ZN(y[232]) );
  OR2_X1 U109bar ( .A1(abar[14]), .A2(bbar[8]), .ZN(ybar[232]) );
  AND2_X1 U110 ( .A1(a[14]), .A2(b[7]), .ZN(y[231]) );
  OR2_X1 U110bar ( .A1(abar[14]), .A2(bbar[7]), .ZN(ybar[231]) );
  AND2_X1 U111 ( .A1(a[14]), .A2(b[6]), .ZN(y[230]) );
  OR2_X1 U111bar ( .A1(abar[14]), .A2(bbar[6]), .ZN(ybar[230]) );
  AND2_X1 U112 ( .A1(a[1]), .A2(b[6]), .ZN(y[22]) );
  OR2_X1 U112bar ( .A1(abar[1]), .A2(bbar[6]), .ZN(ybar[22]) );
  AND2_X1 U113 ( .A1(a[14]), .A2(b[5]), .ZN(y[229]) );
  OR2_X1 U113bar ( .A1(abar[14]), .A2(bbar[5]), .ZN(ybar[229]) );
  AND2_X1 U114 ( .A1(a[14]), .A2(b[4]), .ZN(y[228]) );
  OR2_X1 U114bar ( .A1(abar[14]), .A2(bbar[4]), .ZN(ybar[228]) );
  AND2_X1 U115 ( .A1(a[14]), .A2(b[3]), .ZN(y[227]) );
  OR2_X1 U115bar ( .A1(abar[14]), .A2(bbar[3]), .ZN(ybar[227]) );
  AND2_X1 U116 ( .A1(a[14]), .A2(b[2]), .ZN(y[226]) );
  OR2_X1 U116bar ( .A1(abar[14]), .A2(bbar[2]), .ZN(ybar[226]) );
  AND2_X1 U117 ( .A1(a[14]), .A2(b[1]), .ZN(y[225]) );
  OR2_X1 U117bar ( .A1(abar[14]), .A2(bbar[1]), .ZN(ybar[225]) );
  AND2_X1 U118 ( .A1(a[14]), .A2(b[0]), .ZN(y[224]) );
  OR2_X1 U118bar ( .A1(abar[14]), .A2(bbar[0]), .ZN(ybar[224]) );
  AND2_X1 U119 ( .A1(a[13]), .A2(b[15]), .ZN(y[223]) );
  OR2_X1 U119bar ( .A1(abar[13]), .A2(bbar[15]), .ZN(ybar[223]) );
  AND2_X1 U120 ( .A1(a[13]), .A2(b[14]), .ZN(y[222]) );
  OR2_X1 U120bar ( .A1(abar[13]), .A2(bbar[14]), .ZN(ybar[222]) );
  AND2_X1 U121 ( .A1(a[13]), .A2(b[13]), .ZN(y[221]) );
  OR2_X1 U121bar ( .A1(abar[13]), .A2(bbar[13]), .ZN(ybar[221]) );
  AND2_X1 U122 ( .A1(a[13]), .A2(b[12]), .ZN(y[220]) );
  OR2_X1 U122bar ( .A1(abar[13]), .A2(bbar[12]), .ZN(ybar[220]) );
  AND2_X1 U123 ( .A1(a[1]), .A2(b[5]), .ZN(y[21]) );
  OR2_X1 U123bar ( .A1(abar[1]), .A2(bbar[5]), .ZN(ybar[21]) );
  AND2_X1 U124 ( .A1(a[13]), .A2(b[11]), .ZN(y[219]) );
  OR2_X1 U124bar ( .A1(abar[13]), .A2(bbar[11]), .ZN(ybar[219]) );
  AND2_X1 U125 ( .A1(a[13]), .A2(b[10]), .ZN(y[218]) );
  OR2_X1 U125bar ( .A1(abar[13]), .A2(bbar[10]), .ZN(ybar[218]) );
  AND2_X1 U126 ( .A1(a[13]), .A2(b[9]), .ZN(y[217]) );
  OR2_X1 U126bar ( .A1(abar[13]), .A2(bbar[9]), .ZN(ybar[217]) );
  AND2_X1 U127 ( .A1(a[13]), .A2(b[8]), .ZN(y[216]) );
  OR2_X1 U127bar ( .A1(abar[13]), .A2(bbar[8]), .ZN(ybar[216]) );
  AND2_X1 U128 ( .A1(a[13]), .A2(b[7]), .ZN(y[215]) );
  OR2_X1 U128bar ( .A1(abar[13]), .A2(bbar[7]), .ZN(ybar[215]) );
  AND2_X1 U129 ( .A1(a[13]), .A2(b[6]), .ZN(y[214]) );
  OR2_X1 U129bar ( .A1(abar[13]), .A2(bbar[6]), .ZN(ybar[214]) );
  AND2_X1 U130 ( .A1(a[13]), .A2(b[5]), .ZN(y[213]) );
  OR2_X1 U130bar ( .A1(abar[13]), .A2(bbar[5]), .ZN(ybar[213]) );
  AND2_X1 U131 ( .A1(a[13]), .A2(b[4]), .ZN(y[212]) );
  OR2_X1 U131bar ( .A1(abar[13]), .A2(bbar[4]), .ZN(ybar[212]) );
  AND2_X1 U132 ( .A1(a[13]), .A2(b[3]), .ZN(y[211]) );
  OR2_X1 U132bar ( .A1(abar[13]), .A2(bbar[3]), .ZN(ybar[211]) );
  AND2_X1 U133 ( .A1(a[13]), .A2(b[2]), .ZN(y[210]) );
  OR2_X1 U133bar ( .A1(abar[13]), .A2(bbar[2]), .ZN(ybar[210]) );
  AND2_X1 U134 ( .A1(a[1]), .A2(b[4]), .ZN(y[20]) );
  OR2_X1 U134bar ( .A1(abar[1]), .A2(bbar[4]), .ZN(ybar[20]) );
  AND2_X1 U135 ( .A1(a[13]), .A2(b[1]), .ZN(y[209]) );
  OR2_X1 U135bar ( .A1(abar[13]), .A2(bbar[1]), .ZN(ybar[209]) );
  AND2_X1 U136 ( .A1(a[13]), .A2(b[0]), .ZN(y[208]) );
  OR2_X1 U136bar ( .A1(abar[13]), .A2(bbar[0]), .ZN(ybar[208]) );
  AND2_X1 U137 ( .A1(a[12]), .A2(b[15]), .ZN(y[207]) );
  OR2_X1 U137bar ( .A1(abar[12]), .A2(bbar[15]), .ZN(ybar[207]) );
  AND2_X1 U138 ( .A1(a[12]), .A2(b[14]), .ZN(y[206]) );
  OR2_X1 U138bar ( .A1(abar[12]), .A2(bbar[14]), .ZN(ybar[206]) );
  AND2_X1 U139 ( .A1(a[12]), .A2(b[13]), .ZN(y[205]) );
  OR2_X1 U139bar ( .A1(abar[12]), .A2(bbar[13]), .ZN(ybar[205]) );
  AND2_X1 U140 ( .A1(a[12]), .A2(b[12]), .ZN(y[204]) );
  OR2_X1 U140bar ( .A1(abar[12]), .A2(bbar[12]), .ZN(ybar[204]) );
  AND2_X1 U141 ( .A1(a[12]), .A2(b[11]), .ZN(y[203]) );
  OR2_X1 U141bar ( .A1(abar[12]), .A2(bbar[11]), .ZN(ybar[203]) );
  AND2_X1 U142 ( .A1(a[12]), .A2(b[10]), .ZN(y[202]) );
  OR2_X1 U142bar ( .A1(abar[12]), .A2(bbar[10]), .ZN(ybar[202]) );
  AND2_X1 U143 ( .A1(a[12]), .A2(b[9]), .ZN(y[201]) );
  OR2_X1 U143bar ( .A1(abar[12]), .A2(bbar[9]), .ZN(ybar[201]) );
  AND2_X1 U144 ( .A1(a[12]), .A2(b[8]), .ZN(y[200]) );
  OR2_X1 U144bar ( .A1(abar[12]), .A2(bbar[8]), .ZN(ybar[200]) );
  AND2_X1 U145 ( .A1(b[1]), .A2(a[0]), .ZN(y[1]) );
  OR2_X1 U145bar ( .A1(bbar[1]), .A2(abar[0]), .ZN(ybar[1]) );
  AND2_X1 U146 ( .A1(a[1]), .A2(b[3]), .ZN(y[19]) );
  OR2_X1 U146bar ( .A1(abar[1]), .A2(bbar[3]), .ZN(ybar[19]) );
  AND2_X1 U147 ( .A1(a[12]), .A2(b[7]), .ZN(y[199]) );
  OR2_X1 U147bar ( .A1(abar[12]), .A2(bbar[7]), .ZN(ybar[199]) );
  AND2_X1 U148 ( .A1(a[12]), .A2(b[6]), .ZN(y[198]) );
  OR2_X1 U148bar ( .A1(abar[12]), .A2(bbar[6]), .ZN(ybar[198]) );
  AND2_X1 U149 ( .A1(a[12]), .A2(b[5]), .ZN(y[197]) );
  OR2_X1 U149bar ( .A1(abar[12]), .A2(bbar[5]), .ZN(ybar[197]) );
  AND2_X1 U150 ( .A1(a[12]), .A2(b[4]), .ZN(y[196]) );
  OR2_X1 U150bar ( .A1(abar[12]), .A2(bbar[4]), .ZN(ybar[196]) );
  AND2_X1 U151 ( .A1(a[12]), .A2(b[3]), .ZN(y[195]) );
  OR2_X1 U151bar ( .A1(abar[12]), .A2(bbar[3]), .ZN(ybar[195]) );
  AND2_X1 U152 ( .A1(a[12]), .A2(b[2]), .ZN(y[194]) );
  OR2_X1 U152bar ( .A1(abar[12]), .A2(bbar[2]), .ZN(ybar[194]) );
  AND2_X1 U153 ( .A1(a[12]), .A2(b[1]), .ZN(y[193]) );
  OR2_X1 U153bar ( .A1(abar[12]), .A2(bbar[1]), .ZN(ybar[193]) );
  AND2_X1 U154 ( .A1(a[12]), .A2(b[0]), .ZN(y[192]) );
  OR2_X1 U154bar ( .A1(abar[12]), .A2(bbar[0]), .ZN(ybar[192]) );
  AND2_X1 U155 ( .A1(a[11]), .A2(b[15]), .ZN(y[191]) );
  OR2_X1 U155bar ( .A1(abar[11]), .A2(bbar[15]), .ZN(ybar[191]) );
  AND2_X1 U156 ( .A1(a[11]), .A2(b[14]), .ZN(y[190]) );
  OR2_X1 U156bar ( .A1(abar[11]), .A2(bbar[14]), .ZN(ybar[190]) );
  AND2_X1 U157 ( .A1(a[1]), .A2(b[2]), .ZN(y[18]) );
  OR2_X1 U157bar ( .A1(abar[1]), .A2(bbar[2]), .ZN(ybar[18]) );
  AND2_X1 U158 ( .A1(a[11]), .A2(b[13]), .ZN(y[189]) );
  OR2_X1 U158bar ( .A1(abar[11]), .A2(bbar[13]), .ZN(ybar[189]) );
  AND2_X1 U159 ( .A1(a[11]), .A2(b[12]), .ZN(y[188]) );
  OR2_X1 U159bar ( .A1(abar[11]), .A2(bbar[12]), .ZN(ybar[188]) );
  AND2_X1 U160 ( .A1(a[11]), .A2(b[11]), .ZN(y[187]) );
  OR2_X1 U160bar ( .A1(abar[11]), .A2(bbar[11]), .ZN(ybar[187]) );
  AND2_X1 U161 ( .A1(a[11]), .A2(b[10]), .ZN(y[186]) );
  OR2_X1 U161bar ( .A1(abar[11]), .A2(bbar[10]), .ZN(ybar[186]) );
  AND2_X1 U162 ( .A1(a[11]), .A2(b[9]), .ZN(y[185]) );
  OR2_X1 U162bar ( .A1(abar[11]), .A2(bbar[9]), .ZN(ybar[185]) );
  AND2_X1 U163 ( .A1(a[11]), .A2(b[8]), .ZN(y[184]) );
  OR2_X1 U163bar ( .A1(abar[11]), .A2(bbar[8]), .ZN(ybar[184]) );
  AND2_X1 U164 ( .A1(a[11]), .A2(b[7]), .ZN(y[183]) );
  OR2_X1 U164bar ( .A1(abar[11]), .A2(bbar[7]), .ZN(ybar[183]) );
  AND2_X1 U165 ( .A1(a[11]), .A2(b[6]), .ZN(y[182]) );
  OR2_X1 U165bar ( .A1(abar[11]), .A2(bbar[6]), .ZN(ybar[182]) );
  AND2_X1 U166 ( .A1(a[11]), .A2(b[5]), .ZN(y[181]) );
  OR2_X1 U166bar ( .A1(abar[11]), .A2(bbar[5]), .ZN(ybar[181]) );
  AND2_X1 U167 ( .A1(a[11]), .A2(b[4]), .ZN(y[180]) );
  OR2_X1 U167bar ( .A1(abar[11]), .A2(bbar[4]), .ZN(ybar[180]) );
  AND2_X1 U168 ( .A1(a[1]), .A2(b[1]), .ZN(y[17]) );
  OR2_X1 U168bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[17]) );
  AND2_X1 U169 ( .A1(a[11]), .A2(b[3]), .ZN(y[179]) );
  OR2_X1 U169bar ( .A1(abar[11]), .A2(bbar[3]), .ZN(ybar[179]) );
  AND2_X1 U170 ( .A1(a[11]), .A2(b[2]), .ZN(y[178]) );
  OR2_X1 U170bar ( .A1(abar[11]), .A2(bbar[2]), .ZN(ybar[178]) );
  AND2_X1 U171 ( .A1(a[11]), .A2(b[1]), .ZN(y[177]) );
  OR2_X1 U171bar ( .A1(abar[11]), .A2(bbar[1]), .ZN(ybar[177]) );
  AND2_X1 U172 ( .A1(a[11]), .A2(b[0]), .ZN(y[176]) );
  OR2_X1 U172bar ( .A1(abar[11]), .A2(bbar[0]), .ZN(ybar[176]) );
  AND2_X1 U173 ( .A1(a[10]), .A2(b[15]), .ZN(y[175]) );
  OR2_X1 U173bar ( .A1(abar[10]), .A2(bbar[15]), .ZN(ybar[175]) );
  AND2_X1 U174 ( .A1(a[10]), .A2(b[14]), .ZN(y[174]) );
  OR2_X1 U174bar ( .A1(abar[10]), .A2(bbar[14]), .ZN(ybar[174]) );
  AND2_X1 U175 ( .A1(a[10]), .A2(b[13]), .ZN(y[173]) );
  OR2_X1 U175bar ( .A1(abar[10]), .A2(bbar[13]), .ZN(ybar[173]) );
  AND2_X1 U176 ( .A1(a[10]), .A2(b[12]), .ZN(y[172]) );
  OR2_X1 U176bar ( .A1(abar[10]), .A2(bbar[12]), .ZN(ybar[172]) );
  AND2_X1 U177 ( .A1(a[10]), .A2(b[11]), .ZN(y[171]) );
  OR2_X1 U177bar ( .A1(abar[10]), .A2(bbar[11]), .ZN(ybar[171]) );
  AND2_X1 U178 ( .A1(a[10]), .A2(b[10]), .ZN(y[170]) );
  OR2_X1 U178bar ( .A1(abar[10]), .A2(bbar[10]), .ZN(ybar[170]) );
  AND2_X1 U179 ( .A1(a[1]), .A2(b[0]), .ZN(y[16]) );
  OR2_X1 U179bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[16]) );
  AND2_X1 U180 ( .A1(a[10]), .A2(b[9]), .ZN(y[169]) );
  OR2_X1 U180bar ( .A1(abar[10]), .A2(bbar[9]), .ZN(ybar[169]) );
  AND2_X1 U181 ( .A1(a[10]), .A2(b[8]), .ZN(y[168]) );
  OR2_X1 U181bar ( .A1(abar[10]), .A2(bbar[8]), .ZN(ybar[168]) );
  AND2_X1 U182 ( .A1(a[10]), .A2(b[7]), .ZN(y[167]) );
  OR2_X1 U182bar ( .A1(abar[10]), .A2(bbar[7]), .ZN(ybar[167]) );
  AND2_X1 U183 ( .A1(a[10]), .A2(b[6]), .ZN(y[166]) );
  OR2_X1 U183bar ( .A1(abar[10]), .A2(bbar[6]), .ZN(ybar[166]) );
  AND2_X1 U184 ( .A1(a[10]), .A2(b[5]), .ZN(y[165]) );
  OR2_X1 U184bar ( .A1(abar[10]), .A2(bbar[5]), .ZN(ybar[165]) );
  AND2_X1 U185 ( .A1(a[10]), .A2(b[4]), .ZN(y[164]) );
  OR2_X1 U185bar ( .A1(abar[10]), .A2(bbar[4]), .ZN(ybar[164]) );
  AND2_X1 U186 ( .A1(a[10]), .A2(b[3]), .ZN(y[163]) );
  OR2_X1 U186bar ( .A1(abar[10]), .A2(bbar[3]), .ZN(ybar[163]) );
  AND2_X1 U187 ( .A1(a[10]), .A2(b[2]), .ZN(y[162]) );
  OR2_X1 U187bar ( .A1(abar[10]), .A2(bbar[2]), .ZN(ybar[162]) );
  AND2_X1 U188 ( .A1(a[10]), .A2(b[1]), .ZN(y[161]) );
  OR2_X1 U188bar ( .A1(abar[10]), .A2(bbar[1]), .ZN(ybar[161]) );
  AND2_X1 U189 ( .A1(a[10]), .A2(b[0]), .ZN(y[160]) );
  OR2_X1 U189bar ( .A1(abar[10]), .A2(bbar[0]), .ZN(ybar[160]) );
  AND2_X1 U190 ( .A1(b[15]), .A2(a[0]), .ZN(y[15]) );
  OR2_X1 U190bar ( .A1(bbar[15]), .A2(abar[0]), .ZN(ybar[15]) );
  AND2_X1 U191 ( .A1(a[9]), .A2(b[15]), .ZN(y[159]) );
  OR2_X1 U191bar ( .A1(abar[9]), .A2(bbar[15]), .ZN(ybar[159]) );
  AND2_X1 U192 ( .A1(a[9]), .A2(b[14]), .ZN(y[158]) );
  OR2_X1 U192bar ( .A1(abar[9]), .A2(bbar[14]), .ZN(ybar[158]) );
  AND2_X1 U193 ( .A1(a[9]), .A2(b[13]), .ZN(y[157]) );
  OR2_X1 U193bar ( .A1(abar[9]), .A2(bbar[13]), .ZN(ybar[157]) );
  AND2_X1 U194 ( .A1(a[9]), .A2(b[12]), .ZN(y[156]) );
  OR2_X1 U194bar ( .A1(abar[9]), .A2(bbar[12]), .ZN(ybar[156]) );
  AND2_X1 U195 ( .A1(a[9]), .A2(b[11]), .ZN(y[155]) );
  OR2_X1 U195bar ( .A1(abar[9]), .A2(bbar[11]), .ZN(ybar[155]) );
  AND2_X1 U196 ( .A1(a[9]), .A2(b[10]), .ZN(y[154]) );
  OR2_X1 U196bar ( .A1(abar[9]), .A2(bbar[10]), .ZN(ybar[154]) );
  AND2_X1 U197 ( .A1(a[9]), .A2(b[9]), .ZN(y[153]) );
  OR2_X1 U197bar ( .A1(abar[9]), .A2(bbar[9]), .ZN(ybar[153]) );
  AND2_X1 U198 ( .A1(a[9]), .A2(b[8]), .ZN(y[152]) );
  OR2_X1 U198bar ( .A1(abar[9]), .A2(bbar[8]), .ZN(ybar[152]) );
  AND2_X1 U199 ( .A1(a[9]), .A2(b[7]), .ZN(y[151]) );
  OR2_X1 U199bar ( .A1(abar[9]), .A2(bbar[7]), .ZN(ybar[151]) );
  AND2_X1 U200 ( .A1(a[9]), .A2(b[6]), .ZN(y[150]) );
  OR2_X1 U200bar ( .A1(abar[9]), .A2(bbar[6]), .ZN(ybar[150]) );
  AND2_X1 U201 ( .A1(b[14]), .A2(a[0]), .ZN(y[14]) );
  OR2_X1 U201bar ( .A1(bbar[14]), .A2(abar[0]), .ZN(ybar[14]) );
  AND2_X1 U202 ( .A1(a[9]), .A2(b[5]), .ZN(y[149]) );
  OR2_X1 U202bar ( .A1(abar[9]), .A2(bbar[5]), .ZN(ybar[149]) );
  AND2_X1 U203 ( .A1(a[9]), .A2(b[4]), .ZN(y[148]) );
  OR2_X1 U203bar ( .A1(abar[9]), .A2(bbar[4]), .ZN(ybar[148]) );
  AND2_X1 U204 ( .A1(a[9]), .A2(b[3]), .ZN(y[147]) );
  OR2_X1 U204bar ( .A1(abar[9]), .A2(bbar[3]), .ZN(ybar[147]) );
  AND2_X1 U205 ( .A1(a[9]), .A2(b[2]), .ZN(y[146]) );
  OR2_X1 U205bar ( .A1(abar[9]), .A2(bbar[2]), .ZN(ybar[146]) );
  AND2_X1 U206 ( .A1(a[9]), .A2(b[1]), .ZN(y[145]) );
  OR2_X1 U206bar ( .A1(abar[9]), .A2(bbar[1]), .ZN(ybar[145]) );
  AND2_X1 U207 ( .A1(a[9]), .A2(b[0]), .ZN(y[144]) );
  OR2_X1 U207bar ( .A1(abar[9]), .A2(bbar[0]), .ZN(ybar[144]) );
  AND2_X1 U208 ( .A1(a[8]), .A2(b[15]), .ZN(y[143]) );
  OR2_X1 U208bar ( .A1(abar[8]), .A2(bbar[15]), .ZN(ybar[143]) );
  AND2_X1 U209 ( .A1(a[8]), .A2(b[14]), .ZN(y[142]) );
  OR2_X1 U209bar ( .A1(abar[8]), .A2(bbar[14]), .ZN(ybar[142]) );
  AND2_X1 U210 ( .A1(a[8]), .A2(b[13]), .ZN(y[141]) );
  OR2_X1 U210bar ( .A1(abar[8]), .A2(bbar[13]), .ZN(ybar[141]) );
  AND2_X1 U211 ( .A1(a[8]), .A2(b[12]), .ZN(y[140]) );
  OR2_X1 U211bar ( .A1(abar[8]), .A2(bbar[12]), .ZN(ybar[140]) );
  AND2_X1 U212 ( .A1(b[13]), .A2(a[0]), .ZN(y[13]) );
  OR2_X1 U212bar ( .A1(bbar[13]), .A2(abar[0]), .ZN(ybar[13]) );
  AND2_X1 U213 ( .A1(a[8]), .A2(b[11]), .ZN(y[139]) );
  OR2_X1 U213bar ( .A1(abar[8]), .A2(bbar[11]), .ZN(ybar[139]) );
  AND2_X1 U214 ( .A1(a[8]), .A2(b[10]), .ZN(y[138]) );
  OR2_X1 U214bar ( .A1(abar[8]), .A2(bbar[10]), .ZN(ybar[138]) );
  AND2_X1 U215 ( .A1(a[8]), .A2(b[9]), .ZN(y[137]) );
  OR2_X1 U215bar ( .A1(abar[8]), .A2(bbar[9]), .ZN(ybar[137]) );
  AND2_X1 U216 ( .A1(a[8]), .A2(b[8]), .ZN(y[136]) );
  OR2_X1 U216bar ( .A1(abar[8]), .A2(bbar[8]), .ZN(ybar[136]) );
  AND2_X1 U217 ( .A1(a[8]), .A2(b[7]), .ZN(y[135]) );
  OR2_X1 U217bar ( .A1(abar[8]), .A2(bbar[7]), .ZN(ybar[135]) );
  AND2_X1 U218 ( .A1(a[8]), .A2(b[6]), .ZN(y[134]) );
  OR2_X1 U218bar ( .A1(abar[8]), .A2(bbar[6]), .ZN(ybar[134]) );
  AND2_X1 U219 ( .A1(a[8]), .A2(b[5]), .ZN(y[133]) );
  OR2_X1 U219bar ( .A1(abar[8]), .A2(bbar[5]), .ZN(ybar[133]) );
  AND2_X1 U220 ( .A1(a[8]), .A2(b[4]), .ZN(y[132]) );
  OR2_X1 U220bar ( .A1(abar[8]), .A2(bbar[4]), .ZN(ybar[132]) );
  AND2_X1 U221 ( .A1(a[8]), .A2(b[3]), .ZN(y[131]) );
  OR2_X1 U221bar ( .A1(abar[8]), .A2(bbar[3]), .ZN(ybar[131]) );
  AND2_X1 U222 ( .A1(a[8]), .A2(b[2]), .ZN(y[130]) );
  OR2_X1 U222bar ( .A1(abar[8]), .A2(bbar[2]), .ZN(ybar[130]) );
  AND2_X1 U223 ( .A1(b[12]), .A2(a[0]), .ZN(y[12]) );
  OR2_X1 U223bar ( .A1(bbar[12]), .A2(abar[0]), .ZN(ybar[12]) );
  AND2_X1 U224 ( .A1(a[8]), .A2(b[1]), .ZN(y[129]) );
  OR2_X1 U224bar ( .A1(abar[8]), .A2(bbar[1]), .ZN(ybar[129]) );
  AND2_X1 U225 ( .A1(a[8]), .A2(b[0]), .ZN(y[128]) );
  OR2_X1 U225bar ( .A1(abar[8]), .A2(bbar[0]), .ZN(ybar[128]) );
  AND2_X1 U226 ( .A1(a[7]), .A2(b[15]), .ZN(y[127]) );
  OR2_X1 U226bar ( .A1(abar[7]), .A2(bbar[15]), .ZN(ybar[127]) );
  AND2_X1 U227 ( .A1(a[7]), .A2(b[14]), .ZN(y[126]) );
  OR2_X1 U227bar ( .A1(abar[7]), .A2(bbar[14]), .ZN(ybar[126]) );
  AND2_X1 U228 ( .A1(a[7]), .A2(b[13]), .ZN(y[125]) );
  OR2_X1 U228bar ( .A1(abar[7]), .A2(bbar[13]), .ZN(ybar[125]) );
  AND2_X1 U229 ( .A1(a[7]), .A2(b[12]), .ZN(y[124]) );
  OR2_X1 U229bar ( .A1(abar[7]), .A2(bbar[12]), .ZN(ybar[124]) );
  AND2_X1 U230 ( .A1(a[7]), .A2(b[11]), .ZN(y[123]) );
  OR2_X1 U230bar ( .A1(abar[7]), .A2(bbar[11]), .ZN(ybar[123]) );
  AND2_X1 U231 ( .A1(a[7]), .A2(b[10]), .ZN(y[122]) );
  OR2_X1 U231bar ( .A1(abar[7]), .A2(bbar[10]), .ZN(ybar[122]) );
  AND2_X1 U232 ( .A1(a[7]), .A2(b[9]), .ZN(y[121]) );
  OR2_X1 U232bar ( .A1(abar[7]), .A2(bbar[9]), .ZN(ybar[121]) );
  AND2_X1 U233 ( .A1(a[7]), .A2(b[8]), .ZN(y[120]) );
  OR2_X1 U233bar ( .A1(abar[7]), .A2(bbar[8]), .ZN(ybar[120]) );
  AND2_X1 U234 ( .A1(b[11]), .A2(a[0]), .ZN(y[11]) );
  OR2_X1 U234bar ( .A1(bbar[11]), .A2(abar[0]), .ZN(ybar[11]) );
  AND2_X1 U235 ( .A1(a[7]), .A2(b[7]), .ZN(y[119]) );
  OR2_X1 U235bar ( .A1(abar[7]), .A2(bbar[7]), .ZN(ybar[119]) );
  AND2_X1 U236 ( .A1(a[7]), .A2(b[6]), .ZN(y[118]) );
  OR2_X1 U236bar ( .A1(abar[7]), .A2(bbar[6]), .ZN(ybar[118]) );
  AND2_X1 U237 ( .A1(a[7]), .A2(b[5]), .ZN(y[117]) );
  OR2_X1 U237bar ( .A1(abar[7]), .A2(bbar[5]), .ZN(ybar[117]) );
  AND2_X1 U238 ( .A1(a[7]), .A2(b[4]), .ZN(y[116]) );
  OR2_X1 U238bar ( .A1(abar[7]), .A2(bbar[4]), .ZN(ybar[116]) );
  AND2_X1 U239 ( .A1(a[7]), .A2(b[3]), .ZN(y[115]) );
  OR2_X1 U239bar ( .A1(abar[7]), .A2(bbar[3]), .ZN(ybar[115]) );
  AND2_X1 U240 ( .A1(a[7]), .A2(b[2]), .ZN(y[114]) );
  OR2_X1 U240bar ( .A1(abar[7]), .A2(bbar[2]), .ZN(ybar[114]) );
  AND2_X1 U241 ( .A1(a[7]), .A2(b[1]), .ZN(y[113]) );
  OR2_X1 U241bar ( .A1(abar[7]), .A2(bbar[1]), .ZN(ybar[113]) );
  AND2_X1 U242 ( .A1(a[7]), .A2(b[0]), .ZN(y[112]) );
  OR2_X1 U242bar ( .A1(abar[7]), .A2(bbar[0]), .ZN(ybar[112]) );
  AND2_X1 U243 ( .A1(b[15]), .A2(a[6]), .ZN(y[111]) );
  OR2_X1 U243bar ( .A1(bbar[15]), .A2(abar[6]), .ZN(ybar[111]) );
  AND2_X1 U244 ( .A1(b[14]), .A2(a[6]), .ZN(y[110]) );
  OR2_X1 U244bar ( .A1(bbar[14]), .A2(abar[6]), .ZN(ybar[110]) );
  AND2_X1 U245 ( .A1(b[10]), .A2(a[0]), .ZN(y[10]) );
  OR2_X1 U245bar ( .A1(bbar[10]), .A2(abar[0]), .ZN(ybar[10]) );
  AND2_X1 U246 ( .A1(b[13]), .A2(a[6]), .ZN(y[109]) );
  OR2_X1 U246bar ( .A1(bbar[13]), .A2(abar[6]), .ZN(ybar[109]) );
  AND2_X1 U247 ( .A1(b[12]), .A2(a[6]), .ZN(y[108]) );
  OR2_X1 U247bar ( .A1(bbar[12]), .A2(abar[6]), .ZN(ybar[108]) );
  AND2_X1 U248 ( .A1(b[11]), .A2(a[6]), .ZN(y[107]) );
  OR2_X1 U248bar ( .A1(bbar[11]), .A2(abar[6]), .ZN(ybar[107]) );
  AND2_X1 U249 ( .A1(b[10]), .A2(a[6]), .ZN(y[106]) );
  OR2_X1 U249bar ( .A1(bbar[10]), .A2(abar[6]), .ZN(ybar[106]) );
  AND2_X1 U250 ( .A1(a[6]), .A2(b[9]), .ZN(y[105]) );
  OR2_X1 U250bar ( .A1(abar[6]), .A2(bbar[9]), .ZN(ybar[105]) );
  AND2_X1 U251 ( .A1(b[8]), .A2(a[6]), .ZN(y[104]) );
  OR2_X1 U251bar ( .A1(bbar[8]), .A2(abar[6]), .ZN(ybar[104]) );
  AND2_X1 U252 ( .A1(b[7]), .A2(a[6]), .ZN(y[103]) );
  OR2_X1 U252bar ( .A1(bbar[7]), .A2(abar[6]), .ZN(ybar[103]) );
  AND2_X1 U253 ( .A1(b[6]), .A2(a[6]), .ZN(y[102]) );
  OR2_X1 U253bar ( .A1(bbar[6]), .A2(abar[6]), .ZN(ybar[102]) );
  AND2_X1 U254 ( .A1(b[5]), .A2(a[6]), .ZN(y[101]) );
  OR2_X1 U254bar ( .A1(bbar[5]), .A2(abar[6]), .ZN(ybar[101]) );
  AND2_X1 U255 ( .A1(b[4]), .A2(a[6]), .ZN(y[100]) );
  OR2_X1 U255bar ( .A1(bbar[4]), .A2(abar[6]), .ZN(ybar[100]) );
  AND2_X1 U256 ( .A1(b[0]), .A2(a[0]), .ZN(y[0]) );
  OR2_X1 U256bar ( .A1(bbar[0]), .A2(abar[0]), .ZN(ybar[0]) );
endmodule

module decode_8 ( in, inbar, out, outbar );

  input wire [7:0] in;
  input wire [7:0] inbar;
//input_done

  output wire [255:0] out;
  output wire [255:0] outbar;
//output_done

  wire [15:0] level1;
  wire [31:0] level2;
  wire [15:0] level1bar;
  wire [31:0] level2bar;
//wire_done

  CD2_32 cd_l1_1 ( .a(in[1]), .abar(inbar[1]), .b(in[0]), .bbar(inbar[0]), .y(level1[3:0]), .ybar(level1bar[3:0]) );
  CD2_31 cd_l1_2 ( .a(in[3]), .abar(inbar[3]), .b(in[2]), .bbar(inbar[2]), .y(level1[7:4]), .ybar(level1bar[7:4]) );
  CD2_30 cd_l1_3 ( .a(in[5]), .abar(inbar[5]), .b(in[4]), .bbar(inbar[4]), .y(level1[11:8]), .ybar(level1bar[11:8]) );
  CD2_29 cd_l1_4 ( .a(in[7]), .abar(inbar[7]), .b(in[6]), .bbar(inbar[6]), .y(level1[15:12]), .ybar(level1bar[15:12]) );

  CD4_16 cd_l2_1 ( .a(level1[7:4]), .abar(level1bar[7:4]), .b(level1[3:0]), .bbar(level1bar[3:0]), 
        .y(level2[15:0]), .ybar(level2bar[15:0]) );
  CD4_15 cd_l2_2 ( .a(level1[15:12]), .abar(level1bar[15:12]), .b(level1[11:8]), .bbar(level1bar[11:8]), 
        .y(level2[31:16]), .ybar(level2bar[31:16]) );
  CD16_8 cd_l3 ( .a(level2[31:16]), .abar(level2bar[31:16]), .b(level2[15:0]), .bbar(level2bar[15:0]), 
        .y(out), .ybar(outbar) );
endmodule

module encode_8 ( in, inbar, out, outbar );

  input wire [255:0] in;
  input wire [255:0] inbar;
//input_done

  output wire [7:0] out;
  output wire [7:0] outbar;
//output_done

  wire in_81;
  wire in_80;
  wire in_79;
  wire in_78;
  wire in_77;
  wire in_76;
  wire in_75;
  wire in_74;
  wire in_73;
  wire in_72;
  wire in_71;
  wire in_70;
  wire in_69;
  wire in_68;
  wire in_67;
  wire in_66;
  wire in_65;
  wire in_64;
  wire in_63;
  wire in_62;
  wire in_61;
  wire in_60;
  wire in_59;
  wire in_58;
  wire in_57;
  wire in_56;
  wire in_55;
  wire in_54;
  wire in_53;
  wire in_52;
  wire in_51;
  wire in_50;
  wire in_49;
  wire in_48;
  wire in_47;
  wire in_46;
  wire in_45;
  wire in_44;
  wire in_43;
  wire in_42;
  wire in_41;
  wire in_40;
  wire in_39;
  wire in_38;
  wire in_37;
  wire in_36;
  wire in_35;
  wire in_34;
  wire in_33;
  wire in_32;
  wire in_31;
  wire in_30;
  wire in_29;
  wire in_28;
  wire in_27;
  wire in_26;
  wire in_25;
  wire in_24;
  wire in_23;
  wire in_22;
  wire in_21;
  wire in_20;
  wire in_19;
  wire in_18;
  wire in_17;
  wire in_16;
  wire in_15;
  wire in_14;
  wire in_13;
  wire in_12;
  wire in_11;
  wire in_10;
  wire in_9;
  wire in_8;
  wire in_7;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_3;
  wire in_2;
  wire in_1;
  wire in_0;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire in_81bar;
  wire in_80bar;
  wire in_79bar;
  wire in_78bar;
  wire in_77bar;
  wire in_76bar;
  wire in_75bar;
  wire in_74bar;
  wire in_73bar;
  wire in_72bar;
  wire in_71bar;
  wire in_70bar;
  wire in_69bar;
  wire in_68bar;
  wire in_67bar;
  wire in_66bar;
  wire in_65bar;
  wire in_64bar;
  wire in_63bar;
  wire in_62bar;
  wire in_61bar;
  wire in_60bar;
  wire in_59bar;
  wire in_58bar;
  wire in_57bar;
  wire in_56bar;
  wire in_55bar;
  wire in_54bar;
  wire in_53bar;
  wire in_52bar;
  wire in_51bar;
  wire in_50bar;
  wire in_49bar;
  wire in_48bar;
  wire in_47bar;
  wire in_46bar;
  wire in_45bar;
  wire in_44bar;
  wire in_43bar;
  wire in_42bar;
  wire in_41bar;
  wire in_40bar;
  wire in_39bar;
  wire in_38bar;
  wire in_37bar;
  wire in_36bar;
  wire in_35bar;
  wire in_34bar;
  wire in_33bar;
  wire in_32bar;
  wire in_31bar;
  wire in_30bar;
  wire in_29bar;
  wire in_28bar;
  wire in_27bar;
  wire in_26bar;
  wire in_25bar;
  wire in_24bar;
  wire in_23bar;
  wire in_22bar;
  wire in_21bar;
  wire in_20bar;
  wire in_19bar;
  wire in_18bar;
  wire in_17bar;
  wire in_16bar;
  wire in_15bar;
  wire in_14bar;
  wire in_13bar;
  wire in_12bar;
  wire in_11bar;
  wire in_10bar;
  wire in_9bar;
  wire in_8bar;
  wire in_7bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_3bar;
  wire in_2bar;
  wire in_1bar;
  wire in_0bar;
  wire n487bar;
  wire n488bar;
  wire n489bar;
  wire n490bar;
  wire n491bar;
  wire n492bar;
  wire n493bar;
  wire n494bar;
  wire n495bar;
  wire n496bar;
  wire n497bar;
  wire n498bar;
  wire n499bar;
  wire n500bar;
  wire n501bar;
  wire n502bar;
  wire n503bar;
  wire n504bar;
  wire n505bar;
  wire n506bar;
  wire n507bar;
  wire n508bar;
  wire n509bar;
  wire n510bar;
  wire n511bar;
  wire n512bar;
  wire n513bar;
  wire n514bar;
  wire n515bar;
  wire n516bar;
  wire n517bar;
  wire n518bar;
  wire n519bar;
  wire n520bar;
  wire n521bar;
  wire n522bar;
  wire n523bar;
  wire n524bar;
  wire n525bar;
  wire n526bar;
  wire n527bar;
  wire n528bar;
  wire n529bar;
  wire n530bar;
  wire n531bar;
  wire n532bar;
  wire n533bar;
  wire n534bar;
  wire n535bar;
  wire n536bar;
  wire n537bar;
  wire n538bar;
  wire n539bar;
  wire n540bar;
  wire n541bar;
  wire n542bar;
  wire n543bar;
  wire n544bar;
  wire n545bar;
  wire n546bar;
  wire n547bar;
  wire n548bar;
  wire n549bar;
  wire n550bar;
  wire n551bar;
  wire n552bar;
  wire n553bar;
  wire n554bar;
  wire n555bar;
  wire n556bar;
  wire n557bar;
  wire n558bar;
  wire n559bar;
  wire n560bar;
  wire n561bar;
  wire n562bar;
  wire n563bar;
  wire n564bar;
  wire n565bar;
  wire n566bar;
  wire n567bar;
  wire n568bar;
  wire n569bar;
  wire n570bar;
  wire n571bar;
  wire n572bar;
  wire n573bar;
  wire n574bar;
  wire n575bar;
  wire n576bar;
  wire n577bar;
  wire n578bar;
  wire n579bar;
  wire n580bar;
  wire n581bar;
  wire n582bar;
  wire n583bar;
  wire n584bar;
  wire n585bar;
  wire n586bar;
  wire n587bar;
  wire n588bar;
  wire n589bar;
  wire n590bar;
  wire n591bar;
  wire n592bar;
  wire n593bar;
  wire n594bar;
  wire n595bar;
  wire n596bar;
  wire n597bar;
  wire n598bar;
  wire n599bar;
  wire n600bar;
  wire n601bar;
  wire n602bar;
  wire n603bar;
  wire n604bar;
  wire n605bar;
  wire n606bar;
  wire n607bar;
  wire n608bar;
  wire n609bar;
  wire n610bar;
  wire n611bar;
  wire n612bar;
  wire n613bar;
  wire n614bar;
  wire n615bar;
  wire n616bar;
  wire n617bar;
  wire n618bar;
  wire n619bar;
  wire n620bar;
  wire n621bar;
  wire n622bar;
  wire n623bar;
  wire n624bar;
  wire n625bar;
  wire n626bar;
  wire n627bar;
  wire n628bar;
  wire n629bar;
  wire n630bar;
  wire n631bar;
  wire n632bar;
  wire n633bar;
  wire n634bar;
  wire n635bar;
  wire n636bar;
  wire n637bar;
  wire n638bar;
  wire n639bar;
  wire n640bar;
  wire n641bar;
  wire n642bar;
  wire n643bar;
  wire n644bar;
  wire n645bar;
  wire n646bar;
  wire n647bar;
  wire n648bar;
  wire n649bar;
  wire n650bar;
  wire n651bar;
  wire n652bar;
  wire n653bar;
  wire n654bar;
  wire n655bar;
  wire n656bar;
  wire n657bar;
  wire n658bar;
  wire n659bar;
  wire n660bar;
  wire n661bar;
  wire n662bar;
  wire n663bar;
  wire n664bar;
  wire n665bar;
  wire n666bar;
  wire n667bar;
  wire n668bar;
  wire n669bar;
  wire n670bar;
  wire n671bar;
  wire n672bar;
  wire n673bar;
  wire n674bar;
  wire n675bar;
  wire n676bar;
  wire n677bar;
  wire n678bar;
  wire n679bar;
  wire n680bar;
  wire n681bar;
  wire n682bar;
  wire n683bar;
  wire n684bar;
  wire n685bar;
  wire n686bar;
  wire n687bar;
  wire n688bar;
  wire n689bar;
  wire n690bar;
  wire n691bar;
  wire n692bar;
  wire n693bar;
  wire n694bar;
  wire n695bar;
  wire n696bar;
  wire n697bar;
  wire n698bar;
  wire n699bar;
  wire n700bar;
  wire n701bar;
  wire n702bar;
  wire n703bar;
  wire n704bar;
  wire n705bar;
  wire n706bar;
  wire n707bar;
  wire n708bar;
  wire n709bar;
  wire n710bar;
  wire n711bar;
  wire n712bar;
  wire n713bar;
  wire n714bar;
  wire n715bar;
  wire n716bar;
  wire n717bar;
  wire n718bar;
  wire n719bar;
  wire n720bar;
  wire n721bar;
  wire n722bar;
  wire n723bar;
  wire n724bar;
  wire n725bar;
  wire n726bar;
  wire n727bar;
  wire n728bar;
  wire n729bar;
  wire n730bar;
  wire n731bar;
  wire n732bar;
  wire n733bar;
  wire n734bar;
  wire n735bar;
  wire n736bar;
  wire n737bar;
  wire n738bar;
  wire n739bar;
  wire n740bar;
  wire n741bar;
  wire n742bar;
  wire n743bar;
  wire n744bar;
  wire n745bar;
  wire n746bar;
  wire n747bar;
  wire n748bar;
  wire n749bar;
  wire n750bar;
  wire n751bar;
  wire n752bar;
  wire n753bar;
  wire n754bar;
  wire n755bar;
  wire n756bar;
  wire n757bar;
  wire n758bar;
  wire n759bar;
  wire n760bar;
  wire n761bar;
  wire n762bar;
  wire n763bar;
  wire n764bar;
  wire n765bar;
  wire n766bar;
  wire n767bar;
  wire n768bar;
  wire n769bar;
  wire n770bar;
  wire n771bar;
  wire n772bar;
  wire n773bar;
  wire n774bar;
  wire n775bar;
  wire n776bar;
  wire n777bar;
  wire n778bar;
  wire n779bar;
  wire n780bar;
  wire n781bar;
  wire n782bar;
  wire n783bar;
  wire n784bar;
  wire n785bar;
  wire n786bar;
  wire n787bar;
  wire n788bar;
  wire n789bar;
  wire n790bar;
  wire n791bar;
  wire n792bar;
  wire n793bar;
  wire n794bar;
  wire n795bar;
  wire n796bar;
  wire n797bar;
  wire n798bar;
  wire n799bar;
  wire n800bar;
  wire n801bar;
  wire n802bar;
  wire n803bar;
  wire n804bar;
  wire n805bar;
  wire n806bar;
  wire n807bar;
  wire n808bar;
  wire n809bar;
  wire n810bar;
  wire n811bar;
  wire n812bar;
  wire n813bar;
  wire n814bar;
  wire n815bar;
  wire n816bar;
  wire n817bar;
  wire n818bar;
  wire n819bar;
  wire n820bar;
  wire n821bar;
  wire n822bar;
  wire n823bar;
  wire n824bar;
  wire n825bar;
  wire n826bar;
  wire n827bar;
  wire n828bar;
  wire n829bar;
  wire n830bar;
  wire n831bar;
  wire n832bar;
  wire n833bar;
  wire n834bar;
  wire n835bar;
  wire n836bar;
  wire n837bar;
  wire n838bar;
  wire n839bar;
  wire n840bar;
  wire n841bar;
  wire n842bar;
  wire n843bar;
  wire n844bar;
  wire n845bar;
  wire n846bar;
  wire n847bar;
  wire n848bar;
  wire n849bar;
  wire n850bar;
  wire n851bar;
  wire n852bar;
  wire n853bar;
  wire n854bar;
  wire n855bar;
  wire n856bar;
  wire n857bar;
  wire n858bar;
  wire n859bar;
  wire n860bar;
  wire n861bar;
  wire n862bar;
  wire n863bar;
  wire n864bar;
  wire n865bar;
  wire n866bar;
  wire n867bar;
  wire n868bar;
  wire n869bar;
  wire n870bar;
  wire n871bar;
  wire n872bar;
  wire n873bar;
  wire n874bar;
  wire n875bar;
  wire n876bar;
  wire n877bar;
  wire n878bar;
  wire n879bar;
  wire n880bar;
  wire n881bar;
  wire n882bar;
  wire n883bar;
  wire n884bar;
  wire n885bar;
  wire n886bar;
  wire n887bar;
  wire n888bar;
  wire n889bar;
  wire n890bar;
  wire n891bar;
  wire n892bar;
  wire n893bar;
  wire n894bar;
  wire n895bar;
  wire n896bar;
  wire n897bar;
  wire n898bar;
  wire n899bar;
  wire n900bar;
  wire n901bar;
  wire n902bar;
  wire n903bar;
  wire n904bar;
  wire n905bar;
  wire n906bar;
  wire n907bar;
  wire n908bar;
  wire n909bar;
  wire n910bar;
  wire n911bar;
  wire n912bar;
  wire n913bar;
  wire n914bar;
  wire n915bar;
  wire n916bar;
  wire n917bar;
  wire n918bar;
  wire n919bar;
  wire n920bar;
  wire n921bar;
  wire n922bar;
  wire n923bar;
  wire n924bar;
  wire n925bar;
  wire n926bar;
  wire n927bar;
  wire n928bar;
  wire n929bar;
  wire n930bar;
  wire n931bar;
  wire n932bar;
  wire n933bar;
  wire n934bar;
  wire n935bar;
  wire n936bar;
  wire n937bar;
  wire n938bar;
  wire n939bar;
  wire n940bar;
  wire n941bar;
  wire n942bar;
  wire n943bar;
  wire n944bar;
  wire n945bar;
  wire n946bar;
  wire n947bar;
  wire n948bar;
  wire n949bar;
  wire n950bar;
  wire n951bar;
  wire n952bar;
  wire n953bar;
  wire n954bar;
  wire n955bar;
  wire n956bar;
  wire n957bar;
  wire n958bar;
  wire n959bar;
  wire n960bar;
  wire n961bar;
  wire n962bar;
  wire n963bar;
  wire n964bar;
  wire n965bar;
  wire n966bar;
  wire n967bar;
  wire n968bar;
  wire n969bar;
  wire n970bar;
  wire n971bar;
  wire n972bar;
//wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];
  assign in_81bar = inbar[81];
  assign in_80bar = inbar[80];
  assign in_79bar = inbar[79];
  assign in_78bar = inbar[78];
  assign in_77bar = inbar[77];
  assign in_76bar = inbar[76];
  assign in_75bar = inbar[75];
  assign in_74bar = inbar[74];
  assign in_73bar = inbar[73];
  assign in_72bar = inbar[72];
  assign in_71bar = inbar[71];
  assign in_70bar = inbar[70];
  assign in_69bar = inbar[69];
  assign in_68bar = inbar[68];
  assign in_67bar = inbar[67];
  assign in_66bar = inbar[66];
  assign in_65bar = inbar[65];
  assign in_64bar = inbar[64];
  assign in_63bar = inbar[63];
  assign in_62bar = inbar[62];
  assign in_61bar = inbar[61];
  assign in_60bar = inbar[60];
  assign in_59bar = inbar[59];
  assign in_58bar = inbar[58];
  assign in_57bar = inbar[57];
  assign in_56bar = inbar[56];
  assign in_55bar = inbar[55];
  assign in_54bar = inbar[54];
  assign in_53bar = inbar[53];
  assign in_52bar = inbar[52];
  assign in_51bar = inbar[51];
  assign in_50bar = inbar[50];
  assign in_49bar = inbar[49];
  assign in_48bar = inbar[48];
  assign in_47bar = inbar[47];
  assign in_46bar = inbar[46];
  assign in_45bar = inbar[45];
  assign in_44bar = inbar[44];
  assign in_43bar = inbar[43];
  assign in_42bar = inbar[42];
  assign in_41bar = inbar[41];
  assign in_40bar = inbar[40];
  assign in_39bar = inbar[39];
  assign in_38bar = inbar[38];
  assign in_37bar = inbar[37];
  assign in_36bar = inbar[36];
  assign in_35bar = inbar[35];
  assign in_34bar = inbar[34];
  assign in_33bar = inbar[33];
  assign in_32bar = inbar[32];
  assign in_31bar = inbar[31];
  assign in_30bar = inbar[30];
  assign in_29bar = inbar[29];
  assign in_28bar = inbar[28];
  assign in_27bar = inbar[27];
  assign in_26bar = inbar[26];
  assign in_25bar = inbar[25];
  assign in_24bar = inbar[24];
  assign in_23bar = inbar[23];
  assign in_22bar = inbar[22];
  assign in_21bar = inbar[21];
  assign in_20bar = inbar[20];
  assign in_19bar = inbar[19];
  assign in_18bar = inbar[18];
  assign in_17bar = inbar[17];
  assign in_16bar = inbar[16];
  assign in_15bar = inbar[15];
  assign in_14bar = inbar[14];
  assign in_13bar = inbar[13];
  assign in_12bar = inbar[12];
  assign in_11bar = inbar[11];
  assign in_10bar = inbar[10];
  assign in_9bar = inbar[9];
  assign in_8bar = inbar[8];
  assign in_7bar = inbar[7];
  assign in_6bar = inbar[6];
  assign in_5bar = inbar[5];
  assign in_4bar = inbar[4];
  assign in_3bar = inbar[3];
  assign in_2bar = inbar[2];
  assign in_1bar = inbar[1];
  assign in_0bar = inbar[0];
//assign_done

  OR2_X1 U1 ( .A1(n972), .A2(n971), .ZN(out[7]) );
  AND2_X1 U1bar ( .A1(n972bar), .A2(n971bar), .ZN(outbar[7]) );
  OR2_X1 U2 ( .A1(n970), .A2(n969), .ZN(n971) );
  AND2_X1 U2bar ( .A1(n970bar), .A2(n969bar), .ZN(n971bar) );
  OR2_X1 U3 ( .A1(n968), .A2(n967), .ZN(n969) );
  AND2_X1 U3bar ( .A1(n968bar), .A2(n967bar), .ZN(n969bar) );
  OR2_X1 U4 ( .A1(n966), .A2(n965), .ZN(n967) );
  AND2_X1 U4bar ( .A1(n966bar), .A2(n965bar), .ZN(n967bar) );
  OR2_X1 U5 ( .A1(n964), .A2(n963), .ZN(n968) );
  AND2_X1 U5bar ( .A1(n964bar), .A2(n963bar), .ZN(n968bar) );
  OR2_X1 U6 ( .A1(in[116]), .A2(n962), .ZN(n963) );
  AND2_X1 U6bar ( .A1(inbar[116]), .A2(n962bar), .ZN(n963bar) );
  OR2_X1 U7 ( .A1(n961), .A2(n960), .ZN(n970) );
  AND2_X1 U7bar ( .A1(n961bar), .A2(n960bar), .ZN(n970bar) );
  OR2_X1 U8 ( .A1(in[150]), .A2(in[127]), .ZN(n960) );
  AND2_X1 U8bar ( .A1(inbar[150]), .A2(inbar[127]), .ZN(n960bar) );
  OR2_X1 U9 ( .A1(in[160]), .A2(n959), .ZN(n961) );
  AND2_X1 U9bar ( .A1(inbar[160]), .A2(n959bar), .ZN(n961bar) );
  OR2_X1 U10 ( .A1(in[252]), .A2(in[168]), .ZN(n959) );
  AND2_X1 U10bar ( .A1(inbar[252]), .A2(inbar[168]), .ZN(n959bar) );
  OR2_X1 U11 ( .A1(n958), .A2(n957), .ZN(n972) );
  AND2_X1 U11bar ( .A1(n958bar), .A2(n957bar), .ZN(n972bar) );
  OR2_X1 U12 ( .A1(n956), .A2(n955), .ZN(n957) );
  AND2_X1 U12bar ( .A1(n956bar), .A2(n955bar), .ZN(n957bar) );
  OR2_X1 U13 ( .A1(in_17), .A2(in[96]), .ZN(n955) );
  AND2_X1 U13bar ( .A1(in_17bar), .A2(inbar[96]), .ZN(n955bar) );
  OR2_X1 U14 ( .A1(in_23), .A2(n954), .ZN(n956) );
  AND2_X1 U14bar ( .A1(in_23bar), .A2(n954bar), .ZN(n956bar) );
  OR2_X1 U15 ( .A1(in_31), .A2(in_26), .ZN(n954) );
  AND2_X1 U15bar ( .A1(in_31bar), .A2(in_26bar), .ZN(n954bar) );
  OR2_X1 U16 ( .A1(n953), .A2(n952), .ZN(n958) );
  AND2_X1 U16bar ( .A1(n953bar), .A2(n952bar), .ZN(n958bar) );
  OR2_X1 U17 ( .A1(in_58), .A2(in_4), .ZN(n952) );
  AND2_X1 U17bar ( .A1(in_58bar), .A2(in_4bar), .ZN(n952bar) );
  OR2_X1 U18 ( .A1(in_59), .A2(n951), .ZN(n953) );
  AND2_X1 U18bar ( .A1(in_59bar), .A2(n951bar), .ZN(n953bar) );
  OR2_X1 U19 ( .A1(in_71), .A2(in_62), .ZN(n951) );
  AND2_X1 U19bar ( .A1(in_71bar), .A2(in_62bar), .ZN(n951bar) );
  OR2_X1 U20 ( .A1(n950), .A2(n949), .ZN(out[6]) );
  AND2_X1 U20bar ( .A1(n950bar), .A2(n949bar), .ZN(outbar[6]) );
  OR2_X1 U21 ( .A1(n948), .A2(n947), .ZN(n949) );
  AND2_X1 U21bar ( .A1(n948bar), .A2(n947bar), .ZN(n949bar) );
  OR2_X1 U22 ( .A1(n946), .A2(n945), .ZN(n947) );
  AND2_X1 U22bar ( .A1(n946bar), .A2(n945bar), .ZN(n947bar) );
  OR2_X1 U23 ( .A1(n944), .A2(n943), .ZN(n945) );
  AND2_X1 U23bar ( .A1(n944bar), .A2(n943bar), .ZN(n945bar) );
  OR2_X1 U24 ( .A1(n942), .A2(n941), .ZN(n946) );
  AND2_X1 U24bar ( .A1(n942bar), .A2(n941bar), .ZN(n946bar) );
  OR2_X1 U25 ( .A1(in[101]), .A2(n940), .ZN(n941) );
  AND2_X1 U25bar ( .A1(inbar[101]), .A2(n940bar), .ZN(n941bar) );
  OR2_X1 U26 ( .A1(n939), .A2(n938), .ZN(n948) );
  AND2_X1 U26bar ( .A1(n939bar), .A2(n938bar), .ZN(n948bar) );
  OR2_X1 U27 ( .A1(in[114]), .A2(in[104]), .ZN(n938) );
  AND2_X1 U27bar ( .A1(inbar[114]), .A2(inbar[104]), .ZN(n938bar) );
  OR2_X1 U28 ( .A1(in[128]), .A2(n937), .ZN(n939) );
  AND2_X1 U28bar ( .A1(inbar[128]), .A2(n937bar), .ZN(n939bar) );
  OR2_X1 U29 ( .A1(in[136]), .A2(in[134]), .ZN(n937) );
  AND2_X1 U29bar ( .A1(inbar[136]), .A2(inbar[134]), .ZN(n937bar) );
  OR2_X1 U30 ( .A1(n936), .A2(n935), .ZN(n950) );
  AND2_X1 U30bar ( .A1(n936bar), .A2(n935bar), .ZN(n950bar) );
  OR2_X1 U31 ( .A1(n934), .A2(n933), .ZN(n935) );
  AND2_X1 U31bar ( .A1(n934bar), .A2(n933bar), .ZN(n935bar) );
  OR2_X1 U32 ( .A1(in[177]), .A2(in[164]), .ZN(n933) );
  AND2_X1 U32bar ( .A1(inbar[177]), .A2(inbar[164]), .ZN(n933bar) );
  OR2_X1 U33 ( .A1(in[212]), .A2(n932), .ZN(n934) );
  AND2_X1 U33bar ( .A1(inbar[212]), .A2(n932bar), .ZN(n934bar) );
  OR2_X1 U34 ( .A1(in[248]), .A2(in[221]), .ZN(n932) );
  AND2_X1 U34bar ( .A1(inbar[248]), .A2(inbar[221]), .ZN(n932bar) );
  OR2_X1 U35 ( .A1(n931), .A2(n930), .ZN(n936) );
  AND2_X1 U35bar ( .A1(n931bar), .A2(n930bar), .ZN(n936bar) );
  OR2_X1 U36 ( .A1(in_18), .A2(in[93]), .ZN(n930) );
  AND2_X1 U36bar ( .A1(in_18bar), .A2(inbar[93]), .ZN(n930bar) );
  OR2_X1 U37 ( .A1(in_31), .A2(n929), .ZN(n931) );
  AND2_X1 U37bar ( .A1(in_31bar), .A2(n929bar), .ZN(n931bar) );
  OR2_X1 U38 ( .A1(in_7), .A2(in_39), .ZN(n929) );
  AND2_X1 U38bar ( .A1(in_7bar), .A2(in_39bar), .ZN(n929bar) );
  OR2_X1 U39 ( .A1(n928), .A2(n927), .ZN(out[5]) );
  AND2_X1 U39bar ( .A1(n928bar), .A2(n927bar), .ZN(outbar[5]) );
  OR2_X1 U40 ( .A1(n926), .A2(n925), .ZN(n927) );
  AND2_X1 U40bar ( .A1(n926bar), .A2(n925bar), .ZN(n927bar) );
  OR2_X1 U41 ( .A1(n924), .A2(n923), .ZN(n925) );
  AND2_X1 U41bar ( .A1(n924bar), .A2(n923bar), .ZN(n925bar) );
  OR2_X1 U42 ( .A1(n922), .A2(n921), .ZN(n923) );
  AND2_X1 U42bar ( .A1(n922bar), .A2(n921bar), .ZN(n923bar) );
  OR2_X1 U43 ( .A1(n940), .A2(n920), .ZN(n924) );
  AND2_X1 U43bar ( .A1(n940bar), .A2(n920bar), .ZN(n924bar) );
  OR2_X1 U44 ( .A1(in[111]), .A2(n919), .ZN(n920) );
  AND2_X1 U44bar ( .A1(inbar[111]), .A2(n919bar), .ZN(n920bar) );
  OR2_X1 U45 ( .A1(n918), .A2(n917), .ZN(n940) );
  AND2_X1 U45bar ( .A1(n918bar), .A2(n917bar), .ZN(n940bar) );
  OR2_X1 U46 ( .A1(n916), .A2(n915), .ZN(n917) );
  AND2_X1 U46bar ( .A1(n916bar), .A2(n915bar), .ZN(n917bar) );
  OR2_X1 U47 ( .A1(n914), .A2(n913), .ZN(n915) );
  AND2_X1 U47bar ( .A1(n914bar), .A2(n913bar), .ZN(n915bar) );
  OR2_X1 U48 ( .A1(in[140]), .A2(in[131]), .ZN(n913) );
  AND2_X1 U48bar ( .A1(inbar[140]), .A2(inbar[131]), .ZN(n913bar) );
  OR2_X1 U49 ( .A1(in[160]), .A2(in[144]), .ZN(n914) );
  AND2_X1 U49bar ( .A1(inbar[160]), .A2(inbar[144]), .ZN(n914bar) );
  OR2_X1 U50 ( .A1(n912), .A2(n911), .ZN(n916) );
  AND2_X1 U50bar ( .A1(n912bar), .A2(n911bar), .ZN(n916bar) );
  OR2_X1 U51 ( .A1(in[179]), .A2(in[174]), .ZN(n911) );
  AND2_X1 U51bar ( .A1(inbar[179]), .A2(inbar[174]), .ZN(n911bar) );
  OR2_X1 U52 ( .A1(in[188]), .A2(in[184]), .ZN(n912) );
  AND2_X1 U52bar ( .A1(inbar[188]), .A2(inbar[184]), .ZN(n912bar) );
  OR2_X1 U53 ( .A1(n910), .A2(n909), .ZN(n918) );
  AND2_X1 U53bar ( .A1(n910bar), .A2(n909bar), .ZN(n918bar) );
  OR2_X1 U54 ( .A1(n908), .A2(n907), .ZN(n909) );
  AND2_X1 U54bar ( .A1(n908bar), .A2(n907bar), .ZN(n909bar) );
  OR2_X1 U55 ( .A1(in[216]), .A2(in[200]), .ZN(n907) );
  AND2_X1 U55bar ( .A1(inbar[216]), .A2(inbar[200]), .ZN(n907bar) );
  OR2_X1 U56 ( .A1(in[228]), .A2(in[224]), .ZN(n908) );
  AND2_X1 U56bar ( .A1(inbar[228]), .A2(inbar[224]), .ZN(n908bar) );
  OR2_X1 U57 ( .A1(n906), .A2(n905), .ZN(n910) );
  AND2_X1 U57bar ( .A1(n906bar), .A2(n905bar), .ZN(n910bar) );
  OR2_X1 U58 ( .A1(in[247]), .A2(in[235]), .ZN(n905) );
  AND2_X1 U58bar ( .A1(inbar[247]), .A2(inbar[235]), .ZN(n905bar) );
  OR2_X1 U59 ( .A1(in_42), .A2(in[83]), .ZN(n906) );
  AND2_X1 U59bar ( .A1(in_42bar), .A2(inbar[83]), .ZN(n906bar) );
  OR2_X1 U60 ( .A1(n904), .A2(n903), .ZN(n926) );
  AND2_X1 U60bar ( .A1(n904bar), .A2(n903bar), .ZN(n926bar) );
  OR2_X1 U61 ( .A1(in[166]), .A2(in[123]), .ZN(n903) );
  AND2_X1 U61bar ( .A1(inbar[166]), .A2(inbar[123]), .ZN(n903bar) );
  OR2_X1 U62 ( .A1(in[170]), .A2(n902), .ZN(n904) );
  AND2_X1 U62bar ( .A1(inbar[170]), .A2(n902bar), .ZN(n904bar) );
  OR2_X1 U63 ( .A1(in[194]), .A2(in[183]), .ZN(n902) );
  AND2_X1 U63bar ( .A1(inbar[194]), .A2(inbar[183]), .ZN(n902bar) );
  OR2_X1 U64 ( .A1(n901), .A2(n900), .ZN(n928) );
  AND2_X1 U64bar ( .A1(n901bar), .A2(n900bar), .ZN(n928bar) );
  OR2_X1 U65 ( .A1(n899), .A2(n898), .ZN(n900) );
  AND2_X1 U65bar ( .A1(n899bar), .A2(n898bar), .ZN(n900bar) );
  OR2_X1 U66 ( .A1(in[241]), .A2(in[238]), .ZN(n898) );
  AND2_X1 U66bar ( .A1(inbar[241]), .A2(inbar[238]), .ZN(n898bar) );
  OR2_X1 U67 ( .A1(in[250]), .A2(n897), .ZN(n899) );
  AND2_X1 U67bar ( .A1(inbar[250]), .A2(n897bar), .ZN(n899bar) );
  OR2_X1 U68 ( .A1(in_24), .A2(in[84]), .ZN(n897) );
  AND2_X1 U68bar ( .A1(in_24bar), .A2(inbar[84]), .ZN(n897bar) );
  OR2_X1 U69 ( .A1(n896), .A2(n895), .ZN(n901) );
  AND2_X1 U69bar ( .A1(n896bar), .A2(n895bar), .ZN(n901bar) );
  OR2_X1 U70 ( .A1(in_41), .A2(in_29), .ZN(n895) );
  AND2_X1 U70bar ( .A1(in_41bar), .A2(in_29bar), .ZN(n895bar) );
  OR2_X1 U71 ( .A1(in_66), .A2(n894), .ZN(n896) );
  AND2_X1 U71bar ( .A1(in_66bar), .A2(n894bar), .ZN(n896bar) );
  OR2_X1 U72 ( .A1(in_76), .A2(in_71), .ZN(n894) );
  AND2_X1 U72bar ( .A1(in_76bar), .A2(in_71bar), .ZN(n894bar) );
  OR2_X1 U73 ( .A1(n893), .A2(n892), .ZN(out[4]) );
  AND2_X1 U73bar ( .A1(n893bar), .A2(n892bar), .ZN(outbar[4]) );
  OR2_X1 U74 ( .A1(n891), .A2(n890), .ZN(n892) );
  AND2_X1 U74bar ( .A1(n891bar), .A2(n890bar), .ZN(n892bar) );
  OR2_X1 U75 ( .A1(n889), .A2(n888), .ZN(n890) );
  AND2_X1 U75bar ( .A1(n889bar), .A2(n888bar), .ZN(n890bar) );
  OR2_X1 U76 ( .A1(n922), .A2(n887), .ZN(n888) );
  AND2_X1 U76bar ( .A1(n922bar), .A2(n887bar), .ZN(n888bar) );
  OR2_X1 U77 ( .A1(n886), .A2(n885), .ZN(n922) );
  AND2_X1 U77bar ( .A1(n886bar), .A2(n885bar), .ZN(n922bar) );
  OR2_X1 U78 ( .A1(n884), .A2(n883), .ZN(n885) );
  AND2_X1 U78bar ( .A1(n884bar), .A2(n883bar), .ZN(n885bar) );
  OR2_X1 U79 ( .A1(n882), .A2(n881), .ZN(n883) );
  AND2_X1 U79bar ( .A1(n882bar), .A2(n881bar), .ZN(n883bar) );
  OR2_X1 U80 ( .A1(in[118]), .A2(in[109]), .ZN(n881) );
  AND2_X1 U80bar ( .A1(inbar[118]), .A2(inbar[109]), .ZN(n881bar) );
  OR2_X1 U81 ( .A1(in[139]), .A2(in[120]), .ZN(n882) );
  AND2_X1 U81bar ( .A1(inbar[139]), .A2(inbar[120]), .ZN(n882bar) );
  OR2_X1 U82 ( .A1(n880), .A2(n879), .ZN(n884) );
  AND2_X1 U82bar ( .A1(n880bar), .A2(n879bar), .ZN(n884bar) );
  OR2_X1 U83 ( .A1(in[198]), .A2(in[154]), .ZN(n879) );
  AND2_X1 U83bar ( .A1(inbar[198]), .A2(inbar[154]), .ZN(n879bar) );
  OR2_X1 U84 ( .A1(in[210]), .A2(in[205]), .ZN(n880) );
  AND2_X1 U84bar ( .A1(inbar[210]), .A2(inbar[205]), .ZN(n880bar) );
  OR2_X1 U85 ( .A1(n878), .A2(n877), .ZN(n886) );
  AND2_X1 U85bar ( .A1(n878bar), .A2(n877bar), .ZN(n886bar) );
  OR2_X1 U86 ( .A1(n876), .A2(n875), .ZN(n877) );
  AND2_X1 U86bar ( .A1(n876bar), .A2(n875bar), .ZN(n877bar) );
  OR2_X1 U87 ( .A1(in[219]), .A2(in[217]), .ZN(n875) );
  AND2_X1 U87bar ( .A1(inbar[219]), .A2(inbar[217]), .ZN(n875bar) );
  OR2_X1 U88 ( .A1(in[86]), .A2(in[252]), .ZN(n876) );
  AND2_X1 U88bar ( .A1(inbar[86]), .A2(inbar[252]), .ZN(n876bar) );
  OR2_X1 U89 ( .A1(n874), .A2(n873), .ZN(n878) );
  AND2_X1 U89bar ( .A1(n874bar), .A2(n873bar), .ZN(n878bar) );
  OR2_X1 U90 ( .A1(in_40), .A2(in[91]), .ZN(n873) );
  AND2_X1 U90bar ( .A1(in_40bar), .A2(inbar[91]), .ZN(n873bar) );
  OR2_X1 U91 ( .A1(in_8), .A2(in_46), .ZN(n874) );
  AND2_X1 U91bar ( .A1(in_8bar), .A2(in_46bar), .ZN(n874bar) );
  OR2_X1 U92 ( .A1(n872), .A2(n871), .ZN(n889) );
  AND2_X1 U92bar ( .A1(n872bar), .A2(n871bar), .ZN(n889bar) );
  OR2_X1 U93 ( .A1(in[117]), .A2(n943), .ZN(n871) );
  AND2_X1 U93bar ( .A1(inbar[117]), .A2(n943bar), .ZN(n871bar) );
  OR2_X1 U94 ( .A1(n870), .A2(n869), .ZN(n943) );
  AND2_X1 U94bar ( .A1(n870bar), .A2(n869bar), .ZN(n943bar) );
  OR2_X1 U95 ( .A1(n868), .A2(n867), .ZN(n869) );
  AND2_X1 U95bar ( .A1(n868bar), .A2(n867bar), .ZN(n869bar) );
  OR2_X1 U96 ( .A1(n866), .A2(n865), .ZN(n867) );
  AND2_X1 U96bar ( .A1(n866bar), .A2(n865bar), .ZN(n867bar) );
  OR2_X1 U97 ( .A1(n864), .A2(n863), .ZN(n865) );
  AND2_X1 U97bar ( .A1(n864bar), .A2(n863bar), .ZN(n865bar) );
  OR2_X1 U98 ( .A1(in[108]), .A2(n919), .ZN(n866) );
  AND2_X1 U98bar ( .A1(inbar[108]), .A2(n919bar), .ZN(n866bar) );
  OR2_X1 U99 ( .A1(n862), .A2(n861), .ZN(n919) );
  AND2_X1 U99bar ( .A1(n862bar), .A2(n861bar), .ZN(n919bar) );
  OR2_X1 U100 ( .A1(n860), .A2(n859), .ZN(n861) );
  AND2_X1 U100bar ( .A1(n860bar), .A2(n859bar), .ZN(n861bar) );
  OR2_X1 U101 ( .A1(n858), .A2(n857), .ZN(n859) );
  AND2_X1 U101bar ( .A1(n858bar), .A2(n857bar), .ZN(n859bar) );
  OR2_X1 U102 ( .A1(in[119]), .A2(in[105]), .ZN(n857) );
  AND2_X1 U102bar ( .A1(inbar[119]), .A2(inbar[105]), .ZN(n857bar) );
  OR2_X1 U103 ( .A1(in[186]), .A2(in[175]), .ZN(n858) );
  AND2_X1 U103bar ( .A1(inbar[186]), .A2(inbar[175]), .ZN(n858bar) );
  OR2_X1 U104 ( .A1(n856), .A2(n855), .ZN(n860) );
  AND2_X1 U104bar ( .A1(n856bar), .A2(n855bar), .ZN(n860bar) );
  OR2_X1 U105 ( .A1(in[202]), .A2(in[193]), .ZN(n855) );
  AND2_X1 U105bar ( .A1(inbar[202]), .A2(inbar[193]), .ZN(n855bar) );
  OR2_X1 U106 ( .A1(in[225]), .A2(in[208]), .ZN(n856) );
  AND2_X1 U106bar ( .A1(inbar[225]), .A2(inbar[208]), .ZN(n856bar) );
  OR2_X1 U107 ( .A1(n854), .A2(n853), .ZN(n862) );
  AND2_X1 U107bar ( .A1(n854bar), .A2(n853bar), .ZN(n862bar) );
  OR2_X1 U108 ( .A1(n852), .A2(n851), .ZN(n853) );
  AND2_X1 U108bar ( .A1(n852bar), .A2(n851bar), .ZN(n853bar) );
  OR2_X1 U109 ( .A1(in_1), .A2(in[85]), .ZN(n851) );
  AND2_X1 U109bar ( .A1(in_1bar), .A2(inbar[85]), .ZN(n851bar) );
  OR2_X1 U110 ( .A1(in_23), .A2(in_19), .ZN(n852) );
  AND2_X1 U110bar ( .A1(in_23bar), .A2(in_19bar), .ZN(n852bar) );
  OR2_X1 U111 ( .A1(n850), .A2(n849), .ZN(n854) );
  AND2_X1 U111bar ( .A1(n850bar), .A2(n849bar), .ZN(n854bar) );
  OR2_X1 U112 ( .A1(in_43), .A2(in_33), .ZN(n849) );
  AND2_X1 U112bar ( .A1(in_43bar), .A2(in_33bar), .ZN(n849bar) );
  OR2_X1 U113 ( .A1(in_63), .A2(in_44), .ZN(n850) );
  AND2_X1 U113bar ( .A1(in_63bar), .A2(in_44bar), .ZN(n850bar) );
  OR2_X1 U114 ( .A1(n848), .A2(n847), .ZN(n868) );
  AND2_X1 U114bar ( .A1(n848bar), .A2(n847bar), .ZN(n868bar) );
  OR2_X1 U115 ( .A1(in[141]), .A2(in[112]), .ZN(n847) );
  AND2_X1 U115bar ( .A1(inbar[141]), .A2(inbar[112]), .ZN(n847bar) );
  OR2_X1 U116 ( .A1(in[147]), .A2(n846), .ZN(n848) );
  AND2_X1 U116bar ( .A1(inbar[147]), .A2(n846bar), .ZN(n848bar) );
  OR2_X1 U117 ( .A1(in[181]), .A2(in[167]), .ZN(n846) );
  AND2_X1 U117bar ( .A1(inbar[181]), .A2(inbar[167]), .ZN(n846bar) );
  OR2_X1 U118 ( .A1(n845), .A2(n844), .ZN(n870) );
  AND2_X1 U118bar ( .A1(n845bar), .A2(n844bar), .ZN(n870bar) );
  OR2_X1 U119 ( .A1(n843), .A2(n842), .ZN(n844) );
  AND2_X1 U119bar ( .A1(n843bar), .A2(n842bar), .ZN(n844bar) );
  OR2_X1 U120 ( .A1(in[229]), .A2(in[201]), .ZN(n842) );
  AND2_X1 U120bar ( .A1(inbar[229]), .A2(inbar[201]), .ZN(n842bar) );
  OR2_X1 U121 ( .A1(in[237]), .A2(n841), .ZN(n843) );
  AND2_X1 U121bar ( .A1(inbar[237]), .A2(n841bar), .ZN(n843bar) );
  OR2_X1 U122 ( .A1(in[94]), .A2(in[253]), .ZN(n841) );
  AND2_X1 U122bar ( .A1(inbar[94]), .A2(inbar[253]), .ZN(n841bar) );
  OR2_X1 U123 ( .A1(n840), .A2(n839), .ZN(n845) );
  AND2_X1 U123bar ( .A1(n840bar), .A2(n839bar), .ZN(n845bar) );
  OR2_X1 U124 ( .A1(in_21), .A2(in[96]), .ZN(n839) );
  AND2_X1 U124bar ( .A1(in_21bar), .A2(inbar[96]), .ZN(n839bar) );
  OR2_X1 U125 ( .A1(in_25), .A2(n838), .ZN(n840) );
  AND2_X1 U125bar ( .A1(in_25bar), .A2(n838bar), .ZN(n840bar) );
  OR2_X1 U126 ( .A1(in_81), .A2(in_45), .ZN(n838) );
  AND2_X1 U126bar ( .A1(in_81bar), .A2(in_45bar), .ZN(n838bar) );
  OR2_X1 U127 ( .A1(n837), .A2(n836), .ZN(n891) );
  AND2_X1 U127bar ( .A1(n837bar), .A2(n836bar), .ZN(n891bar) );
  OR2_X1 U128 ( .A1(in[142]), .A2(in[124]), .ZN(n836) );
  AND2_X1 U128bar ( .A1(inbar[142]), .A2(inbar[124]), .ZN(n836bar) );
  OR2_X1 U129 ( .A1(in[150]), .A2(n835), .ZN(n837) );
  AND2_X1 U129bar ( .A1(inbar[150]), .A2(n835bar), .ZN(n837bar) );
  OR2_X1 U130 ( .A1(in[172]), .A2(in[155]), .ZN(n835) );
  AND2_X1 U130bar ( .A1(inbar[172]), .A2(inbar[155]), .ZN(n835bar) );
  OR2_X1 U131 ( .A1(n834), .A2(n833), .ZN(n893) );
  AND2_X1 U131bar ( .A1(n834bar), .A2(n833bar), .ZN(n893bar) );
  OR2_X1 U132 ( .A1(n832), .A2(n831), .ZN(n833) );
  AND2_X1 U132bar ( .A1(n832bar), .A2(n831bar), .ZN(n833bar) );
  OR2_X1 U133 ( .A1(in[196]), .A2(in[173]), .ZN(n831) );
  AND2_X1 U133bar ( .A1(inbar[196]), .A2(inbar[173]), .ZN(n831bar) );
  OR2_X1 U134 ( .A1(in[222]), .A2(n830), .ZN(n832) );
  AND2_X1 U134bar ( .A1(inbar[222]), .A2(n830bar), .ZN(n832bar) );
  OR2_X1 U135 ( .A1(in[227]), .A2(in[226]), .ZN(n830) );
  AND2_X1 U135bar ( .A1(inbar[227]), .A2(inbar[226]), .ZN(n830bar) );
  OR2_X1 U136 ( .A1(n829), .A2(n828), .ZN(n834) );
  AND2_X1 U136bar ( .A1(n829bar), .A2(n828bar), .ZN(n834bar) );
  OR2_X1 U137 ( .A1(in[249]), .A2(in[231]), .ZN(n828) );
  AND2_X1 U137bar ( .A1(inbar[249]), .A2(inbar[231]), .ZN(n828bar) );
  OR2_X1 U138 ( .A1(in_28), .A2(n827), .ZN(n829) );
  AND2_X1 U138bar ( .A1(in_28bar), .A2(n827bar), .ZN(n829bar) );
  OR2_X1 U139 ( .A1(in_52), .A2(in_47), .ZN(n827) );
  AND2_X1 U139bar ( .A1(in_52bar), .A2(in_47bar), .ZN(n827bar) );
  OR2_X1 U140 ( .A1(n826), .A2(n825), .ZN(out[3]) );
  AND2_X1 U140bar ( .A1(n826bar), .A2(n825bar), .ZN(outbar[3]) );
  OR2_X1 U141 ( .A1(n824), .A2(n823), .ZN(n825) );
  AND2_X1 U141bar ( .A1(n824bar), .A2(n823bar), .ZN(n825bar) );
  OR2_X1 U142 ( .A1(n822), .A2(n821), .ZN(n823) );
  AND2_X1 U142bar ( .A1(n822bar), .A2(n821bar), .ZN(n823bar) );
  OR2_X1 U143 ( .A1(n820), .A2(n819), .ZN(n821) );
  AND2_X1 U143bar ( .A1(n820bar), .A2(n819bar), .ZN(n821bar) );
  OR2_X1 U144 ( .A1(n964), .A2(n818), .ZN(n822) );
  AND2_X1 U144bar ( .A1(n964bar), .A2(n818bar), .ZN(n822bar) );
  OR2_X1 U145 ( .A1(in[118]), .A2(n817), .ZN(n818) );
  AND2_X1 U145bar ( .A1(inbar[118]), .A2(n817bar), .ZN(n818bar) );
  OR2_X1 U146 ( .A1(n816), .A2(n815), .ZN(n964) );
  AND2_X1 U146bar ( .A1(n816bar), .A2(n815bar), .ZN(n964bar) );
  OR2_X1 U147 ( .A1(n814), .A2(n813), .ZN(n815) );
  AND2_X1 U147bar ( .A1(n814bar), .A2(n813bar), .ZN(n815bar) );
  OR2_X1 U148 ( .A1(n812), .A2(n811), .ZN(n813) );
  AND2_X1 U148bar ( .A1(n812bar), .A2(n811bar), .ZN(n813bar) );
  OR2_X1 U149 ( .A1(in[122]), .A2(in[111]), .ZN(n811) );
  AND2_X1 U149bar ( .A1(inbar[122]), .A2(inbar[111]), .ZN(n811bar) );
  OR2_X1 U150 ( .A1(in[154]), .A2(in[151]), .ZN(n812) );
  AND2_X1 U150bar ( .A1(inbar[154]), .A2(inbar[151]), .ZN(n812bar) );
  OR2_X1 U151 ( .A1(n810), .A2(n809), .ZN(n814) );
  AND2_X1 U151bar ( .A1(n810bar), .A2(n809bar), .ZN(n814bar) );
  OR2_X1 U152 ( .A1(in[187]), .A2(in[177]), .ZN(n809) );
  AND2_X1 U152bar ( .A1(inbar[187]), .A2(inbar[177]), .ZN(n809bar) );
  OR2_X1 U153 ( .A1(in[200]), .A2(in[192]), .ZN(n810) );
  AND2_X1 U153bar ( .A1(inbar[200]), .A2(inbar[192]), .ZN(n810bar) );
  OR2_X1 U154 ( .A1(n808), .A2(n807), .ZN(n816) );
  AND2_X1 U154bar ( .A1(n808bar), .A2(n807bar), .ZN(n816bar) );
  OR2_X1 U155 ( .A1(n806), .A2(n805), .ZN(n807) );
  AND2_X1 U155bar ( .A1(n806bar), .A2(n805bar), .ZN(n807bar) );
  OR2_X1 U156 ( .A1(in[225]), .A2(in[207]), .ZN(n805) );
  AND2_X1 U156bar ( .A1(inbar[225]), .A2(inbar[207]), .ZN(n805bar) );
  OR2_X1 U157 ( .A1(in[98]), .A2(in[226]), .ZN(n806) );
  AND2_X1 U157bar ( .A1(inbar[98]), .A2(inbar[226]), .ZN(n806bar) );
  OR2_X1 U158 ( .A1(n804), .A2(n803), .ZN(n808) );
  AND2_X1 U158bar ( .A1(n804bar), .A2(n803bar), .ZN(n808bar) );
  OR2_X1 U159 ( .A1(in_20), .A2(in_16), .ZN(n803) );
  AND2_X1 U159bar ( .A1(in_20bar), .A2(in_16bar), .ZN(n803bar) );
  OR2_X1 U160 ( .A1(in_55), .A2(in_45), .ZN(n804) );
  AND2_X1 U160bar ( .A1(in_55bar), .A2(in_45bar), .ZN(n804bar) );
  OR2_X1 U161 ( .A1(n802), .A2(n801), .ZN(n824) );
  AND2_X1 U161bar ( .A1(n802bar), .A2(n801bar), .ZN(n824bar) );
  OR2_X1 U162 ( .A1(in[162]), .A2(in[149]), .ZN(n801) );
  AND2_X1 U162bar ( .A1(inbar[162]), .A2(inbar[149]), .ZN(n801bar) );
  OR2_X1 U163 ( .A1(in[163]), .A2(n800), .ZN(n802) );
  AND2_X1 U163bar ( .A1(inbar[163]), .A2(n800bar), .ZN(n802bar) );
  OR2_X1 U164 ( .A1(in[191]), .A2(in[189]), .ZN(n800) );
  AND2_X1 U164bar ( .A1(inbar[191]), .A2(inbar[189]), .ZN(n800bar) );
  OR2_X1 U165 ( .A1(n799), .A2(n798), .ZN(n826) );
  AND2_X1 U165bar ( .A1(n799bar), .A2(n798bar), .ZN(n826bar) );
  OR2_X1 U166 ( .A1(n797), .A2(n796), .ZN(n798) );
  AND2_X1 U166bar ( .A1(n797bar), .A2(n796bar), .ZN(n798bar) );
  OR2_X1 U167 ( .A1(in[212]), .A2(in[193]), .ZN(n796) );
  AND2_X1 U167bar ( .A1(inbar[212]), .A2(inbar[193]), .ZN(n796bar) );
  OR2_X1 U168 ( .A1(in[238]), .A2(n795), .ZN(n797) );
  AND2_X1 U168bar ( .A1(inbar[238]), .A2(n795bar), .ZN(n797bar) );
  OR2_X1 U169 ( .A1(in[88]), .A2(in[247]), .ZN(n795) );
  AND2_X1 U169bar ( .A1(inbar[88]), .A2(inbar[247]), .ZN(n795bar) );
  OR2_X1 U170 ( .A1(n794), .A2(n793), .ZN(n799) );
  AND2_X1 U170bar ( .A1(n794bar), .A2(n793bar), .ZN(n799bar) );
  OR2_X1 U171 ( .A1(in[94]), .A2(in[92]), .ZN(n793) );
  AND2_X1 U171bar ( .A1(inbar[94]), .A2(inbar[92]), .ZN(n793bar) );
  OR2_X1 U172 ( .A1(in_52), .A2(n792), .ZN(n794) );
  AND2_X1 U172bar ( .A1(in_52bar), .A2(n792bar), .ZN(n794bar) );
  OR2_X1 U173 ( .A1(in_70), .A2(in_67), .ZN(n792) );
  AND2_X1 U173bar ( .A1(in_70bar), .A2(in_67bar), .ZN(n792bar) );
  OR2_X1 U174 ( .A1(n791), .A2(n790), .ZN(out[2]) );
  AND2_X1 U174bar ( .A1(n791bar), .A2(n790bar), .ZN(outbar[2]) );
  OR2_X1 U175 ( .A1(n789), .A2(n788), .ZN(n790) );
  AND2_X1 U175bar ( .A1(n789bar), .A2(n788bar), .ZN(n790bar) );
  OR2_X1 U176 ( .A1(n787), .A2(n786), .ZN(n788) );
  AND2_X1 U176bar ( .A1(n787bar), .A2(n786bar), .ZN(n788bar) );
  OR2_X1 U177 ( .A1(n819), .A2(n785), .ZN(n786) );
  AND2_X1 U177bar ( .A1(n819bar), .A2(n785bar), .ZN(n786bar) );
  OR2_X1 U178 ( .A1(n784), .A2(n783), .ZN(n819) );
  AND2_X1 U178bar ( .A1(n784bar), .A2(n783bar), .ZN(n819bar) );
  OR2_X1 U179 ( .A1(n782), .A2(n781), .ZN(n783) );
  AND2_X1 U179bar ( .A1(n782bar), .A2(n781bar), .ZN(n783bar) );
  OR2_X1 U180 ( .A1(n780), .A2(n779), .ZN(n781) );
  AND2_X1 U180bar ( .A1(n780bar), .A2(n779bar), .ZN(n781bar) );
  OR2_X1 U181 ( .A1(n962), .A2(n778), .ZN(n779) );
  AND2_X1 U181bar ( .A1(n962bar), .A2(n778bar), .ZN(n779bar) );
  OR2_X1 U182 ( .A1(n777), .A2(n776), .ZN(n962) );
  AND2_X1 U182bar ( .A1(n777bar), .A2(n776bar), .ZN(n962bar) );
  OR2_X1 U183 ( .A1(n775), .A2(n774), .ZN(n776) );
  AND2_X1 U183bar ( .A1(n775bar), .A2(n774bar), .ZN(n776bar) );
  OR2_X1 U184 ( .A1(n773), .A2(n772), .ZN(n774) );
  AND2_X1 U184bar ( .A1(n773bar), .A2(n772bar), .ZN(n774bar) );
  OR2_X1 U185 ( .A1(in[131]), .A2(in[120]), .ZN(n772) );
  AND2_X1 U185bar ( .A1(inbar[131]), .A2(inbar[120]), .ZN(n772bar) );
  OR2_X1 U186 ( .A1(in[153]), .A2(in[147]), .ZN(n773) );
  AND2_X1 U186bar ( .A1(inbar[153]), .A2(inbar[147]), .ZN(n773bar) );
  OR2_X1 U187 ( .A1(n771), .A2(n770), .ZN(n775) );
  AND2_X1 U187bar ( .A1(n771bar), .A2(n770bar), .ZN(n775bar) );
  OR2_X1 U188 ( .A1(in[170]), .A2(in[156]), .ZN(n770) );
  AND2_X1 U188bar ( .A1(inbar[170]), .A2(inbar[156]), .ZN(n770bar) );
  OR2_X1 U189 ( .A1(in[223]), .A2(in[190]), .ZN(n771) );
  AND2_X1 U189bar ( .A1(inbar[223]), .A2(inbar[190]), .ZN(n771bar) );
  OR2_X1 U190 ( .A1(n769), .A2(n768), .ZN(n777) );
  AND2_X1 U190bar ( .A1(n769bar), .A2(n768bar), .ZN(n777bar) );
  OR2_X1 U191 ( .A1(n767), .A2(n766), .ZN(n768) );
  AND2_X1 U191bar ( .A1(n767bar), .A2(n766bar), .ZN(n768bar) );
  OR2_X1 U192 ( .A1(in[236]), .A2(in[230]), .ZN(n766) );
  AND2_X1 U192bar ( .A1(inbar[236]), .A2(inbar[230]), .ZN(n766bar) );
  OR2_X1 U193 ( .A1(in[85]), .A2(in[240]), .ZN(n767) );
  AND2_X1 U193bar ( .A1(inbar[85]), .A2(inbar[240]), .ZN(n767bar) );
  OR2_X1 U194 ( .A1(n765), .A2(n764), .ZN(n769) );
  AND2_X1 U194bar ( .A1(n765bar), .A2(n764bar), .ZN(n769bar) );
  OR2_X1 U195 ( .A1(in_12), .A2(in[90]), .ZN(n764) );
  AND2_X1 U195bar ( .A1(in_12bar), .A2(inbar[90]), .ZN(n764bar) );
  OR2_X1 U196 ( .A1(in_39), .A2(in_28), .ZN(n765) );
  AND2_X1 U196bar ( .A1(in_39bar), .A2(in_28bar), .ZN(n765bar) );
  OR2_X1 U197 ( .A1(in[109]), .A2(n763), .ZN(n780) );
  AND2_X1 U197bar ( .A1(inbar[109]), .A2(n763bar), .ZN(n780bar) );
  OR2_X1 U198 ( .A1(n762), .A2(n761), .ZN(n782) );
  AND2_X1 U198bar ( .A1(n762bar), .A2(n761bar), .ZN(n782bar) );
  OR2_X1 U199 ( .A1(in[138]), .A2(in[129]), .ZN(n761) );
  AND2_X1 U199bar ( .A1(inbar[138]), .A2(inbar[129]), .ZN(n761bar) );
  OR2_X1 U200 ( .A1(in[157]), .A2(n760), .ZN(n762) );
  AND2_X1 U200bar ( .A1(inbar[157]), .A2(n760bar), .ZN(n762bar) );
  OR2_X1 U201 ( .A1(in[182]), .A2(in[167]), .ZN(n760) );
  AND2_X1 U201bar ( .A1(inbar[182]), .A2(inbar[167]), .ZN(n760bar) );
  OR2_X1 U202 ( .A1(n759), .A2(n758), .ZN(n784) );
  AND2_X1 U202bar ( .A1(n759bar), .A2(n758bar), .ZN(n784bar) );
  OR2_X1 U203 ( .A1(n757), .A2(n756), .ZN(n758) );
  AND2_X1 U203bar ( .A1(n757bar), .A2(n756bar), .ZN(n758bar) );
  OR2_X1 U204 ( .A1(in[195]), .A2(in[184]), .ZN(n756) );
  AND2_X1 U204bar ( .A1(inbar[195]), .A2(inbar[184]), .ZN(n756bar) );
  OR2_X1 U205 ( .A1(in[196]), .A2(n755), .ZN(n757) );
  AND2_X1 U205bar ( .A1(inbar[196]), .A2(n755bar), .ZN(n757bar) );
  OR2_X1 U206 ( .A1(in[215]), .A2(in[209]), .ZN(n755) );
  AND2_X1 U206bar ( .A1(inbar[215]), .A2(inbar[209]), .ZN(n755bar) );
  OR2_X1 U207 ( .A1(n754), .A2(n753), .ZN(n759) );
  AND2_X1 U207bar ( .A1(n754bar), .A2(n753bar), .ZN(n759bar) );
  OR2_X1 U208 ( .A1(in[93]), .A2(in[233]), .ZN(n753) );
  AND2_X1 U208bar ( .A1(inbar[93]), .A2(inbar[233]), .ZN(n753bar) );
  OR2_X1 U209 ( .A1(in_1), .A2(n752), .ZN(n754) );
  AND2_X1 U209bar ( .A1(in_1bar), .A2(n752bar), .ZN(n754bar) );
  OR2_X1 U210 ( .A1(in_69), .A2(in_66), .ZN(n752) );
  AND2_X1 U210bar ( .A1(in_69bar), .A2(in_66bar), .ZN(n752bar) );
  OR2_X1 U211 ( .A1(n966), .A2(n751), .ZN(n787) );
  AND2_X1 U211bar ( .A1(n966bar), .A2(n751bar), .ZN(n787bar) );
  OR2_X1 U212 ( .A1(in[134]), .A2(n750), .ZN(n751) );
  AND2_X1 U212bar ( .A1(inbar[134]), .A2(n750bar), .ZN(n751bar) );
  OR2_X1 U213 ( .A1(n749), .A2(n748), .ZN(n966) );
  AND2_X1 U213bar ( .A1(n749bar), .A2(n748bar), .ZN(n966bar) );
  OR2_X1 U214 ( .A1(n747), .A2(n746), .ZN(n748) );
  AND2_X1 U214bar ( .A1(n747bar), .A2(n746bar), .ZN(n748bar) );
  OR2_X1 U215 ( .A1(n745), .A2(n744), .ZN(n746) );
  AND2_X1 U215bar ( .A1(n745bar), .A2(n744bar), .ZN(n746bar) );
  OR2_X1 U216 ( .A1(in[136]), .A2(in[121]), .ZN(n744) );
  AND2_X1 U216bar ( .A1(inbar[136]), .A2(inbar[121]), .ZN(n744bar) );
  OR2_X1 U217 ( .A1(in[186]), .A2(in[174]), .ZN(n745) );
  AND2_X1 U217bar ( .A1(inbar[186]), .A2(inbar[174]), .ZN(n745bar) );
  OR2_X1 U218 ( .A1(n743), .A2(n742), .ZN(n747) );
  AND2_X1 U218bar ( .A1(n743bar), .A2(n742bar), .ZN(n747bar) );
  OR2_X1 U219 ( .A1(in[198]), .A2(in[197]), .ZN(n742) );
  AND2_X1 U219bar ( .A1(inbar[198]), .A2(inbar[197]), .ZN(n742bar) );
  OR2_X1 U220 ( .A1(in[214]), .A2(in[199]), .ZN(n743) );
  AND2_X1 U220bar ( .A1(inbar[214]), .A2(inbar[199]), .ZN(n743bar) );
  OR2_X1 U221 ( .A1(n741), .A2(n740), .ZN(n749) );
  AND2_X1 U221bar ( .A1(n741bar), .A2(n740bar), .ZN(n749bar) );
  OR2_X1 U222 ( .A1(n739), .A2(n738), .ZN(n740) );
  AND2_X1 U222bar ( .A1(n739bar), .A2(n738bar), .ZN(n740bar) );
  OR2_X1 U223 ( .A1(in[231]), .A2(in[220]), .ZN(n738) );
  AND2_X1 U223bar ( .A1(inbar[231]), .A2(inbar[220]), .ZN(n738bar) );
  OR2_X1 U224 ( .A1(in_25), .A2(in[245]), .ZN(n739) );
  AND2_X1 U224bar ( .A1(in_25bar), .A2(inbar[245]), .ZN(n739bar) );
  OR2_X1 U225 ( .A1(n737), .A2(n736), .ZN(n741) );
  AND2_X1 U225bar ( .A1(n737bar), .A2(n736bar), .ZN(n741bar) );
  OR2_X1 U226 ( .A1(in_53), .A2(in_29), .ZN(n736) );
  AND2_X1 U226bar ( .A1(in_53bar), .A2(in_29bar), .ZN(n736bar) );
  OR2_X1 U227 ( .A1(in_79), .A2(in_74), .ZN(n737) );
  AND2_X1 U227bar ( .A1(in_79bar), .A2(in_74bar), .ZN(n737bar) );
  OR2_X1 U228 ( .A1(n735), .A2(n734), .ZN(n789) );
  AND2_X1 U228bar ( .A1(n735bar), .A2(n734bar), .ZN(n789bar) );
  OR2_X1 U229 ( .A1(in[152]), .A2(in[140]), .ZN(n734) );
  AND2_X1 U229bar ( .A1(inbar[152]), .A2(inbar[140]), .ZN(n734bar) );
  OR2_X1 U230 ( .A1(in[155]), .A2(n733), .ZN(n735) );
  AND2_X1 U230bar ( .A1(inbar[155]), .A2(n733bar), .ZN(n735bar) );
  OR2_X1 U231 ( .A1(in[166]), .A2(in[165]), .ZN(n733) );
  AND2_X1 U231bar ( .A1(inbar[166]), .A2(inbar[165]), .ZN(n733bar) );
  OR2_X1 U232 ( .A1(n732), .A2(n731), .ZN(n791) );
  AND2_X1 U232bar ( .A1(n732bar), .A2(n731bar), .ZN(n791bar) );
  OR2_X1 U233 ( .A1(n730), .A2(n729), .ZN(n731) );
  AND2_X1 U233bar ( .A1(n730bar), .A2(n729bar), .ZN(n731bar) );
  OR2_X1 U234 ( .A1(in[202]), .A2(in[185]), .ZN(n729) );
  AND2_X1 U234bar ( .A1(inbar[202]), .A2(inbar[185]), .ZN(n729bar) );
  OR2_X1 U235 ( .A1(in[211]), .A2(n728), .ZN(n730) );
  AND2_X1 U235bar ( .A1(inbar[211]), .A2(n728bar), .ZN(n730bar) );
  OR2_X1 U236 ( .A1(in[255]), .A2(in[253]), .ZN(n728) );
  AND2_X1 U236bar ( .A1(inbar[255]), .A2(inbar[253]), .ZN(n728bar) );
  OR2_X1 U237 ( .A1(n727), .A2(n726), .ZN(n732) );
  AND2_X1 U237bar ( .A1(n727bar), .A2(n726bar), .ZN(n732bar) );
  OR2_X1 U238 ( .A1(in_35), .A2(in_15), .ZN(n726) );
  AND2_X1 U238bar ( .A1(in_35bar), .A2(in_15bar), .ZN(n726bar) );
  OR2_X1 U239 ( .A1(in_36), .A2(n725), .ZN(n727) );
  AND2_X1 U239bar ( .A1(in_36bar), .A2(n725bar), .ZN(n727bar) );
  OR2_X1 U240 ( .A1(in_48), .A2(in_40), .ZN(n725) );
  AND2_X1 U240bar ( .A1(in_48bar), .A2(in_40bar), .ZN(n725bar) );
  OR2_X1 U241 ( .A1(n724), .A2(n723), .ZN(out[1]) );
  AND2_X1 U241bar ( .A1(n724bar), .A2(n723bar), .ZN(outbar[1]) );
  OR2_X1 U242 ( .A1(n722), .A2(n721), .ZN(n723) );
  AND2_X1 U242bar ( .A1(n722bar), .A2(n721bar), .ZN(n723bar) );
  OR2_X1 U243 ( .A1(n720), .A2(n719), .ZN(n721) );
  AND2_X1 U243bar ( .A1(n720bar), .A2(n719bar), .ZN(n721bar) );
  OR2_X1 U244 ( .A1(n921), .A2(n887), .ZN(n719) );
  AND2_X1 U244bar ( .A1(n921bar), .A2(n887bar), .ZN(n719bar) );
  OR2_X1 U245 ( .A1(n718), .A2(n717), .ZN(n887) );
  AND2_X1 U245bar ( .A1(n718bar), .A2(n717bar), .ZN(n887bar) );
  OR2_X1 U246 ( .A1(n716), .A2(n715), .ZN(n717) );
  AND2_X1 U246bar ( .A1(n716bar), .A2(n715bar), .ZN(n717bar) );
  OR2_X1 U247 ( .A1(n714), .A2(n713), .ZN(n715) );
  AND2_X1 U247bar ( .A1(n714bar), .A2(n713bar), .ZN(n715bar) );
  OR2_X1 U248 ( .A1(in[116]), .A2(in[110]), .ZN(n713) );
  AND2_X1 U248bar ( .A1(inbar[116]), .A2(inbar[110]), .ZN(n713bar) );
  OR2_X1 U249 ( .A1(in[133]), .A2(in[130]), .ZN(n714) );
  AND2_X1 U249bar ( .A1(inbar[133]), .A2(inbar[130]), .ZN(n714bar) );
  OR2_X1 U250 ( .A1(n712), .A2(n711), .ZN(n716) );
  AND2_X1 U250bar ( .A1(n712bar), .A2(n711bar), .ZN(n716bar) );
  OR2_X1 U251 ( .A1(in[203]), .A2(in[135]), .ZN(n711) );
  AND2_X1 U251bar ( .A1(inbar[203]), .A2(inbar[135]), .ZN(n711bar) );
  OR2_X1 U252 ( .A1(in[232]), .A2(in[223]), .ZN(n712) );
  AND2_X1 U252bar ( .A1(inbar[232]), .A2(inbar[223]), .ZN(n712bar) );
  OR2_X1 U253 ( .A1(n710), .A2(n709), .ZN(n718) );
  AND2_X1 U253bar ( .A1(n710bar), .A2(n709bar), .ZN(n718bar) );
  OR2_X1 U254 ( .A1(n708), .A2(n707), .ZN(n709) );
  AND2_X1 U254bar ( .A1(n708bar), .A2(n707bar), .ZN(n709bar) );
  OR2_X1 U255 ( .A1(in[255]), .A2(in[233]), .ZN(n707) );
  AND2_X1 U255bar ( .A1(inbar[255]), .A2(inbar[233]), .ZN(n707bar) );
  OR2_X1 U256 ( .A1(in_53), .A2(in_34), .ZN(n708) );
  AND2_X1 U256bar ( .A1(in_53bar), .A2(in_34bar), .ZN(n708bar) );
  OR2_X1 U257 ( .A1(n706), .A2(n705), .ZN(n710) );
  AND2_X1 U257bar ( .A1(n706bar), .A2(n705bar), .ZN(n710bar) );
  OR2_X1 U258 ( .A1(in_57), .A2(in_55), .ZN(n705) );
  AND2_X1 U258bar ( .A1(in_57bar), .A2(in_55bar), .ZN(n705bar) );
  OR2_X1 U259 ( .A1(in_68), .A2(in_67), .ZN(n706) );
  AND2_X1 U259bar ( .A1(in_68bar), .A2(in_67bar), .ZN(n706bar) );
  OR2_X1 U260 ( .A1(n704), .A2(n703), .ZN(n921) );
  AND2_X1 U260bar ( .A1(n704bar), .A2(n703bar), .ZN(n921bar) );
  OR2_X1 U261 ( .A1(n702), .A2(n701), .ZN(n703) );
  AND2_X1 U261bar ( .A1(n702bar), .A2(n701bar), .ZN(n703bar) );
  OR2_X1 U262 ( .A1(n700), .A2(n699), .ZN(n701) );
  AND2_X1 U262bar ( .A1(n700bar), .A2(n699bar), .ZN(n701bar) );
  OR2_X1 U263 ( .A1(n944), .A2(n872), .ZN(n699) );
  AND2_X1 U263bar ( .A1(n944bar), .A2(n872bar), .ZN(n699bar) );
  OR2_X1 U264 ( .A1(n698), .A2(n697), .ZN(n872) );
  AND2_X1 U264bar ( .A1(n698bar), .A2(n697bar), .ZN(n872bar) );
  OR2_X1 U265 ( .A1(n696), .A2(n695), .ZN(n697) );
  AND2_X1 U265bar ( .A1(n696bar), .A2(n695bar), .ZN(n697bar) );
  OR2_X1 U266 ( .A1(n694), .A2(n693), .ZN(n695) );
  AND2_X1 U266bar ( .A1(n694bar), .A2(n693bar), .ZN(n695bar) );
  OR2_X1 U267 ( .A1(in[121]), .A2(in[102]), .ZN(n693) );
  AND2_X1 U267bar ( .A1(inbar[121]), .A2(inbar[102]), .ZN(n693bar) );
  OR2_X1 U268 ( .A1(in[162]), .A2(in[161]), .ZN(n694) );
  AND2_X1 U268bar ( .A1(inbar[162]), .A2(inbar[161]), .ZN(n694bar) );
  OR2_X1 U269 ( .A1(n692), .A2(n691), .ZN(n696) );
  AND2_X1 U269bar ( .A1(n692bar), .A2(n691bar), .ZN(n696bar) );
  OR2_X1 U270 ( .A1(in[192]), .A2(in[178]), .ZN(n691) );
  AND2_X1 U270bar ( .A1(inbar[192]), .A2(inbar[178]), .ZN(n691bar) );
  OR2_X1 U271 ( .A1(in[244]), .A2(in[209]), .ZN(n692) );
  AND2_X1 U271bar ( .A1(inbar[244]), .A2(inbar[209]), .ZN(n692bar) );
  OR2_X1 U272 ( .A1(n690), .A2(n689), .ZN(n698) );
  AND2_X1 U272bar ( .A1(n690bar), .A2(n689bar), .ZN(n698bar) );
  OR2_X1 U273 ( .A1(n688), .A2(n687), .ZN(n689) );
  AND2_X1 U273bar ( .A1(n688bar), .A2(n687bar), .ZN(n689bar) );
  OR2_X1 U274 ( .A1(in[90]), .A2(in[254]), .ZN(n687) );
  AND2_X1 U274bar ( .A1(inbar[90]), .A2(inbar[254]), .ZN(n687bar) );
  OR2_X1 U275 ( .A1(in_36), .A2(in_32), .ZN(n688) );
  AND2_X1 U275bar ( .A1(in_36bar), .A2(in_32bar), .ZN(n688bar) );
  OR2_X1 U276 ( .A1(n686), .A2(n685), .ZN(n690) );
  AND2_X1 U276bar ( .A1(n686bar), .A2(n685bar), .ZN(n690bar) );
  OR2_X1 U277 ( .A1(in_62), .A2(in_37), .ZN(n685) );
  AND2_X1 U277bar ( .A1(in_62bar), .A2(in_37bar), .ZN(n685bar) );
  OR2_X1 U278 ( .A1(in_75), .A2(in_73), .ZN(n686) );
  AND2_X1 U278bar ( .A1(in_75bar), .A2(in_73bar), .ZN(n686bar) );
  OR2_X1 U279 ( .A1(n684), .A2(n683), .ZN(n944) );
  AND2_X1 U279bar ( .A1(n684bar), .A2(n683bar), .ZN(n944bar) );
  OR2_X1 U280 ( .A1(n682), .A2(n681), .ZN(n683) );
  AND2_X1 U280bar ( .A1(n682bar), .A2(n681bar), .ZN(n683bar) );
  OR2_X1 U281 ( .A1(n680), .A2(n679), .ZN(n681) );
  AND2_X1 U281bar ( .A1(n680bar), .A2(n679bar), .ZN(n681bar) );
  OR2_X1 U282 ( .A1(in[171]), .A2(in[153]), .ZN(n679) );
  AND2_X1 U282bar ( .A1(inbar[171]), .A2(inbar[153]), .ZN(n679bar) );
  OR2_X1 U283 ( .A1(in[187]), .A2(in[176]), .ZN(n680) );
  AND2_X1 U283bar ( .A1(inbar[187]), .A2(inbar[176]), .ZN(n680bar) );
  OR2_X1 U284 ( .A1(n678), .A2(n677), .ZN(n682) );
  AND2_X1 U284bar ( .A1(n678bar), .A2(n677bar), .ZN(n682bar) );
  OR2_X1 U285 ( .A1(in[245]), .A2(in[211]), .ZN(n677) );
  AND2_X1 U285bar ( .A1(inbar[245]), .A2(inbar[211]), .ZN(n677bar) );
  OR2_X1 U286 ( .A1(in[97]), .A2(in[88]), .ZN(n678) );
  AND2_X1 U286bar ( .A1(inbar[97]), .A2(inbar[88]), .ZN(n678bar) );
  OR2_X1 U287 ( .A1(n676), .A2(n675), .ZN(n684) );
  AND2_X1 U287bar ( .A1(n676bar), .A2(n675bar), .ZN(n684bar) );
  OR2_X1 U288 ( .A1(n674), .A2(n673), .ZN(n675) );
  AND2_X1 U288bar ( .A1(n674bar), .A2(n673bar), .ZN(n675bar) );
  OR2_X1 U289 ( .A1(in_10), .A2(in_0), .ZN(n673) );
  AND2_X1 U289bar ( .A1(in_10bar), .A2(in_0bar), .ZN(n673bar) );
  OR2_X1 U290 ( .A1(in_59), .A2(in_5), .ZN(n674) );
  AND2_X1 U290bar ( .A1(in_59bar), .A2(in_5bar), .ZN(n674bar) );
  OR2_X1 U291 ( .A1(n672), .A2(n671), .ZN(n676) );
  AND2_X1 U291bar ( .A1(n672bar), .A2(n671bar), .ZN(n676bar) );
  OR2_X1 U292 ( .A1(in_60), .A2(in_6), .ZN(n671) );
  AND2_X1 U292bar ( .A1(in_60bar), .A2(in_6bar), .ZN(n671bar) );
  OR2_X1 U293 ( .A1(in_77), .A2(in_69), .ZN(n672) );
  AND2_X1 U293bar ( .A1(in_77bar), .A2(in_69bar), .ZN(n672bar) );
  OR2_X1 U294 ( .A1(in[113]), .A2(n864), .ZN(n700) );
  AND2_X1 U294bar ( .A1(inbar[113]), .A2(n864bar), .ZN(n700bar) );
  OR2_X1 U295 ( .A1(n670), .A2(n669), .ZN(n864) );
  AND2_X1 U295bar ( .A1(n670bar), .A2(n669bar), .ZN(n864bar) );
  OR2_X1 U296 ( .A1(n668), .A2(n667), .ZN(n669) );
  AND2_X1 U296bar ( .A1(n668bar), .A2(n667bar), .ZN(n669bar) );
  OR2_X1 U297 ( .A1(n666), .A2(n665), .ZN(n667) );
  AND2_X1 U297bar ( .A1(n666bar), .A2(n665bar), .ZN(n667bar) );
  OR2_X1 U298 ( .A1(in[125]), .A2(in[107]), .ZN(n665) );
  AND2_X1 U298bar ( .A1(inbar[125]), .A2(inbar[107]), .ZN(n665bar) );
  OR2_X1 U299 ( .A1(in[138]), .A2(in[126]), .ZN(n666) );
  AND2_X1 U299bar ( .A1(inbar[138]), .A2(inbar[126]), .ZN(n666bar) );
  OR2_X1 U300 ( .A1(n664), .A2(n663), .ZN(n668) );
  AND2_X1 U300bar ( .A1(n664bar), .A2(n663bar), .ZN(n668bar) );
  OR2_X1 U301 ( .A1(in[189]), .A2(in[143]), .ZN(n663) );
  AND2_X1 U301bar ( .A1(inbar[189]), .A2(inbar[143]), .ZN(n663bar) );
  OR2_X1 U302 ( .A1(in[99]), .A2(in[214]), .ZN(n664) );
  AND2_X1 U302bar ( .A1(inbar[99]), .A2(inbar[214]), .ZN(n664bar) );
  OR2_X1 U303 ( .A1(n662), .A2(n661), .ZN(n670) );
  AND2_X1 U303bar ( .A1(n662bar), .A2(n661bar), .ZN(n670bar) );
  OR2_X1 U304 ( .A1(n660), .A2(n659), .ZN(n661) );
  AND2_X1 U304bar ( .A1(n660bar), .A2(n659bar), .ZN(n661bar) );
  OR2_X1 U305 ( .A1(in_15), .A2(in_12), .ZN(n659) );
  AND2_X1 U305bar ( .A1(in_15bar), .A2(in_12bar), .ZN(n659bar) );
  OR2_X1 U306 ( .A1(in_20), .A2(in_2), .ZN(n660) );
  AND2_X1 U306bar ( .A1(in_20bar), .A2(in_2bar), .ZN(n660bar) );
  OR2_X1 U307 ( .A1(n658), .A2(n657), .ZN(n662) );
  AND2_X1 U307bar ( .A1(n658bar), .A2(n657bar), .ZN(n662bar) );
  OR2_X1 U308 ( .A1(in_30), .A2(in_3), .ZN(n657) );
  AND2_X1 U308bar ( .A1(in_30bar), .A2(in_3bar), .ZN(n657bar) );
  OR2_X1 U309 ( .A1(in_4), .A2(in_38), .ZN(n658) );
  AND2_X1 U309bar ( .A1(in_4bar), .A2(in_38bar), .ZN(n658bar) );
  OR2_X1 U310 ( .A1(n656), .A2(n655), .ZN(n702) );
  AND2_X1 U310bar ( .A1(n656bar), .A2(n655bar), .ZN(n702bar) );
  OR2_X1 U311 ( .A1(in[148]), .A2(in[137]), .ZN(n655) );
  AND2_X1 U311bar ( .A1(inbar[148]), .A2(inbar[137]), .ZN(n655bar) );
  OR2_X1 U312 ( .A1(in[149]), .A2(n654), .ZN(n656) );
  AND2_X1 U312bar ( .A1(inbar[149]), .A2(n654bar), .ZN(n656bar) );
  OR2_X1 U313 ( .A1(in[195]), .A2(in[190]), .ZN(n654) );
  AND2_X1 U313bar ( .A1(inbar[195]), .A2(inbar[190]), .ZN(n654bar) );
  OR2_X1 U314 ( .A1(n653), .A2(n652), .ZN(n704) );
  AND2_X1 U314bar ( .A1(n653bar), .A2(n652bar), .ZN(n704bar) );
  OR2_X1 U315 ( .A1(n651), .A2(n650), .ZN(n652) );
  AND2_X1 U315bar ( .A1(n651bar), .A2(n650bar), .ZN(n652bar) );
  OR2_X1 U316 ( .A1(in[98]), .A2(in[197]), .ZN(n650) );
  AND2_X1 U316bar ( .A1(inbar[98]), .A2(inbar[197]), .ZN(n650bar) );
  OR2_X1 U317 ( .A1(in_11), .A2(n649), .ZN(n651) );
  AND2_X1 U317bar ( .A1(in_11bar), .A2(n649bar), .ZN(n651bar) );
  OR2_X1 U318 ( .A1(in_26), .A2(in_14), .ZN(n649) );
  AND2_X1 U318bar ( .A1(in_26bar), .A2(in_14bar), .ZN(n649bar) );
  OR2_X1 U319 ( .A1(n648), .A2(n647), .ZN(n653) );
  AND2_X1 U319bar ( .A1(n648bar), .A2(n647bar), .ZN(n653bar) );
  OR2_X1 U320 ( .A1(in_35), .A2(in_27), .ZN(n647) );
  AND2_X1 U320bar ( .A1(in_35bar), .A2(in_27bar), .ZN(n647bar) );
  OR2_X1 U321 ( .A1(in_50), .A2(n646), .ZN(n648) );
  AND2_X1 U321bar ( .A1(in_50bar), .A2(n646bar), .ZN(n648bar) );
  OR2_X1 U322 ( .A1(in_78), .A2(in_61), .ZN(n646) );
  AND2_X1 U322bar ( .A1(in_78bar), .A2(in_61bar), .ZN(n646bar) );
  OR2_X1 U323 ( .A1(n942), .A2(n645), .ZN(n720) );
  AND2_X1 U323bar ( .A1(n942bar), .A2(n645bar), .ZN(n720bar) );
  OR2_X1 U324 ( .A1(in[106]), .A2(n863), .ZN(n645) );
  AND2_X1 U324bar ( .A1(inbar[106]), .A2(n863bar), .ZN(n645bar) );
  OR2_X1 U325 ( .A1(n644), .A2(n643), .ZN(n863) );
  AND2_X1 U325bar ( .A1(n644bar), .A2(n643bar), .ZN(n863bar) );
  OR2_X1 U326 ( .A1(n642), .A2(n641), .ZN(n643) );
  AND2_X1 U326bar ( .A1(n642bar), .A2(n641bar), .ZN(n643bar) );
  OR2_X1 U327 ( .A1(n640), .A2(n639), .ZN(n641) );
  AND2_X1 U327bar ( .A1(n640bar), .A2(n639bar), .ZN(n641bar) );
  OR2_X1 U328 ( .A1(in[127]), .A2(in[122]), .ZN(n639) );
  AND2_X1 U328bar ( .A1(inbar[127]), .A2(inbar[122]), .ZN(n639bar) );
  OR2_X1 U329 ( .A1(in[156]), .A2(in[132]), .ZN(n640) );
  AND2_X1 U329bar ( .A1(inbar[156]), .A2(inbar[132]), .ZN(n640bar) );
  OR2_X1 U330 ( .A1(n638), .A2(n637), .ZN(n642) );
  AND2_X1 U330bar ( .A1(n638bar), .A2(n637bar), .ZN(n642bar) );
  OR2_X1 U331 ( .A1(in[159]), .A2(in[157]), .ZN(n637) );
  AND2_X1 U331bar ( .A1(inbar[159]), .A2(inbar[157]), .ZN(n637bar) );
  OR2_X1 U332 ( .A1(in[185]), .A2(in[169]), .ZN(n638) );
  AND2_X1 U332bar ( .A1(inbar[185]), .A2(inbar[169]), .ZN(n638bar) );
  OR2_X1 U333 ( .A1(n636), .A2(n635), .ZN(n644) );
  AND2_X1 U333bar ( .A1(n636bar), .A2(n635bar), .ZN(n644bar) );
  OR2_X1 U334 ( .A1(n634), .A2(n633), .ZN(n635) );
  AND2_X1 U334bar ( .A1(n634bar), .A2(n633bar), .ZN(n635bar) );
  OR2_X1 U335 ( .A1(in[239]), .A2(in[218]), .ZN(n633) );
  AND2_X1 U335bar ( .A1(inbar[239]), .A2(inbar[218]), .ZN(n633bar) );
  OR2_X1 U336 ( .A1(in_13), .A2(in[87]), .ZN(n634) );
  AND2_X1 U336bar ( .A1(in_13bar), .A2(inbar[87]), .ZN(n634bar) );
  OR2_X1 U337 ( .A1(n632), .A2(n631), .ZN(n636) );
  AND2_X1 U337bar ( .A1(n632bar), .A2(n631bar), .ZN(n636bar) );
  OR2_X1 U338 ( .A1(in_72), .A2(in_70), .ZN(n631) );
  AND2_X1 U338bar ( .A1(in_72bar), .A2(in_70bar), .ZN(n631bar) );
  OR2_X1 U339 ( .A1(in_80), .A2(in_74), .ZN(n632) );
  AND2_X1 U339bar ( .A1(in_80bar), .A2(in_74bar), .ZN(n632bar) );
  OR2_X1 U340 ( .A1(n630), .A2(n629), .ZN(n942) );
  AND2_X1 U340bar ( .A1(n630bar), .A2(n629bar), .ZN(n942bar) );
  OR2_X1 U341 ( .A1(n628), .A2(n627), .ZN(n629) );
  AND2_X1 U341bar ( .A1(n628bar), .A2(n627bar), .ZN(n629bar) );
  OR2_X1 U342 ( .A1(n626), .A2(n625), .ZN(n627) );
  AND2_X1 U342bar ( .A1(n626bar), .A2(n625bar), .ZN(n627bar) );
  OR2_X1 U343 ( .A1(in[146]), .A2(in[100]), .ZN(n625) );
  AND2_X1 U343bar ( .A1(inbar[146]), .A2(inbar[100]), .ZN(n625bar) );
  OR2_X1 U344 ( .A1(in[168]), .A2(in[152]), .ZN(n626) );
  AND2_X1 U344bar ( .A1(inbar[168]), .A2(inbar[152]), .ZN(n626bar) );
  OR2_X1 U345 ( .A1(n624), .A2(n623), .ZN(n628) );
  AND2_X1 U345bar ( .A1(n624bar), .A2(n623bar), .ZN(n628bar) );
  OR2_X1 U346 ( .A1(in[199]), .A2(in[182]), .ZN(n623) );
  AND2_X1 U346bar ( .A1(inbar[199]), .A2(inbar[182]), .ZN(n623bar) );
  OR2_X1 U347 ( .A1(in[236]), .A2(in[204]), .ZN(n624) );
  AND2_X1 U347bar ( .A1(inbar[236]), .A2(inbar[204]), .ZN(n624bar) );
  OR2_X1 U348 ( .A1(n622), .A2(n621), .ZN(n630) );
  AND2_X1 U348bar ( .A1(n622bar), .A2(n621bar), .ZN(n630bar) );
  OR2_X1 U349 ( .A1(n620), .A2(n619), .ZN(n621) );
  AND2_X1 U349bar ( .A1(n620bar), .A2(n619bar), .ZN(n621bar) );
  OR2_X1 U350 ( .A1(in[89]), .A2(in[246]), .ZN(n619) );
  AND2_X1 U350bar ( .A1(inbar[89]), .A2(inbar[246]), .ZN(n619bar) );
  OR2_X1 U351 ( .A1(in[95]), .A2(in[92]), .ZN(n620) );
  AND2_X1 U351bar ( .A1(inbar[95]), .A2(inbar[92]), .ZN(n620bar) );
  OR2_X1 U352 ( .A1(n618), .A2(n617), .ZN(n622) );
  AND2_X1 U352bar ( .A1(n618bar), .A2(n617bar), .ZN(n622bar) );
  OR2_X1 U353 ( .A1(in_22), .A2(in_16), .ZN(n617) );
  AND2_X1 U353bar ( .A1(in_22bar), .A2(in_16bar), .ZN(n617bar) );
  OR2_X1 U354 ( .A1(in_51), .A2(in_49), .ZN(n618) );
  AND2_X1 U354bar ( .A1(in_51bar), .A2(in_49bar), .ZN(n618bar) );
  OR2_X1 U355 ( .A1(n616), .A2(n615), .ZN(n722) );
  AND2_X1 U355bar ( .A1(n616bar), .A2(n615bar), .ZN(n722bar) );
  OR2_X1 U356 ( .A1(in[158]), .A2(in[115]), .ZN(n615) );
  AND2_X1 U356bar ( .A1(inbar[158]), .A2(inbar[115]), .ZN(n615bar) );
  OR2_X1 U357 ( .A1(in[163]), .A2(n614), .ZN(n616) );
  AND2_X1 U357bar ( .A1(inbar[163]), .A2(n614bar), .ZN(n616bar) );
  OR2_X1 U358 ( .A1(in[206]), .A2(in[165]), .ZN(n614) );
  AND2_X1 U358bar ( .A1(inbar[206]), .A2(inbar[165]), .ZN(n614bar) );
  OR2_X1 U359 ( .A1(n613), .A2(n612), .ZN(n724) );
  AND2_X1 U359bar ( .A1(n613bar), .A2(n612bar), .ZN(n724bar) );
  OR2_X1 U360 ( .A1(n611), .A2(n610), .ZN(n612) );
  AND2_X1 U360bar ( .A1(n611bar), .A2(n610bar), .ZN(n612bar) );
  OR2_X1 U361 ( .A1(in[213]), .A2(in[207]), .ZN(n610) );
  AND2_X1 U361bar ( .A1(inbar[213]), .A2(inbar[207]), .ZN(n610bar) );
  OR2_X1 U362 ( .A1(in[215]), .A2(n609), .ZN(n611) );
  AND2_X1 U362bar ( .A1(inbar[215]), .A2(n609bar), .ZN(n611bar) );
  OR2_X1 U363 ( .A1(in[230]), .A2(in[220]), .ZN(n609) );
  AND2_X1 U363bar ( .A1(inbar[230]), .A2(inbar[220]), .ZN(n609bar) );
  OR2_X1 U364 ( .A1(n608), .A2(n607), .ZN(n613) );
  AND2_X1 U364bar ( .A1(n608bar), .A2(n607bar), .ZN(n613bar) );
  OR2_X1 U365 ( .A1(in[251]), .A2(in[234]), .ZN(n607) );
  AND2_X1 U365bar ( .A1(inbar[251]), .A2(inbar[234]), .ZN(n607bar) );
  OR2_X1 U366 ( .A1(in_17), .A2(n606), .ZN(n608) );
  AND2_X1 U366bar ( .A1(in_17bar), .A2(n606bar), .ZN(n608bar) );
  OR2_X1 U367 ( .A1(in_65), .A2(in_56), .ZN(n606) );
  AND2_X1 U367bar ( .A1(in_65bar), .A2(in_56bar), .ZN(n606bar) );
  OR2_X1 U368 ( .A1(n605), .A2(n604), .ZN(out[0]) );
  AND2_X1 U368bar ( .A1(n605bar), .A2(n604bar), .ZN(outbar[0]) );
  OR2_X1 U369 ( .A1(n603), .A2(n602), .ZN(n604) );
  AND2_X1 U369bar ( .A1(n603bar), .A2(n602bar), .ZN(n604bar) );
  OR2_X1 U370 ( .A1(n601), .A2(n600), .ZN(n602) );
  AND2_X1 U370bar ( .A1(n601bar), .A2(n600bar), .ZN(n602bar) );
  OR2_X1 U371 ( .A1(n820), .A2(n785), .ZN(n600) );
  AND2_X1 U371bar ( .A1(n820bar), .A2(n785bar), .ZN(n600bar) );
  OR2_X1 U372 ( .A1(n599), .A2(n598), .ZN(n785) );
  AND2_X1 U372bar ( .A1(n599bar), .A2(n598bar), .ZN(n785bar) );
  OR2_X1 U373 ( .A1(n597), .A2(n596), .ZN(n598) );
  AND2_X1 U373bar ( .A1(n597bar), .A2(n596bar), .ZN(n598bar) );
  OR2_X1 U374 ( .A1(n595), .A2(n594), .ZN(n596) );
  AND2_X1 U374bar ( .A1(n595bar), .A2(n594bar), .ZN(n596bar) );
  OR2_X1 U375 ( .A1(in[135]), .A2(in[104]), .ZN(n594) );
  AND2_X1 U375bar ( .A1(inbar[135]), .A2(inbar[104]), .ZN(n594bar) );
  OR2_X1 U376 ( .A1(in[188]), .A2(in[178]), .ZN(n595) );
  AND2_X1 U376bar ( .A1(inbar[188]), .A2(inbar[178]), .ZN(n595bar) );
  OR2_X1 U377 ( .A1(n593), .A2(n592), .ZN(n597) );
  AND2_X1 U377bar ( .A1(n593bar), .A2(n592bar), .ZN(n597bar) );
  OR2_X1 U378 ( .A1(in[217]), .A2(in[194]), .ZN(n592) );
  AND2_X1 U378bar ( .A1(inbar[217]), .A2(inbar[194]), .ZN(n592bar) );
  OR2_X1 U379 ( .A1(in[237]), .A2(in[218]), .ZN(n593) );
  AND2_X1 U379bar ( .A1(inbar[237]), .A2(inbar[218]), .ZN(n593bar) );
  OR2_X1 U380 ( .A1(n591), .A2(n590), .ZN(n599) );
  AND2_X1 U380bar ( .A1(n591bar), .A2(n590bar), .ZN(n599bar) );
  OR2_X1 U381 ( .A1(n589), .A2(n588), .ZN(n590) );
  AND2_X1 U381bar ( .A1(n589bar), .A2(n588bar), .ZN(n590bar) );
  OR2_X1 U382 ( .A1(in_2), .A2(in_10), .ZN(n588) );
  AND2_X1 U382bar ( .A1(in_2bar), .A2(in_10bar), .ZN(n588bar) );
  OR2_X1 U383 ( .A1(in_47), .A2(in_22), .ZN(n589) );
  AND2_X1 U383bar ( .A1(in_47bar), .A2(in_22bar), .ZN(n589bar) );
  OR2_X1 U384 ( .A1(n587), .A2(n586), .ZN(n591) );
  AND2_X1 U384bar ( .A1(n587bar), .A2(n586bar), .ZN(n591bar) );
  OR2_X1 U385 ( .A1(in_56), .A2(in_54), .ZN(n586) );
  AND2_X1 U385bar ( .A1(in_56bar), .A2(in_54bar), .ZN(n586bar) );
  OR2_X1 U386 ( .A1(in_63), .A2(in_61), .ZN(n587) );
  AND2_X1 U386bar ( .A1(in_63bar), .A2(in_61bar), .ZN(n587bar) );
  OR2_X1 U387 ( .A1(n585), .A2(n584), .ZN(n820) );
  AND2_X1 U387bar ( .A1(n585bar), .A2(n584bar), .ZN(n820bar) );
  OR2_X1 U388 ( .A1(n583), .A2(n582), .ZN(n584) );
  AND2_X1 U388bar ( .A1(n583bar), .A2(n582bar), .ZN(n584bar) );
  OR2_X1 U389 ( .A1(n581), .A2(n580), .ZN(n582) );
  AND2_X1 U389bar ( .A1(n581bar), .A2(n580bar), .ZN(n582bar) );
  OR2_X1 U390 ( .A1(in[158]), .A2(in[142]), .ZN(n580) );
  AND2_X1 U390bar ( .A1(inbar[158]), .A2(inbar[142]), .ZN(n580bar) );
  OR2_X1 U391 ( .A1(in[175]), .A2(in[164]), .ZN(n581) );
  AND2_X1 U391bar ( .A1(inbar[175]), .A2(inbar[164]), .ZN(n581bar) );
  OR2_X1 U392 ( .A1(n579), .A2(n578), .ZN(n583) );
  AND2_X1 U392bar ( .A1(n579bar), .A2(n578bar), .ZN(n583bar) );
  OR2_X1 U393 ( .A1(in[228]), .A2(in[204]), .ZN(n578) );
  AND2_X1 U393bar ( .A1(inbar[228]), .A2(inbar[204]), .ZN(n578bar) );
  OR2_X1 U394 ( .A1(in[91]), .A2(in[87]), .ZN(n579) );
  AND2_X1 U394bar ( .A1(inbar[91]), .A2(inbar[87]), .ZN(n579bar) );
  OR2_X1 U395 ( .A1(n577), .A2(n576), .ZN(n585) );
  AND2_X1 U395bar ( .A1(n577bar), .A2(n576bar), .ZN(n585bar) );
  OR2_X1 U396 ( .A1(n575), .A2(n574), .ZN(n576) );
  AND2_X1 U396bar ( .A1(n575bar), .A2(n574bar), .ZN(n576bar) );
  OR2_X1 U397 ( .A1(in_21), .A2(in_11), .ZN(n574) );
  AND2_X1 U397bar ( .A1(in_21bar), .A2(in_11bar), .ZN(n574bar) );
  OR2_X1 U398 ( .A1(in_5), .A2(in_3), .ZN(n575) );
  AND2_X1 U398bar ( .A1(in_5bar), .A2(in_3bar), .ZN(n575bar) );
  OR2_X1 U399 ( .A1(n573), .A2(n572), .ZN(n577) );
  AND2_X1 U399bar ( .A1(n573bar), .A2(n572bar), .ZN(n577bar) );
  OR2_X1 U400 ( .A1(in_68), .A2(in_64), .ZN(n572) );
  AND2_X1 U400bar ( .A1(in_68bar), .A2(in_64bar), .ZN(n572bar) );
  OR2_X1 U401 ( .A1(in_76), .A2(in_73), .ZN(n573) );
  AND2_X1 U401bar ( .A1(in_76bar), .A2(in_73bar), .ZN(n573bar) );
  OR2_X1 U402 ( .A1(n778), .A2(n571), .ZN(n601) );
  AND2_X1 U402bar ( .A1(n778bar), .A2(n571bar), .ZN(n601bar) );
  OR2_X1 U403 ( .A1(in[100]), .A2(n965), .ZN(n571) );
  AND2_X1 U403bar ( .A1(inbar[100]), .A2(n965bar), .ZN(n571bar) );
  OR2_X1 U404 ( .A1(n570), .A2(n569), .ZN(n965) );
  AND2_X1 U404bar ( .A1(n570bar), .A2(n569bar), .ZN(n965bar) );
  OR2_X1 U405 ( .A1(n568), .A2(n567), .ZN(n569) );
  AND2_X1 U405bar ( .A1(n568bar), .A2(n567bar), .ZN(n569bar) );
  OR2_X1 U406 ( .A1(n566), .A2(n565), .ZN(n567) );
  AND2_X1 U406bar ( .A1(n566bar), .A2(n565bar), .ZN(n567bar) );
  OR2_X1 U407 ( .A1(n817), .A2(n750), .ZN(n565) );
  AND2_X1 U407bar ( .A1(n817bar), .A2(n750bar), .ZN(n565bar) );
  OR2_X1 U408 ( .A1(n564), .A2(n563), .ZN(n750) );
  AND2_X1 U408bar ( .A1(n564bar), .A2(n563bar), .ZN(n750bar) );
  OR2_X1 U409 ( .A1(n562), .A2(n561), .ZN(n563) );
  AND2_X1 U409bar ( .A1(n562bar), .A2(n561bar), .ZN(n563bar) );
  OR2_X1 U410 ( .A1(n560), .A2(n559), .ZN(n561) );
  AND2_X1 U410bar ( .A1(n560bar), .A2(n559bar), .ZN(n561bar) );
  OR2_X1 U411 ( .A1(in[119]), .A2(in[103]), .ZN(n559) );
  AND2_X1 U411bar ( .A1(inbar[119]), .A2(inbar[103]), .ZN(n559bar) );
  OR2_X1 U412 ( .A1(in[137]), .A2(in[133]), .ZN(n560) );
  AND2_X1 U412bar ( .A1(inbar[137]), .A2(inbar[133]), .ZN(n560bar) );
  OR2_X1 U413 ( .A1(n558), .A2(n557), .ZN(n562) );
  AND2_X1 U413bar ( .A1(n558bar), .A2(n557bar), .ZN(n562bar) );
  OR2_X1 U414 ( .A1(in[176]), .A2(in[173]), .ZN(n557) );
  AND2_X1 U414bar ( .A1(inbar[176]), .A2(inbar[173]), .ZN(n557bar) );
  OR2_X1 U415 ( .A1(in[210]), .A2(in[181]), .ZN(n558) );
  AND2_X1 U415bar ( .A1(inbar[210]), .A2(inbar[181]), .ZN(n558bar) );
  OR2_X1 U416 ( .A1(n556), .A2(n555), .ZN(n564) );
  AND2_X1 U416bar ( .A1(n556bar), .A2(n555bar), .ZN(n564bar) );
  OR2_X1 U417 ( .A1(n554), .A2(n553), .ZN(n555) );
  AND2_X1 U417bar ( .A1(n554bar), .A2(n553bar), .ZN(n555bar) );
  OR2_X1 U418 ( .A1(in_13), .A2(in[234]), .ZN(n553) );
  AND2_X1 U418bar ( .A1(in_13bar), .A2(inbar[234]), .ZN(n553bar) );
  OR2_X1 U419 ( .A1(in_38), .A2(in_32), .ZN(n554) );
  AND2_X1 U419bar ( .A1(in_38bar), .A2(in_32bar), .ZN(n554bar) );
  OR2_X1 U420 ( .A1(n552), .A2(n551), .ZN(n556) );
  AND2_X1 U420bar ( .A1(n552bar), .A2(n551bar), .ZN(n556bar) );
  OR2_X1 U421 ( .A1(in_42), .A2(in_41), .ZN(n551) );
  AND2_X1 U421bar ( .A1(in_42bar), .A2(in_41bar), .ZN(n551bar) );
  OR2_X1 U422 ( .A1(in_7), .A2(in_49), .ZN(n552) );
  AND2_X1 U422bar ( .A1(in_7bar), .A2(in_49bar), .ZN(n552bar) );
  OR2_X1 U423 ( .A1(n550), .A2(n549), .ZN(n817) );
  AND2_X1 U423bar ( .A1(n550bar), .A2(n549bar), .ZN(n817bar) );
  OR2_X1 U424 ( .A1(n548), .A2(n547), .ZN(n549) );
  AND2_X1 U424bar ( .A1(n548bar), .A2(n547bar), .ZN(n549bar) );
  OR2_X1 U425 ( .A1(n546), .A2(n545), .ZN(n547) );
  AND2_X1 U425bar ( .A1(n546bar), .A2(n545bar), .ZN(n547bar) );
  OR2_X1 U426 ( .A1(in[159]), .A2(in[105]), .ZN(n545) );
  AND2_X1 U426bar ( .A1(inbar[159]), .A2(inbar[105]), .ZN(n545bar) );
  OR2_X1 U427 ( .A1(in[206]), .A2(in[183]), .ZN(n546) );
  AND2_X1 U427bar ( .A1(inbar[206]), .A2(inbar[183]), .ZN(n546bar) );
  OR2_X1 U428 ( .A1(n544), .A2(n543), .ZN(n548) );
  AND2_X1 U428bar ( .A1(n544bar), .A2(n543bar), .ZN(n548bar) );
  OR2_X1 U429 ( .A1(in[229]), .A2(in[219]), .ZN(n543) );
  AND2_X1 U429bar ( .A1(inbar[229]), .A2(inbar[219]), .ZN(n543bar) );
  OR2_X1 U430 ( .A1(in[235]), .A2(in[232]), .ZN(n544) );
  AND2_X1 U430bar ( .A1(inbar[235]), .A2(inbar[232]), .ZN(n544bar) );
  OR2_X1 U431 ( .A1(n542), .A2(n541), .ZN(n550) );
  AND2_X1 U431bar ( .A1(n542bar), .A2(n541bar), .ZN(n550bar) );
  OR2_X1 U432 ( .A1(n540), .A2(n539), .ZN(n541) );
  AND2_X1 U432bar ( .A1(n540bar), .A2(n539bar), .ZN(n541bar) );
  OR2_X1 U433 ( .A1(in[249]), .A2(in[242]), .ZN(n539) );
  AND2_X1 U433bar ( .A1(inbar[249]), .A2(inbar[242]), .ZN(n539bar) );
  OR2_X1 U434 ( .A1(in[89]), .A2(in[254]), .ZN(n540) );
  AND2_X1 U434bar ( .A1(inbar[89]), .A2(inbar[254]), .ZN(n540bar) );
  OR2_X1 U435 ( .A1(n538), .A2(n537), .ZN(n542) );
  AND2_X1 U435bar ( .A1(n538bar), .A2(n537bar), .ZN(n542bar) );
  OR2_X1 U436 ( .A1(in_14), .A2(in[99]), .ZN(n537) );
  AND2_X1 U436bar ( .A1(in_14bar), .A2(inbar[99]), .ZN(n537bar) );
  OR2_X1 U437 ( .A1(in_60), .A2(in_18), .ZN(n538) );
  AND2_X1 U437bar ( .A1(in_60bar), .A2(in_18bar), .ZN(n538bar) );
  OR2_X1 U438 ( .A1(in[113]), .A2(n763), .ZN(n566) );
  AND2_X1 U438bar ( .A1(inbar[113]), .A2(n763bar), .ZN(n566bar) );
  OR2_X1 U439 ( .A1(n536), .A2(n535), .ZN(n763) );
  AND2_X1 U439bar ( .A1(n536bar), .A2(n535bar), .ZN(n763bar) );
  OR2_X1 U440 ( .A1(n534), .A2(n533), .ZN(n535) );
  AND2_X1 U440bar ( .A1(n534bar), .A2(n533bar), .ZN(n535bar) );
  OR2_X1 U441 ( .A1(n532), .A2(n531), .ZN(n533) );
  AND2_X1 U441bar ( .A1(n532bar), .A2(n531bar), .ZN(n533bar) );
  OR2_X1 U442 ( .A1(in[115]), .A2(in[110]), .ZN(n531) );
  AND2_X1 U442bar ( .A1(inbar[115]), .A2(inbar[110]), .ZN(n531bar) );
  OR2_X1 U443 ( .A1(in[125]), .A2(in[117]), .ZN(n532) );
  AND2_X1 U443bar ( .A1(inbar[125]), .A2(inbar[117]), .ZN(n532bar) );
  OR2_X1 U444 ( .A1(n530), .A2(n529), .ZN(n534) );
  AND2_X1 U444bar ( .A1(n530bar), .A2(n529bar), .ZN(n534bar) );
  OR2_X1 U445 ( .A1(in[180]), .A2(in[128]), .ZN(n529) );
  AND2_X1 U445bar ( .A1(inbar[180]), .A2(inbar[128]), .ZN(n529bar) );
  OR2_X1 U446 ( .A1(in[205]), .A2(in[201]), .ZN(n530) );
  AND2_X1 U446bar ( .A1(inbar[205]), .A2(inbar[201]), .ZN(n530bar) );
  OR2_X1 U447 ( .A1(n528), .A2(n527), .ZN(n536) );
  AND2_X1 U447bar ( .A1(n528bar), .A2(n527bar), .ZN(n536bar) );
  OR2_X1 U448 ( .A1(n526), .A2(n525), .ZN(n527) );
  AND2_X1 U448bar ( .A1(n526bar), .A2(n525bar), .ZN(n527bar) );
  OR2_X1 U449 ( .A1(in[244]), .A2(in[239]), .ZN(n525) );
  AND2_X1 U449bar ( .A1(inbar[244]), .A2(inbar[239]), .ZN(n525bar) );
  OR2_X1 U450 ( .A1(in[95]), .A2(in[83]), .ZN(n526) );
  AND2_X1 U450bar ( .A1(inbar[95]), .A2(inbar[83]), .ZN(n526bar) );
  OR2_X1 U451 ( .A1(n524), .A2(n523), .ZN(n528) );
  AND2_X1 U451bar ( .A1(n524bar), .A2(n523bar), .ZN(n528bar) );
  OR2_X1 U452 ( .A1(in_24), .A2(in[97]), .ZN(n523) );
  AND2_X1 U452bar ( .A1(in_24bar), .A2(inbar[97]), .ZN(n523bar) );
  OR2_X1 U453 ( .A1(in_33), .A2(in_27), .ZN(n524) );
  AND2_X1 U453bar ( .A1(in_33bar), .A2(in_27bar), .ZN(n524bar) );
  OR2_X1 U454 ( .A1(n522), .A2(n521), .ZN(n568) );
  AND2_X1 U454bar ( .A1(n522bar), .A2(n521bar), .ZN(n568bar) );
  OR2_X1 U455 ( .A1(in[145]), .A2(in[126]), .ZN(n521) );
  AND2_X1 U455bar ( .A1(inbar[145]), .A2(inbar[126]), .ZN(n521bar) );
  OR2_X1 U456 ( .A1(in[169]), .A2(n520), .ZN(n522) );
  AND2_X1 U456bar ( .A1(inbar[169]), .A2(n520bar), .ZN(n522bar) );
  OR2_X1 U457 ( .A1(in[221]), .A2(in[172]), .ZN(n520) );
  AND2_X1 U457bar ( .A1(inbar[221]), .A2(inbar[172]), .ZN(n520bar) );
  OR2_X1 U458 ( .A1(n519), .A2(n518), .ZN(n570) );
  AND2_X1 U458bar ( .A1(n519bar), .A2(n518bar), .ZN(n570bar) );
  OR2_X1 U459 ( .A1(n517), .A2(n516), .ZN(n518) );
  AND2_X1 U459bar ( .A1(n517bar), .A2(n516bar), .ZN(n518bar) );
  OR2_X1 U460 ( .A1(in[241]), .A2(in[224]), .ZN(n516) );
  AND2_X1 U460bar ( .A1(inbar[241]), .A2(inbar[224]), .ZN(n516bar) );
  OR2_X1 U461 ( .A1(in[86]), .A2(n515), .ZN(n517) );
  AND2_X1 U461bar ( .A1(inbar[86]), .A2(n515bar), .ZN(n517bar) );
  OR2_X1 U462 ( .A1(in_43), .A2(in_34), .ZN(n515) );
  AND2_X1 U462bar ( .A1(in_43bar), .A2(in_34bar), .ZN(n515bar) );
  OR2_X1 U463 ( .A1(n514), .A2(n513), .ZN(n519) );
  AND2_X1 U463bar ( .A1(n514bar), .A2(n513bar), .ZN(n519bar) );
  OR2_X1 U464 ( .A1(in_65), .A2(in_51), .ZN(n513) );
  AND2_X1 U464bar ( .A1(in_65bar), .A2(in_51bar), .ZN(n513bar) );
  OR2_X1 U465 ( .A1(in_75), .A2(n512), .ZN(n514) );
  AND2_X1 U465bar ( .A1(in_75bar), .A2(n512bar), .ZN(n514bar) );
  OR2_X1 U466 ( .A1(in_81), .A2(in_77), .ZN(n512) );
  AND2_X1 U466bar ( .A1(in_81bar), .A2(in_77bar), .ZN(n512bar) );
  OR2_X1 U467 ( .A1(n511), .A2(n510), .ZN(n778) );
  AND2_X1 U467bar ( .A1(n511bar), .A2(n510bar), .ZN(n778bar) );
  OR2_X1 U468 ( .A1(n509), .A2(n508), .ZN(n510) );
  AND2_X1 U468bar ( .A1(n509bar), .A2(n508bar), .ZN(n510bar) );
  OR2_X1 U469 ( .A1(n507), .A2(n506), .ZN(n508) );
  AND2_X1 U469bar ( .A1(n507bar), .A2(n506bar), .ZN(n508bar) );
  OR2_X1 U470 ( .A1(in[107]), .A2(in[101]), .ZN(n506) );
  AND2_X1 U470bar ( .A1(inbar[107]), .A2(inbar[101]), .ZN(n506bar) );
  OR2_X1 U471 ( .A1(in[139]), .A2(in[132]), .ZN(n507) );
  AND2_X1 U471bar ( .A1(inbar[139]), .A2(inbar[132]), .ZN(n507bar) );
  OR2_X1 U472 ( .A1(n505), .A2(n504), .ZN(n509) );
  AND2_X1 U472bar ( .A1(n505bar), .A2(n504bar), .ZN(n509bar) );
  OR2_X1 U473 ( .A1(in[146]), .A2(in[141]), .ZN(n504) );
  AND2_X1 U473bar ( .A1(inbar[146]), .A2(inbar[141]), .ZN(n504bar) );
  OR2_X1 U474 ( .A1(in[203]), .A2(in[179]), .ZN(n505) );
  AND2_X1 U474bar ( .A1(inbar[203]), .A2(inbar[179]), .ZN(n505bar) );
  OR2_X1 U475 ( .A1(n503), .A2(n502), .ZN(n511) );
  AND2_X1 U475bar ( .A1(n503bar), .A2(n502bar), .ZN(n511bar) );
  OR2_X1 U476 ( .A1(n501), .A2(n500), .ZN(n502) );
  AND2_X1 U476bar ( .A1(n501bar), .A2(n500bar), .ZN(n502bar) );
  OR2_X1 U477 ( .A1(in[243]), .A2(in[222]), .ZN(n500) );
  AND2_X1 U477bar ( .A1(inbar[243]), .A2(inbar[222]), .ZN(n500bar) );
  OR2_X1 U478 ( .A1(in[251]), .A2(in[250]), .ZN(n501) );
  AND2_X1 U478bar ( .A1(inbar[251]), .A2(inbar[250]), .ZN(n501bar) );
  OR2_X1 U479 ( .A1(n499), .A2(n498), .ZN(n503) );
  AND2_X1 U479bar ( .A1(n499bar), .A2(n498bar), .ZN(n503bar) );
  OR2_X1 U480 ( .A1(in_37), .A2(in_19), .ZN(n498) );
  AND2_X1 U480bar ( .A1(in_37bar), .A2(in_19bar), .ZN(n498bar) );
  OR2_X1 U481 ( .A1(in_78), .A2(in_6), .ZN(n499) );
  AND2_X1 U481bar ( .A1(in_78bar), .A2(in_6bar), .ZN(n499bar) );
  OR2_X1 U482 ( .A1(n497), .A2(n496), .ZN(n603) );
  AND2_X1 U482bar ( .A1(n497bar), .A2(n496bar), .ZN(n603bar) );
  OR2_X1 U483 ( .A1(in[112]), .A2(in[102]), .ZN(n496) );
  AND2_X1 U483bar ( .A1(inbar[112]), .A2(inbar[102]), .ZN(n496bar) );
  OR2_X1 U484 ( .A1(in[123]), .A2(n495), .ZN(n497) );
  AND2_X1 U484bar ( .A1(inbar[123]), .A2(n495bar), .ZN(n497bar) );
  OR2_X1 U485 ( .A1(in[143]), .A2(in[130]), .ZN(n495) );
  AND2_X1 U485bar ( .A1(inbar[143]), .A2(inbar[130]), .ZN(n495bar) );
  OR2_X1 U486 ( .A1(n494), .A2(n493), .ZN(n605) );
  AND2_X1 U486bar ( .A1(n494bar), .A2(n493bar), .ZN(n605bar) );
  OR2_X1 U487 ( .A1(n492), .A2(n491), .ZN(n493) );
  AND2_X1 U487bar ( .A1(n492bar), .A2(n491bar), .ZN(n493bar) );
  OR2_X1 U488 ( .A1(in[216]), .A2(in[213]), .ZN(n491) );
  AND2_X1 U488bar ( .A1(inbar[216]), .A2(inbar[213]), .ZN(n491bar) );
  OR2_X1 U489 ( .A1(in[227]), .A2(n490), .ZN(n492) );
  AND2_X1 U489bar ( .A1(inbar[227]), .A2(n490bar), .ZN(n492bar) );
  OR2_X1 U490 ( .A1(in_0), .A2(in[248]), .ZN(n490) );
  AND2_X1 U490bar ( .A1(in_0bar), .A2(inbar[248]), .ZN(n490bar) );
  OR2_X1 U491 ( .A1(n489), .A2(n488), .ZN(n494) );
  AND2_X1 U491bar ( .A1(n489bar), .A2(n488bar), .ZN(n494bar) );
  OR2_X1 U492 ( .A1(in_46), .A2(in_44), .ZN(n488) );
  AND2_X1 U492bar ( .A1(in_46bar), .A2(in_44bar), .ZN(n488bar) );
  OR2_X1 U493 ( .A1(in_50), .A2(n487), .ZN(n489) );
  AND2_X1 U493bar ( .A1(in_50bar), .A2(n487bar), .ZN(n489bar) );
  OR2_X1 U494 ( .A1(in_9), .A2(in_80), .ZN(n487) );
  AND2_X1 U494bar ( .A1(in_9bar), .A2(in_80bar), .ZN(n487bar) );
endmodule

module sBox_8 ( in, inbar, out, outbar );

  input wire [7:0] in;
  input wire [7:0] inbar;
//input_done

  output wire [7:0] out;
  output wire [7:0] outbar;
//output_done

  wire [255:0] decodeOut;
  wire [255:0] decodeOutbar;
//wire_done

  decode_8 dec ( .in(in), .inbar(inbar), .out(decodeOut), .outbar(decodeOutbar) );
  encode_8 enc ( .in(decodeOut), .inbar(decodeOutbar), .out(out), .outbar(outbar) );
endmodule

module CD2_33 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD2_34 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD2_35 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD2_36 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD4_17 ( a, abar, b, bbar, y, ybar );

  input wire [3:0] a;
  input wire [3:0] b;
  input wire [3:0] abar;
  input wire [3:0] bbar;
//input_done

  output wire [15:0] y;
  output wire [15:0] ybar;
//output_done

//wire_done

  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]) );
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]) );
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]) );
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]) );
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]) );
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]) );
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]) );
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]) );
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]) );
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]) );
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]) );
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]) );
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]) );
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]) );
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]) );
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]) );
endmodule

module CD4_18 ( a, abar, b, bbar, y, ybar );

  input wire [3:0] a;
  input wire [3:0] b;
  input wire [3:0] abar;
  input wire [3:0] bbar;
//input_done

  output wire [15:0] y;
  output wire [15:0] ybar;
//output_done

//wire_done

  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]) );
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]) );
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]) );
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]) );
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]) );
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]) );
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]) );
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]) );
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]) );
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]) );
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]) );
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]) );
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]) );
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]) );
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]) );
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]) );
endmodule

module CD16_9 ( a, abar, b, bbar, y, ybar );

  input wire [15:0] a;
  input wire [15:0] b;
  input wire [15:0] abar;
  input wire [15:0] bbar;
//input_done

  output wire [255:0] y;
  output wire [255:0] ybar;
//output_done

//wire_done

  AND2_X1 U1 ( .A1(b[9]), .A2(a[0]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[9]), .A2(abar[0]), .ZN(ybar[9]) );
  AND2_X1 U2 ( .A1(b[3]), .A2(a[6]), .ZN(y[99]) );
  OR2_X1 U2bar ( .A1(bbar[3]), .A2(abar[6]), .ZN(ybar[99]) );
  AND2_X1 U3 ( .A1(b[2]), .A2(a[6]), .ZN(y[98]) );
  OR2_X1 U3bar ( .A1(bbar[2]), .A2(abar[6]), .ZN(ybar[98]) );
  AND2_X1 U4 ( .A1(b[1]), .A2(a[6]), .ZN(y[97]) );
  OR2_X1 U4bar ( .A1(bbar[1]), .A2(abar[6]), .ZN(ybar[97]) );
  AND2_X1 U5 ( .A1(b[0]), .A2(a[6]), .ZN(y[96]) );
  OR2_X1 U5bar ( .A1(bbar[0]), .A2(abar[6]), .ZN(ybar[96]) );
  AND2_X1 U6 ( .A1(b[15]), .A2(a[5]), .ZN(y[95]) );
  OR2_X1 U6bar ( .A1(bbar[15]), .A2(abar[5]), .ZN(ybar[95]) );
  AND2_X1 U7 ( .A1(b[14]), .A2(a[5]), .ZN(y[94]) );
  OR2_X1 U7bar ( .A1(bbar[14]), .A2(abar[5]), .ZN(ybar[94]) );
  AND2_X1 U8 ( .A1(b[13]), .A2(a[5]), .ZN(y[93]) );
  OR2_X1 U8bar ( .A1(bbar[13]), .A2(abar[5]), .ZN(ybar[93]) );
  AND2_X1 U9 ( .A1(b[12]), .A2(a[5]), .ZN(y[92]) );
  OR2_X1 U9bar ( .A1(bbar[12]), .A2(abar[5]), .ZN(ybar[92]) );
  AND2_X1 U10 ( .A1(b[11]), .A2(a[5]), .ZN(y[91]) );
  OR2_X1 U10bar ( .A1(bbar[11]), .A2(abar[5]), .ZN(ybar[91]) );
  AND2_X1 U11 ( .A1(b[10]), .A2(a[5]), .ZN(y[90]) );
  OR2_X1 U11bar ( .A1(bbar[10]), .A2(abar[5]), .ZN(ybar[90]) );
  AND2_X1 U12 ( .A1(b[8]), .A2(a[0]), .ZN(y[8]) );
  OR2_X1 U12bar ( .A1(bbar[8]), .A2(abar[0]), .ZN(ybar[8]) );
  AND2_X1 U13 ( .A1(a[5]), .A2(b[9]), .ZN(y[89]) );
  OR2_X1 U13bar ( .A1(abar[5]), .A2(bbar[9]), .ZN(ybar[89]) );
  AND2_X1 U14 ( .A1(b[8]), .A2(a[5]), .ZN(y[88]) );
  OR2_X1 U14bar ( .A1(bbar[8]), .A2(abar[5]), .ZN(ybar[88]) );
  AND2_X1 U15 ( .A1(b[7]), .A2(a[5]), .ZN(y[87]) );
  OR2_X1 U15bar ( .A1(bbar[7]), .A2(abar[5]), .ZN(ybar[87]) );
  AND2_X1 U16 ( .A1(b[6]), .A2(a[5]), .ZN(y[86]) );
  OR2_X1 U16bar ( .A1(bbar[6]), .A2(abar[5]), .ZN(ybar[86]) );
  AND2_X1 U17 ( .A1(b[5]), .A2(a[5]), .ZN(y[85]) );
  OR2_X1 U17bar ( .A1(bbar[5]), .A2(abar[5]), .ZN(ybar[85]) );
  AND2_X1 U18 ( .A1(b[4]), .A2(a[5]), .ZN(y[84]) );
  OR2_X1 U18bar ( .A1(bbar[4]), .A2(abar[5]), .ZN(ybar[84]) );
  AND2_X1 U19 ( .A1(a[5]), .A2(b[3]), .ZN(y[83]) );
  OR2_X1 U19bar ( .A1(abar[5]), .A2(bbar[3]), .ZN(ybar[83]) );
  AND2_X1 U20 ( .A1(a[5]), .A2(b[2]), .ZN(y[82]) );
  OR2_X1 U20bar ( .A1(abar[5]), .A2(bbar[2]), .ZN(ybar[82]) );
  AND2_X1 U21 ( .A1(a[5]), .A2(b[1]), .ZN(y[81]) );
  OR2_X1 U21bar ( .A1(abar[5]), .A2(bbar[1]), .ZN(ybar[81]) );
  AND2_X1 U22 ( .A1(a[5]), .A2(b[0]), .ZN(y[80]) );
  OR2_X1 U22bar ( .A1(abar[5]), .A2(bbar[0]), .ZN(ybar[80]) );
  AND2_X1 U23 ( .A1(b[7]), .A2(a[0]), .ZN(y[7]) );
  OR2_X1 U23bar ( .A1(bbar[7]), .A2(abar[0]), .ZN(ybar[7]) );
  AND2_X1 U24 ( .A1(a[4]), .A2(b[15]), .ZN(y[79]) );
  OR2_X1 U24bar ( .A1(abar[4]), .A2(bbar[15]), .ZN(ybar[79]) );
  AND2_X1 U25 ( .A1(a[4]), .A2(b[14]), .ZN(y[78]) );
  OR2_X1 U25bar ( .A1(abar[4]), .A2(bbar[14]), .ZN(ybar[78]) );
  AND2_X1 U26 ( .A1(a[4]), .A2(b[13]), .ZN(y[77]) );
  OR2_X1 U26bar ( .A1(abar[4]), .A2(bbar[13]), .ZN(ybar[77]) );
  AND2_X1 U27 ( .A1(a[4]), .A2(b[12]), .ZN(y[76]) );
  OR2_X1 U27bar ( .A1(abar[4]), .A2(bbar[12]), .ZN(ybar[76]) );
  AND2_X1 U28 ( .A1(a[4]), .A2(b[11]), .ZN(y[75]) );
  OR2_X1 U28bar ( .A1(abar[4]), .A2(bbar[11]), .ZN(ybar[75]) );
  AND2_X1 U29 ( .A1(a[4]), .A2(b[10]), .ZN(y[74]) );
  OR2_X1 U29bar ( .A1(abar[4]), .A2(bbar[10]), .ZN(ybar[74]) );
  AND2_X1 U30 ( .A1(a[4]), .A2(b[9]), .ZN(y[73]) );
  OR2_X1 U30bar ( .A1(abar[4]), .A2(bbar[9]), .ZN(ybar[73]) );
  AND2_X1 U31 ( .A1(a[4]), .A2(b[8]), .ZN(y[72]) );
  OR2_X1 U31bar ( .A1(abar[4]), .A2(bbar[8]), .ZN(ybar[72]) );
  AND2_X1 U32 ( .A1(a[4]), .A2(b[7]), .ZN(y[71]) );
  OR2_X1 U32bar ( .A1(abar[4]), .A2(bbar[7]), .ZN(ybar[71]) );
  AND2_X1 U33 ( .A1(a[4]), .A2(b[6]), .ZN(y[70]) );
  OR2_X1 U33bar ( .A1(abar[4]), .A2(bbar[6]), .ZN(ybar[70]) );
  AND2_X1 U34 ( .A1(b[6]), .A2(a[0]), .ZN(y[6]) );
  OR2_X1 U34bar ( .A1(bbar[6]), .A2(abar[0]), .ZN(ybar[6]) );
  AND2_X1 U35 ( .A1(a[4]), .A2(b[5]), .ZN(y[69]) );
  OR2_X1 U35bar ( .A1(abar[4]), .A2(bbar[5]), .ZN(ybar[69]) );
  AND2_X1 U36 ( .A1(a[4]), .A2(b[4]), .ZN(y[68]) );
  OR2_X1 U36bar ( .A1(abar[4]), .A2(bbar[4]), .ZN(ybar[68]) );
  AND2_X1 U37 ( .A1(a[4]), .A2(b[3]), .ZN(y[67]) );
  OR2_X1 U37bar ( .A1(abar[4]), .A2(bbar[3]), .ZN(ybar[67]) );
  AND2_X1 U38 ( .A1(a[4]), .A2(b[2]), .ZN(y[66]) );
  OR2_X1 U38bar ( .A1(abar[4]), .A2(bbar[2]), .ZN(ybar[66]) );
  AND2_X1 U39 ( .A1(a[4]), .A2(b[1]), .ZN(y[65]) );
  OR2_X1 U39bar ( .A1(abar[4]), .A2(bbar[1]), .ZN(ybar[65]) );
  AND2_X1 U40 ( .A1(a[4]), .A2(b[0]), .ZN(y[64]) );
  OR2_X1 U40bar ( .A1(abar[4]), .A2(bbar[0]), .ZN(ybar[64]) );
  AND2_X1 U41 ( .A1(a[3]), .A2(b[15]), .ZN(y[63]) );
  OR2_X1 U41bar ( .A1(abar[3]), .A2(bbar[15]), .ZN(ybar[63]) );
  AND2_X1 U42 ( .A1(a[3]), .A2(b[14]), .ZN(y[62]) );
  OR2_X1 U42bar ( .A1(abar[3]), .A2(bbar[14]), .ZN(ybar[62]) );
  AND2_X1 U43 ( .A1(a[3]), .A2(b[13]), .ZN(y[61]) );
  OR2_X1 U43bar ( .A1(abar[3]), .A2(bbar[13]), .ZN(ybar[61]) );
  AND2_X1 U44 ( .A1(a[3]), .A2(b[12]), .ZN(y[60]) );
  OR2_X1 U44bar ( .A1(abar[3]), .A2(bbar[12]), .ZN(ybar[60]) );
  AND2_X1 U45 ( .A1(b[5]), .A2(a[0]), .ZN(y[5]) );
  OR2_X1 U45bar ( .A1(bbar[5]), .A2(abar[0]), .ZN(ybar[5]) );
  AND2_X1 U46 ( .A1(a[3]), .A2(b[11]), .ZN(y[59]) );
  OR2_X1 U46bar ( .A1(abar[3]), .A2(bbar[11]), .ZN(ybar[59]) );
  AND2_X1 U47 ( .A1(a[3]), .A2(b[10]), .ZN(y[58]) );
  OR2_X1 U47bar ( .A1(abar[3]), .A2(bbar[10]), .ZN(ybar[58]) );
  AND2_X1 U48 ( .A1(a[3]), .A2(b[9]), .ZN(y[57]) );
  OR2_X1 U48bar ( .A1(abar[3]), .A2(bbar[9]), .ZN(ybar[57]) );
  AND2_X1 U49 ( .A1(a[3]), .A2(b[8]), .ZN(y[56]) );
  OR2_X1 U49bar ( .A1(abar[3]), .A2(bbar[8]), .ZN(ybar[56]) );
  AND2_X1 U50 ( .A1(a[3]), .A2(b[7]), .ZN(y[55]) );
  OR2_X1 U50bar ( .A1(abar[3]), .A2(bbar[7]), .ZN(ybar[55]) );
  AND2_X1 U51 ( .A1(a[3]), .A2(b[6]), .ZN(y[54]) );
  OR2_X1 U51bar ( .A1(abar[3]), .A2(bbar[6]), .ZN(ybar[54]) );
  AND2_X1 U52 ( .A1(a[3]), .A2(b[5]), .ZN(y[53]) );
  OR2_X1 U52bar ( .A1(abar[3]), .A2(bbar[5]), .ZN(ybar[53]) );
  AND2_X1 U53 ( .A1(a[3]), .A2(b[4]), .ZN(y[52]) );
  OR2_X1 U53bar ( .A1(abar[3]), .A2(bbar[4]), .ZN(ybar[52]) );
  AND2_X1 U54 ( .A1(a[3]), .A2(b[3]), .ZN(y[51]) );
  OR2_X1 U54bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[51]) );
  AND2_X1 U55 ( .A1(a[3]), .A2(b[2]), .ZN(y[50]) );
  OR2_X1 U55bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[50]) );
  AND2_X1 U56 ( .A1(b[4]), .A2(a[0]), .ZN(y[4]) );
  OR2_X1 U56bar ( .A1(bbar[4]), .A2(abar[0]), .ZN(ybar[4]) );
  AND2_X1 U57 ( .A1(a[3]), .A2(b[1]), .ZN(y[49]) );
  OR2_X1 U57bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[49]) );
  AND2_X1 U58 ( .A1(a[3]), .A2(b[0]), .ZN(y[48]) );
  OR2_X1 U58bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[48]) );
  AND2_X1 U59 ( .A1(a[2]), .A2(b[15]), .ZN(y[47]) );
  OR2_X1 U59bar ( .A1(abar[2]), .A2(bbar[15]), .ZN(ybar[47]) );
  AND2_X1 U60 ( .A1(a[2]), .A2(b[14]), .ZN(y[46]) );
  OR2_X1 U60bar ( .A1(abar[2]), .A2(bbar[14]), .ZN(ybar[46]) );
  AND2_X1 U61 ( .A1(a[2]), .A2(b[13]), .ZN(y[45]) );
  OR2_X1 U61bar ( .A1(abar[2]), .A2(bbar[13]), .ZN(ybar[45]) );
  AND2_X1 U62 ( .A1(a[2]), .A2(b[12]), .ZN(y[44]) );
  OR2_X1 U62bar ( .A1(abar[2]), .A2(bbar[12]), .ZN(ybar[44]) );
  AND2_X1 U63 ( .A1(a[2]), .A2(b[11]), .ZN(y[43]) );
  OR2_X1 U63bar ( .A1(abar[2]), .A2(bbar[11]), .ZN(ybar[43]) );
  AND2_X1 U64 ( .A1(a[2]), .A2(b[10]), .ZN(y[42]) );
  OR2_X1 U64bar ( .A1(abar[2]), .A2(bbar[10]), .ZN(ybar[42]) );
  AND2_X1 U65 ( .A1(a[2]), .A2(b[9]), .ZN(y[41]) );
  OR2_X1 U65bar ( .A1(abar[2]), .A2(bbar[9]), .ZN(ybar[41]) );
  AND2_X1 U66 ( .A1(a[2]), .A2(b[8]), .ZN(y[40]) );
  OR2_X1 U66bar ( .A1(abar[2]), .A2(bbar[8]), .ZN(ybar[40]) );
  AND2_X1 U67 ( .A1(b[3]), .A2(a[0]), .ZN(y[3]) );
  OR2_X1 U67bar ( .A1(bbar[3]), .A2(abar[0]), .ZN(ybar[3]) );
  AND2_X1 U68 ( .A1(a[2]), .A2(b[7]), .ZN(y[39]) );
  OR2_X1 U68bar ( .A1(abar[2]), .A2(bbar[7]), .ZN(ybar[39]) );
  AND2_X1 U69 ( .A1(a[2]), .A2(b[6]), .ZN(y[38]) );
  OR2_X1 U69bar ( .A1(abar[2]), .A2(bbar[6]), .ZN(ybar[38]) );
  AND2_X1 U70 ( .A1(a[2]), .A2(b[5]), .ZN(y[37]) );
  OR2_X1 U70bar ( .A1(abar[2]), .A2(bbar[5]), .ZN(ybar[37]) );
  AND2_X1 U71 ( .A1(a[2]), .A2(b[4]), .ZN(y[36]) );
  OR2_X1 U71bar ( .A1(abar[2]), .A2(bbar[4]), .ZN(ybar[36]) );
  AND2_X1 U72 ( .A1(a[2]), .A2(b[3]), .ZN(y[35]) );
  OR2_X1 U72bar ( .A1(abar[2]), .A2(bbar[3]), .ZN(ybar[35]) );
  AND2_X1 U73 ( .A1(a[2]), .A2(b[2]), .ZN(y[34]) );
  OR2_X1 U73bar ( .A1(abar[2]), .A2(bbar[2]), .ZN(ybar[34]) );
  AND2_X1 U74 ( .A1(a[2]), .A2(b[1]), .ZN(y[33]) );
  OR2_X1 U74bar ( .A1(abar[2]), .A2(bbar[1]), .ZN(ybar[33]) );
  AND2_X1 U75 ( .A1(a[2]), .A2(b[0]), .ZN(y[32]) );
  OR2_X1 U75bar ( .A1(abar[2]), .A2(bbar[0]), .ZN(ybar[32]) );
  AND2_X1 U76 ( .A1(a[1]), .A2(b[15]), .ZN(y[31]) );
  OR2_X1 U76bar ( .A1(abar[1]), .A2(bbar[15]), .ZN(ybar[31]) );
  AND2_X1 U77 ( .A1(a[1]), .A2(b[14]), .ZN(y[30]) );
  OR2_X1 U77bar ( .A1(abar[1]), .A2(bbar[14]), .ZN(ybar[30]) );
  AND2_X1 U78 ( .A1(b[2]), .A2(a[0]), .ZN(y[2]) );
  OR2_X1 U78bar ( .A1(bbar[2]), .A2(abar[0]), .ZN(ybar[2]) );
  AND2_X1 U79 ( .A1(a[1]), .A2(b[13]), .ZN(y[29]) );
  OR2_X1 U79bar ( .A1(abar[1]), .A2(bbar[13]), .ZN(ybar[29]) );
  AND2_X1 U80 ( .A1(a[1]), .A2(b[12]), .ZN(y[28]) );
  OR2_X1 U80bar ( .A1(abar[1]), .A2(bbar[12]), .ZN(ybar[28]) );
  AND2_X1 U81 ( .A1(a[1]), .A2(b[11]), .ZN(y[27]) );
  OR2_X1 U81bar ( .A1(abar[1]), .A2(bbar[11]), .ZN(ybar[27]) );
  AND2_X1 U82 ( .A1(a[1]), .A2(b[10]), .ZN(y[26]) );
  OR2_X1 U82bar ( .A1(abar[1]), .A2(bbar[10]), .ZN(ybar[26]) );
  AND2_X1 U83 ( .A1(a[1]), .A2(b[9]), .ZN(y[25]) );
  OR2_X1 U83bar ( .A1(abar[1]), .A2(bbar[9]), .ZN(ybar[25]) );
  AND2_X1 U84 ( .A1(a[15]), .A2(b[15]), .ZN(y[255]) );
  OR2_X1 U84bar ( .A1(abar[15]), .A2(bbar[15]), .ZN(ybar[255]) );
  AND2_X1 U85 ( .A1(a[15]), .A2(b[14]), .ZN(y[254]) );
  OR2_X1 U85bar ( .A1(abar[15]), .A2(bbar[14]), .ZN(ybar[254]) );
  AND2_X1 U86 ( .A1(a[15]), .A2(b[13]), .ZN(y[253]) );
  OR2_X1 U86bar ( .A1(abar[15]), .A2(bbar[13]), .ZN(ybar[253]) );
  AND2_X1 U87 ( .A1(a[15]), .A2(b[12]), .ZN(y[252]) );
  OR2_X1 U87bar ( .A1(abar[15]), .A2(bbar[12]), .ZN(ybar[252]) );
  AND2_X1 U88 ( .A1(a[15]), .A2(b[11]), .ZN(y[251]) );
  OR2_X1 U88bar ( .A1(abar[15]), .A2(bbar[11]), .ZN(ybar[251]) );
  AND2_X1 U89 ( .A1(a[15]), .A2(b[10]), .ZN(y[250]) );
  OR2_X1 U89bar ( .A1(abar[15]), .A2(bbar[10]), .ZN(ybar[250]) );
  AND2_X1 U90 ( .A1(a[1]), .A2(b[8]), .ZN(y[24]) );
  OR2_X1 U90bar ( .A1(abar[1]), .A2(bbar[8]), .ZN(ybar[24]) );
  AND2_X1 U91 ( .A1(a[15]), .A2(b[9]), .ZN(y[249]) );
  OR2_X1 U91bar ( .A1(abar[15]), .A2(bbar[9]), .ZN(ybar[249]) );
  AND2_X1 U92 ( .A1(a[15]), .A2(b[8]), .ZN(y[248]) );
  OR2_X1 U92bar ( .A1(abar[15]), .A2(bbar[8]), .ZN(ybar[248]) );
  AND2_X1 U93 ( .A1(a[15]), .A2(b[7]), .ZN(y[247]) );
  OR2_X1 U93bar ( .A1(abar[15]), .A2(bbar[7]), .ZN(ybar[247]) );
  AND2_X1 U94 ( .A1(a[15]), .A2(b[6]), .ZN(y[246]) );
  OR2_X1 U94bar ( .A1(abar[15]), .A2(bbar[6]), .ZN(ybar[246]) );
  AND2_X1 U95 ( .A1(a[15]), .A2(b[5]), .ZN(y[245]) );
  OR2_X1 U95bar ( .A1(abar[15]), .A2(bbar[5]), .ZN(ybar[245]) );
  AND2_X1 U96 ( .A1(a[15]), .A2(b[4]), .ZN(y[244]) );
  OR2_X1 U96bar ( .A1(abar[15]), .A2(bbar[4]), .ZN(ybar[244]) );
  AND2_X1 U97 ( .A1(a[15]), .A2(b[3]), .ZN(y[243]) );
  OR2_X1 U97bar ( .A1(abar[15]), .A2(bbar[3]), .ZN(ybar[243]) );
  AND2_X1 U98 ( .A1(a[15]), .A2(b[2]), .ZN(y[242]) );
  OR2_X1 U98bar ( .A1(abar[15]), .A2(bbar[2]), .ZN(ybar[242]) );
  AND2_X1 U99 ( .A1(a[15]), .A2(b[1]), .ZN(y[241]) );
  OR2_X1 U99bar ( .A1(abar[15]), .A2(bbar[1]), .ZN(ybar[241]) );
  AND2_X1 U100 ( .A1(a[15]), .A2(b[0]), .ZN(y[240]) );
  OR2_X1 U100bar ( .A1(abar[15]), .A2(bbar[0]), .ZN(ybar[240]) );
  AND2_X1 U101 ( .A1(a[1]), .A2(b[7]), .ZN(y[23]) );
  OR2_X1 U101bar ( .A1(abar[1]), .A2(bbar[7]), .ZN(ybar[23]) );
  AND2_X1 U102 ( .A1(a[14]), .A2(b[15]), .ZN(y[239]) );
  OR2_X1 U102bar ( .A1(abar[14]), .A2(bbar[15]), .ZN(ybar[239]) );
  AND2_X1 U103 ( .A1(a[14]), .A2(b[14]), .ZN(y[238]) );
  OR2_X1 U103bar ( .A1(abar[14]), .A2(bbar[14]), .ZN(ybar[238]) );
  AND2_X1 U104 ( .A1(a[14]), .A2(b[13]), .ZN(y[237]) );
  OR2_X1 U104bar ( .A1(abar[14]), .A2(bbar[13]), .ZN(ybar[237]) );
  AND2_X1 U105 ( .A1(a[14]), .A2(b[12]), .ZN(y[236]) );
  OR2_X1 U105bar ( .A1(abar[14]), .A2(bbar[12]), .ZN(ybar[236]) );
  AND2_X1 U106 ( .A1(a[14]), .A2(b[11]), .ZN(y[235]) );
  OR2_X1 U106bar ( .A1(abar[14]), .A2(bbar[11]), .ZN(ybar[235]) );
  AND2_X1 U107 ( .A1(a[14]), .A2(b[10]), .ZN(y[234]) );
  OR2_X1 U107bar ( .A1(abar[14]), .A2(bbar[10]), .ZN(ybar[234]) );
  AND2_X1 U108 ( .A1(a[14]), .A2(b[9]), .ZN(y[233]) );
  OR2_X1 U108bar ( .A1(abar[14]), .A2(bbar[9]), .ZN(ybar[233]) );
  AND2_X1 U109 ( .A1(a[14]), .A2(b[8]), .ZN(y[232]) );
  OR2_X1 U109bar ( .A1(abar[14]), .A2(bbar[8]), .ZN(ybar[232]) );
  AND2_X1 U110 ( .A1(a[14]), .A2(b[7]), .ZN(y[231]) );
  OR2_X1 U110bar ( .A1(abar[14]), .A2(bbar[7]), .ZN(ybar[231]) );
  AND2_X1 U111 ( .A1(a[14]), .A2(b[6]), .ZN(y[230]) );
  OR2_X1 U111bar ( .A1(abar[14]), .A2(bbar[6]), .ZN(ybar[230]) );
  AND2_X1 U112 ( .A1(a[1]), .A2(b[6]), .ZN(y[22]) );
  OR2_X1 U112bar ( .A1(abar[1]), .A2(bbar[6]), .ZN(ybar[22]) );
  AND2_X1 U113 ( .A1(a[14]), .A2(b[5]), .ZN(y[229]) );
  OR2_X1 U113bar ( .A1(abar[14]), .A2(bbar[5]), .ZN(ybar[229]) );
  AND2_X1 U114 ( .A1(a[14]), .A2(b[4]), .ZN(y[228]) );
  OR2_X1 U114bar ( .A1(abar[14]), .A2(bbar[4]), .ZN(ybar[228]) );
  AND2_X1 U115 ( .A1(a[14]), .A2(b[3]), .ZN(y[227]) );
  OR2_X1 U115bar ( .A1(abar[14]), .A2(bbar[3]), .ZN(ybar[227]) );
  AND2_X1 U116 ( .A1(a[14]), .A2(b[2]), .ZN(y[226]) );
  OR2_X1 U116bar ( .A1(abar[14]), .A2(bbar[2]), .ZN(ybar[226]) );
  AND2_X1 U117 ( .A1(a[14]), .A2(b[1]), .ZN(y[225]) );
  OR2_X1 U117bar ( .A1(abar[14]), .A2(bbar[1]), .ZN(ybar[225]) );
  AND2_X1 U118 ( .A1(a[14]), .A2(b[0]), .ZN(y[224]) );
  OR2_X1 U118bar ( .A1(abar[14]), .A2(bbar[0]), .ZN(ybar[224]) );
  AND2_X1 U119 ( .A1(a[13]), .A2(b[15]), .ZN(y[223]) );
  OR2_X1 U119bar ( .A1(abar[13]), .A2(bbar[15]), .ZN(ybar[223]) );
  AND2_X1 U120 ( .A1(a[13]), .A2(b[14]), .ZN(y[222]) );
  OR2_X1 U120bar ( .A1(abar[13]), .A2(bbar[14]), .ZN(ybar[222]) );
  AND2_X1 U121 ( .A1(a[13]), .A2(b[13]), .ZN(y[221]) );
  OR2_X1 U121bar ( .A1(abar[13]), .A2(bbar[13]), .ZN(ybar[221]) );
  AND2_X1 U122 ( .A1(a[13]), .A2(b[12]), .ZN(y[220]) );
  OR2_X1 U122bar ( .A1(abar[13]), .A2(bbar[12]), .ZN(ybar[220]) );
  AND2_X1 U123 ( .A1(a[1]), .A2(b[5]), .ZN(y[21]) );
  OR2_X1 U123bar ( .A1(abar[1]), .A2(bbar[5]), .ZN(ybar[21]) );
  AND2_X1 U124 ( .A1(a[13]), .A2(b[11]), .ZN(y[219]) );
  OR2_X1 U124bar ( .A1(abar[13]), .A2(bbar[11]), .ZN(ybar[219]) );
  AND2_X1 U125 ( .A1(a[13]), .A2(b[10]), .ZN(y[218]) );
  OR2_X1 U125bar ( .A1(abar[13]), .A2(bbar[10]), .ZN(ybar[218]) );
  AND2_X1 U126 ( .A1(a[13]), .A2(b[9]), .ZN(y[217]) );
  OR2_X1 U126bar ( .A1(abar[13]), .A2(bbar[9]), .ZN(ybar[217]) );
  AND2_X1 U127 ( .A1(a[13]), .A2(b[8]), .ZN(y[216]) );
  OR2_X1 U127bar ( .A1(abar[13]), .A2(bbar[8]), .ZN(ybar[216]) );
  AND2_X1 U128 ( .A1(a[13]), .A2(b[7]), .ZN(y[215]) );
  OR2_X1 U128bar ( .A1(abar[13]), .A2(bbar[7]), .ZN(ybar[215]) );
  AND2_X1 U129 ( .A1(a[13]), .A2(b[6]), .ZN(y[214]) );
  OR2_X1 U129bar ( .A1(abar[13]), .A2(bbar[6]), .ZN(ybar[214]) );
  AND2_X1 U130 ( .A1(a[13]), .A2(b[5]), .ZN(y[213]) );
  OR2_X1 U130bar ( .A1(abar[13]), .A2(bbar[5]), .ZN(ybar[213]) );
  AND2_X1 U131 ( .A1(a[13]), .A2(b[4]), .ZN(y[212]) );
  OR2_X1 U131bar ( .A1(abar[13]), .A2(bbar[4]), .ZN(ybar[212]) );
  AND2_X1 U132 ( .A1(a[13]), .A2(b[3]), .ZN(y[211]) );
  OR2_X1 U132bar ( .A1(abar[13]), .A2(bbar[3]), .ZN(ybar[211]) );
  AND2_X1 U133 ( .A1(a[13]), .A2(b[2]), .ZN(y[210]) );
  OR2_X1 U133bar ( .A1(abar[13]), .A2(bbar[2]), .ZN(ybar[210]) );
  AND2_X1 U134 ( .A1(a[1]), .A2(b[4]), .ZN(y[20]) );
  OR2_X1 U134bar ( .A1(abar[1]), .A2(bbar[4]), .ZN(ybar[20]) );
  AND2_X1 U135 ( .A1(a[13]), .A2(b[1]), .ZN(y[209]) );
  OR2_X1 U135bar ( .A1(abar[13]), .A2(bbar[1]), .ZN(ybar[209]) );
  AND2_X1 U136 ( .A1(a[13]), .A2(b[0]), .ZN(y[208]) );
  OR2_X1 U136bar ( .A1(abar[13]), .A2(bbar[0]), .ZN(ybar[208]) );
  AND2_X1 U137 ( .A1(a[12]), .A2(b[15]), .ZN(y[207]) );
  OR2_X1 U137bar ( .A1(abar[12]), .A2(bbar[15]), .ZN(ybar[207]) );
  AND2_X1 U138 ( .A1(a[12]), .A2(b[14]), .ZN(y[206]) );
  OR2_X1 U138bar ( .A1(abar[12]), .A2(bbar[14]), .ZN(ybar[206]) );
  AND2_X1 U139 ( .A1(a[12]), .A2(b[13]), .ZN(y[205]) );
  OR2_X1 U139bar ( .A1(abar[12]), .A2(bbar[13]), .ZN(ybar[205]) );
  AND2_X1 U140 ( .A1(a[12]), .A2(b[12]), .ZN(y[204]) );
  OR2_X1 U140bar ( .A1(abar[12]), .A2(bbar[12]), .ZN(ybar[204]) );
  AND2_X1 U141 ( .A1(a[12]), .A2(b[11]), .ZN(y[203]) );
  OR2_X1 U141bar ( .A1(abar[12]), .A2(bbar[11]), .ZN(ybar[203]) );
  AND2_X1 U142 ( .A1(a[12]), .A2(b[10]), .ZN(y[202]) );
  OR2_X1 U142bar ( .A1(abar[12]), .A2(bbar[10]), .ZN(ybar[202]) );
  AND2_X1 U143 ( .A1(a[12]), .A2(b[9]), .ZN(y[201]) );
  OR2_X1 U143bar ( .A1(abar[12]), .A2(bbar[9]), .ZN(ybar[201]) );
  AND2_X1 U144 ( .A1(a[12]), .A2(b[8]), .ZN(y[200]) );
  OR2_X1 U144bar ( .A1(abar[12]), .A2(bbar[8]), .ZN(ybar[200]) );
  AND2_X1 U145 ( .A1(b[1]), .A2(a[0]), .ZN(y[1]) );
  OR2_X1 U145bar ( .A1(bbar[1]), .A2(abar[0]), .ZN(ybar[1]) );
  AND2_X1 U146 ( .A1(a[1]), .A2(b[3]), .ZN(y[19]) );
  OR2_X1 U146bar ( .A1(abar[1]), .A2(bbar[3]), .ZN(ybar[19]) );
  AND2_X1 U147 ( .A1(a[12]), .A2(b[7]), .ZN(y[199]) );
  OR2_X1 U147bar ( .A1(abar[12]), .A2(bbar[7]), .ZN(ybar[199]) );
  AND2_X1 U148 ( .A1(a[12]), .A2(b[6]), .ZN(y[198]) );
  OR2_X1 U148bar ( .A1(abar[12]), .A2(bbar[6]), .ZN(ybar[198]) );
  AND2_X1 U149 ( .A1(a[12]), .A2(b[5]), .ZN(y[197]) );
  OR2_X1 U149bar ( .A1(abar[12]), .A2(bbar[5]), .ZN(ybar[197]) );
  AND2_X1 U150 ( .A1(a[12]), .A2(b[4]), .ZN(y[196]) );
  OR2_X1 U150bar ( .A1(abar[12]), .A2(bbar[4]), .ZN(ybar[196]) );
  AND2_X1 U151 ( .A1(a[12]), .A2(b[3]), .ZN(y[195]) );
  OR2_X1 U151bar ( .A1(abar[12]), .A2(bbar[3]), .ZN(ybar[195]) );
  AND2_X1 U152 ( .A1(a[12]), .A2(b[2]), .ZN(y[194]) );
  OR2_X1 U152bar ( .A1(abar[12]), .A2(bbar[2]), .ZN(ybar[194]) );
  AND2_X1 U153 ( .A1(a[12]), .A2(b[1]), .ZN(y[193]) );
  OR2_X1 U153bar ( .A1(abar[12]), .A2(bbar[1]), .ZN(ybar[193]) );
  AND2_X1 U154 ( .A1(a[12]), .A2(b[0]), .ZN(y[192]) );
  OR2_X1 U154bar ( .A1(abar[12]), .A2(bbar[0]), .ZN(ybar[192]) );
  AND2_X1 U155 ( .A1(a[11]), .A2(b[15]), .ZN(y[191]) );
  OR2_X1 U155bar ( .A1(abar[11]), .A2(bbar[15]), .ZN(ybar[191]) );
  AND2_X1 U156 ( .A1(a[11]), .A2(b[14]), .ZN(y[190]) );
  OR2_X1 U156bar ( .A1(abar[11]), .A2(bbar[14]), .ZN(ybar[190]) );
  AND2_X1 U157 ( .A1(a[1]), .A2(b[2]), .ZN(y[18]) );
  OR2_X1 U157bar ( .A1(abar[1]), .A2(bbar[2]), .ZN(ybar[18]) );
  AND2_X1 U158 ( .A1(a[11]), .A2(b[13]), .ZN(y[189]) );
  OR2_X1 U158bar ( .A1(abar[11]), .A2(bbar[13]), .ZN(ybar[189]) );
  AND2_X1 U159 ( .A1(a[11]), .A2(b[12]), .ZN(y[188]) );
  OR2_X1 U159bar ( .A1(abar[11]), .A2(bbar[12]), .ZN(ybar[188]) );
  AND2_X1 U160 ( .A1(a[11]), .A2(b[11]), .ZN(y[187]) );
  OR2_X1 U160bar ( .A1(abar[11]), .A2(bbar[11]), .ZN(ybar[187]) );
  AND2_X1 U161 ( .A1(a[11]), .A2(b[10]), .ZN(y[186]) );
  OR2_X1 U161bar ( .A1(abar[11]), .A2(bbar[10]), .ZN(ybar[186]) );
  AND2_X1 U162 ( .A1(a[11]), .A2(b[9]), .ZN(y[185]) );
  OR2_X1 U162bar ( .A1(abar[11]), .A2(bbar[9]), .ZN(ybar[185]) );
  AND2_X1 U163 ( .A1(a[11]), .A2(b[8]), .ZN(y[184]) );
  OR2_X1 U163bar ( .A1(abar[11]), .A2(bbar[8]), .ZN(ybar[184]) );
  AND2_X1 U164 ( .A1(a[11]), .A2(b[7]), .ZN(y[183]) );
  OR2_X1 U164bar ( .A1(abar[11]), .A2(bbar[7]), .ZN(ybar[183]) );
  AND2_X1 U165 ( .A1(a[11]), .A2(b[6]), .ZN(y[182]) );
  OR2_X1 U165bar ( .A1(abar[11]), .A2(bbar[6]), .ZN(ybar[182]) );
  AND2_X1 U166 ( .A1(a[11]), .A2(b[5]), .ZN(y[181]) );
  OR2_X1 U166bar ( .A1(abar[11]), .A2(bbar[5]), .ZN(ybar[181]) );
  AND2_X1 U167 ( .A1(a[11]), .A2(b[4]), .ZN(y[180]) );
  OR2_X1 U167bar ( .A1(abar[11]), .A2(bbar[4]), .ZN(ybar[180]) );
  AND2_X1 U168 ( .A1(a[1]), .A2(b[1]), .ZN(y[17]) );
  OR2_X1 U168bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[17]) );
  AND2_X1 U169 ( .A1(a[11]), .A2(b[3]), .ZN(y[179]) );
  OR2_X1 U169bar ( .A1(abar[11]), .A2(bbar[3]), .ZN(ybar[179]) );
  AND2_X1 U170 ( .A1(a[11]), .A2(b[2]), .ZN(y[178]) );
  OR2_X1 U170bar ( .A1(abar[11]), .A2(bbar[2]), .ZN(ybar[178]) );
  AND2_X1 U171 ( .A1(a[11]), .A2(b[1]), .ZN(y[177]) );
  OR2_X1 U171bar ( .A1(abar[11]), .A2(bbar[1]), .ZN(ybar[177]) );
  AND2_X1 U172 ( .A1(a[11]), .A2(b[0]), .ZN(y[176]) );
  OR2_X1 U172bar ( .A1(abar[11]), .A2(bbar[0]), .ZN(ybar[176]) );
  AND2_X1 U173 ( .A1(a[10]), .A2(b[15]), .ZN(y[175]) );
  OR2_X1 U173bar ( .A1(abar[10]), .A2(bbar[15]), .ZN(ybar[175]) );
  AND2_X1 U174 ( .A1(a[10]), .A2(b[14]), .ZN(y[174]) );
  OR2_X1 U174bar ( .A1(abar[10]), .A2(bbar[14]), .ZN(ybar[174]) );
  AND2_X1 U175 ( .A1(a[10]), .A2(b[13]), .ZN(y[173]) );
  OR2_X1 U175bar ( .A1(abar[10]), .A2(bbar[13]), .ZN(ybar[173]) );
  AND2_X1 U176 ( .A1(a[10]), .A2(b[12]), .ZN(y[172]) );
  OR2_X1 U176bar ( .A1(abar[10]), .A2(bbar[12]), .ZN(ybar[172]) );
  AND2_X1 U177 ( .A1(a[10]), .A2(b[11]), .ZN(y[171]) );
  OR2_X1 U177bar ( .A1(abar[10]), .A2(bbar[11]), .ZN(ybar[171]) );
  AND2_X1 U178 ( .A1(a[10]), .A2(b[10]), .ZN(y[170]) );
  OR2_X1 U178bar ( .A1(abar[10]), .A2(bbar[10]), .ZN(ybar[170]) );
  AND2_X1 U179 ( .A1(a[1]), .A2(b[0]), .ZN(y[16]) );
  OR2_X1 U179bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[16]) );
  AND2_X1 U180 ( .A1(a[10]), .A2(b[9]), .ZN(y[169]) );
  OR2_X1 U180bar ( .A1(abar[10]), .A2(bbar[9]), .ZN(ybar[169]) );
  AND2_X1 U181 ( .A1(a[10]), .A2(b[8]), .ZN(y[168]) );
  OR2_X1 U181bar ( .A1(abar[10]), .A2(bbar[8]), .ZN(ybar[168]) );
  AND2_X1 U182 ( .A1(a[10]), .A2(b[7]), .ZN(y[167]) );
  OR2_X1 U182bar ( .A1(abar[10]), .A2(bbar[7]), .ZN(ybar[167]) );
  AND2_X1 U183 ( .A1(a[10]), .A2(b[6]), .ZN(y[166]) );
  OR2_X1 U183bar ( .A1(abar[10]), .A2(bbar[6]), .ZN(ybar[166]) );
  AND2_X1 U184 ( .A1(a[10]), .A2(b[5]), .ZN(y[165]) );
  OR2_X1 U184bar ( .A1(abar[10]), .A2(bbar[5]), .ZN(ybar[165]) );
  AND2_X1 U185 ( .A1(a[10]), .A2(b[4]), .ZN(y[164]) );
  OR2_X1 U185bar ( .A1(abar[10]), .A2(bbar[4]), .ZN(ybar[164]) );
  AND2_X1 U186 ( .A1(a[10]), .A2(b[3]), .ZN(y[163]) );
  OR2_X1 U186bar ( .A1(abar[10]), .A2(bbar[3]), .ZN(ybar[163]) );
  AND2_X1 U187 ( .A1(a[10]), .A2(b[2]), .ZN(y[162]) );
  OR2_X1 U187bar ( .A1(abar[10]), .A2(bbar[2]), .ZN(ybar[162]) );
  AND2_X1 U188 ( .A1(a[10]), .A2(b[1]), .ZN(y[161]) );
  OR2_X1 U188bar ( .A1(abar[10]), .A2(bbar[1]), .ZN(ybar[161]) );
  AND2_X1 U189 ( .A1(a[10]), .A2(b[0]), .ZN(y[160]) );
  OR2_X1 U189bar ( .A1(abar[10]), .A2(bbar[0]), .ZN(ybar[160]) );
  AND2_X1 U190 ( .A1(b[15]), .A2(a[0]), .ZN(y[15]) );
  OR2_X1 U190bar ( .A1(bbar[15]), .A2(abar[0]), .ZN(ybar[15]) );
  AND2_X1 U191 ( .A1(a[9]), .A2(b[15]), .ZN(y[159]) );
  OR2_X1 U191bar ( .A1(abar[9]), .A2(bbar[15]), .ZN(ybar[159]) );
  AND2_X1 U192 ( .A1(a[9]), .A2(b[14]), .ZN(y[158]) );
  OR2_X1 U192bar ( .A1(abar[9]), .A2(bbar[14]), .ZN(ybar[158]) );
  AND2_X1 U193 ( .A1(a[9]), .A2(b[13]), .ZN(y[157]) );
  OR2_X1 U193bar ( .A1(abar[9]), .A2(bbar[13]), .ZN(ybar[157]) );
  AND2_X1 U194 ( .A1(a[9]), .A2(b[12]), .ZN(y[156]) );
  OR2_X1 U194bar ( .A1(abar[9]), .A2(bbar[12]), .ZN(ybar[156]) );
  AND2_X1 U195 ( .A1(a[9]), .A2(b[11]), .ZN(y[155]) );
  OR2_X1 U195bar ( .A1(abar[9]), .A2(bbar[11]), .ZN(ybar[155]) );
  AND2_X1 U196 ( .A1(a[9]), .A2(b[10]), .ZN(y[154]) );
  OR2_X1 U196bar ( .A1(abar[9]), .A2(bbar[10]), .ZN(ybar[154]) );
  AND2_X1 U197 ( .A1(a[9]), .A2(b[9]), .ZN(y[153]) );
  OR2_X1 U197bar ( .A1(abar[9]), .A2(bbar[9]), .ZN(ybar[153]) );
  AND2_X1 U198 ( .A1(a[9]), .A2(b[8]), .ZN(y[152]) );
  OR2_X1 U198bar ( .A1(abar[9]), .A2(bbar[8]), .ZN(ybar[152]) );
  AND2_X1 U199 ( .A1(a[9]), .A2(b[7]), .ZN(y[151]) );
  OR2_X1 U199bar ( .A1(abar[9]), .A2(bbar[7]), .ZN(ybar[151]) );
  AND2_X1 U200 ( .A1(a[9]), .A2(b[6]), .ZN(y[150]) );
  OR2_X1 U200bar ( .A1(abar[9]), .A2(bbar[6]), .ZN(ybar[150]) );
  AND2_X1 U201 ( .A1(b[14]), .A2(a[0]), .ZN(y[14]) );
  OR2_X1 U201bar ( .A1(bbar[14]), .A2(abar[0]), .ZN(ybar[14]) );
  AND2_X1 U202 ( .A1(a[9]), .A2(b[5]), .ZN(y[149]) );
  OR2_X1 U202bar ( .A1(abar[9]), .A2(bbar[5]), .ZN(ybar[149]) );
  AND2_X1 U203 ( .A1(a[9]), .A2(b[4]), .ZN(y[148]) );
  OR2_X1 U203bar ( .A1(abar[9]), .A2(bbar[4]), .ZN(ybar[148]) );
  AND2_X1 U204 ( .A1(a[9]), .A2(b[3]), .ZN(y[147]) );
  OR2_X1 U204bar ( .A1(abar[9]), .A2(bbar[3]), .ZN(ybar[147]) );
  AND2_X1 U205 ( .A1(a[9]), .A2(b[2]), .ZN(y[146]) );
  OR2_X1 U205bar ( .A1(abar[9]), .A2(bbar[2]), .ZN(ybar[146]) );
  AND2_X1 U206 ( .A1(a[9]), .A2(b[1]), .ZN(y[145]) );
  OR2_X1 U206bar ( .A1(abar[9]), .A2(bbar[1]), .ZN(ybar[145]) );
  AND2_X1 U207 ( .A1(a[9]), .A2(b[0]), .ZN(y[144]) );
  OR2_X1 U207bar ( .A1(abar[9]), .A2(bbar[0]), .ZN(ybar[144]) );
  AND2_X1 U208 ( .A1(a[8]), .A2(b[15]), .ZN(y[143]) );
  OR2_X1 U208bar ( .A1(abar[8]), .A2(bbar[15]), .ZN(ybar[143]) );
  AND2_X1 U209 ( .A1(a[8]), .A2(b[14]), .ZN(y[142]) );
  OR2_X1 U209bar ( .A1(abar[8]), .A2(bbar[14]), .ZN(ybar[142]) );
  AND2_X1 U210 ( .A1(a[8]), .A2(b[13]), .ZN(y[141]) );
  OR2_X1 U210bar ( .A1(abar[8]), .A2(bbar[13]), .ZN(ybar[141]) );
  AND2_X1 U211 ( .A1(a[8]), .A2(b[12]), .ZN(y[140]) );
  OR2_X1 U211bar ( .A1(abar[8]), .A2(bbar[12]), .ZN(ybar[140]) );
  AND2_X1 U212 ( .A1(b[13]), .A2(a[0]), .ZN(y[13]) );
  OR2_X1 U212bar ( .A1(bbar[13]), .A2(abar[0]), .ZN(ybar[13]) );
  AND2_X1 U213 ( .A1(a[8]), .A2(b[11]), .ZN(y[139]) );
  OR2_X1 U213bar ( .A1(abar[8]), .A2(bbar[11]), .ZN(ybar[139]) );
  AND2_X1 U214 ( .A1(a[8]), .A2(b[10]), .ZN(y[138]) );
  OR2_X1 U214bar ( .A1(abar[8]), .A2(bbar[10]), .ZN(ybar[138]) );
  AND2_X1 U215 ( .A1(a[8]), .A2(b[9]), .ZN(y[137]) );
  OR2_X1 U215bar ( .A1(abar[8]), .A2(bbar[9]), .ZN(ybar[137]) );
  AND2_X1 U216 ( .A1(a[8]), .A2(b[8]), .ZN(y[136]) );
  OR2_X1 U216bar ( .A1(abar[8]), .A2(bbar[8]), .ZN(ybar[136]) );
  AND2_X1 U217 ( .A1(a[8]), .A2(b[7]), .ZN(y[135]) );
  OR2_X1 U217bar ( .A1(abar[8]), .A2(bbar[7]), .ZN(ybar[135]) );
  AND2_X1 U218 ( .A1(a[8]), .A2(b[6]), .ZN(y[134]) );
  OR2_X1 U218bar ( .A1(abar[8]), .A2(bbar[6]), .ZN(ybar[134]) );
  AND2_X1 U219 ( .A1(a[8]), .A2(b[5]), .ZN(y[133]) );
  OR2_X1 U219bar ( .A1(abar[8]), .A2(bbar[5]), .ZN(ybar[133]) );
  AND2_X1 U220 ( .A1(a[8]), .A2(b[4]), .ZN(y[132]) );
  OR2_X1 U220bar ( .A1(abar[8]), .A2(bbar[4]), .ZN(ybar[132]) );
  AND2_X1 U221 ( .A1(a[8]), .A2(b[3]), .ZN(y[131]) );
  OR2_X1 U221bar ( .A1(abar[8]), .A2(bbar[3]), .ZN(ybar[131]) );
  AND2_X1 U222 ( .A1(a[8]), .A2(b[2]), .ZN(y[130]) );
  OR2_X1 U222bar ( .A1(abar[8]), .A2(bbar[2]), .ZN(ybar[130]) );
  AND2_X1 U223 ( .A1(b[12]), .A2(a[0]), .ZN(y[12]) );
  OR2_X1 U223bar ( .A1(bbar[12]), .A2(abar[0]), .ZN(ybar[12]) );
  AND2_X1 U224 ( .A1(a[8]), .A2(b[1]), .ZN(y[129]) );
  OR2_X1 U224bar ( .A1(abar[8]), .A2(bbar[1]), .ZN(ybar[129]) );
  AND2_X1 U225 ( .A1(a[8]), .A2(b[0]), .ZN(y[128]) );
  OR2_X1 U225bar ( .A1(abar[8]), .A2(bbar[0]), .ZN(ybar[128]) );
  AND2_X1 U226 ( .A1(a[7]), .A2(b[15]), .ZN(y[127]) );
  OR2_X1 U226bar ( .A1(abar[7]), .A2(bbar[15]), .ZN(ybar[127]) );
  AND2_X1 U227 ( .A1(a[7]), .A2(b[14]), .ZN(y[126]) );
  OR2_X1 U227bar ( .A1(abar[7]), .A2(bbar[14]), .ZN(ybar[126]) );
  AND2_X1 U228 ( .A1(a[7]), .A2(b[13]), .ZN(y[125]) );
  OR2_X1 U228bar ( .A1(abar[7]), .A2(bbar[13]), .ZN(ybar[125]) );
  AND2_X1 U229 ( .A1(a[7]), .A2(b[12]), .ZN(y[124]) );
  OR2_X1 U229bar ( .A1(abar[7]), .A2(bbar[12]), .ZN(ybar[124]) );
  AND2_X1 U230 ( .A1(a[7]), .A2(b[11]), .ZN(y[123]) );
  OR2_X1 U230bar ( .A1(abar[7]), .A2(bbar[11]), .ZN(ybar[123]) );
  AND2_X1 U231 ( .A1(a[7]), .A2(b[10]), .ZN(y[122]) );
  OR2_X1 U231bar ( .A1(abar[7]), .A2(bbar[10]), .ZN(ybar[122]) );
  AND2_X1 U232 ( .A1(a[7]), .A2(b[9]), .ZN(y[121]) );
  OR2_X1 U232bar ( .A1(abar[7]), .A2(bbar[9]), .ZN(ybar[121]) );
  AND2_X1 U233 ( .A1(a[7]), .A2(b[8]), .ZN(y[120]) );
  OR2_X1 U233bar ( .A1(abar[7]), .A2(bbar[8]), .ZN(ybar[120]) );
  AND2_X1 U234 ( .A1(b[11]), .A2(a[0]), .ZN(y[11]) );
  OR2_X1 U234bar ( .A1(bbar[11]), .A2(abar[0]), .ZN(ybar[11]) );
  AND2_X1 U235 ( .A1(a[7]), .A2(b[7]), .ZN(y[119]) );
  OR2_X1 U235bar ( .A1(abar[7]), .A2(bbar[7]), .ZN(ybar[119]) );
  AND2_X1 U236 ( .A1(a[7]), .A2(b[6]), .ZN(y[118]) );
  OR2_X1 U236bar ( .A1(abar[7]), .A2(bbar[6]), .ZN(ybar[118]) );
  AND2_X1 U237 ( .A1(a[7]), .A2(b[5]), .ZN(y[117]) );
  OR2_X1 U237bar ( .A1(abar[7]), .A2(bbar[5]), .ZN(ybar[117]) );
  AND2_X1 U238 ( .A1(a[7]), .A2(b[4]), .ZN(y[116]) );
  OR2_X1 U238bar ( .A1(abar[7]), .A2(bbar[4]), .ZN(ybar[116]) );
  AND2_X1 U239 ( .A1(a[7]), .A2(b[3]), .ZN(y[115]) );
  OR2_X1 U239bar ( .A1(abar[7]), .A2(bbar[3]), .ZN(ybar[115]) );
  AND2_X1 U240 ( .A1(a[7]), .A2(b[2]), .ZN(y[114]) );
  OR2_X1 U240bar ( .A1(abar[7]), .A2(bbar[2]), .ZN(ybar[114]) );
  AND2_X1 U241 ( .A1(a[7]), .A2(b[1]), .ZN(y[113]) );
  OR2_X1 U241bar ( .A1(abar[7]), .A2(bbar[1]), .ZN(ybar[113]) );
  AND2_X1 U242 ( .A1(a[7]), .A2(b[0]), .ZN(y[112]) );
  OR2_X1 U242bar ( .A1(abar[7]), .A2(bbar[0]), .ZN(ybar[112]) );
  AND2_X1 U243 ( .A1(b[15]), .A2(a[6]), .ZN(y[111]) );
  OR2_X1 U243bar ( .A1(bbar[15]), .A2(abar[6]), .ZN(ybar[111]) );
  AND2_X1 U244 ( .A1(b[14]), .A2(a[6]), .ZN(y[110]) );
  OR2_X1 U244bar ( .A1(bbar[14]), .A2(abar[6]), .ZN(ybar[110]) );
  AND2_X1 U245 ( .A1(b[10]), .A2(a[0]), .ZN(y[10]) );
  OR2_X1 U245bar ( .A1(bbar[10]), .A2(abar[0]), .ZN(ybar[10]) );
  AND2_X1 U246 ( .A1(b[13]), .A2(a[6]), .ZN(y[109]) );
  OR2_X1 U246bar ( .A1(bbar[13]), .A2(abar[6]), .ZN(ybar[109]) );
  AND2_X1 U247 ( .A1(b[12]), .A2(a[6]), .ZN(y[108]) );
  OR2_X1 U247bar ( .A1(bbar[12]), .A2(abar[6]), .ZN(ybar[108]) );
  AND2_X1 U248 ( .A1(b[11]), .A2(a[6]), .ZN(y[107]) );
  OR2_X1 U248bar ( .A1(bbar[11]), .A2(abar[6]), .ZN(ybar[107]) );
  AND2_X1 U249 ( .A1(b[10]), .A2(a[6]), .ZN(y[106]) );
  OR2_X1 U249bar ( .A1(bbar[10]), .A2(abar[6]), .ZN(ybar[106]) );
  AND2_X1 U250 ( .A1(a[6]), .A2(b[9]), .ZN(y[105]) );
  OR2_X1 U250bar ( .A1(abar[6]), .A2(bbar[9]), .ZN(ybar[105]) );
  AND2_X1 U251 ( .A1(b[8]), .A2(a[6]), .ZN(y[104]) );
  OR2_X1 U251bar ( .A1(bbar[8]), .A2(abar[6]), .ZN(ybar[104]) );
  AND2_X1 U252 ( .A1(b[7]), .A2(a[6]), .ZN(y[103]) );
  OR2_X1 U252bar ( .A1(bbar[7]), .A2(abar[6]), .ZN(ybar[103]) );
  AND2_X1 U253 ( .A1(b[6]), .A2(a[6]), .ZN(y[102]) );
  OR2_X1 U253bar ( .A1(bbar[6]), .A2(abar[6]), .ZN(ybar[102]) );
  AND2_X1 U254 ( .A1(b[5]), .A2(a[6]), .ZN(y[101]) );
  OR2_X1 U254bar ( .A1(bbar[5]), .A2(abar[6]), .ZN(ybar[101]) );
  AND2_X1 U255 ( .A1(b[4]), .A2(a[6]), .ZN(y[100]) );
  OR2_X1 U255bar ( .A1(bbar[4]), .A2(abar[6]), .ZN(ybar[100]) );
  AND2_X1 U256 ( .A1(b[0]), .A2(a[0]), .ZN(y[0]) );
  OR2_X1 U256bar ( .A1(bbar[0]), .A2(abar[0]), .ZN(ybar[0]) );
endmodule

module decode_9 ( in, inbar, out, outbar );

  input wire [7:0] in;
  input wire [7:0] inbar;
//input_done

  output wire [255:0] out;
  output wire [255:0] outbar;
//output_done

  wire [15:0] level1;
  wire [31:0] level2;
  wire [15:0] level1bar;
  wire [31:0] level2bar;
//wire_done

  CD2_36 cd_l1_1 ( .a(in[1]), .abar(inbar[1]), .b(in[0]), .bbar(inbar[0]), .y(level1[3:0]), .ybar(level1bar[3:0]) );
  CD2_35 cd_l1_2 ( .a(in[3]), .abar(inbar[3]), .b(in[2]), .bbar(inbar[2]), .y(level1[7:4]), .ybar(level1bar[7:4]) );
  CD2_34 cd_l1_3 ( .a(in[5]), .abar(inbar[5]), .b(in[4]), .bbar(inbar[4]), .y(level1[11:8]), .ybar(level1bar[11:8]) );
  CD2_33 cd_l1_4 ( .a(in[7]), .abar(inbar[7]), .b(in[6]), .bbar(inbar[6]), .y(level1[15:12]), .ybar(level1bar[15:12]) );

  CD4_18 cd_l2_1 ( .a(level1[7:4]), .abar(level1bar[7:4]), .b(level1[3:0]), .bbar(level1bar[3:0]), 
        .y(level2[15:0]), .ybar(level2bar[15:0]) );
  CD4_17 cd_l2_2 ( .a(level1[15:12]), .abar(level1bar[15:12]), .b(level1[11:8]), .bbar(level1bar[11:8]), 
        .y(level2[31:16]), .ybar(level2bar[31:16]) );
  CD16_9 cd_l3 ( .a(level2[31:16]), .abar(level2bar[31:16]), .b(level2[15:0]), .bbar(level2bar[15:0]), 
        .y(out), .ybar(outbar) );
endmodule

module encode_9 ( in, inbar, out, outbar );

  input wire [255:0] in;
  input wire [255:0] inbar;
//input_done

  output wire [7:0] out;
  output wire [7:0] outbar;
//output_done

  wire in_81;
  wire in_80;
  wire in_79;
  wire in_78;
  wire in_77;
  wire in_76;
  wire in_75;
  wire in_74;
  wire in_73;
  wire in_72;
  wire in_71;
  wire in_70;
  wire in_69;
  wire in_68;
  wire in_67;
  wire in_66;
  wire in_65;
  wire in_64;
  wire in_63;
  wire in_62;
  wire in_61;
  wire in_60;
  wire in_59;
  wire in_58;
  wire in_57;
  wire in_56;
  wire in_55;
  wire in_54;
  wire in_53;
  wire in_52;
  wire in_51;
  wire in_50;
  wire in_49;
  wire in_48;
  wire in_47;
  wire in_46;
  wire in_45;
  wire in_44;
  wire in_43;
  wire in_42;
  wire in_41;
  wire in_40;
  wire in_39;
  wire in_38;
  wire in_37;
  wire in_36;
  wire in_35;
  wire in_34;
  wire in_33;
  wire in_32;
  wire in_31;
  wire in_30;
  wire in_29;
  wire in_28;
  wire in_27;
  wire in_26;
  wire in_25;
  wire in_24;
  wire in_23;
  wire in_22;
  wire in_21;
  wire in_20;
  wire in_19;
  wire in_18;
  wire in_17;
  wire in_16;
  wire in_15;
  wire in_14;
  wire in_13;
  wire in_12;
  wire in_11;
  wire in_10;
  wire in_9;
  wire in_8;
  wire in_7;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_3;
  wire in_2;
  wire in_1;
  wire in_0;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire in_81bar;
  wire in_80bar;
  wire in_79bar;
  wire in_78bar;
  wire in_77bar;
  wire in_76bar;
  wire in_75bar;
  wire in_74bar;
  wire in_73bar;
  wire in_72bar;
  wire in_71bar;
  wire in_70bar;
  wire in_69bar;
  wire in_68bar;
  wire in_67bar;
  wire in_66bar;
  wire in_65bar;
  wire in_64bar;
  wire in_63bar;
  wire in_62bar;
  wire in_61bar;
  wire in_60bar;
  wire in_59bar;
  wire in_58bar;
  wire in_57bar;
  wire in_56bar;
  wire in_55bar;
  wire in_54bar;
  wire in_53bar;
  wire in_52bar;
  wire in_51bar;
  wire in_50bar;
  wire in_49bar;
  wire in_48bar;
  wire in_47bar;
  wire in_46bar;
  wire in_45bar;
  wire in_44bar;
  wire in_43bar;
  wire in_42bar;
  wire in_41bar;
  wire in_40bar;
  wire in_39bar;
  wire in_38bar;
  wire in_37bar;
  wire in_36bar;
  wire in_35bar;
  wire in_34bar;
  wire in_33bar;
  wire in_32bar;
  wire in_31bar;
  wire in_30bar;
  wire in_29bar;
  wire in_28bar;
  wire in_27bar;
  wire in_26bar;
  wire in_25bar;
  wire in_24bar;
  wire in_23bar;
  wire in_22bar;
  wire in_21bar;
  wire in_20bar;
  wire in_19bar;
  wire in_18bar;
  wire in_17bar;
  wire in_16bar;
  wire in_15bar;
  wire in_14bar;
  wire in_13bar;
  wire in_12bar;
  wire in_11bar;
  wire in_10bar;
  wire in_9bar;
  wire in_8bar;
  wire in_7bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_3bar;
  wire in_2bar;
  wire in_1bar;
  wire in_0bar;
  wire n487bar;
  wire n488bar;
  wire n489bar;
  wire n490bar;
  wire n491bar;
  wire n492bar;
  wire n493bar;
  wire n494bar;
  wire n495bar;
  wire n496bar;
  wire n497bar;
  wire n498bar;
  wire n499bar;
  wire n500bar;
  wire n501bar;
  wire n502bar;
  wire n503bar;
  wire n504bar;
  wire n505bar;
  wire n506bar;
  wire n507bar;
  wire n508bar;
  wire n509bar;
  wire n510bar;
  wire n511bar;
  wire n512bar;
  wire n513bar;
  wire n514bar;
  wire n515bar;
  wire n516bar;
  wire n517bar;
  wire n518bar;
  wire n519bar;
  wire n520bar;
  wire n521bar;
  wire n522bar;
  wire n523bar;
  wire n524bar;
  wire n525bar;
  wire n526bar;
  wire n527bar;
  wire n528bar;
  wire n529bar;
  wire n530bar;
  wire n531bar;
  wire n532bar;
  wire n533bar;
  wire n534bar;
  wire n535bar;
  wire n536bar;
  wire n537bar;
  wire n538bar;
  wire n539bar;
  wire n540bar;
  wire n541bar;
  wire n542bar;
  wire n543bar;
  wire n544bar;
  wire n545bar;
  wire n546bar;
  wire n547bar;
  wire n548bar;
  wire n549bar;
  wire n550bar;
  wire n551bar;
  wire n552bar;
  wire n553bar;
  wire n554bar;
  wire n555bar;
  wire n556bar;
  wire n557bar;
  wire n558bar;
  wire n559bar;
  wire n560bar;
  wire n561bar;
  wire n562bar;
  wire n563bar;
  wire n564bar;
  wire n565bar;
  wire n566bar;
  wire n567bar;
  wire n568bar;
  wire n569bar;
  wire n570bar;
  wire n571bar;
  wire n572bar;
  wire n573bar;
  wire n574bar;
  wire n575bar;
  wire n576bar;
  wire n577bar;
  wire n578bar;
  wire n579bar;
  wire n580bar;
  wire n581bar;
  wire n582bar;
  wire n583bar;
  wire n584bar;
  wire n585bar;
  wire n586bar;
  wire n587bar;
  wire n588bar;
  wire n589bar;
  wire n590bar;
  wire n591bar;
  wire n592bar;
  wire n593bar;
  wire n594bar;
  wire n595bar;
  wire n596bar;
  wire n597bar;
  wire n598bar;
  wire n599bar;
  wire n600bar;
  wire n601bar;
  wire n602bar;
  wire n603bar;
  wire n604bar;
  wire n605bar;
  wire n606bar;
  wire n607bar;
  wire n608bar;
  wire n609bar;
  wire n610bar;
  wire n611bar;
  wire n612bar;
  wire n613bar;
  wire n614bar;
  wire n615bar;
  wire n616bar;
  wire n617bar;
  wire n618bar;
  wire n619bar;
  wire n620bar;
  wire n621bar;
  wire n622bar;
  wire n623bar;
  wire n624bar;
  wire n625bar;
  wire n626bar;
  wire n627bar;
  wire n628bar;
  wire n629bar;
  wire n630bar;
  wire n631bar;
  wire n632bar;
  wire n633bar;
  wire n634bar;
  wire n635bar;
  wire n636bar;
  wire n637bar;
  wire n638bar;
  wire n639bar;
  wire n640bar;
  wire n641bar;
  wire n642bar;
  wire n643bar;
  wire n644bar;
  wire n645bar;
  wire n646bar;
  wire n647bar;
  wire n648bar;
  wire n649bar;
  wire n650bar;
  wire n651bar;
  wire n652bar;
  wire n653bar;
  wire n654bar;
  wire n655bar;
  wire n656bar;
  wire n657bar;
  wire n658bar;
  wire n659bar;
  wire n660bar;
  wire n661bar;
  wire n662bar;
  wire n663bar;
  wire n664bar;
  wire n665bar;
  wire n666bar;
  wire n667bar;
  wire n668bar;
  wire n669bar;
  wire n670bar;
  wire n671bar;
  wire n672bar;
  wire n673bar;
  wire n674bar;
  wire n675bar;
  wire n676bar;
  wire n677bar;
  wire n678bar;
  wire n679bar;
  wire n680bar;
  wire n681bar;
  wire n682bar;
  wire n683bar;
  wire n684bar;
  wire n685bar;
  wire n686bar;
  wire n687bar;
  wire n688bar;
  wire n689bar;
  wire n690bar;
  wire n691bar;
  wire n692bar;
  wire n693bar;
  wire n694bar;
  wire n695bar;
  wire n696bar;
  wire n697bar;
  wire n698bar;
  wire n699bar;
  wire n700bar;
  wire n701bar;
  wire n702bar;
  wire n703bar;
  wire n704bar;
  wire n705bar;
  wire n706bar;
  wire n707bar;
  wire n708bar;
  wire n709bar;
  wire n710bar;
  wire n711bar;
  wire n712bar;
  wire n713bar;
  wire n714bar;
  wire n715bar;
  wire n716bar;
  wire n717bar;
  wire n718bar;
  wire n719bar;
  wire n720bar;
  wire n721bar;
  wire n722bar;
  wire n723bar;
  wire n724bar;
  wire n725bar;
  wire n726bar;
  wire n727bar;
  wire n728bar;
  wire n729bar;
  wire n730bar;
  wire n731bar;
  wire n732bar;
  wire n733bar;
  wire n734bar;
  wire n735bar;
  wire n736bar;
  wire n737bar;
  wire n738bar;
  wire n739bar;
  wire n740bar;
  wire n741bar;
  wire n742bar;
  wire n743bar;
  wire n744bar;
  wire n745bar;
  wire n746bar;
  wire n747bar;
  wire n748bar;
  wire n749bar;
  wire n750bar;
  wire n751bar;
  wire n752bar;
  wire n753bar;
  wire n754bar;
  wire n755bar;
  wire n756bar;
  wire n757bar;
  wire n758bar;
  wire n759bar;
  wire n760bar;
  wire n761bar;
  wire n762bar;
  wire n763bar;
  wire n764bar;
  wire n765bar;
  wire n766bar;
  wire n767bar;
  wire n768bar;
  wire n769bar;
  wire n770bar;
  wire n771bar;
  wire n772bar;
  wire n773bar;
  wire n774bar;
  wire n775bar;
  wire n776bar;
  wire n777bar;
  wire n778bar;
  wire n779bar;
  wire n780bar;
  wire n781bar;
  wire n782bar;
  wire n783bar;
  wire n784bar;
  wire n785bar;
  wire n786bar;
  wire n787bar;
  wire n788bar;
  wire n789bar;
  wire n790bar;
  wire n791bar;
  wire n792bar;
  wire n793bar;
  wire n794bar;
  wire n795bar;
  wire n796bar;
  wire n797bar;
  wire n798bar;
  wire n799bar;
  wire n800bar;
  wire n801bar;
  wire n802bar;
  wire n803bar;
  wire n804bar;
  wire n805bar;
  wire n806bar;
  wire n807bar;
  wire n808bar;
  wire n809bar;
  wire n810bar;
  wire n811bar;
  wire n812bar;
  wire n813bar;
  wire n814bar;
  wire n815bar;
  wire n816bar;
  wire n817bar;
  wire n818bar;
  wire n819bar;
  wire n820bar;
  wire n821bar;
  wire n822bar;
  wire n823bar;
  wire n824bar;
  wire n825bar;
  wire n826bar;
  wire n827bar;
  wire n828bar;
  wire n829bar;
  wire n830bar;
  wire n831bar;
  wire n832bar;
  wire n833bar;
  wire n834bar;
  wire n835bar;
  wire n836bar;
  wire n837bar;
  wire n838bar;
  wire n839bar;
  wire n840bar;
  wire n841bar;
  wire n842bar;
  wire n843bar;
  wire n844bar;
  wire n845bar;
  wire n846bar;
  wire n847bar;
  wire n848bar;
  wire n849bar;
  wire n850bar;
  wire n851bar;
  wire n852bar;
  wire n853bar;
  wire n854bar;
  wire n855bar;
  wire n856bar;
  wire n857bar;
  wire n858bar;
  wire n859bar;
  wire n860bar;
  wire n861bar;
  wire n862bar;
  wire n863bar;
  wire n864bar;
  wire n865bar;
  wire n866bar;
  wire n867bar;
  wire n868bar;
  wire n869bar;
  wire n870bar;
  wire n871bar;
  wire n872bar;
  wire n873bar;
  wire n874bar;
  wire n875bar;
  wire n876bar;
  wire n877bar;
  wire n878bar;
  wire n879bar;
  wire n880bar;
  wire n881bar;
  wire n882bar;
  wire n883bar;
  wire n884bar;
  wire n885bar;
  wire n886bar;
  wire n887bar;
  wire n888bar;
  wire n889bar;
  wire n890bar;
  wire n891bar;
  wire n892bar;
  wire n893bar;
  wire n894bar;
  wire n895bar;
  wire n896bar;
  wire n897bar;
  wire n898bar;
  wire n899bar;
  wire n900bar;
  wire n901bar;
  wire n902bar;
  wire n903bar;
  wire n904bar;
  wire n905bar;
  wire n906bar;
  wire n907bar;
  wire n908bar;
  wire n909bar;
  wire n910bar;
  wire n911bar;
  wire n912bar;
  wire n913bar;
  wire n914bar;
  wire n915bar;
  wire n916bar;
  wire n917bar;
  wire n918bar;
  wire n919bar;
  wire n920bar;
  wire n921bar;
  wire n922bar;
  wire n923bar;
  wire n924bar;
  wire n925bar;
  wire n926bar;
  wire n927bar;
  wire n928bar;
  wire n929bar;
  wire n930bar;
  wire n931bar;
  wire n932bar;
  wire n933bar;
  wire n934bar;
  wire n935bar;
  wire n936bar;
  wire n937bar;
  wire n938bar;
  wire n939bar;
  wire n940bar;
  wire n941bar;
  wire n942bar;
  wire n943bar;
  wire n944bar;
  wire n945bar;
  wire n946bar;
  wire n947bar;
  wire n948bar;
  wire n949bar;
  wire n950bar;
  wire n951bar;
  wire n952bar;
  wire n953bar;
  wire n954bar;
  wire n955bar;
  wire n956bar;
  wire n957bar;
  wire n958bar;
  wire n959bar;
  wire n960bar;
  wire n961bar;
  wire n962bar;
  wire n963bar;
  wire n964bar;
  wire n965bar;
  wire n966bar;
  wire n967bar;
  wire n968bar;
  wire n969bar;
  wire n970bar;
  wire n971bar;
  wire n972bar;
//wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];
  assign in_81bar = inbar[81];
  assign in_80bar = inbar[80];
  assign in_79bar = inbar[79];
  assign in_78bar = inbar[78];
  assign in_77bar = inbar[77];
  assign in_76bar = inbar[76];
  assign in_75bar = inbar[75];
  assign in_74bar = inbar[74];
  assign in_73bar = inbar[73];
  assign in_72bar = inbar[72];
  assign in_71bar = inbar[71];
  assign in_70bar = inbar[70];
  assign in_69bar = inbar[69];
  assign in_68bar = inbar[68];
  assign in_67bar = inbar[67];
  assign in_66bar = inbar[66];
  assign in_65bar = inbar[65];
  assign in_64bar = inbar[64];
  assign in_63bar = inbar[63];
  assign in_62bar = inbar[62];
  assign in_61bar = inbar[61];
  assign in_60bar = inbar[60];
  assign in_59bar = inbar[59];
  assign in_58bar = inbar[58];
  assign in_57bar = inbar[57];
  assign in_56bar = inbar[56];
  assign in_55bar = inbar[55];
  assign in_54bar = inbar[54];
  assign in_53bar = inbar[53];
  assign in_52bar = inbar[52];
  assign in_51bar = inbar[51];
  assign in_50bar = inbar[50];
  assign in_49bar = inbar[49];
  assign in_48bar = inbar[48];
  assign in_47bar = inbar[47];
  assign in_46bar = inbar[46];
  assign in_45bar = inbar[45];
  assign in_44bar = inbar[44];
  assign in_43bar = inbar[43];
  assign in_42bar = inbar[42];
  assign in_41bar = inbar[41];
  assign in_40bar = inbar[40];
  assign in_39bar = inbar[39];
  assign in_38bar = inbar[38];
  assign in_37bar = inbar[37];
  assign in_36bar = inbar[36];
  assign in_35bar = inbar[35];
  assign in_34bar = inbar[34];
  assign in_33bar = inbar[33];
  assign in_32bar = inbar[32];
  assign in_31bar = inbar[31];
  assign in_30bar = inbar[30];
  assign in_29bar = inbar[29];
  assign in_28bar = inbar[28];
  assign in_27bar = inbar[27];
  assign in_26bar = inbar[26];
  assign in_25bar = inbar[25];
  assign in_24bar = inbar[24];
  assign in_23bar = inbar[23];
  assign in_22bar = inbar[22];
  assign in_21bar = inbar[21];
  assign in_20bar = inbar[20];
  assign in_19bar = inbar[19];
  assign in_18bar = inbar[18];
  assign in_17bar = inbar[17];
  assign in_16bar = inbar[16];
  assign in_15bar = inbar[15];
  assign in_14bar = inbar[14];
  assign in_13bar = inbar[13];
  assign in_12bar = inbar[12];
  assign in_11bar = inbar[11];
  assign in_10bar = inbar[10];
  assign in_9bar = inbar[9];
  assign in_8bar = inbar[8];
  assign in_7bar = inbar[7];
  assign in_6bar = inbar[6];
  assign in_5bar = inbar[5];
  assign in_4bar = inbar[4];
  assign in_3bar = inbar[3];
  assign in_2bar = inbar[2];
  assign in_1bar = inbar[1];
  assign in_0bar = inbar[0];
//assign_done

  OR2_X1 U1 ( .A1(n972), .A2(n971), .ZN(out[7]) );
  AND2_X1 U1bar ( .A1(n972bar), .A2(n971bar), .ZN(outbar[7]) );
  OR2_X1 U2 ( .A1(n970), .A2(n969), .ZN(n971) );
  AND2_X1 U2bar ( .A1(n970bar), .A2(n969bar), .ZN(n971bar) );
  OR2_X1 U3 ( .A1(n968), .A2(n967), .ZN(n969) );
  AND2_X1 U3bar ( .A1(n968bar), .A2(n967bar), .ZN(n969bar) );
  OR2_X1 U4 ( .A1(n966), .A2(n965), .ZN(n967) );
  AND2_X1 U4bar ( .A1(n966bar), .A2(n965bar), .ZN(n967bar) );
  OR2_X1 U5 ( .A1(n964), .A2(n963), .ZN(n968) );
  AND2_X1 U5bar ( .A1(n964bar), .A2(n963bar), .ZN(n968bar) );
  OR2_X1 U6 ( .A1(in[116]), .A2(n962), .ZN(n963) );
  AND2_X1 U6bar ( .A1(inbar[116]), .A2(n962bar), .ZN(n963bar) );
  OR2_X1 U7 ( .A1(n961), .A2(n960), .ZN(n970) );
  AND2_X1 U7bar ( .A1(n961bar), .A2(n960bar), .ZN(n970bar) );
  OR2_X1 U8 ( .A1(in[150]), .A2(in[127]), .ZN(n960) );
  AND2_X1 U8bar ( .A1(inbar[150]), .A2(inbar[127]), .ZN(n960bar) );
  OR2_X1 U9 ( .A1(in[160]), .A2(n959), .ZN(n961) );
  AND2_X1 U9bar ( .A1(inbar[160]), .A2(n959bar), .ZN(n961bar) );
  OR2_X1 U10 ( .A1(in[252]), .A2(in[168]), .ZN(n959) );
  AND2_X1 U10bar ( .A1(inbar[252]), .A2(inbar[168]), .ZN(n959bar) );
  OR2_X1 U11 ( .A1(n958), .A2(n957), .ZN(n972) );
  AND2_X1 U11bar ( .A1(n958bar), .A2(n957bar), .ZN(n972bar) );
  OR2_X1 U12 ( .A1(n956), .A2(n955), .ZN(n957) );
  AND2_X1 U12bar ( .A1(n956bar), .A2(n955bar), .ZN(n957bar) );
  OR2_X1 U13 ( .A1(in_17), .A2(in[96]), .ZN(n955) );
  AND2_X1 U13bar ( .A1(in_17bar), .A2(inbar[96]), .ZN(n955bar) );
  OR2_X1 U14 ( .A1(in_23), .A2(n954), .ZN(n956) );
  AND2_X1 U14bar ( .A1(in_23bar), .A2(n954bar), .ZN(n956bar) );
  OR2_X1 U15 ( .A1(in_31), .A2(in_26), .ZN(n954) );
  AND2_X1 U15bar ( .A1(in_31bar), .A2(in_26bar), .ZN(n954bar) );
  OR2_X1 U16 ( .A1(n953), .A2(n952), .ZN(n958) );
  AND2_X1 U16bar ( .A1(n953bar), .A2(n952bar), .ZN(n958bar) );
  OR2_X1 U17 ( .A1(in_58), .A2(in_4), .ZN(n952) );
  AND2_X1 U17bar ( .A1(in_58bar), .A2(in_4bar), .ZN(n952bar) );
  OR2_X1 U18 ( .A1(in_59), .A2(n951), .ZN(n953) );
  AND2_X1 U18bar ( .A1(in_59bar), .A2(n951bar), .ZN(n953bar) );
  OR2_X1 U19 ( .A1(in_71), .A2(in_62), .ZN(n951) );
  AND2_X1 U19bar ( .A1(in_71bar), .A2(in_62bar), .ZN(n951bar) );
  OR2_X1 U20 ( .A1(n950), .A2(n949), .ZN(out[6]) );
  AND2_X1 U20bar ( .A1(n950bar), .A2(n949bar), .ZN(outbar[6]) );
  OR2_X1 U21 ( .A1(n948), .A2(n947), .ZN(n949) );
  AND2_X1 U21bar ( .A1(n948bar), .A2(n947bar), .ZN(n949bar) );
  OR2_X1 U22 ( .A1(n946), .A2(n945), .ZN(n947) );
  AND2_X1 U22bar ( .A1(n946bar), .A2(n945bar), .ZN(n947bar) );
  OR2_X1 U23 ( .A1(n944), .A2(n943), .ZN(n945) );
  AND2_X1 U23bar ( .A1(n944bar), .A2(n943bar), .ZN(n945bar) );
  OR2_X1 U24 ( .A1(n942), .A2(n941), .ZN(n946) );
  AND2_X1 U24bar ( .A1(n942bar), .A2(n941bar), .ZN(n946bar) );
  OR2_X1 U25 ( .A1(in[101]), .A2(n940), .ZN(n941) );
  AND2_X1 U25bar ( .A1(inbar[101]), .A2(n940bar), .ZN(n941bar) );
  OR2_X1 U26 ( .A1(n939), .A2(n938), .ZN(n948) );
  AND2_X1 U26bar ( .A1(n939bar), .A2(n938bar), .ZN(n948bar) );
  OR2_X1 U27 ( .A1(in[114]), .A2(in[104]), .ZN(n938) );
  AND2_X1 U27bar ( .A1(inbar[114]), .A2(inbar[104]), .ZN(n938bar) );
  OR2_X1 U28 ( .A1(in[128]), .A2(n937), .ZN(n939) );
  AND2_X1 U28bar ( .A1(inbar[128]), .A2(n937bar), .ZN(n939bar) );
  OR2_X1 U29 ( .A1(in[136]), .A2(in[134]), .ZN(n937) );
  AND2_X1 U29bar ( .A1(inbar[136]), .A2(inbar[134]), .ZN(n937bar) );
  OR2_X1 U30 ( .A1(n936), .A2(n935), .ZN(n950) );
  AND2_X1 U30bar ( .A1(n936bar), .A2(n935bar), .ZN(n950bar) );
  OR2_X1 U31 ( .A1(n934), .A2(n933), .ZN(n935) );
  AND2_X1 U31bar ( .A1(n934bar), .A2(n933bar), .ZN(n935bar) );
  OR2_X1 U32 ( .A1(in[177]), .A2(in[164]), .ZN(n933) );
  AND2_X1 U32bar ( .A1(inbar[177]), .A2(inbar[164]), .ZN(n933bar) );
  OR2_X1 U33 ( .A1(in[212]), .A2(n932), .ZN(n934) );
  AND2_X1 U33bar ( .A1(inbar[212]), .A2(n932bar), .ZN(n934bar) );
  OR2_X1 U34 ( .A1(in[248]), .A2(in[221]), .ZN(n932) );
  AND2_X1 U34bar ( .A1(inbar[248]), .A2(inbar[221]), .ZN(n932bar) );
  OR2_X1 U35 ( .A1(n931), .A2(n930), .ZN(n936) );
  AND2_X1 U35bar ( .A1(n931bar), .A2(n930bar), .ZN(n936bar) );
  OR2_X1 U36 ( .A1(in_18), .A2(in[93]), .ZN(n930) );
  AND2_X1 U36bar ( .A1(in_18bar), .A2(inbar[93]), .ZN(n930bar) );
  OR2_X1 U37 ( .A1(in_31), .A2(n929), .ZN(n931) );
  AND2_X1 U37bar ( .A1(in_31bar), .A2(n929bar), .ZN(n931bar) );
  OR2_X1 U38 ( .A1(in_7), .A2(in_39), .ZN(n929) );
  AND2_X1 U38bar ( .A1(in_7bar), .A2(in_39bar), .ZN(n929bar) );
  OR2_X1 U39 ( .A1(n928), .A2(n927), .ZN(out[5]) );
  AND2_X1 U39bar ( .A1(n928bar), .A2(n927bar), .ZN(outbar[5]) );
  OR2_X1 U40 ( .A1(n926), .A2(n925), .ZN(n927) );
  AND2_X1 U40bar ( .A1(n926bar), .A2(n925bar), .ZN(n927bar) );
  OR2_X1 U41 ( .A1(n924), .A2(n923), .ZN(n925) );
  AND2_X1 U41bar ( .A1(n924bar), .A2(n923bar), .ZN(n925bar) );
  OR2_X1 U42 ( .A1(n922), .A2(n921), .ZN(n923) );
  AND2_X1 U42bar ( .A1(n922bar), .A2(n921bar), .ZN(n923bar) );
  OR2_X1 U43 ( .A1(n940), .A2(n920), .ZN(n924) );
  AND2_X1 U43bar ( .A1(n940bar), .A2(n920bar), .ZN(n924bar) );
  OR2_X1 U44 ( .A1(in[111]), .A2(n919), .ZN(n920) );
  AND2_X1 U44bar ( .A1(inbar[111]), .A2(n919bar), .ZN(n920bar) );
  OR2_X1 U45 ( .A1(n918), .A2(n917), .ZN(n940) );
  AND2_X1 U45bar ( .A1(n918bar), .A2(n917bar), .ZN(n940bar) );
  OR2_X1 U46 ( .A1(n916), .A2(n915), .ZN(n917) );
  AND2_X1 U46bar ( .A1(n916bar), .A2(n915bar), .ZN(n917bar) );
  OR2_X1 U47 ( .A1(n914), .A2(n913), .ZN(n915) );
  AND2_X1 U47bar ( .A1(n914bar), .A2(n913bar), .ZN(n915bar) );
  OR2_X1 U48 ( .A1(in[140]), .A2(in[131]), .ZN(n913) );
  AND2_X1 U48bar ( .A1(inbar[140]), .A2(inbar[131]), .ZN(n913bar) );
  OR2_X1 U49 ( .A1(in[160]), .A2(in[144]), .ZN(n914) );
  AND2_X1 U49bar ( .A1(inbar[160]), .A2(inbar[144]), .ZN(n914bar) );
  OR2_X1 U50 ( .A1(n912), .A2(n911), .ZN(n916) );
  AND2_X1 U50bar ( .A1(n912bar), .A2(n911bar), .ZN(n916bar) );
  OR2_X1 U51 ( .A1(in[179]), .A2(in[174]), .ZN(n911) );
  AND2_X1 U51bar ( .A1(inbar[179]), .A2(inbar[174]), .ZN(n911bar) );
  OR2_X1 U52 ( .A1(in[188]), .A2(in[184]), .ZN(n912) );
  AND2_X1 U52bar ( .A1(inbar[188]), .A2(inbar[184]), .ZN(n912bar) );
  OR2_X1 U53 ( .A1(n910), .A2(n909), .ZN(n918) );
  AND2_X1 U53bar ( .A1(n910bar), .A2(n909bar), .ZN(n918bar) );
  OR2_X1 U54 ( .A1(n908), .A2(n907), .ZN(n909) );
  AND2_X1 U54bar ( .A1(n908bar), .A2(n907bar), .ZN(n909bar) );
  OR2_X1 U55 ( .A1(in[216]), .A2(in[200]), .ZN(n907) );
  AND2_X1 U55bar ( .A1(inbar[216]), .A2(inbar[200]), .ZN(n907bar) );
  OR2_X1 U56 ( .A1(in[228]), .A2(in[224]), .ZN(n908) );
  AND2_X1 U56bar ( .A1(inbar[228]), .A2(inbar[224]), .ZN(n908bar) );
  OR2_X1 U57 ( .A1(n906), .A2(n905), .ZN(n910) );
  AND2_X1 U57bar ( .A1(n906bar), .A2(n905bar), .ZN(n910bar) );
  OR2_X1 U58 ( .A1(in[247]), .A2(in[235]), .ZN(n905) );
  AND2_X1 U58bar ( .A1(inbar[247]), .A2(inbar[235]), .ZN(n905bar) );
  OR2_X1 U59 ( .A1(in_42), .A2(in[83]), .ZN(n906) );
  AND2_X1 U59bar ( .A1(in_42bar), .A2(inbar[83]), .ZN(n906bar) );
  OR2_X1 U60 ( .A1(n904), .A2(n903), .ZN(n926) );
  AND2_X1 U60bar ( .A1(n904bar), .A2(n903bar), .ZN(n926bar) );
  OR2_X1 U61 ( .A1(in[166]), .A2(in[123]), .ZN(n903) );
  AND2_X1 U61bar ( .A1(inbar[166]), .A2(inbar[123]), .ZN(n903bar) );
  OR2_X1 U62 ( .A1(in[170]), .A2(n902), .ZN(n904) );
  AND2_X1 U62bar ( .A1(inbar[170]), .A2(n902bar), .ZN(n904bar) );
  OR2_X1 U63 ( .A1(in[194]), .A2(in[183]), .ZN(n902) );
  AND2_X1 U63bar ( .A1(inbar[194]), .A2(inbar[183]), .ZN(n902bar) );
  OR2_X1 U64 ( .A1(n901), .A2(n900), .ZN(n928) );
  AND2_X1 U64bar ( .A1(n901bar), .A2(n900bar), .ZN(n928bar) );
  OR2_X1 U65 ( .A1(n899), .A2(n898), .ZN(n900) );
  AND2_X1 U65bar ( .A1(n899bar), .A2(n898bar), .ZN(n900bar) );
  OR2_X1 U66 ( .A1(in[241]), .A2(in[238]), .ZN(n898) );
  AND2_X1 U66bar ( .A1(inbar[241]), .A2(inbar[238]), .ZN(n898bar) );
  OR2_X1 U67 ( .A1(in[250]), .A2(n897), .ZN(n899) );
  AND2_X1 U67bar ( .A1(inbar[250]), .A2(n897bar), .ZN(n899bar) );
  OR2_X1 U68 ( .A1(in_24), .A2(in[84]), .ZN(n897) );
  AND2_X1 U68bar ( .A1(in_24bar), .A2(inbar[84]), .ZN(n897bar) );
  OR2_X1 U69 ( .A1(n896), .A2(n895), .ZN(n901) );
  AND2_X1 U69bar ( .A1(n896bar), .A2(n895bar), .ZN(n901bar) );
  OR2_X1 U70 ( .A1(in_41), .A2(in_29), .ZN(n895) );
  AND2_X1 U70bar ( .A1(in_41bar), .A2(in_29bar), .ZN(n895bar) );
  OR2_X1 U71 ( .A1(in_66), .A2(n894), .ZN(n896) );
  AND2_X1 U71bar ( .A1(in_66bar), .A2(n894bar), .ZN(n896bar) );
  OR2_X1 U72 ( .A1(in_76), .A2(in_71), .ZN(n894) );
  AND2_X1 U72bar ( .A1(in_76bar), .A2(in_71bar), .ZN(n894bar) );
  OR2_X1 U73 ( .A1(n893), .A2(n892), .ZN(out[4]) );
  AND2_X1 U73bar ( .A1(n893bar), .A2(n892bar), .ZN(outbar[4]) );
  OR2_X1 U74 ( .A1(n891), .A2(n890), .ZN(n892) );
  AND2_X1 U74bar ( .A1(n891bar), .A2(n890bar), .ZN(n892bar) );
  OR2_X1 U75 ( .A1(n889), .A2(n888), .ZN(n890) );
  AND2_X1 U75bar ( .A1(n889bar), .A2(n888bar), .ZN(n890bar) );
  OR2_X1 U76 ( .A1(n922), .A2(n887), .ZN(n888) );
  AND2_X1 U76bar ( .A1(n922bar), .A2(n887bar), .ZN(n888bar) );
  OR2_X1 U77 ( .A1(n886), .A2(n885), .ZN(n922) );
  AND2_X1 U77bar ( .A1(n886bar), .A2(n885bar), .ZN(n922bar) );
  OR2_X1 U78 ( .A1(n884), .A2(n883), .ZN(n885) );
  AND2_X1 U78bar ( .A1(n884bar), .A2(n883bar), .ZN(n885bar) );
  OR2_X1 U79 ( .A1(n882), .A2(n881), .ZN(n883) );
  AND2_X1 U79bar ( .A1(n882bar), .A2(n881bar), .ZN(n883bar) );
  OR2_X1 U80 ( .A1(in[118]), .A2(in[109]), .ZN(n881) );
  AND2_X1 U80bar ( .A1(inbar[118]), .A2(inbar[109]), .ZN(n881bar) );
  OR2_X1 U81 ( .A1(in[139]), .A2(in[120]), .ZN(n882) );
  AND2_X1 U81bar ( .A1(inbar[139]), .A2(inbar[120]), .ZN(n882bar) );
  OR2_X1 U82 ( .A1(n880), .A2(n879), .ZN(n884) );
  AND2_X1 U82bar ( .A1(n880bar), .A2(n879bar), .ZN(n884bar) );
  OR2_X1 U83 ( .A1(in[198]), .A2(in[154]), .ZN(n879) );
  AND2_X1 U83bar ( .A1(inbar[198]), .A2(inbar[154]), .ZN(n879bar) );
  OR2_X1 U84 ( .A1(in[210]), .A2(in[205]), .ZN(n880) );
  AND2_X1 U84bar ( .A1(inbar[210]), .A2(inbar[205]), .ZN(n880bar) );
  OR2_X1 U85 ( .A1(n878), .A2(n877), .ZN(n886) );
  AND2_X1 U85bar ( .A1(n878bar), .A2(n877bar), .ZN(n886bar) );
  OR2_X1 U86 ( .A1(n876), .A2(n875), .ZN(n877) );
  AND2_X1 U86bar ( .A1(n876bar), .A2(n875bar), .ZN(n877bar) );
  OR2_X1 U87 ( .A1(in[219]), .A2(in[217]), .ZN(n875) );
  AND2_X1 U87bar ( .A1(inbar[219]), .A2(inbar[217]), .ZN(n875bar) );
  OR2_X1 U88 ( .A1(in[86]), .A2(in[252]), .ZN(n876) );
  AND2_X1 U88bar ( .A1(inbar[86]), .A2(inbar[252]), .ZN(n876bar) );
  OR2_X1 U89 ( .A1(n874), .A2(n873), .ZN(n878) );
  AND2_X1 U89bar ( .A1(n874bar), .A2(n873bar), .ZN(n878bar) );
  OR2_X1 U90 ( .A1(in_40), .A2(in[91]), .ZN(n873) );
  AND2_X1 U90bar ( .A1(in_40bar), .A2(inbar[91]), .ZN(n873bar) );
  OR2_X1 U91 ( .A1(in_8), .A2(in_46), .ZN(n874) );
  AND2_X1 U91bar ( .A1(in_8bar), .A2(in_46bar), .ZN(n874bar) );
  OR2_X1 U92 ( .A1(n872), .A2(n871), .ZN(n889) );
  AND2_X1 U92bar ( .A1(n872bar), .A2(n871bar), .ZN(n889bar) );
  OR2_X1 U93 ( .A1(in[117]), .A2(n943), .ZN(n871) );
  AND2_X1 U93bar ( .A1(inbar[117]), .A2(n943bar), .ZN(n871bar) );
  OR2_X1 U94 ( .A1(n870), .A2(n869), .ZN(n943) );
  AND2_X1 U94bar ( .A1(n870bar), .A2(n869bar), .ZN(n943bar) );
  OR2_X1 U95 ( .A1(n868), .A2(n867), .ZN(n869) );
  AND2_X1 U95bar ( .A1(n868bar), .A2(n867bar), .ZN(n869bar) );
  OR2_X1 U96 ( .A1(n866), .A2(n865), .ZN(n867) );
  AND2_X1 U96bar ( .A1(n866bar), .A2(n865bar), .ZN(n867bar) );
  OR2_X1 U97 ( .A1(n864), .A2(n863), .ZN(n865) );
  AND2_X1 U97bar ( .A1(n864bar), .A2(n863bar), .ZN(n865bar) );
  OR2_X1 U98 ( .A1(in[108]), .A2(n919), .ZN(n866) );
  AND2_X1 U98bar ( .A1(inbar[108]), .A2(n919bar), .ZN(n866bar) );
  OR2_X1 U99 ( .A1(n862), .A2(n861), .ZN(n919) );
  AND2_X1 U99bar ( .A1(n862bar), .A2(n861bar), .ZN(n919bar) );
  OR2_X1 U100 ( .A1(n860), .A2(n859), .ZN(n861) );
  AND2_X1 U100bar ( .A1(n860bar), .A2(n859bar), .ZN(n861bar) );
  OR2_X1 U101 ( .A1(n858), .A2(n857), .ZN(n859) );
  AND2_X1 U101bar ( .A1(n858bar), .A2(n857bar), .ZN(n859bar) );
  OR2_X1 U102 ( .A1(in[119]), .A2(in[105]), .ZN(n857) );
  AND2_X1 U102bar ( .A1(inbar[119]), .A2(inbar[105]), .ZN(n857bar) );
  OR2_X1 U103 ( .A1(in[186]), .A2(in[175]), .ZN(n858) );
  AND2_X1 U103bar ( .A1(inbar[186]), .A2(inbar[175]), .ZN(n858bar) );
  OR2_X1 U104 ( .A1(n856), .A2(n855), .ZN(n860) );
  AND2_X1 U104bar ( .A1(n856bar), .A2(n855bar), .ZN(n860bar) );
  OR2_X1 U105 ( .A1(in[202]), .A2(in[193]), .ZN(n855) );
  AND2_X1 U105bar ( .A1(inbar[202]), .A2(inbar[193]), .ZN(n855bar) );
  OR2_X1 U106 ( .A1(in[225]), .A2(in[208]), .ZN(n856) );
  AND2_X1 U106bar ( .A1(inbar[225]), .A2(inbar[208]), .ZN(n856bar) );
  OR2_X1 U107 ( .A1(n854), .A2(n853), .ZN(n862) );
  AND2_X1 U107bar ( .A1(n854bar), .A2(n853bar), .ZN(n862bar) );
  OR2_X1 U108 ( .A1(n852), .A2(n851), .ZN(n853) );
  AND2_X1 U108bar ( .A1(n852bar), .A2(n851bar), .ZN(n853bar) );
  OR2_X1 U109 ( .A1(in_1), .A2(in[85]), .ZN(n851) );
  AND2_X1 U109bar ( .A1(in_1bar), .A2(inbar[85]), .ZN(n851bar) );
  OR2_X1 U110 ( .A1(in_23), .A2(in_19), .ZN(n852) );
  AND2_X1 U110bar ( .A1(in_23bar), .A2(in_19bar), .ZN(n852bar) );
  OR2_X1 U111 ( .A1(n850), .A2(n849), .ZN(n854) );
  AND2_X1 U111bar ( .A1(n850bar), .A2(n849bar), .ZN(n854bar) );
  OR2_X1 U112 ( .A1(in_43), .A2(in_33), .ZN(n849) );
  AND2_X1 U112bar ( .A1(in_43bar), .A2(in_33bar), .ZN(n849bar) );
  OR2_X1 U113 ( .A1(in_63), .A2(in_44), .ZN(n850) );
  AND2_X1 U113bar ( .A1(in_63bar), .A2(in_44bar), .ZN(n850bar) );
  OR2_X1 U114 ( .A1(n848), .A2(n847), .ZN(n868) );
  AND2_X1 U114bar ( .A1(n848bar), .A2(n847bar), .ZN(n868bar) );
  OR2_X1 U115 ( .A1(in[141]), .A2(in[112]), .ZN(n847) );
  AND2_X1 U115bar ( .A1(inbar[141]), .A2(inbar[112]), .ZN(n847bar) );
  OR2_X1 U116 ( .A1(in[147]), .A2(n846), .ZN(n848) );
  AND2_X1 U116bar ( .A1(inbar[147]), .A2(n846bar), .ZN(n848bar) );
  OR2_X1 U117 ( .A1(in[181]), .A2(in[167]), .ZN(n846) );
  AND2_X1 U117bar ( .A1(inbar[181]), .A2(inbar[167]), .ZN(n846bar) );
  OR2_X1 U118 ( .A1(n845), .A2(n844), .ZN(n870) );
  AND2_X1 U118bar ( .A1(n845bar), .A2(n844bar), .ZN(n870bar) );
  OR2_X1 U119 ( .A1(n843), .A2(n842), .ZN(n844) );
  AND2_X1 U119bar ( .A1(n843bar), .A2(n842bar), .ZN(n844bar) );
  OR2_X1 U120 ( .A1(in[229]), .A2(in[201]), .ZN(n842) );
  AND2_X1 U120bar ( .A1(inbar[229]), .A2(inbar[201]), .ZN(n842bar) );
  OR2_X1 U121 ( .A1(in[237]), .A2(n841), .ZN(n843) );
  AND2_X1 U121bar ( .A1(inbar[237]), .A2(n841bar), .ZN(n843bar) );
  OR2_X1 U122 ( .A1(in[94]), .A2(in[253]), .ZN(n841) );
  AND2_X1 U122bar ( .A1(inbar[94]), .A2(inbar[253]), .ZN(n841bar) );
  OR2_X1 U123 ( .A1(n840), .A2(n839), .ZN(n845) );
  AND2_X1 U123bar ( .A1(n840bar), .A2(n839bar), .ZN(n845bar) );
  OR2_X1 U124 ( .A1(in_21), .A2(in[96]), .ZN(n839) );
  AND2_X1 U124bar ( .A1(in_21bar), .A2(inbar[96]), .ZN(n839bar) );
  OR2_X1 U125 ( .A1(in_25), .A2(n838), .ZN(n840) );
  AND2_X1 U125bar ( .A1(in_25bar), .A2(n838bar), .ZN(n840bar) );
  OR2_X1 U126 ( .A1(in_81), .A2(in_45), .ZN(n838) );
  AND2_X1 U126bar ( .A1(in_81bar), .A2(in_45bar), .ZN(n838bar) );
  OR2_X1 U127 ( .A1(n837), .A2(n836), .ZN(n891) );
  AND2_X1 U127bar ( .A1(n837bar), .A2(n836bar), .ZN(n891bar) );
  OR2_X1 U128 ( .A1(in[142]), .A2(in[124]), .ZN(n836) );
  AND2_X1 U128bar ( .A1(inbar[142]), .A2(inbar[124]), .ZN(n836bar) );
  OR2_X1 U129 ( .A1(in[150]), .A2(n835), .ZN(n837) );
  AND2_X1 U129bar ( .A1(inbar[150]), .A2(n835bar), .ZN(n837bar) );
  OR2_X1 U130 ( .A1(in[172]), .A2(in[155]), .ZN(n835) );
  AND2_X1 U130bar ( .A1(inbar[172]), .A2(inbar[155]), .ZN(n835bar) );
  OR2_X1 U131 ( .A1(n834), .A2(n833), .ZN(n893) );
  AND2_X1 U131bar ( .A1(n834bar), .A2(n833bar), .ZN(n893bar) );
  OR2_X1 U132 ( .A1(n832), .A2(n831), .ZN(n833) );
  AND2_X1 U132bar ( .A1(n832bar), .A2(n831bar), .ZN(n833bar) );
  OR2_X1 U133 ( .A1(in[196]), .A2(in[173]), .ZN(n831) );
  AND2_X1 U133bar ( .A1(inbar[196]), .A2(inbar[173]), .ZN(n831bar) );
  OR2_X1 U134 ( .A1(in[222]), .A2(n830), .ZN(n832) );
  AND2_X1 U134bar ( .A1(inbar[222]), .A2(n830bar), .ZN(n832bar) );
  OR2_X1 U135 ( .A1(in[227]), .A2(in[226]), .ZN(n830) );
  AND2_X1 U135bar ( .A1(inbar[227]), .A2(inbar[226]), .ZN(n830bar) );
  OR2_X1 U136 ( .A1(n829), .A2(n828), .ZN(n834) );
  AND2_X1 U136bar ( .A1(n829bar), .A2(n828bar), .ZN(n834bar) );
  OR2_X1 U137 ( .A1(in[249]), .A2(in[231]), .ZN(n828) );
  AND2_X1 U137bar ( .A1(inbar[249]), .A2(inbar[231]), .ZN(n828bar) );
  OR2_X1 U138 ( .A1(in_28), .A2(n827), .ZN(n829) );
  AND2_X1 U138bar ( .A1(in_28bar), .A2(n827bar), .ZN(n829bar) );
  OR2_X1 U139 ( .A1(in_52), .A2(in_47), .ZN(n827) );
  AND2_X1 U139bar ( .A1(in_52bar), .A2(in_47bar), .ZN(n827bar) );
  OR2_X1 U140 ( .A1(n826), .A2(n825), .ZN(out[3]) );
  AND2_X1 U140bar ( .A1(n826bar), .A2(n825bar), .ZN(outbar[3]) );
  OR2_X1 U141 ( .A1(n824), .A2(n823), .ZN(n825) );
  AND2_X1 U141bar ( .A1(n824bar), .A2(n823bar), .ZN(n825bar) );
  OR2_X1 U142 ( .A1(n822), .A2(n821), .ZN(n823) );
  AND2_X1 U142bar ( .A1(n822bar), .A2(n821bar), .ZN(n823bar) );
  OR2_X1 U143 ( .A1(n820), .A2(n819), .ZN(n821) );
  AND2_X1 U143bar ( .A1(n820bar), .A2(n819bar), .ZN(n821bar) );
  OR2_X1 U144 ( .A1(n964), .A2(n818), .ZN(n822) );
  AND2_X1 U144bar ( .A1(n964bar), .A2(n818bar), .ZN(n822bar) );
  OR2_X1 U145 ( .A1(in[118]), .A2(n817), .ZN(n818) );
  AND2_X1 U145bar ( .A1(inbar[118]), .A2(n817bar), .ZN(n818bar) );
  OR2_X1 U146 ( .A1(n816), .A2(n815), .ZN(n964) );
  AND2_X1 U146bar ( .A1(n816bar), .A2(n815bar), .ZN(n964bar) );
  OR2_X1 U147 ( .A1(n814), .A2(n813), .ZN(n815) );
  AND2_X1 U147bar ( .A1(n814bar), .A2(n813bar), .ZN(n815bar) );
  OR2_X1 U148 ( .A1(n812), .A2(n811), .ZN(n813) );
  AND2_X1 U148bar ( .A1(n812bar), .A2(n811bar), .ZN(n813bar) );
  OR2_X1 U149 ( .A1(in[122]), .A2(in[111]), .ZN(n811) );
  AND2_X1 U149bar ( .A1(inbar[122]), .A2(inbar[111]), .ZN(n811bar) );
  OR2_X1 U150 ( .A1(in[154]), .A2(in[151]), .ZN(n812) );
  AND2_X1 U150bar ( .A1(inbar[154]), .A2(inbar[151]), .ZN(n812bar) );
  OR2_X1 U151 ( .A1(n810), .A2(n809), .ZN(n814) );
  AND2_X1 U151bar ( .A1(n810bar), .A2(n809bar), .ZN(n814bar) );
  OR2_X1 U152 ( .A1(in[187]), .A2(in[177]), .ZN(n809) );
  AND2_X1 U152bar ( .A1(inbar[187]), .A2(inbar[177]), .ZN(n809bar) );
  OR2_X1 U153 ( .A1(in[200]), .A2(in[192]), .ZN(n810) );
  AND2_X1 U153bar ( .A1(inbar[200]), .A2(inbar[192]), .ZN(n810bar) );
  OR2_X1 U154 ( .A1(n808), .A2(n807), .ZN(n816) );
  AND2_X1 U154bar ( .A1(n808bar), .A2(n807bar), .ZN(n816bar) );
  OR2_X1 U155 ( .A1(n806), .A2(n805), .ZN(n807) );
  AND2_X1 U155bar ( .A1(n806bar), .A2(n805bar), .ZN(n807bar) );
  OR2_X1 U156 ( .A1(in[225]), .A2(in[207]), .ZN(n805) );
  AND2_X1 U156bar ( .A1(inbar[225]), .A2(inbar[207]), .ZN(n805bar) );
  OR2_X1 U157 ( .A1(in[98]), .A2(in[226]), .ZN(n806) );
  AND2_X1 U157bar ( .A1(inbar[98]), .A2(inbar[226]), .ZN(n806bar) );
  OR2_X1 U158 ( .A1(n804), .A2(n803), .ZN(n808) );
  AND2_X1 U158bar ( .A1(n804bar), .A2(n803bar), .ZN(n808bar) );
  OR2_X1 U159 ( .A1(in_20), .A2(in_16), .ZN(n803) );
  AND2_X1 U159bar ( .A1(in_20bar), .A2(in_16bar), .ZN(n803bar) );
  OR2_X1 U160 ( .A1(in_55), .A2(in_45), .ZN(n804) );
  AND2_X1 U160bar ( .A1(in_55bar), .A2(in_45bar), .ZN(n804bar) );
  OR2_X1 U161 ( .A1(n802), .A2(n801), .ZN(n824) );
  AND2_X1 U161bar ( .A1(n802bar), .A2(n801bar), .ZN(n824bar) );
  OR2_X1 U162 ( .A1(in[162]), .A2(in[149]), .ZN(n801) );
  AND2_X1 U162bar ( .A1(inbar[162]), .A2(inbar[149]), .ZN(n801bar) );
  OR2_X1 U163 ( .A1(in[163]), .A2(n800), .ZN(n802) );
  AND2_X1 U163bar ( .A1(inbar[163]), .A2(n800bar), .ZN(n802bar) );
  OR2_X1 U164 ( .A1(in[191]), .A2(in[189]), .ZN(n800) );
  AND2_X1 U164bar ( .A1(inbar[191]), .A2(inbar[189]), .ZN(n800bar) );
  OR2_X1 U165 ( .A1(n799), .A2(n798), .ZN(n826) );
  AND2_X1 U165bar ( .A1(n799bar), .A2(n798bar), .ZN(n826bar) );
  OR2_X1 U166 ( .A1(n797), .A2(n796), .ZN(n798) );
  AND2_X1 U166bar ( .A1(n797bar), .A2(n796bar), .ZN(n798bar) );
  OR2_X1 U167 ( .A1(in[212]), .A2(in[193]), .ZN(n796) );
  AND2_X1 U167bar ( .A1(inbar[212]), .A2(inbar[193]), .ZN(n796bar) );
  OR2_X1 U168 ( .A1(in[238]), .A2(n795), .ZN(n797) );
  AND2_X1 U168bar ( .A1(inbar[238]), .A2(n795bar), .ZN(n797bar) );
  OR2_X1 U169 ( .A1(in[88]), .A2(in[247]), .ZN(n795) );
  AND2_X1 U169bar ( .A1(inbar[88]), .A2(inbar[247]), .ZN(n795bar) );
  OR2_X1 U170 ( .A1(n794), .A2(n793), .ZN(n799) );
  AND2_X1 U170bar ( .A1(n794bar), .A2(n793bar), .ZN(n799bar) );
  OR2_X1 U171 ( .A1(in[94]), .A2(in[92]), .ZN(n793) );
  AND2_X1 U171bar ( .A1(inbar[94]), .A2(inbar[92]), .ZN(n793bar) );
  OR2_X1 U172 ( .A1(in_52), .A2(n792), .ZN(n794) );
  AND2_X1 U172bar ( .A1(in_52bar), .A2(n792bar), .ZN(n794bar) );
  OR2_X1 U173 ( .A1(in_70), .A2(in_67), .ZN(n792) );
  AND2_X1 U173bar ( .A1(in_70bar), .A2(in_67bar), .ZN(n792bar) );
  OR2_X1 U174 ( .A1(n791), .A2(n790), .ZN(out[2]) );
  AND2_X1 U174bar ( .A1(n791bar), .A2(n790bar), .ZN(outbar[2]) );
  OR2_X1 U175 ( .A1(n789), .A2(n788), .ZN(n790) );
  AND2_X1 U175bar ( .A1(n789bar), .A2(n788bar), .ZN(n790bar) );
  OR2_X1 U176 ( .A1(n787), .A2(n786), .ZN(n788) );
  AND2_X1 U176bar ( .A1(n787bar), .A2(n786bar), .ZN(n788bar) );
  OR2_X1 U177 ( .A1(n819), .A2(n785), .ZN(n786) );
  AND2_X1 U177bar ( .A1(n819bar), .A2(n785bar), .ZN(n786bar) );
  OR2_X1 U178 ( .A1(n784), .A2(n783), .ZN(n819) );
  AND2_X1 U178bar ( .A1(n784bar), .A2(n783bar), .ZN(n819bar) );
  OR2_X1 U179 ( .A1(n782), .A2(n781), .ZN(n783) );
  AND2_X1 U179bar ( .A1(n782bar), .A2(n781bar), .ZN(n783bar) );
  OR2_X1 U180 ( .A1(n780), .A2(n779), .ZN(n781) );
  AND2_X1 U180bar ( .A1(n780bar), .A2(n779bar), .ZN(n781bar) );
  OR2_X1 U181 ( .A1(n962), .A2(n778), .ZN(n779) );
  AND2_X1 U181bar ( .A1(n962bar), .A2(n778bar), .ZN(n779bar) );
  OR2_X1 U182 ( .A1(n777), .A2(n776), .ZN(n962) );
  AND2_X1 U182bar ( .A1(n777bar), .A2(n776bar), .ZN(n962bar) );
  OR2_X1 U183 ( .A1(n775), .A2(n774), .ZN(n776) );
  AND2_X1 U183bar ( .A1(n775bar), .A2(n774bar), .ZN(n776bar) );
  OR2_X1 U184 ( .A1(n773), .A2(n772), .ZN(n774) );
  AND2_X1 U184bar ( .A1(n773bar), .A2(n772bar), .ZN(n774bar) );
  OR2_X1 U185 ( .A1(in[131]), .A2(in[120]), .ZN(n772) );
  AND2_X1 U185bar ( .A1(inbar[131]), .A2(inbar[120]), .ZN(n772bar) );
  OR2_X1 U186 ( .A1(in[153]), .A2(in[147]), .ZN(n773) );
  AND2_X1 U186bar ( .A1(inbar[153]), .A2(inbar[147]), .ZN(n773bar) );
  OR2_X1 U187 ( .A1(n771), .A2(n770), .ZN(n775) );
  AND2_X1 U187bar ( .A1(n771bar), .A2(n770bar), .ZN(n775bar) );
  OR2_X1 U188 ( .A1(in[170]), .A2(in[156]), .ZN(n770) );
  AND2_X1 U188bar ( .A1(inbar[170]), .A2(inbar[156]), .ZN(n770bar) );
  OR2_X1 U189 ( .A1(in[223]), .A2(in[190]), .ZN(n771) );
  AND2_X1 U189bar ( .A1(inbar[223]), .A2(inbar[190]), .ZN(n771bar) );
  OR2_X1 U190 ( .A1(n769), .A2(n768), .ZN(n777) );
  AND2_X1 U190bar ( .A1(n769bar), .A2(n768bar), .ZN(n777bar) );
  OR2_X1 U191 ( .A1(n767), .A2(n766), .ZN(n768) );
  AND2_X1 U191bar ( .A1(n767bar), .A2(n766bar), .ZN(n768bar) );
  OR2_X1 U192 ( .A1(in[236]), .A2(in[230]), .ZN(n766) );
  AND2_X1 U192bar ( .A1(inbar[236]), .A2(inbar[230]), .ZN(n766bar) );
  OR2_X1 U193 ( .A1(in[85]), .A2(in[240]), .ZN(n767) );
  AND2_X1 U193bar ( .A1(inbar[85]), .A2(inbar[240]), .ZN(n767bar) );
  OR2_X1 U194 ( .A1(n765), .A2(n764), .ZN(n769) );
  AND2_X1 U194bar ( .A1(n765bar), .A2(n764bar), .ZN(n769bar) );
  OR2_X1 U195 ( .A1(in_12), .A2(in[90]), .ZN(n764) );
  AND2_X1 U195bar ( .A1(in_12bar), .A2(inbar[90]), .ZN(n764bar) );
  OR2_X1 U196 ( .A1(in_39), .A2(in_28), .ZN(n765) );
  AND2_X1 U196bar ( .A1(in_39bar), .A2(in_28bar), .ZN(n765bar) );
  OR2_X1 U197 ( .A1(in[109]), .A2(n763), .ZN(n780) );
  AND2_X1 U197bar ( .A1(inbar[109]), .A2(n763bar), .ZN(n780bar) );
  OR2_X1 U198 ( .A1(n762), .A2(n761), .ZN(n782) );
  AND2_X1 U198bar ( .A1(n762bar), .A2(n761bar), .ZN(n782bar) );
  OR2_X1 U199 ( .A1(in[138]), .A2(in[129]), .ZN(n761) );
  AND2_X1 U199bar ( .A1(inbar[138]), .A2(inbar[129]), .ZN(n761bar) );
  OR2_X1 U200 ( .A1(in[157]), .A2(n760), .ZN(n762) );
  AND2_X1 U200bar ( .A1(inbar[157]), .A2(n760bar), .ZN(n762bar) );
  OR2_X1 U201 ( .A1(in[182]), .A2(in[167]), .ZN(n760) );
  AND2_X1 U201bar ( .A1(inbar[182]), .A2(inbar[167]), .ZN(n760bar) );
  OR2_X1 U202 ( .A1(n759), .A2(n758), .ZN(n784) );
  AND2_X1 U202bar ( .A1(n759bar), .A2(n758bar), .ZN(n784bar) );
  OR2_X1 U203 ( .A1(n757), .A2(n756), .ZN(n758) );
  AND2_X1 U203bar ( .A1(n757bar), .A2(n756bar), .ZN(n758bar) );
  OR2_X1 U204 ( .A1(in[195]), .A2(in[184]), .ZN(n756) );
  AND2_X1 U204bar ( .A1(inbar[195]), .A2(inbar[184]), .ZN(n756bar) );
  OR2_X1 U205 ( .A1(in[196]), .A2(n755), .ZN(n757) );
  AND2_X1 U205bar ( .A1(inbar[196]), .A2(n755bar), .ZN(n757bar) );
  OR2_X1 U206 ( .A1(in[215]), .A2(in[209]), .ZN(n755) );
  AND2_X1 U206bar ( .A1(inbar[215]), .A2(inbar[209]), .ZN(n755bar) );
  OR2_X1 U207 ( .A1(n754), .A2(n753), .ZN(n759) );
  AND2_X1 U207bar ( .A1(n754bar), .A2(n753bar), .ZN(n759bar) );
  OR2_X1 U208 ( .A1(in[93]), .A2(in[233]), .ZN(n753) );
  AND2_X1 U208bar ( .A1(inbar[93]), .A2(inbar[233]), .ZN(n753bar) );
  OR2_X1 U209 ( .A1(in_1), .A2(n752), .ZN(n754) );
  AND2_X1 U209bar ( .A1(in_1bar), .A2(n752bar), .ZN(n754bar) );
  OR2_X1 U210 ( .A1(in_69), .A2(in_66), .ZN(n752) );
  AND2_X1 U210bar ( .A1(in_69bar), .A2(in_66bar), .ZN(n752bar) );
  OR2_X1 U211 ( .A1(n966), .A2(n751), .ZN(n787) );
  AND2_X1 U211bar ( .A1(n966bar), .A2(n751bar), .ZN(n787bar) );
  OR2_X1 U212 ( .A1(in[134]), .A2(n750), .ZN(n751) );
  AND2_X1 U212bar ( .A1(inbar[134]), .A2(n750bar), .ZN(n751bar) );
  OR2_X1 U213 ( .A1(n749), .A2(n748), .ZN(n966) );
  AND2_X1 U213bar ( .A1(n749bar), .A2(n748bar), .ZN(n966bar) );
  OR2_X1 U214 ( .A1(n747), .A2(n746), .ZN(n748) );
  AND2_X1 U214bar ( .A1(n747bar), .A2(n746bar), .ZN(n748bar) );
  OR2_X1 U215 ( .A1(n745), .A2(n744), .ZN(n746) );
  AND2_X1 U215bar ( .A1(n745bar), .A2(n744bar), .ZN(n746bar) );
  OR2_X1 U216 ( .A1(in[136]), .A2(in[121]), .ZN(n744) );
  AND2_X1 U216bar ( .A1(inbar[136]), .A2(inbar[121]), .ZN(n744bar) );
  OR2_X1 U217 ( .A1(in[186]), .A2(in[174]), .ZN(n745) );
  AND2_X1 U217bar ( .A1(inbar[186]), .A2(inbar[174]), .ZN(n745bar) );
  OR2_X1 U218 ( .A1(n743), .A2(n742), .ZN(n747) );
  AND2_X1 U218bar ( .A1(n743bar), .A2(n742bar), .ZN(n747bar) );
  OR2_X1 U219 ( .A1(in[198]), .A2(in[197]), .ZN(n742) );
  AND2_X1 U219bar ( .A1(inbar[198]), .A2(inbar[197]), .ZN(n742bar) );
  OR2_X1 U220 ( .A1(in[214]), .A2(in[199]), .ZN(n743) );
  AND2_X1 U220bar ( .A1(inbar[214]), .A2(inbar[199]), .ZN(n743bar) );
  OR2_X1 U221 ( .A1(n741), .A2(n740), .ZN(n749) );
  AND2_X1 U221bar ( .A1(n741bar), .A2(n740bar), .ZN(n749bar) );
  OR2_X1 U222 ( .A1(n739), .A2(n738), .ZN(n740) );
  AND2_X1 U222bar ( .A1(n739bar), .A2(n738bar), .ZN(n740bar) );
  OR2_X1 U223 ( .A1(in[231]), .A2(in[220]), .ZN(n738) );
  AND2_X1 U223bar ( .A1(inbar[231]), .A2(inbar[220]), .ZN(n738bar) );
  OR2_X1 U224 ( .A1(in_25), .A2(in[245]), .ZN(n739) );
  AND2_X1 U224bar ( .A1(in_25bar), .A2(inbar[245]), .ZN(n739bar) );
  OR2_X1 U225 ( .A1(n737), .A2(n736), .ZN(n741) );
  AND2_X1 U225bar ( .A1(n737bar), .A2(n736bar), .ZN(n741bar) );
  OR2_X1 U226 ( .A1(in_53), .A2(in_29), .ZN(n736) );
  AND2_X1 U226bar ( .A1(in_53bar), .A2(in_29bar), .ZN(n736bar) );
  OR2_X1 U227 ( .A1(in_79), .A2(in_74), .ZN(n737) );
  AND2_X1 U227bar ( .A1(in_79bar), .A2(in_74bar), .ZN(n737bar) );
  OR2_X1 U228 ( .A1(n735), .A2(n734), .ZN(n789) );
  AND2_X1 U228bar ( .A1(n735bar), .A2(n734bar), .ZN(n789bar) );
  OR2_X1 U229 ( .A1(in[152]), .A2(in[140]), .ZN(n734) );
  AND2_X1 U229bar ( .A1(inbar[152]), .A2(inbar[140]), .ZN(n734bar) );
  OR2_X1 U230 ( .A1(in[155]), .A2(n733), .ZN(n735) );
  AND2_X1 U230bar ( .A1(inbar[155]), .A2(n733bar), .ZN(n735bar) );
  OR2_X1 U231 ( .A1(in[166]), .A2(in[165]), .ZN(n733) );
  AND2_X1 U231bar ( .A1(inbar[166]), .A2(inbar[165]), .ZN(n733bar) );
  OR2_X1 U232 ( .A1(n732), .A2(n731), .ZN(n791) );
  AND2_X1 U232bar ( .A1(n732bar), .A2(n731bar), .ZN(n791bar) );
  OR2_X1 U233 ( .A1(n730), .A2(n729), .ZN(n731) );
  AND2_X1 U233bar ( .A1(n730bar), .A2(n729bar), .ZN(n731bar) );
  OR2_X1 U234 ( .A1(in[202]), .A2(in[185]), .ZN(n729) );
  AND2_X1 U234bar ( .A1(inbar[202]), .A2(inbar[185]), .ZN(n729bar) );
  OR2_X1 U235 ( .A1(in[211]), .A2(n728), .ZN(n730) );
  AND2_X1 U235bar ( .A1(inbar[211]), .A2(n728bar), .ZN(n730bar) );
  OR2_X1 U236 ( .A1(in[255]), .A2(in[253]), .ZN(n728) );
  AND2_X1 U236bar ( .A1(inbar[255]), .A2(inbar[253]), .ZN(n728bar) );
  OR2_X1 U237 ( .A1(n727), .A2(n726), .ZN(n732) );
  AND2_X1 U237bar ( .A1(n727bar), .A2(n726bar), .ZN(n732bar) );
  OR2_X1 U238 ( .A1(in_35), .A2(in_15), .ZN(n726) );
  AND2_X1 U238bar ( .A1(in_35bar), .A2(in_15bar), .ZN(n726bar) );
  OR2_X1 U239 ( .A1(in_36), .A2(n725), .ZN(n727) );
  AND2_X1 U239bar ( .A1(in_36bar), .A2(n725bar), .ZN(n727bar) );
  OR2_X1 U240 ( .A1(in_48), .A2(in_40), .ZN(n725) );
  AND2_X1 U240bar ( .A1(in_48bar), .A2(in_40bar), .ZN(n725bar) );
  OR2_X1 U241 ( .A1(n724), .A2(n723), .ZN(out[1]) );
  AND2_X1 U241bar ( .A1(n724bar), .A2(n723bar), .ZN(outbar[1]) );
  OR2_X1 U242 ( .A1(n722), .A2(n721), .ZN(n723) );
  AND2_X1 U242bar ( .A1(n722bar), .A2(n721bar), .ZN(n723bar) );
  OR2_X1 U243 ( .A1(n720), .A2(n719), .ZN(n721) );
  AND2_X1 U243bar ( .A1(n720bar), .A2(n719bar), .ZN(n721bar) );
  OR2_X1 U244 ( .A1(n921), .A2(n887), .ZN(n719) );
  AND2_X1 U244bar ( .A1(n921bar), .A2(n887bar), .ZN(n719bar) );
  OR2_X1 U245 ( .A1(n718), .A2(n717), .ZN(n887) );
  AND2_X1 U245bar ( .A1(n718bar), .A2(n717bar), .ZN(n887bar) );
  OR2_X1 U246 ( .A1(n716), .A2(n715), .ZN(n717) );
  AND2_X1 U246bar ( .A1(n716bar), .A2(n715bar), .ZN(n717bar) );
  OR2_X1 U247 ( .A1(n714), .A2(n713), .ZN(n715) );
  AND2_X1 U247bar ( .A1(n714bar), .A2(n713bar), .ZN(n715bar) );
  OR2_X1 U248 ( .A1(in[116]), .A2(in[110]), .ZN(n713) );
  AND2_X1 U248bar ( .A1(inbar[116]), .A2(inbar[110]), .ZN(n713bar) );
  OR2_X1 U249 ( .A1(in[133]), .A2(in[130]), .ZN(n714) );
  AND2_X1 U249bar ( .A1(inbar[133]), .A2(inbar[130]), .ZN(n714bar) );
  OR2_X1 U250 ( .A1(n712), .A2(n711), .ZN(n716) );
  AND2_X1 U250bar ( .A1(n712bar), .A2(n711bar), .ZN(n716bar) );
  OR2_X1 U251 ( .A1(in[203]), .A2(in[135]), .ZN(n711) );
  AND2_X1 U251bar ( .A1(inbar[203]), .A2(inbar[135]), .ZN(n711bar) );
  OR2_X1 U252 ( .A1(in[232]), .A2(in[223]), .ZN(n712) );
  AND2_X1 U252bar ( .A1(inbar[232]), .A2(inbar[223]), .ZN(n712bar) );
  OR2_X1 U253 ( .A1(n710), .A2(n709), .ZN(n718) );
  AND2_X1 U253bar ( .A1(n710bar), .A2(n709bar), .ZN(n718bar) );
  OR2_X1 U254 ( .A1(n708), .A2(n707), .ZN(n709) );
  AND2_X1 U254bar ( .A1(n708bar), .A2(n707bar), .ZN(n709bar) );
  OR2_X1 U255 ( .A1(in[255]), .A2(in[233]), .ZN(n707) );
  AND2_X1 U255bar ( .A1(inbar[255]), .A2(inbar[233]), .ZN(n707bar) );
  OR2_X1 U256 ( .A1(in_53), .A2(in_34), .ZN(n708) );
  AND2_X1 U256bar ( .A1(in_53bar), .A2(in_34bar), .ZN(n708bar) );
  OR2_X1 U257 ( .A1(n706), .A2(n705), .ZN(n710) );
  AND2_X1 U257bar ( .A1(n706bar), .A2(n705bar), .ZN(n710bar) );
  OR2_X1 U258 ( .A1(in_57), .A2(in_55), .ZN(n705) );
  AND2_X1 U258bar ( .A1(in_57bar), .A2(in_55bar), .ZN(n705bar) );
  OR2_X1 U259 ( .A1(in_68), .A2(in_67), .ZN(n706) );
  AND2_X1 U259bar ( .A1(in_68bar), .A2(in_67bar), .ZN(n706bar) );
  OR2_X1 U260 ( .A1(n704), .A2(n703), .ZN(n921) );
  AND2_X1 U260bar ( .A1(n704bar), .A2(n703bar), .ZN(n921bar) );
  OR2_X1 U261 ( .A1(n702), .A2(n701), .ZN(n703) );
  AND2_X1 U261bar ( .A1(n702bar), .A2(n701bar), .ZN(n703bar) );
  OR2_X1 U262 ( .A1(n700), .A2(n699), .ZN(n701) );
  AND2_X1 U262bar ( .A1(n700bar), .A2(n699bar), .ZN(n701bar) );
  OR2_X1 U263 ( .A1(n944), .A2(n872), .ZN(n699) );
  AND2_X1 U263bar ( .A1(n944bar), .A2(n872bar), .ZN(n699bar) );
  OR2_X1 U264 ( .A1(n698), .A2(n697), .ZN(n872) );
  AND2_X1 U264bar ( .A1(n698bar), .A2(n697bar), .ZN(n872bar) );
  OR2_X1 U265 ( .A1(n696), .A2(n695), .ZN(n697) );
  AND2_X1 U265bar ( .A1(n696bar), .A2(n695bar), .ZN(n697bar) );
  OR2_X1 U266 ( .A1(n694), .A2(n693), .ZN(n695) );
  AND2_X1 U266bar ( .A1(n694bar), .A2(n693bar), .ZN(n695bar) );
  OR2_X1 U267 ( .A1(in[121]), .A2(in[102]), .ZN(n693) );
  AND2_X1 U267bar ( .A1(inbar[121]), .A2(inbar[102]), .ZN(n693bar) );
  OR2_X1 U268 ( .A1(in[162]), .A2(in[161]), .ZN(n694) );
  AND2_X1 U268bar ( .A1(inbar[162]), .A2(inbar[161]), .ZN(n694bar) );
  OR2_X1 U269 ( .A1(n692), .A2(n691), .ZN(n696) );
  AND2_X1 U269bar ( .A1(n692bar), .A2(n691bar), .ZN(n696bar) );
  OR2_X1 U270 ( .A1(in[192]), .A2(in[178]), .ZN(n691) );
  AND2_X1 U270bar ( .A1(inbar[192]), .A2(inbar[178]), .ZN(n691bar) );
  OR2_X1 U271 ( .A1(in[244]), .A2(in[209]), .ZN(n692) );
  AND2_X1 U271bar ( .A1(inbar[244]), .A2(inbar[209]), .ZN(n692bar) );
  OR2_X1 U272 ( .A1(n690), .A2(n689), .ZN(n698) );
  AND2_X1 U272bar ( .A1(n690bar), .A2(n689bar), .ZN(n698bar) );
  OR2_X1 U273 ( .A1(n688), .A2(n687), .ZN(n689) );
  AND2_X1 U273bar ( .A1(n688bar), .A2(n687bar), .ZN(n689bar) );
  OR2_X1 U274 ( .A1(in[90]), .A2(in[254]), .ZN(n687) );
  AND2_X1 U274bar ( .A1(inbar[90]), .A2(inbar[254]), .ZN(n687bar) );
  OR2_X1 U275 ( .A1(in_36), .A2(in_32), .ZN(n688) );
  AND2_X1 U275bar ( .A1(in_36bar), .A2(in_32bar), .ZN(n688bar) );
  OR2_X1 U276 ( .A1(n686), .A2(n685), .ZN(n690) );
  AND2_X1 U276bar ( .A1(n686bar), .A2(n685bar), .ZN(n690bar) );
  OR2_X1 U277 ( .A1(in_62), .A2(in_37), .ZN(n685) );
  AND2_X1 U277bar ( .A1(in_62bar), .A2(in_37bar), .ZN(n685bar) );
  OR2_X1 U278 ( .A1(in_75), .A2(in_73), .ZN(n686) );
  AND2_X1 U278bar ( .A1(in_75bar), .A2(in_73bar), .ZN(n686bar) );
  OR2_X1 U279 ( .A1(n684), .A2(n683), .ZN(n944) );
  AND2_X1 U279bar ( .A1(n684bar), .A2(n683bar), .ZN(n944bar) );
  OR2_X1 U280 ( .A1(n682), .A2(n681), .ZN(n683) );
  AND2_X1 U280bar ( .A1(n682bar), .A2(n681bar), .ZN(n683bar) );
  OR2_X1 U281 ( .A1(n680), .A2(n679), .ZN(n681) );
  AND2_X1 U281bar ( .A1(n680bar), .A2(n679bar), .ZN(n681bar) );
  OR2_X1 U282 ( .A1(in[171]), .A2(in[153]), .ZN(n679) );
  AND2_X1 U282bar ( .A1(inbar[171]), .A2(inbar[153]), .ZN(n679bar) );
  OR2_X1 U283 ( .A1(in[187]), .A2(in[176]), .ZN(n680) );
  AND2_X1 U283bar ( .A1(inbar[187]), .A2(inbar[176]), .ZN(n680bar) );
  OR2_X1 U284 ( .A1(n678), .A2(n677), .ZN(n682) );
  AND2_X1 U284bar ( .A1(n678bar), .A2(n677bar), .ZN(n682bar) );
  OR2_X1 U285 ( .A1(in[245]), .A2(in[211]), .ZN(n677) );
  AND2_X1 U285bar ( .A1(inbar[245]), .A2(inbar[211]), .ZN(n677bar) );
  OR2_X1 U286 ( .A1(in[97]), .A2(in[88]), .ZN(n678) );
  AND2_X1 U286bar ( .A1(inbar[97]), .A2(inbar[88]), .ZN(n678bar) );
  OR2_X1 U287 ( .A1(n676), .A2(n675), .ZN(n684) );
  AND2_X1 U287bar ( .A1(n676bar), .A2(n675bar), .ZN(n684bar) );
  OR2_X1 U288 ( .A1(n674), .A2(n673), .ZN(n675) );
  AND2_X1 U288bar ( .A1(n674bar), .A2(n673bar), .ZN(n675bar) );
  OR2_X1 U289 ( .A1(in_10), .A2(in_0), .ZN(n673) );
  AND2_X1 U289bar ( .A1(in_10bar), .A2(in_0bar), .ZN(n673bar) );
  OR2_X1 U290 ( .A1(in_59), .A2(in_5), .ZN(n674) );
  AND2_X1 U290bar ( .A1(in_59bar), .A2(in_5bar), .ZN(n674bar) );
  OR2_X1 U291 ( .A1(n672), .A2(n671), .ZN(n676) );
  AND2_X1 U291bar ( .A1(n672bar), .A2(n671bar), .ZN(n676bar) );
  OR2_X1 U292 ( .A1(in_60), .A2(in_6), .ZN(n671) );
  AND2_X1 U292bar ( .A1(in_60bar), .A2(in_6bar), .ZN(n671bar) );
  OR2_X1 U293 ( .A1(in_77), .A2(in_69), .ZN(n672) );
  AND2_X1 U293bar ( .A1(in_77bar), .A2(in_69bar), .ZN(n672bar) );
  OR2_X1 U294 ( .A1(in[113]), .A2(n864), .ZN(n700) );
  AND2_X1 U294bar ( .A1(inbar[113]), .A2(n864bar), .ZN(n700bar) );
  OR2_X1 U295 ( .A1(n670), .A2(n669), .ZN(n864) );
  AND2_X1 U295bar ( .A1(n670bar), .A2(n669bar), .ZN(n864bar) );
  OR2_X1 U296 ( .A1(n668), .A2(n667), .ZN(n669) );
  AND2_X1 U296bar ( .A1(n668bar), .A2(n667bar), .ZN(n669bar) );
  OR2_X1 U297 ( .A1(n666), .A2(n665), .ZN(n667) );
  AND2_X1 U297bar ( .A1(n666bar), .A2(n665bar), .ZN(n667bar) );
  OR2_X1 U298 ( .A1(in[125]), .A2(in[107]), .ZN(n665) );
  AND2_X1 U298bar ( .A1(inbar[125]), .A2(inbar[107]), .ZN(n665bar) );
  OR2_X1 U299 ( .A1(in[138]), .A2(in[126]), .ZN(n666) );
  AND2_X1 U299bar ( .A1(inbar[138]), .A2(inbar[126]), .ZN(n666bar) );
  OR2_X1 U300 ( .A1(n664), .A2(n663), .ZN(n668) );
  AND2_X1 U300bar ( .A1(n664bar), .A2(n663bar), .ZN(n668bar) );
  OR2_X1 U301 ( .A1(in[189]), .A2(in[143]), .ZN(n663) );
  AND2_X1 U301bar ( .A1(inbar[189]), .A2(inbar[143]), .ZN(n663bar) );
  OR2_X1 U302 ( .A1(in[99]), .A2(in[214]), .ZN(n664) );
  AND2_X1 U302bar ( .A1(inbar[99]), .A2(inbar[214]), .ZN(n664bar) );
  OR2_X1 U303 ( .A1(n662), .A2(n661), .ZN(n670) );
  AND2_X1 U303bar ( .A1(n662bar), .A2(n661bar), .ZN(n670bar) );
  OR2_X1 U304 ( .A1(n660), .A2(n659), .ZN(n661) );
  AND2_X1 U304bar ( .A1(n660bar), .A2(n659bar), .ZN(n661bar) );
  OR2_X1 U305 ( .A1(in_15), .A2(in_12), .ZN(n659) );
  AND2_X1 U305bar ( .A1(in_15bar), .A2(in_12bar), .ZN(n659bar) );
  OR2_X1 U306 ( .A1(in_20), .A2(in_2), .ZN(n660) );
  AND2_X1 U306bar ( .A1(in_20bar), .A2(in_2bar), .ZN(n660bar) );
  OR2_X1 U307 ( .A1(n658), .A2(n657), .ZN(n662) );
  AND2_X1 U307bar ( .A1(n658bar), .A2(n657bar), .ZN(n662bar) );
  OR2_X1 U308 ( .A1(in_30), .A2(in_3), .ZN(n657) );
  AND2_X1 U308bar ( .A1(in_30bar), .A2(in_3bar), .ZN(n657bar) );
  OR2_X1 U309 ( .A1(in_4), .A2(in_38), .ZN(n658) );
  AND2_X1 U309bar ( .A1(in_4bar), .A2(in_38bar), .ZN(n658bar) );
  OR2_X1 U310 ( .A1(n656), .A2(n655), .ZN(n702) );
  AND2_X1 U310bar ( .A1(n656bar), .A2(n655bar), .ZN(n702bar) );
  OR2_X1 U311 ( .A1(in[148]), .A2(in[137]), .ZN(n655) );
  AND2_X1 U311bar ( .A1(inbar[148]), .A2(inbar[137]), .ZN(n655bar) );
  OR2_X1 U312 ( .A1(in[149]), .A2(n654), .ZN(n656) );
  AND2_X1 U312bar ( .A1(inbar[149]), .A2(n654bar), .ZN(n656bar) );
  OR2_X1 U313 ( .A1(in[195]), .A2(in[190]), .ZN(n654) );
  AND2_X1 U313bar ( .A1(inbar[195]), .A2(inbar[190]), .ZN(n654bar) );
  OR2_X1 U314 ( .A1(n653), .A2(n652), .ZN(n704) );
  AND2_X1 U314bar ( .A1(n653bar), .A2(n652bar), .ZN(n704bar) );
  OR2_X1 U315 ( .A1(n651), .A2(n650), .ZN(n652) );
  AND2_X1 U315bar ( .A1(n651bar), .A2(n650bar), .ZN(n652bar) );
  OR2_X1 U316 ( .A1(in[98]), .A2(in[197]), .ZN(n650) );
  AND2_X1 U316bar ( .A1(inbar[98]), .A2(inbar[197]), .ZN(n650bar) );
  OR2_X1 U317 ( .A1(in_11), .A2(n649), .ZN(n651) );
  AND2_X1 U317bar ( .A1(in_11bar), .A2(n649bar), .ZN(n651bar) );
  OR2_X1 U318 ( .A1(in_26), .A2(in_14), .ZN(n649) );
  AND2_X1 U318bar ( .A1(in_26bar), .A2(in_14bar), .ZN(n649bar) );
  OR2_X1 U319 ( .A1(n648), .A2(n647), .ZN(n653) );
  AND2_X1 U319bar ( .A1(n648bar), .A2(n647bar), .ZN(n653bar) );
  OR2_X1 U320 ( .A1(in_35), .A2(in_27), .ZN(n647) );
  AND2_X1 U320bar ( .A1(in_35bar), .A2(in_27bar), .ZN(n647bar) );
  OR2_X1 U321 ( .A1(in_50), .A2(n646), .ZN(n648) );
  AND2_X1 U321bar ( .A1(in_50bar), .A2(n646bar), .ZN(n648bar) );
  OR2_X1 U322 ( .A1(in_78), .A2(in_61), .ZN(n646) );
  AND2_X1 U322bar ( .A1(in_78bar), .A2(in_61bar), .ZN(n646bar) );
  OR2_X1 U323 ( .A1(n942), .A2(n645), .ZN(n720) );
  AND2_X1 U323bar ( .A1(n942bar), .A2(n645bar), .ZN(n720bar) );
  OR2_X1 U324 ( .A1(in[106]), .A2(n863), .ZN(n645) );
  AND2_X1 U324bar ( .A1(inbar[106]), .A2(n863bar), .ZN(n645bar) );
  OR2_X1 U325 ( .A1(n644), .A2(n643), .ZN(n863) );
  AND2_X1 U325bar ( .A1(n644bar), .A2(n643bar), .ZN(n863bar) );
  OR2_X1 U326 ( .A1(n642), .A2(n641), .ZN(n643) );
  AND2_X1 U326bar ( .A1(n642bar), .A2(n641bar), .ZN(n643bar) );
  OR2_X1 U327 ( .A1(n640), .A2(n639), .ZN(n641) );
  AND2_X1 U327bar ( .A1(n640bar), .A2(n639bar), .ZN(n641bar) );
  OR2_X1 U328 ( .A1(in[127]), .A2(in[122]), .ZN(n639) );
  AND2_X1 U328bar ( .A1(inbar[127]), .A2(inbar[122]), .ZN(n639bar) );
  OR2_X1 U329 ( .A1(in[156]), .A2(in[132]), .ZN(n640) );
  AND2_X1 U329bar ( .A1(inbar[156]), .A2(inbar[132]), .ZN(n640bar) );
  OR2_X1 U330 ( .A1(n638), .A2(n637), .ZN(n642) );
  AND2_X1 U330bar ( .A1(n638bar), .A2(n637bar), .ZN(n642bar) );
  OR2_X1 U331 ( .A1(in[159]), .A2(in[157]), .ZN(n637) );
  AND2_X1 U331bar ( .A1(inbar[159]), .A2(inbar[157]), .ZN(n637bar) );
  OR2_X1 U332 ( .A1(in[185]), .A2(in[169]), .ZN(n638) );
  AND2_X1 U332bar ( .A1(inbar[185]), .A2(inbar[169]), .ZN(n638bar) );
  OR2_X1 U333 ( .A1(n636), .A2(n635), .ZN(n644) );
  AND2_X1 U333bar ( .A1(n636bar), .A2(n635bar), .ZN(n644bar) );
  OR2_X1 U334 ( .A1(n634), .A2(n633), .ZN(n635) );
  AND2_X1 U334bar ( .A1(n634bar), .A2(n633bar), .ZN(n635bar) );
  OR2_X1 U335 ( .A1(in[239]), .A2(in[218]), .ZN(n633) );
  AND2_X1 U335bar ( .A1(inbar[239]), .A2(inbar[218]), .ZN(n633bar) );
  OR2_X1 U336 ( .A1(in_13), .A2(in[87]), .ZN(n634) );
  AND2_X1 U336bar ( .A1(in_13bar), .A2(inbar[87]), .ZN(n634bar) );
  OR2_X1 U337 ( .A1(n632), .A2(n631), .ZN(n636) );
  AND2_X1 U337bar ( .A1(n632bar), .A2(n631bar), .ZN(n636bar) );
  OR2_X1 U338 ( .A1(in_72), .A2(in_70), .ZN(n631) );
  AND2_X1 U338bar ( .A1(in_72bar), .A2(in_70bar), .ZN(n631bar) );
  OR2_X1 U339 ( .A1(in_80), .A2(in_74), .ZN(n632) );
  AND2_X1 U339bar ( .A1(in_80bar), .A2(in_74bar), .ZN(n632bar) );
  OR2_X1 U340 ( .A1(n630), .A2(n629), .ZN(n942) );
  AND2_X1 U340bar ( .A1(n630bar), .A2(n629bar), .ZN(n942bar) );
  OR2_X1 U341 ( .A1(n628), .A2(n627), .ZN(n629) );
  AND2_X1 U341bar ( .A1(n628bar), .A2(n627bar), .ZN(n629bar) );
  OR2_X1 U342 ( .A1(n626), .A2(n625), .ZN(n627) );
  AND2_X1 U342bar ( .A1(n626bar), .A2(n625bar), .ZN(n627bar) );
  OR2_X1 U343 ( .A1(in[146]), .A2(in[100]), .ZN(n625) );
  AND2_X1 U343bar ( .A1(inbar[146]), .A2(inbar[100]), .ZN(n625bar) );
  OR2_X1 U344 ( .A1(in[168]), .A2(in[152]), .ZN(n626) );
  AND2_X1 U344bar ( .A1(inbar[168]), .A2(inbar[152]), .ZN(n626bar) );
  OR2_X1 U345 ( .A1(n624), .A2(n623), .ZN(n628) );
  AND2_X1 U345bar ( .A1(n624bar), .A2(n623bar), .ZN(n628bar) );
  OR2_X1 U346 ( .A1(in[199]), .A2(in[182]), .ZN(n623) );
  AND2_X1 U346bar ( .A1(inbar[199]), .A2(inbar[182]), .ZN(n623bar) );
  OR2_X1 U347 ( .A1(in[236]), .A2(in[204]), .ZN(n624) );
  AND2_X1 U347bar ( .A1(inbar[236]), .A2(inbar[204]), .ZN(n624bar) );
  OR2_X1 U348 ( .A1(n622), .A2(n621), .ZN(n630) );
  AND2_X1 U348bar ( .A1(n622bar), .A2(n621bar), .ZN(n630bar) );
  OR2_X1 U349 ( .A1(n620), .A2(n619), .ZN(n621) );
  AND2_X1 U349bar ( .A1(n620bar), .A2(n619bar), .ZN(n621bar) );
  OR2_X1 U350 ( .A1(in[89]), .A2(in[246]), .ZN(n619) );
  AND2_X1 U350bar ( .A1(inbar[89]), .A2(inbar[246]), .ZN(n619bar) );
  OR2_X1 U351 ( .A1(in[95]), .A2(in[92]), .ZN(n620) );
  AND2_X1 U351bar ( .A1(inbar[95]), .A2(inbar[92]), .ZN(n620bar) );
  OR2_X1 U352 ( .A1(n618), .A2(n617), .ZN(n622) );
  AND2_X1 U352bar ( .A1(n618bar), .A2(n617bar), .ZN(n622bar) );
  OR2_X1 U353 ( .A1(in_22), .A2(in_16), .ZN(n617) );
  AND2_X1 U353bar ( .A1(in_22bar), .A2(in_16bar), .ZN(n617bar) );
  OR2_X1 U354 ( .A1(in_51), .A2(in_49), .ZN(n618) );
  AND2_X1 U354bar ( .A1(in_51bar), .A2(in_49bar), .ZN(n618bar) );
  OR2_X1 U355 ( .A1(n616), .A2(n615), .ZN(n722) );
  AND2_X1 U355bar ( .A1(n616bar), .A2(n615bar), .ZN(n722bar) );
  OR2_X1 U356 ( .A1(in[158]), .A2(in[115]), .ZN(n615) );
  AND2_X1 U356bar ( .A1(inbar[158]), .A2(inbar[115]), .ZN(n615bar) );
  OR2_X1 U357 ( .A1(in[163]), .A2(n614), .ZN(n616) );
  AND2_X1 U357bar ( .A1(inbar[163]), .A2(n614bar), .ZN(n616bar) );
  OR2_X1 U358 ( .A1(in[206]), .A2(in[165]), .ZN(n614) );
  AND2_X1 U358bar ( .A1(inbar[206]), .A2(inbar[165]), .ZN(n614bar) );
  OR2_X1 U359 ( .A1(n613), .A2(n612), .ZN(n724) );
  AND2_X1 U359bar ( .A1(n613bar), .A2(n612bar), .ZN(n724bar) );
  OR2_X1 U360 ( .A1(n611), .A2(n610), .ZN(n612) );
  AND2_X1 U360bar ( .A1(n611bar), .A2(n610bar), .ZN(n612bar) );
  OR2_X1 U361 ( .A1(in[213]), .A2(in[207]), .ZN(n610) );
  AND2_X1 U361bar ( .A1(inbar[213]), .A2(inbar[207]), .ZN(n610bar) );
  OR2_X1 U362 ( .A1(in[215]), .A2(n609), .ZN(n611) );
  AND2_X1 U362bar ( .A1(inbar[215]), .A2(n609bar), .ZN(n611bar) );
  OR2_X1 U363 ( .A1(in[230]), .A2(in[220]), .ZN(n609) );
  AND2_X1 U363bar ( .A1(inbar[230]), .A2(inbar[220]), .ZN(n609bar) );
  OR2_X1 U364 ( .A1(n608), .A2(n607), .ZN(n613) );
  AND2_X1 U364bar ( .A1(n608bar), .A2(n607bar), .ZN(n613bar) );
  OR2_X1 U365 ( .A1(in[251]), .A2(in[234]), .ZN(n607) );
  AND2_X1 U365bar ( .A1(inbar[251]), .A2(inbar[234]), .ZN(n607bar) );
  OR2_X1 U366 ( .A1(in_17), .A2(n606), .ZN(n608) );
  AND2_X1 U366bar ( .A1(in_17bar), .A2(n606bar), .ZN(n608bar) );
  OR2_X1 U367 ( .A1(in_65), .A2(in_56), .ZN(n606) );
  AND2_X1 U367bar ( .A1(in_65bar), .A2(in_56bar), .ZN(n606bar) );
  OR2_X1 U368 ( .A1(n605), .A2(n604), .ZN(out[0]) );
  AND2_X1 U368bar ( .A1(n605bar), .A2(n604bar), .ZN(outbar[0]) );
  OR2_X1 U369 ( .A1(n603), .A2(n602), .ZN(n604) );
  AND2_X1 U369bar ( .A1(n603bar), .A2(n602bar), .ZN(n604bar) );
  OR2_X1 U370 ( .A1(n601), .A2(n600), .ZN(n602) );
  AND2_X1 U370bar ( .A1(n601bar), .A2(n600bar), .ZN(n602bar) );
  OR2_X1 U371 ( .A1(n820), .A2(n785), .ZN(n600) );
  AND2_X1 U371bar ( .A1(n820bar), .A2(n785bar), .ZN(n600bar) );
  OR2_X1 U372 ( .A1(n599), .A2(n598), .ZN(n785) );
  AND2_X1 U372bar ( .A1(n599bar), .A2(n598bar), .ZN(n785bar) );
  OR2_X1 U373 ( .A1(n597), .A2(n596), .ZN(n598) );
  AND2_X1 U373bar ( .A1(n597bar), .A2(n596bar), .ZN(n598bar) );
  OR2_X1 U374 ( .A1(n595), .A2(n594), .ZN(n596) );
  AND2_X1 U374bar ( .A1(n595bar), .A2(n594bar), .ZN(n596bar) );
  OR2_X1 U375 ( .A1(in[135]), .A2(in[104]), .ZN(n594) );
  AND2_X1 U375bar ( .A1(inbar[135]), .A2(inbar[104]), .ZN(n594bar) );
  OR2_X1 U376 ( .A1(in[188]), .A2(in[178]), .ZN(n595) );
  AND2_X1 U376bar ( .A1(inbar[188]), .A2(inbar[178]), .ZN(n595bar) );
  OR2_X1 U377 ( .A1(n593), .A2(n592), .ZN(n597) );
  AND2_X1 U377bar ( .A1(n593bar), .A2(n592bar), .ZN(n597bar) );
  OR2_X1 U378 ( .A1(in[217]), .A2(in[194]), .ZN(n592) );
  AND2_X1 U378bar ( .A1(inbar[217]), .A2(inbar[194]), .ZN(n592bar) );
  OR2_X1 U379 ( .A1(in[237]), .A2(in[218]), .ZN(n593) );
  AND2_X1 U379bar ( .A1(inbar[237]), .A2(inbar[218]), .ZN(n593bar) );
  OR2_X1 U380 ( .A1(n591), .A2(n590), .ZN(n599) );
  AND2_X1 U380bar ( .A1(n591bar), .A2(n590bar), .ZN(n599bar) );
  OR2_X1 U381 ( .A1(n589), .A2(n588), .ZN(n590) );
  AND2_X1 U381bar ( .A1(n589bar), .A2(n588bar), .ZN(n590bar) );
  OR2_X1 U382 ( .A1(in_2), .A2(in_10), .ZN(n588) );
  AND2_X1 U382bar ( .A1(in_2bar), .A2(in_10bar), .ZN(n588bar) );
  OR2_X1 U383 ( .A1(in_47), .A2(in_22), .ZN(n589) );
  AND2_X1 U383bar ( .A1(in_47bar), .A2(in_22bar), .ZN(n589bar) );
  OR2_X1 U384 ( .A1(n587), .A2(n586), .ZN(n591) );
  AND2_X1 U384bar ( .A1(n587bar), .A2(n586bar), .ZN(n591bar) );
  OR2_X1 U385 ( .A1(in_56), .A2(in_54), .ZN(n586) );
  AND2_X1 U385bar ( .A1(in_56bar), .A2(in_54bar), .ZN(n586bar) );
  OR2_X1 U386 ( .A1(in_63), .A2(in_61), .ZN(n587) );
  AND2_X1 U386bar ( .A1(in_63bar), .A2(in_61bar), .ZN(n587bar) );
  OR2_X1 U387 ( .A1(n585), .A2(n584), .ZN(n820) );
  AND2_X1 U387bar ( .A1(n585bar), .A2(n584bar), .ZN(n820bar) );
  OR2_X1 U388 ( .A1(n583), .A2(n582), .ZN(n584) );
  AND2_X1 U388bar ( .A1(n583bar), .A2(n582bar), .ZN(n584bar) );
  OR2_X1 U389 ( .A1(n581), .A2(n580), .ZN(n582) );
  AND2_X1 U389bar ( .A1(n581bar), .A2(n580bar), .ZN(n582bar) );
  OR2_X1 U390 ( .A1(in[158]), .A2(in[142]), .ZN(n580) );
  AND2_X1 U390bar ( .A1(inbar[158]), .A2(inbar[142]), .ZN(n580bar) );
  OR2_X1 U391 ( .A1(in[175]), .A2(in[164]), .ZN(n581) );
  AND2_X1 U391bar ( .A1(inbar[175]), .A2(inbar[164]), .ZN(n581bar) );
  OR2_X1 U392 ( .A1(n579), .A2(n578), .ZN(n583) );
  AND2_X1 U392bar ( .A1(n579bar), .A2(n578bar), .ZN(n583bar) );
  OR2_X1 U393 ( .A1(in[228]), .A2(in[204]), .ZN(n578) );
  AND2_X1 U393bar ( .A1(inbar[228]), .A2(inbar[204]), .ZN(n578bar) );
  OR2_X1 U394 ( .A1(in[91]), .A2(in[87]), .ZN(n579) );
  AND2_X1 U394bar ( .A1(inbar[91]), .A2(inbar[87]), .ZN(n579bar) );
  OR2_X1 U395 ( .A1(n577), .A2(n576), .ZN(n585) );
  AND2_X1 U395bar ( .A1(n577bar), .A2(n576bar), .ZN(n585bar) );
  OR2_X1 U396 ( .A1(n575), .A2(n574), .ZN(n576) );
  AND2_X1 U396bar ( .A1(n575bar), .A2(n574bar), .ZN(n576bar) );
  OR2_X1 U397 ( .A1(in_21), .A2(in_11), .ZN(n574) );
  AND2_X1 U397bar ( .A1(in_21bar), .A2(in_11bar), .ZN(n574bar) );
  OR2_X1 U398 ( .A1(in_5), .A2(in_3), .ZN(n575) );
  AND2_X1 U398bar ( .A1(in_5bar), .A2(in_3bar), .ZN(n575bar) );
  OR2_X1 U399 ( .A1(n573), .A2(n572), .ZN(n577) );
  AND2_X1 U399bar ( .A1(n573bar), .A2(n572bar), .ZN(n577bar) );
  OR2_X1 U400 ( .A1(in_68), .A2(in_64), .ZN(n572) );
  AND2_X1 U400bar ( .A1(in_68bar), .A2(in_64bar), .ZN(n572bar) );
  OR2_X1 U401 ( .A1(in_76), .A2(in_73), .ZN(n573) );
  AND2_X1 U401bar ( .A1(in_76bar), .A2(in_73bar), .ZN(n573bar) );
  OR2_X1 U402 ( .A1(n778), .A2(n571), .ZN(n601) );
  AND2_X1 U402bar ( .A1(n778bar), .A2(n571bar), .ZN(n601bar) );
  OR2_X1 U403 ( .A1(in[100]), .A2(n965), .ZN(n571) );
  AND2_X1 U403bar ( .A1(inbar[100]), .A2(n965bar), .ZN(n571bar) );
  OR2_X1 U404 ( .A1(n570), .A2(n569), .ZN(n965) );
  AND2_X1 U404bar ( .A1(n570bar), .A2(n569bar), .ZN(n965bar) );
  OR2_X1 U405 ( .A1(n568), .A2(n567), .ZN(n569) );
  AND2_X1 U405bar ( .A1(n568bar), .A2(n567bar), .ZN(n569bar) );
  OR2_X1 U406 ( .A1(n566), .A2(n565), .ZN(n567) );
  AND2_X1 U406bar ( .A1(n566bar), .A2(n565bar), .ZN(n567bar) );
  OR2_X1 U407 ( .A1(n817), .A2(n750), .ZN(n565) );
  AND2_X1 U407bar ( .A1(n817bar), .A2(n750bar), .ZN(n565bar) );
  OR2_X1 U408 ( .A1(n564), .A2(n563), .ZN(n750) );
  AND2_X1 U408bar ( .A1(n564bar), .A2(n563bar), .ZN(n750bar) );
  OR2_X1 U409 ( .A1(n562), .A2(n561), .ZN(n563) );
  AND2_X1 U409bar ( .A1(n562bar), .A2(n561bar), .ZN(n563bar) );
  OR2_X1 U410 ( .A1(n560), .A2(n559), .ZN(n561) );
  AND2_X1 U410bar ( .A1(n560bar), .A2(n559bar), .ZN(n561bar) );
  OR2_X1 U411 ( .A1(in[119]), .A2(in[103]), .ZN(n559) );
  AND2_X1 U411bar ( .A1(inbar[119]), .A2(inbar[103]), .ZN(n559bar) );
  OR2_X1 U412 ( .A1(in[137]), .A2(in[133]), .ZN(n560) );
  AND2_X1 U412bar ( .A1(inbar[137]), .A2(inbar[133]), .ZN(n560bar) );
  OR2_X1 U413 ( .A1(n558), .A2(n557), .ZN(n562) );
  AND2_X1 U413bar ( .A1(n558bar), .A2(n557bar), .ZN(n562bar) );
  OR2_X1 U414 ( .A1(in[176]), .A2(in[173]), .ZN(n557) );
  AND2_X1 U414bar ( .A1(inbar[176]), .A2(inbar[173]), .ZN(n557bar) );
  OR2_X1 U415 ( .A1(in[210]), .A2(in[181]), .ZN(n558) );
  AND2_X1 U415bar ( .A1(inbar[210]), .A2(inbar[181]), .ZN(n558bar) );
  OR2_X1 U416 ( .A1(n556), .A2(n555), .ZN(n564) );
  AND2_X1 U416bar ( .A1(n556bar), .A2(n555bar), .ZN(n564bar) );
  OR2_X1 U417 ( .A1(n554), .A2(n553), .ZN(n555) );
  AND2_X1 U417bar ( .A1(n554bar), .A2(n553bar), .ZN(n555bar) );
  OR2_X1 U418 ( .A1(in_13), .A2(in[234]), .ZN(n553) );
  AND2_X1 U418bar ( .A1(in_13bar), .A2(inbar[234]), .ZN(n553bar) );
  OR2_X1 U419 ( .A1(in_38), .A2(in_32), .ZN(n554) );
  AND2_X1 U419bar ( .A1(in_38bar), .A2(in_32bar), .ZN(n554bar) );
  OR2_X1 U420 ( .A1(n552), .A2(n551), .ZN(n556) );
  AND2_X1 U420bar ( .A1(n552bar), .A2(n551bar), .ZN(n556bar) );
  OR2_X1 U421 ( .A1(in_42), .A2(in_41), .ZN(n551) );
  AND2_X1 U421bar ( .A1(in_42bar), .A2(in_41bar), .ZN(n551bar) );
  OR2_X1 U422 ( .A1(in_7), .A2(in_49), .ZN(n552) );
  AND2_X1 U422bar ( .A1(in_7bar), .A2(in_49bar), .ZN(n552bar) );
  OR2_X1 U423 ( .A1(n550), .A2(n549), .ZN(n817) );
  AND2_X1 U423bar ( .A1(n550bar), .A2(n549bar), .ZN(n817bar) );
  OR2_X1 U424 ( .A1(n548), .A2(n547), .ZN(n549) );
  AND2_X1 U424bar ( .A1(n548bar), .A2(n547bar), .ZN(n549bar) );
  OR2_X1 U425 ( .A1(n546), .A2(n545), .ZN(n547) );
  AND2_X1 U425bar ( .A1(n546bar), .A2(n545bar), .ZN(n547bar) );
  OR2_X1 U426 ( .A1(in[159]), .A2(in[105]), .ZN(n545) );
  AND2_X1 U426bar ( .A1(inbar[159]), .A2(inbar[105]), .ZN(n545bar) );
  OR2_X1 U427 ( .A1(in[206]), .A2(in[183]), .ZN(n546) );
  AND2_X1 U427bar ( .A1(inbar[206]), .A2(inbar[183]), .ZN(n546bar) );
  OR2_X1 U428 ( .A1(n544), .A2(n543), .ZN(n548) );
  AND2_X1 U428bar ( .A1(n544bar), .A2(n543bar), .ZN(n548bar) );
  OR2_X1 U429 ( .A1(in[229]), .A2(in[219]), .ZN(n543) );
  AND2_X1 U429bar ( .A1(inbar[229]), .A2(inbar[219]), .ZN(n543bar) );
  OR2_X1 U430 ( .A1(in[235]), .A2(in[232]), .ZN(n544) );
  AND2_X1 U430bar ( .A1(inbar[235]), .A2(inbar[232]), .ZN(n544bar) );
  OR2_X1 U431 ( .A1(n542), .A2(n541), .ZN(n550) );
  AND2_X1 U431bar ( .A1(n542bar), .A2(n541bar), .ZN(n550bar) );
  OR2_X1 U432 ( .A1(n540), .A2(n539), .ZN(n541) );
  AND2_X1 U432bar ( .A1(n540bar), .A2(n539bar), .ZN(n541bar) );
  OR2_X1 U433 ( .A1(in[249]), .A2(in[242]), .ZN(n539) );
  AND2_X1 U433bar ( .A1(inbar[249]), .A2(inbar[242]), .ZN(n539bar) );
  OR2_X1 U434 ( .A1(in[89]), .A2(in[254]), .ZN(n540) );
  AND2_X1 U434bar ( .A1(inbar[89]), .A2(inbar[254]), .ZN(n540bar) );
  OR2_X1 U435 ( .A1(n538), .A2(n537), .ZN(n542) );
  AND2_X1 U435bar ( .A1(n538bar), .A2(n537bar), .ZN(n542bar) );
  OR2_X1 U436 ( .A1(in_14), .A2(in[99]), .ZN(n537) );
  AND2_X1 U436bar ( .A1(in_14bar), .A2(inbar[99]), .ZN(n537bar) );
  OR2_X1 U437 ( .A1(in_60), .A2(in_18), .ZN(n538) );
  AND2_X1 U437bar ( .A1(in_60bar), .A2(in_18bar), .ZN(n538bar) );
  OR2_X1 U438 ( .A1(in[113]), .A2(n763), .ZN(n566) );
  AND2_X1 U438bar ( .A1(inbar[113]), .A2(n763bar), .ZN(n566bar) );
  OR2_X1 U439 ( .A1(n536), .A2(n535), .ZN(n763) );
  AND2_X1 U439bar ( .A1(n536bar), .A2(n535bar), .ZN(n763bar) );
  OR2_X1 U440 ( .A1(n534), .A2(n533), .ZN(n535) );
  AND2_X1 U440bar ( .A1(n534bar), .A2(n533bar), .ZN(n535bar) );
  OR2_X1 U441 ( .A1(n532), .A2(n531), .ZN(n533) );
  AND2_X1 U441bar ( .A1(n532bar), .A2(n531bar), .ZN(n533bar) );
  OR2_X1 U442 ( .A1(in[115]), .A2(in[110]), .ZN(n531) );
  AND2_X1 U442bar ( .A1(inbar[115]), .A2(inbar[110]), .ZN(n531bar) );
  OR2_X1 U443 ( .A1(in[125]), .A2(in[117]), .ZN(n532) );
  AND2_X1 U443bar ( .A1(inbar[125]), .A2(inbar[117]), .ZN(n532bar) );
  OR2_X1 U444 ( .A1(n530), .A2(n529), .ZN(n534) );
  AND2_X1 U444bar ( .A1(n530bar), .A2(n529bar), .ZN(n534bar) );
  OR2_X1 U445 ( .A1(in[180]), .A2(in[128]), .ZN(n529) );
  AND2_X1 U445bar ( .A1(inbar[180]), .A2(inbar[128]), .ZN(n529bar) );
  OR2_X1 U446 ( .A1(in[205]), .A2(in[201]), .ZN(n530) );
  AND2_X1 U446bar ( .A1(inbar[205]), .A2(inbar[201]), .ZN(n530bar) );
  OR2_X1 U447 ( .A1(n528), .A2(n527), .ZN(n536) );
  AND2_X1 U447bar ( .A1(n528bar), .A2(n527bar), .ZN(n536bar) );
  OR2_X1 U448 ( .A1(n526), .A2(n525), .ZN(n527) );
  AND2_X1 U448bar ( .A1(n526bar), .A2(n525bar), .ZN(n527bar) );
  OR2_X1 U449 ( .A1(in[244]), .A2(in[239]), .ZN(n525) );
  AND2_X1 U449bar ( .A1(inbar[244]), .A2(inbar[239]), .ZN(n525bar) );
  OR2_X1 U450 ( .A1(in[95]), .A2(in[83]), .ZN(n526) );
  AND2_X1 U450bar ( .A1(inbar[95]), .A2(inbar[83]), .ZN(n526bar) );
  OR2_X1 U451 ( .A1(n524), .A2(n523), .ZN(n528) );
  AND2_X1 U451bar ( .A1(n524bar), .A2(n523bar), .ZN(n528bar) );
  OR2_X1 U452 ( .A1(in_24), .A2(in[97]), .ZN(n523) );
  AND2_X1 U452bar ( .A1(in_24bar), .A2(inbar[97]), .ZN(n523bar) );
  OR2_X1 U453 ( .A1(in_33), .A2(in_27), .ZN(n524) );
  AND2_X1 U453bar ( .A1(in_33bar), .A2(in_27bar), .ZN(n524bar) );
  OR2_X1 U454 ( .A1(n522), .A2(n521), .ZN(n568) );
  AND2_X1 U454bar ( .A1(n522bar), .A2(n521bar), .ZN(n568bar) );
  OR2_X1 U455 ( .A1(in[145]), .A2(in[126]), .ZN(n521) );
  AND2_X1 U455bar ( .A1(inbar[145]), .A2(inbar[126]), .ZN(n521bar) );
  OR2_X1 U456 ( .A1(in[169]), .A2(n520), .ZN(n522) );
  AND2_X1 U456bar ( .A1(inbar[169]), .A2(n520bar), .ZN(n522bar) );
  OR2_X1 U457 ( .A1(in[221]), .A2(in[172]), .ZN(n520) );
  AND2_X1 U457bar ( .A1(inbar[221]), .A2(inbar[172]), .ZN(n520bar) );
  OR2_X1 U458 ( .A1(n519), .A2(n518), .ZN(n570) );
  AND2_X1 U458bar ( .A1(n519bar), .A2(n518bar), .ZN(n570bar) );
  OR2_X1 U459 ( .A1(n517), .A2(n516), .ZN(n518) );
  AND2_X1 U459bar ( .A1(n517bar), .A2(n516bar), .ZN(n518bar) );
  OR2_X1 U460 ( .A1(in[241]), .A2(in[224]), .ZN(n516) );
  AND2_X1 U460bar ( .A1(inbar[241]), .A2(inbar[224]), .ZN(n516bar) );
  OR2_X1 U461 ( .A1(in[86]), .A2(n515), .ZN(n517) );
  AND2_X1 U461bar ( .A1(inbar[86]), .A2(n515bar), .ZN(n517bar) );
  OR2_X1 U462 ( .A1(in_43), .A2(in_34), .ZN(n515) );
  AND2_X1 U462bar ( .A1(in_43bar), .A2(in_34bar), .ZN(n515bar) );
  OR2_X1 U463 ( .A1(n514), .A2(n513), .ZN(n519) );
  AND2_X1 U463bar ( .A1(n514bar), .A2(n513bar), .ZN(n519bar) );
  OR2_X1 U464 ( .A1(in_65), .A2(in_51), .ZN(n513) );
  AND2_X1 U464bar ( .A1(in_65bar), .A2(in_51bar), .ZN(n513bar) );
  OR2_X1 U465 ( .A1(in_75), .A2(n512), .ZN(n514) );
  AND2_X1 U465bar ( .A1(in_75bar), .A2(n512bar), .ZN(n514bar) );
  OR2_X1 U466 ( .A1(in_81), .A2(in_77), .ZN(n512) );
  AND2_X1 U466bar ( .A1(in_81bar), .A2(in_77bar), .ZN(n512bar) );
  OR2_X1 U467 ( .A1(n511), .A2(n510), .ZN(n778) );
  AND2_X1 U467bar ( .A1(n511bar), .A2(n510bar), .ZN(n778bar) );
  OR2_X1 U468 ( .A1(n509), .A2(n508), .ZN(n510) );
  AND2_X1 U468bar ( .A1(n509bar), .A2(n508bar), .ZN(n510bar) );
  OR2_X1 U469 ( .A1(n507), .A2(n506), .ZN(n508) );
  AND2_X1 U469bar ( .A1(n507bar), .A2(n506bar), .ZN(n508bar) );
  OR2_X1 U470 ( .A1(in[107]), .A2(in[101]), .ZN(n506) );
  AND2_X1 U470bar ( .A1(inbar[107]), .A2(inbar[101]), .ZN(n506bar) );
  OR2_X1 U471 ( .A1(in[139]), .A2(in[132]), .ZN(n507) );
  AND2_X1 U471bar ( .A1(inbar[139]), .A2(inbar[132]), .ZN(n507bar) );
  OR2_X1 U472 ( .A1(n505), .A2(n504), .ZN(n509) );
  AND2_X1 U472bar ( .A1(n505bar), .A2(n504bar), .ZN(n509bar) );
  OR2_X1 U473 ( .A1(in[146]), .A2(in[141]), .ZN(n504) );
  AND2_X1 U473bar ( .A1(inbar[146]), .A2(inbar[141]), .ZN(n504bar) );
  OR2_X1 U474 ( .A1(in[203]), .A2(in[179]), .ZN(n505) );
  AND2_X1 U474bar ( .A1(inbar[203]), .A2(inbar[179]), .ZN(n505bar) );
  OR2_X1 U475 ( .A1(n503), .A2(n502), .ZN(n511) );
  AND2_X1 U475bar ( .A1(n503bar), .A2(n502bar), .ZN(n511bar) );
  OR2_X1 U476 ( .A1(n501), .A2(n500), .ZN(n502) );
  AND2_X1 U476bar ( .A1(n501bar), .A2(n500bar), .ZN(n502bar) );
  OR2_X1 U477 ( .A1(in[243]), .A2(in[222]), .ZN(n500) );
  AND2_X1 U477bar ( .A1(inbar[243]), .A2(inbar[222]), .ZN(n500bar) );
  OR2_X1 U478 ( .A1(in[251]), .A2(in[250]), .ZN(n501) );
  AND2_X1 U478bar ( .A1(inbar[251]), .A2(inbar[250]), .ZN(n501bar) );
  OR2_X1 U479 ( .A1(n499), .A2(n498), .ZN(n503) );
  AND2_X1 U479bar ( .A1(n499bar), .A2(n498bar), .ZN(n503bar) );
  OR2_X1 U480 ( .A1(in_37), .A2(in_19), .ZN(n498) );
  AND2_X1 U480bar ( .A1(in_37bar), .A2(in_19bar), .ZN(n498bar) );
  OR2_X1 U481 ( .A1(in_78), .A2(in_6), .ZN(n499) );
  AND2_X1 U481bar ( .A1(in_78bar), .A2(in_6bar), .ZN(n499bar) );
  OR2_X1 U482 ( .A1(n497), .A2(n496), .ZN(n603) );
  AND2_X1 U482bar ( .A1(n497bar), .A2(n496bar), .ZN(n603bar) );
  OR2_X1 U483 ( .A1(in[112]), .A2(in[102]), .ZN(n496) );
  AND2_X1 U483bar ( .A1(inbar[112]), .A2(inbar[102]), .ZN(n496bar) );
  OR2_X1 U484 ( .A1(in[123]), .A2(n495), .ZN(n497) );
  AND2_X1 U484bar ( .A1(inbar[123]), .A2(n495bar), .ZN(n497bar) );
  OR2_X1 U485 ( .A1(in[143]), .A2(in[130]), .ZN(n495) );
  AND2_X1 U485bar ( .A1(inbar[143]), .A2(inbar[130]), .ZN(n495bar) );
  OR2_X1 U486 ( .A1(n494), .A2(n493), .ZN(n605) );
  AND2_X1 U486bar ( .A1(n494bar), .A2(n493bar), .ZN(n605bar) );
  OR2_X1 U487 ( .A1(n492), .A2(n491), .ZN(n493) );
  AND2_X1 U487bar ( .A1(n492bar), .A2(n491bar), .ZN(n493bar) );
  OR2_X1 U488 ( .A1(in[216]), .A2(in[213]), .ZN(n491) );
  AND2_X1 U488bar ( .A1(inbar[216]), .A2(inbar[213]), .ZN(n491bar) );
  OR2_X1 U489 ( .A1(in[227]), .A2(n490), .ZN(n492) );
  AND2_X1 U489bar ( .A1(inbar[227]), .A2(n490bar), .ZN(n492bar) );
  OR2_X1 U490 ( .A1(in_0), .A2(in[248]), .ZN(n490) );
  AND2_X1 U490bar ( .A1(in_0bar), .A2(inbar[248]), .ZN(n490bar) );
  OR2_X1 U491 ( .A1(n489), .A2(n488), .ZN(n494) );
  AND2_X1 U491bar ( .A1(n489bar), .A2(n488bar), .ZN(n494bar) );
  OR2_X1 U492 ( .A1(in_46), .A2(in_44), .ZN(n488) );
  AND2_X1 U492bar ( .A1(in_46bar), .A2(in_44bar), .ZN(n488bar) );
  OR2_X1 U493 ( .A1(in_50), .A2(n487), .ZN(n489) );
  AND2_X1 U493bar ( .A1(in_50bar), .A2(n487bar), .ZN(n489bar) );
  OR2_X1 U494 ( .A1(in_9), .A2(in_80), .ZN(n487) );
  AND2_X1 U494bar ( .A1(in_9bar), .A2(in_80bar), .ZN(n487bar) );
endmodule

module sBox_9 ( in, inbar, out, outbar );

  input wire [7:0] in;
  input wire [7:0] inbar;
//input_done

  output wire [7:0] out;
  output wire [7:0] outbar;
//output_done

  wire [255:0] decodeOut;
  wire [255:0] decodeOutbar;
//wire_done

  decode_9 dec ( .in(in), .inbar(inbar), .out(decodeOut), .outbar(decodeOutbar) );
  encode_9 enc ( .in(decodeOut), .inbar(decodeOutbar), .out(out), .outbar(outbar) );
endmodule

module CD2_37 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD2_38 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD2_39 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD2_40 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD4_19 ( a, abar, b, bbar, y, ybar );

  input wire [3:0] a;
  input wire [3:0] b;
  input wire [3:0] abar;
  input wire [3:0] bbar;
//input_done

  output wire [15:0] y;
  output wire [15:0] ybar;
//output_done

//wire_done

  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]) );
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]) );
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]) );
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]) );
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]) );
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]) );
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]) );
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]) );
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]) );
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]) );
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]) );
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]) );
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]) );
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]) );
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]) );
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]) );
endmodule

module CD4_20 ( a, abar, b, bbar, y, ybar );

  input wire [3:0] a;
  input wire [3:0] b;
  input wire [3:0] abar;
  input wire [3:0] bbar;
//input_done

  output wire [15:0] y;
  output wire [15:0] ybar;
//output_done

//wire_done

  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]) );
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]) );
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]) );
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]) );
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]) );
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]) );
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]) );
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]) );
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]) );
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]) );
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]) );
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]) );
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]) );
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]) );
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]) );
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]) );
endmodule

module CD16_10 ( a, abar, b, bbar, y, ybar );

  input wire [15:0] a;
  input wire [15:0] b;
  input wire [15:0] abar;
  input wire [15:0] bbar;
//input_done

  output wire [255:0] y;
  output wire [255:0] ybar;
//output_done

//wire_done

  AND2_X1 U1 ( .A1(b[9]), .A2(a[0]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[9]), .A2(abar[0]), .ZN(ybar[9]) );
  AND2_X1 U2 ( .A1(b[3]), .A2(a[6]), .ZN(y[99]) );
  OR2_X1 U2bar ( .A1(bbar[3]), .A2(abar[6]), .ZN(ybar[99]) );
  AND2_X1 U3 ( .A1(b[2]), .A2(a[6]), .ZN(y[98]) );
  OR2_X1 U3bar ( .A1(bbar[2]), .A2(abar[6]), .ZN(ybar[98]) );
  AND2_X1 U4 ( .A1(b[1]), .A2(a[6]), .ZN(y[97]) );
  OR2_X1 U4bar ( .A1(bbar[1]), .A2(abar[6]), .ZN(ybar[97]) );
  AND2_X1 U5 ( .A1(b[0]), .A2(a[6]), .ZN(y[96]) );
  OR2_X1 U5bar ( .A1(bbar[0]), .A2(abar[6]), .ZN(ybar[96]) );
  AND2_X1 U6 ( .A1(b[15]), .A2(a[5]), .ZN(y[95]) );
  OR2_X1 U6bar ( .A1(bbar[15]), .A2(abar[5]), .ZN(ybar[95]) );
  AND2_X1 U7 ( .A1(b[14]), .A2(a[5]), .ZN(y[94]) );
  OR2_X1 U7bar ( .A1(bbar[14]), .A2(abar[5]), .ZN(ybar[94]) );
  AND2_X1 U8 ( .A1(b[13]), .A2(a[5]), .ZN(y[93]) );
  OR2_X1 U8bar ( .A1(bbar[13]), .A2(abar[5]), .ZN(ybar[93]) );
  AND2_X1 U9 ( .A1(b[12]), .A2(a[5]), .ZN(y[92]) );
  OR2_X1 U9bar ( .A1(bbar[12]), .A2(abar[5]), .ZN(ybar[92]) );
  AND2_X1 U10 ( .A1(b[11]), .A2(a[5]), .ZN(y[91]) );
  OR2_X1 U10bar ( .A1(bbar[11]), .A2(abar[5]), .ZN(ybar[91]) );
  AND2_X1 U11 ( .A1(b[10]), .A2(a[5]), .ZN(y[90]) );
  OR2_X1 U11bar ( .A1(bbar[10]), .A2(abar[5]), .ZN(ybar[90]) );
  AND2_X1 U12 ( .A1(b[8]), .A2(a[0]), .ZN(y[8]) );
  OR2_X1 U12bar ( .A1(bbar[8]), .A2(abar[0]), .ZN(ybar[8]) );
  AND2_X1 U13 ( .A1(a[5]), .A2(b[9]), .ZN(y[89]) );
  OR2_X1 U13bar ( .A1(abar[5]), .A2(bbar[9]), .ZN(ybar[89]) );
  AND2_X1 U14 ( .A1(b[8]), .A2(a[5]), .ZN(y[88]) );
  OR2_X1 U14bar ( .A1(bbar[8]), .A2(abar[5]), .ZN(ybar[88]) );
  AND2_X1 U15 ( .A1(b[7]), .A2(a[5]), .ZN(y[87]) );
  OR2_X1 U15bar ( .A1(bbar[7]), .A2(abar[5]), .ZN(ybar[87]) );
  AND2_X1 U16 ( .A1(b[6]), .A2(a[5]), .ZN(y[86]) );
  OR2_X1 U16bar ( .A1(bbar[6]), .A2(abar[5]), .ZN(ybar[86]) );
  AND2_X1 U17 ( .A1(b[5]), .A2(a[5]), .ZN(y[85]) );
  OR2_X1 U17bar ( .A1(bbar[5]), .A2(abar[5]), .ZN(ybar[85]) );
  AND2_X1 U18 ( .A1(b[4]), .A2(a[5]), .ZN(y[84]) );
  OR2_X1 U18bar ( .A1(bbar[4]), .A2(abar[5]), .ZN(ybar[84]) );
  AND2_X1 U19 ( .A1(a[5]), .A2(b[3]), .ZN(y[83]) );
  OR2_X1 U19bar ( .A1(abar[5]), .A2(bbar[3]), .ZN(ybar[83]) );
  AND2_X1 U20 ( .A1(a[5]), .A2(b[2]), .ZN(y[82]) );
  OR2_X1 U20bar ( .A1(abar[5]), .A2(bbar[2]), .ZN(ybar[82]) );
  AND2_X1 U21 ( .A1(a[5]), .A2(b[1]), .ZN(y[81]) );
  OR2_X1 U21bar ( .A1(abar[5]), .A2(bbar[1]), .ZN(ybar[81]) );
  AND2_X1 U22 ( .A1(a[5]), .A2(b[0]), .ZN(y[80]) );
  OR2_X1 U22bar ( .A1(abar[5]), .A2(bbar[0]), .ZN(ybar[80]) );
  AND2_X1 U23 ( .A1(b[7]), .A2(a[0]), .ZN(y[7]) );
  OR2_X1 U23bar ( .A1(bbar[7]), .A2(abar[0]), .ZN(ybar[7]) );
  AND2_X1 U24 ( .A1(a[4]), .A2(b[15]), .ZN(y[79]) );
  OR2_X1 U24bar ( .A1(abar[4]), .A2(bbar[15]), .ZN(ybar[79]) );
  AND2_X1 U25 ( .A1(a[4]), .A2(b[14]), .ZN(y[78]) );
  OR2_X1 U25bar ( .A1(abar[4]), .A2(bbar[14]), .ZN(ybar[78]) );
  AND2_X1 U26 ( .A1(a[4]), .A2(b[13]), .ZN(y[77]) );
  OR2_X1 U26bar ( .A1(abar[4]), .A2(bbar[13]), .ZN(ybar[77]) );
  AND2_X1 U27 ( .A1(a[4]), .A2(b[12]), .ZN(y[76]) );
  OR2_X1 U27bar ( .A1(abar[4]), .A2(bbar[12]), .ZN(ybar[76]) );
  AND2_X1 U28 ( .A1(a[4]), .A2(b[11]), .ZN(y[75]) );
  OR2_X1 U28bar ( .A1(abar[4]), .A2(bbar[11]), .ZN(ybar[75]) );
  AND2_X1 U29 ( .A1(a[4]), .A2(b[10]), .ZN(y[74]) );
  OR2_X1 U29bar ( .A1(abar[4]), .A2(bbar[10]), .ZN(ybar[74]) );
  AND2_X1 U30 ( .A1(a[4]), .A2(b[9]), .ZN(y[73]) );
  OR2_X1 U30bar ( .A1(abar[4]), .A2(bbar[9]), .ZN(ybar[73]) );
  AND2_X1 U31 ( .A1(a[4]), .A2(b[8]), .ZN(y[72]) );
  OR2_X1 U31bar ( .A1(abar[4]), .A2(bbar[8]), .ZN(ybar[72]) );
  AND2_X1 U32 ( .A1(a[4]), .A2(b[7]), .ZN(y[71]) );
  OR2_X1 U32bar ( .A1(abar[4]), .A2(bbar[7]), .ZN(ybar[71]) );
  AND2_X1 U33 ( .A1(a[4]), .A2(b[6]), .ZN(y[70]) );
  OR2_X1 U33bar ( .A1(abar[4]), .A2(bbar[6]), .ZN(ybar[70]) );
  AND2_X1 U34 ( .A1(b[6]), .A2(a[0]), .ZN(y[6]) );
  OR2_X1 U34bar ( .A1(bbar[6]), .A2(abar[0]), .ZN(ybar[6]) );
  AND2_X1 U35 ( .A1(a[4]), .A2(b[5]), .ZN(y[69]) );
  OR2_X1 U35bar ( .A1(abar[4]), .A2(bbar[5]), .ZN(ybar[69]) );
  AND2_X1 U36 ( .A1(a[4]), .A2(b[4]), .ZN(y[68]) );
  OR2_X1 U36bar ( .A1(abar[4]), .A2(bbar[4]), .ZN(ybar[68]) );
  AND2_X1 U37 ( .A1(a[4]), .A2(b[3]), .ZN(y[67]) );
  OR2_X1 U37bar ( .A1(abar[4]), .A2(bbar[3]), .ZN(ybar[67]) );
  AND2_X1 U38 ( .A1(a[4]), .A2(b[2]), .ZN(y[66]) );
  OR2_X1 U38bar ( .A1(abar[4]), .A2(bbar[2]), .ZN(ybar[66]) );
  AND2_X1 U39 ( .A1(a[4]), .A2(b[1]), .ZN(y[65]) );
  OR2_X1 U39bar ( .A1(abar[4]), .A2(bbar[1]), .ZN(ybar[65]) );
  AND2_X1 U40 ( .A1(a[4]), .A2(b[0]), .ZN(y[64]) );
  OR2_X1 U40bar ( .A1(abar[4]), .A2(bbar[0]), .ZN(ybar[64]) );
  AND2_X1 U41 ( .A1(a[3]), .A2(b[15]), .ZN(y[63]) );
  OR2_X1 U41bar ( .A1(abar[3]), .A2(bbar[15]), .ZN(ybar[63]) );
  AND2_X1 U42 ( .A1(a[3]), .A2(b[14]), .ZN(y[62]) );
  OR2_X1 U42bar ( .A1(abar[3]), .A2(bbar[14]), .ZN(ybar[62]) );
  AND2_X1 U43 ( .A1(a[3]), .A2(b[13]), .ZN(y[61]) );
  OR2_X1 U43bar ( .A1(abar[3]), .A2(bbar[13]), .ZN(ybar[61]) );
  AND2_X1 U44 ( .A1(a[3]), .A2(b[12]), .ZN(y[60]) );
  OR2_X1 U44bar ( .A1(abar[3]), .A2(bbar[12]), .ZN(ybar[60]) );
  AND2_X1 U45 ( .A1(b[5]), .A2(a[0]), .ZN(y[5]) );
  OR2_X1 U45bar ( .A1(bbar[5]), .A2(abar[0]), .ZN(ybar[5]) );
  AND2_X1 U46 ( .A1(a[3]), .A2(b[11]), .ZN(y[59]) );
  OR2_X1 U46bar ( .A1(abar[3]), .A2(bbar[11]), .ZN(ybar[59]) );
  AND2_X1 U47 ( .A1(a[3]), .A2(b[10]), .ZN(y[58]) );
  OR2_X1 U47bar ( .A1(abar[3]), .A2(bbar[10]), .ZN(ybar[58]) );
  AND2_X1 U48 ( .A1(a[3]), .A2(b[9]), .ZN(y[57]) );
  OR2_X1 U48bar ( .A1(abar[3]), .A2(bbar[9]), .ZN(ybar[57]) );
  AND2_X1 U49 ( .A1(a[3]), .A2(b[8]), .ZN(y[56]) );
  OR2_X1 U49bar ( .A1(abar[3]), .A2(bbar[8]), .ZN(ybar[56]) );
  AND2_X1 U50 ( .A1(a[3]), .A2(b[7]), .ZN(y[55]) );
  OR2_X1 U50bar ( .A1(abar[3]), .A2(bbar[7]), .ZN(ybar[55]) );
  AND2_X1 U51 ( .A1(a[3]), .A2(b[6]), .ZN(y[54]) );
  OR2_X1 U51bar ( .A1(abar[3]), .A2(bbar[6]), .ZN(ybar[54]) );
  AND2_X1 U52 ( .A1(a[3]), .A2(b[5]), .ZN(y[53]) );
  OR2_X1 U52bar ( .A1(abar[3]), .A2(bbar[5]), .ZN(ybar[53]) );
  AND2_X1 U53 ( .A1(a[3]), .A2(b[4]), .ZN(y[52]) );
  OR2_X1 U53bar ( .A1(abar[3]), .A2(bbar[4]), .ZN(ybar[52]) );
  AND2_X1 U54 ( .A1(a[3]), .A2(b[3]), .ZN(y[51]) );
  OR2_X1 U54bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[51]) );
  AND2_X1 U55 ( .A1(a[3]), .A2(b[2]), .ZN(y[50]) );
  OR2_X1 U55bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[50]) );
  AND2_X1 U56 ( .A1(b[4]), .A2(a[0]), .ZN(y[4]) );
  OR2_X1 U56bar ( .A1(bbar[4]), .A2(abar[0]), .ZN(ybar[4]) );
  AND2_X1 U57 ( .A1(a[3]), .A2(b[1]), .ZN(y[49]) );
  OR2_X1 U57bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[49]) );
  AND2_X1 U58 ( .A1(a[3]), .A2(b[0]), .ZN(y[48]) );
  OR2_X1 U58bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[48]) );
  AND2_X1 U59 ( .A1(a[2]), .A2(b[15]), .ZN(y[47]) );
  OR2_X1 U59bar ( .A1(abar[2]), .A2(bbar[15]), .ZN(ybar[47]) );
  AND2_X1 U60 ( .A1(a[2]), .A2(b[14]), .ZN(y[46]) );
  OR2_X1 U60bar ( .A1(abar[2]), .A2(bbar[14]), .ZN(ybar[46]) );
  AND2_X1 U61 ( .A1(a[2]), .A2(b[13]), .ZN(y[45]) );
  OR2_X1 U61bar ( .A1(abar[2]), .A2(bbar[13]), .ZN(ybar[45]) );
  AND2_X1 U62 ( .A1(a[2]), .A2(b[12]), .ZN(y[44]) );
  OR2_X1 U62bar ( .A1(abar[2]), .A2(bbar[12]), .ZN(ybar[44]) );
  AND2_X1 U63 ( .A1(a[2]), .A2(b[11]), .ZN(y[43]) );
  OR2_X1 U63bar ( .A1(abar[2]), .A2(bbar[11]), .ZN(ybar[43]) );
  AND2_X1 U64 ( .A1(a[2]), .A2(b[10]), .ZN(y[42]) );
  OR2_X1 U64bar ( .A1(abar[2]), .A2(bbar[10]), .ZN(ybar[42]) );
  AND2_X1 U65 ( .A1(a[2]), .A2(b[9]), .ZN(y[41]) );
  OR2_X1 U65bar ( .A1(abar[2]), .A2(bbar[9]), .ZN(ybar[41]) );
  AND2_X1 U66 ( .A1(a[2]), .A2(b[8]), .ZN(y[40]) );
  OR2_X1 U66bar ( .A1(abar[2]), .A2(bbar[8]), .ZN(ybar[40]) );
  AND2_X1 U67 ( .A1(b[3]), .A2(a[0]), .ZN(y[3]) );
  OR2_X1 U67bar ( .A1(bbar[3]), .A2(abar[0]), .ZN(ybar[3]) );
  AND2_X1 U68 ( .A1(a[2]), .A2(b[7]), .ZN(y[39]) );
  OR2_X1 U68bar ( .A1(abar[2]), .A2(bbar[7]), .ZN(ybar[39]) );
  AND2_X1 U69 ( .A1(a[2]), .A2(b[6]), .ZN(y[38]) );
  OR2_X1 U69bar ( .A1(abar[2]), .A2(bbar[6]), .ZN(ybar[38]) );
  AND2_X1 U70 ( .A1(a[2]), .A2(b[5]), .ZN(y[37]) );
  OR2_X1 U70bar ( .A1(abar[2]), .A2(bbar[5]), .ZN(ybar[37]) );
  AND2_X1 U71 ( .A1(a[2]), .A2(b[4]), .ZN(y[36]) );
  OR2_X1 U71bar ( .A1(abar[2]), .A2(bbar[4]), .ZN(ybar[36]) );
  AND2_X1 U72 ( .A1(a[2]), .A2(b[3]), .ZN(y[35]) );
  OR2_X1 U72bar ( .A1(abar[2]), .A2(bbar[3]), .ZN(ybar[35]) );
  AND2_X1 U73 ( .A1(a[2]), .A2(b[2]), .ZN(y[34]) );
  OR2_X1 U73bar ( .A1(abar[2]), .A2(bbar[2]), .ZN(ybar[34]) );
  AND2_X1 U74 ( .A1(a[2]), .A2(b[1]), .ZN(y[33]) );
  OR2_X1 U74bar ( .A1(abar[2]), .A2(bbar[1]), .ZN(ybar[33]) );
  AND2_X1 U75 ( .A1(a[2]), .A2(b[0]), .ZN(y[32]) );
  OR2_X1 U75bar ( .A1(abar[2]), .A2(bbar[0]), .ZN(ybar[32]) );
  AND2_X1 U76 ( .A1(a[1]), .A2(b[15]), .ZN(y[31]) );
  OR2_X1 U76bar ( .A1(abar[1]), .A2(bbar[15]), .ZN(ybar[31]) );
  AND2_X1 U77 ( .A1(a[1]), .A2(b[14]), .ZN(y[30]) );
  OR2_X1 U77bar ( .A1(abar[1]), .A2(bbar[14]), .ZN(ybar[30]) );
  AND2_X1 U78 ( .A1(b[2]), .A2(a[0]), .ZN(y[2]) );
  OR2_X1 U78bar ( .A1(bbar[2]), .A2(abar[0]), .ZN(ybar[2]) );
  AND2_X1 U79 ( .A1(a[1]), .A2(b[13]), .ZN(y[29]) );
  OR2_X1 U79bar ( .A1(abar[1]), .A2(bbar[13]), .ZN(ybar[29]) );
  AND2_X1 U80 ( .A1(a[1]), .A2(b[12]), .ZN(y[28]) );
  OR2_X1 U80bar ( .A1(abar[1]), .A2(bbar[12]), .ZN(ybar[28]) );
  AND2_X1 U81 ( .A1(a[1]), .A2(b[11]), .ZN(y[27]) );
  OR2_X1 U81bar ( .A1(abar[1]), .A2(bbar[11]), .ZN(ybar[27]) );
  AND2_X1 U82 ( .A1(a[1]), .A2(b[10]), .ZN(y[26]) );
  OR2_X1 U82bar ( .A1(abar[1]), .A2(bbar[10]), .ZN(ybar[26]) );
  AND2_X1 U83 ( .A1(a[1]), .A2(b[9]), .ZN(y[25]) );
  OR2_X1 U83bar ( .A1(abar[1]), .A2(bbar[9]), .ZN(ybar[25]) );
  AND2_X1 U84 ( .A1(a[15]), .A2(b[15]), .ZN(y[255]) );
  OR2_X1 U84bar ( .A1(abar[15]), .A2(bbar[15]), .ZN(ybar[255]) );
  AND2_X1 U85 ( .A1(a[15]), .A2(b[14]), .ZN(y[254]) );
  OR2_X1 U85bar ( .A1(abar[15]), .A2(bbar[14]), .ZN(ybar[254]) );
  AND2_X1 U86 ( .A1(a[15]), .A2(b[13]), .ZN(y[253]) );
  OR2_X1 U86bar ( .A1(abar[15]), .A2(bbar[13]), .ZN(ybar[253]) );
  AND2_X1 U87 ( .A1(a[15]), .A2(b[12]), .ZN(y[252]) );
  OR2_X1 U87bar ( .A1(abar[15]), .A2(bbar[12]), .ZN(ybar[252]) );
  AND2_X1 U88 ( .A1(a[15]), .A2(b[11]), .ZN(y[251]) );
  OR2_X1 U88bar ( .A1(abar[15]), .A2(bbar[11]), .ZN(ybar[251]) );
  AND2_X1 U89 ( .A1(a[15]), .A2(b[10]), .ZN(y[250]) );
  OR2_X1 U89bar ( .A1(abar[15]), .A2(bbar[10]), .ZN(ybar[250]) );
  AND2_X1 U90 ( .A1(a[1]), .A2(b[8]), .ZN(y[24]) );
  OR2_X1 U90bar ( .A1(abar[1]), .A2(bbar[8]), .ZN(ybar[24]) );
  AND2_X1 U91 ( .A1(a[15]), .A2(b[9]), .ZN(y[249]) );
  OR2_X1 U91bar ( .A1(abar[15]), .A2(bbar[9]), .ZN(ybar[249]) );
  AND2_X1 U92 ( .A1(a[15]), .A2(b[8]), .ZN(y[248]) );
  OR2_X1 U92bar ( .A1(abar[15]), .A2(bbar[8]), .ZN(ybar[248]) );
  AND2_X1 U93 ( .A1(a[15]), .A2(b[7]), .ZN(y[247]) );
  OR2_X1 U93bar ( .A1(abar[15]), .A2(bbar[7]), .ZN(ybar[247]) );
  AND2_X1 U94 ( .A1(a[15]), .A2(b[6]), .ZN(y[246]) );
  OR2_X1 U94bar ( .A1(abar[15]), .A2(bbar[6]), .ZN(ybar[246]) );
  AND2_X1 U95 ( .A1(a[15]), .A2(b[5]), .ZN(y[245]) );
  OR2_X1 U95bar ( .A1(abar[15]), .A2(bbar[5]), .ZN(ybar[245]) );
  AND2_X1 U96 ( .A1(a[15]), .A2(b[4]), .ZN(y[244]) );
  OR2_X1 U96bar ( .A1(abar[15]), .A2(bbar[4]), .ZN(ybar[244]) );
  AND2_X1 U97 ( .A1(a[15]), .A2(b[3]), .ZN(y[243]) );
  OR2_X1 U97bar ( .A1(abar[15]), .A2(bbar[3]), .ZN(ybar[243]) );
  AND2_X1 U98 ( .A1(a[15]), .A2(b[2]), .ZN(y[242]) );
  OR2_X1 U98bar ( .A1(abar[15]), .A2(bbar[2]), .ZN(ybar[242]) );
  AND2_X1 U99 ( .A1(a[15]), .A2(b[1]), .ZN(y[241]) );
  OR2_X1 U99bar ( .A1(abar[15]), .A2(bbar[1]), .ZN(ybar[241]) );
  AND2_X1 U100 ( .A1(a[15]), .A2(b[0]), .ZN(y[240]) );
  OR2_X1 U100bar ( .A1(abar[15]), .A2(bbar[0]), .ZN(ybar[240]) );
  AND2_X1 U101 ( .A1(a[1]), .A2(b[7]), .ZN(y[23]) );
  OR2_X1 U101bar ( .A1(abar[1]), .A2(bbar[7]), .ZN(ybar[23]) );
  AND2_X1 U102 ( .A1(a[14]), .A2(b[15]), .ZN(y[239]) );
  OR2_X1 U102bar ( .A1(abar[14]), .A2(bbar[15]), .ZN(ybar[239]) );
  AND2_X1 U103 ( .A1(a[14]), .A2(b[14]), .ZN(y[238]) );
  OR2_X1 U103bar ( .A1(abar[14]), .A2(bbar[14]), .ZN(ybar[238]) );
  AND2_X1 U104 ( .A1(a[14]), .A2(b[13]), .ZN(y[237]) );
  OR2_X1 U104bar ( .A1(abar[14]), .A2(bbar[13]), .ZN(ybar[237]) );
  AND2_X1 U105 ( .A1(a[14]), .A2(b[12]), .ZN(y[236]) );
  OR2_X1 U105bar ( .A1(abar[14]), .A2(bbar[12]), .ZN(ybar[236]) );
  AND2_X1 U106 ( .A1(a[14]), .A2(b[11]), .ZN(y[235]) );
  OR2_X1 U106bar ( .A1(abar[14]), .A2(bbar[11]), .ZN(ybar[235]) );
  AND2_X1 U107 ( .A1(a[14]), .A2(b[10]), .ZN(y[234]) );
  OR2_X1 U107bar ( .A1(abar[14]), .A2(bbar[10]), .ZN(ybar[234]) );
  AND2_X1 U108 ( .A1(a[14]), .A2(b[9]), .ZN(y[233]) );
  OR2_X1 U108bar ( .A1(abar[14]), .A2(bbar[9]), .ZN(ybar[233]) );
  AND2_X1 U109 ( .A1(a[14]), .A2(b[8]), .ZN(y[232]) );
  OR2_X1 U109bar ( .A1(abar[14]), .A2(bbar[8]), .ZN(ybar[232]) );
  AND2_X1 U110 ( .A1(a[14]), .A2(b[7]), .ZN(y[231]) );
  OR2_X1 U110bar ( .A1(abar[14]), .A2(bbar[7]), .ZN(ybar[231]) );
  AND2_X1 U111 ( .A1(a[14]), .A2(b[6]), .ZN(y[230]) );
  OR2_X1 U111bar ( .A1(abar[14]), .A2(bbar[6]), .ZN(ybar[230]) );
  AND2_X1 U112 ( .A1(a[1]), .A2(b[6]), .ZN(y[22]) );
  OR2_X1 U112bar ( .A1(abar[1]), .A2(bbar[6]), .ZN(ybar[22]) );
  AND2_X1 U113 ( .A1(a[14]), .A2(b[5]), .ZN(y[229]) );
  OR2_X1 U113bar ( .A1(abar[14]), .A2(bbar[5]), .ZN(ybar[229]) );
  AND2_X1 U114 ( .A1(a[14]), .A2(b[4]), .ZN(y[228]) );
  OR2_X1 U114bar ( .A1(abar[14]), .A2(bbar[4]), .ZN(ybar[228]) );
  AND2_X1 U115 ( .A1(a[14]), .A2(b[3]), .ZN(y[227]) );
  OR2_X1 U115bar ( .A1(abar[14]), .A2(bbar[3]), .ZN(ybar[227]) );
  AND2_X1 U116 ( .A1(a[14]), .A2(b[2]), .ZN(y[226]) );
  OR2_X1 U116bar ( .A1(abar[14]), .A2(bbar[2]), .ZN(ybar[226]) );
  AND2_X1 U117 ( .A1(a[14]), .A2(b[1]), .ZN(y[225]) );
  OR2_X1 U117bar ( .A1(abar[14]), .A2(bbar[1]), .ZN(ybar[225]) );
  AND2_X1 U118 ( .A1(a[14]), .A2(b[0]), .ZN(y[224]) );
  OR2_X1 U118bar ( .A1(abar[14]), .A2(bbar[0]), .ZN(ybar[224]) );
  AND2_X1 U119 ( .A1(a[13]), .A2(b[15]), .ZN(y[223]) );
  OR2_X1 U119bar ( .A1(abar[13]), .A2(bbar[15]), .ZN(ybar[223]) );
  AND2_X1 U120 ( .A1(a[13]), .A2(b[14]), .ZN(y[222]) );
  OR2_X1 U120bar ( .A1(abar[13]), .A2(bbar[14]), .ZN(ybar[222]) );
  AND2_X1 U121 ( .A1(a[13]), .A2(b[13]), .ZN(y[221]) );
  OR2_X1 U121bar ( .A1(abar[13]), .A2(bbar[13]), .ZN(ybar[221]) );
  AND2_X1 U122 ( .A1(a[13]), .A2(b[12]), .ZN(y[220]) );
  OR2_X1 U122bar ( .A1(abar[13]), .A2(bbar[12]), .ZN(ybar[220]) );
  AND2_X1 U123 ( .A1(a[1]), .A2(b[5]), .ZN(y[21]) );
  OR2_X1 U123bar ( .A1(abar[1]), .A2(bbar[5]), .ZN(ybar[21]) );
  AND2_X1 U124 ( .A1(a[13]), .A2(b[11]), .ZN(y[219]) );
  OR2_X1 U124bar ( .A1(abar[13]), .A2(bbar[11]), .ZN(ybar[219]) );
  AND2_X1 U125 ( .A1(a[13]), .A2(b[10]), .ZN(y[218]) );
  OR2_X1 U125bar ( .A1(abar[13]), .A2(bbar[10]), .ZN(ybar[218]) );
  AND2_X1 U126 ( .A1(a[13]), .A2(b[9]), .ZN(y[217]) );
  OR2_X1 U126bar ( .A1(abar[13]), .A2(bbar[9]), .ZN(ybar[217]) );
  AND2_X1 U127 ( .A1(a[13]), .A2(b[8]), .ZN(y[216]) );
  OR2_X1 U127bar ( .A1(abar[13]), .A2(bbar[8]), .ZN(ybar[216]) );
  AND2_X1 U128 ( .A1(a[13]), .A2(b[7]), .ZN(y[215]) );
  OR2_X1 U128bar ( .A1(abar[13]), .A2(bbar[7]), .ZN(ybar[215]) );
  AND2_X1 U129 ( .A1(a[13]), .A2(b[6]), .ZN(y[214]) );
  OR2_X1 U129bar ( .A1(abar[13]), .A2(bbar[6]), .ZN(ybar[214]) );
  AND2_X1 U130 ( .A1(a[13]), .A2(b[5]), .ZN(y[213]) );
  OR2_X1 U130bar ( .A1(abar[13]), .A2(bbar[5]), .ZN(ybar[213]) );
  AND2_X1 U131 ( .A1(a[13]), .A2(b[4]), .ZN(y[212]) );
  OR2_X1 U131bar ( .A1(abar[13]), .A2(bbar[4]), .ZN(ybar[212]) );
  AND2_X1 U132 ( .A1(a[13]), .A2(b[3]), .ZN(y[211]) );
  OR2_X1 U132bar ( .A1(abar[13]), .A2(bbar[3]), .ZN(ybar[211]) );
  AND2_X1 U133 ( .A1(a[13]), .A2(b[2]), .ZN(y[210]) );
  OR2_X1 U133bar ( .A1(abar[13]), .A2(bbar[2]), .ZN(ybar[210]) );
  AND2_X1 U134 ( .A1(a[1]), .A2(b[4]), .ZN(y[20]) );
  OR2_X1 U134bar ( .A1(abar[1]), .A2(bbar[4]), .ZN(ybar[20]) );
  AND2_X1 U135 ( .A1(a[13]), .A2(b[1]), .ZN(y[209]) );
  OR2_X1 U135bar ( .A1(abar[13]), .A2(bbar[1]), .ZN(ybar[209]) );
  AND2_X1 U136 ( .A1(a[13]), .A2(b[0]), .ZN(y[208]) );
  OR2_X1 U136bar ( .A1(abar[13]), .A2(bbar[0]), .ZN(ybar[208]) );
  AND2_X1 U137 ( .A1(a[12]), .A2(b[15]), .ZN(y[207]) );
  OR2_X1 U137bar ( .A1(abar[12]), .A2(bbar[15]), .ZN(ybar[207]) );
  AND2_X1 U138 ( .A1(a[12]), .A2(b[14]), .ZN(y[206]) );
  OR2_X1 U138bar ( .A1(abar[12]), .A2(bbar[14]), .ZN(ybar[206]) );
  AND2_X1 U139 ( .A1(a[12]), .A2(b[13]), .ZN(y[205]) );
  OR2_X1 U139bar ( .A1(abar[12]), .A2(bbar[13]), .ZN(ybar[205]) );
  AND2_X1 U140 ( .A1(a[12]), .A2(b[12]), .ZN(y[204]) );
  OR2_X1 U140bar ( .A1(abar[12]), .A2(bbar[12]), .ZN(ybar[204]) );
  AND2_X1 U141 ( .A1(a[12]), .A2(b[11]), .ZN(y[203]) );
  OR2_X1 U141bar ( .A1(abar[12]), .A2(bbar[11]), .ZN(ybar[203]) );
  AND2_X1 U142 ( .A1(a[12]), .A2(b[10]), .ZN(y[202]) );
  OR2_X1 U142bar ( .A1(abar[12]), .A2(bbar[10]), .ZN(ybar[202]) );
  AND2_X1 U143 ( .A1(a[12]), .A2(b[9]), .ZN(y[201]) );
  OR2_X1 U143bar ( .A1(abar[12]), .A2(bbar[9]), .ZN(ybar[201]) );
  AND2_X1 U144 ( .A1(a[12]), .A2(b[8]), .ZN(y[200]) );
  OR2_X1 U144bar ( .A1(abar[12]), .A2(bbar[8]), .ZN(ybar[200]) );
  AND2_X1 U145 ( .A1(b[1]), .A2(a[0]), .ZN(y[1]) );
  OR2_X1 U145bar ( .A1(bbar[1]), .A2(abar[0]), .ZN(ybar[1]) );
  AND2_X1 U146 ( .A1(a[1]), .A2(b[3]), .ZN(y[19]) );
  OR2_X1 U146bar ( .A1(abar[1]), .A2(bbar[3]), .ZN(ybar[19]) );
  AND2_X1 U147 ( .A1(a[12]), .A2(b[7]), .ZN(y[199]) );
  OR2_X1 U147bar ( .A1(abar[12]), .A2(bbar[7]), .ZN(ybar[199]) );
  AND2_X1 U148 ( .A1(a[12]), .A2(b[6]), .ZN(y[198]) );
  OR2_X1 U148bar ( .A1(abar[12]), .A2(bbar[6]), .ZN(ybar[198]) );
  AND2_X1 U149 ( .A1(a[12]), .A2(b[5]), .ZN(y[197]) );
  OR2_X1 U149bar ( .A1(abar[12]), .A2(bbar[5]), .ZN(ybar[197]) );
  AND2_X1 U150 ( .A1(a[12]), .A2(b[4]), .ZN(y[196]) );
  OR2_X1 U150bar ( .A1(abar[12]), .A2(bbar[4]), .ZN(ybar[196]) );
  AND2_X1 U151 ( .A1(a[12]), .A2(b[3]), .ZN(y[195]) );
  OR2_X1 U151bar ( .A1(abar[12]), .A2(bbar[3]), .ZN(ybar[195]) );
  AND2_X1 U152 ( .A1(a[12]), .A2(b[2]), .ZN(y[194]) );
  OR2_X1 U152bar ( .A1(abar[12]), .A2(bbar[2]), .ZN(ybar[194]) );
  AND2_X1 U153 ( .A1(a[12]), .A2(b[1]), .ZN(y[193]) );
  OR2_X1 U153bar ( .A1(abar[12]), .A2(bbar[1]), .ZN(ybar[193]) );
  AND2_X1 U154 ( .A1(a[12]), .A2(b[0]), .ZN(y[192]) );
  OR2_X1 U154bar ( .A1(abar[12]), .A2(bbar[0]), .ZN(ybar[192]) );
  AND2_X1 U155 ( .A1(a[11]), .A2(b[15]), .ZN(y[191]) );
  OR2_X1 U155bar ( .A1(abar[11]), .A2(bbar[15]), .ZN(ybar[191]) );
  AND2_X1 U156 ( .A1(a[11]), .A2(b[14]), .ZN(y[190]) );
  OR2_X1 U156bar ( .A1(abar[11]), .A2(bbar[14]), .ZN(ybar[190]) );
  AND2_X1 U157 ( .A1(a[1]), .A2(b[2]), .ZN(y[18]) );
  OR2_X1 U157bar ( .A1(abar[1]), .A2(bbar[2]), .ZN(ybar[18]) );
  AND2_X1 U158 ( .A1(a[11]), .A2(b[13]), .ZN(y[189]) );
  OR2_X1 U158bar ( .A1(abar[11]), .A2(bbar[13]), .ZN(ybar[189]) );
  AND2_X1 U159 ( .A1(a[11]), .A2(b[12]), .ZN(y[188]) );
  OR2_X1 U159bar ( .A1(abar[11]), .A2(bbar[12]), .ZN(ybar[188]) );
  AND2_X1 U160 ( .A1(a[11]), .A2(b[11]), .ZN(y[187]) );
  OR2_X1 U160bar ( .A1(abar[11]), .A2(bbar[11]), .ZN(ybar[187]) );
  AND2_X1 U161 ( .A1(a[11]), .A2(b[10]), .ZN(y[186]) );
  OR2_X1 U161bar ( .A1(abar[11]), .A2(bbar[10]), .ZN(ybar[186]) );
  AND2_X1 U162 ( .A1(a[11]), .A2(b[9]), .ZN(y[185]) );
  OR2_X1 U162bar ( .A1(abar[11]), .A2(bbar[9]), .ZN(ybar[185]) );
  AND2_X1 U163 ( .A1(a[11]), .A2(b[8]), .ZN(y[184]) );
  OR2_X1 U163bar ( .A1(abar[11]), .A2(bbar[8]), .ZN(ybar[184]) );
  AND2_X1 U164 ( .A1(a[11]), .A2(b[7]), .ZN(y[183]) );
  OR2_X1 U164bar ( .A1(abar[11]), .A2(bbar[7]), .ZN(ybar[183]) );
  AND2_X1 U165 ( .A1(a[11]), .A2(b[6]), .ZN(y[182]) );
  OR2_X1 U165bar ( .A1(abar[11]), .A2(bbar[6]), .ZN(ybar[182]) );
  AND2_X1 U166 ( .A1(a[11]), .A2(b[5]), .ZN(y[181]) );
  OR2_X1 U166bar ( .A1(abar[11]), .A2(bbar[5]), .ZN(ybar[181]) );
  AND2_X1 U167 ( .A1(a[11]), .A2(b[4]), .ZN(y[180]) );
  OR2_X1 U167bar ( .A1(abar[11]), .A2(bbar[4]), .ZN(ybar[180]) );
  AND2_X1 U168 ( .A1(a[1]), .A2(b[1]), .ZN(y[17]) );
  OR2_X1 U168bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[17]) );
  AND2_X1 U169 ( .A1(a[11]), .A2(b[3]), .ZN(y[179]) );
  OR2_X1 U169bar ( .A1(abar[11]), .A2(bbar[3]), .ZN(ybar[179]) );
  AND2_X1 U170 ( .A1(a[11]), .A2(b[2]), .ZN(y[178]) );
  OR2_X1 U170bar ( .A1(abar[11]), .A2(bbar[2]), .ZN(ybar[178]) );
  AND2_X1 U171 ( .A1(a[11]), .A2(b[1]), .ZN(y[177]) );
  OR2_X1 U171bar ( .A1(abar[11]), .A2(bbar[1]), .ZN(ybar[177]) );
  AND2_X1 U172 ( .A1(a[11]), .A2(b[0]), .ZN(y[176]) );
  OR2_X1 U172bar ( .A1(abar[11]), .A2(bbar[0]), .ZN(ybar[176]) );
  AND2_X1 U173 ( .A1(a[10]), .A2(b[15]), .ZN(y[175]) );
  OR2_X1 U173bar ( .A1(abar[10]), .A2(bbar[15]), .ZN(ybar[175]) );
  AND2_X1 U174 ( .A1(a[10]), .A2(b[14]), .ZN(y[174]) );
  OR2_X1 U174bar ( .A1(abar[10]), .A2(bbar[14]), .ZN(ybar[174]) );
  AND2_X1 U175 ( .A1(a[10]), .A2(b[13]), .ZN(y[173]) );
  OR2_X1 U175bar ( .A1(abar[10]), .A2(bbar[13]), .ZN(ybar[173]) );
  AND2_X1 U176 ( .A1(a[10]), .A2(b[12]), .ZN(y[172]) );
  OR2_X1 U176bar ( .A1(abar[10]), .A2(bbar[12]), .ZN(ybar[172]) );
  AND2_X1 U177 ( .A1(a[10]), .A2(b[11]), .ZN(y[171]) );
  OR2_X1 U177bar ( .A1(abar[10]), .A2(bbar[11]), .ZN(ybar[171]) );
  AND2_X1 U178 ( .A1(a[10]), .A2(b[10]), .ZN(y[170]) );
  OR2_X1 U178bar ( .A1(abar[10]), .A2(bbar[10]), .ZN(ybar[170]) );
  AND2_X1 U179 ( .A1(a[1]), .A2(b[0]), .ZN(y[16]) );
  OR2_X1 U179bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[16]) );
  AND2_X1 U180 ( .A1(a[10]), .A2(b[9]), .ZN(y[169]) );
  OR2_X1 U180bar ( .A1(abar[10]), .A2(bbar[9]), .ZN(ybar[169]) );
  AND2_X1 U181 ( .A1(a[10]), .A2(b[8]), .ZN(y[168]) );
  OR2_X1 U181bar ( .A1(abar[10]), .A2(bbar[8]), .ZN(ybar[168]) );
  AND2_X1 U182 ( .A1(a[10]), .A2(b[7]), .ZN(y[167]) );
  OR2_X1 U182bar ( .A1(abar[10]), .A2(bbar[7]), .ZN(ybar[167]) );
  AND2_X1 U183 ( .A1(a[10]), .A2(b[6]), .ZN(y[166]) );
  OR2_X1 U183bar ( .A1(abar[10]), .A2(bbar[6]), .ZN(ybar[166]) );
  AND2_X1 U184 ( .A1(a[10]), .A2(b[5]), .ZN(y[165]) );
  OR2_X1 U184bar ( .A1(abar[10]), .A2(bbar[5]), .ZN(ybar[165]) );
  AND2_X1 U185 ( .A1(a[10]), .A2(b[4]), .ZN(y[164]) );
  OR2_X1 U185bar ( .A1(abar[10]), .A2(bbar[4]), .ZN(ybar[164]) );
  AND2_X1 U186 ( .A1(a[10]), .A2(b[3]), .ZN(y[163]) );
  OR2_X1 U186bar ( .A1(abar[10]), .A2(bbar[3]), .ZN(ybar[163]) );
  AND2_X1 U187 ( .A1(a[10]), .A2(b[2]), .ZN(y[162]) );
  OR2_X1 U187bar ( .A1(abar[10]), .A2(bbar[2]), .ZN(ybar[162]) );
  AND2_X1 U188 ( .A1(a[10]), .A2(b[1]), .ZN(y[161]) );
  OR2_X1 U188bar ( .A1(abar[10]), .A2(bbar[1]), .ZN(ybar[161]) );
  AND2_X1 U189 ( .A1(a[10]), .A2(b[0]), .ZN(y[160]) );
  OR2_X1 U189bar ( .A1(abar[10]), .A2(bbar[0]), .ZN(ybar[160]) );
  AND2_X1 U190 ( .A1(b[15]), .A2(a[0]), .ZN(y[15]) );
  OR2_X1 U190bar ( .A1(bbar[15]), .A2(abar[0]), .ZN(ybar[15]) );
  AND2_X1 U191 ( .A1(a[9]), .A2(b[15]), .ZN(y[159]) );
  OR2_X1 U191bar ( .A1(abar[9]), .A2(bbar[15]), .ZN(ybar[159]) );
  AND2_X1 U192 ( .A1(a[9]), .A2(b[14]), .ZN(y[158]) );
  OR2_X1 U192bar ( .A1(abar[9]), .A2(bbar[14]), .ZN(ybar[158]) );
  AND2_X1 U193 ( .A1(a[9]), .A2(b[13]), .ZN(y[157]) );
  OR2_X1 U193bar ( .A1(abar[9]), .A2(bbar[13]), .ZN(ybar[157]) );
  AND2_X1 U194 ( .A1(a[9]), .A2(b[12]), .ZN(y[156]) );
  OR2_X1 U194bar ( .A1(abar[9]), .A2(bbar[12]), .ZN(ybar[156]) );
  AND2_X1 U195 ( .A1(a[9]), .A2(b[11]), .ZN(y[155]) );
  OR2_X1 U195bar ( .A1(abar[9]), .A2(bbar[11]), .ZN(ybar[155]) );
  AND2_X1 U196 ( .A1(a[9]), .A2(b[10]), .ZN(y[154]) );
  OR2_X1 U196bar ( .A1(abar[9]), .A2(bbar[10]), .ZN(ybar[154]) );
  AND2_X1 U197 ( .A1(a[9]), .A2(b[9]), .ZN(y[153]) );
  OR2_X1 U197bar ( .A1(abar[9]), .A2(bbar[9]), .ZN(ybar[153]) );
  AND2_X1 U198 ( .A1(a[9]), .A2(b[8]), .ZN(y[152]) );
  OR2_X1 U198bar ( .A1(abar[9]), .A2(bbar[8]), .ZN(ybar[152]) );
  AND2_X1 U199 ( .A1(a[9]), .A2(b[7]), .ZN(y[151]) );
  OR2_X1 U199bar ( .A1(abar[9]), .A2(bbar[7]), .ZN(ybar[151]) );
  AND2_X1 U200 ( .A1(a[9]), .A2(b[6]), .ZN(y[150]) );
  OR2_X1 U200bar ( .A1(abar[9]), .A2(bbar[6]), .ZN(ybar[150]) );
  AND2_X1 U201 ( .A1(b[14]), .A2(a[0]), .ZN(y[14]) );
  OR2_X1 U201bar ( .A1(bbar[14]), .A2(abar[0]), .ZN(ybar[14]) );
  AND2_X1 U202 ( .A1(a[9]), .A2(b[5]), .ZN(y[149]) );
  OR2_X1 U202bar ( .A1(abar[9]), .A2(bbar[5]), .ZN(ybar[149]) );
  AND2_X1 U203 ( .A1(a[9]), .A2(b[4]), .ZN(y[148]) );
  OR2_X1 U203bar ( .A1(abar[9]), .A2(bbar[4]), .ZN(ybar[148]) );
  AND2_X1 U204 ( .A1(a[9]), .A2(b[3]), .ZN(y[147]) );
  OR2_X1 U204bar ( .A1(abar[9]), .A2(bbar[3]), .ZN(ybar[147]) );
  AND2_X1 U205 ( .A1(a[9]), .A2(b[2]), .ZN(y[146]) );
  OR2_X1 U205bar ( .A1(abar[9]), .A2(bbar[2]), .ZN(ybar[146]) );
  AND2_X1 U206 ( .A1(a[9]), .A2(b[1]), .ZN(y[145]) );
  OR2_X1 U206bar ( .A1(abar[9]), .A2(bbar[1]), .ZN(ybar[145]) );
  AND2_X1 U207 ( .A1(a[9]), .A2(b[0]), .ZN(y[144]) );
  OR2_X1 U207bar ( .A1(abar[9]), .A2(bbar[0]), .ZN(ybar[144]) );
  AND2_X1 U208 ( .A1(a[8]), .A2(b[15]), .ZN(y[143]) );
  OR2_X1 U208bar ( .A1(abar[8]), .A2(bbar[15]), .ZN(ybar[143]) );
  AND2_X1 U209 ( .A1(a[8]), .A2(b[14]), .ZN(y[142]) );
  OR2_X1 U209bar ( .A1(abar[8]), .A2(bbar[14]), .ZN(ybar[142]) );
  AND2_X1 U210 ( .A1(a[8]), .A2(b[13]), .ZN(y[141]) );
  OR2_X1 U210bar ( .A1(abar[8]), .A2(bbar[13]), .ZN(ybar[141]) );
  AND2_X1 U211 ( .A1(a[8]), .A2(b[12]), .ZN(y[140]) );
  OR2_X1 U211bar ( .A1(abar[8]), .A2(bbar[12]), .ZN(ybar[140]) );
  AND2_X1 U212 ( .A1(b[13]), .A2(a[0]), .ZN(y[13]) );
  OR2_X1 U212bar ( .A1(bbar[13]), .A2(abar[0]), .ZN(ybar[13]) );
  AND2_X1 U213 ( .A1(a[8]), .A2(b[11]), .ZN(y[139]) );
  OR2_X1 U213bar ( .A1(abar[8]), .A2(bbar[11]), .ZN(ybar[139]) );
  AND2_X1 U214 ( .A1(a[8]), .A2(b[10]), .ZN(y[138]) );
  OR2_X1 U214bar ( .A1(abar[8]), .A2(bbar[10]), .ZN(ybar[138]) );
  AND2_X1 U215 ( .A1(a[8]), .A2(b[9]), .ZN(y[137]) );
  OR2_X1 U215bar ( .A1(abar[8]), .A2(bbar[9]), .ZN(ybar[137]) );
  AND2_X1 U216 ( .A1(a[8]), .A2(b[8]), .ZN(y[136]) );
  OR2_X1 U216bar ( .A1(abar[8]), .A2(bbar[8]), .ZN(ybar[136]) );
  AND2_X1 U217 ( .A1(a[8]), .A2(b[7]), .ZN(y[135]) );
  OR2_X1 U217bar ( .A1(abar[8]), .A2(bbar[7]), .ZN(ybar[135]) );
  AND2_X1 U218 ( .A1(a[8]), .A2(b[6]), .ZN(y[134]) );
  OR2_X1 U218bar ( .A1(abar[8]), .A2(bbar[6]), .ZN(ybar[134]) );
  AND2_X1 U219 ( .A1(a[8]), .A2(b[5]), .ZN(y[133]) );
  OR2_X1 U219bar ( .A1(abar[8]), .A2(bbar[5]), .ZN(ybar[133]) );
  AND2_X1 U220 ( .A1(a[8]), .A2(b[4]), .ZN(y[132]) );
  OR2_X1 U220bar ( .A1(abar[8]), .A2(bbar[4]), .ZN(ybar[132]) );
  AND2_X1 U221 ( .A1(a[8]), .A2(b[3]), .ZN(y[131]) );
  OR2_X1 U221bar ( .A1(abar[8]), .A2(bbar[3]), .ZN(ybar[131]) );
  AND2_X1 U222 ( .A1(a[8]), .A2(b[2]), .ZN(y[130]) );
  OR2_X1 U222bar ( .A1(abar[8]), .A2(bbar[2]), .ZN(ybar[130]) );
  AND2_X1 U223 ( .A1(b[12]), .A2(a[0]), .ZN(y[12]) );
  OR2_X1 U223bar ( .A1(bbar[12]), .A2(abar[0]), .ZN(ybar[12]) );
  AND2_X1 U224 ( .A1(a[8]), .A2(b[1]), .ZN(y[129]) );
  OR2_X1 U224bar ( .A1(abar[8]), .A2(bbar[1]), .ZN(ybar[129]) );
  AND2_X1 U225 ( .A1(a[8]), .A2(b[0]), .ZN(y[128]) );
  OR2_X1 U225bar ( .A1(abar[8]), .A2(bbar[0]), .ZN(ybar[128]) );
  AND2_X1 U226 ( .A1(a[7]), .A2(b[15]), .ZN(y[127]) );
  OR2_X1 U226bar ( .A1(abar[7]), .A2(bbar[15]), .ZN(ybar[127]) );
  AND2_X1 U227 ( .A1(a[7]), .A2(b[14]), .ZN(y[126]) );
  OR2_X1 U227bar ( .A1(abar[7]), .A2(bbar[14]), .ZN(ybar[126]) );
  AND2_X1 U228 ( .A1(a[7]), .A2(b[13]), .ZN(y[125]) );
  OR2_X1 U228bar ( .A1(abar[7]), .A2(bbar[13]), .ZN(ybar[125]) );
  AND2_X1 U229 ( .A1(a[7]), .A2(b[12]), .ZN(y[124]) );
  OR2_X1 U229bar ( .A1(abar[7]), .A2(bbar[12]), .ZN(ybar[124]) );
  AND2_X1 U230 ( .A1(a[7]), .A2(b[11]), .ZN(y[123]) );
  OR2_X1 U230bar ( .A1(abar[7]), .A2(bbar[11]), .ZN(ybar[123]) );
  AND2_X1 U231 ( .A1(a[7]), .A2(b[10]), .ZN(y[122]) );
  OR2_X1 U231bar ( .A1(abar[7]), .A2(bbar[10]), .ZN(ybar[122]) );
  AND2_X1 U232 ( .A1(a[7]), .A2(b[9]), .ZN(y[121]) );
  OR2_X1 U232bar ( .A1(abar[7]), .A2(bbar[9]), .ZN(ybar[121]) );
  AND2_X1 U233 ( .A1(a[7]), .A2(b[8]), .ZN(y[120]) );
  OR2_X1 U233bar ( .A1(abar[7]), .A2(bbar[8]), .ZN(ybar[120]) );
  AND2_X1 U234 ( .A1(b[11]), .A2(a[0]), .ZN(y[11]) );
  OR2_X1 U234bar ( .A1(bbar[11]), .A2(abar[0]), .ZN(ybar[11]) );
  AND2_X1 U235 ( .A1(a[7]), .A2(b[7]), .ZN(y[119]) );
  OR2_X1 U235bar ( .A1(abar[7]), .A2(bbar[7]), .ZN(ybar[119]) );
  AND2_X1 U236 ( .A1(a[7]), .A2(b[6]), .ZN(y[118]) );
  OR2_X1 U236bar ( .A1(abar[7]), .A2(bbar[6]), .ZN(ybar[118]) );
  AND2_X1 U237 ( .A1(a[7]), .A2(b[5]), .ZN(y[117]) );
  OR2_X1 U237bar ( .A1(abar[7]), .A2(bbar[5]), .ZN(ybar[117]) );
  AND2_X1 U238 ( .A1(a[7]), .A2(b[4]), .ZN(y[116]) );
  OR2_X1 U238bar ( .A1(abar[7]), .A2(bbar[4]), .ZN(ybar[116]) );
  AND2_X1 U239 ( .A1(a[7]), .A2(b[3]), .ZN(y[115]) );
  OR2_X1 U239bar ( .A1(abar[7]), .A2(bbar[3]), .ZN(ybar[115]) );
  AND2_X1 U240 ( .A1(a[7]), .A2(b[2]), .ZN(y[114]) );
  OR2_X1 U240bar ( .A1(abar[7]), .A2(bbar[2]), .ZN(ybar[114]) );
  AND2_X1 U241 ( .A1(a[7]), .A2(b[1]), .ZN(y[113]) );
  OR2_X1 U241bar ( .A1(abar[7]), .A2(bbar[1]), .ZN(ybar[113]) );
  AND2_X1 U242 ( .A1(a[7]), .A2(b[0]), .ZN(y[112]) );
  OR2_X1 U242bar ( .A1(abar[7]), .A2(bbar[0]), .ZN(ybar[112]) );
  AND2_X1 U243 ( .A1(b[15]), .A2(a[6]), .ZN(y[111]) );
  OR2_X1 U243bar ( .A1(bbar[15]), .A2(abar[6]), .ZN(ybar[111]) );
  AND2_X1 U244 ( .A1(b[14]), .A2(a[6]), .ZN(y[110]) );
  OR2_X1 U244bar ( .A1(bbar[14]), .A2(abar[6]), .ZN(ybar[110]) );
  AND2_X1 U245 ( .A1(b[10]), .A2(a[0]), .ZN(y[10]) );
  OR2_X1 U245bar ( .A1(bbar[10]), .A2(abar[0]), .ZN(ybar[10]) );
  AND2_X1 U246 ( .A1(b[13]), .A2(a[6]), .ZN(y[109]) );
  OR2_X1 U246bar ( .A1(bbar[13]), .A2(abar[6]), .ZN(ybar[109]) );
  AND2_X1 U247 ( .A1(b[12]), .A2(a[6]), .ZN(y[108]) );
  OR2_X1 U247bar ( .A1(bbar[12]), .A2(abar[6]), .ZN(ybar[108]) );
  AND2_X1 U248 ( .A1(b[11]), .A2(a[6]), .ZN(y[107]) );
  OR2_X1 U248bar ( .A1(bbar[11]), .A2(abar[6]), .ZN(ybar[107]) );
  AND2_X1 U249 ( .A1(b[10]), .A2(a[6]), .ZN(y[106]) );
  OR2_X1 U249bar ( .A1(bbar[10]), .A2(abar[6]), .ZN(ybar[106]) );
  AND2_X1 U250 ( .A1(a[6]), .A2(b[9]), .ZN(y[105]) );
  OR2_X1 U250bar ( .A1(abar[6]), .A2(bbar[9]), .ZN(ybar[105]) );
  AND2_X1 U251 ( .A1(b[8]), .A2(a[6]), .ZN(y[104]) );
  OR2_X1 U251bar ( .A1(bbar[8]), .A2(abar[6]), .ZN(ybar[104]) );
  AND2_X1 U252 ( .A1(b[7]), .A2(a[6]), .ZN(y[103]) );
  OR2_X1 U252bar ( .A1(bbar[7]), .A2(abar[6]), .ZN(ybar[103]) );
  AND2_X1 U253 ( .A1(b[6]), .A2(a[6]), .ZN(y[102]) );
  OR2_X1 U253bar ( .A1(bbar[6]), .A2(abar[6]), .ZN(ybar[102]) );
  AND2_X1 U254 ( .A1(b[5]), .A2(a[6]), .ZN(y[101]) );
  OR2_X1 U254bar ( .A1(bbar[5]), .A2(abar[6]), .ZN(ybar[101]) );
  AND2_X1 U255 ( .A1(b[4]), .A2(a[6]), .ZN(y[100]) );
  OR2_X1 U255bar ( .A1(bbar[4]), .A2(abar[6]), .ZN(ybar[100]) );
  AND2_X1 U256 ( .A1(b[0]), .A2(a[0]), .ZN(y[0]) );
  OR2_X1 U256bar ( .A1(bbar[0]), .A2(abar[0]), .ZN(ybar[0]) );
endmodule

module decode_10 ( in, inbar, out, outbar );

  input wire [7:0] in;
  input wire [7:0] inbar;
//input_done

  output wire [255:0] out;
  output wire [255:0] outbar;
//output_done

  wire [15:0] level1;
  wire [31:0] level2;
  wire [15:0] level1bar;
  wire [31:0] level2bar;
//wire_done

  CD2_40 cd_l1_1 ( .a(in[1]), .abar(inbar[1]), .b(in[0]), .bbar(inbar[0]), .y(level1[3:0]), .ybar(level1bar[3:0]) );
  CD2_39 cd_l1_2 ( .a(in[3]), .abar(inbar[3]), .b(in[2]), .bbar(inbar[2]), .y(level1[7:4]), .ybar(level1bar[7:4]) );
  CD2_38 cd_l1_3 ( .a(in[5]), .abar(inbar[5]), .b(in[4]), .bbar(inbar[4]), .y(level1[11:8]), .ybar(level1bar[11:8]) );
  CD2_37 cd_l1_4 ( .a(in[7]), .abar(inbar[7]), .b(in[6]), .bbar(inbar[6]), .y(level1[15:12]), .ybar(level1bar[15:12]) );

  CD4_20 cd_l2_1 ( .a(level1[7:4]), .abar(level1bar[7:4]), .b(level1[3:0]), .bbar(level1bar[3:0]), 
        .y(level2[15:0]), .ybar(level2bar[15:0]) );
  CD4_19 cd_l2_2 ( .a(level1[15:12]), .abar(level1bar[15:12]), .b(level1[11:8]), .bbar(level1bar[11:8]), 
        .y(level2[31:16]), .ybar(level2bar[31:16]) );
  CD16_10 cd_l3 ( .a(level2[31:16]), .abar(level2bar[31:16]), .b(level2[15:0]), .bbar(level2bar[15:0]), 
        .y(out), .ybar(outbar) );
endmodule

module encode_10 ( in, inbar, out, outbar );

  input wire [255:0] in;
  input wire [255:0] inbar;
//input_done

  output wire [7:0] out;
  output wire [7:0] outbar;
//output_done

  wire in_81;
  wire in_80;
  wire in_79;
  wire in_78;
  wire in_77;
  wire in_76;
  wire in_75;
  wire in_74;
  wire in_73;
  wire in_72;
  wire in_71;
  wire in_70;
  wire in_69;
  wire in_68;
  wire in_67;
  wire in_66;
  wire in_65;
  wire in_64;
  wire in_63;
  wire in_62;
  wire in_61;
  wire in_60;
  wire in_59;
  wire in_58;
  wire in_57;
  wire in_56;
  wire in_55;
  wire in_54;
  wire in_53;
  wire in_52;
  wire in_51;
  wire in_50;
  wire in_49;
  wire in_48;
  wire in_47;
  wire in_46;
  wire in_45;
  wire in_44;
  wire in_43;
  wire in_42;
  wire in_41;
  wire in_40;
  wire in_39;
  wire in_38;
  wire in_37;
  wire in_36;
  wire in_35;
  wire in_34;
  wire in_33;
  wire in_32;
  wire in_31;
  wire in_30;
  wire in_29;
  wire in_28;
  wire in_27;
  wire in_26;
  wire in_25;
  wire in_24;
  wire in_23;
  wire in_22;
  wire in_21;
  wire in_20;
  wire in_19;
  wire in_18;
  wire in_17;
  wire in_16;
  wire in_15;
  wire in_14;
  wire in_13;
  wire in_12;
  wire in_11;
  wire in_10;
  wire in_9;
  wire in_8;
  wire in_7;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_3;
  wire in_2;
  wire in_1;
  wire in_0;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire in_81bar;
  wire in_80bar;
  wire in_79bar;
  wire in_78bar;
  wire in_77bar;
  wire in_76bar;
  wire in_75bar;
  wire in_74bar;
  wire in_73bar;
  wire in_72bar;
  wire in_71bar;
  wire in_70bar;
  wire in_69bar;
  wire in_68bar;
  wire in_67bar;
  wire in_66bar;
  wire in_65bar;
  wire in_64bar;
  wire in_63bar;
  wire in_62bar;
  wire in_61bar;
  wire in_60bar;
  wire in_59bar;
  wire in_58bar;
  wire in_57bar;
  wire in_56bar;
  wire in_55bar;
  wire in_54bar;
  wire in_53bar;
  wire in_52bar;
  wire in_51bar;
  wire in_50bar;
  wire in_49bar;
  wire in_48bar;
  wire in_47bar;
  wire in_46bar;
  wire in_45bar;
  wire in_44bar;
  wire in_43bar;
  wire in_42bar;
  wire in_41bar;
  wire in_40bar;
  wire in_39bar;
  wire in_38bar;
  wire in_37bar;
  wire in_36bar;
  wire in_35bar;
  wire in_34bar;
  wire in_33bar;
  wire in_32bar;
  wire in_31bar;
  wire in_30bar;
  wire in_29bar;
  wire in_28bar;
  wire in_27bar;
  wire in_26bar;
  wire in_25bar;
  wire in_24bar;
  wire in_23bar;
  wire in_22bar;
  wire in_21bar;
  wire in_20bar;
  wire in_19bar;
  wire in_18bar;
  wire in_17bar;
  wire in_16bar;
  wire in_15bar;
  wire in_14bar;
  wire in_13bar;
  wire in_12bar;
  wire in_11bar;
  wire in_10bar;
  wire in_9bar;
  wire in_8bar;
  wire in_7bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_3bar;
  wire in_2bar;
  wire in_1bar;
  wire in_0bar;
  wire n487bar;
  wire n488bar;
  wire n489bar;
  wire n490bar;
  wire n491bar;
  wire n492bar;
  wire n493bar;
  wire n494bar;
  wire n495bar;
  wire n496bar;
  wire n497bar;
  wire n498bar;
  wire n499bar;
  wire n500bar;
  wire n501bar;
  wire n502bar;
  wire n503bar;
  wire n504bar;
  wire n505bar;
  wire n506bar;
  wire n507bar;
  wire n508bar;
  wire n509bar;
  wire n510bar;
  wire n511bar;
  wire n512bar;
  wire n513bar;
  wire n514bar;
  wire n515bar;
  wire n516bar;
  wire n517bar;
  wire n518bar;
  wire n519bar;
  wire n520bar;
  wire n521bar;
  wire n522bar;
  wire n523bar;
  wire n524bar;
  wire n525bar;
  wire n526bar;
  wire n527bar;
  wire n528bar;
  wire n529bar;
  wire n530bar;
  wire n531bar;
  wire n532bar;
  wire n533bar;
  wire n534bar;
  wire n535bar;
  wire n536bar;
  wire n537bar;
  wire n538bar;
  wire n539bar;
  wire n540bar;
  wire n541bar;
  wire n542bar;
  wire n543bar;
  wire n544bar;
  wire n545bar;
  wire n546bar;
  wire n547bar;
  wire n548bar;
  wire n549bar;
  wire n550bar;
  wire n551bar;
  wire n552bar;
  wire n553bar;
  wire n554bar;
  wire n555bar;
  wire n556bar;
  wire n557bar;
  wire n558bar;
  wire n559bar;
  wire n560bar;
  wire n561bar;
  wire n562bar;
  wire n563bar;
  wire n564bar;
  wire n565bar;
  wire n566bar;
  wire n567bar;
  wire n568bar;
  wire n569bar;
  wire n570bar;
  wire n571bar;
  wire n572bar;
  wire n573bar;
  wire n574bar;
  wire n575bar;
  wire n576bar;
  wire n577bar;
  wire n578bar;
  wire n579bar;
  wire n580bar;
  wire n581bar;
  wire n582bar;
  wire n583bar;
  wire n584bar;
  wire n585bar;
  wire n586bar;
  wire n587bar;
  wire n588bar;
  wire n589bar;
  wire n590bar;
  wire n591bar;
  wire n592bar;
  wire n593bar;
  wire n594bar;
  wire n595bar;
  wire n596bar;
  wire n597bar;
  wire n598bar;
  wire n599bar;
  wire n600bar;
  wire n601bar;
  wire n602bar;
  wire n603bar;
  wire n604bar;
  wire n605bar;
  wire n606bar;
  wire n607bar;
  wire n608bar;
  wire n609bar;
  wire n610bar;
  wire n611bar;
  wire n612bar;
  wire n613bar;
  wire n614bar;
  wire n615bar;
  wire n616bar;
  wire n617bar;
  wire n618bar;
  wire n619bar;
  wire n620bar;
  wire n621bar;
  wire n622bar;
  wire n623bar;
  wire n624bar;
  wire n625bar;
  wire n626bar;
  wire n627bar;
  wire n628bar;
  wire n629bar;
  wire n630bar;
  wire n631bar;
  wire n632bar;
  wire n633bar;
  wire n634bar;
  wire n635bar;
  wire n636bar;
  wire n637bar;
  wire n638bar;
  wire n639bar;
  wire n640bar;
  wire n641bar;
  wire n642bar;
  wire n643bar;
  wire n644bar;
  wire n645bar;
  wire n646bar;
  wire n647bar;
  wire n648bar;
  wire n649bar;
  wire n650bar;
  wire n651bar;
  wire n652bar;
  wire n653bar;
  wire n654bar;
  wire n655bar;
  wire n656bar;
  wire n657bar;
  wire n658bar;
  wire n659bar;
  wire n660bar;
  wire n661bar;
  wire n662bar;
  wire n663bar;
  wire n664bar;
  wire n665bar;
  wire n666bar;
  wire n667bar;
  wire n668bar;
  wire n669bar;
  wire n670bar;
  wire n671bar;
  wire n672bar;
  wire n673bar;
  wire n674bar;
  wire n675bar;
  wire n676bar;
  wire n677bar;
  wire n678bar;
  wire n679bar;
  wire n680bar;
  wire n681bar;
  wire n682bar;
  wire n683bar;
  wire n684bar;
  wire n685bar;
  wire n686bar;
  wire n687bar;
  wire n688bar;
  wire n689bar;
  wire n690bar;
  wire n691bar;
  wire n692bar;
  wire n693bar;
  wire n694bar;
  wire n695bar;
  wire n696bar;
  wire n697bar;
  wire n698bar;
  wire n699bar;
  wire n700bar;
  wire n701bar;
  wire n702bar;
  wire n703bar;
  wire n704bar;
  wire n705bar;
  wire n706bar;
  wire n707bar;
  wire n708bar;
  wire n709bar;
  wire n710bar;
  wire n711bar;
  wire n712bar;
  wire n713bar;
  wire n714bar;
  wire n715bar;
  wire n716bar;
  wire n717bar;
  wire n718bar;
  wire n719bar;
  wire n720bar;
  wire n721bar;
  wire n722bar;
  wire n723bar;
  wire n724bar;
  wire n725bar;
  wire n726bar;
  wire n727bar;
  wire n728bar;
  wire n729bar;
  wire n730bar;
  wire n731bar;
  wire n732bar;
  wire n733bar;
  wire n734bar;
  wire n735bar;
  wire n736bar;
  wire n737bar;
  wire n738bar;
  wire n739bar;
  wire n740bar;
  wire n741bar;
  wire n742bar;
  wire n743bar;
  wire n744bar;
  wire n745bar;
  wire n746bar;
  wire n747bar;
  wire n748bar;
  wire n749bar;
  wire n750bar;
  wire n751bar;
  wire n752bar;
  wire n753bar;
  wire n754bar;
  wire n755bar;
  wire n756bar;
  wire n757bar;
  wire n758bar;
  wire n759bar;
  wire n760bar;
  wire n761bar;
  wire n762bar;
  wire n763bar;
  wire n764bar;
  wire n765bar;
  wire n766bar;
  wire n767bar;
  wire n768bar;
  wire n769bar;
  wire n770bar;
  wire n771bar;
  wire n772bar;
  wire n773bar;
  wire n774bar;
  wire n775bar;
  wire n776bar;
  wire n777bar;
  wire n778bar;
  wire n779bar;
  wire n780bar;
  wire n781bar;
  wire n782bar;
  wire n783bar;
  wire n784bar;
  wire n785bar;
  wire n786bar;
  wire n787bar;
  wire n788bar;
  wire n789bar;
  wire n790bar;
  wire n791bar;
  wire n792bar;
  wire n793bar;
  wire n794bar;
  wire n795bar;
  wire n796bar;
  wire n797bar;
  wire n798bar;
  wire n799bar;
  wire n800bar;
  wire n801bar;
  wire n802bar;
  wire n803bar;
  wire n804bar;
  wire n805bar;
  wire n806bar;
  wire n807bar;
  wire n808bar;
  wire n809bar;
  wire n810bar;
  wire n811bar;
  wire n812bar;
  wire n813bar;
  wire n814bar;
  wire n815bar;
  wire n816bar;
  wire n817bar;
  wire n818bar;
  wire n819bar;
  wire n820bar;
  wire n821bar;
  wire n822bar;
  wire n823bar;
  wire n824bar;
  wire n825bar;
  wire n826bar;
  wire n827bar;
  wire n828bar;
  wire n829bar;
  wire n830bar;
  wire n831bar;
  wire n832bar;
  wire n833bar;
  wire n834bar;
  wire n835bar;
  wire n836bar;
  wire n837bar;
  wire n838bar;
  wire n839bar;
  wire n840bar;
  wire n841bar;
  wire n842bar;
  wire n843bar;
  wire n844bar;
  wire n845bar;
  wire n846bar;
  wire n847bar;
  wire n848bar;
  wire n849bar;
  wire n850bar;
  wire n851bar;
  wire n852bar;
  wire n853bar;
  wire n854bar;
  wire n855bar;
  wire n856bar;
  wire n857bar;
  wire n858bar;
  wire n859bar;
  wire n860bar;
  wire n861bar;
  wire n862bar;
  wire n863bar;
  wire n864bar;
  wire n865bar;
  wire n866bar;
  wire n867bar;
  wire n868bar;
  wire n869bar;
  wire n870bar;
  wire n871bar;
  wire n872bar;
  wire n873bar;
  wire n874bar;
  wire n875bar;
  wire n876bar;
  wire n877bar;
  wire n878bar;
  wire n879bar;
  wire n880bar;
  wire n881bar;
  wire n882bar;
  wire n883bar;
  wire n884bar;
  wire n885bar;
  wire n886bar;
  wire n887bar;
  wire n888bar;
  wire n889bar;
  wire n890bar;
  wire n891bar;
  wire n892bar;
  wire n893bar;
  wire n894bar;
  wire n895bar;
  wire n896bar;
  wire n897bar;
  wire n898bar;
  wire n899bar;
  wire n900bar;
  wire n901bar;
  wire n902bar;
  wire n903bar;
  wire n904bar;
  wire n905bar;
  wire n906bar;
  wire n907bar;
  wire n908bar;
  wire n909bar;
  wire n910bar;
  wire n911bar;
  wire n912bar;
  wire n913bar;
  wire n914bar;
  wire n915bar;
  wire n916bar;
  wire n917bar;
  wire n918bar;
  wire n919bar;
  wire n920bar;
  wire n921bar;
  wire n922bar;
  wire n923bar;
  wire n924bar;
  wire n925bar;
  wire n926bar;
  wire n927bar;
  wire n928bar;
  wire n929bar;
  wire n930bar;
  wire n931bar;
  wire n932bar;
  wire n933bar;
  wire n934bar;
  wire n935bar;
  wire n936bar;
  wire n937bar;
  wire n938bar;
  wire n939bar;
  wire n940bar;
  wire n941bar;
  wire n942bar;
  wire n943bar;
  wire n944bar;
  wire n945bar;
  wire n946bar;
  wire n947bar;
  wire n948bar;
  wire n949bar;
  wire n950bar;
  wire n951bar;
  wire n952bar;
  wire n953bar;
  wire n954bar;
  wire n955bar;
  wire n956bar;
  wire n957bar;
  wire n958bar;
  wire n959bar;
  wire n960bar;
  wire n961bar;
  wire n962bar;
  wire n963bar;
  wire n964bar;
  wire n965bar;
  wire n966bar;
  wire n967bar;
  wire n968bar;
  wire n969bar;
  wire n970bar;
  wire n971bar;
  wire n972bar;
//wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];
  assign in_81bar = inbar[81];
  assign in_80bar = inbar[80];
  assign in_79bar = inbar[79];
  assign in_78bar = inbar[78];
  assign in_77bar = inbar[77];
  assign in_76bar = inbar[76];
  assign in_75bar = inbar[75];
  assign in_74bar = inbar[74];
  assign in_73bar = inbar[73];
  assign in_72bar = inbar[72];
  assign in_71bar = inbar[71];
  assign in_70bar = inbar[70];
  assign in_69bar = inbar[69];
  assign in_68bar = inbar[68];
  assign in_67bar = inbar[67];
  assign in_66bar = inbar[66];
  assign in_65bar = inbar[65];
  assign in_64bar = inbar[64];
  assign in_63bar = inbar[63];
  assign in_62bar = inbar[62];
  assign in_61bar = inbar[61];
  assign in_60bar = inbar[60];
  assign in_59bar = inbar[59];
  assign in_58bar = inbar[58];
  assign in_57bar = inbar[57];
  assign in_56bar = inbar[56];
  assign in_55bar = inbar[55];
  assign in_54bar = inbar[54];
  assign in_53bar = inbar[53];
  assign in_52bar = inbar[52];
  assign in_51bar = inbar[51];
  assign in_50bar = inbar[50];
  assign in_49bar = inbar[49];
  assign in_48bar = inbar[48];
  assign in_47bar = inbar[47];
  assign in_46bar = inbar[46];
  assign in_45bar = inbar[45];
  assign in_44bar = inbar[44];
  assign in_43bar = inbar[43];
  assign in_42bar = inbar[42];
  assign in_41bar = inbar[41];
  assign in_40bar = inbar[40];
  assign in_39bar = inbar[39];
  assign in_38bar = inbar[38];
  assign in_37bar = inbar[37];
  assign in_36bar = inbar[36];
  assign in_35bar = inbar[35];
  assign in_34bar = inbar[34];
  assign in_33bar = inbar[33];
  assign in_32bar = inbar[32];
  assign in_31bar = inbar[31];
  assign in_30bar = inbar[30];
  assign in_29bar = inbar[29];
  assign in_28bar = inbar[28];
  assign in_27bar = inbar[27];
  assign in_26bar = inbar[26];
  assign in_25bar = inbar[25];
  assign in_24bar = inbar[24];
  assign in_23bar = inbar[23];
  assign in_22bar = inbar[22];
  assign in_21bar = inbar[21];
  assign in_20bar = inbar[20];
  assign in_19bar = inbar[19];
  assign in_18bar = inbar[18];
  assign in_17bar = inbar[17];
  assign in_16bar = inbar[16];
  assign in_15bar = inbar[15];
  assign in_14bar = inbar[14];
  assign in_13bar = inbar[13];
  assign in_12bar = inbar[12];
  assign in_11bar = inbar[11];
  assign in_10bar = inbar[10];
  assign in_9bar = inbar[9];
  assign in_8bar = inbar[8];
  assign in_7bar = inbar[7];
  assign in_6bar = inbar[6];
  assign in_5bar = inbar[5];
  assign in_4bar = inbar[4];
  assign in_3bar = inbar[3];
  assign in_2bar = inbar[2];
  assign in_1bar = inbar[1];
  assign in_0bar = inbar[0];
//assign_done

  OR2_X1 U1 ( .A1(n972), .A2(n971), .ZN(out[7]) );
  AND2_X1 U1bar ( .A1(n972bar), .A2(n971bar), .ZN(outbar[7]) );
  OR2_X1 U2 ( .A1(n970), .A2(n969), .ZN(n971) );
  AND2_X1 U2bar ( .A1(n970bar), .A2(n969bar), .ZN(n971bar) );
  OR2_X1 U3 ( .A1(n968), .A2(n967), .ZN(n969) );
  AND2_X1 U3bar ( .A1(n968bar), .A2(n967bar), .ZN(n969bar) );
  OR2_X1 U4 ( .A1(n966), .A2(n965), .ZN(n967) );
  AND2_X1 U4bar ( .A1(n966bar), .A2(n965bar), .ZN(n967bar) );
  OR2_X1 U5 ( .A1(n964), .A2(n963), .ZN(n968) );
  AND2_X1 U5bar ( .A1(n964bar), .A2(n963bar), .ZN(n968bar) );
  OR2_X1 U6 ( .A1(in[116]), .A2(n962), .ZN(n963) );
  AND2_X1 U6bar ( .A1(inbar[116]), .A2(n962bar), .ZN(n963bar) );
  OR2_X1 U7 ( .A1(n961), .A2(n960), .ZN(n970) );
  AND2_X1 U7bar ( .A1(n961bar), .A2(n960bar), .ZN(n970bar) );
  OR2_X1 U8 ( .A1(in[150]), .A2(in[127]), .ZN(n960) );
  AND2_X1 U8bar ( .A1(inbar[150]), .A2(inbar[127]), .ZN(n960bar) );
  OR2_X1 U9 ( .A1(in[160]), .A2(n959), .ZN(n961) );
  AND2_X1 U9bar ( .A1(inbar[160]), .A2(n959bar), .ZN(n961bar) );
  OR2_X1 U10 ( .A1(in[252]), .A2(in[168]), .ZN(n959) );
  AND2_X1 U10bar ( .A1(inbar[252]), .A2(inbar[168]), .ZN(n959bar) );
  OR2_X1 U11 ( .A1(n958), .A2(n957), .ZN(n972) );
  AND2_X1 U11bar ( .A1(n958bar), .A2(n957bar), .ZN(n972bar) );
  OR2_X1 U12 ( .A1(n956), .A2(n955), .ZN(n957) );
  AND2_X1 U12bar ( .A1(n956bar), .A2(n955bar), .ZN(n957bar) );
  OR2_X1 U13 ( .A1(in_17), .A2(in[96]), .ZN(n955) );
  AND2_X1 U13bar ( .A1(in_17bar), .A2(inbar[96]), .ZN(n955bar) );
  OR2_X1 U14 ( .A1(in_23), .A2(n954), .ZN(n956) );
  AND2_X1 U14bar ( .A1(in_23bar), .A2(n954bar), .ZN(n956bar) );
  OR2_X1 U15 ( .A1(in_31), .A2(in_26), .ZN(n954) );
  AND2_X1 U15bar ( .A1(in_31bar), .A2(in_26bar), .ZN(n954bar) );
  OR2_X1 U16 ( .A1(n953), .A2(n952), .ZN(n958) );
  AND2_X1 U16bar ( .A1(n953bar), .A2(n952bar), .ZN(n958bar) );
  OR2_X1 U17 ( .A1(in_58), .A2(in_4), .ZN(n952) );
  AND2_X1 U17bar ( .A1(in_58bar), .A2(in_4bar), .ZN(n952bar) );
  OR2_X1 U18 ( .A1(in_59), .A2(n951), .ZN(n953) );
  AND2_X1 U18bar ( .A1(in_59bar), .A2(n951bar), .ZN(n953bar) );
  OR2_X1 U19 ( .A1(in_71), .A2(in_62), .ZN(n951) );
  AND2_X1 U19bar ( .A1(in_71bar), .A2(in_62bar), .ZN(n951bar) );
  OR2_X1 U20 ( .A1(n950), .A2(n949), .ZN(out[6]) );
  AND2_X1 U20bar ( .A1(n950bar), .A2(n949bar), .ZN(outbar[6]) );
  OR2_X1 U21 ( .A1(n948), .A2(n947), .ZN(n949) );
  AND2_X1 U21bar ( .A1(n948bar), .A2(n947bar), .ZN(n949bar) );
  OR2_X1 U22 ( .A1(n946), .A2(n945), .ZN(n947) );
  AND2_X1 U22bar ( .A1(n946bar), .A2(n945bar), .ZN(n947bar) );
  OR2_X1 U23 ( .A1(n944), .A2(n943), .ZN(n945) );
  AND2_X1 U23bar ( .A1(n944bar), .A2(n943bar), .ZN(n945bar) );
  OR2_X1 U24 ( .A1(n942), .A2(n941), .ZN(n946) );
  AND2_X1 U24bar ( .A1(n942bar), .A2(n941bar), .ZN(n946bar) );
  OR2_X1 U25 ( .A1(in[101]), .A2(n940), .ZN(n941) );
  AND2_X1 U25bar ( .A1(inbar[101]), .A2(n940bar), .ZN(n941bar) );
  OR2_X1 U26 ( .A1(n939), .A2(n938), .ZN(n948) );
  AND2_X1 U26bar ( .A1(n939bar), .A2(n938bar), .ZN(n948bar) );
  OR2_X1 U27 ( .A1(in[114]), .A2(in[104]), .ZN(n938) );
  AND2_X1 U27bar ( .A1(inbar[114]), .A2(inbar[104]), .ZN(n938bar) );
  OR2_X1 U28 ( .A1(in[128]), .A2(n937), .ZN(n939) );
  AND2_X1 U28bar ( .A1(inbar[128]), .A2(n937bar), .ZN(n939bar) );
  OR2_X1 U29 ( .A1(in[136]), .A2(in[134]), .ZN(n937) );
  AND2_X1 U29bar ( .A1(inbar[136]), .A2(inbar[134]), .ZN(n937bar) );
  OR2_X1 U30 ( .A1(n936), .A2(n935), .ZN(n950) );
  AND2_X1 U30bar ( .A1(n936bar), .A2(n935bar), .ZN(n950bar) );
  OR2_X1 U31 ( .A1(n934), .A2(n933), .ZN(n935) );
  AND2_X1 U31bar ( .A1(n934bar), .A2(n933bar), .ZN(n935bar) );
  OR2_X1 U32 ( .A1(in[177]), .A2(in[164]), .ZN(n933) );
  AND2_X1 U32bar ( .A1(inbar[177]), .A2(inbar[164]), .ZN(n933bar) );
  OR2_X1 U33 ( .A1(in[212]), .A2(n932), .ZN(n934) );
  AND2_X1 U33bar ( .A1(inbar[212]), .A2(n932bar), .ZN(n934bar) );
  OR2_X1 U34 ( .A1(in[248]), .A2(in[221]), .ZN(n932) );
  AND2_X1 U34bar ( .A1(inbar[248]), .A2(inbar[221]), .ZN(n932bar) );
  OR2_X1 U35 ( .A1(n931), .A2(n930), .ZN(n936) );
  AND2_X1 U35bar ( .A1(n931bar), .A2(n930bar), .ZN(n936bar) );
  OR2_X1 U36 ( .A1(in_18), .A2(in[93]), .ZN(n930) );
  AND2_X1 U36bar ( .A1(in_18bar), .A2(inbar[93]), .ZN(n930bar) );
  OR2_X1 U37 ( .A1(in_31), .A2(n929), .ZN(n931) );
  AND2_X1 U37bar ( .A1(in_31bar), .A2(n929bar), .ZN(n931bar) );
  OR2_X1 U38 ( .A1(in_7), .A2(in_39), .ZN(n929) );
  AND2_X1 U38bar ( .A1(in_7bar), .A2(in_39bar), .ZN(n929bar) );
  OR2_X1 U39 ( .A1(n928), .A2(n927), .ZN(out[5]) );
  AND2_X1 U39bar ( .A1(n928bar), .A2(n927bar), .ZN(outbar[5]) );
  OR2_X1 U40 ( .A1(n926), .A2(n925), .ZN(n927) );
  AND2_X1 U40bar ( .A1(n926bar), .A2(n925bar), .ZN(n927bar) );
  OR2_X1 U41 ( .A1(n924), .A2(n923), .ZN(n925) );
  AND2_X1 U41bar ( .A1(n924bar), .A2(n923bar), .ZN(n925bar) );
  OR2_X1 U42 ( .A1(n922), .A2(n921), .ZN(n923) );
  AND2_X1 U42bar ( .A1(n922bar), .A2(n921bar), .ZN(n923bar) );
  OR2_X1 U43 ( .A1(n940), .A2(n920), .ZN(n924) );
  AND2_X1 U43bar ( .A1(n940bar), .A2(n920bar), .ZN(n924bar) );
  OR2_X1 U44 ( .A1(in[111]), .A2(n919), .ZN(n920) );
  AND2_X1 U44bar ( .A1(inbar[111]), .A2(n919bar), .ZN(n920bar) );
  OR2_X1 U45 ( .A1(n918), .A2(n917), .ZN(n940) );
  AND2_X1 U45bar ( .A1(n918bar), .A2(n917bar), .ZN(n940bar) );
  OR2_X1 U46 ( .A1(n916), .A2(n915), .ZN(n917) );
  AND2_X1 U46bar ( .A1(n916bar), .A2(n915bar), .ZN(n917bar) );
  OR2_X1 U47 ( .A1(n914), .A2(n913), .ZN(n915) );
  AND2_X1 U47bar ( .A1(n914bar), .A2(n913bar), .ZN(n915bar) );
  OR2_X1 U48 ( .A1(in[140]), .A2(in[131]), .ZN(n913) );
  AND2_X1 U48bar ( .A1(inbar[140]), .A2(inbar[131]), .ZN(n913bar) );
  OR2_X1 U49 ( .A1(in[160]), .A2(in[144]), .ZN(n914) );
  AND2_X1 U49bar ( .A1(inbar[160]), .A2(inbar[144]), .ZN(n914bar) );
  OR2_X1 U50 ( .A1(n912), .A2(n911), .ZN(n916) );
  AND2_X1 U50bar ( .A1(n912bar), .A2(n911bar), .ZN(n916bar) );
  OR2_X1 U51 ( .A1(in[179]), .A2(in[174]), .ZN(n911) );
  AND2_X1 U51bar ( .A1(inbar[179]), .A2(inbar[174]), .ZN(n911bar) );
  OR2_X1 U52 ( .A1(in[188]), .A2(in[184]), .ZN(n912) );
  AND2_X1 U52bar ( .A1(inbar[188]), .A2(inbar[184]), .ZN(n912bar) );
  OR2_X1 U53 ( .A1(n910), .A2(n909), .ZN(n918) );
  AND2_X1 U53bar ( .A1(n910bar), .A2(n909bar), .ZN(n918bar) );
  OR2_X1 U54 ( .A1(n908), .A2(n907), .ZN(n909) );
  AND2_X1 U54bar ( .A1(n908bar), .A2(n907bar), .ZN(n909bar) );
  OR2_X1 U55 ( .A1(in[216]), .A2(in[200]), .ZN(n907) );
  AND2_X1 U55bar ( .A1(inbar[216]), .A2(inbar[200]), .ZN(n907bar) );
  OR2_X1 U56 ( .A1(in[228]), .A2(in[224]), .ZN(n908) );
  AND2_X1 U56bar ( .A1(inbar[228]), .A2(inbar[224]), .ZN(n908bar) );
  OR2_X1 U57 ( .A1(n906), .A2(n905), .ZN(n910) );
  AND2_X1 U57bar ( .A1(n906bar), .A2(n905bar), .ZN(n910bar) );
  OR2_X1 U58 ( .A1(in[247]), .A2(in[235]), .ZN(n905) );
  AND2_X1 U58bar ( .A1(inbar[247]), .A2(inbar[235]), .ZN(n905bar) );
  OR2_X1 U59 ( .A1(in_42), .A2(in[83]), .ZN(n906) );
  AND2_X1 U59bar ( .A1(in_42bar), .A2(inbar[83]), .ZN(n906bar) );
  OR2_X1 U60 ( .A1(n904), .A2(n903), .ZN(n926) );
  AND2_X1 U60bar ( .A1(n904bar), .A2(n903bar), .ZN(n926bar) );
  OR2_X1 U61 ( .A1(in[166]), .A2(in[123]), .ZN(n903) );
  AND2_X1 U61bar ( .A1(inbar[166]), .A2(inbar[123]), .ZN(n903bar) );
  OR2_X1 U62 ( .A1(in[170]), .A2(n902), .ZN(n904) );
  AND2_X1 U62bar ( .A1(inbar[170]), .A2(n902bar), .ZN(n904bar) );
  OR2_X1 U63 ( .A1(in[194]), .A2(in[183]), .ZN(n902) );
  AND2_X1 U63bar ( .A1(inbar[194]), .A2(inbar[183]), .ZN(n902bar) );
  OR2_X1 U64 ( .A1(n901), .A2(n900), .ZN(n928) );
  AND2_X1 U64bar ( .A1(n901bar), .A2(n900bar), .ZN(n928bar) );
  OR2_X1 U65 ( .A1(n899), .A2(n898), .ZN(n900) );
  AND2_X1 U65bar ( .A1(n899bar), .A2(n898bar), .ZN(n900bar) );
  OR2_X1 U66 ( .A1(in[241]), .A2(in[238]), .ZN(n898) );
  AND2_X1 U66bar ( .A1(inbar[241]), .A2(inbar[238]), .ZN(n898bar) );
  OR2_X1 U67 ( .A1(in[250]), .A2(n897), .ZN(n899) );
  AND2_X1 U67bar ( .A1(inbar[250]), .A2(n897bar), .ZN(n899bar) );
  OR2_X1 U68 ( .A1(in_24), .A2(in[84]), .ZN(n897) );
  AND2_X1 U68bar ( .A1(in_24bar), .A2(inbar[84]), .ZN(n897bar) );
  OR2_X1 U69 ( .A1(n896), .A2(n895), .ZN(n901) );
  AND2_X1 U69bar ( .A1(n896bar), .A2(n895bar), .ZN(n901bar) );
  OR2_X1 U70 ( .A1(in_41), .A2(in_29), .ZN(n895) );
  AND2_X1 U70bar ( .A1(in_41bar), .A2(in_29bar), .ZN(n895bar) );
  OR2_X1 U71 ( .A1(in_66), .A2(n894), .ZN(n896) );
  AND2_X1 U71bar ( .A1(in_66bar), .A2(n894bar), .ZN(n896bar) );
  OR2_X1 U72 ( .A1(in_76), .A2(in_71), .ZN(n894) );
  AND2_X1 U72bar ( .A1(in_76bar), .A2(in_71bar), .ZN(n894bar) );
  OR2_X1 U73 ( .A1(n893), .A2(n892), .ZN(out[4]) );
  AND2_X1 U73bar ( .A1(n893bar), .A2(n892bar), .ZN(outbar[4]) );
  OR2_X1 U74 ( .A1(n891), .A2(n890), .ZN(n892) );
  AND2_X1 U74bar ( .A1(n891bar), .A2(n890bar), .ZN(n892bar) );
  OR2_X1 U75 ( .A1(n889), .A2(n888), .ZN(n890) );
  AND2_X1 U75bar ( .A1(n889bar), .A2(n888bar), .ZN(n890bar) );
  OR2_X1 U76 ( .A1(n922), .A2(n887), .ZN(n888) );
  AND2_X1 U76bar ( .A1(n922bar), .A2(n887bar), .ZN(n888bar) );
  OR2_X1 U77 ( .A1(n886), .A2(n885), .ZN(n922) );
  AND2_X1 U77bar ( .A1(n886bar), .A2(n885bar), .ZN(n922bar) );
  OR2_X1 U78 ( .A1(n884), .A2(n883), .ZN(n885) );
  AND2_X1 U78bar ( .A1(n884bar), .A2(n883bar), .ZN(n885bar) );
  OR2_X1 U79 ( .A1(n882), .A2(n881), .ZN(n883) );
  AND2_X1 U79bar ( .A1(n882bar), .A2(n881bar), .ZN(n883bar) );
  OR2_X1 U80 ( .A1(in[118]), .A2(in[109]), .ZN(n881) );
  AND2_X1 U80bar ( .A1(inbar[118]), .A2(inbar[109]), .ZN(n881bar) );
  OR2_X1 U81 ( .A1(in[139]), .A2(in[120]), .ZN(n882) );
  AND2_X1 U81bar ( .A1(inbar[139]), .A2(inbar[120]), .ZN(n882bar) );
  OR2_X1 U82 ( .A1(n880), .A2(n879), .ZN(n884) );
  AND2_X1 U82bar ( .A1(n880bar), .A2(n879bar), .ZN(n884bar) );
  OR2_X1 U83 ( .A1(in[198]), .A2(in[154]), .ZN(n879) );
  AND2_X1 U83bar ( .A1(inbar[198]), .A2(inbar[154]), .ZN(n879bar) );
  OR2_X1 U84 ( .A1(in[210]), .A2(in[205]), .ZN(n880) );
  AND2_X1 U84bar ( .A1(inbar[210]), .A2(inbar[205]), .ZN(n880bar) );
  OR2_X1 U85 ( .A1(n878), .A2(n877), .ZN(n886) );
  AND2_X1 U85bar ( .A1(n878bar), .A2(n877bar), .ZN(n886bar) );
  OR2_X1 U86 ( .A1(n876), .A2(n875), .ZN(n877) );
  AND2_X1 U86bar ( .A1(n876bar), .A2(n875bar), .ZN(n877bar) );
  OR2_X1 U87 ( .A1(in[219]), .A2(in[217]), .ZN(n875) );
  AND2_X1 U87bar ( .A1(inbar[219]), .A2(inbar[217]), .ZN(n875bar) );
  OR2_X1 U88 ( .A1(in[86]), .A2(in[252]), .ZN(n876) );
  AND2_X1 U88bar ( .A1(inbar[86]), .A2(inbar[252]), .ZN(n876bar) );
  OR2_X1 U89 ( .A1(n874), .A2(n873), .ZN(n878) );
  AND2_X1 U89bar ( .A1(n874bar), .A2(n873bar), .ZN(n878bar) );
  OR2_X1 U90 ( .A1(in_40), .A2(in[91]), .ZN(n873) );
  AND2_X1 U90bar ( .A1(in_40bar), .A2(inbar[91]), .ZN(n873bar) );
  OR2_X1 U91 ( .A1(in_8), .A2(in_46), .ZN(n874) );
  AND2_X1 U91bar ( .A1(in_8bar), .A2(in_46bar), .ZN(n874bar) );
  OR2_X1 U92 ( .A1(n872), .A2(n871), .ZN(n889) );
  AND2_X1 U92bar ( .A1(n872bar), .A2(n871bar), .ZN(n889bar) );
  OR2_X1 U93 ( .A1(in[117]), .A2(n943), .ZN(n871) );
  AND2_X1 U93bar ( .A1(inbar[117]), .A2(n943bar), .ZN(n871bar) );
  OR2_X1 U94 ( .A1(n870), .A2(n869), .ZN(n943) );
  AND2_X1 U94bar ( .A1(n870bar), .A2(n869bar), .ZN(n943bar) );
  OR2_X1 U95 ( .A1(n868), .A2(n867), .ZN(n869) );
  AND2_X1 U95bar ( .A1(n868bar), .A2(n867bar), .ZN(n869bar) );
  OR2_X1 U96 ( .A1(n866), .A2(n865), .ZN(n867) );
  AND2_X1 U96bar ( .A1(n866bar), .A2(n865bar), .ZN(n867bar) );
  OR2_X1 U97 ( .A1(n864), .A2(n863), .ZN(n865) );
  AND2_X1 U97bar ( .A1(n864bar), .A2(n863bar), .ZN(n865bar) );
  OR2_X1 U98 ( .A1(in[108]), .A2(n919), .ZN(n866) );
  AND2_X1 U98bar ( .A1(inbar[108]), .A2(n919bar), .ZN(n866bar) );
  OR2_X1 U99 ( .A1(n862), .A2(n861), .ZN(n919) );
  AND2_X1 U99bar ( .A1(n862bar), .A2(n861bar), .ZN(n919bar) );
  OR2_X1 U100 ( .A1(n860), .A2(n859), .ZN(n861) );
  AND2_X1 U100bar ( .A1(n860bar), .A2(n859bar), .ZN(n861bar) );
  OR2_X1 U101 ( .A1(n858), .A2(n857), .ZN(n859) );
  AND2_X1 U101bar ( .A1(n858bar), .A2(n857bar), .ZN(n859bar) );
  OR2_X1 U102 ( .A1(in[119]), .A2(in[105]), .ZN(n857) );
  AND2_X1 U102bar ( .A1(inbar[119]), .A2(inbar[105]), .ZN(n857bar) );
  OR2_X1 U103 ( .A1(in[186]), .A2(in[175]), .ZN(n858) );
  AND2_X1 U103bar ( .A1(inbar[186]), .A2(inbar[175]), .ZN(n858bar) );
  OR2_X1 U104 ( .A1(n856), .A2(n855), .ZN(n860) );
  AND2_X1 U104bar ( .A1(n856bar), .A2(n855bar), .ZN(n860bar) );
  OR2_X1 U105 ( .A1(in[202]), .A2(in[193]), .ZN(n855) );
  AND2_X1 U105bar ( .A1(inbar[202]), .A2(inbar[193]), .ZN(n855bar) );
  OR2_X1 U106 ( .A1(in[225]), .A2(in[208]), .ZN(n856) );
  AND2_X1 U106bar ( .A1(inbar[225]), .A2(inbar[208]), .ZN(n856bar) );
  OR2_X1 U107 ( .A1(n854), .A2(n853), .ZN(n862) );
  AND2_X1 U107bar ( .A1(n854bar), .A2(n853bar), .ZN(n862bar) );
  OR2_X1 U108 ( .A1(n852), .A2(n851), .ZN(n853) );
  AND2_X1 U108bar ( .A1(n852bar), .A2(n851bar), .ZN(n853bar) );
  OR2_X1 U109 ( .A1(in_1), .A2(in[85]), .ZN(n851) );
  AND2_X1 U109bar ( .A1(in_1bar), .A2(inbar[85]), .ZN(n851bar) );
  OR2_X1 U110 ( .A1(in_23), .A2(in_19), .ZN(n852) );
  AND2_X1 U110bar ( .A1(in_23bar), .A2(in_19bar), .ZN(n852bar) );
  OR2_X1 U111 ( .A1(n850), .A2(n849), .ZN(n854) );
  AND2_X1 U111bar ( .A1(n850bar), .A2(n849bar), .ZN(n854bar) );
  OR2_X1 U112 ( .A1(in_43), .A2(in_33), .ZN(n849) );
  AND2_X1 U112bar ( .A1(in_43bar), .A2(in_33bar), .ZN(n849bar) );
  OR2_X1 U113 ( .A1(in_63), .A2(in_44), .ZN(n850) );
  AND2_X1 U113bar ( .A1(in_63bar), .A2(in_44bar), .ZN(n850bar) );
  OR2_X1 U114 ( .A1(n848), .A2(n847), .ZN(n868) );
  AND2_X1 U114bar ( .A1(n848bar), .A2(n847bar), .ZN(n868bar) );
  OR2_X1 U115 ( .A1(in[141]), .A2(in[112]), .ZN(n847) );
  AND2_X1 U115bar ( .A1(inbar[141]), .A2(inbar[112]), .ZN(n847bar) );
  OR2_X1 U116 ( .A1(in[147]), .A2(n846), .ZN(n848) );
  AND2_X1 U116bar ( .A1(inbar[147]), .A2(n846bar), .ZN(n848bar) );
  OR2_X1 U117 ( .A1(in[181]), .A2(in[167]), .ZN(n846) );
  AND2_X1 U117bar ( .A1(inbar[181]), .A2(inbar[167]), .ZN(n846bar) );
  OR2_X1 U118 ( .A1(n845), .A2(n844), .ZN(n870) );
  AND2_X1 U118bar ( .A1(n845bar), .A2(n844bar), .ZN(n870bar) );
  OR2_X1 U119 ( .A1(n843), .A2(n842), .ZN(n844) );
  AND2_X1 U119bar ( .A1(n843bar), .A2(n842bar), .ZN(n844bar) );
  OR2_X1 U120 ( .A1(in[229]), .A2(in[201]), .ZN(n842) );
  AND2_X1 U120bar ( .A1(inbar[229]), .A2(inbar[201]), .ZN(n842bar) );
  OR2_X1 U121 ( .A1(in[237]), .A2(n841), .ZN(n843) );
  AND2_X1 U121bar ( .A1(inbar[237]), .A2(n841bar), .ZN(n843bar) );
  OR2_X1 U122 ( .A1(in[94]), .A2(in[253]), .ZN(n841) );
  AND2_X1 U122bar ( .A1(inbar[94]), .A2(inbar[253]), .ZN(n841bar) );
  OR2_X1 U123 ( .A1(n840), .A2(n839), .ZN(n845) );
  AND2_X1 U123bar ( .A1(n840bar), .A2(n839bar), .ZN(n845bar) );
  OR2_X1 U124 ( .A1(in_21), .A2(in[96]), .ZN(n839) );
  AND2_X1 U124bar ( .A1(in_21bar), .A2(inbar[96]), .ZN(n839bar) );
  OR2_X1 U125 ( .A1(in_25), .A2(n838), .ZN(n840) );
  AND2_X1 U125bar ( .A1(in_25bar), .A2(n838bar), .ZN(n840bar) );
  OR2_X1 U126 ( .A1(in_81), .A2(in_45), .ZN(n838) );
  AND2_X1 U126bar ( .A1(in_81bar), .A2(in_45bar), .ZN(n838bar) );
  OR2_X1 U127 ( .A1(n837), .A2(n836), .ZN(n891) );
  AND2_X1 U127bar ( .A1(n837bar), .A2(n836bar), .ZN(n891bar) );
  OR2_X1 U128 ( .A1(in[142]), .A2(in[124]), .ZN(n836) );
  AND2_X1 U128bar ( .A1(inbar[142]), .A2(inbar[124]), .ZN(n836bar) );
  OR2_X1 U129 ( .A1(in[150]), .A2(n835), .ZN(n837) );
  AND2_X1 U129bar ( .A1(inbar[150]), .A2(n835bar), .ZN(n837bar) );
  OR2_X1 U130 ( .A1(in[172]), .A2(in[155]), .ZN(n835) );
  AND2_X1 U130bar ( .A1(inbar[172]), .A2(inbar[155]), .ZN(n835bar) );
  OR2_X1 U131 ( .A1(n834), .A2(n833), .ZN(n893) );
  AND2_X1 U131bar ( .A1(n834bar), .A2(n833bar), .ZN(n893bar) );
  OR2_X1 U132 ( .A1(n832), .A2(n831), .ZN(n833) );
  AND2_X1 U132bar ( .A1(n832bar), .A2(n831bar), .ZN(n833bar) );
  OR2_X1 U133 ( .A1(in[196]), .A2(in[173]), .ZN(n831) );
  AND2_X1 U133bar ( .A1(inbar[196]), .A2(inbar[173]), .ZN(n831bar) );
  OR2_X1 U134 ( .A1(in[222]), .A2(n830), .ZN(n832) );
  AND2_X1 U134bar ( .A1(inbar[222]), .A2(n830bar), .ZN(n832bar) );
  OR2_X1 U135 ( .A1(in[227]), .A2(in[226]), .ZN(n830) );
  AND2_X1 U135bar ( .A1(inbar[227]), .A2(inbar[226]), .ZN(n830bar) );
  OR2_X1 U136 ( .A1(n829), .A2(n828), .ZN(n834) );
  AND2_X1 U136bar ( .A1(n829bar), .A2(n828bar), .ZN(n834bar) );
  OR2_X1 U137 ( .A1(in[249]), .A2(in[231]), .ZN(n828) );
  AND2_X1 U137bar ( .A1(inbar[249]), .A2(inbar[231]), .ZN(n828bar) );
  OR2_X1 U138 ( .A1(in_28), .A2(n827), .ZN(n829) );
  AND2_X1 U138bar ( .A1(in_28bar), .A2(n827bar), .ZN(n829bar) );
  OR2_X1 U139 ( .A1(in_52), .A2(in_47), .ZN(n827) );
  AND2_X1 U139bar ( .A1(in_52bar), .A2(in_47bar), .ZN(n827bar) );
  OR2_X1 U140 ( .A1(n826), .A2(n825), .ZN(out[3]) );
  AND2_X1 U140bar ( .A1(n826bar), .A2(n825bar), .ZN(outbar[3]) );
  OR2_X1 U141 ( .A1(n824), .A2(n823), .ZN(n825) );
  AND2_X1 U141bar ( .A1(n824bar), .A2(n823bar), .ZN(n825bar) );
  OR2_X1 U142 ( .A1(n822), .A2(n821), .ZN(n823) );
  AND2_X1 U142bar ( .A1(n822bar), .A2(n821bar), .ZN(n823bar) );
  OR2_X1 U143 ( .A1(n820), .A2(n819), .ZN(n821) );
  AND2_X1 U143bar ( .A1(n820bar), .A2(n819bar), .ZN(n821bar) );
  OR2_X1 U144 ( .A1(n964), .A2(n818), .ZN(n822) );
  AND2_X1 U144bar ( .A1(n964bar), .A2(n818bar), .ZN(n822bar) );
  OR2_X1 U145 ( .A1(in[118]), .A2(n817), .ZN(n818) );
  AND2_X1 U145bar ( .A1(inbar[118]), .A2(n817bar), .ZN(n818bar) );
  OR2_X1 U146 ( .A1(n816), .A2(n815), .ZN(n964) );
  AND2_X1 U146bar ( .A1(n816bar), .A2(n815bar), .ZN(n964bar) );
  OR2_X1 U147 ( .A1(n814), .A2(n813), .ZN(n815) );
  AND2_X1 U147bar ( .A1(n814bar), .A2(n813bar), .ZN(n815bar) );
  OR2_X1 U148 ( .A1(n812), .A2(n811), .ZN(n813) );
  AND2_X1 U148bar ( .A1(n812bar), .A2(n811bar), .ZN(n813bar) );
  OR2_X1 U149 ( .A1(in[122]), .A2(in[111]), .ZN(n811) );
  AND2_X1 U149bar ( .A1(inbar[122]), .A2(inbar[111]), .ZN(n811bar) );
  OR2_X1 U150 ( .A1(in[154]), .A2(in[151]), .ZN(n812) );
  AND2_X1 U150bar ( .A1(inbar[154]), .A2(inbar[151]), .ZN(n812bar) );
  OR2_X1 U151 ( .A1(n810), .A2(n809), .ZN(n814) );
  AND2_X1 U151bar ( .A1(n810bar), .A2(n809bar), .ZN(n814bar) );
  OR2_X1 U152 ( .A1(in[187]), .A2(in[177]), .ZN(n809) );
  AND2_X1 U152bar ( .A1(inbar[187]), .A2(inbar[177]), .ZN(n809bar) );
  OR2_X1 U153 ( .A1(in[200]), .A2(in[192]), .ZN(n810) );
  AND2_X1 U153bar ( .A1(inbar[200]), .A2(inbar[192]), .ZN(n810bar) );
  OR2_X1 U154 ( .A1(n808), .A2(n807), .ZN(n816) );
  AND2_X1 U154bar ( .A1(n808bar), .A2(n807bar), .ZN(n816bar) );
  OR2_X1 U155 ( .A1(n806), .A2(n805), .ZN(n807) );
  AND2_X1 U155bar ( .A1(n806bar), .A2(n805bar), .ZN(n807bar) );
  OR2_X1 U156 ( .A1(in[225]), .A2(in[207]), .ZN(n805) );
  AND2_X1 U156bar ( .A1(inbar[225]), .A2(inbar[207]), .ZN(n805bar) );
  OR2_X1 U157 ( .A1(in[98]), .A2(in[226]), .ZN(n806) );
  AND2_X1 U157bar ( .A1(inbar[98]), .A2(inbar[226]), .ZN(n806bar) );
  OR2_X1 U158 ( .A1(n804), .A2(n803), .ZN(n808) );
  AND2_X1 U158bar ( .A1(n804bar), .A2(n803bar), .ZN(n808bar) );
  OR2_X1 U159 ( .A1(in_20), .A2(in_16), .ZN(n803) );
  AND2_X1 U159bar ( .A1(in_20bar), .A2(in_16bar), .ZN(n803bar) );
  OR2_X1 U160 ( .A1(in_55), .A2(in_45), .ZN(n804) );
  AND2_X1 U160bar ( .A1(in_55bar), .A2(in_45bar), .ZN(n804bar) );
  OR2_X1 U161 ( .A1(n802), .A2(n801), .ZN(n824) );
  AND2_X1 U161bar ( .A1(n802bar), .A2(n801bar), .ZN(n824bar) );
  OR2_X1 U162 ( .A1(in[162]), .A2(in[149]), .ZN(n801) );
  AND2_X1 U162bar ( .A1(inbar[162]), .A2(inbar[149]), .ZN(n801bar) );
  OR2_X1 U163 ( .A1(in[163]), .A2(n800), .ZN(n802) );
  AND2_X1 U163bar ( .A1(inbar[163]), .A2(n800bar), .ZN(n802bar) );
  OR2_X1 U164 ( .A1(in[191]), .A2(in[189]), .ZN(n800) );
  AND2_X1 U164bar ( .A1(inbar[191]), .A2(inbar[189]), .ZN(n800bar) );
  OR2_X1 U165 ( .A1(n799), .A2(n798), .ZN(n826) );
  AND2_X1 U165bar ( .A1(n799bar), .A2(n798bar), .ZN(n826bar) );
  OR2_X1 U166 ( .A1(n797), .A2(n796), .ZN(n798) );
  AND2_X1 U166bar ( .A1(n797bar), .A2(n796bar), .ZN(n798bar) );
  OR2_X1 U167 ( .A1(in[212]), .A2(in[193]), .ZN(n796) );
  AND2_X1 U167bar ( .A1(inbar[212]), .A2(inbar[193]), .ZN(n796bar) );
  OR2_X1 U168 ( .A1(in[238]), .A2(n795), .ZN(n797) );
  AND2_X1 U168bar ( .A1(inbar[238]), .A2(n795bar), .ZN(n797bar) );
  OR2_X1 U169 ( .A1(in[88]), .A2(in[247]), .ZN(n795) );
  AND2_X1 U169bar ( .A1(inbar[88]), .A2(inbar[247]), .ZN(n795bar) );
  OR2_X1 U170 ( .A1(n794), .A2(n793), .ZN(n799) );
  AND2_X1 U170bar ( .A1(n794bar), .A2(n793bar), .ZN(n799bar) );
  OR2_X1 U171 ( .A1(in[94]), .A2(in[92]), .ZN(n793) );
  AND2_X1 U171bar ( .A1(inbar[94]), .A2(inbar[92]), .ZN(n793bar) );
  OR2_X1 U172 ( .A1(in_52), .A2(n792), .ZN(n794) );
  AND2_X1 U172bar ( .A1(in_52bar), .A2(n792bar), .ZN(n794bar) );
  OR2_X1 U173 ( .A1(in_70), .A2(in_67), .ZN(n792) );
  AND2_X1 U173bar ( .A1(in_70bar), .A2(in_67bar), .ZN(n792bar) );
  OR2_X1 U174 ( .A1(n791), .A2(n790), .ZN(out[2]) );
  AND2_X1 U174bar ( .A1(n791bar), .A2(n790bar), .ZN(outbar[2]) );
  OR2_X1 U175 ( .A1(n789), .A2(n788), .ZN(n790) );
  AND2_X1 U175bar ( .A1(n789bar), .A2(n788bar), .ZN(n790bar) );
  OR2_X1 U176 ( .A1(n787), .A2(n786), .ZN(n788) );
  AND2_X1 U176bar ( .A1(n787bar), .A2(n786bar), .ZN(n788bar) );
  OR2_X1 U177 ( .A1(n819), .A2(n785), .ZN(n786) );
  AND2_X1 U177bar ( .A1(n819bar), .A2(n785bar), .ZN(n786bar) );
  OR2_X1 U178 ( .A1(n784), .A2(n783), .ZN(n819) );
  AND2_X1 U178bar ( .A1(n784bar), .A2(n783bar), .ZN(n819bar) );
  OR2_X1 U179 ( .A1(n782), .A2(n781), .ZN(n783) );
  AND2_X1 U179bar ( .A1(n782bar), .A2(n781bar), .ZN(n783bar) );
  OR2_X1 U180 ( .A1(n780), .A2(n779), .ZN(n781) );
  AND2_X1 U180bar ( .A1(n780bar), .A2(n779bar), .ZN(n781bar) );
  OR2_X1 U181 ( .A1(n962), .A2(n778), .ZN(n779) );
  AND2_X1 U181bar ( .A1(n962bar), .A2(n778bar), .ZN(n779bar) );
  OR2_X1 U182 ( .A1(n777), .A2(n776), .ZN(n962) );
  AND2_X1 U182bar ( .A1(n777bar), .A2(n776bar), .ZN(n962bar) );
  OR2_X1 U183 ( .A1(n775), .A2(n774), .ZN(n776) );
  AND2_X1 U183bar ( .A1(n775bar), .A2(n774bar), .ZN(n776bar) );
  OR2_X1 U184 ( .A1(n773), .A2(n772), .ZN(n774) );
  AND2_X1 U184bar ( .A1(n773bar), .A2(n772bar), .ZN(n774bar) );
  OR2_X1 U185 ( .A1(in[131]), .A2(in[120]), .ZN(n772) );
  AND2_X1 U185bar ( .A1(inbar[131]), .A2(inbar[120]), .ZN(n772bar) );
  OR2_X1 U186 ( .A1(in[153]), .A2(in[147]), .ZN(n773) );
  AND2_X1 U186bar ( .A1(inbar[153]), .A2(inbar[147]), .ZN(n773bar) );
  OR2_X1 U187 ( .A1(n771), .A2(n770), .ZN(n775) );
  AND2_X1 U187bar ( .A1(n771bar), .A2(n770bar), .ZN(n775bar) );
  OR2_X1 U188 ( .A1(in[170]), .A2(in[156]), .ZN(n770) );
  AND2_X1 U188bar ( .A1(inbar[170]), .A2(inbar[156]), .ZN(n770bar) );
  OR2_X1 U189 ( .A1(in[223]), .A2(in[190]), .ZN(n771) );
  AND2_X1 U189bar ( .A1(inbar[223]), .A2(inbar[190]), .ZN(n771bar) );
  OR2_X1 U190 ( .A1(n769), .A2(n768), .ZN(n777) );
  AND2_X1 U190bar ( .A1(n769bar), .A2(n768bar), .ZN(n777bar) );
  OR2_X1 U191 ( .A1(n767), .A2(n766), .ZN(n768) );
  AND2_X1 U191bar ( .A1(n767bar), .A2(n766bar), .ZN(n768bar) );
  OR2_X1 U192 ( .A1(in[236]), .A2(in[230]), .ZN(n766) );
  AND2_X1 U192bar ( .A1(inbar[236]), .A2(inbar[230]), .ZN(n766bar) );
  OR2_X1 U193 ( .A1(in[85]), .A2(in[240]), .ZN(n767) );
  AND2_X1 U193bar ( .A1(inbar[85]), .A2(inbar[240]), .ZN(n767bar) );
  OR2_X1 U194 ( .A1(n765), .A2(n764), .ZN(n769) );
  AND2_X1 U194bar ( .A1(n765bar), .A2(n764bar), .ZN(n769bar) );
  OR2_X1 U195 ( .A1(in_12), .A2(in[90]), .ZN(n764) );
  AND2_X1 U195bar ( .A1(in_12bar), .A2(inbar[90]), .ZN(n764bar) );
  OR2_X1 U196 ( .A1(in_39), .A2(in_28), .ZN(n765) );
  AND2_X1 U196bar ( .A1(in_39bar), .A2(in_28bar), .ZN(n765bar) );
  OR2_X1 U197 ( .A1(in[109]), .A2(n763), .ZN(n780) );
  AND2_X1 U197bar ( .A1(inbar[109]), .A2(n763bar), .ZN(n780bar) );
  OR2_X1 U198 ( .A1(n762), .A2(n761), .ZN(n782) );
  AND2_X1 U198bar ( .A1(n762bar), .A2(n761bar), .ZN(n782bar) );
  OR2_X1 U199 ( .A1(in[138]), .A2(in[129]), .ZN(n761) );
  AND2_X1 U199bar ( .A1(inbar[138]), .A2(inbar[129]), .ZN(n761bar) );
  OR2_X1 U200 ( .A1(in[157]), .A2(n760), .ZN(n762) );
  AND2_X1 U200bar ( .A1(inbar[157]), .A2(n760bar), .ZN(n762bar) );
  OR2_X1 U201 ( .A1(in[182]), .A2(in[167]), .ZN(n760) );
  AND2_X1 U201bar ( .A1(inbar[182]), .A2(inbar[167]), .ZN(n760bar) );
  OR2_X1 U202 ( .A1(n759), .A2(n758), .ZN(n784) );
  AND2_X1 U202bar ( .A1(n759bar), .A2(n758bar), .ZN(n784bar) );
  OR2_X1 U203 ( .A1(n757), .A2(n756), .ZN(n758) );
  AND2_X1 U203bar ( .A1(n757bar), .A2(n756bar), .ZN(n758bar) );
  OR2_X1 U204 ( .A1(in[195]), .A2(in[184]), .ZN(n756) );
  AND2_X1 U204bar ( .A1(inbar[195]), .A2(inbar[184]), .ZN(n756bar) );
  OR2_X1 U205 ( .A1(in[196]), .A2(n755), .ZN(n757) );
  AND2_X1 U205bar ( .A1(inbar[196]), .A2(n755bar), .ZN(n757bar) );
  OR2_X1 U206 ( .A1(in[215]), .A2(in[209]), .ZN(n755) );
  AND2_X1 U206bar ( .A1(inbar[215]), .A2(inbar[209]), .ZN(n755bar) );
  OR2_X1 U207 ( .A1(n754), .A2(n753), .ZN(n759) );
  AND2_X1 U207bar ( .A1(n754bar), .A2(n753bar), .ZN(n759bar) );
  OR2_X1 U208 ( .A1(in[93]), .A2(in[233]), .ZN(n753) );
  AND2_X1 U208bar ( .A1(inbar[93]), .A2(inbar[233]), .ZN(n753bar) );
  OR2_X1 U209 ( .A1(in_1), .A2(n752), .ZN(n754) );
  AND2_X1 U209bar ( .A1(in_1bar), .A2(n752bar), .ZN(n754bar) );
  OR2_X1 U210 ( .A1(in_69), .A2(in_66), .ZN(n752) );
  AND2_X1 U210bar ( .A1(in_69bar), .A2(in_66bar), .ZN(n752bar) );
  OR2_X1 U211 ( .A1(n966), .A2(n751), .ZN(n787) );
  AND2_X1 U211bar ( .A1(n966bar), .A2(n751bar), .ZN(n787bar) );
  OR2_X1 U212 ( .A1(in[134]), .A2(n750), .ZN(n751) );
  AND2_X1 U212bar ( .A1(inbar[134]), .A2(n750bar), .ZN(n751bar) );
  OR2_X1 U213 ( .A1(n749), .A2(n748), .ZN(n966) );
  AND2_X1 U213bar ( .A1(n749bar), .A2(n748bar), .ZN(n966bar) );
  OR2_X1 U214 ( .A1(n747), .A2(n746), .ZN(n748) );
  AND2_X1 U214bar ( .A1(n747bar), .A2(n746bar), .ZN(n748bar) );
  OR2_X1 U215 ( .A1(n745), .A2(n744), .ZN(n746) );
  AND2_X1 U215bar ( .A1(n745bar), .A2(n744bar), .ZN(n746bar) );
  OR2_X1 U216 ( .A1(in[136]), .A2(in[121]), .ZN(n744) );
  AND2_X1 U216bar ( .A1(inbar[136]), .A2(inbar[121]), .ZN(n744bar) );
  OR2_X1 U217 ( .A1(in[186]), .A2(in[174]), .ZN(n745) );
  AND2_X1 U217bar ( .A1(inbar[186]), .A2(inbar[174]), .ZN(n745bar) );
  OR2_X1 U218 ( .A1(n743), .A2(n742), .ZN(n747) );
  AND2_X1 U218bar ( .A1(n743bar), .A2(n742bar), .ZN(n747bar) );
  OR2_X1 U219 ( .A1(in[198]), .A2(in[197]), .ZN(n742) );
  AND2_X1 U219bar ( .A1(inbar[198]), .A2(inbar[197]), .ZN(n742bar) );
  OR2_X1 U220 ( .A1(in[214]), .A2(in[199]), .ZN(n743) );
  AND2_X1 U220bar ( .A1(inbar[214]), .A2(inbar[199]), .ZN(n743bar) );
  OR2_X1 U221 ( .A1(n741), .A2(n740), .ZN(n749) );
  AND2_X1 U221bar ( .A1(n741bar), .A2(n740bar), .ZN(n749bar) );
  OR2_X1 U222 ( .A1(n739), .A2(n738), .ZN(n740) );
  AND2_X1 U222bar ( .A1(n739bar), .A2(n738bar), .ZN(n740bar) );
  OR2_X1 U223 ( .A1(in[231]), .A2(in[220]), .ZN(n738) );
  AND2_X1 U223bar ( .A1(inbar[231]), .A2(inbar[220]), .ZN(n738bar) );
  OR2_X1 U224 ( .A1(in_25), .A2(in[245]), .ZN(n739) );
  AND2_X1 U224bar ( .A1(in_25bar), .A2(inbar[245]), .ZN(n739bar) );
  OR2_X1 U225 ( .A1(n737), .A2(n736), .ZN(n741) );
  AND2_X1 U225bar ( .A1(n737bar), .A2(n736bar), .ZN(n741bar) );
  OR2_X1 U226 ( .A1(in_53), .A2(in_29), .ZN(n736) );
  AND2_X1 U226bar ( .A1(in_53bar), .A2(in_29bar), .ZN(n736bar) );
  OR2_X1 U227 ( .A1(in_79), .A2(in_74), .ZN(n737) );
  AND2_X1 U227bar ( .A1(in_79bar), .A2(in_74bar), .ZN(n737bar) );
  OR2_X1 U228 ( .A1(n735), .A2(n734), .ZN(n789) );
  AND2_X1 U228bar ( .A1(n735bar), .A2(n734bar), .ZN(n789bar) );
  OR2_X1 U229 ( .A1(in[152]), .A2(in[140]), .ZN(n734) );
  AND2_X1 U229bar ( .A1(inbar[152]), .A2(inbar[140]), .ZN(n734bar) );
  OR2_X1 U230 ( .A1(in[155]), .A2(n733), .ZN(n735) );
  AND2_X1 U230bar ( .A1(inbar[155]), .A2(n733bar), .ZN(n735bar) );
  OR2_X1 U231 ( .A1(in[166]), .A2(in[165]), .ZN(n733) );
  AND2_X1 U231bar ( .A1(inbar[166]), .A2(inbar[165]), .ZN(n733bar) );
  OR2_X1 U232 ( .A1(n732), .A2(n731), .ZN(n791) );
  AND2_X1 U232bar ( .A1(n732bar), .A2(n731bar), .ZN(n791bar) );
  OR2_X1 U233 ( .A1(n730), .A2(n729), .ZN(n731) );
  AND2_X1 U233bar ( .A1(n730bar), .A2(n729bar), .ZN(n731bar) );
  OR2_X1 U234 ( .A1(in[202]), .A2(in[185]), .ZN(n729) );
  AND2_X1 U234bar ( .A1(inbar[202]), .A2(inbar[185]), .ZN(n729bar) );
  OR2_X1 U235 ( .A1(in[211]), .A2(n728), .ZN(n730) );
  AND2_X1 U235bar ( .A1(inbar[211]), .A2(n728bar), .ZN(n730bar) );
  OR2_X1 U236 ( .A1(in[255]), .A2(in[253]), .ZN(n728) );
  AND2_X1 U236bar ( .A1(inbar[255]), .A2(inbar[253]), .ZN(n728bar) );
  OR2_X1 U237 ( .A1(n727), .A2(n726), .ZN(n732) );
  AND2_X1 U237bar ( .A1(n727bar), .A2(n726bar), .ZN(n732bar) );
  OR2_X1 U238 ( .A1(in_35), .A2(in_15), .ZN(n726) );
  AND2_X1 U238bar ( .A1(in_35bar), .A2(in_15bar), .ZN(n726bar) );
  OR2_X1 U239 ( .A1(in_36), .A2(n725), .ZN(n727) );
  AND2_X1 U239bar ( .A1(in_36bar), .A2(n725bar), .ZN(n727bar) );
  OR2_X1 U240 ( .A1(in_48), .A2(in_40), .ZN(n725) );
  AND2_X1 U240bar ( .A1(in_48bar), .A2(in_40bar), .ZN(n725bar) );
  OR2_X1 U241 ( .A1(n724), .A2(n723), .ZN(out[1]) );
  AND2_X1 U241bar ( .A1(n724bar), .A2(n723bar), .ZN(outbar[1]) );
  OR2_X1 U242 ( .A1(n722), .A2(n721), .ZN(n723) );
  AND2_X1 U242bar ( .A1(n722bar), .A2(n721bar), .ZN(n723bar) );
  OR2_X1 U243 ( .A1(n720), .A2(n719), .ZN(n721) );
  AND2_X1 U243bar ( .A1(n720bar), .A2(n719bar), .ZN(n721bar) );
  OR2_X1 U244 ( .A1(n921), .A2(n887), .ZN(n719) );
  AND2_X1 U244bar ( .A1(n921bar), .A2(n887bar), .ZN(n719bar) );
  OR2_X1 U245 ( .A1(n718), .A2(n717), .ZN(n887) );
  AND2_X1 U245bar ( .A1(n718bar), .A2(n717bar), .ZN(n887bar) );
  OR2_X1 U246 ( .A1(n716), .A2(n715), .ZN(n717) );
  AND2_X1 U246bar ( .A1(n716bar), .A2(n715bar), .ZN(n717bar) );
  OR2_X1 U247 ( .A1(n714), .A2(n713), .ZN(n715) );
  AND2_X1 U247bar ( .A1(n714bar), .A2(n713bar), .ZN(n715bar) );
  OR2_X1 U248 ( .A1(in[116]), .A2(in[110]), .ZN(n713) );
  AND2_X1 U248bar ( .A1(inbar[116]), .A2(inbar[110]), .ZN(n713bar) );
  OR2_X1 U249 ( .A1(in[133]), .A2(in[130]), .ZN(n714) );
  AND2_X1 U249bar ( .A1(inbar[133]), .A2(inbar[130]), .ZN(n714bar) );
  OR2_X1 U250 ( .A1(n712), .A2(n711), .ZN(n716) );
  AND2_X1 U250bar ( .A1(n712bar), .A2(n711bar), .ZN(n716bar) );
  OR2_X1 U251 ( .A1(in[203]), .A2(in[135]), .ZN(n711) );
  AND2_X1 U251bar ( .A1(inbar[203]), .A2(inbar[135]), .ZN(n711bar) );
  OR2_X1 U252 ( .A1(in[232]), .A2(in[223]), .ZN(n712) );
  AND2_X1 U252bar ( .A1(inbar[232]), .A2(inbar[223]), .ZN(n712bar) );
  OR2_X1 U253 ( .A1(n710), .A2(n709), .ZN(n718) );
  AND2_X1 U253bar ( .A1(n710bar), .A2(n709bar), .ZN(n718bar) );
  OR2_X1 U254 ( .A1(n708), .A2(n707), .ZN(n709) );
  AND2_X1 U254bar ( .A1(n708bar), .A2(n707bar), .ZN(n709bar) );
  OR2_X1 U255 ( .A1(in[255]), .A2(in[233]), .ZN(n707) );
  AND2_X1 U255bar ( .A1(inbar[255]), .A2(inbar[233]), .ZN(n707bar) );
  OR2_X1 U256 ( .A1(in_53), .A2(in_34), .ZN(n708) );
  AND2_X1 U256bar ( .A1(in_53bar), .A2(in_34bar), .ZN(n708bar) );
  OR2_X1 U257 ( .A1(n706), .A2(n705), .ZN(n710) );
  AND2_X1 U257bar ( .A1(n706bar), .A2(n705bar), .ZN(n710bar) );
  OR2_X1 U258 ( .A1(in_57), .A2(in_55), .ZN(n705) );
  AND2_X1 U258bar ( .A1(in_57bar), .A2(in_55bar), .ZN(n705bar) );
  OR2_X1 U259 ( .A1(in_68), .A2(in_67), .ZN(n706) );
  AND2_X1 U259bar ( .A1(in_68bar), .A2(in_67bar), .ZN(n706bar) );
  OR2_X1 U260 ( .A1(n704), .A2(n703), .ZN(n921) );
  AND2_X1 U260bar ( .A1(n704bar), .A2(n703bar), .ZN(n921bar) );
  OR2_X1 U261 ( .A1(n702), .A2(n701), .ZN(n703) );
  AND2_X1 U261bar ( .A1(n702bar), .A2(n701bar), .ZN(n703bar) );
  OR2_X1 U262 ( .A1(n700), .A2(n699), .ZN(n701) );
  AND2_X1 U262bar ( .A1(n700bar), .A2(n699bar), .ZN(n701bar) );
  OR2_X1 U263 ( .A1(n944), .A2(n872), .ZN(n699) );
  AND2_X1 U263bar ( .A1(n944bar), .A2(n872bar), .ZN(n699bar) );
  OR2_X1 U264 ( .A1(n698), .A2(n697), .ZN(n872) );
  AND2_X1 U264bar ( .A1(n698bar), .A2(n697bar), .ZN(n872bar) );
  OR2_X1 U265 ( .A1(n696), .A2(n695), .ZN(n697) );
  AND2_X1 U265bar ( .A1(n696bar), .A2(n695bar), .ZN(n697bar) );
  OR2_X1 U266 ( .A1(n694), .A2(n693), .ZN(n695) );
  AND2_X1 U266bar ( .A1(n694bar), .A2(n693bar), .ZN(n695bar) );
  OR2_X1 U267 ( .A1(in[121]), .A2(in[102]), .ZN(n693) );
  AND2_X1 U267bar ( .A1(inbar[121]), .A2(inbar[102]), .ZN(n693bar) );
  OR2_X1 U268 ( .A1(in[162]), .A2(in[161]), .ZN(n694) );
  AND2_X1 U268bar ( .A1(inbar[162]), .A2(inbar[161]), .ZN(n694bar) );
  OR2_X1 U269 ( .A1(n692), .A2(n691), .ZN(n696) );
  AND2_X1 U269bar ( .A1(n692bar), .A2(n691bar), .ZN(n696bar) );
  OR2_X1 U270 ( .A1(in[192]), .A2(in[178]), .ZN(n691) );
  AND2_X1 U270bar ( .A1(inbar[192]), .A2(inbar[178]), .ZN(n691bar) );
  OR2_X1 U271 ( .A1(in[244]), .A2(in[209]), .ZN(n692) );
  AND2_X1 U271bar ( .A1(inbar[244]), .A2(inbar[209]), .ZN(n692bar) );
  OR2_X1 U272 ( .A1(n690), .A2(n689), .ZN(n698) );
  AND2_X1 U272bar ( .A1(n690bar), .A2(n689bar), .ZN(n698bar) );
  OR2_X1 U273 ( .A1(n688), .A2(n687), .ZN(n689) );
  AND2_X1 U273bar ( .A1(n688bar), .A2(n687bar), .ZN(n689bar) );
  OR2_X1 U274 ( .A1(in[90]), .A2(in[254]), .ZN(n687) );
  AND2_X1 U274bar ( .A1(inbar[90]), .A2(inbar[254]), .ZN(n687bar) );
  OR2_X1 U275 ( .A1(in_36), .A2(in_32), .ZN(n688) );
  AND2_X1 U275bar ( .A1(in_36bar), .A2(in_32bar), .ZN(n688bar) );
  OR2_X1 U276 ( .A1(n686), .A2(n685), .ZN(n690) );
  AND2_X1 U276bar ( .A1(n686bar), .A2(n685bar), .ZN(n690bar) );
  OR2_X1 U277 ( .A1(in_62), .A2(in_37), .ZN(n685) );
  AND2_X1 U277bar ( .A1(in_62bar), .A2(in_37bar), .ZN(n685bar) );
  OR2_X1 U278 ( .A1(in_75), .A2(in_73), .ZN(n686) );
  AND2_X1 U278bar ( .A1(in_75bar), .A2(in_73bar), .ZN(n686bar) );
  OR2_X1 U279 ( .A1(n684), .A2(n683), .ZN(n944) );
  AND2_X1 U279bar ( .A1(n684bar), .A2(n683bar), .ZN(n944bar) );
  OR2_X1 U280 ( .A1(n682), .A2(n681), .ZN(n683) );
  AND2_X1 U280bar ( .A1(n682bar), .A2(n681bar), .ZN(n683bar) );
  OR2_X1 U281 ( .A1(n680), .A2(n679), .ZN(n681) );
  AND2_X1 U281bar ( .A1(n680bar), .A2(n679bar), .ZN(n681bar) );
  OR2_X1 U282 ( .A1(in[171]), .A2(in[153]), .ZN(n679) );
  AND2_X1 U282bar ( .A1(inbar[171]), .A2(inbar[153]), .ZN(n679bar) );
  OR2_X1 U283 ( .A1(in[187]), .A2(in[176]), .ZN(n680) );
  AND2_X1 U283bar ( .A1(inbar[187]), .A2(inbar[176]), .ZN(n680bar) );
  OR2_X1 U284 ( .A1(n678), .A2(n677), .ZN(n682) );
  AND2_X1 U284bar ( .A1(n678bar), .A2(n677bar), .ZN(n682bar) );
  OR2_X1 U285 ( .A1(in[245]), .A2(in[211]), .ZN(n677) );
  AND2_X1 U285bar ( .A1(inbar[245]), .A2(inbar[211]), .ZN(n677bar) );
  OR2_X1 U286 ( .A1(in[97]), .A2(in[88]), .ZN(n678) );
  AND2_X1 U286bar ( .A1(inbar[97]), .A2(inbar[88]), .ZN(n678bar) );
  OR2_X1 U287 ( .A1(n676), .A2(n675), .ZN(n684) );
  AND2_X1 U287bar ( .A1(n676bar), .A2(n675bar), .ZN(n684bar) );
  OR2_X1 U288 ( .A1(n674), .A2(n673), .ZN(n675) );
  AND2_X1 U288bar ( .A1(n674bar), .A2(n673bar), .ZN(n675bar) );
  OR2_X1 U289 ( .A1(in_10), .A2(in_0), .ZN(n673) );
  AND2_X1 U289bar ( .A1(in_10bar), .A2(in_0bar), .ZN(n673bar) );
  OR2_X1 U290 ( .A1(in_59), .A2(in_5), .ZN(n674) );
  AND2_X1 U290bar ( .A1(in_59bar), .A2(in_5bar), .ZN(n674bar) );
  OR2_X1 U291 ( .A1(n672), .A2(n671), .ZN(n676) );
  AND2_X1 U291bar ( .A1(n672bar), .A2(n671bar), .ZN(n676bar) );
  OR2_X1 U292 ( .A1(in_60), .A2(in_6), .ZN(n671) );
  AND2_X1 U292bar ( .A1(in_60bar), .A2(in_6bar), .ZN(n671bar) );
  OR2_X1 U293 ( .A1(in_77), .A2(in_69), .ZN(n672) );
  AND2_X1 U293bar ( .A1(in_77bar), .A2(in_69bar), .ZN(n672bar) );
  OR2_X1 U294 ( .A1(in[113]), .A2(n864), .ZN(n700) );
  AND2_X1 U294bar ( .A1(inbar[113]), .A2(n864bar), .ZN(n700bar) );
  OR2_X1 U295 ( .A1(n670), .A2(n669), .ZN(n864) );
  AND2_X1 U295bar ( .A1(n670bar), .A2(n669bar), .ZN(n864bar) );
  OR2_X1 U296 ( .A1(n668), .A2(n667), .ZN(n669) );
  AND2_X1 U296bar ( .A1(n668bar), .A2(n667bar), .ZN(n669bar) );
  OR2_X1 U297 ( .A1(n666), .A2(n665), .ZN(n667) );
  AND2_X1 U297bar ( .A1(n666bar), .A2(n665bar), .ZN(n667bar) );
  OR2_X1 U298 ( .A1(in[125]), .A2(in[107]), .ZN(n665) );
  AND2_X1 U298bar ( .A1(inbar[125]), .A2(inbar[107]), .ZN(n665bar) );
  OR2_X1 U299 ( .A1(in[138]), .A2(in[126]), .ZN(n666) );
  AND2_X1 U299bar ( .A1(inbar[138]), .A2(inbar[126]), .ZN(n666bar) );
  OR2_X1 U300 ( .A1(n664), .A2(n663), .ZN(n668) );
  AND2_X1 U300bar ( .A1(n664bar), .A2(n663bar), .ZN(n668bar) );
  OR2_X1 U301 ( .A1(in[189]), .A2(in[143]), .ZN(n663) );
  AND2_X1 U301bar ( .A1(inbar[189]), .A2(inbar[143]), .ZN(n663bar) );
  OR2_X1 U302 ( .A1(in[99]), .A2(in[214]), .ZN(n664) );
  AND2_X1 U302bar ( .A1(inbar[99]), .A2(inbar[214]), .ZN(n664bar) );
  OR2_X1 U303 ( .A1(n662), .A2(n661), .ZN(n670) );
  AND2_X1 U303bar ( .A1(n662bar), .A2(n661bar), .ZN(n670bar) );
  OR2_X1 U304 ( .A1(n660), .A2(n659), .ZN(n661) );
  AND2_X1 U304bar ( .A1(n660bar), .A2(n659bar), .ZN(n661bar) );
  OR2_X1 U305 ( .A1(in_15), .A2(in_12), .ZN(n659) );
  AND2_X1 U305bar ( .A1(in_15bar), .A2(in_12bar), .ZN(n659bar) );
  OR2_X1 U306 ( .A1(in_20), .A2(in_2), .ZN(n660) );
  AND2_X1 U306bar ( .A1(in_20bar), .A2(in_2bar), .ZN(n660bar) );
  OR2_X1 U307 ( .A1(n658), .A2(n657), .ZN(n662) );
  AND2_X1 U307bar ( .A1(n658bar), .A2(n657bar), .ZN(n662bar) );
  OR2_X1 U308 ( .A1(in_30), .A2(in_3), .ZN(n657) );
  AND2_X1 U308bar ( .A1(in_30bar), .A2(in_3bar), .ZN(n657bar) );
  OR2_X1 U309 ( .A1(in_4), .A2(in_38), .ZN(n658) );
  AND2_X1 U309bar ( .A1(in_4bar), .A2(in_38bar), .ZN(n658bar) );
  OR2_X1 U310 ( .A1(n656), .A2(n655), .ZN(n702) );
  AND2_X1 U310bar ( .A1(n656bar), .A2(n655bar), .ZN(n702bar) );
  OR2_X1 U311 ( .A1(in[148]), .A2(in[137]), .ZN(n655) );
  AND2_X1 U311bar ( .A1(inbar[148]), .A2(inbar[137]), .ZN(n655bar) );
  OR2_X1 U312 ( .A1(in[149]), .A2(n654), .ZN(n656) );
  AND2_X1 U312bar ( .A1(inbar[149]), .A2(n654bar), .ZN(n656bar) );
  OR2_X1 U313 ( .A1(in[195]), .A2(in[190]), .ZN(n654) );
  AND2_X1 U313bar ( .A1(inbar[195]), .A2(inbar[190]), .ZN(n654bar) );
  OR2_X1 U314 ( .A1(n653), .A2(n652), .ZN(n704) );
  AND2_X1 U314bar ( .A1(n653bar), .A2(n652bar), .ZN(n704bar) );
  OR2_X1 U315 ( .A1(n651), .A2(n650), .ZN(n652) );
  AND2_X1 U315bar ( .A1(n651bar), .A2(n650bar), .ZN(n652bar) );
  OR2_X1 U316 ( .A1(in[98]), .A2(in[197]), .ZN(n650) );
  AND2_X1 U316bar ( .A1(inbar[98]), .A2(inbar[197]), .ZN(n650bar) );
  OR2_X1 U317 ( .A1(in_11), .A2(n649), .ZN(n651) );
  AND2_X1 U317bar ( .A1(in_11bar), .A2(n649bar), .ZN(n651bar) );
  OR2_X1 U318 ( .A1(in_26), .A2(in_14), .ZN(n649) );
  AND2_X1 U318bar ( .A1(in_26bar), .A2(in_14bar), .ZN(n649bar) );
  OR2_X1 U319 ( .A1(n648), .A2(n647), .ZN(n653) );
  AND2_X1 U319bar ( .A1(n648bar), .A2(n647bar), .ZN(n653bar) );
  OR2_X1 U320 ( .A1(in_35), .A2(in_27), .ZN(n647) );
  AND2_X1 U320bar ( .A1(in_35bar), .A2(in_27bar), .ZN(n647bar) );
  OR2_X1 U321 ( .A1(in_50), .A2(n646), .ZN(n648) );
  AND2_X1 U321bar ( .A1(in_50bar), .A2(n646bar), .ZN(n648bar) );
  OR2_X1 U322 ( .A1(in_78), .A2(in_61), .ZN(n646) );
  AND2_X1 U322bar ( .A1(in_78bar), .A2(in_61bar), .ZN(n646bar) );
  OR2_X1 U323 ( .A1(n942), .A2(n645), .ZN(n720) );
  AND2_X1 U323bar ( .A1(n942bar), .A2(n645bar), .ZN(n720bar) );
  OR2_X1 U324 ( .A1(in[106]), .A2(n863), .ZN(n645) );
  AND2_X1 U324bar ( .A1(inbar[106]), .A2(n863bar), .ZN(n645bar) );
  OR2_X1 U325 ( .A1(n644), .A2(n643), .ZN(n863) );
  AND2_X1 U325bar ( .A1(n644bar), .A2(n643bar), .ZN(n863bar) );
  OR2_X1 U326 ( .A1(n642), .A2(n641), .ZN(n643) );
  AND2_X1 U326bar ( .A1(n642bar), .A2(n641bar), .ZN(n643bar) );
  OR2_X1 U327 ( .A1(n640), .A2(n639), .ZN(n641) );
  AND2_X1 U327bar ( .A1(n640bar), .A2(n639bar), .ZN(n641bar) );
  OR2_X1 U328 ( .A1(in[127]), .A2(in[122]), .ZN(n639) );
  AND2_X1 U328bar ( .A1(inbar[127]), .A2(inbar[122]), .ZN(n639bar) );
  OR2_X1 U329 ( .A1(in[156]), .A2(in[132]), .ZN(n640) );
  AND2_X1 U329bar ( .A1(inbar[156]), .A2(inbar[132]), .ZN(n640bar) );
  OR2_X1 U330 ( .A1(n638), .A2(n637), .ZN(n642) );
  AND2_X1 U330bar ( .A1(n638bar), .A2(n637bar), .ZN(n642bar) );
  OR2_X1 U331 ( .A1(in[159]), .A2(in[157]), .ZN(n637) );
  AND2_X1 U331bar ( .A1(inbar[159]), .A2(inbar[157]), .ZN(n637bar) );
  OR2_X1 U332 ( .A1(in[185]), .A2(in[169]), .ZN(n638) );
  AND2_X1 U332bar ( .A1(inbar[185]), .A2(inbar[169]), .ZN(n638bar) );
  OR2_X1 U333 ( .A1(n636), .A2(n635), .ZN(n644) );
  AND2_X1 U333bar ( .A1(n636bar), .A2(n635bar), .ZN(n644bar) );
  OR2_X1 U334 ( .A1(n634), .A2(n633), .ZN(n635) );
  AND2_X1 U334bar ( .A1(n634bar), .A2(n633bar), .ZN(n635bar) );
  OR2_X1 U335 ( .A1(in[239]), .A2(in[218]), .ZN(n633) );
  AND2_X1 U335bar ( .A1(inbar[239]), .A2(inbar[218]), .ZN(n633bar) );
  OR2_X1 U336 ( .A1(in_13), .A2(in[87]), .ZN(n634) );
  AND2_X1 U336bar ( .A1(in_13bar), .A2(inbar[87]), .ZN(n634bar) );
  OR2_X1 U337 ( .A1(n632), .A2(n631), .ZN(n636) );
  AND2_X1 U337bar ( .A1(n632bar), .A2(n631bar), .ZN(n636bar) );
  OR2_X1 U338 ( .A1(in_72), .A2(in_70), .ZN(n631) );
  AND2_X1 U338bar ( .A1(in_72bar), .A2(in_70bar), .ZN(n631bar) );
  OR2_X1 U339 ( .A1(in_80), .A2(in_74), .ZN(n632) );
  AND2_X1 U339bar ( .A1(in_80bar), .A2(in_74bar), .ZN(n632bar) );
  OR2_X1 U340 ( .A1(n630), .A2(n629), .ZN(n942) );
  AND2_X1 U340bar ( .A1(n630bar), .A2(n629bar), .ZN(n942bar) );
  OR2_X1 U341 ( .A1(n628), .A2(n627), .ZN(n629) );
  AND2_X1 U341bar ( .A1(n628bar), .A2(n627bar), .ZN(n629bar) );
  OR2_X1 U342 ( .A1(n626), .A2(n625), .ZN(n627) );
  AND2_X1 U342bar ( .A1(n626bar), .A2(n625bar), .ZN(n627bar) );
  OR2_X1 U343 ( .A1(in[146]), .A2(in[100]), .ZN(n625) );
  AND2_X1 U343bar ( .A1(inbar[146]), .A2(inbar[100]), .ZN(n625bar) );
  OR2_X1 U344 ( .A1(in[168]), .A2(in[152]), .ZN(n626) );
  AND2_X1 U344bar ( .A1(inbar[168]), .A2(inbar[152]), .ZN(n626bar) );
  OR2_X1 U345 ( .A1(n624), .A2(n623), .ZN(n628) );
  AND2_X1 U345bar ( .A1(n624bar), .A2(n623bar), .ZN(n628bar) );
  OR2_X1 U346 ( .A1(in[199]), .A2(in[182]), .ZN(n623) );
  AND2_X1 U346bar ( .A1(inbar[199]), .A2(inbar[182]), .ZN(n623bar) );
  OR2_X1 U347 ( .A1(in[236]), .A2(in[204]), .ZN(n624) );
  AND2_X1 U347bar ( .A1(inbar[236]), .A2(inbar[204]), .ZN(n624bar) );
  OR2_X1 U348 ( .A1(n622), .A2(n621), .ZN(n630) );
  AND2_X1 U348bar ( .A1(n622bar), .A2(n621bar), .ZN(n630bar) );
  OR2_X1 U349 ( .A1(n620), .A2(n619), .ZN(n621) );
  AND2_X1 U349bar ( .A1(n620bar), .A2(n619bar), .ZN(n621bar) );
  OR2_X1 U350 ( .A1(in[89]), .A2(in[246]), .ZN(n619) );
  AND2_X1 U350bar ( .A1(inbar[89]), .A2(inbar[246]), .ZN(n619bar) );
  OR2_X1 U351 ( .A1(in[95]), .A2(in[92]), .ZN(n620) );
  AND2_X1 U351bar ( .A1(inbar[95]), .A2(inbar[92]), .ZN(n620bar) );
  OR2_X1 U352 ( .A1(n618), .A2(n617), .ZN(n622) );
  AND2_X1 U352bar ( .A1(n618bar), .A2(n617bar), .ZN(n622bar) );
  OR2_X1 U353 ( .A1(in_22), .A2(in_16), .ZN(n617) );
  AND2_X1 U353bar ( .A1(in_22bar), .A2(in_16bar), .ZN(n617bar) );
  OR2_X1 U354 ( .A1(in_51), .A2(in_49), .ZN(n618) );
  AND2_X1 U354bar ( .A1(in_51bar), .A2(in_49bar), .ZN(n618bar) );
  OR2_X1 U355 ( .A1(n616), .A2(n615), .ZN(n722) );
  AND2_X1 U355bar ( .A1(n616bar), .A2(n615bar), .ZN(n722bar) );
  OR2_X1 U356 ( .A1(in[158]), .A2(in[115]), .ZN(n615) );
  AND2_X1 U356bar ( .A1(inbar[158]), .A2(inbar[115]), .ZN(n615bar) );
  OR2_X1 U357 ( .A1(in[163]), .A2(n614), .ZN(n616) );
  AND2_X1 U357bar ( .A1(inbar[163]), .A2(n614bar), .ZN(n616bar) );
  OR2_X1 U358 ( .A1(in[206]), .A2(in[165]), .ZN(n614) );
  AND2_X1 U358bar ( .A1(inbar[206]), .A2(inbar[165]), .ZN(n614bar) );
  OR2_X1 U359 ( .A1(n613), .A2(n612), .ZN(n724) );
  AND2_X1 U359bar ( .A1(n613bar), .A2(n612bar), .ZN(n724bar) );
  OR2_X1 U360 ( .A1(n611), .A2(n610), .ZN(n612) );
  AND2_X1 U360bar ( .A1(n611bar), .A2(n610bar), .ZN(n612bar) );
  OR2_X1 U361 ( .A1(in[213]), .A2(in[207]), .ZN(n610) );
  AND2_X1 U361bar ( .A1(inbar[213]), .A2(inbar[207]), .ZN(n610bar) );
  OR2_X1 U362 ( .A1(in[215]), .A2(n609), .ZN(n611) );
  AND2_X1 U362bar ( .A1(inbar[215]), .A2(n609bar), .ZN(n611bar) );
  OR2_X1 U363 ( .A1(in[230]), .A2(in[220]), .ZN(n609) );
  AND2_X1 U363bar ( .A1(inbar[230]), .A2(inbar[220]), .ZN(n609bar) );
  OR2_X1 U364 ( .A1(n608), .A2(n607), .ZN(n613) );
  AND2_X1 U364bar ( .A1(n608bar), .A2(n607bar), .ZN(n613bar) );
  OR2_X1 U365 ( .A1(in[251]), .A2(in[234]), .ZN(n607) );
  AND2_X1 U365bar ( .A1(inbar[251]), .A2(inbar[234]), .ZN(n607bar) );
  OR2_X1 U366 ( .A1(in_17), .A2(n606), .ZN(n608) );
  AND2_X1 U366bar ( .A1(in_17bar), .A2(n606bar), .ZN(n608bar) );
  OR2_X1 U367 ( .A1(in_65), .A2(in_56), .ZN(n606) );
  AND2_X1 U367bar ( .A1(in_65bar), .A2(in_56bar), .ZN(n606bar) );
  OR2_X1 U368 ( .A1(n605), .A2(n604), .ZN(out[0]) );
  AND2_X1 U368bar ( .A1(n605bar), .A2(n604bar), .ZN(outbar[0]) );
  OR2_X1 U369 ( .A1(n603), .A2(n602), .ZN(n604) );
  AND2_X1 U369bar ( .A1(n603bar), .A2(n602bar), .ZN(n604bar) );
  OR2_X1 U370 ( .A1(n601), .A2(n600), .ZN(n602) );
  AND2_X1 U370bar ( .A1(n601bar), .A2(n600bar), .ZN(n602bar) );
  OR2_X1 U371 ( .A1(n820), .A2(n785), .ZN(n600) );
  AND2_X1 U371bar ( .A1(n820bar), .A2(n785bar), .ZN(n600bar) );
  OR2_X1 U372 ( .A1(n599), .A2(n598), .ZN(n785) );
  AND2_X1 U372bar ( .A1(n599bar), .A2(n598bar), .ZN(n785bar) );
  OR2_X1 U373 ( .A1(n597), .A2(n596), .ZN(n598) );
  AND2_X1 U373bar ( .A1(n597bar), .A2(n596bar), .ZN(n598bar) );
  OR2_X1 U374 ( .A1(n595), .A2(n594), .ZN(n596) );
  AND2_X1 U374bar ( .A1(n595bar), .A2(n594bar), .ZN(n596bar) );
  OR2_X1 U375 ( .A1(in[135]), .A2(in[104]), .ZN(n594) );
  AND2_X1 U375bar ( .A1(inbar[135]), .A2(inbar[104]), .ZN(n594bar) );
  OR2_X1 U376 ( .A1(in[188]), .A2(in[178]), .ZN(n595) );
  AND2_X1 U376bar ( .A1(inbar[188]), .A2(inbar[178]), .ZN(n595bar) );
  OR2_X1 U377 ( .A1(n593), .A2(n592), .ZN(n597) );
  AND2_X1 U377bar ( .A1(n593bar), .A2(n592bar), .ZN(n597bar) );
  OR2_X1 U378 ( .A1(in[217]), .A2(in[194]), .ZN(n592) );
  AND2_X1 U378bar ( .A1(inbar[217]), .A2(inbar[194]), .ZN(n592bar) );
  OR2_X1 U379 ( .A1(in[237]), .A2(in[218]), .ZN(n593) );
  AND2_X1 U379bar ( .A1(inbar[237]), .A2(inbar[218]), .ZN(n593bar) );
  OR2_X1 U380 ( .A1(n591), .A2(n590), .ZN(n599) );
  AND2_X1 U380bar ( .A1(n591bar), .A2(n590bar), .ZN(n599bar) );
  OR2_X1 U381 ( .A1(n589), .A2(n588), .ZN(n590) );
  AND2_X1 U381bar ( .A1(n589bar), .A2(n588bar), .ZN(n590bar) );
  OR2_X1 U382 ( .A1(in_2), .A2(in_10), .ZN(n588) );
  AND2_X1 U382bar ( .A1(in_2bar), .A2(in_10bar), .ZN(n588bar) );
  OR2_X1 U383 ( .A1(in_47), .A2(in_22), .ZN(n589) );
  AND2_X1 U383bar ( .A1(in_47bar), .A2(in_22bar), .ZN(n589bar) );
  OR2_X1 U384 ( .A1(n587), .A2(n586), .ZN(n591) );
  AND2_X1 U384bar ( .A1(n587bar), .A2(n586bar), .ZN(n591bar) );
  OR2_X1 U385 ( .A1(in_56), .A2(in_54), .ZN(n586) );
  AND2_X1 U385bar ( .A1(in_56bar), .A2(in_54bar), .ZN(n586bar) );
  OR2_X1 U386 ( .A1(in_63), .A2(in_61), .ZN(n587) );
  AND2_X1 U386bar ( .A1(in_63bar), .A2(in_61bar), .ZN(n587bar) );
  OR2_X1 U387 ( .A1(n585), .A2(n584), .ZN(n820) );
  AND2_X1 U387bar ( .A1(n585bar), .A2(n584bar), .ZN(n820bar) );
  OR2_X1 U388 ( .A1(n583), .A2(n582), .ZN(n584) );
  AND2_X1 U388bar ( .A1(n583bar), .A2(n582bar), .ZN(n584bar) );
  OR2_X1 U389 ( .A1(n581), .A2(n580), .ZN(n582) );
  AND2_X1 U389bar ( .A1(n581bar), .A2(n580bar), .ZN(n582bar) );
  OR2_X1 U390 ( .A1(in[158]), .A2(in[142]), .ZN(n580) );
  AND2_X1 U390bar ( .A1(inbar[158]), .A2(inbar[142]), .ZN(n580bar) );
  OR2_X1 U391 ( .A1(in[175]), .A2(in[164]), .ZN(n581) );
  AND2_X1 U391bar ( .A1(inbar[175]), .A2(inbar[164]), .ZN(n581bar) );
  OR2_X1 U392 ( .A1(n579), .A2(n578), .ZN(n583) );
  AND2_X1 U392bar ( .A1(n579bar), .A2(n578bar), .ZN(n583bar) );
  OR2_X1 U393 ( .A1(in[228]), .A2(in[204]), .ZN(n578) );
  AND2_X1 U393bar ( .A1(inbar[228]), .A2(inbar[204]), .ZN(n578bar) );
  OR2_X1 U394 ( .A1(in[91]), .A2(in[87]), .ZN(n579) );
  AND2_X1 U394bar ( .A1(inbar[91]), .A2(inbar[87]), .ZN(n579bar) );
  OR2_X1 U395 ( .A1(n577), .A2(n576), .ZN(n585) );
  AND2_X1 U395bar ( .A1(n577bar), .A2(n576bar), .ZN(n585bar) );
  OR2_X1 U396 ( .A1(n575), .A2(n574), .ZN(n576) );
  AND2_X1 U396bar ( .A1(n575bar), .A2(n574bar), .ZN(n576bar) );
  OR2_X1 U397 ( .A1(in_21), .A2(in_11), .ZN(n574) );
  AND2_X1 U397bar ( .A1(in_21bar), .A2(in_11bar), .ZN(n574bar) );
  OR2_X1 U398 ( .A1(in_5), .A2(in_3), .ZN(n575) );
  AND2_X1 U398bar ( .A1(in_5bar), .A2(in_3bar), .ZN(n575bar) );
  OR2_X1 U399 ( .A1(n573), .A2(n572), .ZN(n577) );
  AND2_X1 U399bar ( .A1(n573bar), .A2(n572bar), .ZN(n577bar) );
  OR2_X1 U400 ( .A1(in_68), .A2(in_64), .ZN(n572) );
  AND2_X1 U400bar ( .A1(in_68bar), .A2(in_64bar), .ZN(n572bar) );
  OR2_X1 U401 ( .A1(in_76), .A2(in_73), .ZN(n573) );
  AND2_X1 U401bar ( .A1(in_76bar), .A2(in_73bar), .ZN(n573bar) );
  OR2_X1 U402 ( .A1(n778), .A2(n571), .ZN(n601) );
  AND2_X1 U402bar ( .A1(n778bar), .A2(n571bar), .ZN(n601bar) );
  OR2_X1 U403 ( .A1(in[100]), .A2(n965), .ZN(n571) );
  AND2_X1 U403bar ( .A1(inbar[100]), .A2(n965bar), .ZN(n571bar) );
  OR2_X1 U404 ( .A1(n570), .A2(n569), .ZN(n965) );
  AND2_X1 U404bar ( .A1(n570bar), .A2(n569bar), .ZN(n965bar) );
  OR2_X1 U405 ( .A1(n568), .A2(n567), .ZN(n569) );
  AND2_X1 U405bar ( .A1(n568bar), .A2(n567bar), .ZN(n569bar) );
  OR2_X1 U406 ( .A1(n566), .A2(n565), .ZN(n567) );
  AND2_X1 U406bar ( .A1(n566bar), .A2(n565bar), .ZN(n567bar) );
  OR2_X1 U407 ( .A1(n817), .A2(n750), .ZN(n565) );
  AND2_X1 U407bar ( .A1(n817bar), .A2(n750bar), .ZN(n565bar) );
  OR2_X1 U408 ( .A1(n564), .A2(n563), .ZN(n750) );
  AND2_X1 U408bar ( .A1(n564bar), .A2(n563bar), .ZN(n750bar) );
  OR2_X1 U409 ( .A1(n562), .A2(n561), .ZN(n563) );
  AND2_X1 U409bar ( .A1(n562bar), .A2(n561bar), .ZN(n563bar) );
  OR2_X1 U410 ( .A1(n560), .A2(n559), .ZN(n561) );
  AND2_X1 U410bar ( .A1(n560bar), .A2(n559bar), .ZN(n561bar) );
  OR2_X1 U411 ( .A1(in[119]), .A2(in[103]), .ZN(n559) );
  AND2_X1 U411bar ( .A1(inbar[119]), .A2(inbar[103]), .ZN(n559bar) );
  OR2_X1 U412 ( .A1(in[137]), .A2(in[133]), .ZN(n560) );
  AND2_X1 U412bar ( .A1(inbar[137]), .A2(inbar[133]), .ZN(n560bar) );
  OR2_X1 U413 ( .A1(n558), .A2(n557), .ZN(n562) );
  AND2_X1 U413bar ( .A1(n558bar), .A2(n557bar), .ZN(n562bar) );
  OR2_X1 U414 ( .A1(in[176]), .A2(in[173]), .ZN(n557) );
  AND2_X1 U414bar ( .A1(inbar[176]), .A2(inbar[173]), .ZN(n557bar) );
  OR2_X1 U415 ( .A1(in[210]), .A2(in[181]), .ZN(n558) );
  AND2_X1 U415bar ( .A1(inbar[210]), .A2(inbar[181]), .ZN(n558bar) );
  OR2_X1 U416 ( .A1(n556), .A2(n555), .ZN(n564) );
  AND2_X1 U416bar ( .A1(n556bar), .A2(n555bar), .ZN(n564bar) );
  OR2_X1 U417 ( .A1(n554), .A2(n553), .ZN(n555) );
  AND2_X1 U417bar ( .A1(n554bar), .A2(n553bar), .ZN(n555bar) );
  OR2_X1 U418 ( .A1(in_13), .A2(in[234]), .ZN(n553) );
  AND2_X1 U418bar ( .A1(in_13bar), .A2(inbar[234]), .ZN(n553bar) );
  OR2_X1 U419 ( .A1(in_38), .A2(in_32), .ZN(n554) );
  AND2_X1 U419bar ( .A1(in_38bar), .A2(in_32bar), .ZN(n554bar) );
  OR2_X1 U420 ( .A1(n552), .A2(n551), .ZN(n556) );
  AND2_X1 U420bar ( .A1(n552bar), .A2(n551bar), .ZN(n556bar) );
  OR2_X1 U421 ( .A1(in_42), .A2(in_41), .ZN(n551) );
  AND2_X1 U421bar ( .A1(in_42bar), .A2(in_41bar), .ZN(n551bar) );
  OR2_X1 U422 ( .A1(in_7), .A2(in_49), .ZN(n552) );
  AND2_X1 U422bar ( .A1(in_7bar), .A2(in_49bar), .ZN(n552bar) );
  OR2_X1 U423 ( .A1(n550), .A2(n549), .ZN(n817) );
  AND2_X1 U423bar ( .A1(n550bar), .A2(n549bar), .ZN(n817bar) );
  OR2_X1 U424 ( .A1(n548), .A2(n547), .ZN(n549) );
  AND2_X1 U424bar ( .A1(n548bar), .A2(n547bar), .ZN(n549bar) );
  OR2_X1 U425 ( .A1(n546), .A2(n545), .ZN(n547) );
  AND2_X1 U425bar ( .A1(n546bar), .A2(n545bar), .ZN(n547bar) );
  OR2_X1 U426 ( .A1(in[159]), .A2(in[105]), .ZN(n545) );
  AND2_X1 U426bar ( .A1(inbar[159]), .A2(inbar[105]), .ZN(n545bar) );
  OR2_X1 U427 ( .A1(in[206]), .A2(in[183]), .ZN(n546) );
  AND2_X1 U427bar ( .A1(inbar[206]), .A2(inbar[183]), .ZN(n546bar) );
  OR2_X1 U428 ( .A1(n544), .A2(n543), .ZN(n548) );
  AND2_X1 U428bar ( .A1(n544bar), .A2(n543bar), .ZN(n548bar) );
  OR2_X1 U429 ( .A1(in[229]), .A2(in[219]), .ZN(n543) );
  AND2_X1 U429bar ( .A1(inbar[229]), .A2(inbar[219]), .ZN(n543bar) );
  OR2_X1 U430 ( .A1(in[235]), .A2(in[232]), .ZN(n544) );
  AND2_X1 U430bar ( .A1(inbar[235]), .A2(inbar[232]), .ZN(n544bar) );
  OR2_X1 U431 ( .A1(n542), .A2(n541), .ZN(n550) );
  AND2_X1 U431bar ( .A1(n542bar), .A2(n541bar), .ZN(n550bar) );
  OR2_X1 U432 ( .A1(n540), .A2(n539), .ZN(n541) );
  AND2_X1 U432bar ( .A1(n540bar), .A2(n539bar), .ZN(n541bar) );
  OR2_X1 U433 ( .A1(in[249]), .A2(in[242]), .ZN(n539) );
  AND2_X1 U433bar ( .A1(inbar[249]), .A2(inbar[242]), .ZN(n539bar) );
  OR2_X1 U434 ( .A1(in[89]), .A2(in[254]), .ZN(n540) );
  AND2_X1 U434bar ( .A1(inbar[89]), .A2(inbar[254]), .ZN(n540bar) );
  OR2_X1 U435 ( .A1(n538), .A2(n537), .ZN(n542) );
  AND2_X1 U435bar ( .A1(n538bar), .A2(n537bar), .ZN(n542bar) );
  OR2_X1 U436 ( .A1(in_14), .A2(in[99]), .ZN(n537) );
  AND2_X1 U436bar ( .A1(in_14bar), .A2(inbar[99]), .ZN(n537bar) );
  OR2_X1 U437 ( .A1(in_60), .A2(in_18), .ZN(n538) );
  AND2_X1 U437bar ( .A1(in_60bar), .A2(in_18bar), .ZN(n538bar) );
  OR2_X1 U438 ( .A1(in[113]), .A2(n763), .ZN(n566) );
  AND2_X1 U438bar ( .A1(inbar[113]), .A2(n763bar), .ZN(n566bar) );
  OR2_X1 U439 ( .A1(n536), .A2(n535), .ZN(n763) );
  AND2_X1 U439bar ( .A1(n536bar), .A2(n535bar), .ZN(n763bar) );
  OR2_X1 U440 ( .A1(n534), .A2(n533), .ZN(n535) );
  AND2_X1 U440bar ( .A1(n534bar), .A2(n533bar), .ZN(n535bar) );
  OR2_X1 U441 ( .A1(n532), .A2(n531), .ZN(n533) );
  AND2_X1 U441bar ( .A1(n532bar), .A2(n531bar), .ZN(n533bar) );
  OR2_X1 U442 ( .A1(in[115]), .A2(in[110]), .ZN(n531) );
  AND2_X1 U442bar ( .A1(inbar[115]), .A2(inbar[110]), .ZN(n531bar) );
  OR2_X1 U443 ( .A1(in[125]), .A2(in[117]), .ZN(n532) );
  AND2_X1 U443bar ( .A1(inbar[125]), .A2(inbar[117]), .ZN(n532bar) );
  OR2_X1 U444 ( .A1(n530), .A2(n529), .ZN(n534) );
  AND2_X1 U444bar ( .A1(n530bar), .A2(n529bar), .ZN(n534bar) );
  OR2_X1 U445 ( .A1(in[180]), .A2(in[128]), .ZN(n529) );
  AND2_X1 U445bar ( .A1(inbar[180]), .A2(inbar[128]), .ZN(n529bar) );
  OR2_X1 U446 ( .A1(in[205]), .A2(in[201]), .ZN(n530) );
  AND2_X1 U446bar ( .A1(inbar[205]), .A2(inbar[201]), .ZN(n530bar) );
  OR2_X1 U447 ( .A1(n528), .A2(n527), .ZN(n536) );
  AND2_X1 U447bar ( .A1(n528bar), .A2(n527bar), .ZN(n536bar) );
  OR2_X1 U448 ( .A1(n526), .A2(n525), .ZN(n527) );
  AND2_X1 U448bar ( .A1(n526bar), .A2(n525bar), .ZN(n527bar) );
  OR2_X1 U449 ( .A1(in[244]), .A2(in[239]), .ZN(n525) );
  AND2_X1 U449bar ( .A1(inbar[244]), .A2(inbar[239]), .ZN(n525bar) );
  OR2_X1 U450 ( .A1(in[95]), .A2(in[83]), .ZN(n526) );
  AND2_X1 U450bar ( .A1(inbar[95]), .A2(inbar[83]), .ZN(n526bar) );
  OR2_X1 U451 ( .A1(n524), .A2(n523), .ZN(n528) );
  AND2_X1 U451bar ( .A1(n524bar), .A2(n523bar), .ZN(n528bar) );
  OR2_X1 U452 ( .A1(in_24), .A2(in[97]), .ZN(n523) );
  AND2_X1 U452bar ( .A1(in_24bar), .A2(inbar[97]), .ZN(n523bar) );
  OR2_X1 U453 ( .A1(in_33), .A2(in_27), .ZN(n524) );
  AND2_X1 U453bar ( .A1(in_33bar), .A2(in_27bar), .ZN(n524bar) );
  OR2_X1 U454 ( .A1(n522), .A2(n521), .ZN(n568) );
  AND2_X1 U454bar ( .A1(n522bar), .A2(n521bar), .ZN(n568bar) );
  OR2_X1 U455 ( .A1(in[145]), .A2(in[126]), .ZN(n521) );
  AND2_X1 U455bar ( .A1(inbar[145]), .A2(inbar[126]), .ZN(n521bar) );
  OR2_X1 U456 ( .A1(in[169]), .A2(n520), .ZN(n522) );
  AND2_X1 U456bar ( .A1(inbar[169]), .A2(n520bar), .ZN(n522bar) );
  OR2_X1 U457 ( .A1(in[221]), .A2(in[172]), .ZN(n520) );
  AND2_X1 U457bar ( .A1(inbar[221]), .A2(inbar[172]), .ZN(n520bar) );
  OR2_X1 U458 ( .A1(n519), .A2(n518), .ZN(n570) );
  AND2_X1 U458bar ( .A1(n519bar), .A2(n518bar), .ZN(n570bar) );
  OR2_X1 U459 ( .A1(n517), .A2(n516), .ZN(n518) );
  AND2_X1 U459bar ( .A1(n517bar), .A2(n516bar), .ZN(n518bar) );
  OR2_X1 U460 ( .A1(in[241]), .A2(in[224]), .ZN(n516) );
  AND2_X1 U460bar ( .A1(inbar[241]), .A2(inbar[224]), .ZN(n516bar) );
  OR2_X1 U461 ( .A1(in[86]), .A2(n515), .ZN(n517) );
  AND2_X1 U461bar ( .A1(inbar[86]), .A2(n515bar), .ZN(n517bar) );
  OR2_X1 U462 ( .A1(in_43), .A2(in_34), .ZN(n515) );
  AND2_X1 U462bar ( .A1(in_43bar), .A2(in_34bar), .ZN(n515bar) );
  OR2_X1 U463 ( .A1(n514), .A2(n513), .ZN(n519) );
  AND2_X1 U463bar ( .A1(n514bar), .A2(n513bar), .ZN(n519bar) );
  OR2_X1 U464 ( .A1(in_65), .A2(in_51), .ZN(n513) );
  AND2_X1 U464bar ( .A1(in_65bar), .A2(in_51bar), .ZN(n513bar) );
  OR2_X1 U465 ( .A1(in_75), .A2(n512), .ZN(n514) );
  AND2_X1 U465bar ( .A1(in_75bar), .A2(n512bar), .ZN(n514bar) );
  OR2_X1 U466 ( .A1(in_81), .A2(in_77), .ZN(n512) );
  AND2_X1 U466bar ( .A1(in_81bar), .A2(in_77bar), .ZN(n512bar) );
  OR2_X1 U467 ( .A1(n511), .A2(n510), .ZN(n778) );
  AND2_X1 U467bar ( .A1(n511bar), .A2(n510bar), .ZN(n778bar) );
  OR2_X1 U468 ( .A1(n509), .A2(n508), .ZN(n510) );
  AND2_X1 U468bar ( .A1(n509bar), .A2(n508bar), .ZN(n510bar) );
  OR2_X1 U469 ( .A1(n507), .A2(n506), .ZN(n508) );
  AND2_X1 U469bar ( .A1(n507bar), .A2(n506bar), .ZN(n508bar) );
  OR2_X1 U470 ( .A1(in[107]), .A2(in[101]), .ZN(n506) );
  AND2_X1 U470bar ( .A1(inbar[107]), .A2(inbar[101]), .ZN(n506bar) );
  OR2_X1 U471 ( .A1(in[139]), .A2(in[132]), .ZN(n507) );
  AND2_X1 U471bar ( .A1(inbar[139]), .A2(inbar[132]), .ZN(n507bar) );
  OR2_X1 U472 ( .A1(n505), .A2(n504), .ZN(n509) );
  AND2_X1 U472bar ( .A1(n505bar), .A2(n504bar), .ZN(n509bar) );
  OR2_X1 U473 ( .A1(in[146]), .A2(in[141]), .ZN(n504) );
  AND2_X1 U473bar ( .A1(inbar[146]), .A2(inbar[141]), .ZN(n504bar) );
  OR2_X1 U474 ( .A1(in[203]), .A2(in[179]), .ZN(n505) );
  AND2_X1 U474bar ( .A1(inbar[203]), .A2(inbar[179]), .ZN(n505bar) );
  OR2_X1 U475 ( .A1(n503), .A2(n502), .ZN(n511) );
  AND2_X1 U475bar ( .A1(n503bar), .A2(n502bar), .ZN(n511bar) );
  OR2_X1 U476 ( .A1(n501), .A2(n500), .ZN(n502) );
  AND2_X1 U476bar ( .A1(n501bar), .A2(n500bar), .ZN(n502bar) );
  OR2_X1 U477 ( .A1(in[243]), .A2(in[222]), .ZN(n500) );
  AND2_X1 U477bar ( .A1(inbar[243]), .A2(inbar[222]), .ZN(n500bar) );
  OR2_X1 U478 ( .A1(in[251]), .A2(in[250]), .ZN(n501) );
  AND2_X1 U478bar ( .A1(inbar[251]), .A2(inbar[250]), .ZN(n501bar) );
  OR2_X1 U479 ( .A1(n499), .A2(n498), .ZN(n503) );
  AND2_X1 U479bar ( .A1(n499bar), .A2(n498bar), .ZN(n503bar) );
  OR2_X1 U480 ( .A1(in_37), .A2(in_19), .ZN(n498) );
  AND2_X1 U480bar ( .A1(in_37bar), .A2(in_19bar), .ZN(n498bar) );
  OR2_X1 U481 ( .A1(in_78), .A2(in_6), .ZN(n499) );
  AND2_X1 U481bar ( .A1(in_78bar), .A2(in_6bar), .ZN(n499bar) );
  OR2_X1 U482 ( .A1(n497), .A2(n496), .ZN(n603) );
  AND2_X1 U482bar ( .A1(n497bar), .A2(n496bar), .ZN(n603bar) );
  OR2_X1 U483 ( .A1(in[112]), .A2(in[102]), .ZN(n496) );
  AND2_X1 U483bar ( .A1(inbar[112]), .A2(inbar[102]), .ZN(n496bar) );
  OR2_X1 U484 ( .A1(in[123]), .A2(n495), .ZN(n497) );
  AND2_X1 U484bar ( .A1(inbar[123]), .A2(n495bar), .ZN(n497bar) );
  OR2_X1 U485 ( .A1(in[143]), .A2(in[130]), .ZN(n495) );
  AND2_X1 U485bar ( .A1(inbar[143]), .A2(inbar[130]), .ZN(n495bar) );
  OR2_X1 U486 ( .A1(n494), .A2(n493), .ZN(n605) );
  AND2_X1 U486bar ( .A1(n494bar), .A2(n493bar), .ZN(n605bar) );
  OR2_X1 U487 ( .A1(n492), .A2(n491), .ZN(n493) );
  AND2_X1 U487bar ( .A1(n492bar), .A2(n491bar), .ZN(n493bar) );
  OR2_X1 U488 ( .A1(in[216]), .A2(in[213]), .ZN(n491) );
  AND2_X1 U488bar ( .A1(inbar[216]), .A2(inbar[213]), .ZN(n491bar) );
  OR2_X1 U489 ( .A1(in[227]), .A2(n490), .ZN(n492) );
  AND2_X1 U489bar ( .A1(inbar[227]), .A2(n490bar), .ZN(n492bar) );
  OR2_X1 U490 ( .A1(in_0), .A2(in[248]), .ZN(n490) );
  AND2_X1 U490bar ( .A1(in_0bar), .A2(inbar[248]), .ZN(n490bar) );
  OR2_X1 U491 ( .A1(n489), .A2(n488), .ZN(n494) );
  AND2_X1 U491bar ( .A1(n489bar), .A2(n488bar), .ZN(n494bar) );
  OR2_X1 U492 ( .A1(in_46), .A2(in_44), .ZN(n488) );
  AND2_X1 U492bar ( .A1(in_46bar), .A2(in_44bar), .ZN(n488bar) );
  OR2_X1 U493 ( .A1(in_50), .A2(n487), .ZN(n489) );
  AND2_X1 U493bar ( .A1(in_50bar), .A2(n487bar), .ZN(n489bar) );
  OR2_X1 U494 ( .A1(in_9), .A2(in_80), .ZN(n487) );
  AND2_X1 U494bar ( .A1(in_9bar), .A2(in_80bar), .ZN(n487bar) );
endmodule

module sBox_10 ( in, inbar, out, outbar );

  input wire [7:0] in;
  input wire [7:0] inbar;
//input_done

  output wire [7:0] out;
  output wire [7:0] outbar;
//output_done

  wire [255:0] decodeOut;
  wire [255:0] decodeOutbar;
//wire_done

  decode_10 dec ( .in(in), .inbar(inbar), .out(decodeOut), .outbar(decodeOutbar) );
  encode_10 enc ( .in(decodeOut), .inbar(decodeOutbar), .out(out), .outbar(outbar) );
endmodule

module CD2_41 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD2_42 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD2_43 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD2_44 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD4_21 ( a, abar, b, bbar, y, ybar );

  input wire [3:0] a;
  input wire [3:0] b;
  input wire [3:0] abar;
  input wire [3:0] bbar;
//input_done

  output wire [15:0] y;
  output wire [15:0] ybar;
//output_done

//wire_done

  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]) );
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]) );
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]) );
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]) );
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]) );
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]) );
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]) );
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]) );
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]) );
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]) );
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]) );
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]) );
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]) );
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]) );
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]) );
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]) );
endmodule

module CD4_22 ( a, abar, b, bbar, y, ybar );

  input wire [3:0] a;
  input wire [3:0] b;
  input wire [3:0] abar;
  input wire [3:0] bbar;
//input_done

  output wire [15:0] y;
  output wire [15:0] ybar;
//output_done

//wire_done

  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]) );
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]) );
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]) );
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]) );
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]) );
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]) );
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]) );
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]) );
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]) );
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]) );
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]) );
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]) );
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]) );
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]) );
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]) );
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]) );
endmodule

module CD16_11 ( a, abar, b, bbar, y, ybar );

  input wire [15:0] a;
  input wire [15:0] b;
  input wire [15:0] abar;
  input wire [15:0] bbar;
//input_done

  output wire [255:0] y;
  output wire [255:0] ybar;
//output_done

//wire_done

  AND2_X1 U1 ( .A1(b[9]), .A2(a[0]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[9]), .A2(abar[0]), .ZN(ybar[9]) );
  AND2_X1 U2 ( .A1(b[3]), .A2(a[6]), .ZN(y[99]) );
  OR2_X1 U2bar ( .A1(bbar[3]), .A2(abar[6]), .ZN(ybar[99]) );
  AND2_X1 U3 ( .A1(b[2]), .A2(a[6]), .ZN(y[98]) );
  OR2_X1 U3bar ( .A1(bbar[2]), .A2(abar[6]), .ZN(ybar[98]) );
  AND2_X1 U4 ( .A1(b[1]), .A2(a[6]), .ZN(y[97]) );
  OR2_X1 U4bar ( .A1(bbar[1]), .A2(abar[6]), .ZN(ybar[97]) );
  AND2_X1 U5 ( .A1(b[0]), .A2(a[6]), .ZN(y[96]) );
  OR2_X1 U5bar ( .A1(bbar[0]), .A2(abar[6]), .ZN(ybar[96]) );
  AND2_X1 U6 ( .A1(b[15]), .A2(a[5]), .ZN(y[95]) );
  OR2_X1 U6bar ( .A1(bbar[15]), .A2(abar[5]), .ZN(ybar[95]) );
  AND2_X1 U7 ( .A1(b[14]), .A2(a[5]), .ZN(y[94]) );
  OR2_X1 U7bar ( .A1(bbar[14]), .A2(abar[5]), .ZN(ybar[94]) );
  AND2_X1 U8 ( .A1(b[13]), .A2(a[5]), .ZN(y[93]) );
  OR2_X1 U8bar ( .A1(bbar[13]), .A2(abar[5]), .ZN(ybar[93]) );
  AND2_X1 U9 ( .A1(b[12]), .A2(a[5]), .ZN(y[92]) );
  OR2_X1 U9bar ( .A1(bbar[12]), .A2(abar[5]), .ZN(ybar[92]) );
  AND2_X1 U10 ( .A1(b[11]), .A2(a[5]), .ZN(y[91]) );
  OR2_X1 U10bar ( .A1(bbar[11]), .A2(abar[5]), .ZN(ybar[91]) );
  AND2_X1 U11 ( .A1(b[10]), .A2(a[5]), .ZN(y[90]) );
  OR2_X1 U11bar ( .A1(bbar[10]), .A2(abar[5]), .ZN(ybar[90]) );
  AND2_X1 U12 ( .A1(b[8]), .A2(a[0]), .ZN(y[8]) );
  OR2_X1 U12bar ( .A1(bbar[8]), .A2(abar[0]), .ZN(ybar[8]) );
  AND2_X1 U13 ( .A1(a[5]), .A2(b[9]), .ZN(y[89]) );
  OR2_X1 U13bar ( .A1(abar[5]), .A2(bbar[9]), .ZN(ybar[89]) );
  AND2_X1 U14 ( .A1(b[8]), .A2(a[5]), .ZN(y[88]) );
  OR2_X1 U14bar ( .A1(bbar[8]), .A2(abar[5]), .ZN(ybar[88]) );
  AND2_X1 U15 ( .A1(b[7]), .A2(a[5]), .ZN(y[87]) );
  OR2_X1 U15bar ( .A1(bbar[7]), .A2(abar[5]), .ZN(ybar[87]) );
  AND2_X1 U16 ( .A1(b[6]), .A2(a[5]), .ZN(y[86]) );
  OR2_X1 U16bar ( .A1(bbar[6]), .A2(abar[5]), .ZN(ybar[86]) );
  AND2_X1 U17 ( .A1(b[5]), .A2(a[5]), .ZN(y[85]) );
  OR2_X1 U17bar ( .A1(bbar[5]), .A2(abar[5]), .ZN(ybar[85]) );
  AND2_X1 U18 ( .A1(b[4]), .A2(a[5]), .ZN(y[84]) );
  OR2_X1 U18bar ( .A1(bbar[4]), .A2(abar[5]), .ZN(ybar[84]) );
  AND2_X1 U19 ( .A1(a[5]), .A2(b[3]), .ZN(y[83]) );
  OR2_X1 U19bar ( .A1(abar[5]), .A2(bbar[3]), .ZN(ybar[83]) );
  AND2_X1 U20 ( .A1(a[5]), .A2(b[2]), .ZN(y[82]) );
  OR2_X1 U20bar ( .A1(abar[5]), .A2(bbar[2]), .ZN(ybar[82]) );
  AND2_X1 U21 ( .A1(a[5]), .A2(b[1]), .ZN(y[81]) );
  OR2_X1 U21bar ( .A1(abar[5]), .A2(bbar[1]), .ZN(ybar[81]) );
  AND2_X1 U22 ( .A1(a[5]), .A2(b[0]), .ZN(y[80]) );
  OR2_X1 U22bar ( .A1(abar[5]), .A2(bbar[0]), .ZN(ybar[80]) );
  AND2_X1 U23 ( .A1(b[7]), .A2(a[0]), .ZN(y[7]) );
  OR2_X1 U23bar ( .A1(bbar[7]), .A2(abar[0]), .ZN(ybar[7]) );
  AND2_X1 U24 ( .A1(a[4]), .A2(b[15]), .ZN(y[79]) );
  OR2_X1 U24bar ( .A1(abar[4]), .A2(bbar[15]), .ZN(ybar[79]) );
  AND2_X1 U25 ( .A1(a[4]), .A2(b[14]), .ZN(y[78]) );
  OR2_X1 U25bar ( .A1(abar[4]), .A2(bbar[14]), .ZN(ybar[78]) );
  AND2_X1 U26 ( .A1(a[4]), .A2(b[13]), .ZN(y[77]) );
  OR2_X1 U26bar ( .A1(abar[4]), .A2(bbar[13]), .ZN(ybar[77]) );
  AND2_X1 U27 ( .A1(a[4]), .A2(b[12]), .ZN(y[76]) );
  OR2_X1 U27bar ( .A1(abar[4]), .A2(bbar[12]), .ZN(ybar[76]) );
  AND2_X1 U28 ( .A1(a[4]), .A2(b[11]), .ZN(y[75]) );
  OR2_X1 U28bar ( .A1(abar[4]), .A2(bbar[11]), .ZN(ybar[75]) );
  AND2_X1 U29 ( .A1(a[4]), .A2(b[10]), .ZN(y[74]) );
  OR2_X1 U29bar ( .A1(abar[4]), .A2(bbar[10]), .ZN(ybar[74]) );
  AND2_X1 U30 ( .A1(a[4]), .A2(b[9]), .ZN(y[73]) );
  OR2_X1 U30bar ( .A1(abar[4]), .A2(bbar[9]), .ZN(ybar[73]) );
  AND2_X1 U31 ( .A1(a[4]), .A2(b[8]), .ZN(y[72]) );
  OR2_X1 U31bar ( .A1(abar[4]), .A2(bbar[8]), .ZN(ybar[72]) );
  AND2_X1 U32 ( .A1(a[4]), .A2(b[7]), .ZN(y[71]) );
  OR2_X1 U32bar ( .A1(abar[4]), .A2(bbar[7]), .ZN(ybar[71]) );
  AND2_X1 U33 ( .A1(a[4]), .A2(b[6]), .ZN(y[70]) );
  OR2_X1 U33bar ( .A1(abar[4]), .A2(bbar[6]), .ZN(ybar[70]) );
  AND2_X1 U34 ( .A1(b[6]), .A2(a[0]), .ZN(y[6]) );
  OR2_X1 U34bar ( .A1(bbar[6]), .A2(abar[0]), .ZN(ybar[6]) );
  AND2_X1 U35 ( .A1(a[4]), .A2(b[5]), .ZN(y[69]) );
  OR2_X1 U35bar ( .A1(abar[4]), .A2(bbar[5]), .ZN(ybar[69]) );
  AND2_X1 U36 ( .A1(a[4]), .A2(b[4]), .ZN(y[68]) );
  OR2_X1 U36bar ( .A1(abar[4]), .A2(bbar[4]), .ZN(ybar[68]) );
  AND2_X1 U37 ( .A1(a[4]), .A2(b[3]), .ZN(y[67]) );
  OR2_X1 U37bar ( .A1(abar[4]), .A2(bbar[3]), .ZN(ybar[67]) );
  AND2_X1 U38 ( .A1(a[4]), .A2(b[2]), .ZN(y[66]) );
  OR2_X1 U38bar ( .A1(abar[4]), .A2(bbar[2]), .ZN(ybar[66]) );
  AND2_X1 U39 ( .A1(a[4]), .A2(b[1]), .ZN(y[65]) );
  OR2_X1 U39bar ( .A1(abar[4]), .A2(bbar[1]), .ZN(ybar[65]) );
  AND2_X1 U40 ( .A1(a[4]), .A2(b[0]), .ZN(y[64]) );
  OR2_X1 U40bar ( .A1(abar[4]), .A2(bbar[0]), .ZN(ybar[64]) );
  AND2_X1 U41 ( .A1(a[3]), .A2(b[15]), .ZN(y[63]) );
  OR2_X1 U41bar ( .A1(abar[3]), .A2(bbar[15]), .ZN(ybar[63]) );
  AND2_X1 U42 ( .A1(a[3]), .A2(b[14]), .ZN(y[62]) );
  OR2_X1 U42bar ( .A1(abar[3]), .A2(bbar[14]), .ZN(ybar[62]) );
  AND2_X1 U43 ( .A1(a[3]), .A2(b[13]), .ZN(y[61]) );
  OR2_X1 U43bar ( .A1(abar[3]), .A2(bbar[13]), .ZN(ybar[61]) );
  AND2_X1 U44 ( .A1(a[3]), .A2(b[12]), .ZN(y[60]) );
  OR2_X1 U44bar ( .A1(abar[3]), .A2(bbar[12]), .ZN(ybar[60]) );
  AND2_X1 U45 ( .A1(b[5]), .A2(a[0]), .ZN(y[5]) );
  OR2_X1 U45bar ( .A1(bbar[5]), .A2(abar[0]), .ZN(ybar[5]) );
  AND2_X1 U46 ( .A1(a[3]), .A2(b[11]), .ZN(y[59]) );
  OR2_X1 U46bar ( .A1(abar[3]), .A2(bbar[11]), .ZN(ybar[59]) );
  AND2_X1 U47 ( .A1(a[3]), .A2(b[10]), .ZN(y[58]) );
  OR2_X1 U47bar ( .A1(abar[3]), .A2(bbar[10]), .ZN(ybar[58]) );
  AND2_X1 U48 ( .A1(a[3]), .A2(b[9]), .ZN(y[57]) );
  OR2_X1 U48bar ( .A1(abar[3]), .A2(bbar[9]), .ZN(ybar[57]) );
  AND2_X1 U49 ( .A1(a[3]), .A2(b[8]), .ZN(y[56]) );
  OR2_X1 U49bar ( .A1(abar[3]), .A2(bbar[8]), .ZN(ybar[56]) );
  AND2_X1 U50 ( .A1(a[3]), .A2(b[7]), .ZN(y[55]) );
  OR2_X1 U50bar ( .A1(abar[3]), .A2(bbar[7]), .ZN(ybar[55]) );
  AND2_X1 U51 ( .A1(a[3]), .A2(b[6]), .ZN(y[54]) );
  OR2_X1 U51bar ( .A1(abar[3]), .A2(bbar[6]), .ZN(ybar[54]) );
  AND2_X1 U52 ( .A1(a[3]), .A2(b[5]), .ZN(y[53]) );
  OR2_X1 U52bar ( .A1(abar[3]), .A2(bbar[5]), .ZN(ybar[53]) );
  AND2_X1 U53 ( .A1(a[3]), .A2(b[4]), .ZN(y[52]) );
  OR2_X1 U53bar ( .A1(abar[3]), .A2(bbar[4]), .ZN(ybar[52]) );
  AND2_X1 U54 ( .A1(a[3]), .A2(b[3]), .ZN(y[51]) );
  OR2_X1 U54bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[51]) );
  AND2_X1 U55 ( .A1(a[3]), .A2(b[2]), .ZN(y[50]) );
  OR2_X1 U55bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[50]) );
  AND2_X1 U56 ( .A1(b[4]), .A2(a[0]), .ZN(y[4]) );
  OR2_X1 U56bar ( .A1(bbar[4]), .A2(abar[0]), .ZN(ybar[4]) );
  AND2_X1 U57 ( .A1(a[3]), .A2(b[1]), .ZN(y[49]) );
  OR2_X1 U57bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[49]) );
  AND2_X1 U58 ( .A1(a[3]), .A2(b[0]), .ZN(y[48]) );
  OR2_X1 U58bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[48]) );
  AND2_X1 U59 ( .A1(a[2]), .A2(b[15]), .ZN(y[47]) );
  OR2_X1 U59bar ( .A1(abar[2]), .A2(bbar[15]), .ZN(ybar[47]) );
  AND2_X1 U60 ( .A1(a[2]), .A2(b[14]), .ZN(y[46]) );
  OR2_X1 U60bar ( .A1(abar[2]), .A2(bbar[14]), .ZN(ybar[46]) );
  AND2_X1 U61 ( .A1(a[2]), .A2(b[13]), .ZN(y[45]) );
  OR2_X1 U61bar ( .A1(abar[2]), .A2(bbar[13]), .ZN(ybar[45]) );
  AND2_X1 U62 ( .A1(a[2]), .A2(b[12]), .ZN(y[44]) );
  OR2_X1 U62bar ( .A1(abar[2]), .A2(bbar[12]), .ZN(ybar[44]) );
  AND2_X1 U63 ( .A1(a[2]), .A2(b[11]), .ZN(y[43]) );
  OR2_X1 U63bar ( .A1(abar[2]), .A2(bbar[11]), .ZN(ybar[43]) );
  AND2_X1 U64 ( .A1(a[2]), .A2(b[10]), .ZN(y[42]) );
  OR2_X1 U64bar ( .A1(abar[2]), .A2(bbar[10]), .ZN(ybar[42]) );
  AND2_X1 U65 ( .A1(a[2]), .A2(b[9]), .ZN(y[41]) );
  OR2_X1 U65bar ( .A1(abar[2]), .A2(bbar[9]), .ZN(ybar[41]) );
  AND2_X1 U66 ( .A1(a[2]), .A2(b[8]), .ZN(y[40]) );
  OR2_X1 U66bar ( .A1(abar[2]), .A2(bbar[8]), .ZN(ybar[40]) );
  AND2_X1 U67 ( .A1(b[3]), .A2(a[0]), .ZN(y[3]) );
  OR2_X1 U67bar ( .A1(bbar[3]), .A2(abar[0]), .ZN(ybar[3]) );
  AND2_X1 U68 ( .A1(a[2]), .A2(b[7]), .ZN(y[39]) );
  OR2_X1 U68bar ( .A1(abar[2]), .A2(bbar[7]), .ZN(ybar[39]) );
  AND2_X1 U69 ( .A1(a[2]), .A2(b[6]), .ZN(y[38]) );
  OR2_X1 U69bar ( .A1(abar[2]), .A2(bbar[6]), .ZN(ybar[38]) );
  AND2_X1 U70 ( .A1(a[2]), .A2(b[5]), .ZN(y[37]) );
  OR2_X1 U70bar ( .A1(abar[2]), .A2(bbar[5]), .ZN(ybar[37]) );
  AND2_X1 U71 ( .A1(a[2]), .A2(b[4]), .ZN(y[36]) );
  OR2_X1 U71bar ( .A1(abar[2]), .A2(bbar[4]), .ZN(ybar[36]) );
  AND2_X1 U72 ( .A1(a[2]), .A2(b[3]), .ZN(y[35]) );
  OR2_X1 U72bar ( .A1(abar[2]), .A2(bbar[3]), .ZN(ybar[35]) );
  AND2_X1 U73 ( .A1(a[2]), .A2(b[2]), .ZN(y[34]) );
  OR2_X1 U73bar ( .A1(abar[2]), .A2(bbar[2]), .ZN(ybar[34]) );
  AND2_X1 U74 ( .A1(a[2]), .A2(b[1]), .ZN(y[33]) );
  OR2_X1 U74bar ( .A1(abar[2]), .A2(bbar[1]), .ZN(ybar[33]) );
  AND2_X1 U75 ( .A1(a[2]), .A2(b[0]), .ZN(y[32]) );
  OR2_X1 U75bar ( .A1(abar[2]), .A2(bbar[0]), .ZN(ybar[32]) );
  AND2_X1 U76 ( .A1(a[1]), .A2(b[15]), .ZN(y[31]) );
  OR2_X1 U76bar ( .A1(abar[1]), .A2(bbar[15]), .ZN(ybar[31]) );
  AND2_X1 U77 ( .A1(a[1]), .A2(b[14]), .ZN(y[30]) );
  OR2_X1 U77bar ( .A1(abar[1]), .A2(bbar[14]), .ZN(ybar[30]) );
  AND2_X1 U78 ( .A1(b[2]), .A2(a[0]), .ZN(y[2]) );
  OR2_X1 U78bar ( .A1(bbar[2]), .A2(abar[0]), .ZN(ybar[2]) );
  AND2_X1 U79 ( .A1(a[1]), .A2(b[13]), .ZN(y[29]) );
  OR2_X1 U79bar ( .A1(abar[1]), .A2(bbar[13]), .ZN(ybar[29]) );
  AND2_X1 U80 ( .A1(a[1]), .A2(b[12]), .ZN(y[28]) );
  OR2_X1 U80bar ( .A1(abar[1]), .A2(bbar[12]), .ZN(ybar[28]) );
  AND2_X1 U81 ( .A1(a[1]), .A2(b[11]), .ZN(y[27]) );
  OR2_X1 U81bar ( .A1(abar[1]), .A2(bbar[11]), .ZN(ybar[27]) );
  AND2_X1 U82 ( .A1(a[1]), .A2(b[10]), .ZN(y[26]) );
  OR2_X1 U82bar ( .A1(abar[1]), .A2(bbar[10]), .ZN(ybar[26]) );
  AND2_X1 U83 ( .A1(a[1]), .A2(b[9]), .ZN(y[25]) );
  OR2_X1 U83bar ( .A1(abar[1]), .A2(bbar[9]), .ZN(ybar[25]) );
  AND2_X1 U84 ( .A1(a[15]), .A2(b[15]), .ZN(y[255]) );
  OR2_X1 U84bar ( .A1(abar[15]), .A2(bbar[15]), .ZN(ybar[255]) );
  AND2_X1 U85 ( .A1(a[15]), .A2(b[14]), .ZN(y[254]) );
  OR2_X1 U85bar ( .A1(abar[15]), .A2(bbar[14]), .ZN(ybar[254]) );
  AND2_X1 U86 ( .A1(a[15]), .A2(b[13]), .ZN(y[253]) );
  OR2_X1 U86bar ( .A1(abar[15]), .A2(bbar[13]), .ZN(ybar[253]) );
  AND2_X1 U87 ( .A1(a[15]), .A2(b[12]), .ZN(y[252]) );
  OR2_X1 U87bar ( .A1(abar[15]), .A2(bbar[12]), .ZN(ybar[252]) );
  AND2_X1 U88 ( .A1(a[15]), .A2(b[11]), .ZN(y[251]) );
  OR2_X1 U88bar ( .A1(abar[15]), .A2(bbar[11]), .ZN(ybar[251]) );
  AND2_X1 U89 ( .A1(a[15]), .A2(b[10]), .ZN(y[250]) );
  OR2_X1 U89bar ( .A1(abar[15]), .A2(bbar[10]), .ZN(ybar[250]) );
  AND2_X1 U90 ( .A1(a[1]), .A2(b[8]), .ZN(y[24]) );
  OR2_X1 U90bar ( .A1(abar[1]), .A2(bbar[8]), .ZN(ybar[24]) );
  AND2_X1 U91 ( .A1(a[15]), .A2(b[9]), .ZN(y[249]) );
  OR2_X1 U91bar ( .A1(abar[15]), .A2(bbar[9]), .ZN(ybar[249]) );
  AND2_X1 U92 ( .A1(a[15]), .A2(b[8]), .ZN(y[248]) );
  OR2_X1 U92bar ( .A1(abar[15]), .A2(bbar[8]), .ZN(ybar[248]) );
  AND2_X1 U93 ( .A1(a[15]), .A2(b[7]), .ZN(y[247]) );
  OR2_X1 U93bar ( .A1(abar[15]), .A2(bbar[7]), .ZN(ybar[247]) );
  AND2_X1 U94 ( .A1(a[15]), .A2(b[6]), .ZN(y[246]) );
  OR2_X1 U94bar ( .A1(abar[15]), .A2(bbar[6]), .ZN(ybar[246]) );
  AND2_X1 U95 ( .A1(a[15]), .A2(b[5]), .ZN(y[245]) );
  OR2_X1 U95bar ( .A1(abar[15]), .A2(bbar[5]), .ZN(ybar[245]) );
  AND2_X1 U96 ( .A1(a[15]), .A2(b[4]), .ZN(y[244]) );
  OR2_X1 U96bar ( .A1(abar[15]), .A2(bbar[4]), .ZN(ybar[244]) );
  AND2_X1 U97 ( .A1(a[15]), .A2(b[3]), .ZN(y[243]) );
  OR2_X1 U97bar ( .A1(abar[15]), .A2(bbar[3]), .ZN(ybar[243]) );
  AND2_X1 U98 ( .A1(a[15]), .A2(b[2]), .ZN(y[242]) );
  OR2_X1 U98bar ( .A1(abar[15]), .A2(bbar[2]), .ZN(ybar[242]) );
  AND2_X1 U99 ( .A1(a[15]), .A2(b[1]), .ZN(y[241]) );
  OR2_X1 U99bar ( .A1(abar[15]), .A2(bbar[1]), .ZN(ybar[241]) );
  AND2_X1 U100 ( .A1(a[15]), .A2(b[0]), .ZN(y[240]) );
  OR2_X1 U100bar ( .A1(abar[15]), .A2(bbar[0]), .ZN(ybar[240]) );
  AND2_X1 U101 ( .A1(a[1]), .A2(b[7]), .ZN(y[23]) );
  OR2_X1 U101bar ( .A1(abar[1]), .A2(bbar[7]), .ZN(ybar[23]) );
  AND2_X1 U102 ( .A1(a[14]), .A2(b[15]), .ZN(y[239]) );
  OR2_X1 U102bar ( .A1(abar[14]), .A2(bbar[15]), .ZN(ybar[239]) );
  AND2_X1 U103 ( .A1(a[14]), .A2(b[14]), .ZN(y[238]) );
  OR2_X1 U103bar ( .A1(abar[14]), .A2(bbar[14]), .ZN(ybar[238]) );
  AND2_X1 U104 ( .A1(a[14]), .A2(b[13]), .ZN(y[237]) );
  OR2_X1 U104bar ( .A1(abar[14]), .A2(bbar[13]), .ZN(ybar[237]) );
  AND2_X1 U105 ( .A1(a[14]), .A2(b[12]), .ZN(y[236]) );
  OR2_X1 U105bar ( .A1(abar[14]), .A2(bbar[12]), .ZN(ybar[236]) );
  AND2_X1 U106 ( .A1(a[14]), .A2(b[11]), .ZN(y[235]) );
  OR2_X1 U106bar ( .A1(abar[14]), .A2(bbar[11]), .ZN(ybar[235]) );
  AND2_X1 U107 ( .A1(a[14]), .A2(b[10]), .ZN(y[234]) );
  OR2_X1 U107bar ( .A1(abar[14]), .A2(bbar[10]), .ZN(ybar[234]) );
  AND2_X1 U108 ( .A1(a[14]), .A2(b[9]), .ZN(y[233]) );
  OR2_X1 U108bar ( .A1(abar[14]), .A2(bbar[9]), .ZN(ybar[233]) );
  AND2_X1 U109 ( .A1(a[14]), .A2(b[8]), .ZN(y[232]) );
  OR2_X1 U109bar ( .A1(abar[14]), .A2(bbar[8]), .ZN(ybar[232]) );
  AND2_X1 U110 ( .A1(a[14]), .A2(b[7]), .ZN(y[231]) );
  OR2_X1 U110bar ( .A1(abar[14]), .A2(bbar[7]), .ZN(ybar[231]) );
  AND2_X1 U111 ( .A1(a[14]), .A2(b[6]), .ZN(y[230]) );
  OR2_X1 U111bar ( .A1(abar[14]), .A2(bbar[6]), .ZN(ybar[230]) );
  AND2_X1 U112 ( .A1(a[1]), .A2(b[6]), .ZN(y[22]) );
  OR2_X1 U112bar ( .A1(abar[1]), .A2(bbar[6]), .ZN(ybar[22]) );
  AND2_X1 U113 ( .A1(a[14]), .A2(b[5]), .ZN(y[229]) );
  OR2_X1 U113bar ( .A1(abar[14]), .A2(bbar[5]), .ZN(ybar[229]) );
  AND2_X1 U114 ( .A1(a[14]), .A2(b[4]), .ZN(y[228]) );
  OR2_X1 U114bar ( .A1(abar[14]), .A2(bbar[4]), .ZN(ybar[228]) );
  AND2_X1 U115 ( .A1(a[14]), .A2(b[3]), .ZN(y[227]) );
  OR2_X1 U115bar ( .A1(abar[14]), .A2(bbar[3]), .ZN(ybar[227]) );
  AND2_X1 U116 ( .A1(a[14]), .A2(b[2]), .ZN(y[226]) );
  OR2_X1 U116bar ( .A1(abar[14]), .A2(bbar[2]), .ZN(ybar[226]) );
  AND2_X1 U117 ( .A1(a[14]), .A2(b[1]), .ZN(y[225]) );
  OR2_X1 U117bar ( .A1(abar[14]), .A2(bbar[1]), .ZN(ybar[225]) );
  AND2_X1 U118 ( .A1(a[14]), .A2(b[0]), .ZN(y[224]) );
  OR2_X1 U118bar ( .A1(abar[14]), .A2(bbar[0]), .ZN(ybar[224]) );
  AND2_X1 U119 ( .A1(a[13]), .A2(b[15]), .ZN(y[223]) );
  OR2_X1 U119bar ( .A1(abar[13]), .A2(bbar[15]), .ZN(ybar[223]) );
  AND2_X1 U120 ( .A1(a[13]), .A2(b[14]), .ZN(y[222]) );
  OR2_X1 U120bar ( .A1(abar[13]), .A2(bbar[14]), .ZN(ybar[222]) );
  AND2_X1 U121 ( .A1(a[13]), .A2(b[13]), .ZN(y[221]) );
  OR2_X1 U121bar ( .A1(abar[13]), .A2(bbar[13]), .ZN(ybar[221]) );
  AND2_X1 U122 ( .A1(a[13]), .A2(b[12]), .ZN(y[220]) );
  OR2_X1 U122bar ( .A1(abar[13]), .A2(bbar[12]), .ZN(ybar[220]) );
  AND2_X1 U123 ( .A1(a[1]), .A2(b[5]), .ZN(y[21]) );
  OR2_X1 U123bar ( .A1(abar[1]), .A2(bbar[5]), .ZN(ybar[21]) );
  AND2_X1 U124 ( .A1(a[13]), .A2(b[11]), .ZN(y[219]) );
  OR2_X1 U124bar ( .A1(abar[13]), .A2(bbar[11]), .ZN(ybar[219]) );
  AND2_X1 U125 ( .A1(a[13]), .A2(b[10]), .ZN(y[218]) );
  OR2_X1 U125bar ( .A1(abar[13]), .A2(bbar[10]), .ZN(ybar[218]) );
  AND2_X1 U126 ( .A1(a[13]), .A2(b[9]), .ZN(y[217]) );
  OR2_X1 U126bar ( .A1(abar[13]), .A2(bbar[9]), .ZN(ybar[217]) );
  AND2_X1 U127 ( .A1(a[13]), .A2(b[8]), .ZN(y[216]) );
  OR2_X1 U127bar ( .A1(abar[13]), .A2(bbar[8]), .ZN(ybar[216]) );
  AND2_X1 U128 ( .A1(a[13]), .A2(b[7]), .ZN(y[215]) );
  OR2_X1 U128bar ( .A1(abar[13]), .A2(bbar[7]), .ZN(ybar[215]) );
  AND2_X1 U129 ( .A1(a[13]), .A2(b[6]), .ZN(y[214]) );
  OR2_X1 U129bar ( .A1(abar[13]), .A2(bbar[6]), .ZN(ybar[214]) );
  AND2_X1 U130 ( .A1(a[13]), .A2(b[5]), .ZN(y[213]) );
  OR2_X1 U130bar ( .A1(abar[13]), .A2(bbar[5]), .ZN(ybar[213]) );
  AND2_X1 U131 ( .A1(a[13]), .A2(b[4]), .ZN(y[212]) );
  OR2_X1 U131bar ( .A1(abar[13]), .A2(bbar[4]), .ZN(ybar[212]) );
  AND2_X1 U132 ( .A1(a[13]), .A2(b[3]), .ZN(y[211]) );
  OR2_X1 U132bar ( .A1(abar[13]), .A2(bbar[3]), .ZN(ybar[211]) );
  AND2_X1 U133 ( .A1(a[13]), .A2(b[2]), .ZN(y[210]) );
  OR2_X1 U133bar ( .A1(abar[13]), .A2(bbar[2]), .ZN(ybar[210]) );
  AND2_X1 U134 ( .A1(a[1]), .A2(b[4]), .ZN(y[20]) );
  OR2_X1 U134bar ( .A1(abar[1]), .A2(bbar[4]), .ZN(ybar[20]) );
  AND2_X1 U135 ( .A1(a[13]), .A2(b[1]), .ZN(y[209]) );
  OR2_X1 U135bar ( .A1(abar[13]), .A2(bbar[1]), .ZN(ybar[209]) );
  AND2_X1 U136 ( .A1(a[13]), .A2(b[0]), .ZN(y[208]) );
  OR2_X1 U136bar ( .A1(abar[13]), .A2(bbar[0]), .ZN(ybar[208]) );
  AND2_X1 U137 ( .A1(a[12]), .A2(b[15]), .ZN(y[207]) );
  OR2_X1 U137bar ( .A1(abar[12]), .A2(bbar[15]), .ZN(ybar[207]) );
  AND2_X1 U138 ( .A1(a[12]), .A2(b[14]), .ZN(y[206]) );
  OR2_X1 U138bar ( .A1(abar[12]), .A2(bbar[14]), .ZN(ybar[206]) );
  AND2_X1 U139 ( .A1(a[12]), .A2(b[13]), .ZN(y[205]) );
  OR2_X1 U139bar ( .A1(abar[12]), .A2(bbar[13]), .ZN(ybar[205]) );
  AND2_X1 U140 ( .A1(a[12]), .A2(b[12]), .ZN(y[204]) );
  OR2_X1 U140bar ( .A1(abar[12]), .A2(bbar[12]), .ZN(ybar[204]) );
  AND2_X1 U141 ( .A1(a[12]), .A2(b[11]), .ZN(y[203]) );
  OR2_X1 U141bar ( .A1(abar[12]), .A2(bbar[11]), .ZN(ybar[203]) );
  AND2_X1 U142 ( .A1(a[12]), .A2(b[10]), .ZN(y[202]) );
  OR2_X1 U142bar ( .A1(abar[12]), .A2(bbar[10]), .ZN(ybar[202]) );
  AND2_X1 U143 ( .A1(a[12]), .A2(b[9]), .ZN(y[201]) );
  OR2_X1 U143bar ( .A1(abar[12]), .A2(bbar[9]), .ZN(ybar[201]) );
  AND2_X1 U144 ( .A1(a[12]), .A2(b[8]), .ZN(y[200]) );
  OR2_X1 U144bar ( .A1(abar[12]), .A2(bbar[8]), .ZN(ybar[200]) );
  AND2_X1 U145 ( .A1(b[1]), .A2(a[0]), .ZN(y[1]) );
  OR2_X1 U145bar ( .A1(bbar[1]), .A2(abar[0]), .ZN(ybar[1]) );
  AND2_X1 U146 ( .A1(a[1]), .A2(b[3]), .ZN(y[19]) );
  OR2_X1 U146bar ( .A1(abar[1]), .A2(bbar[3]), .ZN(ybar[19]) );
  AND2_X1 U147 ( .A1(a[12]), .A2(b[7]), .ZN(y[199]) );
  OR2_X1 U147bar ( .A1(abar[12]), .A2(bbar[7]), .ZN(ybar[199]) );
  AND2_X1 U148 ( .A1(a[12]), .A2(b[6]), .ZN(y[198]) );
  OR2_X1 U148bar ( .A1(abar[12]), .A2(bbar[6]), .ZN(ybar[198]) );
  AND2_X1 U149 ( .A1(a[12]), .A2(b[5]), .ZN(y[197]) );
  OR2_X1 U149bar ( .A1(abar[12]), .A2(bbar[5]), .ZN(ybar[197]) );
  AND2_X1 U150 ( .A1(a[12]), .A2(b[4]), .ZN(y[196]) );
  OR2_X1 U150bar ( .A1(abar[12]), .A2(bbar[4]), .ZN(ybar[196]) );
  AND2_X1 U151 ( .A1(a[12]), .A2(b[3]), .ZN(y[195]) );
  OR2_X1 U151bar ( .A1(abar[12]), .A2(bbar[3]), .ZN(ybar[195]) );
  AND2_X1 U152 ( .A1(a[12]), .A2(b[2]), .ZN(y[194]) );
  OR2_X1 U152bar ( .A1(abar[12]), .A2(bbar[2]), .ZN(ybar[194]) );
  AND2_X1 U153 ( .A1(a[12]), .A2(b[1]), .ZN(y[193]) );
  OR2_X1 U153bar ( .A1(abar[12]), .A2(bbar[1]), .ZN(ybar[193]) );
  AND2_X1 U154 ( .A1(a[12]), .A2(b[0]), .ZN(y[192]) );
  OR2_X1 U154bar ( .A1(abar[12]), .A2(bbar[0]), .ZN(ybar[192]) );
  AND2_X1 U155 ( .A1(a[11]), .A2(b[15]), .ZN(y[191]) );
  OR2_X1 U155bar ( .A1(abar[11]), .A2(bbar[15]), .ZN(ybar[191]) );
  AND2_X1 U156 ( .A1(a[11]), .A2(b[14]), .ZN(y[190]) );
  OR2_X1 U156bar ( .A1(abar[11]), .A2(bbar[14]), .ZN(ybar[190]) );
  AND2_X1 U157 ( .A1(a[1]), .A2(b[2]), .ZN(y[18]) );
  OR2_X1 U157bar ( .A1(abar[1]), .A2(bbar[2]), .ZN(ybar[18]) );
  AND2_X1 U158 ( .A1(a[11]), .A2(b[13]), .ZN(y[189]) );
  OR2_X1 U158bar ( .A1(abar[11]), .A2(bbar[13]), .ZN(ybar[189]) );
  AND2_X1 U159 ( .A1(a[11]), .A2(b[12]), .ZN(y[188]) );
  OR2_X1 U159bar ( .A1(abar[11]), .A2(bbar[12]), .ZN(ybar[188]) );
  AND2_X1 U160 ( .A1(a[11]), .A2(b[11]), .ZN(y[187]) );
  OR2_X1 U160bar ( .A1(abar[11]), .A2(bbar[11]), .ZN(ybar[187]) );
  AND2_X1 U161 ( .A1(a[11]), .A2(b[10]), .ZN(y[186]) );
  OR2_X1 U161bar ( .A1(abar[11]), .A2(bbar[10]), .ZN(ybar[186]) );
  AND2_X1 U162 ( .A1(a[11]), .A2(b[9]), .ZN(y[185]) );
  OR2_X1 U162bar ( .A1(abar[11]), .A2(bbar[9]), .ZN(ybar[185]) );
  AND2_X1 U163 ( .A1(a[11]), .A2(b[8]), .ZN(y[184]) );
  OR2_X1 U163bar ( .A1(abar[11]), .A2(bbar[8]), .ZN(ybar[184]) );
  AND2_X1 U164 ( .A1(a[11]), .A2(b[7]), .ZN(y[183]) );
  OR2_X1 U164bar ( .A1(abar[11]), .A2(bbar[7]), .ZN(ybar[183]) );
  AND2_X1 U165 ( .A1(a[11]), .A2(b[6]), .ZN(y[182]) );
  OR2_X1 U165bar ( .A1(abar[11]), .A2(bbar[6]), .ZN(ybar[182]) );
  AND2_X1 U166 ( .A1(a[11]), .A2(b[5]), .ZN(y[181]) );
  OR2_X1 U166bar ( .A1(abar[11]), .A2(bbar[5]), .ZN(ybar[181]) );
  AND2_X1 U167 ( .A1(a[11]), .A2(b[4]), .ZN(y[180]) );
  OR2_X1 U167bar ( .A1(abar[11]), .A2(bbar[4]), .ZN(ybar[180]) );
  AND2_X1 U168 ( .A1(a[1]), .A2(b[1]), .ZN(y[17]) );
  OR2_X1 U168bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[17]) );
  AND2_X1 U169 ( .A1(a[11]), .A2(b[3]), .ZN(y[179]) );
  OR2_X1 U169bar ( .A1(abar[11]), .A2(bbar[3]), .ZN(ybar[179]) );
  AND2_X1 U170 ( .A1(a[11]), .A2(b[2]), .ZN(y[178]) );
  OR2_X1 U170bar ( .A1(abar[11]), .A2(bbar[2]), .ZN(ybar[178]) );
  AND2_X1 U171 ( .A1(a[11]), .A2(b[1]), .ZN(y[177]) );
  OR2_X1 U171bar ( .A1(abar[11]), .A2(bbar[1]), .ZN(ybar[177]) );
  AND2_X1 U172 ( .A1(a[11]), .A2(b[0]), .ZN(y[176]) );
  OR2_X1 U172bar ( .A1(abar[11]), .A2(bbar[0]), .ZN(ybar[176]) );
  AND2_X1 U173 ( .A1(a[10]), .A2(b[15]), .ZN(y[175]) );
  OR2_X1 U173bar ( .A1(abar[10]), .A2(bbar[15]), .ZN(ybar[175]) );
  AND2_X1 U174 ( .A1(a[10]), .A2(b[14]), .ZN(y[174]) );
  OR2_X1 U174bar ( .A1(abar[10]), .A2(bbar[14]), .ZN(ybar[174]) );
  AND2_X1 U175 ( .A1(a[10]), .A2(b[13]), .ZN(y[173]) );
  OR2_X1 U175bar ( .A1(abar[10]), .A2(bbar[13]), .ZN(ybar[173]) );
  AND2_X1 U176 ( .A1(a[10]), .A2(b[12]), .ZN(y[172]) );
  OR2_X1 U176bar ( .A1(abar[10]), .A2(bbar[12]), .ZN(ybar[172]) );
  AND2_X1 U177 ( .A1(a[10]), .A2(b[11]), .ZN(y[171]) );
  OR2_X1 U177bar ( .A1(abar[10]), .A2(bbar[11]), .ZN(ybar[171]) );
  AND2_X1 U178 ( .A1(a[10]), .A2(b[10]), .ZN(y[170]) );
  OR2_X1 U178bar ( .A1(abar[10]), .A2(bbar[10]), .ZN(ybar[170]) );
  AND2_X1 U179 ( .A1(a[1]), .A2(b[0]), .ZN(y[16]) );
  OR2_X1 U179bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[16]) );
  AND2_X1 U180 ( .A1(a[10]), .A2(b[9]), .ZN(y[169]) );
  OR2_X1 U180bar ( .A1(abar[10]), .A2(bbar[9]), .ZN(ybar[169]) );
  AND2_X1 U181 ( .A1(a[10]), .A2(b[8]), .ZN(y[168]) );
  OR2_X1 U181bar ( .A1(abar[10]), .A2(bbar[8]), .ZN(ybar[168]) );
  AND2_X1 U182 ( .A1(a[10]), .A2(b[7]), .ZN(y[167]) );
  OR2_X1 U182bar ( .A1(abar[10]), .A2(bbar[7]), .ZN(ybar[167]) );
  AND2_X1 U183 ( .A1(a[10]), .A2(b[6]), .ZN(y[166]) );
  OR2_X1 U183bar ( .A1(abar[10]), .A2(bbar[6]), .ZN(ybar[166]) );
  AND2_X1 U184 ( .A1(a[10]), .A2(b[5]), .ZN(y[165]) );
  OR2_X1 U184bar ( .A1(abar[10]), .A2(bbar[5]), .ZN(ybar[165]) );
  AND2_X1 U185 ( .A1(a[10]), .A2(b[4]), .ZN(y[164]) );
  OR2_X1 U185bar ( .A1(abar[10]), .A2(bbar[4]), .ZN(ybar[164]) );
  AND2_X1 U186 ( .A1(a[10]), .A2(b[3]), .ZN(y[163]) );
  OR2_X1 U186bar ( .A1(abar[10]), .A2(bbar[3]), .ZN(ybar[163]) );
  AND2_X1 U187 ( .A1(a[10]), .A2(b[2]), .ZN(y[162]) );
  OR2_X1 U187bar ( .A1(abar[10]), .A2(bbar[2]), .ZN(ybar[162]) );
  AND2_X1 U188 ( .A1(a[10]), .A2(b[1]), .ZN(y[161]) );
  OR2_X1 U188bar ( .A1(abar[10]), .A2(bbar[1]), .ZN(ybar[161]) );
  AND2_X1 U189 ( .A1(a[10]), .A2(b[0]), .ZN(y[160]) );
  OR2_X1 U189bar ( .A1(abar[10]), .A2(bbar[0]), .ZN(ybar[160]) );
  AND2_X1 U190 ( .A1(b[15]), .A2(a[0]), .ZN(y[15]) );
  OR2_X1 U190bar ( .A1(bbar[15]), .A2(abar[0]), .ZN(ybar[15]) );
  AND2_X1 U191 ( .A1(a[9]), .A2(b[15]), .ZN(y[159]) );
  OR2_X1 U191bar ( .A1(abar[9]), .A2(bbar[15]), .ZN(ybar[159]) );
  AND2_X1 U192 ( .A1(a[9]), .A2(b[14]), .ZN(y[158]) );
  OR2_X1 U192bar ( .A1(abar[9]), .A2(bbar[14]), .ZN(ybar[158]) );
  AND2_X1 U193 ( .A1(a[9]), .A2(b[13]), .ZN(y[157]) );
  OR2_X1 U193bar ( .A1(abar[9]), .A2(bbar[13]), .ZN(ybar[157]) );
  AND2_X1 U194 ( .A1(a[9]), .A2(b[12]), .ZN(y[156]) );
  OR2_X1 U194bar ( .A1(abar[9]), .A2(bbar[12]), .ZN(ybar[156]) );
  AND2_X1 U195 ( .A1(a[9]), .A2(b[11]), .ZN(y[155]) );
  OR2_X1 U195bar ( .A1(abar[9]), .A2(bbar[11]), .ZN(ybar[155]) );
  AND2_X1 U196 ( .A1(a[9]), .A2(b[10]), .ZN(y[154]) );
  OR2_X1 U196bar ( .A1(abar[9]), .A2(bbar[10]), .ZN(ybar[154]) );
  AND2_X1 U197 ( .A1(a[9]), .A2(b[9]), .ZN(y[153]) );
  OR2_X1 U197bar ( .A1(abar[9]), .A2(bbar[9]), .ZN(ybar[153]) );
  AND2_X1 U198 ( .A1(a[9]), .A2(b[8]), .ZN(y[152]) );
  OR2_X1 U198bar ( .A1(abar[9]), .A2(bbar[8]), .ZN(ybar[152]) );
  AND2_X1 U199 ( .A1(a[9]), .A2(b[7]), .ZN(y[151]) );
  OR2_X1 U199bar ( .A1(abar[9]), .A2(bbar[7]), .ZN(ybar[151]) );
  AND2_X1 U200 ( .A1(a[9]), .A2(b[6]), .ZN(y[150]) );
  OR2_X1 U200bar ( .A1(abar[9]), .A2(bbar[6]), .ZN(ybar[150]) );
  AND2_X1 U201 ( .A1(b[14]), .A2(a[0]), .ZN(y[14]) );
  OR2_X1 U201bar ( .A1(bbar[14]), .A2(abar[0]), .ZN(ybar[14]) );
  AND2_X1 U202 ( .A1(a[9]), .A2(b[5]), .ZN(y[149]) );
  OR2_X1 U202bar ( .A1(abar[9]), .A2(bbar[5]), .ZN(ybar[149]) );
  AND2_X1 U203 ( .A1(a[9]), .A2(b[4]), .ZN(y[148]) );
  OR2_X1 U203bar ( .A1(abar[9]), .A2(bbar[4]), .ZN(ybar[148]) );
  AND2_X1 U204 ( .A1(a[9]), .A2(b[3]), .ZN(y[147]) );
  OR2_X1 U204bar ( .A1(abar[9]), .A2(bbar[3]), .ZN(ybar[147]) );
  AND2_X1 U205 ( .A1(a[9]), .A2(b[2]), .ZN(y[146]) );
  OR2_X1 U205bar ( .A1(abar[9]), .A2(bbar[2]), .ZN(ybar[146]) );
  AND2_X1 U206 ( .A1(a[9]), .A2(b[1]), .ZN(y[145]) );
  OR2_X1 U206bar ( .A1(abar[9]), .A2(bbar[1]), .ZN(ybar[145]) );
  AND2_X1 U207 ( .A1(a[9]), .A2(b[0]), .ZN(y[144]) );
  OR2_X1 U207bar ( .A1(abar[9]), .A2(bbar[0]), .ZN(ybar[144]) );
  AND2_X1 U208 ( .A1(a[8]), .A2(b[15]), .ZN(y[143]) );
  OR2_X1 U208bar ( .A1(abar[8]), .A2(bbar[15]), .ZN(ybar[143]) );
  AND2_X1 U209 ( .A1(a[8]), .A2(b[14]), .ZN(y[142]) );
  OR2_X1 U209bar ( .A1(abar[8]), .A2(bbar[14]), .ZN(ybar[142]) );
  AND2_X1 U210 ( .A1(a[8]), .A2(b[13]), .ZN(y[141]) );
  OR2_X1 U210bar ( .A1(abar[8]), .A2(bbar[13]), .ZN(ybar[141]) );
  AND2_X1 U211 ( .A1(a[8]), .A2(b[12]), .ZN(y[140]) );
  OR2_X1 U211bar ( .A1(abar[8]), .A2(bbar[12]), .ZN(ybar[140]) );
  AND2_X1 U212 ( .A1(b[13]), .A2(a[0]), .ZN(y[13]) );
  OR2_X1 U212bar ( .A1(bbar[13]), .A2(abar[0]), .ZN(ybar[13]) );
  AND2_X1 U213 ( .A1(a[8]), .A2(b[11]), .ZN(y[139]) );
  OR2_X1 U213bar ( .A1(abar[8]), .A2(bbar[11]), .ZN(ybar[139]) );
  AND2_X1 U214 ( .A1(a[8]), .A2(b[10]), .ZN(y[138]) );
  OR2_X1 U214bar ( .A1(abar[8]), .A2(bbar[10]), .ZN(ybar[138]) );
  AND2_X1 U215 ( .A1(a[8]), .A2(b[9]), .ZN(y[137]) );
  OR2_X1 U215bar ( .A1(abar[8]), .A2(bbar[9]), .ZN(ybar[137]) );
  AND2_X1 U216 ( .A1(a[8]), .A2(b[8]), .ZN(y[136]) );
  OR2_X1 U216bar ( .A1(abar[8]), .A2(bbar[8]), .ZN(ybar[136]) );
  AND2_X1 U217 ( .A1(a[8]), .A2(b[7]), .ZN(y[135]) );
  OR2_X1 U217bar ( .A1(abar[8]), .A2(bbar[7]), .ZN(ybar[135]) );
  AND2_X1 U218 ( .A1(a[8]), .A2(b[6]), .ZN(y[134]) );
  OR2_X1 U218bar ( .A1(abar[8]), .A2(bbar[6]), .ZN(ybar[134]) );
  AND2_X1 U219 ( .A1(a[8]), .A2(b[5]), .ZN(y[133]) );
  OR2_X1 U219bar ( .A1(abar[8]), .A2(bbar[5]), .ZN(ybar[133]) );
  AND2_X1 U220 ( .A1(a[8]), .A2(b[4]), .ZN(y[132]) );
  OR2_X1 U220bar ( .A1(abar[8]), .A2(bbar[4]), .ZN(ybar[132]) );
  AND2_X1 U221 ( .A1(a[8]), .A2(b[3]), .ZN(y[131]) );
  OR2_X1 U221bar ( .A1(abar[8]), .A2(bbar[3]), .ZN(ybar[131]) );
  AND2_X1 U222 ( .A1(a[8]), .A2(b[2]), .ZN(y[130]) );
  OR2_X1 U222bar ( .A1(abar[8]), .A2(bbar[2]), .ZN(ybar[130]) );
  AND2_X1 U223 ( .A1(b[12]), .A2(a[0]), .ZN(y[12]) );
  OR2_X1 U223bar ( .A1(bbar[12]), .A2(abar[0]), .ZN(ybar[12]) );
  AND2_X1 U224 ( .A1(a[8]), .A2(b[1]), .ZN(y[129]) );
  OR2_X1 U224bar ( .A1(abar[8]), .A2(bbar[1]), .ZN(ybar[129]) );
  AND2_X1 U225 ( .A1(a[8]), .A2(b[0]), .ZN(y[128]) );
  OR2_X1 U225bar ( .A1(abar[8]), .A2(bbar[0]), .ZN(ybar[128]) );
  AND2_X1 U226 ( .A1(a[7]), .A2(b[15]), .ZN(y[127]) );
  OR2_X1 U226bar ( .A1(abar[7]), .A2(bbar[15]), .ZN(ybar[127]) );
  AND2_X1 U227 ( .A1(a[7]), .A2(b[14]), .ZN(y[126]) );
  OR2_X1 U227bar ( .A1(abar[7]), .A2(bbar[14]), .ZN(ybar[126]) );
  AND2_X1 U228 ( .A1(a[7]), .A2(b[13]), .ZN(y[125]) );
  OR2_X1 U228bar ( .A1(abar[7]), .A2(bbar[13]), .ZN(ybar[125]) );
  AND2_X1 U229 ( .A1(a[7]), .A2(b[12]), .ZN(y[124]) );
  OR2_X1 U229bar ( .A1(abar[7]), .A2(bbar[12]), .ZN(ybar[124]) );
  AND2_X1 U230 ( .A1(a[7]), .A2(b[11]), .ZN(y[123]) );
  OR2_X1 U230bar ( .A1(abar[7]), .A2(bbar[11]), .ZN(ybar[123]) );
  AND2_X1 U231 ( .A1(a[7]), .A2(b[10]), .ZN(y[122]) );
  OR2_X1 U231bar ( .A1(abar[7]), .A2(bbar[10]), .ZN(ybar[122]) );
  AND2_X1 U232 ( .A1(a[7]), .A2(b[9]), .ZN(y[121]) );
  OR2_X1 U232bar ( .A1(abar[7]), .A2(bbar[9]), .ZN(ybar[121]) );
  AND2_X1 U233 ( .A1(a[7]), .A2(b[8]), .ZN(y[120]) );
  OR2_X1 U233bar ( .A1(abar[7]), .A2(bbar[8]), .ZN(ybar[120]) );
  AND2_X1 U234 ( .A1(b[11]), .A2(a[0]), .ZN(y[11]) );
  OR2_X1 U234bar ( .A1(bbar[11]), .A2(abar[0]), .ZN(ybar[11]) );
  AND2_X1 U235 ( .A1(a[7]), .A2(b[7]), .ZN(y[119]) );
  OR2_X1 U235bar ( .A1(abar[7]), .A2(bbar[7]), .ZN(ybar[119]) );
  AND2_X1 U236 ( .A1(a[7]), .A2(b[6]), .ZN(y[118]) );
  OR2_X1 U236bar ( .A1(abar[7]), .A2(bbar[6]), .ZN(ybar[118]) );
  AND2_X1 U237 ( .A1(a[7]), .A2(b[5]), .ZN(y[117]) );
  OR2_X1 U237bar ( .A1(abar[7]), .A2(bbar[5]), .ZN(ybar[117]) );
  AND2_X1 U238 ( .A1(a[7]), .A2(b[4]), .ZN(y[116]) );
  OR2_X1 U238bar ( .A1(abar[7]), .A2(bbar[4]), .ZN(ybar[116]) );
  AND2_X1 U239 ( .A1(a[7]), .A2(b[3]), .ZN(y[115]) );
  OR2_X1 U239bar ( .A1(abar[7]), .A2(bbar[3]), .ZN(ybar[115]) );
  AND2_X1 U240 ( .A1(a[7]), .A2(b[2]), .ZN(y[114]) );
  OR2_X1 U240bar ( .A1(abar[7]), .A2(bbar[2]), .ZN(ybar[114]) );
  AND2_X1 U241 ( .A1(a[7]), .A2(b[1]), .ZN(y[113]) );
  OR2_X1 U241bar ( .A1(abar[7]), .A2(bbar[1]), .ZN(ybar[113]) );
  AND2_X1 U242 ( .A1(a[7]), .A2(b[0]), .ZN(y[112]) );
  OR2_X1 U242bar ( .A1(abar[7]), .A2(bbar[0]), .ZN(ybar[112]) );
  AND2_X1 U243 ( .A1(b[15]), .A2(a[6]), .ZN(y[111]) );
  OR2_X1 U243bar ( .A1(bbar[15]), .A2(abar[6]), .ZN(ybar[111]) );
  AND2_X1 U244 ( .A1(b[14]), .A2(a[6]), .ZN(y[110]) );
  OR2_X1 U244bar ( .A1(bbar[14]), .A2(abar[6]), .ZN(ybar[110]) );
  AND2_X1 U245 ( .A1(b[10]), .A2(a[0]), .ZN(y[10]) );
  OR2_X1 U245bar ( .A1(bbar[10]), .A2(abar[0]), .ZN(ybar[10]) );
  AND2_X1 U246 ( .A1(b[13]), .A2(a[6]), .ZN(y[109]) );
  OR2_X1 U246bar ( .A1(bbar[13]), .A2(abar[6]), .ZN(ybar[109]) );
  AND2_X1 U247 ( .A1(b[12]), .A2(a[6]), .ZN(y[108]) );
  OR2_X1 U247bar ( .A1(bbar[12]), .A2(abar[6]), .ZN(ybar[108]) );
  AND2_X1 U248 ( .A1(b[11]), .A2(a[6]), .ZN(y[107]) );
  OR2_X1 U248bar ( .A1(bbar[11]), .A2(abar[6]), .ZN(ybar[107]) );
  AND2_X1 U249 ( .A1(b[10]), .A2(a[6]), .ZN(y[106]) );
  OR2_X1 U249bar ( .A1(bbar[10]), .A2(abar[6]), .ZN(ybar[106]) );
  AND2_X1 U250 ( .A1(a[6]), .A2(b[9]), .ZN(y[105]) );
  OR2_X1 U250bar ( .A1(abar[6]), .A2(bbar[9]), .ZN(ybar[105]) );
  AND2_X1 U251 ( .A1(b[8]), .A2(a[6]), .ZN(y[104]) );
  OR2_X1 U251bar ( .A1(bbar[8]), .A2(abar[6]), .ZN(ybar[104]) );
  AND2_X1 U252 ( .A1(b[7]), .A2(a[6]), .ZN(y[103]) );
  OR2_X1 U252bar ( .A1(bbar[7]), .A2(abar[6]), .ZN(ybar[103]) );
  AND2_X1 U253 ( .A1(b[6]), .A2(a[6]), .ZN(y[102]) );
  OR2_X1 U253bar ( .A1(bbar[6]), .A2(abar[6]), .ZN(ybar[102]) );
  AND2_X1 U254 ( .A1(b[5]), .A2(a[6]), .ZN(y[101]) );
  OR2_X1 U254bar ( .A1(bbar[5]), .A2(abar[6]), .ZN(ybar[101]) );
  AND2_X1 U255 ( .A1(b[4]), .A2(a[6]), .ZN(y[100]) );
  OR2_X1 U255bar ( .A1(bbar[4]), .A2(abar[6]), .ZN(ybar[100]) );
  AND2_X1 U256 ( .A1(b[0]), .A2(a[0]), .ZN(y[0]) );
  OR2_X1 U256bar ( .A1(bbar[0]), .A2(abar[0]), .ZN(ybar[0]) );
endmodule

module decode_11 ( in, inbar, out, outbar );

  input wire [7:0] in;
  input wire [7:0] inbar;
//input_done

  output wire [255:0] out;
  output wire [255:0] outbar;
//output_done

  wire [15:0] level1;
  wire [31:0] level2;
  wire [15:0] level1bar;
  wire [31:0] level2bar;
//wire_done

  CD2_44 cd_l1_1 ( .a(in[1]), .abar(inbar[1]), .b(in[0]), .bbar(inbar[0]), .y(level1[3:0]), .ybar(level1bar[3:0]) );
  CD2_43 cd_l1_2 ( .a(in[3]), .abar(inbar[3]), .b(in[2]), .bbar(inbar[2]), .y(level1[7:4]), .ybar(level1bar[7:4]) );
  CD2_42 cd_l1_3 ( .a(in[5]), .abar(inbar[5]), .b(in[4]), .bbar(inbar[4]), .y(level1[11:8]), .ybar(level1bar[11:8]) );
  CD2_41 cd_l1_4 ( .a(in[7]), .abar(inbar[7]), .b(in[6]), .bbar(inbar[6]), .y(level1[15:12]), .ybar(level1bar[15:12]) );

  CD4_22 cd_l2_1 ( .a(level1[7:4]), .abar(level1bar[7:4]), .b(level1[3:0]), .bbar(level1bar[3:0]), 
        .y(level2[15:0]), .ybar(level2bar[15:0]) );
  CD4_21 cd_l2_2 ( .a(level1[15:12]), .abar(level1bar[15:12]), .b(level1[11:8]), .bbar(level1bar[11:8]), 
        .y(level2[31:16]), .ybar(level2bar[31:16]) );
  CD16_11 cd_l3 ( .a(level2[31:16]), .abar(level2bar[31:16]), .b(level2[15:0]), .bbar(level2bar[15:0]), 
        .y(out), .ybar(outbar) );
endmodule

module encode_11 ( in, inbar, out, outbar );

  input wire [255:0] in;
  input wire [255:0] inbar;
//input_done

  output wire [7:0] out;
  output wire [7:0] outbar;
//output_done

  wire in_81;
  wire in_80;
  wire in_79;
  wire in_78;
  wire in_77;
  wire in_76;
  wire in_75;
  wire in_74;
  wire in_73;
  wire in_72;
  wire in_71;
  wire in_70;
  wire in_69;
  wire in_68;
  wire in_67;
  wire in_66;
  wire in_65;
  wire in_64;
  wire in_63;
  wire in_62;
  wire in_61;
  wire in_60;
  wire in_59;
  wire in_58;
  wire in_57;
  wire in_56;
  wire in_55;
  wire in_54;
  wire in_53;
  wire in_52;
  wire in_51;
  wire in_50;
  wire in_49;
  wire in_48;
  wire in_47;
  wire in_46;
  wire in_45;
  wire in_44;
  wire in_43;
  wire in_42;
  wire in_41;
  wire in_40;
  wire in_39;
  wire in_38;
  wire in_37;
  wire in_36;
  wire in_35;
  wire in_34;
  wire in_33;
  wire in_32;
  wire in_31;
  wire in_30;
  wire in_29;
  wire in_28;
  wire in_27;
  wire in_26;
  wire in_25;
  wire in_24;
  wire in_23;
  wire in_22;
  wire in_21;
  wire in_20;
  wire in_19;
  wire in_18;
  wire in_17;
  wire in_16;
  wire in_15;
  wire in_14;
  wire in_13;
  wire in_12;
  wire in_11;
  wire in_10;
  wire in_9;
  wire in_8;
  wire in_7;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_3;
  wire in_2;
  wire in_1;
  wire in_0;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire in_81bar;
  wire in_80bar;
  wire in_79bar;
  wire in_78bar;
  wire in_77bar;
  wire in_76bar;
  wire in_75bar;
  wire in_74bar;
  wire in_73bar;
  wire in_72bar;
  wire in_71bar;
  wire in_70bar;
  wire in_69bar;
  wire in_68bar;
  wire in_67bar;
  wire in_66bar;
  wire in_65bar;
  wire in_64bar;
  wire in_63bar;
  wire in_62bar;
  wire in_61bar;
  wire in_60bar;
  wire in_59bar;
  wire in_58bar;
  wire in_57bar;
  wire in_56bar;
  wire in_55bar;
  wire in_54bar;
  wire in_53bar;
  wire in_52bar;
  wire in_51bar;
  wire in_50bar;
  wire in_49bar;
  wire in_48bar;
  wire in_47bar;
  wire in_46bar;
  wire in_45bar;
  wire in_44bar;
  wire in_43bar;
  wire in_42bar;
  wire in_41bar;
  wire in_40bar;
  wire in_39bar;
  wire in_38bar;
  wire in_37bar;
  wire in_36bar;
  wire in_35bar;
  wire in_34bar;
  wire in_33bar;
  wire in_32bar;
  wire in_31bar;
  wire in_30bar;
  wire in_29bar;
  wire in_28bar;
  wire in_27bar;
  wire in_26bar;
  wire in_25bar;
  wire in_24bar;
  wire in_23bar;
  wire in_22bar;
  wire in_21bar;
  wire in_20bar;
  wire in_19bar;
  wire in_18bar;
  wire in_17bar;
  wire in_16bar;
  wire in_15bar;
  wire in_14bar;
  wire in_13bar;
  wire in_12bar;
  wire in_11bar;
  wire in_10bar;
  wire in_9bar;
  wire in_8bar;
  wire in_7bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_3bar;
  wire in_2bar;
  wire in_1bar;
  wire in_0bar;
  wire n487bar;
  wire n488bar;
  wire n489bar;
  wire n490bar;
  wire n491bar;
  wire n492bar;
  wire n493bar;
  wire n494bar;
  wire n495bar;
  wire n496bar;
  wire n497bar;
  wire n498bar;
  wire n499bar;
  wire n500bar;
  wire n501bar;
  wire n502bar;
  wire n503bar;
  wire n504bar;
  wire n505bar;
  wire n506bar;
  wire n507bar;
  wire n508bar;
  wire n509bar;
  wire n510bar;
  wire n511bar;
  wire n512bar;
  wire n513bar;
  wire n514bar;
  wire n515bar;
  wire n516bar;
  wire n517bar;
  wire n518bar;
  wire n519bar;
  wire n520bar;
  wire n521bar;
  wire n522bar;
  wire n523bar;
  wire n524bar;
  wire n525bar;
  wire n526bar;
  wire n527bar;
  wire n528bar;
  wire n529bar;
  wire n530bar;
  wire n531bar;
  wire n532bar;
  wire n533bar;
  wire n534bar;
  wire n535bar;
  wire n536bar;
  wire n537bar;
  wire n538bar;
  wire n539bar;
  wire n540bar;
  wire n541bar;
  wire n542bar;
  wire n543bar;
  wire n544bar;
  wire n545bar;
  wire n546bar;
  wire n547bar;
  wire n548bar;
  wire n549bar;
  wire n550bar;
  wire n551bar;
  wire n552bar;
  wire n553bar;
  wire n554bar;
  wire n555bar;
  wire n556bar;
  wire n557bar;
  wire n558bar;
  wire n559bar;
  wire n560bar;
  wire n561bar;
  wire n562bar;
  wire n563bar;
  wire n564bar;
  wire n565bar;
  wire n566bar;
  wire n567bar;
  wire n568bar;
  wire n569bar;
  wire n570bar;
  wire n571bar;
  wire n572bar;
  wire n573bar;
  wire n574bar;
  wire n575bar;
  wire n576bar;
  wire n577bar;
  wire n578bar;
  wire n579bar;
  wire n580bar;
  wire n581bar;
  wire n582bar;
  wire n583bar;
  wire n584bar;
  wire n585bar;
  wire n586bar;
  wire n587bar;
  wire n588bar;
  wire n589bar;
  wire n590bar;
  wire n591bar;
  wire n592bar;
  wire n593bar;
  wire n594bar;
  wire n595bar;
  wire n596bar;
  wire n597bar;
  wire n598bar;
  wire n599bar;
  wire n600bar;
  wire n601bar;
  wire n602bar;
  wire n603bar;
  wire n604bar;
  wire n605bar;
  wire n606bar;
  wire n607bar;
  wire n608bar;
  wire n609bar;
  wire n610bar;
  wire n611bar;
  wire n612bar;
  wire n613bar;
  wire n614bar;
  wire n615bar;
  wire n616bar;
  wire n617bar;
  wire n618bar;
  wire n619bar;
  wire n620bar;
  wire n621bar;
  wire n622bar;
  wire n623bar;
  wire n624bar;
  wire n625bar;
  wire n626bar;
  wire n627bar;
  wire n628bar;
  wire n629bar;
  wire n630bar;
  wire n631bar;
  wire n632bar;
  wire n633bar;
  wire n634bar;
  wire n635bar;
  wire n636bar;
  wire n637bar;
  wire n638bar;
  wire n639bar;
  wire n640bar;
  wire n641bar;
  wire n642bar;
  wire n643bar;
  wire n644bar;
  wire n645bar;
  wire n646bar;
  wire n647bar;
  wire n648bar;
  wire n649bar;
  wire n650bar;
  wire n651bar;
  wire n652bar;
  wire n653bar;
  wire n654bar;
  wire n655bar;
  wire n656bar;
  wire n657bar;
  wire n658bar;
  wire n659bar;
  wire n660bar;
  wire n661bar;
  wire n662bar;
  wire n663bar;
  wire n664bar;
  wire n665bar;
  wire n666bar;
  wire n667bar;
  wire n668bar;
  wire n669bar;
  wire n670bar;
  wire n671bar;
  wire n672bar;
  wire n673bar;
  wire n674bar;
  wire n675bar;
  wire n676bar;
  wire n677bar;
  wire n678bar;
  wire n679bar;
  wire n680bar;
  wire n681bar;
  wire n682bar;
  wire n683bar;
  wire n684bar;
  wire n685bar;
  wire n686bar;
  wire n687bar;
  wire n688bar;
  wire n689bar;
  wire n690bar;
  wire n691bar;
  wire n692bar;
  wire n693bar;
  wire n694bar;
  wire n695bar;
  wire n696bar;
  wire n697bar;
  wire n698bar;
  wire n699bar;
  wire n700bar;
  wire n701bar;
  wire n702bar;
  wire n703bar;
  wire n704bar;
  wire n705bar;
  wire n706bar;
  wire n707bar;
  wire n708bar;
  wire n709bar;
  wire n710bar;
  wire n711bar;
  wire n712bar;
  wire n713bar;
  wire n714bar;
  wire n715bar;
  wire n716bar;
  wire n717bar;
  wire n718bar;
  wire n719bar;
  wire n720bar;
  wire n721bar;
  wire n722bar;
  wire n723bar;
  wire n724bar;
  wire n725bar;
  wire n726bar;
  wire n727bar;
  wire n728bar;
  wire n729bar;
  wire n730bar;
  wire n731bar;
  wire n732bar;
  wire n733bar;
  wire n734bar;
  wire n735bar;
  wire n736bar;
  wire n737bar;
  wire n738bar;
  wire n739bar;
  wire n740bar;
  wire n741bar;
  wire n742bar;
  wire n743bar;
  wire n744bar;
  wire n745bar;
  wire n746bar;
  wire n747bar;
  wire n748bar;
  wire n749bar;
  wire n750bar;
  wire n751bar;
  wire n752bar;
  wire n753bar;
  wire n754bar;
  wire n755bar;
  wire n756bar;
  wire n757bar;
  wire n758bar;
  wire n759bar;
  wire n760bar;
  wire n761bar;
  wire n762bar;
  wire n763bar;
  wire n764bar;
  wire n765bar;
  wire n766bar;
  wire n767bar;
  wire n768bar;
  wire n769bar;
  wire n770bar;
  wire n771bar;
  wire n772bar;
  wire n773bar;
  wire n774bar;
  wire n775bar;
  wire n776bar;
  wire n777bar;
  wire n778bar;
  wire n779bar;
  wire n780bar;
  wire n781bar;
  wire n782bar;
  wire n783bar;
  wire n784bar;
  wire n785bar;
  wire n786bar;
  wire n787bar;
  wire n788bar;
  wire n789bar;
  wire n790bar;
  wire n791bar;
  wire n792bar;
  wire n793bar;
  wire n794bar;
  wire n795bar;
  wire n796bar;
  wire n797bar;
  wire n798bar;
  wire n799bar;
  wire n800bar;
  wire n801bar;
  wire n802bar;
  wire n803bar;
  wire n804bar;
  wire n805bar;
  wire n806bar;
  wire n807bar;
  wire n808bar;
  wire n809bar;
  wire n810bar;
  wire n811bar;
  wire n812bar;
  wire n813bar;
  wire n814bar;
  wire n815bar;
  wire n816bar;
  wire n817bar;
  wire n818bar;
  wire n819bar;
  wire n820bar;
  wire n821bar;
  wire n822bar;
  wire n823bar;
  wire n824bar;
  wire n825bar;
  wire n826bar;
  wire n827bar;
  wire n828bar;
  wire n829bar;
  wire n830bar;
  wire n831bar;
  wire n832bar;
  wire n833bar;
  wire n834bar;
  wire n835bar;
  wire n836bar;
  wire n837bar;
  wire n838bar;
  wire n839bar;
  wire n840bar;
  wire n841bar;
  wire n842bar;
  wire n843bar;
  wire n844bar;
  wire n845bar;
  wire n846bar;
  wire n847bar;
  wire n848bar;
  wire n849bar;
  wire n850bar;
  wire n851bar;
  wire n852bar;
  wire n853bar;
  wire n854bar;
  wire n855bar;
  wire n856bar;
  wire n857bar;
  wire n858bar;
  wire n859bar;
  wire n860bar;
  wire n861bar;
  wire n862bar;
  wire n863bar;
  wire n864bar;
  wire n865bar;
  wire n866bar;
  wire n867bar;
  wire n868bar;
  wire n869bar;
  wire n870bar;
  wire n871bar;
  wire n872bar;
  wire n873bar;
  wire n874bar;
  wire n875bar;
  wire n876bar;
  wire n877bar;
  wire n878bar;
  wire n879bar;
  wire n880bar;
  wire n881bar;
  wire n882bar;
  wire n883bar;
  wire n884bar;
  wire n885bar;
  wire n886bar;
  wire n887bar;
  wire n888bar;
  wire n889bar;
  wire n890bar;
  wire n891bar;
  wire n892bar;
  wire n893bar;
  wire n894bar;
  wire n895bar;
  wire n896bar;
  wire n897bar;
  wire n898bar;
  wire n899bar;
  wire n900bar;
  wire n901bar;
  wire n902bar;
  wire n903bar;
  wire n904bar;
  wire n905bar;
  wire n906bar;
  wire n907bar;
  wire n908bar;
  wire n909bar;
  wire n910bar;
  wire n911bar;
  wire n912bar;
  wire n913bar;
  wire n914bar;
  wire n915bar;
  wire n916bar;
  wire n917bar;
  wire n918bar;
  wire n919bar;
  wire n920bar;
  wire n921bar;
  wire n922bar;
  wire n923bar;
  wire n924bar;
  wire n925bar;
  wire n926bar;
  wire n927bar;
  wire n928bar;
  wire n929bar;
  wire n930bar;
  wire n931bar;
  wire n932bar;
  wire n933bar;
  wire n934bar;
  wire n935bar;
  wire n936bar;
  wire n937bar;
  wire n938bar;
  wire n939bar;
  wire n940bar;
  wire n941bar;
  wire n942bar;
  wire n943bar;
  wire n944bar;
  wire n945bar;
  wire n946bar;
  wire n947bar;
  wire n948bar;
  wire n949bar;
  wire n950bar;
  wire n951bar;
  wire n952bar;
  wire n953bar;
  wire n954bar;
  wire n955bar;
  wire n956bar;
  wire n957bar;
  wire n958bar;
  wire n959bar;
  wire n960bar;
  wire n961bar;
  wire n962bar;
  wire n963bar;
  wire n964bar;
  wire n965bar;
  wire n966bar;
  wire n967bar;
  wire n968bar;
  wire n969bar;
  wire n970bar;
  wire n971bar;
  wire n972bar;
//wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];
  assign in_81bar = inbar[81];
  assign in_80bar = inbar[80];
  assign in_79bar = inbar[79];
  assign in_78bar = inbar[78];
  assign in_77bar = inbar[77];
  assign in_76bar = inbar[76];
  assign in_75bar = inbar[75];
  assign in_74bar = inbar[74];
  assign in_73bar = inbar[73];
  assign in_72bar = inbar[72];
  assign in_71bar = inbar[71];
  assign in_70bar = inbar[70];
  assign in_69bar = inbar[69];
  assign in_68bar = inbar[68];
  assign in_67bar = inbar[67];
  assign in_66bar = inbar[66];
  assign in_65bar = inbar[65];
  assign in_64bar = inbar[64];
  assign in_63bar = inbar[63];
  assign in_62bar = inbar[62];
  assign in_61bar = inbar[61];
  assign in_60bar = inbar[60];
  assign in_59bar = inbar[59];
  assign in_58bar = inbar[58];
  assign in_57bar = inbar[57];
  assign in_56bar = inbar[56];
  assign in_55bar = inbar[55];
  assign in_54bar = inbar[54];
  assign in_53bar = inbar[53];
  assign in_52bar = inbar[52];
  assign in_51bar = inbar[51];
  assign in_50bar = inbar[50];
  assign in_49bar = inbar[49];
  assign in_48bar = inbar[48];
  assign in_47bar = inbar[47];
  assign in_46bar = inbar[46];
  assign in_45bar = inbar[45];
  assign in_44bar = inbar[44];
  assign in_43bar = inbar[43];
  assign in_42bar = inbar[42];
  assign in_41bar = inbar[41];
  assign in_40bar = inbar[40];
  assign in_39bar = inbar[39];
  assign in_38bar = inbar[38];
  assign in_37bar = inbar[37];
  assign in_36bar = inbar[36];
  assign in_35bar = inbar[35];
  assign in_34bar = inbar[34];
  assign in_33bar = inbar[33];
  assign in_32bar = inbar[32];
  assign in_31bar = inbar[31];
  assign in_30bar = inbar[30];
  assign in_29bar = inbar[29];
  assign in_28bar = inbar[28];
  assign in_27bar = inbar[27];
  assign in_26bar = inbar[26];
  assign in_25bar = inbar[25];
  assign in_24bar = inbar[24];
  assign in_23bar = inbar[23];
  assign in_22bar = inbar[22];
  assign in_21bar = inbar[21];
  assign in_20bar = inbar[20];
  assign in_19bar = inbar[19];
  assign in_18bar = inbar[18];
  assign in_17bar = inbar[17];
  assign in_16bar = inbar[16];
  assign in_15bar = inbar[15];
  assign in_14bar = inbar[14];
  assign in_13bar = inbar[13];
  assign in_12bar = inbar[12];
  assign in_11bar = inbar[11];
  assign in_10bar = inbar[10];
  assign in_9bar = inbar[9];
  assign in_8bar = inbar[8];
  assign in_7bar = inbar[7];
  assign in_6bar = inbar[6];
  assign in_5bar = inbar[5];
  assign in_4bar = inbar[4];
  assign in_3bar = inbar[3];
  assign in_2bar = inbar[2];
  assign in_1bar = inbar[1];
  assign in_0bar = inbar[0];
//assign_done

  OR2_X1 U1 ( .A1(n972), .A2(n971), .ZN(out[7]) );
  AND2_X1 U1bar ( .A1(n972bar), .A2(n971bar), .ZN(outbar[7]) );
  OR2_X1 U2 ( .A1(n970), .A2(n969), .ZN(n971) );
  AND2_X1 U2bar ( .A1(n970bar), .A2(n969bar), .ZN(n971bar) );
  OR2_X1 U3 ( .A1(n968), .A2(n967), .ZN(n969) );
  AND2_X1 U3bar ( .A1(n968bar), .A2(n967bar), .ZN(n969bar) );
  OR2_X1 U4 ( .A1(n966), .A2(n965), .ZN(n967) );
  AND2_X1 U4bar ( .A1(n966bar), .A2(n965bar), .ZN(n967bar) );
  OR2_X1 U5 ( .A1(n964), .A2(n963), .ZN(n968) );
  AND2_X1 U5bar ( .A1(n964bar), .A2(n963bar), .ZN(n968bar) );
  OR2_X1 U6 ( .A1(in[116]), .A2(n962), .ZN(n963) );
  AND2_X1 U6bar ( .A1(inbar[116]), .A2(n962bar), .ZN(n963bar) );
  OR2_X1 U7 ( .A1(n961), .A2(n960), .ZN(n970) );
  AND2_X1 U7bar ( .A1(n961bar), .A2(n960bar), .ZN(n970bar) );
  OR2_X1 U8 ( .A1(in[150]), .A2(in[127]), .ZN(n960) );
  AND2_X1 U8bar ( .A1(inbar[150]), .A2(inbar[127]), .ZN(n960bar) );
  OR2_X1 U9 ( .A1(in[160]), .A2(n959), .ZN(n961) );
  AND2_X1 U9bar ( .A1(inbar[160]), .A2(n959bar), .ZN(n961bar) );
  OR2_X1 U10 ( .A1(in[252]), .A2(in[168]), .ZN(n959) );
  AND2_X1 U10bar ( .A1(inbar[252]), .A2(inbar[168]), .ZN(n959bar) );
  OR2_X1 U11 ( .A1(n958), .A2(n957), .ZN(n972) );
  AND2_X1 U11bar ( .A1(n958bar), .A2(n957bar), .ZN(n972bar) );
  OR2_X1 U12 ( .A1(n956), .A2(n955), .ZN(n957) );
  AND2_X1 U12bar ( .A1(n956bar), .A2(n955bar), .ZN(n957bar) );
  OR2_X1 U13 ( .A1(in_17), .A2(in[96]), .ZN(n955) );
  AND2_X1 U13bar ( .A1(in_17bar), .A2(inbar[96]), .ZN(n955bar) );
  OR2_X1 U14 ( .A1(in_23), .A2(n954), .ZN(n956) );
  AND2_X1 U14bar ( .A1(in_23bar), .A2(n954bar), .ZN(n956bar) );
  OR2_X1 U15 ( .A1(in_31), .A2(in_26), .ZN(n954) );
  AND2_X1 U15bar ( .A1(in_31bar), .A2(in_26bar), .ZN(n954bar) );
  OR2_X1 U16 ( .A1(n953), .A2(n952), .ZN(n958) );
  AND2_X1 U16bar ( .A1(n953bar), .A2(n952bar), .ZN(n958bar) );
  OR2_X1 U17 ( .A1(in_58), .A2(in_4), .ZN(n952) );
  AND2_X1 U17bar ( .A1(in_58bar), .A2(in_4bar), .ZN(n952bar) );
  OR2_X1 U18 ( .A1(in_59), .A2(n951), .ZN(n953) );
  AND2_X1 U18bar ( .A1(in_59bar), .A2(n951bar), .ZN(n953bar) );
  OR2_X1 U19 ( .A1(in_71), .A2(in_62), .ZN(n951) );
  AND2_X1 U19bar ( .A1(in_71bar), .A2(in_62bar), .ZN(n951bar) );
  OR2_X1 U20 ( .A1(n950), .A2(n949), .ZN(out[6]) );
  AND2_X1 U20bar ( .A1(n950bar), .A2(n949bar), .ZN(outbar[6]) );
  OR2_X1 U21 ( .A1(n948), .A2(n947), .ZN(n949) );
  AND2_X1 U21bar ( .A1(n948bar), .A2(n947bar), .ZN(n949bar) );
  OR2_X1 U22 ( .A1(n946), .A2(n945), .ZN(n947) );
  AND2_X1 U22bar ( .A1(n946bar), .A2(n945bar), .ZN(n947bar) );
  OR2_X1 U23 ( .A1(n944), .A2(n943), .ZN(n945) );
  AND2_X1 U23bar ( .A1(n944bar), .A2(n943bar), .ZN(n945bar) );
  OR2_X1 U24 ( .A1(n942), .A2(n941), .ZN(n946) );
  AND2_X1 U24bar ( .A1(n942bar), .A2(n941bar), .ZN(n946bar) );
  OR2_X1 U25 ( .A1(in[101]), .A2(n940), .ZN(n941) );
  AND2_X1 U25bar ( .A1(inbar[101]), .A2(n940bar), .ZN(n941bar) );
  OR2_X1 U26 ( .A1(n939), .A2(n938), .ZN(n948) );
  AND2_X1 U26bar ( .A1(n939bar), .A2(n938bar), .ZN(n948bar) );
  OR2_X1 U27 ( .A1(in[114]), .A2(in[104]), .ZN(n938) );
  AND2_X1 U27bar ( .A1(inbar[114]), .A2(inbar[104]), .ZN(n938bar) );
  OR2_X1 U28 ( .A1(in[128]), .A2(n937), .ZN(n939) );
  AND2_X1 U28bar ( .A1(inbar[128]), .A2(n937bar), .ZN(n939bar) );
  OR2_X1 U29 ( .A1(in[136]), .A2(in[134]), .ZN(n937) );
  AND2_X1 U29bar ( .A1(inbar[136]), .A2(inbar[134]), .ZN(n937bar) );
  OR2_X1 U30 ( .A1(n936), .A2(n935), .ZN(n950) );
  AND2_X1 U30bar ( .A1(n936bar), .A2(n935bar), .ZN(n950bar) );
  OR2_X1 U31 ( .A1(n934), .A2(n933), .ZN(n935) );
  AND2_X1 U31bar ( .A1(n934bar), .A2(n933bar), .ZN(n935bar) );
  OR2_X1 U32 ( .A1(in[177]), .A2(in[164]), .ZN(n933) );
  AND2_X1 U32bar ( .A1(inbar[177]), .A2(inbar[164]), .ZN(n933bar) );
  OR2_X1 U33 ( .A1(in[212]), .A2(n932), .ZN(n934) );
  AND2_X1 U33bar ( .A1(inbar[212]), .A2(n932bar), .ZN(n934bar) );
  OR2_X1 U34 ( .A1(in[248]), .A2(in[221]), .ZN(n932) );
  AND2_X1 U34bar ( .A1(inbar[248]), .A2(inbar[221]), .ZN(n932bar) );
  OR2_X1 U35 ( .A1(n931), .A2(n930), .ZN(n936) );
  AND2_X1 U35bar ( .A1(n931bar), .A2(n930bar), .ZN(n936bar) );
  OR2_X1 U36 ( .A1(in_18), .A2(in[93]), .ZN(n930) );
  AND2_X1 U36bar ( .A1(in_18bar), .A2(inbar[93]), .ZN(n930bar) );
  OR2_X1 U37 ( .A1(in_31), .A2(n929), .ZN(n931) );
  AND2_X1 U37bar ( .A1(in_31bar), .A2(n929bar), .ZN(n931bar) );
  OR2_X1 U38 ( .A1(in_7), .A2(in_39), .ZN(n929) );
  AND2_X1 U38bar ( .A1(in_7bar), .A2(in_39bar), .ZN(n929bar) );
  OR2_X1 U39 ( .A1(n928), .A2(n927), .ZN(out[5]) );
  AND2_X1 U39bar ( .A1(n928bar), .A2(n927bar), .ZN(outbar[5]) );
  OR2_X1 U40 ( .A1(n926), .A2(n925), .ZN(n927) );
  AND2_X1 U40bar ( .A1(n926bar), .A2(n925bar), .ZN(n927bar) );
  OR2_X1 U41 ( .A1(n924), .A2(n923), .ZN(n925) );
  AND2_X1 U41bar ( .A1(n924bar), .A2(n923bar), .ZN(n925bar) );
  OR2_X1 U42 ( .A1(n922), .A2(n921), .ZN(n923) );
  AND2_X1 U42bar ( .A1(n922bar), .A2(n921bar), .ZN(n923bar) );
  OR2_X1 U43 ( .A1(n940), .A2(n920), .ZN(n924) );
  AND2_X1 U43bar ( .A1(n940bar), .A2(n920bar), .ZN(n924bar) );
  OR2_X1 U44 ( .A1(in[111]), .A2(n919), .ZN(n920) );
  AND2_X1 U44bar ( .A1(inbar[111]), .A2(n919bar), .ZN(n920bar) );
  OR2_X1 U45 ( .A1(n918), .A2(n917), .ZN(n940) );
  AND2_X1 U45bar ( .A1(n918bar), .A2(n917bar), .ZN(n940bar) );
  OR2_X1 U46 ( .A1(n916), .A2(n915), .ZN(n917) );
  AND2_X1 U46bar ( .A1(n916bar), .A2(n915bar), .ZN(n917bar) );
  OR2_X1 U47 ( .A1(n914), .A2(n913), .ZN(n915) );
  AND2_X1 U47bar ( .A1(n914bar), .A2(n913bar), .ZN(n915bar) );
  OR2_X1 U48 ( .A1(in[140]), .A2(in[131]), .ZN(n913) );
  AND2_X1 U48bar ( .A1(inbar[140]), .A2(inbar[131]), .ZN(n913bar) );
  OR2_X1 U49 ( .A1(in[160]), .A2(in[144]), .ZN(n914) );
  AND2_X1 U49bar ( .A1(inbar[160]), .A2(inbar[144]), .ZN(n914bar) );
  OR2_X1 U50 ( .A1(n912), .A2(n911), .ZN(n916) );
  AND2_X1 U50bar ( .A1(n912bar), .A2(n911bar), .ZN(n916bar) );
  OR2_X1 U51 ( .A1(in[179]), .A2(in[174]), .ZN(n911) );
  AND2_X1 U51bar ( .A1(inbar[179]), .A2(inbar[174]), .ZN(n911bar) );
  OR2_X1 U52 ( .A1(in[188]), .A2(in[184]), .ZN(n912) );
  AND2_X1 U52bar ( .A1(inbar[188]), .A2(inbar[184]), .ZN(n912bar) );
  OR2_X1 U53 ( .A1(n910), .A2(n909), .ZN(n918) );
  AND2_X1 U53bar ( .A1(n910bar), .A2(n909bar), .ZN(n918bar) );
  OR2_X1 U54 ( .A1(n908), .A2(n907), .ZN(n909) );
  AND2_X1 U54bar ( .A1(n908bar), .A2(n907bar), .ZN(n909bar) );
  OR2_X1 U55 ( .A1(in[216]), .A2(in[200]), .ZN(n907) );
  AND2_X1 U55bar ( .A1(inbar[216]), .A2(inbar[200]), .ZN(n907bar) );
  OR2_X1 U56 ( .A1(in[228]), .A2(in[224]), .ZN(n908) );
  AND2_X1 U56bar ( .A1(inbar[228]), .A2(inbar[224]), .ZN(n908bar) );
  OR2_X1 U57 ( .A1(n906), .A2(n905), .ZN(n910) );
  AND2_X1 U57bar ( .A1(n906bar), .A2(n905bar), .ZN(n910bar) );
  OR2_X1 U58 ( .A1(in[247]), .A2(in[235]), .ZN(n905) );
  AND2_X1 U58bar ( .A1(inbar[247]), .A2(inbar[235]), .ZN(n905bar) );
  OR2_X1 U59 ( .A1(in_42), .A2(in[83]), .ZN(n906) );
  AND2_X1 U59bar ( .A1(in_42bar), .A2(inbar[83]), .ZN(n906bar) );
  OR2_X1 U60 ( .A1(n904), .A2(n903), .ZN(n926) );
  AND2_X1 U60bar ( .A1(n904bar), .A2(n903bar), .ZN(n926bar) );
  OR2_X1 U61 ( .A1(in[166]), .A2(in[123]), .ZN(n903) );
  AND2_X1 U61bar ( .A1(inbar[166]), .A2(inbar[123]), .ZN(n903bar) );
  OR2_X1 U62 ( .A1(in[170]), .A2(n902), .ZN(n904) );
  AND2_X1 U62bar ( .A1(inbar[170]), .A2(n902bar), .ZN(n904bar) );
  OR2_X1 U63 ( .A1(in[194]), .A2(in[183]), .ZN(n902) );
  AND2_X1 U63bar ( .A1(inbar[194]), .A2(inbar[183]), .ZN(n902bar) );
  OR2_X1 U64 ( .A1(n901), .A2(n900), .ZN(n928) );
  AND2_X1 U64bar ( .A1(n901bar), .A2(n900bar), .ZN(n928bar) );
  OR2_X1 U65 ( .A1(n899), .A2(n898), .ZN(n900) );
  AND2_X1 U65bar ( .A1(n899bar), .A2(n898bar), .ZN(n900bar) );
  OR2_X1 U66 ( .A1(in[241]), .A2(in[238]), .ZN(n898) );
  AND2_X1 U66bar ( .A1(inbar[241]), .A2(inbar[238]), .ZN(n898bar) );
  OR2_X1 U67 ( .A1(in[250]), .A2(n897), .ZN(n899) );
  AND2_X1 U67bar ( .A1(inbar[250]), .A2(n897bar), .ZN(n899bar) );
  OR2_X1 U68 ( .A1(in_24), .A2(in[84]), .ZN(n897) );
  AND2_X1 U68bar ( .A1(in_24bar), .A2(inbar[84]), .ZN(n897bar) );
  OR2_X1 U69 ( .A1(n896), .A2(n895), .ZN(n901) );
  AND2_X1 U69bar ( .A1(n896bar), .A2(n895bar), .ZN(n901bar) );
  OR2_X1 U70 ( .A1(in_41), .A2(in_29), .ZN(n895) );
  AND2_X1 U70bar ( .A1(in_41bar), .A2(in_29bar), .ZN(n895bar) );
  OR2_X1 U71 ( .A1(in_66), .A2(n894), .ZN(n896) );
  AND2_X1 U71bar ( .A1(in_66bar), .A2(n894bar), .ZN(n896bar) );
  OR2_X1 U72 ( .A1(in_76), .A2(in_71), .ZN(n894) );
  AND2_X1 U72bar ( .A1(in_76bar), .A2(in_71bar), .ZN(n894bar) );
  OR2_X1 U73 ( .A1(n893), .A2(n892), .ZN(out[4]) );
  AND2_X1 U73bar ( .A1(n893bar), .A2(n892bar), .ZN(outbar[4]) );
  OR2_X1 U74 ( .A1(n891), .A2(n890), .ZN(n892) );
  AND2_X1 U74bar ( .A1(n891bar), .A2(n890bar), .ZN(n892bar) );
  OR2_X1 U75 ( .A1(n889), .A2(n888), .ZN(n890) );
  AND2_X1 U75bar ( .A1(n889bar), .A2(n888bar), .ZN(n890bar) );
  OR2_X1 U76 ( .A1(n922), .A2(n887), .ZN(n888) );
  AND2_X1 U76bar ( .A1(n922bar), .A2(n887bar), .ZN(n888bar) );
  OR2_X1 U77 ( .A1(n886), .A2(n885), .ZN(n922) );
  AND2_X1 U77bar ( .A1(n886bar), .A2(n885bar), .ZN(n922bar) );
  OR2_X1 U78 ( .A1(n884), .A2(n883), .ZN(n885) );
  AND2_X1 U78bar ( .A1(n884bar), .A2(n883bar), .ZN(n885bar) );
  OR2_X1 U79 ( .A1(n882), .A2(n881), .ZN(n883) );
  AND2_X1 U79bar ( .A1(n882bar), .A2(n881bar), .ZN(n883bar) );
  OR2_X1 U80 ( .A1(in[118]), .A2(in[109]), .ZN(n881) );
  AND2_X1 U80bar ( .A1(inbar[118]), .A2(inbar[109]), .ZN(n881bar) );
  OR2_X1 U81 ( .A1(in[139]), .A2(in[120]), .ZN(n882) );
  AND2_X1 U81bar ( .A1(inbar[139]), .A2(inbar[120]), .ZN(n882bar) );
  OR2_X1 U82 ( .A1(n880), .A2(n879), .ZN(n884) );
  AND2_X1 U82bar ( .A1(n880bar), .A2(n879bar), .ZN(n884bar) );
  OR2_X1 U83 ( .A1(in[198]), .A2(in[154]), .ZN(n879) );
  AND2_X1 U83bar ( .A1(inbar[198]), .A2(inbar[154]), .ZN(n879bar) );
  OR2_X1 U84 ( .A1(in[210]), .A2(in[205]), .ZN(n880) );
  AND2_X1 U84bar ( .A1(inbar[210]), .A2(inbar[205]), .ZN(n880bar) );
  OR2_X1 U85 ( .A1(n878), .A2(n877), .ZN(n886) );
  AND2_X1 U85bar ( .A1(n878bar), .A2(n877bar), .ZN(n886bar) );
  OR2_X1 U86 ( .A1(n876), .A2(n875), .ZN(n877) );
  AND2_X1 U86bar ( .A1(n876bar), .A2(n875bar), .ZN(n877bar) );
  OR2_X1 U87 ( .A1(in[219]), .A2(in[217]), .ZN(n875) );
  AND2_X1 U87bar ( .A1(inbar[219]), .A2(inbar[217]), .ZN(n875bar) );
  OR2_X1 U88 ( .A1(in[86]), .A2(in[252]), .ZN(n876) );
  AND2_X1 U88bar ( .A1(inbar[86]), .A2(inbar[252]), .ZN(n876bar) );
  OR2_X1 U89 ( .A1(n874), .A2(n873), .ZN(n878) );
  AND2_X1 U89bar ( .A1(n874bar), .A2(n873bar), .ZN(n878bar) );
  OR2_X1 U90 ( .A1(in_40), .A2(in[91]), .ZN(n873) );
  AND2_X1 U90bar ( .A1(in_40bar), .A2(inbar[91]), .ZN(n873bar) );
  OR2_X1 U91 ( .A1(in_8), .A2(in_46), .ZN(n874) );
  AND2_X1 U91bar ( .A1(in_8bar), .A2(in_46bar), .ZN(n874bar) );
  OR2_X1 U92 ( .A1(n872), .A2(n871), .ZN(n889) );
  AND2_X1 U92bar ( .A1(n872bar), .A2(n871bar), .ZN(n889bar) );
  OR2_X1 U93 ( .A1(in[117]), .A2(n943), .ZN(n871) );
  AND2_X1 U93bar ( .A1(inbar[117]), .A2(n943bar), .ZN(n871bar) );
  OR2_X1 U94 ( .A1(n870), .A2(n869), .ZN(n943) );
  AND2_X1 U94bar ( .A1(n870bar), .A2(n869bar), .ZN(n943bar) );
  OR2_X1 U95 ( .A1(n868), .A2(n867), .ZN(n869) );
  AND2_X1 U95bar ( .A1(n868bar), .A2(n867bar), .ZN(n869bar) );
  OR2_X1 U96 ( .A1(n866), .A2(n865), .ZN(n867) );
  AND2_X1 U96bar ( .A1(n866bar), .A2(n865bar), .ZN(n867bar) );
  OR2_X1 U97 ( .A1(n864), .A2(n863), .ZN(n865) );
  AND2_X1 U97bar ( .A1(n864bar), .A2(n863bar), .ZN(n865bar) );
  OR2_X1 U98 ( .A1(in[108]), .A2(n919), .ZN(n866) );
  AND2_X1 U98bar ( .A1(inbar[108]), .A2(n919bar), .ZN(n866bar) );
  OR2_X1 U99 ( .A1(n862), .A2(n861), .ZN(n919) );
  AND2_X1 U99bar ( .A1(n862bar), .A2(n861bar), .ZN(n919bar) );
  OR2_X1 U100 ( .A1(n860), .A2(n859), .ZN(n861) );
  AND2_X1 U100bar ( .A1(n860bar), .A2(n859bar), .ZN(n861bar) );
  OR2_X1 U101 ( .A1(n858), .A2(n857), .ZN(n859) );
  AND2_X1 U101bar ( .A1(n858bar), .A2(n857bar), .ZN(n859bar) );
  OR2_X1 U102 ( .A1(in[119]), .A2(in[105]), .ZN(n857) );
  AND2_X1 U102bar ( .A1(inbar[119]), .A2(inbar[105]), .ZN(n857bar) );
  OR2_X1 U103 ( .A1(in[186]), .A2(in[175]), .ZN(n858) );
  AND2_X1 U103bar ( .A1(inbar[186]), .A2(inbar[175]), .ZN(n858bar) );
  OR2_X1 U104 ( .A1(n856), .A2(n855), .ZN(n860) );
  AND2_X1 U104bar ( .A1(n856bar), .A2(n855bar), .ZN(n860bar) );
  OR2_X1 U105 ( .A1(in[202]), .A2(in[193]), .ZN(n855) );
  AND2_X1 U105bar ( .A1(inbar[202]), .A2(inbar[193]), .ZN(n855bar) );
  OR2_X1 U106 ( .A1(in[225]), .A2(in[208]), .ZN(n856) );
  AND2_X1 U106bar ( .A1(inbar[225]), .A2(inbar[208]), .ZN(n856bar) );
  OR2_X1 U107 ( .A1(n854), .A2(n853), .ZN(n862) );
  AND2_X1 U107bar ( .A1(n854bar), .A2(n853bar), .ZN(n862bar) );
  OR2_X1 U108 ( .A1(n852), .A2(n851), .ZN(n853) );
  AND2_X1 U108bar ( .A1(n852bar), .A2(n851bar), .ZN(n853bar) );
  OR2_X1 U109 ( .A1(in_1), .A2(in[85]), .ZN(n851) );
  AND2_X1 U109bar ( .A1(in_1bar), .A2(inbar[85]), .ZN(n851bar) );
  OR2_X1 U110 ( .A1(in_23), .A2(in_19), .ZN(n852) );
  AND2_X1 U110bar ( .A1(in_23bar), .A2(in_19bar), .ZN(n852bar) );
  OR2_X1 U111 ( .A1(n850), .A2(n849), .ZN(n854) );
  AND2_X1 U111bar ( .A1(n850bar), .A2(n849bar), .ZN(n854bar) );
  OR2_X1 U112 ( .A1(in_43), .A2(in_33), .ZN(n849) );
  AND2_X1 U112bar ( .A1(in_43bar), .A2(in_33bar), .ZN(n849bar) );
  OR2_X1 U113 ( .A1(in_63), .A2(in_44), .ZN(n850) );
  AND2_X1 U113bar ( .A1(in_63bar), .A2(in_44bar), .ZN(n850bar) );
  OR2_X1 U114 ( .A1(n848), .A2(n847), .ZN(n868) );
  AND2_X1 U114bar ( .A1(n848bar), .A2(n847bar), .ZN(n868bar) );
  OR2_X1 U115 ( .A1(in[141]), .A2(in[112]), .ZN(n847) );
  AND2_X1 U115bar ( .A1(inbar[141]), .A2(inbar[112]), .ZN(n847bar) );
  OR2_X1 U116 ( .A1(in[147]), .A2(n846), .ZN(n848) );
  AND2_X1 U116bar ( .A1(inbar[147]), .A2(n846bar), .ZN(n848bar) );
  OR2_X1 U117 ( .A1(in[181]), .A2(in[167]), .ZN(n846) );
  AND2_X1 U117bar ( .A1(inbar[181]), .A2(inbar[167]), .ZN(n846bar) );
  OR2_X1 U118 ( .A1(n845), .A2(n844), .ZN(n870) );
  AND2_X1 U118bar ( .A1(n845bar), .A2(n844bar), .ZN(n870bar) );
  OR2_X1 U119 ( .A1(n843), .A2(n842), .ZN(n844) );
  AND2_X1 U119bar ( .A1(n843bar), .A2(n842bar), .ZN(n844bar) );
  OR2_X1 U120 ( .A1(in[229]), .A2(in[201]), .ZN(n842) );
  AND2_X1 U120bar ( .A1(inbar[229]), .A2(inbar[201]), .ZN(n842bar) );
  OR2_X1 U121 ( .A1(in[237]), .A2(n841), .ZN(n843) );
  AND2_X1 U121bar ( .A1(inbar[237]), .A2(n841bar), .ZN(n843bar) );
  OR2_X1 U122 ( .A1(in[94]), .A2(in[253]), .ZN(n841) );
  AND2_X1 U122bar ( .A1(inbar[94]), .A2(inbar[253]), .ZN(n841bar) );
  OR2_X1 U123 ( .A1(n840), .A2(n839), .ZN(n845) );
  AND2_X1 U123bar ( .A1(n840bar), .A2(n839bar), .ZN(n845bar) );
  OR2_X1 U124 ( .A1(in_21), .A2(in[96]), .ZN(n839) );
  AND2_X1 U124bar ( .A1(in_21bar), .A2(inbar[96]), .ZN(n839bar) );
  OR2_X1 U125 ( .A1(in_25), .A2(n838), .ZN(n840) );
  AND2_X1 U125bar ( .A1(in_25bar), .A2(n838bar), .ZN(n840bar) );
  OR2_X1 U126 ( .A1(in_81), .A2(in_45), .ZN(n838) );
  AND2_X1 U126bar ( .A1(in_81bar), .A2(in_45bar), .ZN(n838bar) );
  OR2_X1 U127 ( .A1(n837), .A2(n836), .ZN(n891) );
  AND2_X1 U127bar ( .A1(n837bar), .A2(n836bar), .ZN(n891bar) );
  OR2_X1 U128 ( .A1(in[142]), .A2(in[124]), .ZN(n836) );
  AND2_X1 U128bar ( .A1(inbar[142]), .A2(inbar[124]), .ZN(n836bar) );
  OR2_X1 U129 ( .A1(in[150]), .A2(n835), .ZN(n837) );
  AND2_X1 U129bar ( .A1(inbar[150]), .A2(n835bar), .ZN(n837bar) );
  OR2_X1 U130 ( .A1(in[172]), .A2(in[155]), .ZN(n835) );
  AND2_X1 U130bar ( .A1(inbar[172]), .A2(inbar[155]), .ZN(n835bar) );
  OR2_X1 U131 ( .A1(n834), .A2(n833), .ZN(n893) );
  AND2_X1 U131bar ( .A1(n834bar), .A2(n833bar), .ZN(n893bar) );
  OR2_X1 U132 ( .A1(n832), .A2(n831), .ZN(n833) );
  AND2_X1 U132bar ( .A1(n832bar), .A2(n831bar), .ZN(n833bar) );
  OR2_X1 U133 ( .A1(in[196]), .A2(in[173]), .ZN(n831) );
  AND2_X1 U133bar ( .A1(inbar[196]), .A2(inbar[173]), .ZN(n831bar) );
  OR2_X1 U134 ( .A1(in[222]), .A2(n830), .ZN(n832) );
  AND2_X1 U134bar ( .A1(inbar[222]), .A2(n830bar), .ZN(n832bar) );
  OR2_X1 U135 ( .A1(in[227]), .A2(in[226]), .ZN(n830) );
  AND2_X1 U135bar ( .A1(inbar[227]), .A2(inbar[226]), .ZN(n830bar) );
  OR2_X1 U136 ( .A1(n829), .A2(n828), .ZN(n834) );
  AND2_X1 U136bar ( .A1(n829bar), .A2(n828bar), .ZN(n834bar) );
  OR2_X1 U137 ( .A1(in[249]), .A2(in[231]), .ZN(n828) );
  AND2_X1 U137bar ( .A1(inbar[249]), .A2(inbar[231]), .ZN(n828bar) );
  OR2_X1 U138 ( .A1(in_28), .A2(n827), .ZN(n829) );
  AND2_X1 U138bar ( .A1(in_28bar), .A2(n827bar), .ZN(n829bar) );
  OR2_X1 U139 ( .A1(in_52), .A2(in_47), .ZN(n827) );
  AND2_X1 U139bar ( .A1(in_52bar), .A2(in_47bar), .ZN(n827bar) );
  OR2_X1 U140 ( .A1(n826), .A2(n825), .ZN(out[3]) );
  AND2_X1 U140bar ( .A1(n826bar), .A2(n825bar), .ZN(outbar[3]) );
  OR2_X1 U141 ( .A1(n824), .A2(n823), .ZN(n825) );
  AND2_X1 U141bar ( .A1(n824bar), .A2(n823bar), .ZN(n825bar) );
  OR2_X1 U142 ( .A1(n822), .A2(n821), .ZN(n823) );
  AND2_X1 U142bar ( .A1(n822bar), .A2(n821bar), .ZN(n823bar) );
  OR2_X1 U143 ( .A1(n820), .A2(n819), .ZN(n821) );
  AND2_X1 U143bar ( .A1(n820bar), .A2(n819bar), .ZN(n821bar) );
  OR2_X1 U144 ( .A1(n964), .A2(n818), .ZN(n822) );
  AND2_X1 U144bar ( .A1(n964bar), .A2(n818bar), .ZN(n822bar) );
  OR2_X1 U145 ( .A1(in[118]), .A2(n817), .ZN(n818) );
  AND2_X1 U145bar ( .A1(inbar[118]), .A2(n817bar), .ZN(n818bar) );
  OR2_X1 U146 ( .A1(n816), .A2(n815), .ZN(n964) );
  AND2_X1 U146bar ( .A1(n816bar), .A2(n815bar), .ZN(n964bar) );
  OR2_X1 U147 ( .A1(n814), .A2(n813), .ZN(n815) );
  AND2_X1 U147bar ( .A1(n814bar), .A2(n813bar), .ZN(n815bar) );
  OR2_X1 U148 ( .A1(n812), .A2(n811), .ZN(n813) );
  AND2_X1 U148bar ( .A1(n812bar), .A2(n811bar), .ZN(n813bar) );
  OR2_X1 U149 ( .A1(in[122]), .A2(in[111]), .ZN(n811) );
  AND2_X1 U149bar ( .A1(inbar[122]), .A2(inbar[111]), .ZN(n811bar) );
  OR2_X1 U150 ( .A1(in[154]), .A2(in[151]), .ZN(n812) );
  AND2_X1 U150bar ( .A1(inbar[154]), .A2(inbar[151]), .ZN(n812bar) );
  OR2_X1 U151 ( .A1(n810), .A2(n809), .ZN(n814) );
  AND2_X1 U151bar ( .A1(n810bar), .A2(n809bar), .ZN(n814bar) );
  OR2_X1 U152 ( .A1(in[187]), .A2(in[177]), .ZN(n809) );
  AND2_X1 U152bar ( .A1(inbar[187]), .A2(inbar[177]), .ZN(n809bar) );
  OR2_X1 U153 ( .A1(in[200]), .A2(in[192]), .ZN(n810) );
  AND2_X1 U153bar ( .A1(inbar[200]), .A2(inbar[192]), .ZN(n810bar) );
  OR2_X1 U154 ( .A1(n808), .A2(n807), .ZN(n816) );
  AND2_X1 U154bar ( .A1(n808bar), .A2(n807bar), .ZN(n816bar) );
  OR2_X1 U155 ( .A1(n806), .A2(n805), .ZN(n807) );
  AND2_X1 U155bar ( .A1(n806bar), .A2(n805bar), .ZN(n807bar) );
  OR2_X1 U156 ( .A1(in[225]), .A2(in[207]), .ZN(n805) );
  AND2_X1 U156bar ( .A1(inbar[225]), .A2(inbar[207]), .ZN(n805bar) );
  OR2_X1 U157 ( .A1(in[98]), .A2(in[226]), .ZN(n806) );
  AND2_X1 U157bar ( .A1(inbar[98]), .A2(inbar[226]), .ZN(n806bar) );
  OR2_X1 U158 ( .A1(n804), .A2(n803), .ZN(n808) );
  AND2_X1 U158bar ( .A1(n804bar), .A2(n803bar), .ZN(n808bar) );
  OR2_X1 U159 ( .A1(in_20), .A2(in_16), .ZN(n803) );
  AND2_X1 U159bar ( .A1(in_20bar), .A2(in_16bar), .ZN(n803bar) );
  OR2_X1 U160 ( .A1(in_55), .A2(in_45), .ZN(n804) );
  AND2_X1 U160bar ( .A1(in_55bar), .A2(in_45bar), .ZN(n804bar) );
  OR2_X1 U161 ( .A1(n802), .A2(n801), .ZN(n824) );
  AND2_X1 U161bar ( .A1(n802bar), .A2(n801bar), .ZN(n824bar) );
  OR2_X1 U162 ( .A1(in[162]), .A2(in[149]), .ZN(n801) );
  AND2_X1 U162bar ( .A1(inbar[162]), .A2(inbar[149]), .ZN(n801bar) );
  OR2_X1 U163 ( .A1(in[163]), .A2(n800), .ZN(n802) );
  AND2_X1 U163bar ( .A1(inbar[163]), .A2(n800bar), .ZN(n802bar) );
  OR2_X1 U164 ( .A1(in[191]), .A2(in[189]), .ZN(n800) );
  AND2_X1 U164bar ( .A1(inbar[191]), .A2(inbar[189]), .ZN(n800bar) );
  OR2_X1 U165 ( .A1(n799), .A2(n798), .ZN(n826) );
  AND2_X1 U165bar ( .A1(n799bar), .A2(n798bar), .ZN(n826bar) );
  OR2_X1 U166 ( .A1(n797), .A2(n796), .ZN(n798) );
  AND2_X1 U166bar ( .A1(n797bar), .A2(n796bar), .ZN(n798bar) );
  OR2_X1 U167 ( .A1(in[212]), .A2(in[193]), .ZN(n796) );
  AND2_X1 U167bar ( .A1(inbar[212]), .A2(inbar[193]), .ZN(n796bar) );
  OR2_X1 U168 ( .A1(in[238]), .A2(n795), .ZN(n797) );
  AND2_X1 U168bar ( .A1(inbar[238]), .A2(n795bar), .ZN(n797bar) );
  OR2_X1 U169 ( .A1(in[88]), .A2(in[247]), .ZN(n795) );
  AND2_X1 U169bar ( .A1(inbar[88]), .A2(inbar[247]), .ZN(n795bar) );
  OR2_X1 U170 ( .A1(n794), .A2(n793), .ZN(n799) );
  AND2_X1 U170bar ( .A1(n794bar), .A2(n793bar), .ZN(n799bar) );
  OR2_X1 U171 ( .A1(in[94]), .A2(in[92]), .ZN(n793) );
  AND2_X1 U171bar ( .A1(inbar[94]), .A2(inbar[92]), .ZN(n793bar) );
  OR2_X1 U172 ( .A1(in_52), .A2(n792), .ZN(n794) );
  AND2_X1 U172bar ( .A1(in_52bar), .A2(n792bar), .ZN(n794bar) );
  OR2_X1 U173 ( .A1(in_70), .A2(in_67), .ZN(n792) );
  AND2_X1 U173bar ( .A1(in_70bar), .A2(in_67bar), .ZN(n792bar) );
  OR2_X1 U174 ( .A1(n791), .A2(n790), .ZN(out[2]) );
  AND2_X1 U174bar ( .A1(n791bar), .A2(n790bar), .ZN(outbar[2]) );
  OR2_X1 U175 ( .A1(n789), .A2(n788), .ZN(n790) );
  AND2_X1 U175bar ( .A1(n789bar), .A2(n788bar), .ZN(n790bar) );
  OR2_X1 U176 ( .A1(n787), .A2(n786), .ZN(n788) );
  AND2_X1 U176bar ( .A1(n787bar), .A2(n786bar), .ZN(n788bar) );
  OR2_X1 U177 ( .A1(n819), .A2(n785), .ZN(n786) );
  AND2_X1 U177bar ( .A1(n819bar), .A2(n785bar), .ZN(n786bar) );
  OR2_X1 U178 ( .A1(n784), .A2(n783), .ZN(n819) );
  AND2_X1 U178bar ( .A1(n784bar), .A2(n783bar), .ZN(n819bar) );
  OR2_X1 U179 ( .A1(n782), .A2(n781), .ZN(n783) );
  AND2_X1 U179bar ( .A1(n782bar), .A2(n781bar), .ZN(n783bar) );
  OR2_X1 U180 ( .A1(n780), .A2(n779), .ZN(n781) );
  AND2_X1 U180bar ( .A1(n780bar), .A2(n779bar), .ZN(n781bar) );
  OR2_X1 U181 ( .A1(n962), .A2(n778), .ZN(n779) );
  AND2_X1 U181bar ( .A1(n962bar), .A2(n778bar), .ZN(n779bar) );
  OR2_X1 U182 ( .A1(n777), .A2(n776), .ZN(n962) );
  AND2_X1 U182bar ( .A1(n777bar), .A2(n776bar), .ZN(n962bar) );
  OR2_X1 U183 ( .A1(n775), .A2(n774), .ZN(n776) );
  AND2_X1 U183bar ( .A1(n775bar), .A2(n774bar), .ZN(n776bar) );
  OR2_X1 U184 ( .A1(n773), .A2(n772), .ZN(n774) );
  AND2_X1 U184bar ( .A1(n773bar), .A2(n772bar), .ZN(n774bar) );
  OR2_X1 U185 ( .A1(in[131]), .A2(in[120]), .ZN(n772) );
  AND2_X1 U185bar ( .A1(inbar[131]), .A2(inbar[120]), .ZN(n772bar) );
  OR2_X1 U186 ( .A1(in[153]), .A2(in[147]), .ZN(n773) );
  AND2_X1 U186bar ( .A1(inbar[153]), .A2(inbar[147]), .ZN(n773bar) );
  OR2_X1 U187 ( .A1(n771), .A2(n770), .ZN(n775) );
  AND2_X1 U187bar ( .A1(n771bar), .A2(n770bar), .ZN(n775bar) );
  OR2_X1 U188 ( .A1(in[170]), .A2(in[156]), .ZN(n770) );
  AND2_X1 U188bar ( .A1(inbar[170]), .A2(inbar[156]), .ZN(n770bar) );
  OR2_X1 U189 ( .A1(in[223]), .A2(in[190]), .ZN(n771) );
  AND2_X1 U189bar ( .A1(inbar[223]), .A2(inbar[190]), .ZN(n771bar) );
  OR2_X1 U190 ( .A1(n769), .A2(n768), .ZN(n777) );
  AND2_X1 U190bar ( .A1(n769bar), .A2(n768bar), .ZN(n777bar) );
  OR2_X1 U191 ( .A1(n767), .A2(n766), .ZN(n768) );
  AND2_X1 U191bar ( .A1(n767bar), .A2(n766bar), .ZN(n768bar) );
  OR2_X1 U192 ( .A1(in[236]), .A2(in[230]), .ZN(n766) );
  AND2_X1 U192bar ( .A1(inbar[236]), .A2(inbar[230]), .ZN(n766bar) );
  OR2_X1 U193 ( .A1(in[85]), .A2(in[240]), .ZN(n767) );
  AND2_X1 U193bar ( .A1(inbar[85]), .A2(inbar[240]), .ZN(n767bar) );
  OR2_X1 U194 ( .A1(n765), .A2(n764), .ZN(n769) );
  AND2_X1 U194bar ( .A1(n765bar), .A2(n764bar), .ZN(n769bar) );
  OR2_X1 U195 ( .A1(in_12), .A2(in[90]), .ZN(n764) );
  AND2_X1 U195bar ( .A1(in_12bar), .A2(inbar[90]), .ZN(n764bar) );
  OR2_X1 U196 ( .A1(in_39), .A2(in_28), .ZN(n765) );
  AND2_X1 U196bar ( .A1(in_39bar), .A2(in_28bar), .ZN(n765bar) );
  OR2_X1 U197 ( .A1(in[109]), .A2(n763), .ZN(n780) );
  AND2_X1 U197bar ( .A1(inbar[109]), .A2(n763bar), .ZN(n780bar) );
  OR2_X1 U198 ( .A1(n762), .A2(n761), .ZN(n782) );
  AND2_X1 U198bar ( .A1(n762bar), .A2(n761bar), .ZN(n782bar) );
  OR2_X1 U199 ( .A1(in[138]), .A2(in[129]), .ZN(n761) );
  AND2_X1 U199bar ( .A1(inbar[138]), .A2(inbar[129]), .ZN(n761bar) );
  OR2_X1 U200 ( .A1(in[157]), .A2(n760), .ZN(n762) );
  AND2_X1 U200bar ( .A1(inbar[157]), .A2(n760bar), .ZN(n762bar) );
  OR2_X1 U201 ( .A1(in[182]), .A2(in[167]), .ZN(n760) );
  AND2_X1 U201bar ( .A1(inbar[182]), .A2(inbar[167]), .ZN(n760bar) );
  OR2_X1 U202 ( .A1(n759), .A2(n758), .ZN(n784) );
  AND2_X1 U202bar ( .A1(n759bar), .A2(n758bar), .ZN(n784bar) );
  OR2_X1 U203 ( .A1(n757), .A2(n756), .ZN(n758) );
  AND2_X1 U203bar ( .A1(n757bar), .A2(n756bar), .ZN(n758bar) );
  OR2_X1 U204 ( .A1(in[195]), .A2(in[184]), .ZN(n756) );
  AND2_X1 U204bar ( .A1(inbar[195]), .A2(inbar[184]), .ZN(n756bar) );
  OR2_X1 U205 ( .A1(in[196]), .A2(n755), .ZN(n757) );
  AND2_X1 U205bar ( .A1(inbar[196]), .A2(n755bar), .ZN(n757bar) );
  OR2_X1 U206 ( .A1(in[215]), .A2(in[209]), .ZN(n755) );
  AND2_X1 U206bar ( .A1(inbar[215]), .A2(inbar[209]), .ZN(n755bar) );
  OR2_X1 U207 ( .A1(n754), .A2(n753), .ZN(n759) );
  AND2_X1 U207bar ( .A1(n754bar), .A2(n753bar), .ZN(n759bar) );
  OR2_X1 U208 ( .A1(in[93]), .A2(in[233]), .ZN(n753) );
  AND2_X1 U208bar ( .A1(inbar[93]), .A2(inbar[233]), .ZN(n753bar) );
  OR2_X1 U209 ( .A1(in_1), .A2(n752), .ZN(n754) );
  AND2_X1 U209bar ( .A1(in_1bar), .A2(n752bar), .ZN(n754bar) );
  OR2_X1 U210 ( .A1(in_69), .A2(in_66), .ZN(n752) );
  AND2_X1 U210bar ( .A1(in_69bar), .A2(in_66bar), .ZN(n752bar) );
  OR2_X1 U211 ( .A1(n966), .A2(n751), .ZN(n787) );
  AND2_X1 U211bar ( .A1(n966bar), .A2(n751bar), .ZN(n787bar) );
  OR2_X1 U212 ( .A1(in[134]), .A2(n750), .ZN(n751) );
  AND2_X1 U212bar ( .A1(inbar[134]), .A2(n750bar), .ZN(n751bar) );
  OR2_X1 U213 ( .A1(n749), .A2(n748), .ZN(n966) );
  AND2_X1 U213bar ( .A1(n749bar), .A2(n748bar), .ZN(n966bar) );
  OR2_X1 U214 ( .A1(n747), .A2(n746), .ZN(n748) );
  AND2_X1 U214bar ( .A1(n747bar), .A2(n746bar), .ZN(n748bar) );
  OR2_X1 U215 ( .A1(n745), .A2(n744), .ZN(n746) );
  AND2_X1 U215bar ( .A1(n745bar), .A2(n744bar), .ZN(n746bar) );
  OR2_X1 U216 ( .A1(in[136]), .A2(in[121]), .ZN(n744) );
  AND2_X1 U216bar ( .A1(inbar[136]), .A2(inbar[121]), .ZN(n744bar) );
  OR2_X1 U217 ( .A1(in[186]), .A2(in[174]), .ZN(n745) );
  AND2_X1 U217bar ( .A1(inbar[186]), .A2(inbar[174]), .ZN(n745bar) );
  OR2_X1 U218 ( .A1(n743), .A2(n742), .ZN(n747) );
  AND2_X1 U218bar ( .A1(n743bar), .A2(n742bar), .ZN(n747bar) );
  OR2_X1 U219 ( .A1(in[198]), .A2(in[197]), .ZN(n742) );
  AND2_X1 U219bar ( .A1(inbar[198]), .A2(inbar[197]), .ZN(n742bar) );
  OR2_X1 U220 ( .A1(in[214]), .A2(in[199]), .ZN(n743) );
  AND2_X1 U220bar ( .A1(inbar[214]), .A2(inbar[199]), .ZN(n743bar) );
  OR2_X1 U221 ( .A1(n741), .A2(n740), .ZN(n749) );
  AND2_X1 U221bar ( .A1(n741bar), .A2(n740bar), .ZN(n749bar) );
  OR2_X1 U222 ( .A1(n739), .A2(n738), .ZN(n740) );
  AND2_X1 U222bar ( .A1(n739bar), .A2(n738bar), .ZN(n740bar) );
  OR2_X1 U223 ( .A1(in[231]), .A2(in[220]), .ZN(n738) );
  AND2_X1 U223bar ( .A1(inbar[231]), .A2(inbar[220]), .ZN(n738bar) );
  OR2_X1 U224 ( .A1(in_25), .A2(in[245]), .ZN(n739) );
  AND2_X1 U224bar ( .A1(in_25bar), .A2(inbar[245]), .ZN(n739bar) );
  OR2_X1 U225 ( .A1(n737), .A2(n736), .ZN(n741) );
  AND2_X1 U225bar ( .A1(n737bar), .A2(n736bar), .ZN(n741bar) );
  OR2_X1 U226 ( .A1(in_53), .A2(in_29), .ZN(n736) );
  AND2_X1 U226bar ( .A1(in_53bar), .A2(in_29bar), .ZN(n736bar) );
  OR2_X1 U227 ( .A1(in_79), .A2(in_74), .ZN(n737) );
  AND2_X1 U227bar ( .A1(in_79bar), .A2(in_74bar), .ZN(n737bar) );
  OR2_X1 U228 ( .A1(n735), .A2(n734), .ZN(n789) );
  AND2_X1 U228bar ( .A1(n735bar), .A2(n734bar), .ZN(n789bar) );
  OR2_X1 U229 ( .A1(in[152]), .A2(in[140]), .ZN(n734) );
  AND2_X1 U229bar ( .A1(inbar[152]), .A2(inbar[140]), .ZN(n734bar) );
  OR2_X1 U230 ( .A1(in[155]), .A2(n733), .ZN(n735) );
  AND2_X1 U230bar ( .A1(inbar[155]), .A2(n733bar), .ZN(n735bar) );
  OR2_X1 U231 ( .A1(in[166]), .A2(in[165]), .ZN(n733) );
  AND2_X1 U231bar ( .A1(inbar[166]), .A2(inbar[165]), .ZN(n733bar) );
  OR2_X1 U232 ( .A1(n732), .A2(n731), .ZN(n791) );
  AND2_X1 U232bar ( .A1(n732bar), .A2(n731bar), .ZN(n791bar) );
  OR2_X1 U233 ( .A1(n730), .A2(n729), .ZN(n731) );
  AND2_X1 U233bar ( .A1(n730bar), .A2(n729bar), .ZN(n731bar) );
  OR2_X1 U234 ( .A1(in[202]), .A2(in[185]), .ZN(n729) );
  AND2_X1 U234bar ( .A1(inbar[202]), .A2(inbar[185]), .ZN(n729bar) );
  OR2_X1 U235 ( .A1(in[211]), .A2(n728), .ZN(n730) );
  AND2_X1 U235bar ( .A1(inbar[211]), .A2(n728bar), .ZN(n730bar) );
  OR2_X1 U236 ( .A1(in[255]), .A2(in[253]), .ZN(n728) );
  AND2_X1 U236bar ( .A1(inbar[255]), .A2(inbar[253]), .ZN(n728bar) );
  OR2_X1 U237 ( .A1(n727), .A2(n726), .ZN(n732) );
  AND2_X1 U237bar ( .A1(n727bar), .A2(n726bar), .ZN(n732bar) );
  OR2_X1 U238 ( .A1(in_35), .A2(in_15), .ZN(n726) );
  AND2_X1 U238bar ( .A1(in_35bar), .A2(in_15bar), .ZN(n726bar) );
  OR2_X1 U239 ( .A1(in_36), .A2(n725), .ZN(n727) );
  AND2_X1 U239bar ( .A1(in_36bar), .A2(n725bar), .ZN(n727bar) );
  OR2_X1 U240 ( .A1(in_48), .A2(in_40), .ZN(n725) );
  AND2_X1 U240bar ( .A1(in_48bar), .A2(in_40bar), .ZN(n725bar) );
  OR2_X1 U241 ( .A1(n724), .A2(n723), .ZN(out[1]) );
  AND2_X1 U241bar ( .A1(n724bar), .A2(n723bar), .ZN(outbar[1]) );
  OR2_X1 U242 ( .A1(n722), .A2(n721), .ZN(n723) );
  AND2_X1 U242bar ( .A1(n722bar), .A2(n721bar), .ZN(n723bar) );
  OR2_X1 U243 ( .A1(n720), .A2(n719), .ZN(n721) );
  AND2_X1 U243bar ( .A1(n720bar), .A2(n719bar), .ZN(n721bar) );
  OR2_X1 U244 ( .A1(n921), .A2(n887), .ZN(n719) );
  AND2_X1 U244bar ( .A1(n921bar), .A2(n887bar), .ZN(n719bar) );
  OR2_X1 U245 ( .A1(n718), .A2(n717), .ZN(n887) );
  AND2_X1 U245bar ( .A1(n718bar), .A2(n717bar), .ZN(n887bar) );
  OR2_X1 U246 ( .A1(n716), .A2(n715), .ZN(n717) );
  AND2_X1 U246bar ( .A1(n716bar), .A2(n715bar), .ZN(n717bar) );
  OR2_X1 U247 ( .A1(n714), .A2(n713), .ZN(n715) );
  AND2_X1 U247bar ( .A1(n714bar), .A2(n713bar), .ZN(n715bar) );
  OR2_X1 U248 ( .A1(in[116]), .A2(in[110]), .ZN(n713) );
  AND2_X1 U248bar ( .A1(inbar[116]), .A2(inbar[110]), .ZN(n713bar) );
  OR2_X1 U249 ( .A1(in[133]), .A2(in[130]), .ZN(n714) );
  AND2_X1 U249bar ( .A1(inbar[133]), .A2(inbar[130]), .ZN(n714bar) );
  OR2_X1 U250 ( .A1(n712), .A2(n711), .ZN(n716) );
  AND2_X1 U250bar ( .A1(n712bar), .A2(n711bar), .ZN(n716bar) );
  OR2_X1 U251 ( .A1(in[203]), .A2(in[135]), .ZN(n711) );
  AND2_X1 U251bar ( .A1(inbar[203]), .A2(inbar[135]), .ZN(n711bar) );
  OR2_X1 U252 ( .A1(in[232]), .A2(in[223]), .ZN(n712) );
  AND2_X1 U252bar ( .A1(inbar[232]), .A2(inbar[223]), .ZN(n712bar) );
  OR2_X1 U253 ( .A1(n710), .A2(n709), .ZN(n718) );
  AND2_X1 U253bar ( .A1(n710bar), .A2(n709bar), .ZN(n718bar) );
  OR2_X1 U254 ( .A1(n708), .A2(n707), .ZN(n709) );
  AND2_X1 U254bar ( .A1(n708bar), .A2(n707bar), .ZN(n709bar) );
  OR2_X1 U255 ( .A1(in[255]), .A2(in[233]), .ZN(n707) );
  AND2_X1 U255bar ( .A1(inbar[255]), .A2(inbar[233]), .ZN(n707bar) );
  OR2_X1 U256 ( .A1(in_53), .A2(in_34), .ZN(n708) );
  AND2_X1 U256bar ( .A1(in_53bar), .A2(in_34bar), .ZN(n708bar) );
  OR2_X1 U257 ( .A1(n706), .A2(n705), .ZN(n710) );
  AND2_X1 U257bar ( .A1(n706bar), .A2(n705bar), .ZN(n710bar) );
  OR2_X1 U258 ( .A1(in_57), .A2(in_55), .ZN(n705) );
  AND2_X1 U258bar ( .A1(in_57bar), .A2(in_55bar), .ZN(n705bar) );
  OR2_X1 U259 ( .A1(in_68), .A2(in_67), .ZN(n706) );
  AND2_X1 U259bar ( .A1(in_68bar), .A2(in_67bar), .ZN(n706bar) );
  OR2_X1 U260 ( .A1(n704), .A2(n703), .ZN(n921) );
  AND2_X1 U260bar ( .A1(n704bar), .A2(n703bar), .ZN(n921bar) );
  OR2_X1 U261 ( .A1(n702), .A2(n701), .ZN(n703) );
  AND2_X1 U261bar ( .A1(n702bar), .A2(n701bar), .ZN(n703bar) );
  OR2_X1 U262 ( .A1(n700), .A2(n699), .ZN(n701) );
  AND2_X1 U262bar ( .A1(n700bar), .A2(n699bar), .ZN(n701bar) );
  OR2_X1 U263 ( .A1(n944), .A2(n872), .ZN(n699) );
  AND2_X1 U263bar ( .A1(n944bar), .A2(n872bar), .ZN(n699bar) );
  OR2_X1 U264 ( .A1(n698), .A2(n697), .ZN(n872) );
  AND2_X1 U264bar ( .A1(n698bar), .A2(n697bar), .ZN(n872bar) );
  OR2_X1 U265 ( .A1(n696), .A2(n695), .ZN(n697) );
  AND2_X1 U265bar ( .A1(n696bar), .A2(n695bar), .ZN(n697bar) );
  OR2_X1 U266 ( .A1(n694), .A2(n693), .ZN(n695) );
  AND2_X1 U266bar ( .A1(n694bar), .A2(n693bar), .ZN(n695bar) );
  OR2_X1 U267 ( .A1(in[121]), .A2(in[102]), .ZN(n693) );
  AND2_X1 U267bar ( .A1(inbar[121]), .A2(inbar[102]), .ZN(n693bar) );
  OR2_X1 U268 ( .A1(in[162]), .A2(in[161]), .ZN(n694) );
  AND2_X1 U268bar ( .A1(inbar[162]), .A2(inbar[161]), .ZN(n694bar) );
  OR2_X1 U269 ( .A1(n692), .A2(n691), .ZN(n696) );
  AND2_X1 U269bar ( .A1(n692bar), .A2(n691bar), .ZN(n696bar) );
  OR2_X1 U270 ( .A1(in[192]), .A2(in[178]), .ZN(n691) );
  AND2_X1 U270bar ( .A1(inbar[192]), .A2(inbar[178]), .ZN(n691bar) );
  OR2_X1 U271 ( .A1(in[244]), .A2(in[209]), .ZN(n692) );
  AND2_X1 U271bar ( .A1(inbar[244]), .A2(inbar[209]), .ZN(n692bar) );
  OR2_X1 U272 ( .A1(n690), .A2(n689), .ZN(n698) );
  AND2_X1 U272bar ( .A1(n690bar), .A2(n689bar), .ZN(n698bar) );
  OR2_X1 U273 ( .A1(n688), .A2(n687), .ZN(n689) );
  AND2_X1 U273bar ( .A1(n688bar), .A2(n687bar), .ZN(n689bar) );
  OR2_X1 U274 ( .A1(in[90]), .A2(in[254]), .ZN(n687) );
  AND2_X1 U274bar ( .A1(inbar[90]), .A2(inbar[254]), .ZN(n687bar) );
  OR2_X1 U275 ( .A1(in_36), .A2(in_32), .ZN(n688) );
  AND2_X1 U275bar ( .A1(in_36bar), .A2(in_32bar), .ZN(n688bar) );
  OR2_X1 U276 ( .A1(n686), .A2(n685), .ZN(n690) );
  AND2_X1 U276bar ( .A1(n686bar), .A2(n685bar), .ZN(n690bar) );
  OR2_X1 U277 ( .A1(in_62), .A2(in_37), .ZN(n685) );
  AND2_X1 U277bar ( .A1(in_62bar), .A2(in_37bar), .ZN(n685bar) );
  OR2_X1 U278 ( .A1(in_75), .A2(in_73), .ZN(n686) );
  AND2_X1 U278bar ( .A1(in_75bar), .A2(in_73bar), .ZN(n686bar) );
  OR2_X1 U279 ( .A1(n684), .A2(n683), .ZN(n944) );
  AND2_X1 U279bar ( .A1(n684bar), .A2(n683bar), .ZN(n944bar) );
  OR2_X1 U280 ( .A1(n682), .A2(n681), .ZN(n683) );
  AND2_X1 U280bar ( .A1(n682bar), .A2(n681bar), .ZN(n683bar) );
  OR2_X1 U281 ( .A1(n680), .A2(n679), .ZN(n681) );
  AND2_X1 U281bar ( .A1(n680bar), .A2(n679bar), .ZN(n681bar) );
  OR2_X1 U282 ( .A1(in[171]), .A2(in[153]), .ZN(n679) );
  AND2_X1 U282bar ( .A1(inbar[171]), .A2(inbar[153]), .ZN(n679bar) );
  OR2_X1 U283 ( .A1(in[187]), .A2(in[176]), .ZN(n680) );
  AND2_X1 U283bar ( .A1(inbar[187]), .A2(inbar[176]), .ZN(n680bar) );
  OR2_X1 U284 ( .A1(n678), .A2(n677), .ZN(n682) );
  AND2_X1 U284bar ( .A1(n678bar), .A2(n677bar), .ZN(n682bar) );
  OR2_X1 U285 ( .A1(in[245]), .A2(in[211]), .ZN(n677) );
  AND2_X1 U285bar ( .A1(inbar[245]), .A2(inbar[211]), .ZN(n677bar) );
  OR2_X1 U286 ( .A1(in[97]), .A2(in[88]), .ZN(n678) );
  AND2_X1 U286bar ( .A1(inbar[97]), .A2(inbar[88]), .ZN(n678bar) );
  OR2_X1 U287 ( .A1(n676), .A2(n675), .ZN(n684) );
  AND2_X1 U287bar ( .A1(n676bar), .A2(n675bar), .ZN(n684bar) );
  OR2_X1 U288 ( .A1(n674), .A2(n673), .ZN(n675) );
  AND2_X1 U288bar ( .A1(n674bar), .A2(n673bar), .ZN(n675bar) );
  OR2_X1 U289 ( .A1(in_10), .A2(in_0), .ZN(n673) );
  AND2_X1 U289bar ( .A1(in_10bar), .A2(in_0bar), .ZN(n673bar) );
  OR2_X1 U290 ( .A1(in_59), .A2(in_5), .ZN(n674) );
  AND2_X1 U290bar ( .A1(in_59bar), .A2(in_5bar), .ZN(n674bar) );
  OR2_X1 U291 ( .A1(n672), .A2(n671), .ZN(n676) );
  AND2_X1 U291bar ( .A1(n672bar), .A2(n671bar), .ZN(n676bar) );
  OR2_X1 U292 ( .A1(in_60), .A2(in_6), .ZN(n671) );
  AND2_X1 U292bar ( .A1(in_60bar), .A2(in_6bar), .ZN(n671bar) );
  OR2_X1 U293 ( .A1(in_77), .A2(in_69), .ZN(n672) );
  AND2_X1 U293bar ( .A1(in_77bar), .A2(in_69bar), .ZN(n672bar) );
  OR2_X1 U294 ( .A1(in[113]), .A2(n864), .ZN(n700) );
  AND2_X1 U294bar ( .A1(inbar[113]), .A2(n864bar), .ZN(n700bar) );
  OR2_X1 U295 ( .A1(n670), .A2(n669), .ZN(n864) );
  AND2_X1 U295bar ( .A1(n670bar), .A2(n669bar), .ZN(n864bar) );
  OR2_X1 U296 ( .A1(n668), .A2(n667), .ZN(n669) );
  AND2_X1 U296bar ( .A1(n668bar), .A2(n667bar), .ZN(n669bar) );
  OR2_X1 U297 ( .A1(n666), .A2(n665), .ZN(n667) );
  AND2_X1 U297bar ( .A1(n666bar), .A2(n665bar), .ZN(n667bar) );
  OR2_X1 U298 ( .A1(in[125]), .A2(in[107]), .ZN(n665) );
  AND2_X1 U298bar ( .A1(inbar[125]), .A2(inbar[107]), .ZN(n665bar) );
  OR2_X1 U299 ( .A1(in[138]), .A2(in[126]), .ZN(n666) );
  AND2_X1 U299bar ( .A1(inbar[138]), .A2(inbar[126]), .ZN(n666bar) );
  OR2_X1 U300 ( .A1(n664), .A2(n663), .ZN(n668) );
  AND2_X1 U300bar ( .A1(n664bar), .A2(n663bar), .ZN(n668bar) );
  OR2_X1 U301 ( .A1(in[189]), .A2(in[143]), .ZN(n663) );
  AND2_X1 U301bar ( .A1(inbar[189]), .A2(inbar[143]), .ZN(n663bar) );
  OR2_X1 U302 ( .A1(in[99]), .A2(in[214]), .ZN(n664) );
  AND2_X1 U302bar ( .A1(inbar[99]), .A2(inbar[214]), .ZN(n664bar) );
  OR2_X1 U303 ( .A1(n662), .A2(n661), .ZN(n670) );
  AND2_X1 U303bar ( .A1(n662bar), .A2(n661bar), .ZN(n670bar) );
  OR2_X1 U304 ( .A1(n660), .A2(n659), .ZN(n661) );
  AND2_X1 U304bar ( .A1(n660bar), .A2(n659bar), .ZN(n661bar) );
  OR2_X1 U305 ( .A1(in_15), .A2(in_12), .ZN(n659) );
  AND2_X1 U305bar ( .A1(in_15bar), .A2(in_12bar), .ZN(n659bar) );
  OR2_X1 U306 ( .A1(in_20), .A2(in_2), .ZN(n660) );
  AND2_X1 U306bar ( .A1(in_20bar), .A2(in_2bar), .ZN(n660bar) );
  OR2_X1 U307 ( .A1(n658), .A2(n657), .ZN(n662) );
  AND2_X1 U307bar ( .A1(n658bar), .A2(n657bar), .ZN(n662bar) );
  OR2_X1 U308 ( .A1(in_30), .A2(in_3), .ZN(n657) );
  AND2_X1 U308bar ( .A1(in_30bar), .A2(in_3bar), .ZN(n657bar) );
  OR2_X1 U309 ( .A1(in_4), .A2(in_38), .ZN(n658) );
  AND2_X1 U309bar ( .A1(in_4bar), .A2(in_38bar), .ZN(n658bar) );
  OR2_X1 U310 ( .A1(n656), .A2(n655), .ZN(n702) );
  AND2_X1 U310bar ( .A1(n656bar), .A2(n655bar), .ZN(n702bar) );
  OR2_X1 U311 ( .A1(in[148]), .A2(in[137]), .ZN(n655) );
  AND2_X1 U311bar ( .A1(inbar[148]), .A2(inbar[137]), .ZN(n655bar) );
  OR2_X1 U312 ( .A1(in[149]), .A2(n654), .ZN(n656) );
  AND2_X1 U312bar ( .A1(inbar[149]), .A2(n654bar), .ZN(n656bar) );
  OR2_X1 U313 ( .A1(in[195]), .A2(in[190]), .ZN(n654) );
  AND2_X1 U313bar ( .A1(inbar[195]), .A2(inbar[190]), .ZN(n654bar) );
  OR2_X1 U314 ( .A1(n653), .A2(n652), .ZN(n704) );
  AND2_X1 U314bar ( .A1(n653bar), .A2(n652bar), .ZN(n704bar) );
  OR2_X1 U315 ( .A1(n651), .A2(n650), .ZN(n652) );
  AND2_X1 U315bar ( .A1(n651bar), .A2(n650bar), .ZN(n652bar) );
  OR2_X1 U316 ( .A1(in[98]), .A2(in[197]), .ZN(n650) );
  AND2_X1 U316bar ( .A1(inbar[98]), .A2(inbar[197]), .ZN(n650bar) );
  OR2_X1 U317 ( .A1(in_11), .A2(n649), .ZN(n651) );
  AND2_X1 U317bar ( .A1(in_11bar), .A2(n649bar), .ZN(n651bar) );
  OR2_X1 U318 ( .A1(in_26), .A2(in_14), .ZN(n649) );
  AND2_X1 U318bar ( .A1(in_26bar), .A2(in_14bar), .ZN(n649bar) );
  OR2_X1 U319 ( .A1(n648), .A2(n647), .ZN(n653) );
  AND2_X1 U319bar ( .A1(n648bar), .A2(n647bar), .ZN(n653bar) );
  OR2_X1 U320 ( .A1(in_35), .A2(in_27), .ZN(n647) );
  AND2_X1 U320bar ( .A1(in_35bar), .A2(in_27bar), .ZN(n647bar) );
  OR2_X1 U321 ( .A1(in_50), .A2(n646), .ZN(n648) );
  AND2_X1 U321bar ( .A1(in_50bar), .A2(n646bar), .ZN(n648bar) );
  OR2_X1 U322 ( .A1(in_78), .A2(in_61), .ZN(n646) );
  AND2_X1 U322bar ( .A1(in_78bar), .A2(in_61bar), .ZN(n646bar) );
  OR2_X1 U323 ( .A1(n942), .A2(n645), .ZN(n720) );
  AND2_X1 U323bar ( .A1(n942bar), .A2(n645bar), .ZN(n720bar) );
  OR2_X1 U324 ( .A1(in[106]), .A2(n863), .ZN(n645) );
  AND2_X1 U324bar ( .A1(inbar[106]), .A2(n863bar), .ZN(n645bar) );
  OR2_X1 U325 ( .A1(n644), .A2(n643), .ZN(n863) );
  AND2_X1 U325bar ( .A1(n644bar), .A2(n643bar), .ZN(n863bar) );
  OR2_X1 U326 ( .A1(n642), .A2(n641), .ZN(n643) );
  AND2_X1 U326bar ( .A1(n642bar), .A2(n641bar), .ZN(n643bar) );
  OR2_X1 U327 ( .A1(n640), .A2(n639), .ZN(n641) );
  AND2_X1 U327bar ( .A1(n640bar), .A2(n639bar), .ZN(n641bar) );
  OR2_X1 U328 ( .A1(in[127]), .A2(in[122]), .ZN(n639) );
  AND2_X1 U328bar ( .A1(inbar[127]), .A2(inbar[122]), .ZN(n639bar) );
  OR2_X1 U329 ( .A1(in[156]), .A2(in[132]), .ZN(n640) );
  AND2_X1 U329bar ( .A1(inbar[156]), .A2(inbar[132]), .ZN(n640bar) );
  OR2_X1 U330 ( .A1(n638), .A2(n637), .ZN(n642) );
  AND2_X1 U330bar ( .A1(n638bar), .A2(n637bar), .ZN(n642bar) );
  OR2_X1 U331 ( .A1(in[159]), .A2(in[157]), .ZN(n637) );
  AND2_X1 U331bar ( .A1(inbar[159]), .A2(inbar[157]), .ZN(n637bar) );
  OR2_X1 U332 ( .A1(in[185]), .A2(in[169]), .ZN(n638) );
  AND2_X1 U332bar ( .A1(inbar[185]), .A2(inbar[169]), .ZN(n638bar) );
  OR2_X1 U333 ( .A1(n636), .A2(n635), .ZN(n644) );
  AND2_X1 U333bar ( .A1(n636bar), .A2(n635bar), .ZN(n644bar) );
  OR2_X1 U334 ( .A1(n634), .A2(n633), .ZN(n635) );
  AND2_X1 U334bar ( .A1(n634bar), .A2(n633bar), .ZN(n635bar) );
  OR2_X1 U335 ( .A1(in[239]), .A2(in[218]), .ZN(n633) );
  AND2_X1 U335bar ( .A1(inbar[239]), .A2(inbar[218]), .ZN(n633bar) );
  OR2_X1 U336 ( .A1(in_13), .A2(in[87]), .ZN(n634) );
  AND2_X1 U336bar ( .A1(in_13bar), .A2(inbar[87]), .ZN(n634bar) );
  OR2_X1 U337 ( .A1(n632), .A2(n631), .ZN(n636) );
  AND2_X1 U337bar ( .A1(n632bar), .A2(n631bar), .ZN(n636bar) );
  OR2_X1 U338 ( .A1(in_72), .A2(in_70), .ZN(n631) );
  AND2_X1 U338bar ( .A1(in_72bar), .A2(in_70bar), .ZN(n631bar) );
  OR2_X1 U339 ( .A1(in_80), .A2(in_74), .ZN(n632) );
  AND2_X1 U339bar ( .A1(in_80bar), .A2(in_74bar), .ZN(n632bar) );
  OR2_X1 U340 ( .A1(n630), .A2(n629), .ZN(n942) );
  AND2_X1 U340bar ( .A1(n630bar), .A2(n629bar), .ZN(n942bar) );
  OR2_X1 U341 ( .A1(n628), .A2(n627), .ZN(n629) );
  AND2_X1 U341bar ( .A1(n628bar), .A2(n627bar), .ZN(n629bar) );
  OR2_X1 U342 ( .A1(n626), .A2(n625), .ZN(n627) );
  AND2_X1 U342bar ( .A1(n626bar), .A2(n625bar), .ZN(n627bar) );
  OR2_X1 U343 ( .A1(in[146]), .A2(in[100]), .ZN(n625) );
  AND2_X1 U343bar ( .A1(inbar[146]), .A2(inbar[100]), .ZN(n625bar) );
  OR2_X1 U344 ( .A1(in[168]), .A2(in[152]), .ZN(n626) );
  AND2_X1 U344bar ( .A1(inbar[168]), .A2(inbar[152]), .ZN(n626bar) );
  OR2_X1 U345 ( .A1(n624), .A2(n623), .ZN(n628) );
  AND2_X1 U345bar ( .A1(n624bar), .A2(n623bar), .ZN(n628bar) );
  OR2_X1 U346 ( .A1(in[199]), .A2(in[182]), .ZN(n623) );
  AND2_X1 U346bar ( .A1(inbar[199]), .A2(inbar[182]), .ZN(n623bar) );
  OR2_X1 U347 ( .A1(in[236]), .A2(in[204]), .ZN(n624) );
  AND2_X1 U347bar ( .A1(inbar[236]), .A2(inbar[204]), .ZN(n624bar) );
  OR2_X1 U348 ( .A1(n622), .A2(n621), .ZN(n630) );
  AND2_X1 U348bar ( .A1(n622bar), .A2(n621bar), .ZN(n630bar) );
  OR2_X1 U349 ( .A1(n620), .A2(n619), .ZN(n621) );
  AND2_X1 U349bar ( .A1(n620bar), .A2(n619bar), .ZN(n621bar) );
  OR2_X1 U350 ( .A1(in[89]), .A2(in[246]), .ZN(n619) );
  AND2_X1 U350bar ( .A1(inbar[89]), .A2(inbar[246]), .ZN(n619bar) );
  OR2_X1 U351 ( .A1(in[95]), .A2(in[92]), .ZN(n620) );
  AND2_X1 U351bar ( .A1(inbar[95]), .A2(inbar[92]), .ZN(n620bar) );
  OR2_X1 U352 ( .A1(n618), .A2(n617), .ZN(n622) );
  AND2_X1 U352bar ( .A1(n618bar), .A2(n617bar), .ZN(n622bar) );
  OR2_X1 U353 ( .A1(in_22), .A2(in_16), .ZN(n617) );
  AND2_X1 U353bar ( .A1(in_22bar), .A2(in_16bar), .ZN(n617bar) );
  OR2_X1 U354 ( .A1(in_51), .A2(in_49), .ZN(n618) );
  AND2_X1 U354bar ( .A1(in_51bar), .A2(in_49bar), .ZN(n618bar) );
  OR2_X1 U355 ( .A1(n616), .A2(n615), .ZN(n722) );
  AND2_X1 U355bar ( .A1(n616bar), .A2(n615bar), .ZN(n722bar) );
  OR2_X1 U356 ( .A1(in[158]), .A2(in[115]), .ZN(n615) );
  AND2_X1 U356bar ( .A1(inbar[158]), .A2(inbar[115]), .ZN(n615bar) );
  OR2_X1 U357 ( .A1(in[163]), .A2(n614), .ZN(n616) );
  AND2_X1 U357bar ( .A1(inbar[163]), .A2(n614bar), .ZN(n616bar) );
  OR2_X1 U358 ( .A1(in[206]), .A2(in[165]), .ZN(n614) );
  AND2_X1 U358bar ( .A1(inbar[206]), .A2(inbar[165]), .ZN(n614bar) );
  OR2_X1 U359 ( .A1(n613), .A2(n612), .ZN(n724) );
  AND2_X1 U359bar ( .A1(n613bar), .A2(n612bar), .ZN(n724bar) );
  OR2_X1 U360 ( .A1(n611), .A2(n610), .ZN(n612) );
  AND2_X1 U360bar ( .A1(n611bar), .A2(n610bar), .ZN(n612bar) );
  OR2_X1 U361 ( .A1(in[213]), .A2(in[207]), .ZN(n610) );
  AND2_X1 U361bar ( .A1(inbar[213]), .A2(inbar[207]), .ZN(n610bar) );
  OR2_X1 U362 ( .A1(in[215]), .A2(n609), .ZN(n611) );
  AND2_X1 U362bar ( .A1(inbar[215]), .A2(n609bar), .ZN(n611bar) );
  OR2_X1 U363 ( .A1(in[230]), .A2(in[220]), .ZN(n609) );
  AND2_X1 U363bar ( .A1(inbar[230]), .A2(inbar[220]), .ZN(n609bar) );
  OR2_X1 U364 ( .A1(n608), .A2(n607), .ZN(n613) );
  AND2_X1 U364bar ( .A1(n608bar), .A2(n607bar), .ZN(n613bar) );
  OR2_X1 U365 ( .A1(in[251]), .A2(in[234]), .ZN(n607) );
  AND2_X1 U365bar ( .A1(inbar[251]), .A2(inbar[234]), .ZN(n607bar) );
  OR2_X1 U366 ( .A1(in_17), .A2(n606), .ZN(n608) );
  AND2_X1 U366bar ( .A1(in_17bar), .A2(n606bar), .ZN(n608bar) );
  OR2_X1 U367 ( .A1(in_65), .A2(in_56), .ZN(n606) );
  AND2_X1 U367bar ( .A1(in_65bar), .A2(in_56bar), .ZN(n606bar) );
  OR2_X1 U368 ( .A1(n605), .A2(n604), .ZN(out[0]) );
  AND2_X1 U368bar ( .A1(n605bar), .A2(n604bar), .ZN(outbar[0]) );
  OR2_X1 U369 ( .A1(n603), .A2(n602), .ZN(n604) );
  AND2_X1 U369bar ( .A1(n603bar), .A2(n602bar), .ZN(n604bar) );
  OR2_X1 U370 ( .A1(n601), .A2(n600), .ZN(n602) );
  AND2_X1 U370bar ( .A1(n601bar), .A2(n600bar), .ZN(n602bar) );
  OR2_X1 U371 ( .A1(n820), .A2(n785), .ZN(n600) );
  AND2_X1 U371bar ( .A1(n820bar), .A2(n785bar), .ZN(n600bar) );
  OR2_X1 U372 ( .A1(n599), .A2(n598), .ZN(n785) );
  AND2_X1 U372bar ( .A1(n599bar), .A2(n598bar), .ZN(n785bar) );
  OR2_X1 U373 ( .A1(n597), .A2(n596), .ZN(n598) );
  AND2_X1 U373bar ( .A1(n597bar), .A2(n596bar), .ZN(n598bar) );
  OR2_X1 U374 ( .A1(n595), .A2(n594), .ZN(n596) );
  AND2_X1 U374bar ( .A1(n595bar), .A2(n594bar), .ZN(n596bar) );
  OR2_X1 U375 ( .A1(in[135]), .A2(in[104]), .ZN(n594) );
  AND2_X1 U375bar ( .A1(inbar[135]), .A2(inbar[104]), .ZN(n594bar) );
  OR2_X1 U376 ( .A1(in[188]), .A2(in[178]), .ZN(n595) );
  AND2_X1 U376bar ( .A1(inbar[188]), .A2(inbar[178]), .ZN(n595bar) );
  OR2_X1 U377 ( .A1(n593), .A2(n592), .ZN(n597) );
  AND2_X1 U377bar ( .A1(n593bar), .A2(n592bar), .ZN(n597bar) );
  OR2_X1 U378 ( .A1(in[217]), .A2(in[194]), .ZN(n592) );
  AND2_X1 U378bar ( .A1(inbar[217]), .A2(inbar[194]), .ZN(n592bar) );
  OR2_X1 U379 ( .A1(in[237]), .A2(in[218]), .ZN(n593) );
  AND2_X1 U379bar ( .A1(inbar[237]), .A2(inbar[218]), .ZN(n593bar) );
  OR2_X1 U380 ( .A1(n591), .A2(n590), .ZN(n599) );
  AND2_X1 U380bar ( .A1(n591bar), .A2(n590bar), .ZN(n599bar) );
  OR2_X1 U381 ( .A1(n589), .A2(n588), .ZN(n590) );
  AND2_X1 U381bar ( .A1(n589bar), .A2(n588bar), .ZN(n590bar) );
  OR2_X1 U382 ( .A1(in_2), .A2(in_10), .ZN(n588) );
  AND2_X1 U382bar ( .A1(in_2bar), .A2(in_10bar), .ZN(n588bar) );
  OR2_X1 U383 ( .A1(in_47), .A2(in_22), .ZN(n589) );
  AND2_X1 U383bar ( .A1(in_47bar), .A2(in_22bar), .ZN(n589bar) );
  OR2_X1 U384 ( .A1(n587), .A2(n586), .ZN(n591) );
  AND2_X1 U384bar ( .A1(n587bar), .A2(n586bar), .ZN(n591bar) );
  OR2_X1 U385 ( .A1(in_56), .A2(in_54), .ZN(n586) );
  AND2_X1 U385bar ( .A1(in_56bar), .A2(in_54bar), .ZN(n586bar) );
  OR2_X1 U386 ( .A1(in_63), .A2(in_61), .ZN(n587) );
  AND2_X1 U386bar ( .A1(in_63bar), .A2(in_61bar), .ZN(n587bar) );
  OR2_X1 U387 ( .A1(n585), .A2(n584), .ZN(n820) );
  AND2_X1 U387bar ( .A1(n585bar), .A2(n584bar), .ZN(n820bar) );
  OR2_X1 U388 ( .A1(n583), .A2(n582), .ZN(n584) );
  AND2_X1 U388bar ( .A1(n583bar), .A2(n582bar), .ZN(n584bar) );
  OR2_X1 U389 ( .A1(n581), .A2(n580), .ZN(n582) );
  AND2_X1 U389bar ( .A1(n581bar), .A2(n580bar), .ZN(n582bar) );
  OR2_X1 U390 ( .A1(in[158]), .A2(in[142]), .ZN(n580) );
  AND2_X1 U390bar ( .A1(inbar[158]), .A2(inbar[142]), .ZN(n580bar) );
  OR2_X1 U391 ( .A1(in[175]), .A2(in[164]), .ZN(n581) );
  AND2_X1 U391bar ( .A1(inbar[175]), .A2(inbar[164]), .ZN(n581bar) );
  OR2_X1 U392 ( .A1(n579), .A2(n578), .ZN(n583) );
  AND2_X1 U392bar ( .A1(n579bar), .A2(n578bar), .ZN(n583bar) );
  OR2_X1 U393 ( .A1(in[228]), .A2(in[204]), .ZN(n578) );
  AND2_X1 U393bar ( .A1(inbar[228]), .A2(inbar[204]), .ZN(n578bar) );
  OR2_X1 U394 ( .A1(in[91]), .A2(in[87]), .ZN(n579) );
  AND2_X1 U394bar ( .A1(inbar[91]), .A2(inbar[87]), .ZN(n579bar) );
  OR2_X1 U395 ( .A1(n577), .A2(n576), .ZN(n585) );
  AND2_X1 U395bar ( .A1(n577bar), .A2(n576bar), .ZN(n585bar) );
  OR2_X1 U396 ( .A1(n575), .A2(n574), .ZN(n576) );
  AND2_X1 U396bar ( .A1(n575bar), .A2(n574bar), .ZN(n576bar) );
  OR2_X1 U397 ( .A1(in_21), .A2(in_11), .ZN(n574) );
  AND2_X1 U397bar ( .A1(in_21bar), .A2(in_11bar), .ZN(n574bar) );
  OR2_X1 U398 ( .A1(in_5), .A2(in_3), .ZN(n575) );
  AND2_X1 U398bar ( .A1(in_5bar), .A2(in_3bar), .ZN(n575bar) );
  OR2_X1 U399 ( .A1(n573), .A2(n572), .ZN(n577) );
  AND2_X1 U399bar ( .A1(n573bar), .A2(n572bar), .ZN(n577bar) );
  OR2_X1 U400 ( .A1(in_68), .A2(in_64), .ZN(n572) );
  AND2_X1 U400bar ( .A1(in_68bar), .A2(in_64bar), .ZN(n572bar) );
  OR2_X1 U401 ( .A1(in_76), .A2(in_73), .ZN(n573) );
  AND2_X1 U401bar ( .A1(in_76bar), .A2(in_73bar), .ZN(n573bar) );
  OR2_X1 U402 ( .A1(n778), .A2(n571), .ZN(n601) );
  AND2_X1 U402bar ( .A1(n778bar), .A2(n571bar), .ZN(n601bar) );
  OR2_X1 U403 ( .A1(in[100]), .A2(n965), .ZN(n571) );
  AND2_X1 U403bar ( .A1(inbar[100]), .A2(n965bar), .ZN(n571bar) );
  OR2_X1 U404 ( .A1(n570), .A2(n569), .ZN(n965) );
  AND2_X1 U404bar ( .A1(n570bar), .A2(n569bar), .ZN(n965bar) );
  OR2_X1 U405 ( .A1(n568), .A2(n567), .ZN(n569) );
  AND2_X1 U405bar ( .A1(n568bar), .A2(n567bar), .ZN(n569bar) );
  OR2_X1 U406 ( .A1(n566), .A2(n565), .ZN(n567) );
  AND2_X1 U406bar ( .A1(n566bar), .A2(n565bar), .ZN(n567bar) );
  OR2_X1 U407 ( .A1(n817), .A2(n750), .ZN(n565) );
  AND2_X1 U407bar ( .A1(n817bar), .A2(n750bar), .ZN(n565bar) );
  OR2_X1 U408 ( .A1(n564), .A2(n563), .ZN(n750) );
  AND2_X1 U408bar ( .A1(n564bar), .A2(n563bar), .ZN(n750bar) );
  OR2_X1 U409 ( .A1(n562), .A2(n561), .ZN(n563) );
  AND2_X1 U409bar ( .A1(n562bar), .A2(n561bar), .ZN(n563bar) );
  OR2_X1 U410 ( .A1(n560), .A2(n559), .ZN(n561) );
  AND2_X1 U410bar ( .A1(n560bar), .A2(n559bar), .ZN(n561bar) );
  OR2_X1 U411 ( .A1(in[119]), .A2(in[103]), .ZN(n559) );
  AND2_X1 U411bar ( .A1(inbar[119]), .A2(inbar[103]), .ZN(n559bar) );
  OR2_X1 U412 ( .A1(in[137]), .A2(in[133]), .ZN(n560) );
  AND2_X1 U412bar ( .A1(inbar[137]), .A2(inbar[133]), .ZN(n560bar) );
  OR2_X1 U413 ( .A1(n558), .A2(n557), .ZN(n562) );
  AND2_X1 U413bar ( .A1(n558bar), .A2(n557bar), .ZN(n562bar) );
  OR2_X1 U414 ( .A1(in[176]), .A2(in[173]), .ZN(n557) );
  AND2_X1 U414bar ( .A1(inbar[176]), .A2(inbar[173]), .ZN(n557bar) );
  OR2_X1 U415 ( .A1(in[210]), .A2(in[181]), .ZN(n558) );
  AND2_X1 U415bar ( .A1(inbar[210]), .A2(inbar[181]), .ZN(n558bar) );
  OR2_X1 U416 ( .A1(n556), .A2(n555), .ZN(n564) );
  AND2_X1 U416bar ( .A1(n556bar), .A2(n555bar), .ZN(n564bar) );
  OR2_X1 U417 ( .A1(n554), .A2(n553), .ZN(n555) );
  AND2_X1 U417bar ( .A1(n554bar), .A2(n553bar), .ZN(n555bar) );
  OR2_X1 U418 ( .A1(in_13), .A2(in[234]), .ZN(n553) );
  AND2_X1 U418bar ( .A1(in_13bar), .A2(inbar[234]), .ZN(n553bar) );
  OR2_X1 U419 ( .A1(in_38), .A2(in_32), .ZN(n554) );
  AND2_X1 U419bar ( .A1(in_38bar), .A2(in_32bar), .ZN(n554bar) );
  OR2_X1 U420 ( .A1(n552), .A2(n551), .ZN(n556) );
  AND2_X1 U420bar ( .A1(n552bar), .A2(n551bar), .ZN(n556bar) );
  OR2_X1 U421 ( .A1(in_42), .A2(in_41), .ZN(n551) );
  AND2_X1 U421bar ( .A1(in_42bar), .A2(in_41bar), .ZN(n551bar) );
  OR2_X1 U422 ( .A1(in_7), .A2(in_49), .ZN(n552) );
  AND2_X1 U422bar ( .A1(in_7bar), .A2(in_49bar), .ZN(n552bar) );
  OR2_X1 U423 ( .A1(n550), .A2(n549), .ZN(n817) );
  AND2_X1 U423bar ( .A1(n550bar), .A2(n549bar), .ZN(n817bar) );
  OR2_X1 U424 ( .A1(n548), .A2(n547), .ZN(n549) );
  AND2_X1 U424bar ( .A1(n548bar), .A2(n547bar), .ZN(n549bar) );
  OR2_X1 U425 ( .A1(n546), .A2(n545), .ZN(n547) );
  AND2_X1 U425bar ( .A1(n546bar), .A2(n545bar), .ZN(n547bar) );
  OR2_X1 U426 ( .A1(in[159]), .A2(in[105]), .ZN(n545) );
  AND2_X1 U426bar ( .A1(inbar[159]), .A2(inbar[105]), .ZN(n545bar) );
  OR2_X1 U427 ( .A1(in[206]), .A2(in[183]), .ZN(n546) );
  AND2_X1 U427bar ( .A1(inbar[206]), .A2(inbar[183]), .ZN(n546bar) );
  OR2_X1 U428 ( .A1(n544), .A2(n543), .ZN(n548) );
  AND2_X1 U428bar ( .A1(n544bar), .A2(n543bar), .ZN(n548bar) );
  OR2_X1 U429 ( .A1(in[229]), .A2(in[219]), .ZN(n543) );
  AND2_X1 U429bar ( .A1(inbar[229]), .A2(inbar[219]), .ZN(n543bar) );
  OR2_X1 U430 ( .A1(in[235]), .A2(in[232]), .ZN(n544) );
  AND2_X1 U430bar ( .A1(inbar[235]), .A2(inbar[232]), .ZN(n544bar) );
  OR2_X1 U431 ( .A1(n542), .A2(n541), .ZN(n550) );
  AND2_X1 U431bar ( .A1(n542bar), .A2(n541bar), .ZN(n550bar) );
  OR2_X1 U432 ( .A1(n540), .A2(n539), .ZN(n541) );
  AND2_X1 U432bar ( .A1(n540bar), .A2(n539bar), .ZN(n541bar) );
  OR2_X1 U433 ( .A1(in[249]), .A2(in[242]), .ZN(n539) );
  AND2_X1 U433bar ( .A1(inbar[249]), .A2(inbar[242]), .ZN(n539bar) );
  OR2_X1 U434 ( .A1(in[89]), .A2(in[254]), .ZN(n540) );
  AND2_X1 U434bar ( .A1(inbar[89]), .A2(inbar[254]), .ZN(n540bar) );
  OR2_X1 U435 ( .A1(n538), .A2(n537), .ZN(n542) );
  AND2_X1 U435bar ( .A1(n538bar), .A2(n537bar), .ZN(n542bar) );
  OR2_X1 U436 ( .A1(in_14), .A2(in[99]), .ZN(n537) );
  AND2_X1 U436bar ( .A1(in_14bar), .A2(inbar[99]), .ZN(n537bar) );
  OR2_X1 U437 ( .A1(in_60), .A2(in_18), .ZN(n538) );
  AND2_X1 U437bar ( .A1(in_60bar), .A2(in_18bar), .ZN(n538bar) );
  OR2_X1 U438 ( .A1(in[113]), .A2(n763), .ZN(n566) );
  AND2_X1 U438bar ( .A1(inbar[113]), .A2(n763bar), .ZN(n566bar) );
  OR2_X1 U439 ( .A1(n536), .A2(n535), .ZN(n763) );
  AND2_X1 U439bar ( .A1(n536bar), .A2(n535bar), .ZN(n763bar) );
  OR2_X1 U440 ( .A1(n534), .A2(n533), .ZN(n535) );
  AND2_X1 U440bar ( .A1(n534bar), .A2(n533bar), .ZN(n535bar) );
  OR2_X1 U441 ( .A1(n532), .A2(n531), .ZN(n533) );
  AND2_X1 U441bar ( .A1(n532bar), .A2(n531bar), .ZN(n533bar) );
  OR2_X1 U442 ( .A1(in[115]), .A2(in[110]), .ZN(n531) );
  AND2_X1 U442bar ( .A1(inbar[115]), .A2(inbar[110]), .ZN(n531bar) );
  OR2_X1 U443 ( .A1(in[125]), .A2(in[117]), .ZN(n532) );
  AND2_X1 U443bar ( .A1(inbar[125]), .A2(inbar[117]), .ZN(n532bar) );
  OR2_X1 U444 ( .A1(n530), .A2(n529), .ZN(n534) );
  AND2_X1 U444bar ( .A1(n530bar), .A2(n529bar), .ZN(n534bar) );
  OR2_X1 U445 ( .A1(in[180]), .A2(in[128]), .ZN(n529) );
  AND2_X1 U445bar ( .A1(inbar[180]), .A2(inbar[128]), .ZN(n529bar) );
  OR2_X1 U446 ( .A1(in[205]), .A2(in[201]), .ZN(n530) );
  AND2_X1 U446bar ( .A1(inbar[205]), .A2(inbar[201]), .ZN(n530bar) );
  OR2_X1 U447 ( .A1(n528), .A2(n527), .ZN(n536) );
  AND2_X1 U447bar ( .A1(n528bar), .A2(n527bar), .ZN(n536bar) );
  OR2_X1 U448 ( .A1(n526), .A2(n525), .ZN(n527) );
  AND2_X1 U448bar ( .A1(n526bar), .A2(n525bar), .ZN(n527bar) );
  OR2_X1 U449 ( .A1(in[244]), .A2(in[239]), .ZN(n525) );
  AND2_X1 U449bar ( .A1(inbar[244]), .A2(inbar[239]), .ZN(n525bar) );
  OR2_X1 U450 ( .A1(in[95]), .A2(in[83]), .ZN(n526) );
  AND2_X1 U450bar ( .A1(inbar[95]), .A2(inbar[83]), .ZN(n526bar) );
  OR2_X1 U451 ( .A1(n524), .A2(n523), .ZN(n528) );
  AND2_X1 U451bar ( .A1(n524bar), .A2(n523bar), .ZN(n528bar) );
  OR2_X1 U452 ( .A1(in_24), .A2(in[97]), .ZN(n523) );
  AND2_X1 U452bar ( .A1(in_24bar), .A2(inbar[97]), .ZN(n523bar) );
  OR2_X1 U453 ( .A1(in_33), .A2(in_27), .ZN(n524) );
  AND2_X1 U453bar ( .A1(in_33bar), .A2(in_27bar), .ZN(n524bar) );
  OR2_X1 U454 ( .A1(n522), .A2(n521), .ZN(n568) );
  AND2_X1 U454bar ( .A1(n522bar), .A2(n521bar), .ZN(n568bar) );
  OR2_X1 U455 ( .A1(in[145]), .A2(in[126]), .ZN(n521) );
  AND2_X1 U455bar ( .A1(inbar[145]), .A2(inbar[126]), .ZN(n521bar) );
  OR2_X1 U456 ( .A1(in[169]), .A2(n520), .ZN(n522) );
  AND2_X1 U456bar ( .A1(inbar[169]), .A2(n520bar), .ZN(n522bar) );
  OR2_X1 U457 ( .A1(in[221]), .A2(in[172]), .ZN(n520) );
  AND2_X1 U457bar ( .A1(inbar[221]), .A2(inbar[172]), .ZN(n520bar) );
  OR2_X1 U458 ( .A1(n519), .A2(n518), .ZN(n570) );
  AND2_X1 U458bar ( .A1(n519bar), .A2(n518bar), .ZN(n570bar) );
  OR2_X1 U459 ( .A1(n517), .A2(n516), .ZN(n518) );
  AND2_X1 U459bar ( .A1(n517bar), .A2(n516bar), .ZN(n518bar) );
  OR2_X1 U460 ( .A1(in[241]), .A2(in[224]), .ZN(n516) );
  AND2_X1 U460bar ( .A1(inbar[241]), .A2(inbar[224]), .ZN(n516bar) );
  OR2_X1 U461 ( .A1(in[86]), .A2(n515), .ZN(n517) );
  AND2_X1 U461bar ( .A1(inbar[86]), .A2(n515bar), .ZN(n517bar) );
  OR2_X1 U462 ( .A1(in_43), .A2(in_34), .ZN(n515) );
  AND2_X1 U462bar ( .A1(in_43bar), .A2(in_34bar), .ZN(n515bar) );
  OR2_X1 U463 ( .A1(n514), .A2(n513), .ZN(n519) );
  AND2_X1 U463bar ( .A1(n514bar), .A2(n513bar), .ZN(n519bar) );
  OR2_X1 U464 ( .A1(in_65), .A2(in_51), .ZN(n513) );
  AND2_X1 U464bar ( .A1(in_65bar), .A2(in_51bar), .ZN(n513bar) );
  OR2_X1 U465 ( .A1(in_75), .A2(n512), .ZN(n514) );
  AND2_X1 U465bar ( .A1(in_75bar), .A2(n512bar), .ZN(n514bar) );
  OR2_X1 U466 ( .A1(in_81), .A2(in_77), .ZN(n512) );
  AND2_X1 U466bar ( .A1(in_81bar), .A2(in_77bar), .ZN(n512bar) );
  OR2_X1 U467 ( .A1(n511), .A2(n510), .ZN(n778) );
  AND2_X1 U467bar ( .A1(n511bar), .A2(n510bar), .ZN(n778bar) );
  OR2_X1 U468 ( .A1(n509), .A2(n508), .ZN(n510) );
  AND2_X1 U468bar ( .A1(n509bar), .A2(n508bar), .ZN(n510bar) );
  OR2_X1 U469 ( .A1(n507), .A2(n506), .ZN(n508) );
  AND2_X1 U469bar ( .A1(n507bar), .A2(n506bar), .ZN(n508bar) );
  OR2_X1 U470 ( .A1(in[107]), .A2(in[101]), .ZN(n506) );
  AND2_X1 U470bar ( .A1(inbar[107]), .A2(inbar[101]), .ZN(n506bar) );
  OR2_X1 U471 ( .A1(in[139]), .A2(in[132]), .ZN(n507) );
  AND2_X1 U471bar ( .A1(inbar[139]), .A2(inbar[132]), .ZN(n507bar) );
  OR2_X1 U472 ( .A1(n505), .A2(n504), .ZN(n509) );
  AND2_X1 U472bar ( .A1(n505bar), .A2(n504bar), .ZN(n509bar) );
  OR2_X1 U473 ( .A1(in[146]), .A2(in[141]), .ZN(n504) );
  AND2_X1 U473bar ( .A1(inbar[146]), .A2(inbar[141]), .ZN(n504bar) );
  OR2_X1 U474 ( .A1(in[203]), .A2(in[179]), .ZN(n505) );
  AND2_X1 U474bar ( .A1(inbar[203]), .A2(inbar[179]), .ZN(n505bar) );
  OR2_X1 U475 ( .A1(n503), .A2(n502), .ZN(n511) );
  AND2_X1 U475bar ( .A1(n503bar), .A2(n502bar), .ZN(n511bar) );
  OR2_X1 U476 ( .A1(n501), .A2(n500), .ZN(n502) );
  AND2_X1 U476bar ( .A1(n501bar), .A2(n500bar), .ZN(n502bar) );
  OR2_X1 U477 ( .A1(in[243]), .A2(in[222]), .ZN(n500) );
  AND2_X1 U477bar ( .A1(inbar[243]), .A2(inbar[222]), .ZN(n500bar) );
  OR2_X1 U478 ( .A1(in[251]), .A2(in[250]), .ZN(n501) );
  AND2_X1 U478bar ( .A1(inbar[251]), .A2(inbar[250]), .ZN(n501bar) );
  OR2_X1 U479 ( .A1(n499), .A2(n498), .ZN(n503) );
  AND2_X1 U479bar ( .A1(n499bar), .A2(n498bar), .ZN(n503bar) );
  OR2_X1 U480 ( .A1(in_37), .A2(in_19), .ZN(n498) );
  AND2_X1 U480bar ( .A1(in_37bar), .A2(in_19bar), .ZN(n498bar) );
  OR2_X1 U481 ( .A1(in_78), .A2(in_6), .ZN(n499) );
  AND2_X1 U481bar ( .A1(in_78bar), .A2(in_6bar), .ZN(n499bar) );
  OR2_X1 U482 ( .A1(n497), .A2(n496), .ZN(n603) );
  AND2_X1 U482bar ( .A1(n497bar), .A2(n496bar), .ZN(n603bar) );
  OR2_X1 U483 ( .A1(in[112]), .A2(in[102]), .ZN(n496) );
  AND2_X1 U483bar ( .A1(inbar[112]), .A2(inbar[102]), .ZN(n496bar) );
  OR2_X1 U484 ( .A1(in[123]), .A2(n495), .ZN(n497) );
  AND2_X1 U484bar ( .A1(inbar[123]), .A2(n495bar), .ZN(n497bar) );
  OR2_X1 U485 ( .A1(in[143]), .A2(in[130]), .ZN(n495) );
  AND2_X1 U485bar ( .A1(inbar[143]), .A2(inbar[130]), .ZN(n495bar) );
  OR2_X1 U486 ( .A1(n494), .A2(n493), .ZN(n605) );
  AND2_X1 U486bar ( .A1(n494bar), .A2(n493bar), .ZN(n605bar) );
  OR2_X1 U487 ( .A1(n492), .A2(n491), .ZN(n493) );
  AND2_X1 U487bar ( .A1(n492bar), .A2(n491bar), .ZN(n493bar) );
  OR2_X1 U488 ( .A1(in[216]), .A2(in[213]), .ZN(n491) );
  AND2_X1 U488bar ( .A1(inbar[216]), .A2(inbar[213]), .ZN(n491bar) );
  OR2_X1 U489 ( .A1(in[227]), .A2(n490), .ZN(n492) );
  AND2_X1 U489bar ( .A1(inbar[227]), .A2(n490bar), .ZN(n492bar) );
  OR2_X1 U490 ( .A1(in_0), .A2(in[248]), .ZN(n490) );
  AND2_X1 U490bar ( .A1(in_0bar), .A2(inbar[248]), .ZN(n490bar) );
  OR2_X1 U491 ( .A1(n489), .A2(n488), .ZN(n494) );
  AND2_X1 U491bar ( .A1(n489bar), .A2(n488bar), .ZN(n494bar) );
  OR2_X1 U492 ( .A1(in_46), .A2(in_44), .ZN(n488) );
  AND2_X1 U492bar ( .A1(in_46bar), .A2(in_44bar), .ZN(n488bar) );
  OR2_X1 U493 ( .A1(in_50), .A2(n487), .ZN(n489) );
  AND2_X1 U493bar ( .A1(in_50bar), .A2(n487bar), .ZN(n489bar) );
  OR2_X1 U494 ( .A1(in_9), .A2(in_80), .ZN(n487) );
  AND2_X1 U494bar ( .A1(in_9bar), .A2(in_80bar), .ZN(n487bar) );
endmodule

module sBox_11 ( in, inbar, out, outbar );

  input wire [7:0] in;
  input wire [7:0] inbar;
//input_done

  output wire [7:0] out;
  output wire [7:0] outbar;
//output_done

  wire [255:0] decodeOut;
  wire [255:0] decodeOutbar;
//wire_done

  decode_11 dec ( .in(in), .inbar(inbar), .out(decodeOut), .outbar(decodeOutbar) );
  encode_11 enc ( .in(decodeOut), .inbar(decodeOutbar), .out(out), .outbar(outbar) );
endmodule

module CD2_45 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD2_46 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD2_47 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD2_48 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD4_23 ( a, abar, b, bbar, y, ybar );

  input wire [3:0] a;
  input wire [3:0] b;
  input wire [3:0] abar;
  input wire [3:0] bbar;
//input_done

  output wire [15:0] y;
  output wire [15:0] ybar;
//output_done

//wire_done

  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]) );
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]) );
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]) );
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]) );
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]) );
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]) );
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]) );
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]) );
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]) );
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]) );
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]) );
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]) );
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]) );
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]) );
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]) );
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]) );
endmodule

module CD4_24 ( a, abar, b, bbar, y, ybar );

  input wire [3:0] a;
  input wire [3:0] b;
  input wire [3:0] abar;
  input wire [3:0] bbar;
//input_done

  output wire [15:0] y;
  output wire [15:0] ybar;
//output_done

//wire_done

  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]) );
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]) );
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]) );
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]) );
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]) );
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]) );
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]) );
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]) );
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]) );
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]) );
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]) );
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]) );
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]) );
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]) );
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]) );
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]) );
endmodule

module CD16_12 ( a, abar, b, bbar, y, ybar );

  input wire [15:0] a;
  input wire [15:0] b;
  input wire [15:0] abar;
  input wire [15:0] bbar;
//input_done

  output wire [255:0] y;
  output wire [255:0] ybar;
//output_done

//wire_done

  AND2_X1 U1 ( .A1(b[9]), .A2(a[0]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[9]), .A2(abar[0]), .ZN(ybar[9]) );
  AND2_X1 U2 ( .A1(b[3]), .A2(a[6]), .ZN(y[99]) );
  OR2_X1 U2bar ( .A1(bbar[3]), .A2(abar[6]), .ZN(ybar[99]) );
  AND2_X1 U3 ( .A1(b[2]), .A2(a[6]), .ZN(y[98]) );
  OR2_X1 U3bar ( .A1(bbar[2]), .A2(abar[6]), .ZN(ybar[98]) );
  AND2_X1 U4 ( .A1(b[1]), .A2(a[6]), .ZN(y[97]) );
  OR2_X1 U4bar ( .A1(bbar[1]), .A2(abar[6]), .ZN(ybar[97]) );
  AND2_X1 U5 ( .A1(b[0]), .A2(a[6]), .ZN(y[96]) );
  OR2_X1 U5bar ( .A1(bbar[0]), .A2(abar[6]), .ZN(ybar[96]) );
  AND2_X1 U6 ( .A1(b[15]), .A2(a[5]), .ZN(y[95]) );
  OR2_X1 U6bar ( .A1(bbar[15]), .A2(abar[5]), .ZN(ybar[95]) );
  AND2_X1 U7 ( .A1(b[14]), .A2(a[5]), .ZN(y[94]) );
  OR2_X1 U7bar ( .A1(bbar[14]), .A2(abar[5]), .ZN(ybar[94]) );
  AND2_X1 U8 ( .A1(b[13]), .A2(a[5]), .ZN(y[93]) );
  OR2_X1 U8bar ( .A1(bbar[13]), .A2(abar[5]), .ZN(ybar[93]) );
  AND2_X1 U9 ( .A1(b[12]), .A2(a[5]), .ZN(y[92]) );
  OR2_X1 U9bar ( .A1(bbar[12]), .A2(abar[5]), .ZN(ybar[92]) );
  AND2_X1 U10 ( .A1(b[11]), .A2(a[5]), .ZN(y[91]) );
  OR2_X1 U10bar ( .A1(bbar[11]), .A2(abar[5]), .ZN(ybar[91]) );
  AND2_X1 U11 ( .A1(b[10]), .A2(a[5]), .ZN(y[90]) );
  OR2_X1 U11bar ( .A1(bbar[10]), .A2(abar[5]), .ZN(ybar[90]) );
  AND2_X1 U12 ( .A1(b[8]), .A2(a[0]), .ZN(y[8]) );
  OR2_X1 U12bar ( .A1(bbar[8]), .A2(abar[0]), .ZN(ybar[8]) );
  AND2_X1 U13 ( .A1(a[5]), .A2(b[9]), .ZN(y[89]) );
  OR2_X1 U13bar ( .A1(abar[5]), .A2(bbar[9]), .ZN(ybar[89]) );
  AND2_X1 U14 ( .A1(b[8]), .A2(a[5]), .ZN(y[88]) );
  OR2_X1 U14bar ( .A1(bbar[8]), .A2(abar[5]), .ZN(ybar[88]) );
  AND2_X1 U15 ( .A1(b[7]), .A2(a[5]), .ZN(y[87]) );
  OR2_X1 U15bar ( .A1(bbar[7]), .A2(abar[5]), .ZN(ybar[87]) );
  AND2_X1 U16 ( .A1(b[6]), .A2(a[5]), .ZN(y[86]) );
  OR2_X1 U16bar ( .A1(bbar[6]), .A2(abar[5]), .ZN(ybar[86]) );
  AND2_X1 U17 ( .A1(b[5]), .A2(a[5]), .ZN(y[85]) );
  OR2_X1 U17bar ( .A1(bbar[5]), .A2(abar[5]), .ZN(ybar[85]) );
  AND2_X1 U18 ( .A1(b[4]), .A2(a[5]), .ZN(y[84]) );
  OR2_X1 U18bar ( .A1(bbar[4]), .A2(abar[5]), .ZN(ybar[84]) );
  AND2_X1 U19 ( .A1(a[5]), .A2(b[3]), .ZN(y[83]) );
  OR2_X1 U19bar ( .A1(abar[5]), .A2(bbar[3]), .ZN(ybar[83]) );
  AND2_X1 U20 ( .A1(a[5]), .A2(b[2]), .ZN(y[82]) );
  OR2_X1 U20bar ( .A1(abar[5]), .A2(bbar[2]), .ZN(ybar[82]) );
  AND2_X1 U21 ( .A1(a[5]), .A2(b[1]), .ZN(y[81]) );
  OR2_X1 U21bar ( .A1(abar[5]), .A2(bbar[1]), .ZN(ybar[81]) );
  AND2_X1 U22 ( .A1(a[5]), .A2(b[0]), .ZN(y[80]) );
  OR2_X1 U22bar ( .A1(abar[5]), .A2(bbar[0]), .ZN(ybar[80]) );
  AND2_X1 U23 ( .A1(b[7]), .A2(a[0]), .ZN(y[7]) );
  OR2_X1 U23bar ( .A1(bbar[7]), .A2(abar[0]), .ZN(ybar[7]) );
  AND2_X1 U24 ( .A1(a[4]), .A2(b[15]), .ZN(y[79]) );
  OR2_X1 U24bar ( .A1(abar[4]), .A2(bbar[15]), .ZN(ybar[79]) );
  AND2_X1 U25 ( .A1(a[4]), .A2(b[14]), .ZN(y[78]) );
  OR2_X1 U25bar ( .A1(abar[4]), .A2(bbar[14]), .ZN(ybar[78]) );
  AND2_X1 U26 ( .A1(a[4]), .A2(b[13]), .ZN(y[77]) );
  OR2_X1 U26bar ( .A1(abar[4]), .A2(bbar[13]), .ZN(ybar[77]) );
  AND2_X1 U27 ( .A1(a[4]), .A2(b[12]), .ZN(y[76]) );
  OR2_X1 U27bar ( .A1(abar[4]), .A2(bbar[12]), .ZN(ybar[76]) );
  AND2_X1 U28 ( .A1(a[4]), .A2(b[11]), .ZN(y[75]) );
  OR2_X1 U28bar ( .A1(abar[4]), .A2(bbar[11]), .ZN(ybar[75]) );
  AND2_X1 U29 ( .A1(a[4]), .A2(b[10]), .ZN(y[74]) );
  OR2_X1 U29bar ( .A1(abar[4]), .A2(bbar[10]), .ZN(ybar[74]) );
  AND2_X1 U30 ( .A1(a[4]), .A2(b[9]), .ZN(y[73]) );
  OR2_X1 U30bar ( .A1(abar[4]), .A2(bbar[9]), .ZN(ybar[73]) );
  AND2_X1 U31 ( .A1(a[4]), .A2(b[8]), .ZN(y[72]) );
  OR2_X1 U31bar ( .A1(abar[4]), .A2(bbar[8]), .ZN(ybar[72]) );
  AND2_X1 U32 ( .A1(a[4]), .A2(b[7]), .ZN(y[71]) );
  OR2_X1 U32bar ( .A1(abar[4]), .A2(bbar[7]), .ZN(ybar[71]) );
  AND2_X1 U33 ( .A1(a[4]), .A2(b[6]), .ZN(y[70]) );
  OR2_X1 U33bar ( .A1(abar[4]), .A2(bbar[6]), .ZN(ybar[70]) );
  AND2_X1 U34 ( .A1(b[6]), .A2(a[0]), .ZN(y[6]) );
  OR2_X1 U34bar ( .A1(bbar[6]), .A2(abar[0]), .ZN(ybar[6]) );
  AND2_X1 U35 ( .A1(a[4]), .A2(b[5]), .ZN(y[69]) );
  OR2_X1 U35bar ( .A1(abar[4]), .A2(bbar[5]), .ZN(ybar[69]) );
  AND2_X1 U36 ( .A1(a[4]), .A2(b[4]), .ZN(y[68]) );
  OR2_X1 U36bar ( .A1(abar[4]), .A2(bbar[4]), .ZN(ybar[68]) );
  AND2_X1 U37 ( .A1(a[4]), .A2(b[3]), .ZN(y[67]) );
  OR2_X1 U37bar ( .A1(abar[4]), .A2(bbar[3]), .ZN(ybar[67]) );
  AND2_X1 U38 ( .A1(a[4]), .A2(b[2]), .ZN(y[66]) );
  OR2_X1 U38bar ( .A1(abar[4]), .A2(bbar[2]), .ZN(ybar[66]) );
  AND2_X1 U39 ( .A1(a[4]), .A2(b[1]), .ZN(y[65]) );
  OR2_X1 U39bar ( .A1(abar[4]), .A2(bbar[1]), .ZN(ybar[65]) );
  AND2_X1 U40 ( .A1(a[4]), .A2(b[0]), .ZN(y[64]) );
  OR2_X1 U40bar ( .A1(abar[4]), .A2(bbar[0]), .ZN(ybar[64]) );
  AND2_X1 U41 ( .A1(a[3]), .A2(b[15]), .ZN(y[63]) );
  OR2_X1 U41bar ( .A1(abar[3]), .A2(bbar[15]), .ZN(ybar[63]) );
  AND2_X1 U42 ( .A1(a[3]), .A2(b[14]), .ZN(y[62]) );
  OR2_X1 U42bar ( .A1(abar[3]), .A2(bbar[14]), .ZN(ybar[62]) );
  AND2_X1 U43 ( .A1(a[3]), .A2(b[13]), .ZN(y[61]) );
  OR2_X1 U43bar ( .A1(abar[3]), .A2(bbar[13]), .ZN(ybar[61]) );
  AND2_X1 U44 ( .A1(a[3]), .A2(b[12]), .ZN(y[60]) );
  OR2_X1 U44bar ( .A1(abar[3]), .A2(bbar[12]), .ZN(ybar[60]) );
  AND2_X1 U45 ( .A1(b[5]), .A2(a[0]), .ZN(y[5]) );
  OR2_X1 U45bar ( .A1(bbar[5]), .A2(abar[0]), .ZN(ybar[5]) );
  AND2_X1 U46 ( .A1(a[3]), .A2(b[11]), .ZN(y[59]) );
  OR2_X1 U46bar ( .A1(abar[3]), .A2(bbar[11]), .ZN(ybar[59]) );
  AND2_X1 U47 ( .A1(a[3]), .A2(b[10]), .ZN(y[58]) );
  OR2_X1 U47bar ( .A1(abar[3]), .A2(bbar[10]), .ZN(ybar[58]) );
  AND2_X1 U48 ( .A1(a[3]), .A2(b[9]), .ZN(y[57]) );
  OR2_X1 U48bar ( .A1(abar[3]), .A2(bbar[9]), .ZN(ybar[57]) );
  AND2_X1 U49 ( .A1(a[3]), .A2(b[8]), .ZN(y[56]) );
  OR2_X1 U49bar ( .A1(abar[3]), .A2(bbar[8]), .ZN(ybar[56]) );
  AND2_X1 U50 ( .A1(a[3]), .A2(b[7]), .ZN(y[55]) );
  OR2_X1 U50bar ( .A1(abar[3]), .A2(bbar[7]), .ZN(ybar[55]) );
  AND2_X1 U51 ( .A1(a[3]), .A2(b[6]), .ZN(y[54]) );
  OR2_X1 U51bar ( .A1(abar[3]), .A2(bbar[6]), .ZN(ybar[54]) );
  AND2_X1 U52 ( .A1(a[3]), .A2(b[5]), .ZN(y[53]) );
  OR2_X1 U52bar ( .A1(abar[3]), .A2(bbar[5]), .ZN(ybar[53]) );
  AND2_X1 U53 ( .A1(a[3]), .A2(b[4]), .ZN(y[52]) );
  OR2_X1 U53bar ( .A1(abar[3]), .A2(bbar[4]), .ZN(ybar[52]) );
  AND2_X1 U54 ( .A1(a[3]), .A2(b[3]), .ZN(y[51]) );
  OR2_X1 U54bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[51]) );
  AND2_X1 U55 ( .A1(a[3]), .A2(b[2]), .ZN(y[50]) );
  OR2_X1 U55bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[50]) );
  AND2_X1 U56 ( .A1(b[4]), .A2(a[0]), .ZN(y[4]) );
  OR2_X1 U56bar ( .A1(bbar[4]), .A2(abar[0]), .ZN(ybar[4]) );
  AND2_X1 U57 ( .A1(a[3]), .A2(b[1]), .ZN(y[49]) );
  OR2_X1 U57bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[49]) );
  AND2_X1 U58 ( .A1(a[3]), .A2(b[0]), .ZN(y[48]) );
  OR2_X1 U58bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[48]) );
  AND2_X1 U59 ( .A1(a[2]), .A2(b[15]), .ZN(y[47]) );
  OR2_X1 U59bar ( .A1(abar[2]), .A2(bbar[15]), .ZN(ybar[47]) );
  AND2_X1 U60 ( .A1(a[2]), .A2(b[14]), .ZN(y[46]) );
  OR2_X1 U60bar ( .A1(abar[2]), .A2(bbar[14]), .ZN(ybar[46]) );
  AND2_X1 U61 ( .A1(a[2]), .A2(b[13]), .ZN(y[45]) );
  OR2_X1 U61bar ( .A1(abar[2]), .A2(bbar[13]), .ZN(ybar[45]) );
  AND2_X1 U62 ( .A1(a[2]), .A2(b[12]), .ZN(y[44]) );
  OR2_X1 U62bar ( .A1(abar[2]), .A2(bbar[12]), .ZN(ybar[44]) );
  AND2_X1 U63 ( .A1(a[2]), .A2(b[11]), .ZN(y[43]) );
  OR2_X1 U63bar ( .A1(abar[2]), .A2(bbar[11]), .ZN(ybar[43]) );
  AND2_X1 U64 ( .A1(a[2]), .A2(b[10]), .ZN(y[42]) );
  OR2_X1 U64bar ( .A1(abar[2]), .A2(bbar[10]), .ZN(ybar[42]) );
  AND2_X1 U65 ( .A1(a[2]), .A2(b[9]), .ZN(y[41]) );
  OR2_X1 U65bar ( .A1(abar[2]), .A2(bbar[9]), .ZN(ybar[41]) );
  AND2_X1 U66 ( .A1(a[2]), .A2(b[8]), .ZN(y[40]) );
  OR2_X1 U66bar ( .A1(abar[2]), .A2(bbar[8]), .ZN(ybar[40]) );
  AND2_X1 U67 ( .A1(b[3]), .A2(a[0]), .ZN(y[3]) );
  OR2_X1 U67bar ( .A1(bbar[3]), .A2(abar[0]), .ZN(ybar[3]) );
  AND2_X1 U68 ( .A1(a[2]), .A2(b[7]), .ZN(y[39]) );
  OR2_X1 U68bar ( .A1(abar[2]), .A2(bbar[7]), .ZN(ybar[39]) );
  AND2_X1 U69 ( .A1(a[2]), .A2(b[6]), .ZN(y[38]) );
  OR2_X1 U69bar ( .A1(abar[2]), .A2(bbar[6]), .ZN(ybar[38]) );
  AND2_X1 U70 ( .A1(a[2]), .A2(b[5]), .ZN(y[37]) );
  OR2_X1 U70bar ( .A1(abar[2]), .A2(bbar[5]), .ZN(ybar[37]) );
  AND2_X1 U71 ( .A1(a[2]), .A2(b[4]), .ZN(y[36]) );
  OR2_X1 U71bar ( .A1(abar[2]), .A2(bbar[4]), .ZN(ybar[36]) );
  AND2_X1 U72 ( .A1(a[2]), .A2(b[3]), .ZN(y[35]) );
  OR2_X1 U72bar ( .A1(abar[2]), .A2(bbar[3]), .ZN(ybar[35]) );
  AND2_X1 U73 ( .A1(a[2]), .A2(b[2]), .ZN(y[34]) );
  OR2_X1 U73bar ( .A1(abar[2]), .A2(bbar[2]), .ZN(ybar[34]) );
  AND2_X1 U74 ( .A1(a[2]), .A2(b[1]), .ZN(y[33]) );
  OR2_X1 U74bar ( .A1(abar[2]), .A2(bbar[1]), .ZN(ybar[33]) );
  AND2_X1 U75 ( .A1(a[2]), .A2(b[0]), .ZN(y[32]) );
  OR2_X1 U75bar ( .A1(abar[2]), .A2(bbar[0]), .ZN(ybar[32]) );
  AND2_X1 U76 ( .A1(a[1]), .A2(b[15]), .ZN(y[31]) );
  OR2_X1 U76bar ( .A1(abar[1]), .A2(bbar[15]), .ZN(ybar[31]) );
  AND2_X1 U77 ( .A1(a[1]), .A2(b[14]), .ZN(y[30]) );
  OR2_X1 U77bar ( .A1(abar[1]), .A2(bbar[14]), .ZN(ybar[30]) );
  AND2_X1 U78 ( .A1(b[2]), .A2(a[0]), .ZN(y[2]) );
  OR2_X1 U78bar ( .A1(bbar[2]), .A2(abar[0]), .ZN(ybar[2]) );
  AND2_X1 U79 ( .A1(a[1]), .A2(b[13]), .ZN(y[29]) );
  OR2_X1 U79bar ( .A1(abar[1]), .A2(bbar[13]), .ZN(ybar[29]) );
  AND2_X1 U80 ( .A1(a[1]), .A2(b[12]), .ZN(y[28]) );
  OR2_X1 U80bar ( .A1(abar[1]), .A2(bbar[12]), .ZN(ybar[28]) );
  AND2_X1 U81 ( .A1(a[1]), .A2(b[11]), .ZN(y[27]) );
  OR2_X1 U81bar ( .A1(abar[1]), .A2(bbar[11]), .ZN(ybar[27]) );
  AND2_X1 U82 ( .A1(a[1]), .A2(b[10]), .ZN(y[26]) );
  OR2_X1 U82bar ( .A1(abar[1]), .A2(bbar[10]), .ZN(ybar[26]) );
  AND2_X1 U83 ( .A1(a[1]), .A2(b[9]), .ZN(y[25]) );
  OR2_X1 U83bar ( .A1(abar[1]), .A2(bbar[9]), .ZN(ybar[25]) );
  AND2_X1 U84 ( .A1(a[15]), .A2(b[15]), .ZN(y[255]) );
  OR2_X1 U84bar ( .A1(abar[15]), .A2(bbar[15]), .ZN(ybar[255]) );
  AND2_X1 U85 ( .A1(a[15]), .A2(b[14]), .ZN(y[254]) );
  OR2_X1 U85bar ( .A1(abar[15]), .A2(bbar[14]), .ZN(ybar[254]) );
  AND2_X1 U86 ( .A1(a[15]), .A2(b[13]), .ZN(y[253]) );
  OR2_X1 U86bar ( .A1(abar[15]), .A2(bbar[13]), .ZN(ybar[253]) );
  AND2_X1 U87 ( .A1(a[15]), .A2(b[12]), .ZN(y[252]) );
  OR2_X1 U87bar ( .A1(abar[15]), .A2(bbar[12]), .ZN(ybar[252]) );
  AND2_X1 U88 ( .A1(a[15]), .A2(b[11]), .ZN(y[251]) );
  OR2_X1 U88bar ( .A1(abar[15]), .A2(bbar[11]), .ZN(ybar[251]) );
  AND2_X1 U89 ( .A1(a[15]), .A2(b[10]), .ZN(y[250]) );
  OR2_X1 U89bar ( .A1(abar[15]), .A2(bbar[10]), .ZN(ybar[250]) );
  AND2_X1 U90 ( .A1(a[1]), .A2(b[8]), .ZN(y[24]) );
  OR2_X1 U90bar ( .A1(abar[1]), .A2(bbar[8]), .ZN(ybar[24]) );
  AND2_X1 U91 ( .A1(a[15]), .A2(b[9]), .ZN(y[249]) );
  OR2_X1 U91bar ( .A1(abar[15]), .A2(bbar[9]), .ZN(ybar[249]) );
  AND2_X1 U92 ( .A1(a[15]), .A2(b[8]), .ZN(y[248]) );
  OR2_X1 U92bar ( .A1(abar[15]), .A2(bbar[8]), .ZN(ybar[248]) );
  AND2_X1 U93 ( .A1(a[15]), .A2(b[7]), .ZN(y[247]) );
  OR2_X1 U93bar ( .A1(abar[15]), .A2(bbar[7]), .ZN(ybar[247]) );
  AND2_X1 U94 ( .A1(a[15]), .A2(b[6]), .ZN(y[246]) );
  OR2_X1 U94bar ( .A1(abar[15]), .A2(bbar[6]), .ZN(ybar[246]) );
  AND2_X1 U95 ( .A1(a[15]), .A2(b[5]), .ZN(y[245]) );
  OR2_X1 U95bar ( .A1(abar[15]), .A2(bbar[5]), .ZN(ybar[245]) );
  AND2_X1 U96 ( .A1(a[15]), .A2(b[4]), .ZN(y[244]) );
  OR2_X1 U96bar ( .A1(abar[15]), .A2(bbar[4]), .ZN(ybar[244]) );
  AND2_X1 U97 ( .A1(a[15]), .A2(b[3]), .ZN(y[243]) );
  OR2_X1 U97bar ( .A1(abar[15]), .A2(bbar[3]), .ZN(ybar[243]) );
  AND2_X1 U98 ( .A1(a[15]), .A2(b[2]), .ZN(y[242]) );
  OR2_X1 U98bar ( .A1(abar[15]), .A2(bbar[2]), .ZN(ybar[242]) );
  AND2_X1 U99 ( .A1(a[15]), .A2(b[1]), .ZN(y[241]) );
  OR2_X1 U99bar ( .A1(abar[15]), .A2(bbar[1]), .ZN(ybar[241]) );
  AND2_X1 U100 ( .A1(a[15]), .A2(b[0]), .ZN(y[240]) );
  OR2_X1 U100bar ( .A1(abar[15]), .A2(bbar[0]), .ZN(ybar[240]) );
  AND2_X1 U101 ( .A1(a[1]), .A2(b[7]), .ZN(y[23]) );
  OR2_X1 U101bar ( .A1(abar[1]), .A2(bbar[7]), .ZN(ybar[23]) );
  AND2_X1 U102 ( .A1(a[14]), .A2(b[15]), .ZN(y[239]) );
  OR2_X1 U102bar ( .A1(abar[14]), .A2(bbar[15]), .ZN(ybar[239]) );
  AND2_X1 U103 ( .A1(a[14]), .A2(b[14]), .ZN(y[238]) );
  OR2_X1 U103bar ( .A1(abar[14]), .A2(bbar[14]), .ZN(ybar[238]) );
  AND2_X1 U104 ( .A1(a[14]), .A2(b[13]), .ZN(y[237]) );
  OR2_X1 U104bar ( .A1(abar[14]), .A2(bbar[13]), .ZN(ybar[237]) );
  AND2_X1 U105 ( .A1(a[14]), .A2(b[12]), .ZN(y[236]) );
  OR2_X1 U105bar ( .A1(abar[14]), .A2(bbar[12]), .ZN(ybar[236]) );
  AND2_X1 U106 ( .A1(a[14]), .A2(b[11]), .ZN(y[235]) );
  OR2_X1 U106bar ( .A1(abar[14]), .A2(bbar[11]), .ZN(ybar[235]) );
  AND2_X1 U107 ( .A1(a[14]), .A2(b[10]), .ZN(y[234]) );
  OR2_X1 U107bar ( .A1(abar[14]), .A2(bbar[10]), .ZN(ybar[234]) );
  AND2_X1 U108 ( .A1(a[14]), .A2(b[9]), .ZN(y[233]) );
  OR2_X1 U108bar ( .A1(abar[14]), .A2(bbar[9]), .ZN(ybar[233]) );
  AND2_X1 U109 ( .A1(a[14]), .A2(b[8]), .ZN(y[232]) );
  OR2_X1 U109bar ( .A1(abar[14]), .A2(bbar[8]), .ZN(ybar[232]) );
  AND2_X1 U110 ( .A1(a[14]), .A2(b[7]), .ZN(y[231]) );
  OR2_X1 U110bar ( .A1(abar[14]), .A2(bbar[7]), .ZN(ybar[231]) );
  AND2_X1 U111 ( .A1(a[14]), .A2(b[6]), .ZN(y[230]) );
  OR2_X1 U111bar ( .A1(abar[14]), .A2(bbar[6]), .ZN(ybar[230]) );
  AND2_X1 U112 ( .A1(a[1]), .A2(b[6]), .ZN(y[22]) );
  OR2_X1 U112bar ( .A1(abar[1]), .A2(bbar[6]), .ZN(ybar[22]) );
  AND2_X1 U113 ( .A1(a[14]), .A2(b[5]), .ZN(y[229]) );
  OR2_X1 U113bar ( .A1(abar[14]), .A2(bbar[5]), .ZN(ybar[229]) );
  AND2_X1 U114 ( .A1(a[14]), .A2(b[4]), .ZN(y[228]) );
  OR2_X1 U114bar ( .A1(abar[14]), .A2(bbar[4]), .ZN(ybar[228]) );
  AND2_X1 U115 ( .A1(a[14]), .A2(b[3]), .ZN(y[227]) );
  OR2_X1 U115bar ( .A1(abar[14]), .A2(bbar[3]), .ZN(ybar[227]) );
  AND2_X1 U116 ( .A1(a[14]), .A2(b[2]), .ZN(y[226]) );
  OR2_X1 U116bar ( .A1(abar[14]), .A2(bbar[2]), .ZN(ybar[226]) );
  AND2_X1 U117 ( .A1(a[14]), .A2(b[1]), .ZN(y[225]) );
  OR2_X1 U117bar ( .A1(abar[14]), .A2(bbar[1]), .ZN(ybar[225]) );
  AND2_X1 U118 ( .A1(a[14]), .A2(b[0]), .ZN(y[224]) );
  OR2_X1 U118bar ( .A1(abar[14]), .A2(bbar[0]), .ZN(ybar[224]) );
  AND2_X1 U119 ( .A1(a[13]), .A2(b[15]), .ZN(y[223]) );
  OR2_X1 U119bar ( .A1(abar[13]), .A2(bbar[15]), .ZN(ybar[223]) );
  AND2_X1 U120 ( .A1(a[13]), .A2(b[14]), .ZN(y[222]) );
  OR2_X1 U120bar ( .A1(abar[13]), .A2(bbar[14]), .ZN(ybar[222]) );
  AND2_X1 U121 ( .A1(a[13]), .A2(b[13]), .ZN(y[221]) );
  OR2_X1 U121bar ( .A1(abar[13]), .A2(bbar[13]), .ZN(ybar[221]) );
  AND2_X1 U122 ( .A1(a[13]), .A2(b[12]), .ZN(y[220]) );
  OR2_X1 U122bar ( .A1(abar[13]), .A2(bbar[12]), .ZN(ybar[220]) );
  AND2_X1 U123 ( .A1(a[1]), .A2(b[5]), .ZN(y[21]) );
  OR2_X1 U123bar ( .A1(abar[1]), .A2(bbar[5]), .ZN(ybar[21]) );
  AND2_X1 U124 ( .A1(a[13]), .A2(b[11]), .ZN(y[219]) );
  OR2_X1 U124bar ( .A1(abar[13]), .A2(bbar[11]), .ZN(ybar[219]) );
  AND2_X1 U125 ( .A1(a[13]), .A2(b[10]), .ZN(y[218]) );
  OR2_X1 U125bar ( .A1(abar[13]), .A2(bbar[10]), .ZN(ybar[218]) );
  AND2_X1 U126 ( .A1(a[13]), .A2(b[9]), .ZN(y[217]) );
  OR2_X1 U126bar ( .A1(abar[13]), .A2(bbar[9]), .ZN(ybar[217]) );
  AND2_X1 U127 ( .A1(a[13]), .A2(b[8]), .ZN(y[216]) );
  OR2_X1 U127bar ( .A1(abar[13]), .A2(bbar[8]), .ZN(ybar[216]) );
  AND2_X1 U128 ( .A1(a[13]), .A2(b[7]), .ZN(y[215]) );
  OR2_X1 U128bar ( .A1(abar[13]), .A2(bbar[7]), .ZN(ybar[215]) );
  AND2_X1 U129 ( .A1(a[13]), .A2(b[6]), .ZN(y[214]) );
  OR2_X1 U129bar ( .A1(abar[13]), .A2(bbar[6]), .ZN(ybar[214]) );
  AND2_X1 U130 ( .A1(a[13]), .A2(b[5]), .ZN(y[213]) );
  OR2_X1 U130bar ( .A1(abar[13]), .A2(bbar[5]), .ZN(ybar[213]) );
  AND2_X1 U131 ( .A1(a[13]), .A2(b[4]), .ZN(y[212]) );
  OR2_X1 U131bar ( .A1(abar[13]), .A2(bbar[4]), .ZN(ybar[212]) );
  AND2_X1 U132 ( .A1(a[13]), .A2(b[3]), .ZN(y[211]) );
  OR2_X1 U132bar ( .A1(abar[13]), .A2(bbar[3]), .ZN(ybar[211]) );
  AND2_X1 U133 ( .A1(a[13]), .A2(b[2]), .ZN(y[210]) );
  OR2_X1 U133bar ( .A1(abar[13]), .A2(bbar[2]), .ZN(ybar[210]) );
  AND2_X1 U134 ( .A1(a[1]), .A2(b[4]), .ZN(y[20]) );
  OR2_X1 U134bar ( .A1(abar[1]), .A2(bbar[4]), .ZN(ybar[20]) );
  AND2_X1 U135 ( .A1(a[13]), .A2(b[1]), .ZN(y[209]) );
  OR2_X1 U135bar ( .A1(abar[13]), .A2(bbar[1]), .ZN(ybar[209]) );
  AND2_X1 U136 ( .A1(a[13]), .A2(b[0]), .ZN(y[208]) );
  OR2_X1 U136bar ( .A1(abar[13]), .A2(bbar[0]), .ZN(ybar[208]) );
  AND2_X1 U137 ( .A1(a[12]), .A2(b[15]), .ZN(y[207]) );
  OR2_X1 U137bar ( .A1(abar[12]), .A2(bbar[15]), .ZN(ybar[207]) );
  AND2_X1 U138 ( .A1(a[12]), .A2(b[14]), .ZN(y[206]) );
  OR2_X1 U138bar ( .A1(abar[12]), .A2(bbar[14]), .ZN(ybar[206]) );
  AND2_X1 U139 ( .A1(a[12]), .A2(b[13]), .ZN(y[205]) );
  OR2_X1 U139bar ( .A1(abar[12]), .A2(bbar[13]), .ZN(ybar[205]) );
  AND2_X1 U140 ( .A1(a[12]), .A2(b[12]), .ZN(y[204]) );
  OR2_X1 U140bar ( .A1(abar[12]), .A2(bbar[12]), .ZN(ybar[204]) );
  AND2_X1 U141 ( .A1(a[12]), .A2(b[11]), .ZN(y[203]) );
  OR2_X1 U141bar ( .A1(abar[12]), .A2(bbar[11]), .ZN(ybar[203]) );
  AND2_X1 U142 ( .A1(a[12]), .A2(b[10]), .ZN(y[202]) );
  OR2_X1 U142bar ( .A1(abar[12]), .A2(bbar[10]), .ZN(ybar[202]) );
  AND2_X1 U143 ( .A1(a[12]), .A2(b[9]), .ZN(y[201]) );
  OR2_X1 U143bar ( .A1(abar[12]), .A2(bbar[9]), .ZN(ybar[201]) );
  AND2_X1 U144 ( .A1(a[12]), .A2(b[8]), .ZN(y[200]) );
  OR2_X1 U144bar ( .A1(abar[12]), .A2(bbar[8]), .ZN(ybar[200]) );
  AND2_X1 U145 ( .A1(b[1]), .A2(a[0]), .ZN(y[1]) );
  OR2_X1 U145bar ( .A1(bbar[1]), .A2(abar[0]), .ZN(ybar[1]) );
  AND2_X1 U146 ( .A1(a[1]), .A2(b[3]), .ZN(y[19]) );
  OR2_X1 U146bar ( .A1(abar[1]), .A2(bbar[3]), .ZN(ybar[19]) );
  AND2_X1 U147 ( .A1(a[12]), .A2(b[7]), .ZN(y[199]) );
  OR2_X1 U147bar ( .A1(abar[12]), .A2(bbar[7]), .ZN(ybar[199]) );
  AND2_X1 U148 ( .A1(a[12]), .A2(b[6]), .ZN(y[198]) );
  OR2_X1 U148bar ( .A1(abar[12]), .A2(bbar[6]), .ZN(ybar[198]) );
  AND2_X1 U149 ( .A1(a[12]), .A2(b[5]), .ZN(y[197]) );
  OR2_X1 U149bar ( .A1(abar[12]), .A2(bbar[5]), .ZN(ybar[197]) );
  AND2_X1 U150 ( .A1(a[12]), .A2(b[4]), .ZN(y[196]) );
  OR2_X1 U150bar ( .A1(abar[12]), .A2(bbar[4]), .ZN(ybar[196]) );
  AND2_X1 U151 ( .A1(a[12]), .A2(b[3]), .ZN(y[195]) );
  OR2_X1 U151bar ( .A1(abar[12]), .A2(bbar[3]), .ZN(ybar[195]) );
  AND2_X1 U152 ( .A1(a[12]), .A2(b[2]), .ZN(y[194]) );
  OR2_X1 U152bar ( .A1(abar[12]), .A2(bbar[2]), .ZN(ybar[194]) );
  AND2_X1 U153 ( .A1(a[12]), .A2(b[1]), .ZN(y[193]) );
  OR2_X1 U153bar ( .A1(abar[12]), .A2(bbar[1]), .ZN(ybar[193]) );
  AND2_X1 U154 ( .A1(a[12]), .A2(b[0]), .ZN(y[192]) );
  OR2_X1 U154bar ( .A1(abar[12]), .A2(bbar[0]), .ZN(ybar[192]) );
  AND2_X1 U155 ( .A1(a[11]), .A2(b[15]), .ZN(y[191]) );
  OR2_X1 U155bar ( .A1(abar[11]), .A2(bbar[15]), .ZN(ybar[191]) );
  AND2_X1 U156 ( .A1(a[11]), .A2(b[14]), .ZN(y[190]) );
  OR2_X1 U156bar ( .A1(abar[11]), .A2(bbar[14]), .ZN(ybar[190]) );
  AND2_X1 U157 ( .A1(a[1]), .A2(b[2]), .ZN(y[18]) );
  OR2_X1 U157bar ( .A1(abar[1]), .A2(bbar[2]), .ZN(ybar[18]) );
  AND2_X1 U158 ( .A1(a[11]), .A2(b[13]), .ZN(y[189]) );
  OR2_X1 U158bar ( .A1(abar[11]), .A2(bbar[13]), .ZN(ybar[189]) );
  AND2_X1 U159 ( .A1(a[11]), .A2(b[12]), .ZN(y[188]) );
  OR2_X1 U159bar ( .A1(abar[11]), .A2(bbar[12]), .ZN(ybar[188]) );
  AND2_X1 U160 ( .A1(a[11]), .A2(b[11]), .ZN(y[187]) );
  OR2_X1 U160bar ( .A1(abar[11]), .A2(bbar[11]), .ZN(ybar[187]) );
  AND2_X1 U161 ( .A1(a[11]), .A2(b[10]), .ZN(y[186]) );
  OR2_X1 U161bar ( .A1(abar[11]), .A2(bbar[10]), .ZN(ybar[186]) );
  AND2_X1 U162 ( .A1(a[11]), .A2(b[9]), .ZN(y[185]) );
  OR2_X1 U162bar ( .A1(abar[11]), .A2(bbar[9]), .ZN(ybar[185]) );
  AND2_X1 U163 ( .A1(a[11]), .A2(b[8]), .ZN(y[184]) );
  OR2_X1 U163bar ( .A1(abar[11]), .A2(bbar[8]), .ZN(ybar[184]) );
  AND2_X1 U164 ( .A1(a[11]), .A2(b[7]), .ZN(y[183]) );
  OR2_X1 U164bar ( .A1(abar[11]), .A2(bbar[7]), .ZN(ybar[183]) );
  AND2_X1 U165 ( .A1(a[11]), .A2(b[6]), .ZN(y[182]) );
  OR2_X1 U165bar ( .A1(abar[11]), .A2(bbar[6]), .ZN(ybar[182]) );
  AND2_X1 U166 ( .A1(a[11]), .A2(b[5]), .ZN(y[181]) );
  OR2_X1 U166bar ( .A1(abar[11]), .A2(bbar[5]), .ZN(ybar[181]) );
  AND2_X1 U167 ( .A1(a[11]), .A2(b[4]), .ZN(y[180]) );
  OR2_X1 U167bar ( .A1(abar[11]), .A2(bbar[4]), .ZN(ybar[180]) );
  AND2_X1 U168 ( .A1(a[1]), .A2(b[1]), .ZN(y[17]) );
  OR2_X1 U168bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[17]) );
  AND2_X1 U169 ( .A1(a[11]), .A2(b[3]), .ZN(y[179]) );
  OR2_X1 U169bar ( .A1(abar[11]), .A2(bbar[3]), .ZN(ybar[179]) );
  AND2_X1 U170 ( .A1(a[11]), .A2(b[2]), .ZN(y[178]) );
  OR2_X1 U170bar ( .A1(abar[11]), .A2(bbar[2]), .ZN(ybar[178]) );
  AND2_X1 U171 ( .A1(a[11]), .A2(b[1]), .ZN(y[177]) );
  OR2_X1 U171bar ( .A1(abar[11]), .A2(bbar[1]), .ZN(ybar[177]) );
  AND2_X1 U172 ( .A1(a[11]), .A2(b[0]), .ZN(y[176]) );
  OR2_X1 U172bar ( .A1(abar[11]), .A2(bbar[0]), .ZN(ybar[176]) );
  AND2_X1 U173 ( .A1(a[10]), .A2(b[15]), .ZN(y[175]) );
  OR2_X1 U173bar ( .A1(abar[10]), .A2(bbar[15]), .ZN(ybar[175]) );
  AND2_X1 U174 ( .A1(a[10]), .A2(b[14]), .ZN(y[174]) );
  OR2_X1 U174bar ( .A1(abar[10]), .A2(bbar[14]), .ZN(ybar[174]) );
  AND2_X1 U175 ( .A1(a[10]), .A2(b[13]), .ZN(y[173]) );
  OR2_X1 U175bar ( .A1(abar[10]), .A2(bbar[13]), .ZN(ybar[173]) );
  AND2_X1 U176 ( .A1(a[10]), .A2(b[12]), .ZN(y[172]) );
  OR2_X1 U176bar ( .A1(abar[10]), .A2(bbar[12]), .ZN(ybar[172]) );
  AND2_X1 U177 ( .A1(a[10]), .A2(b[11]), .ZN(y[171]) );
  OR2_X1 U177bar ( .A1(abar[10]), .A2(bbar[11]), .ZN(ybar[171]) );
  AND2_X1 U178 ( .A1(a[10]), .A2(b[10]), .ZN(y[170]) );
  OR2_X1 U178bar ( .A1(abar[10]), .A2(bbar[10]), .ZN(ybar[170]) );
  AND2_X1 U179 ( .A1(a[1]), .A2(b[0]), .ZN(y[16]) );
  OR2_X1 U179bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[16]) );
  AND2_X1 U180 ( .A1(a[10]), .A2(b[9]), .ZN(y[169]) );
  OR2_X1 U180bar ( .A1(abar[10]), .A2(bbar[9]), .ZN(ybar[169]) );
  AND2_X1 U181 ( .A1(a[10]), .A2(b[8]), .ZN(y[168]) );
  OR2_X1 U181bar ( .A1(abar[10]), .A2(bbar[8]), .ZN(ybar[168]) );
  AND2_X1 U182 ( .A1(a[10]), .A2(b[7]), .ZN(y[167]) );
  OR2_X1 U182bar ( .A1(abar[10]), .A2(bbar[7]), .ZN(ybar[167]) );
  AND2_X1 U183 ( .A1(a[10]), .A2(b[6]), .ZN(y[166]) );
  OR2_X1 U183bar ( .A1(abar[10]), .A2(bbar[6]), .ZN(ybar[166]) );
  AND2_X1 U184 ( .A1(a[10]), .A2(b[5]), .ZN(y[165]) );
  OR2_X1 U184bar ( .A1(abar[10]), .A2(bbar[5]), .ZN(ybar[165]) );
  AND2_X1 U185 ( .A1(a[10]), .A2(b[4]), .ZN(y[164]) );
  OR2_X1 U185bar ( .A1(abar[10]), .A2(bbar[4]), .ZN(ybar[164]) );
  AND2_X1 U186 ( .A1(a[10]), .A2(b[3]), .ZN(y[163]) );
  OR2_X1 U186bar ( .A1(abar[10]), .A2(bbar[3]), .ZN(ybar[163]) );
  AND2_X1 U187 ( .A1(a[10]), .A2(b[2]), .ZN(y[162]) );
  OR2_X1 U187bar ( .A1(abar[10]), .A2(bbar[2]), .ZN(ybar[162]) );
  AND2_X1 U188 ( .A1(a[10]), .A2(b[1]), .ZN(y[161]) );
  OR2_X1 U188bar ( .A1(abar[10]), .A2(bbar[1]), .ZN(ybar[161]) );
  AND2_X1 U189 ( .A1(a[10]), .A2(b[0]), .ZN(y[160]) );
  OR2_X1 U189bar ( .A1(abar[10]), .A2(bbar[0]), .ZN(ybar[160]) );
  AND2_X1 U190 ( .A1(b[15]), .A2(a[0]), .ZN(y[15]) );
  OR2_X1 U190bar ( .A1(bbar[15]), .A2(abar[0]), .ZN(ybar[15]) );
  AND2_X1 U191 ( .A1(a[9]), .A2(b[15]), .ZN(y[159]) );
  OR2_X1 U191bar ( .A1(abar[9]), .A2(bbar[15]), .ZN(ybar[159]) );
  AND2_X1 U192 ( .A1(a[9]), .A2(b[14]), .ZN(y[158]) );
  OR2_X1 U192bar ( .A1(abar[9]), .A2(bbar[14]), .ZN(ybar[158]) );
  AND2_X1 U193 ( .A1(a[9]), .A2(b[13]), .ZN(y[157]) );
  OR2_X1 U193bar ( .A1(abar[9]), .A2(bbar[13]), .ZN(ybar[157]) );
  AND2_X1 U194 ( .A1(a[9]), .A2(b[12]), .ZN(y[156]) );
  OR2_X1 U194bar ( .A1(abar[9]), .A2(bbar[12]), .ZN(ybar[156]) );
  AND2_X1 U195 ( .A1(a[9]), .A2(b[11]), .ZN(y[155]) );
  OR2_X1 U195bar ( .A1(abar[9]), .A2(bbar[11]), .ZN(ybar[155]) );
  AND2_X1 U196 ( .A1(a[9]), .A2(b[10]), .ZN(y[154]) );
  OR2_X1 U196bar ( .A1(abar[9]), .A2(bbar[10]), .ZN(ybar[154]) );
  AND2_X1 U197 ( .A1(a[9]), .A2(b[9]), .ZN(y[153]) );
  OR2_X1 U197bar ( .A1(abar[9]), .A2(bbar[9]), .ZN(ybar[153]) );
  AND2_X1 U198 ( .A1(a[9]), .A2(b[8]), .ZN(y[152]) );
  OR2_X1 U198bar ( .A1(abar[9]), .A2(bbar[8]), .ZN(ybar[152]) );
  AND2_X1 U199 ( .A1(a[9]), .A2(b[7]), .ZN(y[151]) );
  OR2_X1 U199bar ( .A1(abar[9]), .A2(bbar[7]), .ZN(ybar[151]) );
  AND2_X1 U200 ( .A1(a[9]), .A2(b[6]), .ZN(y[150]) );
  OR2_X1 U200bar ( .A1(abar[9]), .A2(bbar[6]), .ZN(ybar[150]) );
  AND2_X1 U201 ( .A1(b[14]), .A2(a[0]), .ZN(y[14]) );
  OR2_X1 U201bar ( .A1(bbar[14]), .A2(abar[0]), .ZN(ybar[14]) );
  AND2_X1 U202 ( .A1(a[9]), .A2(b[5]), .ZN(y[149]) );
  OR2_X1 U202bar ( .A1(abar[9]), .A2(bbar[5]), .ZN(ybar[149]) );
  AND2_X1 U203 ( .A1(a[9]), .A2(b[4]), .ZN(y[148]) );
  OR2_X1 U203bar ( .A1(abar[9]), .A2(bbar[4]), .ZN(ybar[148]) );
  AND2_X1 U204 ( .A1(a[9]), .A2(b[3]), .ZN(y[147]) );
  OR2_X1 U204bar ( .A1(abar[9]), .A2(bbar[3]), .ZN(ybar[147]) );
  AND2_X1 U205 ( .A1(a[9]), .A2(b[2]), .ZN(y[146]) );
  OR2_X1 U205bar ( .A1(abar[9]), .A2(bbar[2]), .ZN(ybar[146]) );
  AND2_X1 U206 ( .A1(a[9]), .A2(b[1]), .ZN(y[145]) );
  OR2_X1 U206bar ( .A1(abar[9]), .A2(bbar[1]), .ZN(ybar[145]) );
  AND2_X1 U207 ( .A1(a[9]), .A2(b[0]), .ZN(y[144]) );
  OR2_X1 U207bar ( .A1(abar[9]), .A2(bbar[0]), .ZN(ybar[144]) );
  AND2_X1 U208 ( .A1(a[8]), .A2(b[15]), .ZN(y[143]) );
  OR2_X1 U208bar ( .A1(abar[8]), .A2(bbar[15]), .ZN(ybar[143]) );
  AND2_X1 U209 ( .A1(a[8]), .A2(b[14]), .ZN(y[142]) );
  OR2_X1 U209bar ( .A1(abar[8]), .A2(bbar[14]), .ZN(ybar[142]) );
  AND2_X1 U210 ( .A1(a[8]), .A2(b[13]), .ZN(y[141]) );
  OR2_X1 U210bar ( .A1(abar[8]), .A2(bbar[13]), .ZN(ybar[141]) );
  AND2_X1 U211 ( .A1(a[8]), .A2(b[12]), .ZN(y[140]) );
  OR2_X1 U211bar ( .A1(abar[8]), .A2(bbar[12]), .ZN(ybar[140]) );
  AND2_X1 U212 ( .A1(b[13]), .A2(a[0]), .ZN(y[13]) );
  OR2_X1 U212bar ( .A1(bbar[13]), .A2(abar[0]), .ZN(ybar[13]) );
  AND2_X1 U213 ( .A1(a[8]), .A2(b[11]), .ZN(y[139]) );
  OR2_X1 U213bar ( .A1(abar[8]), .A2(bbar[11]), .ZN(ybar[139]) );
  AND2_X1 U214 ( .A1(a[8]), .A2(b[10]), .ZN(y[138]) );
  OR2_X1 U214bar ( .A1(abar[8]), .A2(bbar[10]), .ZN(ybar[138]) );
  AND2_X1 U215 ( .A1(a[8]), .A2(b[9]), .ZN(y[137]) );
  OR2_X1 U215bar ( .A1(abar[8]), .A2(bbar[9]), .ZN(ybar[137]) );
  AND2_X1 U216 ( .A1(a[8]), .A2(b[8]), .ZN(y[136]) );
  OR2_X1 U216bar ( .A1(abar[8]), .A2(bbar[8]), .ZN(ybar[136]) );
  AND2_X1 U217 ( .A1(a[8]), .A2(b[7]), .ZN(y[135]) );
  OR2_X1 U217bar ( .A1(abar[8]), .A2(bbar[7]), .ZN(ybar[135]) );
  AND2_X1 U218 ( .A1(a[8]), .A2(b[6]), .ZN(y[134]) );
  OR2_X1 U218bar ( .A1(abar[8]), .A2(bbar[6]), .ZN(ybar[134]) );
  AND2_X1 U219 ( .A1(a[8]), .A2(b[5]), .ZN(y[133]) );
  OR2_X1 U219bar ( .A1(abar[8]), .A2(bbar[5]), .ZN(ybar[133]) );
  AND2_X1 U220 ( .A1(a[8]), .A2(b[4]), .ZN(y[132]) );
  OR2_X1 U220bar ( .A1(abar[8]), .A2(bbar[4]), .ZN(ybar[132]) );
  AND2_X1 U221 ( .A1(a[8]), .A2(b[3]), .ZN(y[131]) );
  OR2_X1 U221bar ( .A1(abar[8]), .A2(bbar[3]), .ZN(ybar[131]) );
  AND2_X1 U222 ( .A1(a[8]), .A2(b[2]), .ZN(y[130]) );
  OR2_X1 U222bar ( .A1(abar[8]), .A2(bbar[2]), .ZN(ybar[130]) );
  AND2_X1 U223 ( .A1(b[12]), .A2(a[0]), .ZN(y[12]) );
  OR2_X1 U223bar ( .A1(bbar[12]), .A2(abar[0]), .ZN(ybar[12]) );
  AND2_X1 U224 ( .A1(a[8]), .A2(b[1]), .ZN(y[129]) );
  OR2_X1 U224bar ( .A1(abar[8]), .A2(bbar[1]), .ZN(ybar[129]) );
  AND2_X1 U225 ( .A1(a[8]), .A2(b[0]), .ZN(y[128]) );
  OR2_X1 U225bar ( .A1(abar[8]), .A2(bbar[0]), .ZN(ybar[128]) );
  AND2_X1 U226 ( .A1(a[7]), .A2(b[15]), .ZN(y[127]) );
  OR2_X1 U226bar ( .A1(abar[7]), .A2(bbar[15]), .ZN(ybar[127]) );
  AND2_X1 U227 ( .A1(a[7]), .A2(b[14]), .ZN(y[126]) );
  OR2_X1 U227bar ( .A1(abar[7]), .A2(bbar[14]), .ZN(ybar[126]) );
  AND2_X1 U228 ( .A1(a[7]), .A2(b[13]), .ZN(y[125]) );
  OR2_X1 U228bar ( .A1(abar[7]), .A2(bbar[13]), .ZN(ybar[125]) );
  AND2_X1 U229 ( .A1(a[7]), .A2(b[12]), .ZN(y[124]) );
  OR2_X1 U229bar ( .A1(abar[7]), .A2(bbar[12]), .ZN(ybar[124]) );
  AND2_X1 U230 ( .A1(a[7]), .A2(b[11]), .ZN(y[123]) );
  OR2_X1 U230bar ( .A1(abar[7]), .A2(bbar[11]), .ZN(ybar[123]) );
  AND2_X1 U231 ( .A1(a[7]), .A2(b[10]), .ZN(y[122]) );
  OR2_X1 U231bar ( .A1(abar[7]), .A2(bbar[10]), .ZN(ybar[122]) );
  AND2_X1 U232 ( .A1(a[7]), .A2(b[9]), .ZN(y[121]) );
  OR2_X1 U232bar ( .A1(abar[7]), .A2(bbar[9]), .ZN(ybar[121]) );
  AND2_X1 U233 ( .A1(a[7]), .A2(b[8]), .ZN(y[120]) );
  OR2_X1 U233bar ( .A1(abar[7]), .A2(bbar[8]), .ZN(ybar[120]) );
  AND2_X1 U234 ( .A1(b[11]), .A2(a[0]), .ZN(y[11]) );
  OR2_X1 U234bar ( .A1(bbar[11]), .A2(abar[0]), .ZN(ybar[11]) );
  AND2_X1 U235 ( .A1(a[7]), .A2(b[7]), .ZN(y[119]) );
  OR2_X1 U235bar ( .A1(abar[7]), .A2(bbar[7]), .ZN(ybar[119]) );
  AND2_X1 U236 ( .A1(a[7]), .A2(b[6]), .ZN(y[118]) );
  OR2_X1 U236bar ( .A1(abar[7]), .A2(bbar[6]), .ZN(ybar[118]) );
  AND2_X1 U237 ( .A1(a[7]), .A2(b[5]), .ZN(y[117]) );
  OR2_X1 U237bar ( .A1(abar[7]), .A2(bbar[5]), .ZN(ybar[117]) );
  AND2_X1 U238 ( .A1(a[7]), .A2(b[4]), .ZN(y[116]) );
  OR2_X1 U238bar ( .A1(abar[7]), .A2(bbar[4]), .ZN(ybar[116]) );
  AND2_X1 U239 ( .A1(a[7]), .A2(b[3]), .ZN(y[115]) );
  OR2_X1 U239bar ( .A1(abar[7]), .A2(bbar[3]), .ZN(ybar[115]) );
  AND2_X1 U240 ( .A1(a[7]), .A2(b[2]), .ZN(y[114]) );
  OR2_X1 U240bar ( .A1(abar[7]), .A2(bbar[2]), .ZN(ybar[114]) );
  AND2_X1 U241 ( .A1(a[7]), .A2(b[1]), .ZN(y[113]) );
  OR2_X1 U241bar ( .A1(abar[7]), .A2(bbar[1]), .ZN(ybar[113]) );
  AND2_X1 U242 ( .A1(a[7]), .A2(b[0]), .ZN(y[112]) );
  OR2_X1 U242bar ( .A1(abar[7]), .A2(bbar[0]), .ZN(ybar[112]) );
  AND2_X1 U243 ( .A1(b[15]), .A2(a[6]), .ZN(y[111]) );
  OR2_X1 U243bar ( .A1(bbar[15]), .A2(abar[6]), .ZN(ybar[111]) );
  AND2_X1 U244 ( .A1(b[14]), .A2(a[6]), .ZN(y[110]) );
  OR2_X1 U244bar ( .A1(bbar[14]), .A2(abar[6]), .ZN(ybar[110]) );
  AND2_X1 U245 ( .A1(b[10]), .A2(a[0]), .ZN(y[10]) );
  OR2_X1 U245bar ( .A1(bbar[10]), .A2(abar[0]), .ZN(ybar[10]) );
  AND2_X1 U246 ( .A1(b[13]), .A2(a[6]), .ZN(y[109]) );
  OR2_X1 U246bar ( .A1(bbar[13]), .A2(abar[6]), .ZN(ybar[109]) );
  AND2_X1 U247 ( .A1(b[12]), .A2(a[6]), .ZN(y[108]) );
  OR2_X1 U247bar ( .A1(bbar[12]), .A2(abar[6]), .ZN(ybar[108]) );
  AND2_X1 U248 ( .A1(b[11]), .A2(a[6]), .ZN(y[107]) );
  OR2_X1 U248bar ( .A1(bbar[11]), .A2(abar[6]), .ZN(ybar[107]) );
  AND2_X1 U249 ( .A1(b[10]), .A2(a[6]), .ZN(y[106]) );
  OR2_X1 U249bar ( .A1(bbar[10]), .A2(abar[6]), .ZN(ybar[106]) );
  AND2_X1 U250 ( .A1(a[6]), .A2(b[9]), .ZN(y[105]) );
  OR2_X1 U250bar ( .A1(abar[6]), .A2(bbar[9]), .ZN(ybar[105]) );
  AND2_X1 U251 ( .A1(b[8]), .A2(a[6]), .ZN(y[104]) );
  OR2_X1 U251bar ( .A1(bbar[8]), .A2(abar[6]), .ZN(ybar[104]) );
  AND2_X1 U252 ( .A1(b[7]), .A2(a[6]), .ZN(y[103]) );
  OR2_X1 U252bar ( .A1(bbar[7]), .A2(abar[6]), .ZN(ybar[103]) );
  AND2_X1 U253 ( .A1(b[6]), .A2(a[6]), .ZN(y[102]) );
  OR2_X1 U253bar ( .A1(bbar[6]), .A2(abar[6]), .ZN(ybar[102]) );
  AND2_X1 U254 ( .A1(b[5]), .A2(a[6]), .ZN(y[101]) );
  OR2_X1 U254bar ( .A1(bbar[5]), .A2(abar[6]), .ZN(ybar[101]) );
  AND2_X1 U255 ( .A1(b[4]), .A2(a[6]), .ZN(y[100]) );
  OR2_X1 U255bar ( .A1(bbar[4]), .A2(abar[6]), .ZN(ybar[100]) );
  AND2_X1 U256 ( .A1(b[0]), .A2(a[0]), .ZN(y[0]) );
  OR2_X1 U256bar ( .A1(bbar[0]), .A2(abar[0]), .ZN(ybar[0]) );
endmodule

module decode_12 ( in, inbar, out, outbar );

  input wire [7:0] in;
  input wire [7:0] inbar;
//input_done

  output wire [255:0] out;
  output wire [255:0] outbar;
//output_done

  wire [15:0] level1;
  wire [31:0] level2;
  wire [15:0] level1bar;
  wire [31:0] level2bar;
//wire_done

  CD2_48 cd_l1_1 ( .a(in[1]), .abar(inbar[1]), .b(in[0]), .bbar(inbar[0]), .y(level1[3:0]), .ybar(level1bar[3:0]) );
  CD2_47 cd_l1_2 ( .a(in[3]), .abar(inbar[3]), .b(in[2]), .bbar(inbar[2]), .y(level1[7:4]), .ybar(level1bar[7:4]) );
  CD2_46 cd_l1_3 ( .a(in[5]), .abar(inbar[5]), .b(in[4]), .bbar(inbar[4]), .y(level1[11:8]), .ybar(level1bar[11:8]) );
  CD2_45 cd_l1_4 ( .a(in[7]), .abar(inbar[7]), .b(in[6]), .bbar(inbar[6]), .y(level1[15:12]), .ybar(level1bar[15:12]) );

  CD4_24 cd_l2_1 ( .a(level1[7:4]), .abar(level1bar[7:4]), .b(level1[3:0]), .bbar(level1bar[3:0]), 
        .y(level2[15:0]), .ybar(level2bar[15:0]) );
  CD4_23 cd_l2_2 ( .a(level1[15:12]), .abar(level1bar[15:12]), .b(level1[11:8]), .bbar(level1bar[11:8]), 
        .y(level2[31:16]), .ybar(level2bar[31:16]) );
  CD16_12 cd_l3 ( .a(level2[31:16]), .abar(level2bar[31:16]), .b(level2[15:0]), .bbar(level2bar[15:0]), 
        .y(out), .ybar(outbar) );
endmodule

module encode_12 ( in, inbar, out, outbar );

  input wire [255:0] in;
  input wire [255:0] inbar;
//input_done

  output wire [7:0] out;
  output wire [7:0] outbar;
//output_done

  wire in_81;
  wire in_80;
  wire in_79;
  wire in_78;
  wire in_77;
  wire in_76;
  wire in_75;
  wire in_74;
  wire in_73;
  wire in_72;
  wire in_71;
  wire in_70;
  wire in_69;
  wire in_68;
  wire in_67;
  wire in_66;
  wire in_65;
  wire in_64;
  wire in_63;
  wire in_62;
  wire in_61;
  wire in_60;
  wire in_59;
  wire in_58;
  wire in_57;
  wire in_56;
  wire in_55;
  wire in_54;
  wire in_53;
  wire in_52;
  wire in_51;
  wire in_50;
  wire in_49;
  wire in_48;
  wire in_47;
  wire in_46;
  wire in_45;
  wire in_44;
  wire in_43;
  wire in_42;
  wire in_41;
  wire in_40;
  wire in_39;
  wire in_38;
  wire in_37;
  wire in_36;
  wire in_35;
  wire in_34;
  wire in_33;
  wire in_32;
  wire in_31;
  wire in_30;
  wire in_29;
  wire in_28;
  wire in_27;
  wire in_26;
  wire in_25;
  wire in_24;
  wire in_23;
  wire in_22;
  wire in_21;
  wire in_20;
  wire in_19;
  wire in_18;
  wire in_17;
  wire in_16;
  wire in_15;
  wire in_14;
  wire in_13;
  wire in_12;
  wire in_11;
  wire in_10;
  wire in_9;
  wire in_8;
  wire in_7;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_3;
  wire in_2;
  wire in_1;
  wire in_0;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire in_81bar;
  wire in_80bar;
  wire in_79bar;
  wire in_78bar;
  wire in_77bar;
  wire in_76bar;
  wire in_75bar;
  wire in_74bar;
  wire in_73bar;
  wire in_72bar;
  wire in_71bar;
  wire in_70bar;
  wire in_69bar;
  wire in_68bar;
  wire in_67bar;
  wire in_66bar;
  wire in_65bar;
  wire in_64bar;
  wire in_63bar;
  wire in_62bar;
  wire in_61bar;
  wire in_60bar;
  wire in_59bar;
  wire in_58bar;
  wire in_57bar;
  wire in_56bar;
  wire in_55bar;
  wire in_54bar;
  wire in_53bar;
  wire in_52bar;
  wire in_51bar;
  wire in_50bar;
  wire in_49bar;
  wire in_48bar;
  wire in_47bar;
  wire in_46bar;
  wire in_45bar;
  wire in_44bar;
  wire in_43bar;
  wire in_42bar;
  wire in_41bar;
  wire in_40bar;
  wire in_39bar;
  wire in_38bar;
  wire in_37bar;
  wire in_36bar;
  wire in_35bar;
  wire in_34bar;
  wire in_33bar;
  wire in_32bar;
  wire in_31bar;
  wire in_30bar;
  wire in_29bar;
  wire in_28bar;
  wire in_27bar;
  wire in_26bar;
  wire in_25bar;
  wire in_24bar;
  wire in_23bar;
  wire in_22bar;
  wire in_21bar;
  wire in_20bar;
  wire in_19bar;
  wire in_18bar;
  wire in_17bar;
  wire in_16bar;
  wire in_15bar;
  wire in_14bar;
  wire in_13bar;
  wire in_12bar;
  wire in_11bar;
  wire in_10bar;
  wire in_9bar;
  wire in_8bar;
  wire in_7bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_3bar;
  wire in_2bar;
  wire in_1bar;
  wire in_0bar;
  wire n487bar;
  wire n488bar;
  wire n489bar;
  wire n490bar;
  wire n491bar;
  wire n492bar;
  wire n493bar;
  wire n494bar;
  wire n495bar;
  wire n496bar;
  wire n497bar;
  wire n498bar;
  wire n499bar;
  wire n500bar;
  wire n501bar;
  wire n502bar;
  wire n503bar;
  wire n504bar;
  wire n505bar;
  wire n506bar;
  wire n507bar;
  wire n508bar;
  wire n509bar;
  wire n510bar;
  wire n511bar;
  wire n512bar;
  wire n513bar;
  wire n514bar;
  wire n515bar;
  wire n516bar;
  wire n517bar;
  wire n518bar;
  wire n519bar;
  wire n520bar;
  wire n521bar;
  wire n522bar;
  wire n523bar;
  wire n524bar;
  wire n525bar;
  wire n526bar;
  wire n527bar;
  wire n528bar;
  wire n529bar;
  wire n530bar;
  wire n531bar;
  wire n532bar;
  wire n533bar;
  wire n534bar;
  wire n535bar;
  wire n536bar;
  wire n537bar;
  wire n538bar;
  wire n539bar;
  wire n540bar;
  wire n541bar;
  wire n542bar;
  wire n543bar;
  wire n544bar;
  wire n545bar;
  wire n546bar;
  wire n547bar;
  wire n548bar;
  wire n549bar;
  wire n550bar;
  wire n551bar;
  wire n552bar;
  wire n553bar;
  wire n554bar;
  wire n555bar;
  wire n556bar;
  wire n557bar;
  wire n558bar;
  wire n559bar;
  wire n560bar;
  wire n561bar;
  wire n562bar;
  wire n563bar;
  wire n564bar;
  wire n565bar;
  wire n566bar;
  wire n567bar;
  wire n568bar;
  wire n569bar;
  wire n570bar;
  wire n571bar;
  wire n572bar;
  wire n573bar;
  wire n574bar;
  wire n575bar;
  wire n576bar;
  wire n577bar;
  wire n578bar;
  wire n579bar;
  wire n580bar;
  wire n581bar;
  wire n582bar;
  wire n583bar;
  wire n584bar;
  wire n585bar;
  wire n586bar;
  wire n587bar;
  wire n588bar;
  wire n589bar;
  wire n590bar;
  wire n591bar;
  wire n592bar;
  wire n593bar;
  wire n594bar;
  wire n595bar;
  wire n596bar;
  wire n597bar;
  wire n598bar;
  wire n599bar;
  wire n600bar;
  wire n601bar;
  wire n602bar;
  wire n603bar;
  wire n604bar;
  wire n605bar;
  wire n606bar;
  wire n607bar;
  wire n608bar;
  wire n609bar;
  wire n610bar;
  wire n611bar;
  wire n612bar;
  wire n613bar;
  wire n614bar;
  wire n615bar;
  wire n616bar;
  wire n617bar;
  wire n618bar;
  wire n619bar;
  wire n620bar;
  wire n621bar;
  wire n622bar;
  wire n623bar;
  wire n624bar;
  wire n625bar;
  wire n626bar;
  wire n627bar;
  wire n628bar;
  wire n629bar;
  wire n630bar;
  wire n631bar;
  wire n632bar;
  wire n633bar;
  wire n634bar;
  wire n635bar;
  wire n636bar;
  wire n637bar;
  wire n638bar;
  wire n639bar;
  wire n640bar;
  wire n641bar;
  wire n642bar;
  wire n643bar;
  wire n644bar;
  wire n645bar;
  wire n646bar;
  wire n647bar;
  wire n648bar;
  wire n649bar;
  wire n650bar;
  wire n651bar;
  wire n652bar;
  wire n653bar;
  wire n654bar;
  wire n655bar;
  wire n656bar;
  wire n657bar;
  wire n658bar;
  wire n659bar;
  wire n660bar;
  wire n661bar;
  wire n662bar;
  wire n663bar;
  wire n664bar;
  wire n665bar;
  wire n666bar;
  wire n667bar;
  wire n668bar;
  wire n669bar;
  wire n670bar;
  wire n671bar;
  wire n672bar;
  wire n673bar;
  wire n674bar;
  wire n675bar;
  wire n676bar;
  wire n677bar;
  wire n678bar;
  wire n679bar;
  wire n680bar;
  wire n681bar;
  wire n682bar;
  wire n683bar;
  wire n684bar;
  wire n685bar;
  wire n686bar;
  wire n687bar;
  wire n688bar;
  wire n689bar;
  wire n690bar;
  wire n691bar;
  wire n692bar;
  wire n693bar;
  wire n694bar;
  wire n695bar;
  wire n696bar;
  wire n697bar;
  wire n698bar;
  wire n699bar;
  wire n700bar;
  wire n701bar;
  wire n702bar;
  wire n703bar;
  wire n704bar;
  wire n705bar;
  wire n706bar;
  wire n707bar;
  wire n708bar;
  wire n709bar;
  wire n710bar;
  wire n711bar;
  wire n712bar;
  wire n713bar;
  wire n714bar;
  wire n715bar;
  wire n716bar;
  wire n717bar;
  wire n718bar;
  wire n719bar;
  wire n720bar;
  wire n721bar;
  wire n722bar;
  wire n723bar;
  wire n724bar;
  wire n725bar;
  wire n726bar;
  wire n727bar;
  wire n728bar;
  wire n729bar;
  wire n730bar;
  wire n731bar;
  wire n732bar;
  wire n733bar;
  wire n734bar;
  wire n735bar;
  wire n736bar;
  wire n737bar;
  wire n738bar;
  wire n739bar;
  wire n740bar;
  wire n741bar;
  wire n742bar;
  wire n743bar;
  wire n744bar;
  wire n745bar;
  wire n746bar;
  wire n747bar;
  wire n748bar;
  wire n749bar;
  wire n750bar;
  wire n751bar;
  wire n752bar;
  wire n753bar;
  wire n754bar;
  wire n755bar;
  wire n756bar;
  wire n757bar;
  wire n758bar;
  wire n759bar;
  wire n760bar;
  wire n761bar;
  wire n762bar;
  wire n763bar;
  wire n764bar;
  wire n765bar;
  wire n766bar;
  wire n767bar;
  wire n768bar;
  wire n769bar;
  wire n770bar;
  wire n771bar;
  wire n772bar;
  wire n773bar;
  wire n774bar;
  wire n775bar;
  wire n776bar;
  wire n777bar;
  wire n778bar;
  wire n779bar;
  wire n780bar;
  wire n781bar;
  wire n782bar;
  wire n783bar;
  wire n784bar;
  wire n785bar;
  wire n786bar;
  wire n787bar;
  wire n788bar;
  wire n789bar;
  wire n790bar;
  wire n791bar;
  wire n792bar;
  wire n793bar;
  wire n794bar;
  wire n795bar;
  wire n796bar;
  wire n797bar;
  wire n798bar;
  wire n799bar;
  wire n800bar;
  wire n801bar;
  wire n802bar;
  wire n803bar;
  wire n804bar;
  wire n805bar;
  wire n806bar;
  wire n807bar;
  wire n808bar;
  wire n809bar;
  wire n810bar;
  wire n811bar;
  wire n812bar;
  wire n813bar;
  wire n814bar;
  wire n815bar;
  wire n816bar;
  wire n817bar;
  wire n818bar;
  wire n819bar;
  wire n820bar;
  wire n821bar;
  wire n822bar;
  wire n823bar;
  wire n824bar;
  wire n825bar;
  wire n826bar;
  wire n827bar;
  wire n828bar;
  wire n829bar;
  wire n830bar;
  wire n831bar;
  wire n832bar;
  wire n833bar;
  wire n834bar;
  wire n835bar;
  wire n836bar;
  wire n837bar;
  wire n838bar;
  wire n839bar;
  wire n840bar;
  wire n841bar;
  wire n842bar;
  wire n843bar;
  wire n844bar;
  wire n845bar;
  wire n846bar;
  wire n847bar;
  wire n848bar;
  wire n849bar;
  wire n850bar;
  wire n851bar;
  wire n852bar;
  wire n853bar;
  wire n854bar;
  wire n855bar;
  wire n856bar;
  wire n857bar;
  wire n858bar;
  wire n859bar;
  wire n860bar;
  wire n861bar;
  wire n862bar;
  wire n863bar;
  wire n864bar;
  wire n865bar;
  wire n866bar;
  wire n867bar;
  wire n868bar;
  wire n869bar;
  wire n870bar;
  wire n871bar;
  wire n872bar;
  wire n873bar;
  wire n874bar;
  wire n875bar;
  wire n876bar;
  wire n877bar;
  wire n878bar;
  wire n879bar;
  wire n880bar;
  wire n881bar;
  wire n882bar;
  wire n883bar;
  wire n884bar;
  wire n885bar;
  wire n886bar;
  wire n887bar;
  wire n888bar;
  wire n889bar;
  wire n890bar;
  wire n891bar;
  wire n892bar;
  wire n893bar;
  wire n894bar;
  wire n895bar;
  wire n896bar;
  wire n897bar;
  wire n898bar;
  wire n899bar;
  wire n900bar;
  wire n901bar;
  wire n902bar;
  wire n903bar;
  wire n904bar;
  wire n905bar;
  wire n906bar;
  wire n907bar;
  wire n908bar;
  wire n909bar;
  wire n910bar;
  wire n911bar;
  wire n912bar;
  wire n913bar;
  wire n914bar;
  wire n915bar;
  wire n916bar;
  wire n917bar;
  wire n918bar;
  wire n919bar;
  wire n920bar;
  wire n921bar;
  wire n922bar;
  wire n923bar;
  wire n924bar;
  wire n925bar;
  wire n926bar;
  wire n927bar;
  wire n928bar;
  wire n929bar;
  wire n930bar;
  wire n931bar;
  wire n932bar;
  wire n933bar;
  wire n934bar;
  wire n935bar;
  wire n936bar;
  wire n937bar;
  wire n938bar;
  wire n939bar;
  wire n940bar;
  wire n941bar;
  wire n942bar;
  wire n943bar;
  wire n944bar;
  wire n945bar;
  wire n946bar;
  wire n947bar;
  wire n948bar;
  wire n949bar;
  wire n950bar;
  wire n951bar;
  wire n952bar;
  wire n953bar;
  wire n954bar;
  wire n955bar;
  wire n956bar;
  wire n957bar;
  wire n958bar;
  wire n959bar;
  wire n960bar;
  wire n961bar;
  wire n962bar;
  wire n963bar;
  wire n964bar;
  wire n965bar;
  wire n966bar;
  wire n967bar;
  wire n968bar;
  wire n969bar;
  wire n970bar;
  wire n971bar;
  wire n972bar;
//wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];
  assign in_81bar = inbar[81];
  assign in_80bar = inbar[80];
  assign in_79bar = inbar[79];
  assign in_78bar = inbar[78];
  assign in_77bar = inbar[77];
  assign in_76bar = inbar[76];
  assign in_75bar = inbar[75];
  assign in_74bar = inbar[74];
  assign in_73bar = inbar[73];
  assign in_72bar = inbar[72];
  assign in_71bar = inbar[71];
  assign in_70bar = inbar[70];
  assign in_69bar = inbar[69];
  assign in_68bar = inbar[68];
  assign in_67bar = inbar[67];
  assign in_66bar = inbar[66];
  assign in_65bar = inbar[65];
  assign in_64bar = inbar[64];
  assign in_63bar = inbar[63];
  assign in_62bar = inbar[62];
  assign in_61bar = inbar[61];
  assign in_60bar = inbar[60];
  assign in_59bar = inbar[59];
  assign in_58bar = inbar[58];
  assign in_57bar = inbar[57];
  assign in_56bar = inbar[56];
  assign in_55bar = inbar[55];
  assign in_54bar = inbar[54];
  assign in_53bar = inbar[53];
  assign in_52bar = inbar[52];
  assign in_51bar = inbar[51];
  assign in_50bar = inbar[50];
  assign in_49bar = inbar[49];
  assign in_48bar = inbar[48];
  assign in_47bar = inbar[47];
  assign in_46bar = inbar[46];
  assign in_45bar = inbar[45];
  assign in_44bar = inbar[44];
  assign in_43bar = inbar[43];
  assign in_42bar = inbar[42];
  assign in_41bar = inbar[41];
  assign in_40bar = inbar[40];
  assign in_39bar = inbar[39];
  assign in_38bar = inbar[38];
  assign in_37bar = inbar[37];
  assign in_36bar = inbar[36];
  assign in_35bar = inbar[35];
  assign in_34bar = inbar[34];
  assign in_33bar = inbar[33];
  assign in_32bar = inbar[32];
  assign in_31bar = inbar[31];
  assign in_30bar = inbar[30];
  assign in_29bar = inbar[29];
  assign in_28bar = inbar[28];
  assign in_27bar = inbar[27];
  assign in_26bar = inbar[26];
  assign in_25bar = inbar[25];
  assign in_24bar = inbar[24];
  assign in_23bar = inbar[23];
  assign in_22bar = inbar[22];
  assign in_21bar = inbar[21];
  assign in_20bar = inbar[20];
  assign in_19bar = inbar[19];
  assign in_18bar = inbar[18];
  assign in_17bar = inbar[17];
  assign in_16bar = inbar[16];
  assign in_15bar = inbar[15];
  assign in_14bar = inbar[14];
  assign in_13bar = inbar[13];
  assign in_12bar = inbar[12];
  assign in_11bar = inbar[11];
  assign in_10bar = inbar[10];
  assign in_9bar = inbar[9];
  assign in_8bar = inbar[8];
  assign in_7bar = inbar[7];
  assign in_6bar = inbar[6];
  assign in_5bar = inbar[5];
  assign in_4bar = inbar[4];
  assign in_3bar = inbar[3];
  assign in_2bar = inbar[2];
  assign in_1bar = inbar[1];
  assign in_0bar = inbar[0];
//assign_done

  OR2_X1 U1 ( .A1(n972), .A2(n971), .ZN(out[7]) );
  AND2_X1 U1bar ( .A1(n972bar), .A2(n971bar), .ZN(outbar[7]) );
  OR2_X1 U2 ( .A1(n970), .A2(n969), .ZN(n971) );
  AND2_X1 U2bar ( .A1(n970bar), .A2(n969bar), .ZN(n971bar) );
  OR2_X1 U3 ( .A1(n968), .A2(n967), .ZN(n969) );
  AND2_X1 U3bar ( .A1(n968bar), .A2(n967bar), .ZN(n969bar) );
  OR2_X1 U4 ( .A1(n966), .A2(n965), .ZN(n967) );
  AND2_X1 U4bar ( .A1(n966bar), .A2(n965bar), .ZN(n967bar) );
  OR2_X1 U5 ( .A1(n964), .A2(n963), .ZN(n968) );
  AND2_X1 U5bar ( .A1(n964bar), .A2(n963bar), .ZN(n968bar) );
  OR2_X1 U6 ( .A1(in[116]), .A2(n962), .ZN(n963) );
  AND2_X1 U6bar ( .A1(inbar[116]), .A2(n962bar), .ZN(n963bar) );
  OR2_X1 U7 ( .A1(n961), .A2(n960), .ZN(n970) );
  AND2_X1 U7bar ( .A1(n961bar), .A2(n960bar), .ZN(n970bar) );
  OR2_X1 U8 ( .A1(in[150]), .A2(in[127]), .ZN(n960) );
  AND2_X1 U8bar ( .A1(inbar[150]), .A2(inbar[127]), .ZN(n960bar) );
  OR2_X1 U9 ( .A1(in[160]), .A2(n959), .ZN(n961) );
  AND2_X1 U9bar ( .A1(inbar[160]), .A2(n959bar), .ZN(n961bar) );
  OR2_X1 U10 ( .A1(in[252]), .A2(in[168]), .ZN(n959) );
  AND2_X1 U10bar ( .A1(inbar[252]), .A2(inbar[168]), .ZN(n959bar) );
  OR2_X1 U11 ( .A1(n958), .A2(n957), .ZN(n972) );
  AND2_X1 U11bar ( .A1(n958bar), .A2(n957bar), .ZN(n972bar) );
  OR2_X1 U12 ( .A1(n956), .A2(n955), .ZN(n957) );
  AND2_X1 U12bar ( .A1(n956bar), .A2(n955bar), .ZN(n957bar) );
  OR2_X1 U13 ( .A1(in_17), .A2(in[96]), .ZN(n955) );
  AND2_X1 U13bar ( .A1(in_17bar), .A2(inbar[96]), .ZN(n955bar) );
  OR2_X1 U14 ( .A1(in_23), .A2(n954), .ZN(n956) );
  AND2_X1 U14bar ( .A1(in_23bar), .A2(n954bar), .ZN(n956bar) );
  OR2_X1 U15 ( .A1(in_31), .A2(in_26), .ZN(n954) );
  AND2_X1 U15bar ( .A1(in_31bar), .A2(in_26bar), .ZN(n954bar) );
  OR2_X1 U16 ( .A1(n953), .A2(n952), .ZN(n958) );
  AND2_X1 U16bar ( .A1(n953bar), .A2(n952bar), .ZN(n958bar) );
  OR2_X1 U17 ( .A1(in_58), .A2(in_4), .ZN(n952) );
  AND2_X1 U17bar ( .A1(in_58bar), .A2(in_4bar), .ZN(n952bar) );
  OR2_X1 U18 ( .A1(in_59), .A2(n951), .ZN(n953) );
  AND2_X1 U18bar ( .A1(in_59bar), .A2(n951bar), .ZN(n953bar) );
  OR2_X1 U19 ( .A1(in_71), .A2(in_62), .ZN(n951) );
  AND2_X1 U19bar ( .A1(in_71bar), .A2(in_62bar), .ZN(n951bar) );
  OR2_X1 U20 ( .A1(n950), .A2(n949), .ZN(out[6]) );
  AND2_X1 U20bar ( .A1(n950bar), .A2(n949bar), .ZN(outbar[6]) );
  OR2_X1 U21 ( .A1(n948), .A2(n947), .ZN(n949) );
  AND2_X1 U21bar ( .A1(n948bar), .A2(n947bar), .ZN(n949bar) );
  OR2_X1 U22 ( .A1(n946), .A2(n945), .ZN(n947) );
  AND2_X1 U22bar ( .A1(n946bar), .A2(n945bar), .ZN(n947bar) );
  OR2_X1 U23 ( .A1(n944), .A2(n943), .ZN(n945) );
  AND2_X1 U23bar ( .A1(n944bar), .A2(n943bar), .ZN(n945bar) );
  OR2_X1 U24 ( .A1(n942), .A2(n941), .ZN(n946) );
  AND2_X1 U24bar ( .A1(n942bar), .A2(n941bar), .ZN(n946bar) );
  OR2_X1 U25 ( .A1(in[101]), .A2(n940), .ZN(n941) );
  AND2_X1 U25bar ( .A1(inbar[101]), .A2(n940bar), .ZN(n941bar) );
  OR2_X1 U26 ( .A1(n939), .A2(n938), .ZN(n948) );
  AND2_X1 U26bar ( .A1(n939bar), .A2(n938bar), .ZN(n948bar) );
  OR2_X1 U27 ( .A1(in[114]), .A2(in[104]), .ZN(n938) );
  AND2_X1 U27bar ( .A1(inbar[114]), .A2(inbar[104]), .ZN(n938bar) );
  OR2_X1 U28 ( .A1(in[128]), .A2(n937), .ZN(n939) );
  AND2_X1 U28bar ( .A1(inbar[128]), .A2(n937bar), .ZN(n939bar) );
  OR2_X1 U29 ( .A1(in[136]), .A2(in[134]), .ZN(n937) );
  AND2_X1 U29bar ( .A1(inbar[136]), .A2(inbar[134]), .ZN(n937bar) );
  OR2_X1 U30 ( .A1(n936), .A2(n935), .ZN(n950) );
  AND2_X1 U30bar ( .A1(n936bar), .A2(n935bar), .ZN(n950bar) );
  OR2_X1 U31 ( .A1(n934), .A2(n933), .ZN(n935) );
  AND2_X1 U31bar ( .A1(n934bar), .A2(n933bar), .ZN(n935bar) );
  OR2_X1 U32 ( .A1(in[177]), .A2(in[164]), .ZN(n933) );
  AND2_X1 U32bar ( .A1(inbar[177]), .A2(inbar[164]), .ZN(n933bar) );
  OR2_X1 U33 ( .A1(in[212]), .A2(n932), .ZN(n934) );
  AND2_X1 U33bar ( .A1(inbar[212]), .A2(n932bar), .ZN(n934bar) );
  OR2_X1 U34 ( .A1(in[248]), .A2(in[221]), .ZN(n932) );
  AND2_X1 U34bar ( .A1(inbar[248]), .A2(inbar[221]), .ZN(n932bar) );
  OR2_X1 U35 ( .A1(n931), .A2(n930), .ZN(n936) );
  AND2_X1 U35bar ( .A1(n931bar), .A2(n930bar), .ZN(n936bar) );
  OR2_X1 U36 ( .A1(in_18), .A2(in[93]), .ZN(n930) );
  AND2_X1 U36bar ( .A1(in_18bar), .A2(inbar[93]), .ZN(n930bar) );
  OR2_X1 U37 ( .A1(in_31), .A2(n929), .ZN(n931) );
  AND2_X1 U37bar ( .A1(in_31bar), .A2(n929bar), .ZN(n931bar) );
  OR2_X1 U38 ( .A1(in_7), .A2(in_39), .ZN(n929) );
  AND2_X1 U38bar ( .A1(in_7bar), .A2(in_39bar), .ZN(n929bar) );
  OR2_X1 U39 ( .A1(n928), .A2(n927), .ZN(out[5]) );
  AND2_X1 U39bar ( .A1(n928bar), .A2(n927bar), .ZN(outbar[5]) );
  OR2_X1 U40 ( .A1(n926), .A2(n925), .ZN(n927) );
  AND2_X1 U40bar ( .A1(n926bar), .A2(n925bar), .ZN(n927bar) );
  OR2_X1 U41 ( .A1(n924), .A2(n923), .ZN(n925) );
  AND2_X1 U41bar ( .A1(n924bar), .A2(n923bar), .ZN(n925bar) );
  OR2_X1 U42 ( .A1(n922), .A2(n921), .ZN(n923) );
  AND2_X1 U42bar ( .A1(n922bar), .A2(n921bar), .ZN(n923bar) );
  OR2_X1 U43 ( .A1(n940), .A2(n920), .ZN(n924) );
  AND2_X1 U43bar ( .A1(n940bar), .A2(n920bar), .ZN(n924bar) );
  OR2_X1 U44 ( .A1(in[111]), .A2(n919), .ZN(n920) );
  AND2_X1 U44bar ( .A1(inbar[111]), .A2(n919bar), .ZN(n920bar) );
  OR2_X1 U45 ( .A1(n918), .A2(n917), .ZN(n940) );
  AND2_X1 U45bar ( .A1(n918bar), .A2(n917bar), .ZN(n940bar) );
  OR2_X1 U46 ( .A1(n916), .A2(n915), .ZN(n917) );
  AND2_X1 U46bar ( .A1(n916bar), .A2(n915bar), .ZN(n917bar) );
  OR2_X1 U47 ( .A1(n914), .A2(n913), .ZN(n915) );
  AND2_X1 U47bar ( .A1(n914bar), .A2(n913bar), .ZN(n915bar) );
  OR2_X1 U48 ( .A1(in[140]), .A2(in[131]), .ZN(n913) );
  AND2_X1 U48bar ( .A1(inbar[140]), .A2(inbar[131]), .ZN(n913bar) );
  OR2_X1 U49 ( .A1(in[160]), .A2(in[144]), .ZN(n914) );
  AND2_X1 U49bar ( .A1(inbar[160]), .A2(inbar[144]), .ZN(n914bar) );
  OR2_X1 U50 ( .A1(n912), .A2(n911), .ZN(n916) );
  AND2_X1 U50bar ( .A1(n912bar), .A2(n911bar), .ZN(n916bar) );
  OR2_X1 U51 ( .A1(in[179]), .A2(in[174]), .ZN(n911) );
  AND2_X1 U51bar ( .A1(inbar[179]), .A2(inbar[174]), .ZN(n911bar) );
  OR2_X1 U52 ( .A1(in[188]), .A2(in[184]), .ZN(n912) );
  AND2_X1 U52bar ( .A1(inbar[188]), .A2(inbar[184]), .ZN(n912bar) );
  OR2_X1 U53 ( .A1(n910), .A2(n909), .ZN(n918) );
  AND2_X1 U53bar ( .A1(n910bar), .A2(n909bar), .ZN(n918bar) );
  OR2_X1 U54 ( .A1(n908), .A2(n907), .ZN(n909) );
  AND2_X1 U54bar ( .A1(n908bar), .A2(n907bar), .ZN(n909bar) );
  OR2_X1 U55 ( .A1(in[216]), .A2(in[200]), .ZN(n907) );
  AND2_X1 U55bar ( .A1(inbar[216]), .A2(inbar[200]), .ZN(n907bar) );
  OR2_X1 U56 ( .A1(in[228]), .A2(in[224]), .ZN(n908) );
  AND2_X1 U56bar ( .A1(inbar[228]), .A2(inbar[224]), .ZN(n908bar) );
  OR2_X1 U57 ( .A1(n906), .A2(n905), .ZN(n910) );
  AND2_X1 U57bar ( .A1(n906bar), .A2(n905bar), .ZN(n910bar) );
  OR2_X1 U58 ( .A1(in[247]), .A2(in[235]), .ZN(n905) );
  AND2_X1 U58bar ( .A1(inbar[247]), .A2(inbar[235]), .ZN(n905bar) );
  OR2_X1 U59 ( .A1(in_42), .A2(in[83]), .ZN(n906) );
  AND2_X1 U59bar ( .A1(in_42bar), .A2(inbar[83]), .ZN(n906bar) );
  OR2_X1 U60 ( .A1(n904), .A2(n903), .ZN(n926) );
  AND2_X1 U60bar ( .A1(n904bar), .A2(n903bar), .ZN(n926bar) );
  OR2_X1 U61 ( .A1(in[166]), .A2(in[123]), .ZN(n903) );
  AND2_X1 U61bar ( .A1(inbar[166]), .A2(inbar[123]), .ZN(n903bar) );
  OR2_X1 U62 ( .A1(in[170]), .A2(n902), .ZN(n904) );
  AND2_X1 U62bar ( .A1(inbar[170]), .A2(n902bar), .ZN(n904bar) );
  OR2_X1 U63 ( .A1(in[194]), .A2(in[183]), .ZN(n902) );
  AND2_X1 U63bar ( .A1(inbar[194]), .A2(inbar[183]), .ZN(n902bar) );
  OR2_X1 U64 ( .A1(n901), .A2(n900), .ZN(n928) );
  AND2_X1 U64bar ( .A1(n901bar), .A2(n900bar), .ZN(n928bar) );
  OR2_X1 U65 ( .A1(n899), .A2(n898), .ZN(n900) );
  AND2_X1 U65bar ( .A1(n899bar), .A2(n898bar), .ZN(n900bar) );
  OR2_X1 U66 ( .A1(in[241]), .A2(in[238]), .ZN(n898) );
  AND2_X1 U66bar ( .A1(inbar[241]), .A2(inbar[238]), .ZN(n898bar) );
  OR2_X1 U67 ( .A1(in[250]), .A2(n897), .ZN(n899) );
  AND2_X1 U67bar ( .A1(inbar[250]), .A2(n897bar), .ZN(n899bar) );
  OR2_X1 U68 ( .A1(in_24), .A2(in[84]), .ZN(n897) );
  AND2_X1 U68bar ( .A1(in_24bar), .A2(inbar[84]), .ZN(n897bar) );
  OR2_X1 U69 ( .A1(n896), .A2(n895), .ZN(n901) );
  AND2_X1 U69bar ( .A1(n896bar), .A2(n895bar), .ZN(n901bar) );
  OR2_X1 U70 ( .A1(in_41), .A2(in_29), .ZN(n895) );
  AND2_X1 U70bar ( .A1(in_41bar), .A2(in_29bar), .ZN(n895bar) );
  OR2_X1 U71 ( .A1(in_66), .A2(n894), .ZN(n896) );
  AND2_X1 U71bar ( .A1(in_66bar), .A2(n894bar), .ZN(n896bar) );
  OR2_X1 U72 ( .A1(in_76), .A2(in_71), .ZN(n894) );
  AND2_X1 U72bar ( .A1(in_76bar), .A2(in_71bar), .ZN(n894bar) );
  OR2_X1 U73 ( .A1(n893), .A2(n892), .ZN(out[4]) );
  AND2_X1 U73bar ( .A1(n893bar), .A2(n892bar), .ZN(outbar[4]) );
  OR2_X1 U74 ( .A1(n891), .A2(n890), .ZN(n892) );
  AND2_X1 U74bar ( .A1(n891bar), .A2(n890bar), .ZN(n892bar) );
  OR2_X1 U75 ( .A1(n889), .A2(n888), .ZN(n890) );
  AND2_X1 U75bar ( .A1(n889bar), .A2(n888bar), .ZN(n890bar) );
  OR2_X1 U76 ( .A1(n922), .A2(n887), .ZN(n888) );
  AND2_X1 U76bar ( .A1(n922bar), .A2(n887bar), .ZN(n888bar) );
  OR2_X1 U77 ( .A1(n886), .A2(n885), .ZN(n922) );
  AND2_X1 U77bar ( .A1(n886bar), .A2(n885bar), .ZN(n922bar) );
  OR2_X1 U78 ( .A1(n884), .A2(n883), .ZN(n885) );
  AND2_X1 U78bar ( .A1(n884bar), .A2(n883bar), .ZN(n885bar) );
  OR2_X1 U79 ( .A1(n882), .A2(n881), .ZN(n883) );
  AND2_X1 U79bar ( .A1(n882bar), .A2(n881bar), .ZN(n883bar) );
  OR2_X1 U80 ( .A1(in[118]), .A2(in[109]), .ZN(n881) );
  AND2_X1 U80bar ( .A1(inbar[118]), .A2(inbar[109]), .ZN(n881bar) );
  OR2_X1 U81 ( .A1(in[139]), .A2(in[120]), .ZN(n882) );
  AND2_X1 U81bar ( .A1(inbar[139]), .A2(inbar[120]), .ZN(n882bar) );
  OR2_X1 U82 ( .A1(n880), .A2(n879), .ZN(n884) );
  AND2_X1 U82bar ( .A1(n880bar), .A2(n879bar), .ZN(n884bar) );
  OR2_X1 U83 ( .A1(in[198]), .A2(in[154]), .ZN(n879) );
  AND2_X1 U83bar ( .A1(inbar[198]), .A2(inbar[154]), .ZN(n879bar) );
  OR2_X1 U84 ( .A1(in[210]), .A2(in[205]), .ZN(n880) );
  AND2_X1 U84bar ( .A1(inbar[210]), .A2(inbar[205]), .ZN(n880bar) );
  OR2_X1 U85 ( .A1(n878), .A2(n877), .ZN(n886) );
  AND2_X1 U85bar ( .A1(n878bar), .A2(n877bar), .ZN(n886bar) );
  OR2_X1 U86 ( .A1(n876), .A2(n875), .ZN(n877) );
  AND2_X1 U86bar ( .A1(n876bar), .A2(n875bar), .ZN(n877bar) );
  OR2_X1 U87 ( .A1(in[219]), .A2(in[217]), .ZN(n875) );
  AND2_X1 U87bar ( .A1(inbar[219]), .A2(inbar[217]), .ZN(n875bar) );
  OR2_X1 U88 ( .A1(in[86]), .A2(in[252]), .ZN(n876) );
  AND2_X1 U88bar ( .A1(inbar[86]), .A2(inbar[252]), .ZN(n876bar) );
  OR2_X1 U89 ( .A1(n874), .A2(n873), .ZN(n878) );
  AND2_X1 U89bar ( .A1(n874bar), .A2(n873bar), .ZN(n878bar) );
  OR2_X1 U90 ( .A1(in_40), .A2(in[91]), .ZN(n873) );
  AND2_X1 U90bar ( .A1(in_40bar), .A2(inbar[91]), .ZN(n873bar) );
  OR2_X1 U91 ( .A1(in_8), .A2(in_46), .ZN(n874) );
  AND2_X1 U91bar ( .A1(in_8bar), .A2(in_46bar), .ZN(n874bar) );
  OR2_X1 U92 ( .A1(n872), .A2(n871), .ZN(n889) );
  AND2_X1 U92bar ( .A1(n872bar), .A2(n871bar), .ZN(n889bar) );
  OR2_X1 U93 ( .A1(in[117]), .A2(n943), .ZN(n871) );
  AND2_X1 U93bar ( .A1(inbar[117]), .A2(n943bar), .ZN(n871bar) );
  OR2_X1 U94 ( .A1(n870), .A2(n869), .ZN(n943) );
  AND2_X1 U94bar ( .A1(n870bar), .A2(n869bar), .ZN(n943bar) );
  OR2_X1 U95 ( .A1(n868), .A2(n867), .ZN(n869) );
  AND2_X1 U95bar ( .A1(n868bar), .A2(n867bar), .ZN(n869bar) );
  OR2_X1 U96 ( .A1(n866), .A2(n865), .ZN(n867) );
  AND2_X1 U96bar ( .A1(n866bar), .A2(n865bar), .ZN(n867bar) );
  OR2_X1 U97 ( .A1(n864), .A2(n863), .ZN(n865) );
  AND2_X1 U97bar ( .A1(n864bar), .A2(n863bar), .ZN(n865bar) );
  OR2_X1 U98 ( .A1(in[108]), .A2(n919), .ZN(n866) );
  AND2_X1 U98bar ( .A1(inbar[108]), .A2(n919bar), .ZN(n866bar) );
  OR2_X1 U99 ( .A1(n862), .A2(n861), .ZN(n919) );
  AND2_X1 U99bar ( .A1(n862bar), .A2(n861bar), .ZN(n919bar) );
  OR2_X1 U100 ( .A1(n860), .A2(n859), .ZN(n861) );
  AND2_X1 U100bar ( .A1(n860bar), .A2(n859bar), .ZN(n861bar) );
  OR2_X1 U101 ( .A1(n858), .A2(n857), .ZN(n859) );
  AND2_X1 U101bar ( .A1(n858bar), .A2(n857bar), .ZN(n859bar) );
  OR2_X1 U102 ( .A1(in[119]), .A2(in[105]), .ZN(n857) );
  AND2_X1 U102bar ( .A1(inbar[119]), .A2(inbar[105]), .ZN(n857bar) );
  OR2_X1 U103 ( .A1(in[186]), .A2(in[175]), .ZN(n858) );
  AND2_X1 U103bar ( .A1(inbar[186]), .A2(inbar[175]), .ZN(n858bar) );
  OR2_X1 U104 ( .A1(n856), .A2(n855), .ZN(n860) );
  AND2_X1 U104bar ( .A1(n856bar), .A2(n855bar), .ZN(n860bar) );
  OR2_X1 U105 ( .A1(in[202]), .A2(in[193]), .ZN(n855) );
  AND2_X1 U105bar ( .A1(inbar[202]), .A2(inbar[193]), .ZN(n855bar) );
  OR2_X1 U106 ( .A1(in[225]), .A2(in[208]), .ZN(n856) );
  AND2_X1 U106bar ( .A1(inbar[225]), .A2(inbar[208]), .ZN(n856bar) );
  OR2_X1 U107 ( .A1(n854), .A2(n853), .ZN(n862) );
  AND2_X1 U107bar ( .A1(n854bar), .A2(n853bar), .ZN(n862bar) );
  OR2_X1 U108 ( .A1(n852), .A2(n851), .ZN(n853) );
  AND2_X1 U108bar ( .A1(n852bar), .A2(n851bar), .ZN(n853bar) );
  OR2_X1 U109 ( .A1(in_1), .A2(in[85]), .ZN(n851) );
  AND2_X1 U109bar ( .A1(in_1bar), .A2(inbar[85]), .ZN(n851bar) );
  OR2_X1 U110 ( .A1(in_23), .A2(in_19), .ZN(n852) );
  AND2_X1 U110bar ( .A1(in_23bar), .A2(in_19bar), .ZN(n852bar) );
  OR2_X1 U111 ( .A1(n850), .A2(n849), .ZN(n854) );
  AND2_X1 U111bar ( .A1(n850bar), .A2(n849bar), .ZN(n854bar) );
  OR2_X1 U112 ( .A1(in_43), .A2(in_33), .ZN(n849) );
  AND2_X1 U112bar ( .A1(in_43bar), .A2(in_33bar), .ZN(n849bar) );
  OR2_X1 U113 ( .A1(in_63), .A2(in_44), .ZN(n850) );
  AND2_X1 U113bar ( .A1(in_63bar), .A2(in_44bar), .ZN(n850bar) );
  OR2_X1 U114 ( .A1(n848), .A2(n847), .ZN(n868) );
  AND2_X1 U114bar ( .A1(n848bar), .A2(n847bar), .ZN(n868bar) );
  OR2_X1 U115 ( .A1(in[141]), .A2(in[112]), .ZN(n847) );
  AND2_X1 U115bar ( .A1(inbar[141]), .A2(inbar[112]), .ZN(n847bar) );
  OR2_X1 U116 ( .A1(in[147]), .A2(n846), .ZN(n848) );
  AND2_X1 U116bar ( .A1(inbar[147]), .A2(n846bar), .ZN(n848bar) );
  OR2_X1 U117 ( .A1(in[181]), .A2(in[167]), .ZN(n846) );
  AND2_X1 U117bar ( .A1(inbar[181]), .A2(inbar[167]), .ZN(n846bar) );
  OR2_X1 U118 ( .A1(n845), .A2(n844), .ZN(n870) );
  AND2_X1 U118bar ( .A1(n845bar), .A2(n844bar), .ZN(n870bar) );
  OR2_X1 U119 ( .A1(n843), .A2(n842), .ZN(n844) );
  AND2_X1 U119bar ( .A1(n843bar), .A2(n842bar), .ZN(n844bar) );
  OR2_X1 U120 ( .A1(in[229]), .A2(in[201]), .ZN(n842) );
  AND2_X1 U120bar ( .A1(inbar[229]), .A2(inbar[201]), .ZN(n842bar) );
  OR2_X1 U121 ( .A1(in[237]), .A2(n841), .ZN(n843) );
  AND2_X1 U121bar ( .A1(inbar[237]), .A2(n841bar), .ZN(n843bar) );
  OR2_X1 U122 ( .A1(in[94]), .A2(in[253]), .ZN(n841) );
  AND2_X1 U122bar ( .A1(inbar[94]), .A2(inbar[253]), .ZN(n841bar) );
  OR2_X1 U123 ( .A1(n840), .A2(n839), .ZN(n845) );
  AND2_X1 U123bar ( .A1(n840bar), .A2(n839bar), .ZN(n845bar) );
  OR2_X1 U124 ( .A1(in_21), .A2(in[96]), .ZN(n839) );
  AND2_X1 U124bar ( .A1(in_21bar), .A2(inbar[96]), .ZN(n839bar) );
  OR2_X1 U125 ( .A1(in_25), .A2(n838), .ZN(n840) );
  AND2_X1 U125bar ( .A1(in_25bar), .A2(n838bar), .ZN(n840bar) );
  OR2_X1 U126 ( .A1(in_81), .A2(in_45), .ZN(n838) );
  AND2_X1 U126bar ( .A1(in_81bar), .A2(in_45bar), .ZN(n838bar) );
  OR2_X1 U127 ( .A1(n837), .A2(n836), .ZN(n891) );
  AND2_X1 U127bar ( .A1(n837bar), .A2(n836bar), .ZN(n891bar) );
  OR2_X1 U128 ( .A1(in[142]), .A2(in[124]), .ZN(n836) );
  AND2_X1 U128bar ( .A1(inbar[142]), .A2(inbar[124]), .ZN(n836bar) );
  OR2_X1 U129 ( .A1(in[150]), .A2(n835), .ZN(n837) );
  AND2_X1 U129bar ( .A1(inbar[150]), .A2(n835bar), .ZN(n837bar) );
  OR2_X1 U130 ( .A1(in[172]), .A2(in[155]), .ZN(n835) );
  AND2_X1 U130bar ( .A1(inbar[172]), .A2(inbar[155]), .ZN(n835bar) );
  OR2_X1 U131 ( .A1(n834), .A2(n833), .ZN(n893) );
  AND2_X1 U131bar ( .A1(n834bar), .A2(n833bar), .ZN(n893bar) );
  OR2_X1 U132 ( .A1(n832), .A2(n831), .ZN(n833) );
  AND2_X1 U132bar ( .A1(n832bar), .A2(n831bar), .ZN(n833bar) );
  OR2_X1 U133 ( .A1(in[196]), .A2(in[173]), .ZN(n831) );
  AND2_X1 U133bar ( .A1(inbar[196]), .A2(inbar[173]), .ZN(n831bar) );
  OR2_X1 U134 ( .A1(in[222]), .A2(n830), .ZN(n832) );
  AND2_X1 U134bar ( .A1(inbar[222]), .A2(n830bar), .ZN(n832bar) );
  OR2_X1 U135 ( .A1(in[227]), .A2(in[226]), .ZN(n830) );
  AND2_X1 U135bar ( .A1(inbar[227]), .A2(inbar[226]), .ZN(n830bar) );
  OR2_X1 U136 ( .A1(n829), .A2(n828), .ZN(n834) );
  AND2_X1 U136bar ( .A1(n829bar), .A2(n828bar), .ZN(n834bar) );
  OR2_X1 U137 ( .A1(in[249]), .A2(in[231]), .ZN(n828) );
  AND2_X1 U137bar ( .A1(inbar[249]), .A2(inbar[231]), .ZN(n828bar) );
  OR2_X1 U138 ( .A1(in_28), .A2(n827), .ZN(n829) );
  AND2_X1 U138bar ( .A1(in_28bar), .A2(n827bar), .ZN(n829bar) );
  OR2_X1 U139 ( .A1(in_52), .A2(in_47), .ZN(n827) );
  AND2_X1 U139bar ( .A1(in_52bar), .A2(in_47bar), .ZN(n827bar) );
  OR2_X1 U140 ( .A1(n826), .A2(n825), .ZN(out[3]) );
  AND2_X1 U140bar ( .A1(n826bar), .A2(n825bar), .ZN(outbar[3]) );
  OR2_X1 U141 ( .A1(n824), .A2(n823), .ZN(n825) );
  AND2_X1 U141bar ( .A1(n824bar), .A2(n823bar), .ZN(n825bar) );
  OR2_X1 U142 ( .A1(n822), .A2(n821), .ZN(n823) );
  AND2_X1 U142bar ( .A1(n822bar), .A2(n821bar), .ZN(n823bar) );
  OR2_X1 U143 ( .A1(n820), .A2(n819), .ZN(n821) );
  AND2_X1 U143bar ( .A1(n820bar), .A2(n819bar), .ZN(n821bar) );
  OR2_X1 U144 ( .A1(n964), .A2(n818), .ZN(n822) );
  AND2_X1 U144bar ( .A1(n964bar), .A2(n818bar), .ZN(n822bar) );
  OR2_X1 U145 ( .A1(in[118]), .A2(n817), .ZN(n818) );
  AND2_X1 U145bar ( .A1(inbar[118]), .A2(n817bar), .ZN(n818bar) );
  OR2_X1 U146 ( .A1(n816), .A2(n815), .ZN(n964) );
  AND2_X1 U146bar ( .A1(n816bar), .A2(n815bar), .ZN(n964bar) );
  OR2_X1 U147 ( .A1(n814), .A2(n813), .ZN(n815) );
  AND2_X1 U147bar ( .A1(n814bar), .A2(n813bar), .ZN(n815bar) );
  OR2_X1 U148 ( .A1(n812), .A2(n811), .ZN(n813) );
  AND2_X1 U148bar ( .A1(n812bar), .A2(n811bar), .ZN(n813bar) );
  OR2_X1 U149 ( .A1(in[122]), .A2(in[111]), .ZN(n811) );
  AND2_X1 U149bar ( .A1(inbar[122]), .A2(inbar[111]), .ZN(n811bar) );
  OR2_X1 U150 ( .A1(in[154]), .A2(in[151]), .ZN(n812) );
  AND2_X1 U150bar ( .A1(inbar[154]), .A2(inbar[151]), .ZN(n812bar) );
  OR2_X1 U151 ( .A1(n810), .A2(n809), .ZN(n814) );
  AND2_X1 U151bar ( .A1(n810bar), .A2(n809bar), .ZN(n814bar) );
  OR2_X1 U152 ( .A1(in[187]), .A2(in[177]), .ZN(n809) );
  AND2_X1 U152bar ( .A1(inbar[187]), .A2(inbar[177]), .ZN(n809bar) );
  OR2_X1 U153 ( .A1(in[200]), .A2(in[192]), .ZN(n810) );
  AND2_X1 U153bar ( .A1(inbar[200]), .A2(inbar[192]), .ZN(n810bar) );
  OR2_X1 U154 ( .A1(n808), .A2(n807), .ZN(n816) );
  AND2_X1 U154bar ( .A1(n808bar), .A2(n807bar), .ZN(n816bar) );
  OR2_X1 U155 ( .A1(n806), .A2(n805), .ZN(n807) );
  AND2_X1 U155bar ( .A1(n806bar), .A2(n805bar), .ZN(n807bar) );
  OR2_X1 U156 ( .A1(in[225]), .A2(in[207]), .ZN(n805) );
  AND2_X1 U156bar ( .A1(inbar[225]), .A2(inbar[207]), .ZN(n805bar) );
  OR2_X1 U157 ( .A1(in[98]), .A2(in[226]), .ZN(n806) );
  AND2_X1 U157bar ( .A1(inbar[98]), .A2(inbar[226]), .ZN(n806bar) );
  OR2_X1 U158 ( .A1(n804), .A2(n803), .ZN(n808) );
  AND2_X1 U158bar ( .A1(n804bar), .A2(n803bar), .ZN(n808bar) );
  OR2_X1 U159 ( .A1(in_20), .A2(in_16), .ZN(n803) );
  AND2_X1 U159bar ( .A1(in_20bar), .A2(in_16bar), .ZN(n803bar) );
  OR2_X1 U160 ( .A1(in_55), .A2(in_45), .ZN(n804) );
  AND2_X1 U160bar ( .A1(in_55bar), .A2(in_45bar), .ZN(n804bar) );
  OR2_X1 U161 ( .A1(n802), .A2(n801), .ZN(n824) );
  AND2_X1 U161bar ( .A1(n802bar), .A2(n801bar), .ZN(n824bar) );
  OR2_X1 U162 ( .A1(in[162]), .A2(in[149]), .ZN(n801) );
  AND2_X1 U162bar ( .A1(inbar[162]), .A2(inbar[149]), .ZN(n801bar) );
  OR2_X1 U163 ( .A1(in[163]), .A2(n800), .ZN(n802) );
  AND2_X1 U163bar ( .A1(inbar[163]), .A2(n800bar), .ZN(n802bar) );
  OR2_X1 U164 ( .A1(in[191]), .A2(in[189]), .ZN(n800) );
  AND2_X1 U164bar ( .A1(inbar[191]), .A2(inbar[189]), .ZN(n800bar) );
  OR2_X1 U165 ( .A1(n799), .A2(n798), .ZN(n826) );
  AND2_X1 U165bar ( .A1(n799bar), .A2(n798bar), .ZN(n826bar) );
  OR2_X1 U166 ( .A1(n797), .A2(n796), .ZN(n798) );
  AND2_X1 U166bar ( .A1(n797bar), .A2(n796bar), .ZN(n798bar) );
  OR2_X1 U167 ( .A1(in[212]), .A2(in[193]), .ZN(n796) );
  AND2_X1 U167bar ( .A1(inbar[212]), .A2(inbar[193]), .ZN(n796bar) );
  OR2_X1 U168 ( .A1(in[238]), .A2(n795), .ZN(n797) );
  AND2_X1 U168bar ( .A1(inbar[238]), .A2(n795bar), .ZN(n797bar) );
  OR2_X1 U169 ( .A1(in[88]), .A2(in[247]), .ZN(n795) );
  AND2_X1 U169bar ( .A1(inbar[88]), .A2(inbar[247]), .ZN(n795bar) );
  OR2_X1 U170 ( .A1(n794), .A2(n793), .ZN(n799) );
  AND2_X1 U170bar ( .A1(n794bar), .A2(n793bar), .ZN(n799bar) );
  OR2_X1 U171 ( .A1(in[94]), .A2(in[92]), .ZN(n793) );
  AND2_X1 U171bar ( .A1(inbar[94]), .A2(inbar[92]), .ZN(n793bar) );
  OR2_X1 U172 ( .A1(in_52), .A2(n792), .ZN(n794) );
  AND2_X1 U172bar ( .A1(in_52bar), .A2(n792bar), .ZN(n794bar) );
  OR2_X1 U173 ( .A1(in_70), .A2(in_67), .ZN(n792) );
  AND2_X1 U173bar ( .A1(in_70bar), .A2(in_67bar), .ZN(n792bar) );
  OR2_X1 U174 ( .A1(n791), .A2(n790), .ZN(out[2]) );
  AND2_X1 U174bar ( .A1(n791bar), .A2(n790bar), .ZN(outbar[2]) );
  OR2_X1 U175 ( .A1(n789), .A2(n788), .ZN(n790) );
  AND2_X1 U175bar ( .A1(n789bar), .A2(n788bar), .ZN(n790bar) );
  OR2_X1 U176 ( .A1(n787), .A2(n786), .ZN(n788) );
  AND2_X1 U176bar ( .A1(n787bar), .A2(n786bar), .ZN(n788bar) );
  OR2_X1 U177 ( .A1(n819), .A2(n785), .ZN(n786) );
  AND2_X1 U177bar ( .A1(n819bar), .A2(n785bar), .ZN(n786bar) );
  OR2_X1 U178 ( .A1(n784), .A2(n783), .ZN(n819) );
  AND2_X1 U178bar ( .A1(n784bar), .A2(n783bar), .ZN(n819bar) );
  OR2_X1 U179 ( .A1(n782), .A2(n781), .ZN(n783) );
  AND2_X1 U179bar ( .A1(n782bar), .A2(n781bar), .ZN(n783bar) );
  OR2_X1 U180 ( .A1(n780), .A2(n779), .ZN(n781) );
  AND2_X1 U180bar ( .A1(n780bar), .A2(n779bar), .ZN(n781bar) );
  OR2_X1 U181 ( .A1(n962), .A2(n778), .ZN(n779) );
  AND2_X1 U181bar ( .A1(n962bar), .A2(n778bar), .ZN(n779bar) );
  OR2_X1 U182 ( .A1(n777), .A2(n776), .ZN(n962) );
  AND2_X1 U182bar ( .A1(n777bar), .A2(n776bar), .ZN(n962bar) );
  OR2_X1 U183 ( .A1(n775), .A2(n774), .ZN(n776) );
  AND2_X1 U183bar ( .A1(n775bar), .A2(n774bar), .ZN(n776bar) );
  OR2_X1 U184 ( .A1(n773), .A2(n772), .ZN(n774) );
  AND2_X1 U184bar ( .A1(n773bar), .A2(n772bar), .ZN(n774bar) );
  OR2_X1 U185 ( .A1(in[131]), .A2(in[120]), .ZN(n772) );
  AND2_X1 U185bar ( .A1(inbar[131]), .A2(inbar[120]), .ZN(n772bar) );
  OR2_X1 U186 ( .A1(in[153]), .A2(in[147]), .ZN(n773) );
  AND2_X1 U186bar ( .A1(inbar[153]), .A2(inbar[147]), .ZN(n773bar) );
  OR2_X1 U187 ( .A1(n771), .A2(n770), .ZN(n775) );
  AND2_X1 U187bar ( .A1(n771bar), .A2(n770bar), .ZN(n775bar) );
  OR2_X1 U188 ( .A1(in[170]), .A2(in[156]), .ZN(n770) );
  AND2_X1 U188bar ( .A1(inbar[170]), .A2(inbar[156]), .ZN(n770bar) );
  OR2_X1 U189 ( .A1(in[223]), .A2(in[190]), .ZN(n771) );
  AND2_X1 U189bar ( .A1(inbar[223]), .A2(inbar[190]), .ZN(n771bar) );
  OR2_X1 U190 ( .A1(n769), .A2(n768), .ZN(n777) );
  AND2_X1 U190bar ( .A1(n769bar), .A2(n768bar), .ZN(n777bar) );
  OR2_X1 U191 ( .A1(n767), .A2(n766), .ZN(n768) );
  AND2_X1 U191bar ( .A1(n767bar), .A2(n766bar), .ZN(n768bar) );
  OR2_X1 U192 ( .A1(in[236]), .A2(in[230]), .ZN(n766) );
  AND2_X1 U192bar ( .A1(inbar[236]), .A2(inbar[230]), .ZN(n766bar) );
  OR2_X1 U193 ( .A1(in[85]), .A2(in[240]), .ZN(n767) );
  AND2_X1 U193bar ( .A1(inbar[85]), .A2(inbar[240]), .ZN(n767bar) );
  OR2_X1 U194 ( .A1(n765), .A2(n764), .ZN(n769) );
  AND2_X1 U194bar ( .A1(n765bar), .A2(n764bar), .ZN(n769bar) );
  OR2_X1 U195 ( .A1(in_12), .A2(in[90]), .ZN(n764) );
  AND2_X1 U195bar ( .A1(in_12bar), .A2(inbar[90]), .ZN(n764bar) );
  OR2_X1 U196 ( .A1(in_39), .A2(in_28), .ZN(n765) );
  AND2_X1 U196bar ( .A1(in_39bar), .A2(in_28bar), .ZN(n765bar) );
  OR2_X1 U197 ( .A1(in[109]), .A2(n763), .ZN(n780) );
  AND2_X1 U197bar ( .A1(inbar[109]), .A2(n763bar), .ZN(n780bar) );
  OR2_X1 U198 ( .A1(n762), .A2(n761), .ZN(n782) );
  AND2_X1 U198bar ( .A1(n762bar), .A2(n761bar), .ZN(n782bar) );
  OR2_X1 U199 ( .A1(in[138]), .A2(in[129]), .ZN(n761) );
  AND2_X1 U199bar ( .A1(inbar[138]), .A2(inbar[129]), .ZN(n761bar) );
  OR2_X1 U200 ( .A1(in[157]), .A2(n760), .ZN(n762) );
  AND2_X1 U200bar ( .A1(inbar[157]), .A2(n760bar), .ZN(n762bar) );
  OR2_X1 U201 ( .A1(in[182]), .A2(in[167]), .ZN(n760) );
  AND2_X1 U201bar ( .A1(inbar[182]), .A2(inbar[167]), .ZN(n760bar) );
  OR2_X1 U202 ( .A1(n759), .A2(n758), .ZN(n784) );
  AND2_X1 U202bar ( .A1(n759bar), .A2(n758bar), .ZN(n784bar) );
  OR2_X1 U203 ( .A1(n757), .A2(n756), .ZN(n758) );
  AND2_X1 U203bar ( .A1(n757bar), .A2(n756bar), .ZN(n758bar) );
  OR2_X1 U204 ( .A1(in[195]), .A2(in[184]), .ZN(n756) );
  AND2_X1 U204bar ( .A1(inbar[195]), .A2(inbar[184]), .ZN(n756bar) );
  OR2_X1 U205 ( .A1(in[196]), .A2(n755), .ZN(n757) );
  AND2_X1 U205bar ( .A1(inbar[196]), .A2(n755bar), .ZN(n757bar) );
  OR2_X1 U206 ( .A1(in[215]), .A2(in[209]), .ZN(n755) );
  AND2_X1 U206bar ( .A1(inbar[215]), .A2(inbar[209]), .ZN(n755bar) );
  OR2_X1 U207 ( .A1(n754), .A2(n753), .ZN(n759) );
  AND2_X1 U207bar ( .A1(n754bar), .A2(n753bar), .ZN(n759bar) );
  OR2_X1 U208 ( .A1(in[93]), .A2(in[233]), .ZN(n753) );
  AND2_X1 U208bar ( .A1(inbar[93]), .A2(inbar[233]), .ZN(n753bar) );
  OR2_X1 U209 ( .A1(in_1), .A2(n752), .ZN(n754) );
  AND2_X1 U209bar ( .A1(in_1bar), .A2(n752bar), .ZN(n754bar) );
  OR2_X1 U210 ( .A1(in_69), .A2(in_66), .ZN(n752) );
  AND2_X1 U210bar ( .A1(in_69bar), .A2(in_66bar), .ZN(n752bar) );
  OR2_X1 U211 ( .A1(n966), .A2(n751), .ZN(n787) );
  AND2_X1 U211bar ( .A1(n966bar), .A2(n751bar), .ZN(n787bar) );
  OR2_X1 U212 ( .A1(in[134]), .A2(n750), .ZN(n751) );
  AND2_X1 U212bar ( .A1(inbar[134]), .A2(n750bar), .ZN(n751bar) );
  OR2_X1 U213 ( .A1(n749), .A2(n748), .ZN(n966) );
  AND2_X1 U213bar ( .A1(n749bar), .A2(n748bar), .ZN(n966bar) );
  OR2_X1 U214 ( .A1(n747), .A2(n746), .ZN(n748) );
  AND2_X1 U214bar ( .A1(n747bar), .A2(n746bar), .ZN(n748bar) );
  OR2_X1 U215 ( .A1(n745), .A2(n744), .ZN(n746) );
  AND2_X1 U215bar ( .A1(n745bar), .A2(n744bar), .ZN(n746bar) );
  OR2_X1 U216 ( .A1(in[136]), .A2(in[121]), .ZN(n744) );
  AND2_X1 U216bar ( .A1(inbar[136]), .A2(inbar[121]), .ZN(n744bar) );
  OR2_X1 U217 ( .A1(in[186]), .A2(in[174]), .ZN(n745) );
  AND2_X1 U217bar ( .A1(inbar[186]), .A2(inbar[174]), .ZN(n745bar) );
  OR2_X1 U218 ( .A1(n743), .A2(n742), .ZN(n747) );
  AND2_X1 U218bar ( .A1(n743bar), .A2(n742bar), .ZN(n747bar) );
  OR2_X1 U219 ( .A1(in[198]), .A2(in[197]), .ZN(n742) );
  AND2_X1 U219bar ( .A1(inbar[198]), .A2(inbar[197]), .ZN(n742bar) );
  OR2_X1 U220 ( .A1(in[214]), .A2(in[199]), .ZN(n743) );
  AND2_X1 U220bar ( .A1(inbar[214]), .A2(inbar[199]), .ZN(n743bar) );
  OR2_X1 U221 ( .A1(n741), .A2(n740), .ZN(n749) );
  AND2_X1 U221bar ( .A1(n741bar), .A2(n740bar), .ZN(n749bar) );
  OR2_X1 U222 ( .A1(n739), .A2(n738), .ZN(n740) );
  AND2_X1 U222bar ( .A1(n739bar), .A2(n738bar), .ZN(n740bar) );
  OR2_X1 U223 ( .A1(in[231]), .A2(in[220]), .ZN(n738) );
  AND2_X1 U223bar ( .A1(inbar[231]), .A2(inbar[220]), .ZN(n738bar) );
  OR2_X1 U224 ( .A1(in_25), .A2(in[245]), .ZN(n739) );
  AND2_X1 U224bar ( .A1(in_25bar), .A2(inbar[245]), .ZN(n739bar) );
  OR2_X1 U225 ( .A1(n737), .A2(n736), .ZN(n741) );
  AND2_X1 U225bar ( .A1(n737bar), .A2(n736bar), .ZN(n741bar) );
  OR2_X1 U226 ( .A1(in_53), .A2(in_29), .ZN(n736) );
  AND2_X1 U226bar ( .A1(in_53bar), .A2(in_29bar), .ZN(n736bar) );
  OR2_X1 U227 ( .A1(in_79), .A2(in_74), .ZN(n737) );
  AND2_X1 U227bar ( .A1(in_79bar), .A2(in_74bar), .ZN(n737bar) );
  OR2_X1 U228 ( .A1(n735), .A2(n734), .ZN(n789) );
  AND2_X1 U228bar ( .A1(n735bar), .A2(n734bar), .ZN(n789bar) );
  OR2_X1 U229 ( .A1(in[152]), .A2(in[140]), .ZN(n734) );
  AND2_X1 U229bar ( .A1(inbar[152]), .A2(inbar[140]), .ZN(n734bar) );
  OR2_X1 U230 ( .A1(in[155]), .A2(n733), .ZN(n735) );
  AND2_X1 U230bar ( .A1(inbar[155]), .A2(n733bar), .ZN(n735bar) );
  OR2_X1 U231 ( .A1(in[166]), .A2(in[165]), .ZN(n733) );
  AND2_X1 U231bar ( .A1(inbar[166]), .A2(inbar[165]), .ZN(n733bar) );
  OR2_X1 U232 ( .A1(n732), .A2(n731), .ZN(n791) );
  AND2_X1 U232bar ( .A1(n732bar), .A2(n731bar), .ZN(n791bar) );
  OR2_X1 U233 ( .A1(n730), .A2(n729), .ZN(n731) );
  AND2_X1 U233bar ( .A1(n730bar), .A2(n729bar), .ZN(n731bar) );
  OR2_X1 U234 ( .A1(in[202]), .A2(in[185]), .ZN(n729) );
  AND2_X1 U234bar ( .A1(inbar[202]), .A2(inbar[185]), .ZN(n729bar) );
  OR2_X1 U235 ( .A1(in[211]), .A2(n728), .ZN(n730) );
  AND2_X1 U235bar ( .A1(inbar[211]), .A2(n728bar), .ZN(n730bar) );
  OR2_X1 U236 ( .A1(in[255]), .A2(in[253]), .ZN(n728) );
  AND2_X1 U236bar ( .A1(inbar[255]), .A2(inbar[253]), .ZN(n728bar) );
  OR2_X1 U237 ( .A1(n727), .A2(n726), .ZN(n732) );
  AND2_X1 U237bar ( .A1(n727bar), .A2(n726bar), .ZN(n732bar) );
  OR2_X1 U238 ( .A1(in_35), .A2(in_15), .ZN(n726) );
  AND2_X1 U238bar ( .A1(in_35bar), .A2(in_15bar), .ZN(n726bar) );
  OR2_X1 U239 ( .A1(in_36), .A2(n725), .ZN(n727) );
  AND2_X1 U239bar ( .A1(in_36bar), .A2(n725bar), .ZN(n727bar) );
  OR2_X1 U240 ( .A1(in_48), .A2(in_40), .ZN(n725) );
  AND2_X1 U240bar ( .A1(in_48bar), .A2(in_40bar), .ZN(n725bar) );
  OR2_X1 U241 ( .A1(n724), .A2(n723), .ZN(out[1]) );
  AND2_X1 U241bar ( .A1(n724bar), .A2(n723bar), .ZN(outbar[1]) );
  OR2_X1 U242 ( .A1(n722), .A2(n721), .ZN(n723) );
  AND2_X1 U242bar ( .A1(n722bar), .A2(n721bar), .ZN(n723bar) );
  OR2_X1 U243 ( .A1(n720), .A2(n719), .ZN(n721) );
  AND2_X1 U243bar ( .A1(n720bar), .A2(n719bar), .ZN(n721bar) );
  OR2_X1 U244 ( .A1(n921), .A2(n887), .ZN(n719) );
  AND2_X1 U244bar ( .A1(n921bar), .A2(n887bar), .ZN(n719bar) );
  OR2_X1 U245 ( .A1(n718), .A2(n717), .ZN(n887) );
  AND2_X1 U245bar ( .A1(n718bar), .A2(n717bar), .ZN(n887bar) );
  OR2_X1 U246 ( .A1(n716), .A2(n715), .ZN(n717) );
  AND2_X1 U246bar ( .A1(n716bar), .A2(n715bar), .ZN(n717bar) );
  OR2_X1 U247 ( .A1(n714), .A2(n713), .ZN(n715) );
  AND2_X1 U247bar ( .A1(n714bar), .A2(n713bar), .ZN(n715bar) );
  OR2_X1 U248 ( .A1(in[116]), .A2(in[110]), .ZN(n713) );
  AND2_X1 U248bar ( .A1(inbar[116]), .A2(inbar[110]), .ZN(n713bar) );
  OR2_X1 U249 ( .A1(in[133]), .A2(in[130]), .ZN(n714) );
  AND2_X1 U249bar ( .A1(inbar[133]), .A2(inbar[130]), .ZN(n714bar) );
  OR2_X1 U250 ( .A1(n712), .A2(n711), .ZN(n716) );
  AND2_X1 U250bar ( .A1(n712bar), .A2(n711bar), .ZN(n716bar) );
  OR2_X1 U251 ( .A1(in[203]), .A2(in[135]), .ZN(n711) );
  AND2_X1 U251bar ( .A1(inbar[203]), .A2(inbar[135]), .ZN(n711bar) );
  OR2_X1 U252 ( .A1(in[232]), .A2(in[223]), .ZN(n712) );
  AND2_X1 U252bar ( .A1(inbar[232]), .A2(inbar[223]), .ZN(n712bar) );
  OR2_X1 U253 ( .A1(n710), .A2(n709), .ZN(n718) );
  AND2_X1 U253bar ( .A1(n710bar), .A2(n709bar), .ZN(n718bar) );
  OR2_X1 U254 ( .A1(n708), .A2(n707), .ZN(n709) );
  AND2_X1 U254bar ( .A1(n708bar), .A2(n707bar), .ZN(n709bar) );
  OR2_X1 U255 ( .A1(in[255]), .A2(in[233]), .ZN(n707) );
  AND2_X1 U255bar ( .A1(inbar[255]), .A2(inbar[233]), .ZN(n707bar) );
  OR2_X1 U256 ( .A1(in_53), .A2(in_34), .ZN(n708) );
  AND2_X1 U256bar ( .A1(in_53bar), .A2(in_34bar), .ZN(n708bar) );
  OR2_X1 U257 ( .A1(n706), .A2(n705), .ZN(n710) );
  AND2_X1 U257bar ( .A1(n706bar), .A2(n705bar), .ZN(n710bar) );
  OR2_X1 U258 ( .A1(in_57), .A2(in_55), .ZN(n705) );
  AND2_X1 U258bar ( .A1(in_57bar), .A2(in_55bar), .ZN(n705bar) );
  OR2_X1 U259 ( .A1(in_68), .A2(in_67), .ZN(n706) );
  AND2_X1 U259bar ( .A1(in_68bar), .A2(in_67bar), .ZN(n706bar) );
  OR2_X1 U260 ( .A1(n704), .A2(n703), .ZN(n921) );
  AND2_X1 U260bar ( .A1(n704bar), .A2(n703bar), .ZN(n921bar) );
  OR2_X1 U261 ( .A1(n702), .A2(n701), .ZN(n703) );
  AND2_X1 U261bar ( .A1(n702bar), .A2(n701bar), .ZN(n703bar) );
  OR2_X1 U262 ( .A1(n700), .A2(n699), .ZN(n701) );
  AND2_X1 U262bar ( .A1(n700bar), .A2(n699bar), .ZN(n701bar) );
  OR2_X1 U263 ( .A1(n944), .A2(n872), .ZN(n699) );
  AND2_X1 U263bar ( .A1(n944bar), .A2(n872bar), .ZN(n699bar) );
  OR2_X1 U264 ( .A1(n698), .A2(n697), .ZN(n872) );
  AND2_X1 U264bar ( .A1(n698bar), .A2(n697bar), .ZN(n872bar) );
  OR2_X1 U265 ( .A1(n696), .A2(n695), .ZN(n697) );
  AND2_X1 U265bar ( .A1(n696bar), .A2(n695bar), .ZN(n697bar) );
  OR2_X1 U266 ( .A1(n694), .A2(n693), .ZN(n695) );
  AND2_X1 U266bar ( .A1(n694bar), .A2(n693bar), .ZN(n695bar) );
  OR2_X1 U267 ( .A1(in[121]), .A2(in[102]), .ZN(n693) );
  AND2_X1 U267bar ( .A1(inbar[121]), .A2(inbar[102]), .ZN(n693bar) );
  OR2_X1 U268 ( .A1(in[162]), .A2(in[161]), .ZN(n694) );
  AND2_X1 U268bar ( .A1(inbar[162]), .A2(inbar[161]), .ZN(n694bar) );
  OR2_X1 U269 ( .A1(n692), .A2(n691), .ZN(n696) );
  AND2_X1 U269bar ( .A1(n692bar), .A2(n691bar), .ZN(n696bar) );
  OR2_X1 U270 ( .A1(in[192]), .A2(in[178]), .ZN(n691) );
  AND2_X1 U270bar ( .A1(inbar[192]), .A2(inbar[178]), .ZN(n691bar) );
  OR2_X1 U271 ( .A1(in[244]), .A2(in[209]), .ZN(n692) );
  AND2_X1 U271bar ( .A1(inbar[244]), .A2(inbar[209]), .ZN(n692bar) );
  OR2_X1 U272 ( .A1(n690), .A2(n689), .ZN(n698) );
  AND2_X1 U272bar ( .A1(n690bar), .A2(n689bar), .ZN(n698bar) );
  OR2_X1 U273 ( .A1(n688), .A2(n687), .ZN(n689) );
  AND2_X1 U273bar ( .A1(n688bar), .A2(n687bar), .ZN(n689bar) );
  OR2_X1 U274 ( .A1(in[90]), .A2(in[254]), .ZN(n687) );
  AND2_X1 U274bar ( .A1(inbar[90]), .A2(inbar[254]), .ZN(n687bar) );
  OR2_X1 U275 ( .A1(in_36), .A2(in_32), .ZN(n688) );
  AND2_X1 U275bar ( .A1(in_36bar), .A2(in_32bar), .ZN(n688bar) );
  OR2_X1 U276 ( .A1(n686), .A2(n685), .ZN(n690) );
  AND2_X1 U276bar ( .A1(n686bar), .A2(n685bar), .ZN(n690bar) );
  OR2_X1 U277 ( .A1(in_62), .A2(in_37), .ZN(n685) );
  AND2_X1 U277bar ( .A1(in_62bar), .A2(in_37bar), .ZN(n685bar) );
  OR2_X1 U278 ( .A1(in_75), .A2(in_73), .ZN(n686) );
  AND2_X1 U278bar ( .A1(in_75bar), .A2(in_73bar), .ZN(n686bar) );
  OR2_X1 U279 ( .A1(n684), .A2(n683), .ZN(n944) );
  AND2_X1 U279bar ( .A1(n684bar), .A2(n683bar), .ZN(n944bar) );
  OR2_X1 U280 ( .A1(n682), .A2(n681), .ZN(n683) );
  AND2_X1 U280bar ( .A1(n682bar), .A2(n681bar), .ZN(n683bar) );
  OR2_X1 U281 ( .A1(n680), .A2(n679), .ZN(n681) );
  AND2_X1 U281bar ( .A1(n680bar), .A2(n679bar), .ZN(n681bar) );
  OR2_X1 U282 ( .A1(in[171]), .A2(in[153]), .ZN(n679) );
  AND2_X1 U282bar ( .A1(inbar[171]), .A2(inbar[153]), .ZN(n679bar) );
  OR2_X1 U283 ( .A1(in[187]), .A2(in[176]), .ZN(n680) );
  AND2_X1 U283bar ( .A1(inbar[187]), .A2(inbar[176]), .ZN(n680bar) );
  OR2_X1 U284 ( .A1(n678), .A2(n677), .ZN(n682) );
  AND2_X1 U284bar ( .A1(n678bar), .A2(n677bar), .ZN(n682bar) );
  OR2_X1 U285 ( .A1(in[245]), .A2(in[211]), .ZN(n677) );
  AND2_X1 U285bar ( .A1(inbar[245]), .A2(inbar[211]), .ZN(n677bar) );
  OR2_X1 U286 ( .A1(in[97]), .A2(in[88]), .ZN(n678) );
  AND2_X1 U286bar ( .A1(inbar[97]), .A2(inbar[88]), .ZN(n678bar) );
  OR2_X1 U287 ( .A1(n676), .A2(n675), .ZN(n684) );
  AND2_X1 U287bar ( .A1(n676bar), .A2(n675bar), .ZN(n684bar) );
  OR2_X1 U288 ( .A1(n674), .A2(n673), .ZN(n675) );
  AND2_X1 U288bar ( .A1(n674bar), .A2(n673bar), .ZN(n675bar) );
  OR2_X1 U289 ( .A1(in_10), .A2(in_0), .ZN(n673) );
  AND2_X1 U289bar ( .A1(in_10bar), .A2(in_0bar), .ZN(n673bar) );
  OR2_X1 U290 ( .A1(in_59), .A2(in_5), .ZN(n674) );
  AND2_X1 U290bar ( .A1(in_59bar), .A2(in_5bar), .ZN(n674bar) );
  OR2_X1 U291 ( .A1(n672), .A2(n671), .ZN(n676) );
  AND2_X1 U291bar ( .A1(n672bar), .A2(n671bar), .ZN(n676bar) );
  OR2_X1 U292 ( .A1(in_60), .A2(in_6), .ZN(n671) );
  AND2_X1 U292bar ( .A1(in_60bar), .A2(in_6bar), .ZN(n671bar) );
  OR2_X1 U293 ( .A1(in_77), .A2(in_69), .ZN(n672) );
  AND2_X1 U293bar ( .A1(in_77bar), .A2(in_69bar), .ZN(n672bar) );
  OR2_X1 U294 ( .A1(in[113]), .A2(n864), .ZN(n700) );
  AND2_X1 U294bar ( .A1(inbar[113]), .A2(n864bar), .ZN(n700bar) );
  OR2_X1 U295 ( .A1(n670), .A2(n669), .ZN(n864) );
  AND2_X1 U295bar ( .A1(n670bar), .A2(n669bar), .ZN(n864bar) );
  OR2_X1 U296 ( .A1(n668), .A2(n667), .ZN(n669) );
  AND2_X1 U296bar ( .A1(n668bar), .A2(n667bar), .ZN(n669bar) );
  OR2_X1 U297 ( .A1(n666), .A2(n665), .ZN(n667) );
  AND2_X1 U297bar ( .A1(n666bar), .A2(n665bar), .ZN(n667bar) );
  OR2_X1 U298 ( .A1(in[125]), .A2(in[107]), .ZN(n665) );
  AND2_X1 U298bar ( .A1(inbar[125]), .A2(inbar[107]), .ZN(n665bar) );
  OR2_X1 U299 ( .A1(in[138]), .A2(in[126]), .ZN(n666) );
  AND2_X1 U299bar ( .A1(inbar[138]), .A2(inbar[126]), .ZN(n666bar) );
  OR2_X1 U300 ( .A1(n664), .A2(n663), .ZN(n668) );
  AND2_X1 U300bar ( .A1(n664bar), .A2(n663bar), .ZN(n668bar) );
  OR2_X1 U301 ( .A1(in[189]), .A2(in[143]), .ZN(n663) );
  AND2_X1 U301bar ( .A1(inbar[189]), .A2(inbar[143]), .ZN(n663bar) );
  OR2_X1 U302 ( .A1(in[99]), .A2(in[214]), .ZN(n664) );
  AND2_X1 U302bar ( .A1(inbar[99]), .A2(inbar[214]), .ZN(n664bar) );
  OR2_X1 U303 ( .A1(n662), .A2(n661), .ZN(n670) );
  AND2_X1 U303bar ( .A1(n662bar), .A2(n661bar), .ZN(n670bar) );
  OR2_X1 U304 ( .A1(n660), .A2(n659), .ZN(n661) );
  AND2_X1 U304bar ( .A1(n660bar), .A2(n659bar), .ZN(n661bar) );
  OR2_X1 U305 ( .A1(in_15), .A2(in_12), .ZN(n659) );
  AND2_X1 U305bar ( .A1(in_15bar), .A2(in_12bar), .ZN(n659bar) );
  OR2_X1 U306 ( .A1(in_20), .A2(in_2), .ZN(n660) );
  AND2_X1 U306bar ( .A1(in_20bar), .A2(in_2bar), .ZN(n660bar) );
  OR2_X1 U307 ( .A1(n658), .A2(n657), .ZN(n662) );
  AND2_X1 U307bar ( .A1(n658bar), .A2(n657bar), .ZN(n662bar) );
  OR2_X1 U308 ( .A1(in_30), .A2(in_3), .ZN(n657) );
  AND2_X1 U308bar ( .A1(in_30bar), .A2(in_3bar), .ZN(n657bar) );
  OR2_X1 U309 ( .A1(in_4), .A2(in_38), .ZN(n658) );
  AND2_X1 U309bar ( .A1(in_4bar), .A2(in_38bar), .ZN(n658bar) );
  OR2_X1 U310 ( .A1(n656), .A2(n655), .ZN(n702) );
  AND2_X1 U310bar ( .A1(n656bar), .A2(n655bar), .ZN(n702bar) );
  OR2_X1 U311 ( .A1(in[148]), .A2(in[137]), .ZN(n655) );
  AND2_X1 U311bar ( .A1(inbar[148]), .A2(inbar[137]), .ZN(n655bar) );
  OR2_X1 U312 ( .A1(in[149]), .A2(n654), .ZN(n656) );
  AND2_X1 U312bar ( .A1(inbar[149]), .A2(n654bar), .ZN(n656bar) );
  OR2_X1 U313 ( .A1(in[195]), .A2(in[190]), .ZN(n654) );
  AND2_X1 U313bar ( .A1(inbar[195]), .A2(inbar[190]), .ZN(n654bar) );
  OR2_X1 U314 ( .A1(n653), .A2(n652), .ZN(n704) );
  AND2_X1 U314bar ( .A1(n653bar), .A2(n652bar), .ZN(n704bar) );
  OR2_X1 U315 ( .A1(n651), .A2(n650), .ZN(n652) );
  AND2_X1 U315bar ( .A1(n651bar), .A2(n650bar), .ZN(n652bar) );
  OR2_X1 U316 ( .A1(in[98]), .A2(in[197]), .ZN(n650) );
  AND2_X1 U316bar ( .A1(inbar[98]), .A2(inbar[197]), .ZN(n650bar) );
  OR2_X1 U317 ( .A1(in_11), .A2(n649), .ZN(n651) );
  AND2_X1 U317bar ( .A1(in_11bar), .A2(n649bar), .ZN(n651bar) );
  OR2_X1 U318 ( .A1(in_26), .A2(in_14), .ZN(n649) );
  AND2_X1 U318bar ( .A1(in_26bar), .A2(in_14bar), .ZN(n649bar) );
  OR2_X1 U319 ( .A1(n648), .A2(n647), .ZN(n653) );
  AND2_X1 U319bar ( .A1(n648bar), .A2(n647bar), .ZN(n653bar) );
  OR2_X1 U320 ( .A1(in_35), .A2(in_27), .ZN(n647) );
  AND2_X1 U320bar ( .A1(in_35bar), .A2(in_27bar), .ZN(n647bar) );
  OR2_X1 U321 ( .A1(in_50), .A2(n646), .ZN(n648) );
  AND2_X1 U321bar ( .A1(in_50bar), .A2(n646bar), .ZN(n648bar) );
  OR2_X1 U322 ( .A1(in_78), .A2(in_61), .ZN(n646) );
  AND2_X1 U322bar ( .A1(in_78bar), .A2(in_61bar), .ZN(n646bar) );
  OR2_X1 U323 ( .A1(n942), .A2(n645), .ZN(n720) );
  AND2_X1 U323bar ( .A1(n942bar), .A2(n645bar), .ZN(n720bar) );
  OR2_X1 U324 ( .A1(in[106]), .A2(n863), .ZN(n645) );
  AND2_X1 U324bar ( .A1(inbar[106]), .A2(n863bar), .ZN(n645bar) );
  OR2_X1 U325 ( .A1(n644), .A2(n643), .ZN(n863) );
  AND2_X1 U325bar ( .A1(n644bar), .A2(n643bar), .ZN(n863bar) );
  OR2_X1 U326 ( .A1(n642), .A2(n641), .ZN(n643) );
  AND2_X1 U326bar ( .A1(n642bar), .A2(n641bar), .ZN(n643bar) );
  OR2_X1 U327 ( .A1(n640), .A2(n639), .ZN(n641) );
  AND2_X1 U327bar ( .A1(n640bar), .A2(n639bar), .ZN(n641bar) );
  OR2_X1 U328 ( .A1(in[127]), .A2(in[122]), .ZN(n639) );
  AND2_X1 U328bar ( .A1(inbar[127]), .A2(inbar[122]), .ZN(n639bar) );
  OR2_X1 U329 ( .A1(in[156]), .A2(in[132]), .ZN(n640) );
  AND2_X1 U329bar ( .A1(inbar[156]), .A2(inbar[132]), .ZN(n640bar) );
  OR2_X1 U330 ( .A1(n638), .A2(n637), .ZN(n642) );
  AND2_X1 U330bar ( .A1(n638bar), .A2(n637bar), .ZN(n642bar) );
  OR2_X1 U331 ( .A1(in[159]), .A2(in[157]), .ZN(n637) );
  AND2_X1 U331bar ( .A1(inbar[159]), .A2(inbar[157]), .ZN(n637bar) );
  OR2_X1 U332 ( .A1(in[185]), .A2(in[169]), .ZN(n638) );
  AND2_X1 U332bar ( .A1(inbar[185]), .A2(inbar[169]), .ZN(n638bar) );
  OR2_X1 U333 ( .A1(n636), .A2(n635), .ZN(n644) );
  AND2_X1 U333bar ( .A1(n636bar), .A2(n635bar), .ZN(n644bar) );
  OR2_X1 U334 ( .A1(n634), .A2(n633), .ZN(n635) );
  AND2_X1 U334bar ( .A1(n634bar), .A2(n633bar), .ZN(n635bar) );
  OR2_X1 U335 ( .A1(in[239]), .A2(in[218]), .ZN(n633) );
  AND2_X1 U335bar ( .A1(inbar[239]), .A2(inbar[218]), .ZN(n633bar) );
  OR2_X1 U336 ( .A1(in_13), .A2(in[87]), .ZN(n634) );
  AND2_X1 U336bar ( .A1(in_13bar), .A2(inbar[87]), .ZN(n634bar) );
  OR2_X1 U337 ( .A1(n632), .A2(n631), .ZN(n636) );
  AND2_X1 U337bar ( .A1(n632bar), .A2(n631bar), .ZN(n636bar) );
  OR2_X1 U338 ( .A1(in_72), .A2(in_70), .ZN(n631) );
  AND2_X1 U338bar ( .A1(in_72bar), .A2(in_70bar), .ZN(n631bar) );
  OR2_X1 U339 ( .A1(in_80), .A2(in_74), .ZN(n632) );
  AND2_X1 U339bar ( .A1(in_80bar), .A2(in_74bar), .ZN(n632bar) );
  OR2_X1 U340 ( .A1(n630), .A2(n629), .ZN(n942) );
  AND2_X1 U340bar ( .A1(n630bar), .A2(n629bar), .ZN(n942bar) );
  OR2_X1 U341 ( .A1(n628), .A2(n627), .ZN(n629) );
  AND2_X1 U341bar ( .A1(n628bar), .A2(n627bar), .ZN(n629bar) );
  OR2_X1 U342 ( .A1(n626), .A2(n625), .ZN(n627) );
  AND2_X1 U342bar ( .A1(n626bar), .A2(n625bar), .ZN(n627bar) );
  OR2_X1 U343 ( .A1(in[146]), .A2(in[100]), .ZN(n625) );
  AND2_X1 U343bar ( .A1(inbar[146]), .A2(inbar[100]), .ZN(n625bar) );
  OR2_X1 U344 ( .A1(in[168]), .A2(in[152]), .ZN(n626) );
  AND2_X1 U344bar ( .A1(inbar[168]), .A2(inbar[152]), .ZN(n626bar) );
  OR2_X1 U345 ( .A1(n624), .A2(n623), .ZN(n628) );
  AND2_X1 U345bar ( .A1(n624bar), .A2(n623bar), .ZN(n628bar) );
  OR2_X1 U346 ( .A1(in[199]), .A2(in[182]), .ZN(n623) );
  AND2_X1 U346bar ( .A1(inbar[199]), .A2(inbar[182]), .ZN(n623bar) );
  OR2_X1 U347 ( .A1(in[236]), .A2(in[204]), .ZN(n624) );
  AND2_X1 U347bar ( .A1(inbar[236]), .A2(inbar[204]), .ZN(n624bar) );
  OR2_X1 U348 ( .A1(n622), .A2(n621), .ZN(n630) );
  AND2_X1 U348bar ( .A1(n622bar), .A2(n621bar), .ZN(n630bar) );
  OR2_X1 U349 ( .A1(n620), .A2(n619), .ZN(n621) );
  AND2_X1 U349bar ( .A1(n620bar), .A2(n619bar), .ZN(n621bar) );
  OR2_X1 U350 ( .A1(in[89]), .A2(in[246]), .ZN(n619) );
  AND2_X1 U350bar ( .A1(inbar[89]), .A2(inbar[246]), .ZN(n619bar) );
  OR2_X1 U351 ( .A1(in[95]), .A2(in[92]), .ZN(n620) );
  AND2_X1 U351bar ( .A1(inbar[95]), .A2(inbar[92]), .ZN(n620bar) );
  OR2_X1 U352 ( .A1(n618), .A2(n617), .ZN(n622) );
  AND2_X1 U352bar ( .A1(n618bar), .A2(n617bar), .ZN(n622bar) );
  OR2_X1 U353 ( .A1(in_22), .A2(in_16), .ZN(n617) );
  AND2_X1 U353bar ( .A1(in_22bar), .A2(in_16bar), .ZN(n617bar) );
  OR2_X1 U354 ( .A1(in_51), .A2(in_49), .ZN(n618) );
  AND2_X1 U354bar ( .A1(in_51bar), .A2(in_49bar), .ZN(n618bar) );
  OR2_X1 U355 ( .A1(n616), .A2(n615), .ZN(n722) );
  AND2_X1 U355bar ( .A1(n616bar), .A2(n615bar), .ZN(n722bar) );
  OR2_X1 U356 ( .A1(in[158]), .A2(in[115]), .ZN(n615) );
  AND2_X1 U356bar ( .A1(inbar[158]), .A2(inbar[115]), .ZN(n615bar) );
  OR2_X1 U357 ( .A1(in[163]), .A2(n614), .ZN(n616) );
  AND2_X1 U357bar ( .A1(inbar[163]), .A2(n614bar), .ZN(n616bar) );
  OR2_X1 U358 ( .A1(in[206]), .A2(in[165]), .ZN(n614) );
  AND2_X1 U358bar ( .A1(inbar[206]), .A2(inbar[165]), .ZN(n614bar) );
  OR2_X1 U359 ( .A1(n613), .A2(n612), .ZN(n724) );
  AND2_X1 U359bar ( .A1(n613bar), .A2(n612bar), .ZN(n724bar) );
  OR2_X1 U360 ( .A1(n611), .A2(n610), .ZN(n612) );
  AND2_X1 U360bar ( .A1(n611bar), .A2(n610bar), .ZN(n612bar) );
  OR2_X1 U361 ( .A1(in[213]), .A2(in[207]), .ZN(n610) );
  AND2_X1 U361bar ( .A1(inbar[213]), .A2(inbar[207]), .ZN(n610bar) );
  OR2_X1 U362 ( .A1(in[215]), .A2(n609), .ZN(n611) );
  AND2_X1 U362bar ( .A1(inbar[215]), .A2(n609bar), .ZN(n611bar) );
  OR2_X1 U363 ( .A1(in[230]), .A2(in[220]), .ZN(n609) );
  AND2_X1 U363bar ( .A1(inbar[230]), .A2(inbar[220]), .ZN(n609bar) );
  OR2_X1 U364 ( .A1(n608), .A2(n607), .ZN(n613) );
  AND2_X1 U364bar ( .A1(n608bar), .A2(n607bar), .ZN(n613bar) );
  OR2_X1 U365 ( .A1(in[251]), .A2(in[234]), .ZN(n607) );
  AND2_X1 U365bar ( .A1(inbar[251]), .A2(inbar[234]), .ZN(n607bar) );
  OR2_X1 U366 ( .A1(in_17), .A2(n606), .ZN(n608) );
  AND2_X1 U366bar ( .A1(in_17bar), .A2(n606bar), .ZN(n608bar) );
  OR2_X1 U367 ( .A1(in_65), .A2(in_56), .ZN(n606) );
  AND2_X1 U367bar ( .A1(in_65bar), .A2(in_56bar), .ZN(n606bar) );
  OR2_X1 U368 ( .A1(n605), .A2(n604), .ZN(out[0]) );
  AND2_X1 U368bar ( .A1(n605bar), .A2(n604bar), .ZN(outbar[0]) );
  OR2_X1 U369 ( .A1(n603), .A2(n602), .ZN(n604) );
  AND2_X1 U369bar ( .A1(n603bar), .A2(n602bar), .ZN(n604bar) );
  OR2_X1 U370 ( .A1(n601), .A2(n600), .ZN(n602) );
  AND2_X1 U370bar ( .A1(n601bar), .A2(n600bar), .ZN(n602bar) );
  OR2_X1 U371 ( .A1(n820), .A2(n785), .ZN(n600) );
  AND2_X1 U371bar ( .A1(n820bar), .A2(n785bar), .ZN(n600bar) );
  OR2_X1 U372 ( .A1(n599), .A2(n598), .ZN(n785) );
  AND2_X1 U372bar ( .A1(n599bar), .A2(n598bar), .ZN(n785bar) );
  OR2_X1 U373 ( .A1(n597), .A2(n596), .ZN(n598) );
  AND2_X1 U373bar ( .A1(n597bar), .A2(n596bar), .ZN(n598bar) );
  OR2_X1 U374 ( .A1(n595), .A2(n594), .ZN(n596) );
  AND2_X1 U374bar ( .A1(n595bar), .A2(n594bar), .ZN(n596bar) );
  OR2_X1 U375 ( .A1(in[135]), .A2(in[104]), .ZN(n594) );
  AND2_X1 U375bar ( .A1(inbar[135]), .A2(inbar[104]), .ZN(n594bar) );
  OR2_X1 U376 ( .A1(in[188]), .A2(in[178]), .ZN(n595) );
  AND2_X1 U376bar ( .A1(inbar[188]), .A2(inbar[178]), .ZN(n595bar) );
  OR2_X1 U377 ( .A1(n593), .A2(n592), .ZN(n597) );
  AND2_X1 U377bar ( .A1(n593bar), .A2(n592bar), .ZN(n597bar) );
  OR2_X1 U378 ( .A1(in[217]), .A2(in[194]), .ZN(n592) );
  AND2_X1 U378bar ( .A1(inbar[217]), .A2(inbar[194]), .ZN(n592bar) );
  OR2_X1 U379 ( .A1(in[237]), .A2(in[218]), .ZN(n593) );
  AND2_X1 U379bar ( .A1(inbar[237]), .A2(inbar[218]), .ZN(n593bar) );
  OR2_X1 U380 ( .A1(n591), .A2(n590), .ZN(n599) );
  AND2_X1 U380bar ( .A1(n591bar), .A2(n590bar), .ZN(n599bar) );
  OR2_X1 U381 ( .A1(n589), .A2(n588), .ZN(n590) );
  AND2_X1 U381bar ( .A1(n589bar), .A2(n588bar), .ZN(n590bar) );
  OR2_X1 U382 ( .A1(in_2), .A2(in_10), .ZN(n588) );
  AND2_X1 U382bar ( .A1(in_2bar), .A2(in_10bar), .ZN(n588bar) );
  OR2_X1 U383 ( .A1(in_47), .A2(in_22), .ZN(n589) );
  AND2_X1 U383bar ( .A1(in_47bar), .A2(in_22bar), .ZN(n589bar) );
  OR2_X1 U384 ( .A1(n587), .A2(n586), .ZN(n591) );
  AND2_X1 U384bar ( .A1(n587bar), .A2(n586bar), .ZN(n591bar) );
  OR2_X1 U385 ( .A1(in_56), .A2(in_54), .ZN(n586) );
  AND2_X1 U385bar ( .A1(in_56bar), .A2(in_54bar), .ZN(n586bar) );
  OR2_X1 U386 ( .A1(in_63), .A2(in_61), .ZN(n587) );
  AND2_X1 U386bar ( .A1(in_63bar), .A2(in_61bar), .ZN(n587bar) );
  OR2_X1 U387 ( .A1(n585), .A2(n584), .ZN(n820) );
  AND2_X1 U387bar ( .A1(n585bar), .A2(n584bar), .ZN(n820bar) );
  OR2_X1 U388 ( .A1(n583), .A2(n582), .ZN(n584) );
  AND2_X1 U388bar ( .A1(n583bar), .A2(n582bar), .ZN(n584bar) );
  OR2_X1 U389 ( .A1(n581), .A2(n580), .ZN(n582) );
  AND2_X1 U389bar ( .A1(n581bar), .A2(n580bar), .ZN(n582bar) );
  OR2_X1 U390 ( .A1(in[158]), .A2(in[142]), .ZN(n580) );
  AND2_X1 U390bar ( .A1(inbar[158]), .A2(inbar[142]), .ZN(n580bar) );
  OR2_X1 U391 ( .A1(in[175]), .A2(in[164]), .ZN(n581) );
  AND2_X1 U391bar ( .A1(inbar[175]), .A2(inbar[164]), .ZN(n581bar) );
  OR2_X1 U392 ( .A1(n579), .A2(n578), .ZN(n583) );
  AND2_X1 U392bar ( .A1(n579bar), .A2(n578bar), .ZN(n583bar) );
  OR2_X1 U393 ( .A1(in[228]), .A2(in[204]), .ZN(n578) );
  AND2_X1 U393bar ( .A1(inbar[228]), .A2(inbar[204]), .ZN(n578bar) );
  OR2_X1 U394 ( .A1(in[91]), .A2(in[87]), .ZN(n579) );
  AND2_X1 U394bar ( .A1(inbar[91]), .A2(inbar[87]), .ZN(n579bar) );
  OR2_X1 U395 ( .A1(n577), .A2(n576), .ZN(n585) );
  AND2_X1 U395bar ( .A1(n577bar), .A2(n576bar), .ZN(n585bar) );
  OR2_X1 U396 ( .A1(n575), .A2(n574), .ZN(n576) );
  AND2_X1 U396bar ( .A1(n575bar), .A2(n574bar), .ZN(n576bar) );
  OR2_X1 U397 ( .A1(in_21), .A2(in_11), .ZN(n574) );
  AND2_X1 U397bar ( .A1(in_21bar), .A2(in_11bar), .ZN(n574bar) );
  OR2_X1 U398 ( .A1(in_5), .A2(in_3), .ZN(n575) );
  AND2_X1 U398bar ( .A1(in_5bar), .A2(in_3bar), .ZN(n575bar) );
  OR2_X1 U399 ( .A1(n573), .A2(n572), .ZN(n577) );
  AND2_X1 U399bar ( .A1(n573bar), .A2(n572bar), .ZN(n577bar) );
  OR2_X1 U400 ( .A1(in_68), .A2(in_64), .ZN(n572) );
  AND2_X1 U400bar ( .A1(in_68bar), .A2(in_64bar), .ZN(n572bar) );
  OR2_X1 U401 ( .A1(in_76), .A2(in_73), .ZN(n573) );
  AND2_X1 U401bar ( .A1(in_76bar), .A2(in_73bar), .ZN(n573bar) );
  OR2_X1 U402 ( .A1(n778), .A2(n571), .ZN(n601) );
  AND2_X1 U402bar ( .A1(n778bar), .A2(n571bar), .ZN(n601bar) );
  OR2_X1 U403 ( .A1(in[100]), .A2(n965), .ZN(n571) );
  AND2_X1 U403bar ( .A1(inbar[100]), .A2(n965bar), .ZN(n571bar) );
  OR2_X1 U404 ( .A1(n570), .A2(n569), .ZN(n965) );
  AND2_X1 U404bar ( .A1(n570bar), .A2(n569bar), .ZN(n965bar) );
  OR2_X1 U405 ( .A1(n568), .A2(n567), .ZN(n569) );
  AND2_X1 U405bar ( .A1(n568bar), .A2(n567bar), .ZN(n569bar) );
  OR2_X1 U406 ( .A1(n566), .A2(n565), .ZN(n567) );
  AND2_X1 U406bar ( .A1(n566bar), .A2(n565bar), .ZN(n567bar) );
  OR2_X1 U407 ( .A1(n817), .A2(n750), .ZN(n565) );
  AND2_X1 U407bar ( .A1(n817bar), .A2(n750bar), .ZN(n565bar) );
  OR2_X1 U408 ( .A1(n564), .A2(n563), .ZN(n750) );
  AND2_X1 U408bar ( .A1(n564bar), .A2(n563bar), .ZN(n750bar) );
  OR2_X1 U409 ( .A1(n562), .A2(n561), .ZN(n563) );
  AND2_X1 U409bar ( .A1(n562bar), .A2(n561bar), .ZN(n563bar) );
  OR2_X1 U410 ( .A1(n560), .A2(n559), .ZN(n561) );
  AND2_X1 U410bar ( .A1(n560bar), .A2(n559bar), .ZN(n561bar) );
  OR2_X1 U411 ( .A1(in[119]), .A2(in[103]), .ZN(n559) );
  AND2_X1 U411bar ( .A1(inbar[119]), .A2(inbar[103]), .ZN(n559bar) );
  OR2_X1 U412 ( .A1(in[137]), .A2(in[133]), .ZN(n560) );
  AND2_X1 U412bar ( .A1(inbar[137]), .A2(inbar[133]), .ZN(n560bar) );
  OR2_X1 U413 ( .A1(n558), .A2(n557), .ZN(n562) );
  AND2_X1 U413bar ( .A1(n558bar), .A2(n557bar), .ZN(n562bar) );
  OR2_X1 U414 ( .A1(in[176]), .A2(in[173]), .ZN(n557) );
  AND2_X1 U414bar ( .A1(inbar[176]), .A2(inbar[173]), .ZN(n557bar) );
  OR2_X1 U415 ( .A1(in[210]), .A2(in[181]), .ZN(n558) );
  AND2_X1 U415bar ( .A1(inbar[210]), .A2(inbar[181]), .ZN(n558bar) );
  OR2_X1 U416 ( .A1(n556), .A2(n555), .ZN(n564) );
  AND2_X1 U416bar ( .A1(n556bar), .A2(n555bar), .ZN(n564bar) );
  OR2_X1 U417 ( .A1(n554), .A2(n553), .ZN(n555) );
  AND2_X1 U417bar ( .A1(n554bar), .A2(n553bar), .ZN(n555bar) );
  OR2_X1 U418 ( .A1(in_13), .A2(in[234]), .ZN(n553) );
  AND2_X1 U418bar ( .A1(in_13bar), .A2(inbar[234]), .ZN(n553bar) );
  OR2_X1 U419 ( .A1(in_38), .A2(in_32), .ZN(n554) );
  AND2_X1 U419bar ( .A1(in_38bar), .A2(in_32bar), .ZN(n554bar) );
  OR2_X1 U420 ( .A1(n552), .A2(n551), .ZN(n556) );
  AND2_X1 U420bar ( .A1(n552bar), .A2(n551bar), .ZN(n556bar) );
  OR2_X1 U421 ( .A1(in_42), .A2(in_41), .ZN(n551) );
  AND2_X1 U421bar ( .A1(in_42bar), .A2(in_41bar), .ZN(n551bar) );
  OR2_X1 U422 ( .A1(in_7), .A2(in_49), .ZN(n552) );
  AND2_X1 U422bar ( .A1(in_7bar), .A2(in_49bar), .ZN(n552bar) );
  OR2_X1 U423 ( .A1(n550), .A2(n549), .ZN(n817) );
  AND2_X1 U423bar ( .A1(n550bar), .A2(n549bar), .ZN(n817bar) );
  OR2_X1 U424 ( .A1(n548), .A2(n547), .ZN(n549) );
  AND2_X1 U424bar ( .A1(n548bar), .A2(n547bar), .ZN(n549bar) );
  OR2_X1 U425 ( .A1(n546), .A2(n545), .ZN(n547) );
  AND2_X1 U425bar ( .A1(n546bar), .A2(n545bar), .ZN(n547bar) );
  OR2_X1 U426 ( .A1(in[159]), .A2(in[105]), .ZN(n545) );
  AND2_X1 U426bar ( .A1(inbar[159]), .A2(inbar[105]), .ZN(n545bar) );
  OR2_X1 U427 ( .A1(in[206]), .A2(in[183]), .ZN(n546) );
  AND2_X1 U427bar ( .A1(inbar[206]), .A2(inbar[183]), .ZN(n546bar) );
  OR2_X1 U428 ( .A1(n544), .A2(n543), .ZN(n548) );
  AND2_X1 U428bar ( .A1(n544bar), .A2(n543bar), .ZN(n548bar) );
  OR2_X1 U429 ( .A1(in[229]), .A2(in[219]), .ZN(n543) );
  AND2_X1 U429bar ( .A1(inbar[229]), .A2(inbar[219]), .ZN(n543bar) );
  OR2_X1 U430 ( .A1(in[235]), .A2(in[232]), .ZN(n544) );
  AND2_X1 U430bar ( .A1(inbar[235]), .A2(inbar[232]), .ZN(n544bar) );
  OR2_X1 U431 ( .A1(n542), .A2(n541), .ZN(n550) );
  AND2_X1 U431bar ( .A1(n542bar), .A2(n541bar), .ZN(n550bar) );
  OR2_X1 U432 ( .A1(n540), .A2(n539), .ZN(n541) );
  AND2_X1 U432bar ( .A1(n540bar), .A2(n539bar), .ZN(n541bar) );
  OR2_X1 U433 ( .A1(in[249]), .A2(in[242]), .ZN(n539) );
  AND2_X1 U433bar ( .A1(inbar[249]), .A2(inbar[242]), .ZN(n539bar) );
  OR2_X1 U434 ( .A1(in[89]), .A2(in[254]), .ZN(n540) );
  AND2_X1 U434bar ( .A1(inbar[89]), .A2(inbar[254]), .ZN(n540bar) );
  OR2_X1 U435 ( .A1(n538), .A2(n537), .ZN(n542) );
  AND2_X1 U435bar ( .A1(n538bar), .A2(n537bar), .ZN(n542bar) );
  OR2_X1 U436 ( .A1(in_14), .A2(in[99]), .ZN(n537) );
  AND2_X1 U436bar ( .A1(in_14bar), .A2(inbar[99]), .ZN(n537bar) );
  OR2_X1 U437 ( .A1(in_60), .A2(in_18), .ZN(n538) );
  AND2_X1 U437bar ( .A1(in_60bar), .A2(in_18bar), .ZN(n538bar) );
  OR2_X1 U438 ( .A1(in[113]), .A2(n763), .ZN(n566) );
  AND2_X1 U438bar ( .A1(inbar[113]), .A2(n763bar), .ZN(n566bar) );
  OR2_X1 U439 ( .A1(n536), .A2(n535), .ZN(n763) );
  AND2_X1 U439bar ( .A1(n536bar), .A2(n535bar), .ZN(n763bar) );
  OR2_X1 U440 ( .A1(n534), .A2(n533), .ZN(n535) );
  AND2_X1 U440bar ( .A1(n534bar), .A2(n533bar), .ZN(n535bar) );
  OR2_X1 U441 ( .A1(n532), .A2(n531), .ZN(n533) );
  AND2_X1 U441bar ( .A1(n532bar), .A2(n531bar), .ZN(n533bar) );
  OR2_X1 U442 ( .A1(in[115]), .A2(in[110]), .ZN(n531) );
  AND2_X1 U442bar ( .A1(inbar[115]), .A2(inbar[110]), .ZN(n531bar) );
  OR2_X1 U443 ( .A1(in[125]), .A2(in[117]), .ZN(n532) );
  AND2_X1 U443bar ( .A1(inbar[125]), .A2(inbar[117]), .ZN(n532bar) );
  OR2_X1 U444 ( .A1(n530), .A2(n529), .ZN(n534) );
  AND2_X1 U444bar ( .A1(n530bar), .A2(n529bar), .ZN(n534bar) );
  OR2_X1 U445 ( .A1(in[180]), .A2(in[128]), .ZN(n529) );
  AND2_X1 U445bar ( .A1(inbar[180]), .A2(inbar[128]), .ZN(n529bar) );
  OR2_X1 U446 ( .A1(in[205]), .A2(in[201]), .ZN(n530) );
  AND2_X1 U446bar ( .A1(inbar[205]), .A2(inbar[201]), .ZN(n530bar) );
  OR2_X1 U447 ( .A1(n528), .A2(n527), .ZN(n536) );
  AND2_X1 U447bar ( .A1(n528bar), .A2(n527bar), .ZN(n536bar) );
  OR2_X1 U448 ( .A1(n526), .A2(n525), .ZN(n527) );
  AND2_X1 U448bar ( .A1(n526bar), .A2(n525bar), .ZN(n527bar) );
  OR2_X1 U449 ( .A1(in[244]), .A2(in[239]), .ZN(n525) );
  AND2_X1 U449bar ( .A1(inbar[244]), .A2(inbar[239]), .ZN(n525bar) );
  OR2_X1 U450 ( .A1(in[95]), .A2(in[83]), .ZN(n526) );
  AND2_X1 U450bar ( .A1(inbar[95]), .A2(inbar[83]), .ZN(n526bar) );
  OR2_X1 U451 ( .A1(n524), .A2(n523), .ZN(n528) );
  AND2_X1 U451bar ( .A1(n524bar), .A2(n523bar), .ZN(n528bar) );
  OR2_X1 U452 ( .A1(in_24), .A2(in[97]), .ZN(n523) );
  AND2_X1 U452bar ( .A1(in_24bar), .A2(inbar[97]), .ZN(n523bar) );
  OR2_X1 U453 ( .A1(in_33), .A2(in_27), .ZN(n524) );
  AND2_X1 U453bar ( .A1(in_33bar), .A2(in_27bar), .ZN(n524bar) );
  OR2_X1 U454 ( .A1(n522), .A2(n521), .ZN(n568) );
  AND2_X1 U454bar ( .A1(n522bar), .A2(n521bar), .ZN(n568bar) );
  OR2_X1 U455 ( .A1(in[145]), .A2(in[126]), .ZN(n521) );
  AND2_X1 U455bar ( .A1(inbar[145]), .A2(inbar[126]), .ZN(n521bar) );
  OR2_X1 U456 ( .A1(in[169]), .A2(n520), .ZN(n522) );
  AND2_X1 U456bar ( .A1(inbar[169]), .A2(n520bar), .ZN(n522bar) );
  OR2_X1 U457 ( .A1(in[221]), .A2(in[172]), .ZN(n520) );
  AND2_X1 U457bar ( .A1(inbar[221]), .A2(inbar[172]), .ZN(n520bar) );
  OR2_X1 U458 ( .A1(n519), .A2(n518), .ZN(n570) );
  AND2_X1 U458bar ( .A1(n519bar), .A2(n518bar), .ZN(n570bar) );
  OR2_X1 U459 ( .A1(n517), .A2(n516), .ZN(n518) );
  AND2_X1 U459bar ( .A1(n517bar), .A2(n516bar), .ZN(n518bar) );
  OR2_X1 U460 ( .A1(in[241]), .A2(in[224]), .ZN(n516) );
  AND2_X1 U460bar ( .A1(inbar[241]), .A2(inbar[224]), .ZN(n516bar) );
  OR2_X1 U461 ( .A1(in[86]), .A2(n515), .ZN(n517) );
  AND2_X1 U461bar ( .A1(inbar[86]), .A2(n515bar), .ZN(n517bar) );
  OR2_X1 U462 ( .A1(in_43), .A2(in_34), .ZN(n515) );
  AND2_X1 U462bar ( .A1(in_43bar), .A2(in_34bar), .ZN(n515bar) );
  OR2_X1 U463 ( .A1(n514), .A2(n513), .ZN(n519) );
  AND2_X1 U463bar ( .A1(n514bar), .A2(n513bar), .ZN(n519bar) );
  OR2_X1 U464 ( .A1(in_65), .A2(in_51), .ZN(n513) );
  AND2_X1 U464bar ( .A1(in_65bar), .A2(in_51bar), .ZN(n513bar) );
  OR2_X1 U465 ( .A1(in_75), .A2(n512), .ZN(n514) );
  AND2_X1 U465bar ( .A1(in_75bar), .A2(n512bar), .ZN(n514bar) );
  OR2_X1 U466 ( .A1(in_81), .A2(in_77), .ZN(n512) );
  AND2_X1 U466bar ( .A1(in_81bar), .A2(in_77bar), .ZN(n512bar) );
  OR2_X1 U467 ( .A1(n511), .A2(n510), .ZN(n778) );
  AND2_X1 U467bar ( .A1(n511bar), .A2(n510bar), .ZN(n778bar) );
  OR2_X1 U468 ( .A1(n509), .A2(n508), .ZN(n510) );
  AND2_X1 U468bar ( .A1(n509bar), .A2(n508bar), .ZN(n510bar) );
  OR2_X1 U469 ( .A1(n507), .A2(n506), .ZN(n508) );
  AND2_X1 U469bar ( .A1(n507bar), .A2(n506bar), .ZN(n508bar) );
  OR2_X1 U470 ( .A1(in[107]), .A2(in[101]), .ZN(n506) );
  AND2_X1 U470bar ( .A1(inbar[107]), .A2(inbar[101]), .ZN(n506bar) );
  OR2_X1 U471 ( .A1(in[139]), .A2(in[132]), .ZN(n507) );
  AND2_X1 U471bar ( .A1(inbar[139]), .A2(inbar[132]), .ZN(n507bar) );
  OR2_X1 U472 ( .A1(n505), .A2(n504), .ZN(n509) );
  AND2_X1 U472bar ( .A1(n505bar), .A2(n504bar), .ZN(n509bar) );
  OR2_X1 U473 ( .A1(in[146]), .A2(in[141]), .ZN(n504) );
  AND2_X1 U473bar ( .A1(inbar[146]), .A2(inbar[141]), .ZN(n504bar) );
  OR2_X1 U474 ( .A1(in[203]), .A2(in[179]), .ZN(n505) );
  AND2_X1 U474bar ( .A1(inbar[203]), .A2(inbar[179]), .ZN(n505bar) );
  OR2_X1 U475 ( .A1(n503), .A2(n502), .ZN(n511) );
  AND2_X1 U475bar ( .A1(n503bar), .A2(n502bar), .ZN(n511bar) );
  OR2_X1 U476 ( .A1(n501), .A2(n500), .ZN(n502) );
  AND2_X1 U476bar ( .A1(n501bar), .A2(n500bar), .ZN(n502bar) );
  OR2_X1 U477 ( .A1(in[243]), .A2(in[222]), .ZN(n500) );
  AND2_X1 U477bar ( .A1(inbar[243]), .A2(inbar[222]), .ZN(n500bar) );
  OR2_X1 U478 ( .A1(in[251]), .A2(in[250]), .ZN(n501) );
  AND2_X1 U478bar ( .A1(inbar[251]), .A2(inbar[250]), .ZN(n501bar) );
  OR2_X1 U479 ( .A1(n499), .A2(n498), .ZN(n503) );
  AND2_X1 U479bar ( .A1(n499bar), .A2(n498bar), .ZN(n503bar) );
  OR2_X1 U480 ( .A1(in_37), .A2(in_19), .ZN(n498) );
  AND2_X1 U480bar ( .A1(in_37bar), .A2(in_19bar), .ZN(n498bar) );
  OR2_X1 U481 ( .A1(in_78), .A2(in_6), .ZN(n499) );
  AND2_X1 U481bar ( .A1(in_78bar), .A2(in_6bar), .ZN(n499bar) );
  OR2_X1 U482 ( .A1(n497), .A2(n496), .ZN(n603) );
  AND2_X1 U482bar ( .A1(n497bar), .A2(n496bar), .ZN(n603bar) );
  OR2_X1 U483 ( .A1(in[112]), .A2(in[102]), .ZN(n496) );
  AND2_X1 U483bar ( .A1(inbar[112]), .A2(inbar[102]), .ZN(n496bar) );
  OR2_X1 U484 ( .A1(in[123]), .A2(n495), .ZN(n497) );
  AND2_X1 U484bar ( .A1(inbar[123]), .A2(n495bar), .ZN(n497bar) );
  OR2_X1 U485 ( .A1(in[143]), .A2(in[130]), .ZN(n495) );
  AND2_X1 U485bar ( .A1(inbar[143]), .A2(inbar[130]), .ZN(n495bar) );
  OR2_X1 U486 ( .A1(n494), .A2(n493), .ZN(n605) );
  AND2_X1 U486bar ( .A1(n494bar), .A2(n493bar), .ZN(n605bar) );
  OR2_X1 U487 ( .A1(n492), .A2(n491), .ZN(n493) );
  AND2_X1 U487bar ( .A1(n492bar), .A2(n491bar), .ZN(n493bar) );
  OR2_X1 U488 ( .A1(in[216]), .A2(in[213]), .ZN(n491) );
  AND2_X1 U488bar ( .A1(inbar[216]), .A2(inbar[213]), .ZN(n491bar) );
  OR2_X1 U489 ( .A1(in[227]), .A2(n490), .ZN(n492) );
  AND2_X1 U489bar ( .A1(inbar[227]), .A2(n490bar), .ZN(n492bar) );
  OR2_X1 U490 ( .A1(in_0), .A2(in[248]), .ZN(n490) );
  AND2_X1 U490bar ( .A1(in_0bar), .A2(inbar[248]), .ZN(n490bar) );
  OR2_X1 U491 ( .A1(n489), .A2(n488), .ZN(n494) );
  AND2_X1 U491bar ( .A1(n489bar), .A2(n488bar), .ZN(n494bar) );
  OR2_X1 U492 ( .A1(in_46), .A2(in_44), .ZN(n488) );
  AND2_X1 U492bar ( .A1(in_46bar), .A2(in_44bar), .ZN(n488bar) );
  OR2_X1 U493 ( .A1(in_50), .A2(n487), .ZN(n489) );
  AND2_X1 U493bar ( .A1(in_50bar), .A2(n487bar), .ZN(n489bar) );
  OR2_X1 U494 ( .A1(in_9), .A2(in_80), .ZN(n487) );
  AND2_X1 U494bar ( .A1(in_9bar), .A2(in_80bar), .ZN(n487bar) );
endmodule

module sBox_12 ( in, inbar, out, outbar );

  input wire [7:0] in;
  input wire [7:0] inbar;
//input_done

  output wire [7:0] out;
  output wire [7:0] outbar;
//output_done

  wire [255:0] decodeOut;
  wire [255:0] decodeOutbar;
//wire_done

  decode_12 dec ( .in(in), .inbar(inbar), .out(decodeOut), .outbar(decodeOutbar) );
  encode_12 enc ( .in(decodeOut), .inbar(decodeOutbar), .out(out), .outbar(outbar) );
endmodule

module CD2_49 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD2_50( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD2_51 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD2_52 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD4_25 ( a, abar, b, bbar, y, ybar );

  input wire [3:0] a;
  input wire [3:0] b;
  input wire [3:0] abar;
  input wire [3:0] bbar;
//input_done

  output wire [15:0] y;
  output wire [15:0] ybar;
//output_done

//wire_done

  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]) );
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]) );
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]) );
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]) );
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]) );
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]) );
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]) );
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]) );
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]) );
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]) );
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]) );
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]) );
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]) );
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]) );
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]) );
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]) );
endmodule

module CD4_26 ( a, abar, b, bbar, y, ybar );

  input wire [3:0] a;
  input wire [3:0] b;
  input wire [3:0] abar;
  input wire [3:0] bbar;
//input_done

  output wire [15:0] y;
  output wire [15:0] ybar;
//output_done

//wire_done

  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]) );
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]) );
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]) );
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]) );
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]) );
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]) );
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]) );
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]) );
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]) );
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]) );
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]) );
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]) );
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]) );
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]) );
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]) );
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]) );
endmodule

module CD16_13 ( a, abar, b, bbar, y, ybar );

  input wire [15:0] a;
  input wire [15:0] b;
  input wire [15:0] abar;
  input wire [15:0] bbar;
//input_done

  output wire [255:0] y;
  output wire [255:0] ybar;
//output_done

//wire_done

  AND2_X1 U1 ( .A1(b[9]), .A2(a[0]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[9]), .A2(abar[0]), .ZN(ybar[9]) );
  AND2_X1 U2 ( .A1(b[3]), .A2(a[6]), .ZN(y[99]) );
  OR2_X1 U2bar ( .A1(bbar[3]), .A2(abar[6]), .ZN(ybar[99]) );
  AND2_X1 U3 ( .A1(b[2]), .A2(a[6]), .ZN(y[98]) );
  OR2_X1 U3bar ( .A1(bbar[2]), .A2(abar[6]), .ZN(ybar[98]) );
  AND2_X1 U4 ( .A1(b[1]), .A2(a[6]), .ZN(y[97]) );
  OR2_X1 U4bar ( .A1(bbar[1]), .A2(abar[6]), .ZN(ybar[97]) );
  AND2_X1 U5 ( .A1(b[0]), .A2(a[6]), .ZN(y[96]) );
  OR2_X1 U5bar ( .A1(bbar[0]), .A2(abar[6]), .ZN(ybar[96]) );
  AND2_X1 U6 ( .A1(b[15]), .A2(a[5]), .ZN(y[95]) );
  OR2_X1 U6bar ( .A1(bbar[15]), .A2(abar[5]), .ZN(ybar[95]) );
  AND2_X1 U7 ( .A1(b[14]), .A2(a[5]), .ZN(y[94]) );
  OR2_X1 U7bar ( .A1(bbar[14]), .A2(abar[5]), .ZN(ybar[94]) );
  AND2_X1 U8 ( .A1(b[13]), .A2(a[5]), .ZN(y[93]) );
  OR2_X1 U8bar ( .A1(bbar[13]), .A2(abar[5]), .ZN(ybar[93]) );
  AND2_X1 U9 ( .A1(b[12]), .A2(a[5]), .ZN(y[92]) );
  OR2_X1 U9bar ( .A1(bbar[12]), .A2(abar[5]), .ZN(ybar[92]) );
  AND2_X1 U10 ( .A1(b[11]), .A2(a[5]), .ZN(y[91]) );
  OR2_X1 U10bar ( .A1(bbar[11]), .A2(abar[5]), .ZN(ybar[91]) );
  AND2_X1 U11 ( .A1(b[10]), .A2(a[5]), .ZN(y[90]) );
  OR2_X1 U11bar ( .A1(bbar[10]), .A2(abar[5]), .ZN(ybar[90]) );
  AND2_X1 U12 ( .A1(b[8]), .A2(a[0]), .ZN(y[8]) );
  OR2_X1 U12bar ( .A1(bbar[8]), .A2(abar[0]), .ZN(ybar[8]) );
  AND2_X1 U13 ( .A1(a[5]), .A2(b[9]), .ZN(y[89]) );
  OR2_X1 U13bar ( .A1(abar[5]), .A2(bbar[9]), .ZN(ybar[89]) );
  AND2_X1 U14 ( .A1(b[8]), .A2(a[5]), .ZN(y[88]) );
  OR2_X1 U14bar ( .A1(bbar[8]), .A2(abar[5]), .ZN(ybar[88]) );
  AND2_X1 U15 ( .A1(b[7]), .A2(a[5]), .ZN(y[87]) );
  OR2_X1 U15bar ( .A1(bbar[7]), .A2(abar[5]), .ZN(ybar[87]) );
  AND2_X1 U16 ( .A1(b[6]), .A2(a[5]), .ZN(y[86]) );
  OR2_X1 U16bar ( .A1(bbar[6]), .A2(abar[5]), .ZN(ybar[86]) );
  AND2_X1 U17 ( .A1(b[5]), .A2(a[5]), .ZN(y[85]) );
  OR2_X1 U17bar ( .A1(bbar[5]), .A2(abar[5]), .ZN(ybar[85]) );
  AND2_X1 U18 ( .A1(b[4]), .A2(a[5]), .ZN(y[84]) );
  OR2_X1 U18bar ( .A1(bbar[4]), .A2(abar[5]), .ZN(ybar[84]) );
  AND2_X1 U19 ( .A1(a[5]), .A2(b[3]), .ZN(y[83]) );
  OR2_X1 U19bar ( .A1(abar[5]), .A2(bbar[3]), .ZN(ybar[83]) );
  AND2_X1 U20 ( .A1(a[5]), .A2(b[2]), .ZN(y[82]) );
  OR2_X1 U20bar ( .A1(abar[5]), .A2(bbar[2]), .ZN(ybar[82]) );
  AND2_X1 U21 ( .A1(a[5]), .A2(b[1]), .ZN(y[81]) );
  OR2_X1 U21bar ( .A1(abar[5]), .A2(bbar[1]), .ZN(ybar[81]) );
  AND2_X1 U22 ( .A1(a[5]), .A2(b[0]), .ZN(y[80]) );
  OR2_X1 U22bar ( .A1(abar[5]), .A2(bbar[0]), .ZN(ybar[80]) );
  AND2_X1 U23 ( .A1(b[7]), .A2(a[0]), .ZN(y[7]) );
  OR2_X1 U23bar ( .A1(bbar[7]), .A2(abar[0]), .ZN(ybar[7]) );
  AND2_X1 U24 ( .A1(a[4]), .A2(b[15]), .ZN(y[79]) );
  OR2_X1 U24bar ( .A1(abar[4]), .A2(bbar[15]), .ZN(ybar[79]) );
  AND2_X1 U25 ( .A1(a[4]), .A2(b[14]), .ZN(y[78]) );
  OR2_X1 U25bar ( .A1(abar[4]), .A2(bbar[14]), .ZN(ybar[78]) );
  AND2_X1 U26 ( .A1(a[4]), .A2(b[13]), .ZN(y[77]) );
  OR2_X1 U26bar ( .A1(abar[4]), .A2(bbar[13]), .ZN(ybar[77]) );
  AND2_X1 U27 ( .A1(a[4]), .A2(b[12]), .ZN(y[76]) );
  OR2_X1 U27bar ( .A1(abar[4]), .A2(bbar[12]), .ZN(ybar[76]) );
  AND2_X1 U28 ( .A1(a[4]), .A2(b[11]), .ZN(y[75]) );
  OR2_X1 U28bar ( .A1(abar[4]), .A2(bbar[11]), .ZN(ybar[75]) );
  AND2_X1 U29 ( .A1(a[4]), .A2(b[10]), .ZN(y[74]) );
  OR2_X1 U29bar ( .A1(abar[4]), .A2(bbar[10]), .ZN(ybar[74]) );
  AND2_X1 U30 ( .A1(a[4]), .A2(b[9]), .ZN(y[73]) );
  OR2_X1 U30bar ( .A1(abar[4]), .A2(bbar[9]), .ZN(ybar[73]) );
  AND2_X1 U31 ( .A1(a[4]), .A2(b[8]), .ZN(y[72]) );
  OR2_X1 U31bar ( .A1(abar[4]), .A2(bbar[8]), .ZN(ybar[72]) );
  AND2_X1 U32 ( .A1(a[4]), .A2(b[7]), .ZN(y[71]) );
  OR2_X1 U32bar ( .A1(abar[4]), .A2(bbar[7]), .ZN(ybar[71]) );
  AND2_X1 U33 ( .A1(a[4]), .A2(b[6]), .ZN(y[70]) );
  OR2_X1 U33bar ( .A1(abar[4]), .A2(bbar[6]), .ZN(ybar[70]) );
  AND2_X1 U34 ( .A1(b[6]), .A2(a[0]), .ZN(y[6]) );
  OR2_X1 U34bar ( .A1(bbar[6]), .A2(abar[0]), .ZN(ybar[6]) );
  AND2_X1 U35 ( .A1(a[4]), .A2(b[5]), .ZN(y[69]) );
  OR2_X1 U35bar ( .A1(abar[4]), .A2(bbar[5]), .ZN(ybar[69]) );
  AND2_X1 U36 ( .A1(a[4]), .A2(b[4]), .ZN(y[68]) );
  OR2_X1 U36bar ( .A1(abar[4]), .A2(bbar[4]), .ZN(ybar[68]) );
  AND2_X1 U37 ( .A1(a[4]), .A2(b[3]), .ZN(y[67]) );
  OR2_X1 U37bar ( .A1(abar[4]), .A2(bbar[3]), .ZN(ybar[67]) );
  AND2_X1 U38 ( .A1(a[4]), .A2(b[2]), .ZN(y[66]) );
  OR2_X1 U38bar ( .A1(abar[4]), .A2(bbar[2]), .ZN(ybar[66]) );
  AND2_X1 U39 ( .A1(a[4]), .A2(b[1]), .ZN(y[65]) );
  OR2_X1 U39bar ( .A1(abar[4]), .A2(bbar[1]), .ZN(ybar[65]) );
  AND2_X1 U40 ( .A1(a[4]), .A2(b[0]), .ZN(y[64]) );
  OR2_X1 U40bar ( .A1(abar[4]), .A2(bbar[0]), .ZN(ybar[64]) );
  AND2_X1 U41 ( .A1(a[3]), .A2(b[15]), .ZN(y[63]) );
  OR2_X1 U41bar ( .A1(abar[3]), .A2(bbar[15]), .ZN(ybar[63]) );
  AND2_X1 U42 ( .A1(a[3]), .A2(b[14]), .ZN(y[62]) );
  OR2_X1 U42bar ( .A1(abar[3]), .A2(bbar[14]), .ZN(ybar[62]) );
  AND2_X1 U43 ( .A1(a[3]), .A2(b[13]), .ZN(y[61]) );
  OR2_X1 U43bar ( .A1(abar[3]), .A2(bbar[13]), .ZN(ybar[61]) );
  AND2_X1 U44 ( .A1(a[3]), .A2(b[12]), .ZN(y[60]) );
  OR2_X1 U44bar ( .A1(abar[3]), .A2(bbar[12]), .ZN(ybar[60]) );
  AND2_X1 U45 ( .A1(b[5]), .A2(a[0]), .ZN(y[5]) );
  OR2_X1 U45bar ( .A1(bbar[5]), .A2(abar[0]), .ZN(ybar[5]) );
  AND2_X1 U46 ( .A1(a[3]), .A2(b[11]), .ZN(y[59]) );
  OR2_X1 U46bar ( .A1(abar[3]), .A2(bbar[11]), .ZN(ybar[59]) );
  AND2_X1 U47 ( .A1(a[3]), .A2(b[10]), .ZN(y[58]) );
  OR2_X1 U47bar ( .A1(abar[3]), .A2(bbar[10]), .ZN(ybar[58]) );
  AND2_X1 U48 ( .A1(a[3]), .A2(b[9]), .ZN(y[57]) );
  OR2_X1 U48bar ( .A1(abar[3]), .A2(bbar[9]), .ZN(ybar[57]) );
  AND2_X1 U49 ( .A1(a[3]), .A2(b[8]), .ZN(y[56]) );
  OR2_X1 U49bar ( .A1(abar[3]), .A2(bbar[8]), .ZN(ybar[56]) );
  AND2_X1 U50 ( .A1(a[3]), .A2(b[7]), .ZN(y[55]) );
  OR2_X1 U50bar ( .A1(abar[3]), .A2(bbar[7]), .ZN(ybar[55]) );
  AND2_X1 U51 ( .A1(a[3]), .A2(b[6]), .ZN(y[54]) );
  OR2_X1 U51bar ( .A1(abar[3]), .A2(bbar[6]), .ZN(ybar[54]) );
  AND2_X1 U52 ( .A1(a[3]), .A2(b[5]), .ZN(y[53]) );
  OR2_X1 U52bar ( .A1(abar[3]), .A2(bbar[5]), .ZN(ybar[53]) );
  AND2_X1 U53 ( .A1(a[3]), .A2(b[4]), .ZN(y[52]) );
  OR2_X1 U53bar ( .A1(abar[3]), .A2(bbar[4]), .ZN(ybar[52]) );
  AND2_X1 U54 ( .A1(a[3]), .A2(b[3]), .ZN(y[51]) );
  OR2_X1 U54bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[51]) );
  AND2_X1 U55 ( .A1(a[3]), .A2(b[2]), .ZN(y[50]) );
  OR2_X1 U55bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[50]) );
  AND2_X1 U56 ( .A1(b[4]), .A2(a[0]), .ZN(y[4]) );
  OR2_X1 U56bar ( .A1(bbar[4]), .A2(abar[0]), .ZN(ybar[4]) );
  AND2_X1 U57 ( .A1(a[3]), .A2(b[1]), .ZN(y[49]) );
  OR2_X1 U57bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[49]) );
  AND2_X1 U58 ( .A1(a[3]), .A2(b[0]), .ZN(y[48]) );
  OR2_X1 U58bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[48]) );
  AND2_X1 U59 ( .A1(a[2]), .A2(b[15]), .ZN(y[47]) );
  OR2_X1 U59bar ( .A1(abar[2]), .A2(bbar[15]), .ZN(ybar[47]) );
  AND2_X1 U60 ( .A1(a[2]), .A2(b[14]), .ZN(y[46]) );
  OR2_X1 U60bar ( .A1(abar[2]), .A2(bbar[14]), .ZN(ybar[46]) );
  AND2_X1 U61 ( .A1(a[2]), .A2(b[13]), .ZN(y[45]) );
  OR2_X1 U61bar ( .A1(abar[2]), .A2(bbar[13]), .ZN(ybar[45]) );
  AND2_X1 U62 ( .A1(a[2]), .A2(b[12]), .ZN(y[44]) );
  OR2_X1 U62bar ( .A1(abar[2]), .A2(bbar[12]), .ZN(ybar[44]) );
  AND2_X1 U63 ( .A1(a[2]), .A2(b[11]), .ZN(y[43]) );
  OR2_X1 U63bar ( .A1(abar[2]), .A2(bbar[11]), .ZN(ybar[43]) );
  AND2_X1 U64 ( .A1(a[2]), .A2(b[10]), .ZN(y[42]) );
  OR2_X1 U64bar ( .A1(abar[2]), .A2(bbar[10]), .ZN(ybar[42]) );
  AND2_X1 U65 ( .A1(a[2]), .A2(b[9]), .ZN(y[41]) );
  OR2_X1 U65bar ( .A1(abar[2]), .A2(bbar[9]), .ZN(ybar[41]) );
  AND2_X1 U66 ( .A1(a[2]), .A2(b[8]), .ZN(y[40]) );
  OR2_X1 U66bar ( .A1(abar[2]), .A2(bbar[8]), .ZN(ybar[40]) );
  AND2_X1 U67 ( .A1(b[3]), .A2(a[0]), .ZN(y[3]) );
  OR2_X1 U67bar ( .A1(bbar[3]), .A2(abar[0]), .ZN(ybar[3]) );
  AND2_X1 U68 ( .A1(a[2]), .A2(b[7]), .ZN(y[39]) );
  OR2_X1 U68bar ( .A1(abar[2]), .A2(bbar[7]), .ZN(ybar[39]) );
  AND2_X1 U69 ( .A1(a[2]), .A2(b[6]), .ZN(y[38]) );
  OR2_X1 U69bar ( .A1(abar[2]), .A2(bbar[6]), .ZN(ybar[38]) );
  AND2_X1 U70 ( .A1(a[2]), .A2(b[5]), .ZN(y[37]) );
  OR2_X1 U70bar ( .A1(abar[2]), .A2(bbar[5]), .ZN(ybar[37]) );
  AND2_X1 U71 ( .A1(a[2]), .A2(b[4]), .ZN(y[36]) );
  OR2_X1 U71bar ( .A1(abar[2]), .A2(bbar[4]), .ZN(ybar[36]) );
  AND2_X1 U72 ( .A1(a[2]), .A2(b[3]), .ZN(y[35]) );
  OR2_X1 U72bar ( .A1(abar[2]), .A2(bbar[3]), .ZN(ybar[35]) );
  AND2_X1 U73 ( .A1(a[2]), .A2(b[2]), .ZN(y[34]) );
  OR2_X1 U73bar ( .A1(abar[2]), .A2(bbar[2]), .ZN(ybar[34]) );
  AND2_X1 U74 ( .A1(a[2]), .A2(b[1]), .ZN(y[33]) );
  OR2_X1 U74bar ( .A1(abar[2]), .A2(bbar[1]), .ZN(ybar[33]) );
  AND2_X1 U75 ( .A1(a[2]), .A2(b[0]), .ZN(y[32]) );
  OR2_X1 U75bar ( .A1(abar[2]), .A2(bbar[0]), .ZN(ybar[32]) );
  AND2_X1 U76 ( .A1(a[1]), .A2(b[15]), .ZN(y[31]) );
  OR2_X1 U76bar ( .A1(abar[1]), .A2(bbar[15]), .ZN(ybar[31]) );
  AND2_X1 U77 ( .A1(a[1]), .A2(b[14]), .ZN(y[30]) );
  OR2_X1 U77bar ( .A1(abar[1]), .A2(bbar[14]), .ZN(ybar[30]) );
  AND2_X1 U78 ( .A1(b[2]), .A2(a[0]), .ZN(y[2]) );
  OR2_X1 U78bar ( .A1(bbar[2]), .A2(abar[0]), .ZN(ybar[2]) );
  AND2_X1 U79 ( .A1(a[1]), .A2(b[13]), .ZN(y[29]) );
  OR2_X1 U79bar ( .A1(abar[1]), .A2(bbar[13]), .ZN(ybar[29]) );
  AND2_X1 U80 ( .A1(a[1]), .A2(b[12]), .ZN(y[28]) );
  OR2_X1 U80bar ( .A1(abar[1]), .A2(bbar[12]), .ZN(ybar[28]) );
  AND2_X1 U81 ( .A1(a[1]), .A2(b[11]), .ZN(y[27]) );
  OR2_X1 U81bar ( .A1(abar[1]), .A2(bbar[11]), .ZN(ybar[27]) );
  AND2_X1 U82 ( .A1(a[1]), .A2(b[10]), .ZN(y[26]) );
  OR2_X1 U82bar ( .A1(abar[1]), .A2(bbar[10]), .ZN(ybar[26]) );
  AND2_X1 U83 ( .A1(a[1]), .A2(b[9]), .ZN(y[25]) );
  OR2_X1 U83bar ( .A1(abar[1]), .A2(bbar[9]), .ZN(ybar[25]) );
  AND2_X1 U84 ( .A1(a[15]), .A2(b[15]), .ZN(y[255]) );
  OR2_X1 U84bar ( .A1(abar[15]), .A2(bbar[15]), .ZN(ybar[255]) );
  AND2_X1 U85 ( .A1(a[15]), .A2(b[14]), .ZN(y[254]) );
  OR2_X1 U85bar ( .A1(abar[15]), .A2(bbar[14]), .ZN(ybar[254]) );
  AND2_X1 U86 ( .A1(a[15]), .A2(b[13]), .ZN(y[253]) );
  OR2_X1 U86bar ( .A1(abar[15]), .A2(bbar[13]), .ZN(ybar[253]) );
  AND2_X1 U87 ( .A1(a[15]), .A2(b[12]), .ZN(y[252]) );
  OR2_X1 U87bar ( .A1(abar[15]), .A2(bbar[12]), .ZN(ybar[252]) );
  AND2_X1 U88 ( .A1(a[15]), .A2(b[11]), .ZN(y[251]) );
  OR2_X1 U88bar ( .A1(abar[15]), .A2(bbar[11]), .ZN(ybar[251]) );
  AND2_X1 U89 ( .A1(a[15]), .A2(b[10]), .ZN(y[250]) );
  OR2_X1 U89bar ( .A1(abar[15]), .A2(bbar[10]), .ZN(ybar[250]) );
  AND2_X1 U90 ( .A1(a[1]), .A2(b[8]), .ZN(y[24]) );
  OR2_X1 U90bar ( .A1(abar[1]), .A2(bbar[8]), .ZN(ybar[24]) );
  AND2_X1 U91 ( .A1(a[15]), .A2(b[9]), .ZN(y[249]) );
  OR2_X1 U91bar ( .A1(abar[15]), .A2(bbar[9]), .ZN(ybar[249]) );
  AND2_X1 U92 ( .A1(a[15]), .A2(b[8]), .ZN(y[248]) );
  OR2_X1 U92bar ( .A1(abar[15]), .A2(bbar[8]), .ZN(ybar[248]) );
  AND2_X1 U93 ( .A1(a[15]), .A2(b[7]), .ZN(y[247]) );
  OR2_X1 U93bar ( .A1(abar[15]), .A2(bbar[7]), .ZN(ybar[247]) );
  AND2_X1 U94 ( .A1(a[15]), .A2(b[6]), .ZN(y[246]) );
  OR2_X1 U94bar ( .A1(abar[15]), .A2(bbar[6]), .ZN(ybar[246]) );
  AND2_X1 U95 ( .A1(a[15]), .A2(b[5]), .ZN(y[245]) );
  OR2_X1 U95bar ( .A1(abar[15]), .A2(bbar[5]), .ZN(ybar[245]) );
  AND2_X1 U96 ( .A1(a[15]), .A2(b[4]), .ZN(y[244]) );
  OR2_X1 U96bar ( .A1(abar[15]), .A2(bbar[4]), .ZN(ybar[244]) );
  AND2_X1 U97 ( .A1(a[15]), .A2(b[3]), .ZN(y[243]) );
  OR2_X1 U97bar ( .A1(abar[15]), .A2(bbar[3]), .ZN(ybar[243]) );
  AND2_X1 U98 ( .A1(a[15]), .A2(b[2]), .ZN(y[242]) );
  OR2_X1 U98bar ( .A1(abar[15]), .A2(bbar[2]), .ZN(ybar[242]) );
  AND2_X1 U99 ( .A1(a[15]), .A2(b[1]), .ZN(y[241]) );
  OR2_X1 U99bar ( .A1(abar[15]), .A2(bbar[1]), .ZN(ybar[241]) );
  AND2_X1 U100 ( .A1(a[15]), .A2(b[0]), .ZN(y[240]) );
  OR2_X1 U100bar ( .A1(abar[15]), .A2(bbar[0]), .ZN(ybar[240]) );
  AND2_X1 U101 ( .A1(a[1]), .A2(b[7]), .ZN(y[23]) );
  OR2_X1 U101bar ( .A1(abar[1]), .A2(bbar[7]), .ZN(ybar[23]) );
  AND2_X1 U102 ( .A1(a[14]), .A2(b[15]), .ZN(y[239]) );
  OR2_X1 U102bar ( .A1(abar[14]), .A2(bbar[15]), .ZN(ybar[239]) );
  AND2_X1 U103 ( .A1(a[14]), .A2(b[14]), .ZN(y[238]) );
  OR2_X1 U103bar ( .A1(abar[14]), .A2(bbar[14]), .ZN(ybar[238]) );
  AND2_X1 U104 ( .A1(a[14]), .A2(b[13]), .ZN(y[237]) );
  OR2_X1 U104bar ( .A1(abar[14]), .A2(bbar[13]), .ZN(ybar[237]) );
  AND2_X1 U105 ( .A1(a[14]), .A2(b[12]), .ZN(y[236]) );
  OR2_X1 U105bar ( .A1(abar[14]), .A2(bbar[12]), .ZN(ybar[236]) );
  AND2_X1 U106 ( .A1(a[14]), .A2(b[11]), .ZN(y[235]) );
  OR2_X1 U106bar ( .A1(abar[14]), .A2(bbar[11]), .ZN(ybar[235]) );
  AND2_X1 U107 ( .A1(a[14]), .A2(b[10]), .ZN(y[234]) );
  OR2_X1 U107bar ( .A1(abar[14]), .A2(bbar[10]), .ZN(ybar[234]) );
  AND2_X1 U108 ( .A1(a[14]), .A2(b[9]), .ZN(y[233]) );
  OR2_X1 U108bar ( .A1(abar[14]), .A2(bbar[9]), .ZN(ybar[233]) );
  AND2_X1 U109 ( .A1(a[14]), .A2(b[8]), .ZN(y[232]) );
  OR2_X1 U109bar ( .A1(abar[14]), .A2(bbar[8]), .ZN(ybar[232]) );
  AND2_X1 U110 ( .A1(a[14]), .A2(b[7]), .ZN(y[231]) );
  OR2_X1 U110bar ( .A1(abar[14]), .A2(bbar[7]), .ZN(ybar[231]) );
  AND2_X1 U111 ( .A1(a[14]), .A2(b[6]), .ZN(y[230]) );
  OR2_X1 U111bar ( .A1(abar[14]), .A2(bbar[6]), .ZN(ybar[230]) );
  AND2_X1 U112 ( .A1(a[1]), .A2(b[6]), .ZN(y[22]) );
  OR2_X1 U112bar ( .A1(abar[1]), .A2(bbar[6]), .ZN(ybar[22]) );
  AND2_X1 U113 ( .A1(a[14]), .A2(b[5]), .ZN(y[229]) );
  OR2_X1 U113bar ( .A1(abar[14]), .A2(bbar[5]), .ZN(ybar[229]) );
  AND2_X1 U114 ( .A1(a[14]), .A2(b[4]), .ZN(y[228]) );
  OR2_X1 U114bar ( .A1(abar[14]), .A2(bbar[4]), .ZN(ybar[228]) );
  AND2_X1 U115 ( .A1(a[14]), .A2(b[3]), .ZN(y[227]) );
  OR2_X1 U115bar ( .A1(abar[14]), .A2(bbar[3]), .ZN(ybar[227]) );
  AND2_X1 U116 ( .A1(a[14]), .A2(b[2]), .ZN(y[226]) );
  OR2_X1 U116bar ( .A1(abar[14]), .A2(bbar[2]), .ZN(ybar[226]) );
  AND2_X1 U117 ( .A1(a[14]), .A2(b[1]), .ZN(y[225]) );
  OR2_X1 U117bar ( .A1(abar[14]), .A2(bbar[1]), .ZN(ybar[225]) );
  AND2_X1 U118 ( .A1(a[14]), .A2(b[0]), .ZN(y[224]) );
  OR2_X1 U118bar ( .A1(abar[14]), .A2(bbar[0]), .ZN(ybar[224]) );
  AND2_X1 U119 ( .A1(a[13]), .A2(b[15]), .ZN(y[223]) );
  OR2_X1 U119bar ( .A1(abar[13]), .A2(bbar[15]), .ZN(ybar[223]) );
  AND2_X1 U120 ( .A1(a[13]), .A2(b[14]), .ZN(y[222]) );
  OR2_X1 U120bar ( .A1(abar[13]), .A2(bbar[14]), .ZN(ybar[222]) );
  AND2_X1 U121 ( .A1(a[13]), .A2(b[13]), .ZN(y[221]) );
  OR2_X1 U121bar ( .A1(abar[13]), .A2(bbar[13]), .ZN(ybar[221]) );
  AND2_X1 U122 ( .A1(a[13]), .A2(b[12]), .ZN(y[220]) );
  OR2_X1 U122bar ( .A1(abar[13]), .A2(bbar[12]), .ZN(ybar[220]) );
  AND2_X1 U123 ( .A1(a[1]), .A2(b[5]), .ZN(y[21]) );
  OR2_X1 U123bar ( .A1(abar[1]), .A2(bbar[5]), .ZN(ybar[21]) );
  AND2_X1 U124 ( .A1(a[13]), .A2(b[11]), .ZN(y[219]) );
  OR2_X1 U124bar ( .A1(abar[13]), .A2(bbar[11]), .ZN(ybar[219]) );
  AND2_X1 U125 ( .A1(a[13]), .A2(b[10]), .ZN(y[218]) );
  OR2_X1 U125bar ( .A1(abar[13]), .A2(bbar[10]), .ZN(ybar[218]) );
  AND2_X1 U126 ( .A1(a[13]), .A2(b[9]), .ZN(y[217]) );
  OR2_X1 U126bar ( .A1(abar[13]), .A2(bbar[9]), .ZN(ybar[217]) );
  AND2_X1 U127 ( .A1(a[13]), .A2(b[8]), .ZN(y[216]) );
  OR2_X1 U127bar ( .A1(abar[13]), .A2(bbar[8]), .ZN(ybar[216]) );
  AND2_X1 U128 ( .A1(a[13]), .A2(b[7]), .ZN(y[215]) );
  OR2_X1 U128bar ( .A1(abar[13]), .A2(bbar[7]), .ZN(ybar[215]) );
  AND2_X1 U129 ( .A1(a[13]), .A2(b[6]), .ZN(y[214]) );
  OR2_X1 U129bar ( .A1(abar[13]), .A2(bbar[6]), .ZN(ybar[214]) );
  AND2_X1 U130 ( .A1(a[13]), .A2(b[5]), .ZN(y[213]) );
  OR2_X1 U130bar ( .A1(abar[13]), .A2(bbar[5]), .ZN(ybar[213]) );
  AND2_X1 U131 ( .A1(a[13]), .A2(b[4]), .ZN(y[212]) );
  OR2_X1 U131bar ( .A1(abar[13]), .A2(bbar[4]), .ZN(ybar[212]) );
  AND2_X1 U132 ( .A1(a[13]), .A2(b[3]), .ZN(y[211]) );
  OR2_X1 U132bar ( .A1(abar[13]), .A2(bbar[3]), .ZN(ybar[211]) );
  AND2_X1 U133 ( .A1(a[13]), .A2(b[2]), .ZN(y[210]) );
  OR2_X1 U133bar ( .A1(abar[13]), .A2(bbar[2]), .ZN(ybar[210]) );
  AND2_X1 U134 ( .A1(a[1]), .A2(b[4]), .ZN(y[20]) );
  OR2_X1 U134bar ( .A1(abar[1]), .A2(bbar[4]), .ZN(ybar[20]) );
  AND2_X1 U135 ( .A1(a[13]), .A2(b[1]), .ZN(y[209]) );
  OR2_X1 U135bar ( .A1(abar[13]), .A2(bbar[1]), .ZN(ybar[209]) );
  AND2_X1 U136 ( .A1(a[13]), .A2(b[0]), .ZN(y[208]) );
  OR2_X1 U136bar ( .A1(abar[13]), .A2(bbar[0]), .ZN(ybar[208]) );
  AND2_X1 U137 ( .A1(a[12]), .A2(b[15]), .ZN(y[207]) );
  OR2_X1 U137bar ( .A1(abar[12]), .A2(bbar[15]), .ZN(ybar[207]) );
  AND2_X1 U138 ( .A1(a[12]), .A2(b[14]), .ZN(y[206]) );
  OR2_X1 U138bar ( .A1(abar[12]), .A2(bbar[14]), .ZN(ybar[206]) );
  AND2_X1 U139 ( .A1(a[12]), .A2(b[13]), .ZN(y[205]) );
  OR2_X1 U139bar ( .A1(abar[12]), .A2(bbar[13]), .ZN(ybar[205]) );
  AND2_X1 U140 ( .A1(a[12]), .A2(b[12]), .ZN(y[204]) );
  OR2_X1 U140bar ( .A1(abar[12]), .A2(bbar[12]), .ZN(ybar[204]) );
  AND2_X1 U141 ( .A1(a[12]), .A2(b[11]), .ZN(y[203]) );
  OR2_X1 U141bar ( .A1(abar[12]), .A2(bbar[11]), .ZN(ybar[203]) );
  AND2_X1 U142 ( .A1(a[12]), .A2(b[10]), .ZN(y[202]) );
  OR2_X1 U142bar ( .A1(abar[12]), .A2(bbar[10]), .ZN(ybar[202]) );
  AND2_X1 U143 ( .A1(a[12]), .A2(b[9]), .ZN(y[201]) );
  OR2_X1 U143bar ( .A1(abar[12]), .A2(bbar[9]), .ZN(ybar[201]) );
  AND2_X1 U144 ( .A1(a[12]), .A2(b[8]), .ZN(y[200]) );
  OR2_X1 U144bar ( .A1(abar[12]), .A2(bbar[8]), .ZN(ybar[200]) );
  AND2_X1 U145 ( .A1(b[1]), .A2(a[0]), .ZN(y[1]) );
  OR2_X1 U145bar ( .A1(bbar[1]), .A2(abar[0]), .ZN(ybar[1]) );
  AND2_X1 U146 ( .A1(a[1]), .A2(b[3]), .ZN(y[19]) );
  OR2_X1 U146bar ( .A1(abar[1]), .A2(bbar[3]), .ZN(ybar[19]) );
  AND2_X1 U147 ( .A1(a[12]), .A2(b[7]), .ZN(y[199]) );
  OR2_X1 U147bar ( .A1(abar[12]), .A2(bbar[7]), .ZN(ybar[199]) );
  AND2_X1 U148 ( .A1(a[12]), .A2(b[6]), .ZN(y[198]) );
  OR2_X1 U148bar ( .A1(abar[12]), .A2(bbar[6]), .ZN(ybar[198]) );
  AND2_X1 U149 ( .A1(a[12]), .A2(b[5]), .ZN(y[197]) );
  OR2_X1 U149bar ( .A1(abar[12]), .A2(bbar[5]), .ZN(ybar[197]) );
  AND2_X1 U150 ( .A1(a[12]), .A2(b[4]), .ZN(y[196]) );
  OR2_X1 U150bar ( .A1(abar[12]), .A2(bbar[4]), .ZN(ybar[196]) );
  AND2_X1 U151 ( .A1(a[12]), .A2(b[3]), .ZN(y[195]) );
  OR2_X1 U151bar ( .A1(abar[12]), .A2(bbar[3]), .ZN(ybar[195]) );
  AND2_X1 U152 ( .A1(a[12]), .A2(b[2]), .ZN(y[194]) );
  OR2_X1 U152bar ( .A1(abar[12]), .A2(bbar[2]), .ZN(ybar[194]) );
  AND2_X1 U153 ( .A1(a[12]), .A2(b[1]), .ZN(y[193]) );
  OR2_X1 U153bar ( .A1(abar[12]), .A2(bbar[1]), .ZN(ybar[193]) );
  AND2_X1 U154 ( .A1(a[12]), .A2(b[0]), .ZN(y[192]) );
  OR2_X1 U154bar ( .A1(abar[12]), .A2(bbar[0]), .ZN(ybar[192]) );
  AND2_X1 U155 ( .A1(a[11]), .A2(b[15]), .ZN(y[191]) );
  OR2_X1 U155bar ( .A1(abar[11]), .A2(bbar[15]), .ZN(ybar[191]) );
  AND2_X1 U156 ( .A1(a[11]), .A2(b[14]), .ZN(y[190]) );
  OR2_X1 U156bar ( .A1(abar[11]), .A2(bbar[14]), .ZN(ybar[190]) );
  AND2_X1 U157 ( .A1(a[1]), .A2(b[2]), .ZN(y[18]) );
  OR2_X1 U157bar ( .A1(abar[1]), .A2(bbar[2]), .ZN(ybar[18]) );
  AND2_X1 U158 ( .A1(a[11]), .A2(b[13]), .ZN(y[189]) );
  OR2_X1 U158bar ( .A1(abar[11]), .A2(bbar[13]), .ZN(ybar[189]) );
  AND2_X1 U159 ( .A1(a[11]), .A2(b[12]), .ZN(y[188]) );
  OR2_X1 U159bar ( .A1(abar[11]), .A2(bbar[12]), .ZN(ybar[188]) );
  AND2_X1 U160 ( .A1(a[11]), .A2(b[11]), .ZN(y[187]) );
  OR2_X1 U160bar ( .A1(abar[11]), .A2(bbar[11]), .ZN(ybar[187]) );
  AND2_X1 U161 ( .A1(a[11]), .A2(b[10]), .ZN(y[186]) );
  OR2_X1 U161bar ( .A1(abar[11]), .A2(bbar[10]), .ZN(ybar[186]) );
  AND2_X1 U162 ( .A1(a[11]), .A2(b[9]), .ZN(y[185]) );
  OR2_X1 U162bar ( .A1(abar[11]), .A2(bbar[9]), .ZN(ybar[185]) );
  AND2_X1 U163 ( .A1(a[11]), .A2(b[8]), .ZN(y[184]) );
  OR2_X1 U163bar ( .A1(abar[11]), .A2(bbar[8]), .ZN(ybar[184]) );
  AND2_X1 U164 ( .A1(a[11]), .A2(b[7]), .ZN(y[183]) );
  OR2_X1 U164bar ( .A1(abar[11]), .A2(bbar[7]), .ZN(ybar[183]) );
  AND2_X1 U165 ( .A1(a[11]), .A2(b[6]), .ZN(y[182]) );
  OR2_X1 U165bar ( .A1(abar[11]), .A2(bbar[6]), .ZN(ybar[182]) );
  AND2_X1 U166 ( .A1(a[11]), .A2(b[5]), .ZN(y[181]) );
  OR2_X1 U166bar ( .A1(abar[11]), .A2(bbar[5]), .ZN(ybar[181]) );
  AND2_X1 U167 ( .A1(a[11]), .A2(b[4]), .ZN(y[180]) );
  OR2_X1 U167bar ( .A1(abar[11]), .A2(bbar[4]), .ZN(ybar[180]) );
  AND2_X1 U168 ( .A1(a[1]), .A2(b[1]), .ZN(y[17]) );
  OR2_X1 U168bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[17]) );
  AND2_X1 U169 ( .A1(a[11]), .A2(b[3]), .ZN(y[179]) );
  OR2_X1 U169bar ( .A1(abar[11]), .A2(bbar[3]), .ZN(ybar[179]) );
  AND2_X1 U170 ( .A1(a[11]), .A2(b[2]), .ZN(y[178]) );
  OR2_X1 U170bar ( .A1(abar[11]), .A2(bbar[2]), .ZN(ybar[178]) );
  AND2_X1 U171 ( .A1(a[11]), .A2(b[1]), .ZN(y[177]) );
  OR2_X1 U171bar ( .A1(abar[11]), .A2(bbar[1]), .ZN(ybar[177]) );
  AND2_X1 U172 ( .A1(a[11]), .A2(b[0]), .ZN(y[176]) );
  OR2_X1 U172bar ( .A1(abar[11]), .A2(bbar[0]), .ZN(ybar[176]) );
  AND2_X1 U173 ( .A1(a[10]), .A2(b[15]), .ZN(y[175]) );
  OR2_X1 U173bar ( .A1(abar[10]), .A2(bbar[15]), .ZN(ybar[175]) );
  AND2_X1 U174 ( .A1(a[10]), .A2(b[14]), .ZN(y[174]) );
  OR2_X1 U174bar ( .A1(abar[10]), .A2(bbar[14]), .ZN(ybar[174]) );
  AND2_X1 U175 ( .A1(a[10]), .A2(b[13]), .ZN(y[173]) );
  OR2_X1 U175bar ( .A1(abar[10]), .A2(bbar[13]), .ZN(ybar[173]) );
  AND2_X1 U176 ( .A1(a[10]), .A2(b[12]), .ZN(y[172]) );
  OR2_X1 U176bar ( .A1(abar[10]), .A2(bbar[12]), .ZN(ybar[172]) );
  AND2_X1 U177 ( .A1(a[10]), .A2(b[11]), .ZN(y[171]) );
  OR2_X1 U177bar ( .A1(abar[10]), .A2(bbar[11]), .ZN(ybar[171]) );
  AND2_X1 U178 ( .A1(a[10]), .A2(b[10]), .ZN(y[170]) );
  OR2_X1 U178bar ( .A1(abar[10]), .A2(bbar[10]), .ZN(ybar[170]) );
  AND2_X1 U179 ( .A1(a[1]), .A2(b[0]), .ZN(y[16]) );
  OR2_X1 U179bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[16]) );
  AND2_X1 U180 ( .A1(a[10]), .A2(b[9]), .ZN(y[169]) );
  OR2_X1 U180bar ( .A1(abar[10]), .A2(bbar[9]), .ZN(ybar[169]) );
  AND2_X1 U181 ( .A1(a[10]), .A2(b[8]), .ZN(y[168]) );
  OR2_X1 U181bar ( .A1(abar[10]), .A2(bbar[8]), .ZN(ybar[168]) );
  AND2_X1 U182 ( .A1(a[10]), .A2(b[7]), .ZN(y[167]) );
  OR2_X1 U182bar ( .A1(abar[10]), .A2(bbar[7]), .ZN(ybar[167]) );
  AND2_X1 U183 ( .A1(a[10]), .A2(b[6]), .ZN(y[166]) );
  OR2_X1 U183bar ( .A1(abar[10]), .A2(bbar[6]), .ZN(ybar[166]) );
  AND2_X1 U184 ( .A1(a[10]), .A2(b[5]), .ZN(y[165]) );
  OR2_X1 U184bar ( .A1(abar[10]), .A2(bbar[5]), .ZN(ybar[165]) );
  AND2_X1 U185 ( .A1(a[10]), .A2(b[4]), .ZN(y[164]) );
  OR2_X1 U185bar ( .A1(abar[10]), .A2(bbar[4]), .ZN(ybar[164]) );
  AND2_X1 U186 ( .A1(a[10]), .A2(b[3]), .ZN(y[163]) );
  OR2_X1 U186bar ( .A1(abar[10]), .A2(bbar[3]), .ZN(ybar[163]) );
  AND2_X1 U187 ( .A1(a[10]), .A2(b[2]), .ZN(y[162]) );
  OR2_X1 U187bar ( .A1(abar[10]), .A2(bbar[2]), .ZN(ybar[162]) );
  AND2_X1 U188 ( .A1(a[10]), .A2(b[1]), .ZN(y[161]) );
  OR2_X1 U188bar ( .A1(abar[10]), .A2(bbar[1]), .ZN(ybar[161]) );
  AND2_X1 U189 ( .A1(a[10]), .A2(b[0]), .ZN(y[160]) );
  OR2_X1 U189bar ( .A1(abar[10]), .A2(bbar[0]), .ZN(ybar[160]) );
  AND2_X1 U190 ( .A1(b[15]), .A2(a[0]), .ZN(y[15]) );
  OR2_X1 U190bar ( .A1(bbar[15]), .A2(abar[0]), .ZN(ybar[15]) );
  AND2_X1 U191 ( .A1(a[9]), .A2(b[15]), .ZN(y[159]) );
  OR2_X1 U191bar ( .A1(abar[9]), .A2(bbar[15]), .ZN(ybar[159]) );
  AND2_X1 U192 ( .A1(a[9]), .A2(b[14]), .ZN(y[158]) );
  OR2_X1 U192bar ( .A1(abar[9]), .A2(bbar[14]), .ZN(ybar[158]) );
  AND2_X1 U193 ( .A1(a[9]), .A2(b[13]), .ZN(y[157]) );
  OR2_X1 U193bar ( .A1(abar[9]), .A2(bbar[13]), .ZN(ybar[157]) );
  AND2_X1 U194 ( .A1(a[9]), .A2(b[12]), .ZN(y[156]) );
  OR2_X1 U194bar ( .A1(abar[9]), .A2(bbar[12]), .ZN(ybar[156]) );
  AND2_X1 U195 ( .A1(a[9]), .A2(b[11]), .ZN(y[155]) );
  OR2_X1 U195bar ( .A1(abar[9]), .A2(bbar[11]), .ZN(ybar[155]) );
  AND2_X1 U196 ( .A1(a[9]), .A2(b[10]), .ZN(y[154]) );
  OR2_X1 U196bar ( .A1(abar[9]), .A2(bbar[10]), .ZN(ybar[154]) );
  AND2_X1 U197 ( .A1(a[9]), .A2(b[9]), .ZN(y[153]) );
  OR2_X1 U197bar ( .A1(abar[9]), .A2(bbar[9]), .ZN(ybar[153]) );
  AND2_X1 U198 ( .A1(a[9]), .A2(b[8]), .ZN(y[152]) );
  OR2_X1 U198bar ( .A1(abar[9]), .A2(bbar[8]), .ZN(ybar[152]) );
  AND2_X1 U199 ( .A1(a[9]), .A2(b[7]), .ZN(y[151]) );
  OR2_X1 U199bar ( .A1(abar[9]), .A2(bbar[7]), .ZN(ybar[151]) );
  AND2_X1 U200 ( .A1(a[9]), .A2(b[6]), .ZN(y[150]) );
  OR2_X1 U200bar ( .A1(abar[9]), .A2(bbar[6]), .ZN(ybar[150]) );
  AND2_X1 U201 ( .A1(b[14]), .A2(a[0]), .ZN(y[14]) );
  OR2_X1 U201bar ( .A1(bbar[14]), .A2(abar[0]), .ZN(ybar[14]) );
  AND2_X1 U202 ( .A1(a[9]), .A2(b[5]), .ZN(y[149]) );
  OR2_X1 U202bar ( .A1(abar[9]), .A2(bbar[5]), .ZN(ybar[149]) );
  AND2_X1 U203 ( .A1(a[9]), .A2(b[4]), .ZN(y[148]) );
  OR2_X1 U203bar ( .A1(abar[9]), .A2(bbar[4]), .ZN(ybar[148]) );
  AND2_X1 U204 ( .A1(a[9]), .A2(b[3]), .ZN(y[147]) );
  OR2_X1 U204bar ( .A1(abar[9]), .A2(bbar[3]), .ZN(ybar[147]) );
  AND2_X1 U205 ( .A1(a[9]), .A2(b[2]), .ZN(y[146]) );
  OR2_X1 U205bar ( .A1(abar[9]), .A2(bbar[2]), .ZN(ybar[146]) );
  AND2_X1 U206 ( .A1(a[9]), .A2(b[1]), .ZN(y[145]) );
  OR2_X1 U206bar ( .A1(abar[9]), .A2(bbar[1]), .ZN(ybar[145]) );
  AND2_X1 U207 ( .A1(a[9]), .A2(b[0]), .ZN(y[144]) );
  OR2_X1 U207bar ( .A1(abar[9]), .A2(bbar[0]), .ZN(ybar[144]) );
  AND2_X1 U208 ( .A1(a[8]), .A2(b[15]), .ZN(y[143]) );
  OR2_X1 U208bar ( .A1(abar[8]), .A2(bbar[15]), .ZN(ybar[143]) );
  AND2_X1 U209 ( .A1(a[8]), .A2(b[14]), .ZN(y[142]) );
  OR2_X1 U209bar ( .A1(abar[8]), .A2(bbar[14]), .ZN(ybar[142]) );
  AND2_X1 U210 ( .A1(a[8]), .A2(b[13]), .ZN(y[141]) );
  OR2_X1 U210bar ( .A1(abar[8]), .A2(bbar[13]), .ZN(ybar[141]) );
  AND2_X1 U211 ( .A1(a[8]), .A2(b[12]), .ZN(y[140]) );
  OR2_X1 U211bar ( .A1(abar[8]), .A2(bbar[12]), .ZN(ybar[140]) );
  AND2_X1 U212 ( .A1(b[13]), .A2(a[0]), .ZN(y[13]) );
  OR2_X1 U212bar ( .A1(bbar[13]), .A2(abar[0]), .ZN(ybar[13]) );
  AND2_X1 U213 ( .A1(a[8]), .A2(b[11]), .ZN(y[139]) );
  OR2_X1 U213bar ( .A1(abar[8]), .A2(bbar[11]), .ZN(ybar[139]) );
  AND2_X1 U214 ( .A1(a[8]), .A2(b[10]), .ZN(y[138]) );
  OR2_X1 U214bar ( .A1(abar[8]), .A2(bbar[10]), .ZN(ybar[138]) );
  AND2_X1 U215 ( .A1(a[8]), .A2(b[9]), .ZN(y[137]) );
  OR2_X1 U215bar ( .A1(abar[8]), .A2(bbar[9]), .ZN(ybar[137]) );
  AND2_X1 U216 ( .A1(a[8]), .A2(b[8]), .ZN(y[136]) );
  OR2_X1 U216bar ( .A1(abar[8]), .A2(bbar[8]), .ZN(ybar[136]) );
  AND2_X1 U217 ( .A1(a[8]), .A2(b[7]), .ZN(y[135]) );
  OR2_X1 U217bar ( .A1(abar[8]), .A2(bbar[7]), .ZN(ybar[135]) );
  AND2_X1 U218 ( .A1(a[8]), .A2(b[6]), .ZN(y[134]) );
  OR2_X1 U218bar ( .A1(abar[8]), .A2(bbar[6]), .ZN(ybar[134]) );
  AND2_X1 U219 ( .A1(a[8]), .A2(b[5]), .ZN(y[133]) );
  OR2_X1 U219bar ( .A1(abar[8]), .A2(bbar[5]), .ZN(ybar[133]) );
  AND2_X1 U220 ( .A1(a[8]), .A2(b[4]), .ZN(y[132]) );
  OR2_X1 U220bar ( .A1(abar[8]), .A2(bbar[4]), .ZN(ybar[132]) );
  AND2_X1 U221 ( .A1(a[8]), .A2(b[3]), .ZN(y[131]) );
  OR2_X1 U221bar ( .A1(abar[8]), .A2(bbar[3]), .ZN(ybar[131]) );
  AND2_X1 U222 ( .A1(a[8]), .A2(b[2]), .ZN(y[130]) );
  OR2_X1 U222bar ( .A1(abar[8]), .A2(bbar[2]), .ZN(ybar[130]) );
  AND2_X1 U223 ( .A1(b[12]), .A2(a[0]), .ZN(y[12]) );
  OR2_X1 U223bar ( .A1(bbar[12]), .A2(abar[0]), .ZN(ybar[12]) );
  AND2_X1 U224 ( .A1(a[8]), .A2(b[1]), .ZN(y[129]) );
  OR2_X1 U224bar ( .A1(abar[8]), .A2(bbar[1]), .ZN(ybar[129]) );
  AND2_X1 U225 ( .A1(a[8]), .A2(b[0]), .ZN(y[128]) );
  OR2_X1 U225bar ( .A1(abar[8]), .A2(bbar[0]), .ZN(ybar[128]) );
  AND2_X1 U226 ( .A1(a[7]), .A2(b[15]), .ZN(y[127]) );
  OR2_X1 U226bar ( .A1(abar[7]), .A2(bbar[15]), .ZN(ybar[127]) );
  AND2_X1 U227 ( .A1(a[7]), .A2(b[14]), .ZN(y[126]) );
  OR2_X1 U227bar ( .A1(abar[7]), .A2(bbar[14]), .ZN(ybar[126]) );
  AND2_X1 U228 ( .A1(a[7]), .A2(b[13]), .ZN(y[125]) );
  OR2_X1 U228bar ( .A1(abar[7]), .A2(bbar[13]), .ZN(ybar[125]) );
  AND2_X1 U229 ( .A1(a[7]), .A2(b[12]), .ZN(y[124]) );
  OR2_X1 U229bar ( .A1(abar[7]), .A2(bbar[12]), .ZN(ybar[124]) );
  AND2_X1 U230 ( .A1(a[7]), .A2(b[11]), .ZN(y[123]) );
  OR2_X1 U230bar ( .A1(abar[7]), .A2(bbar[11]), .ZN(ybar[123]) );
  AND2_X1 U231 ( .A1(a[7]), .A2(b[10]), .ZN(y[122]) );
  OR2_X1 U231bar ( .A1(abar[7]), .A2(bbar[10]), .ZN(ybar[122]) );
  AND2_X1 U232 ( .A1(a[7]), .A2(b[9]), .ZN(y[121]) );
  OR2_X1 U232bar ( .A1(abar[7]), .A2(bbar[9]), .ZN(ybar[121]) );
  AND2_X1 U233 ( .A1(a[7]), .A2(b[8]), .ZN(y[120]) );
  OR2_X1 U233bar ( .A1(abar[7]), .A2(bbar[8]), .ZN(ybar[120]) );
  AND2_X1 U234 ( .A1(b[11]), .A2(a[0]), .ZN(y[11]) );
  OR2_X1 U234bar ( .A1(bbar[11]), .A2(abar[0]), .ZN(ybar[11]) );
  AND2_X1 U235 ( .A1(a[7]), .A2(b[7]), .ZN(y[119]) );
  OR2_X1 U235bar ( .A1(abar[7]), .A2(bbar[7]), .ZN(ybar[119]) );
  AND2_X1 U236 ( .A1(a[7]), .A2(b[6]), .ZN(y[118]) );
  OR2_X1 U236bar ( .A1(abar[7]), .A2(bbar[6]), .ZN(ybar[118]) );
  AND2_X1 U237 ( .A1(a[7]), .A2(b[5]), .ZN(y[117]) );
  OR2_X1 U237bar ( .A1(abar[7]), .A2(bbar[5]), .ZN(ybar[117]) );
  AND2_X1 U238 ( .A1(a[7]), .A2(b[4]), .ZN(y[116]) );
  OR2_X1 U238bar ( .A1(abar[7]), .A2(bbar[4]), .ZN(ybar[116]) );
  AND2_X1 U239 ( .A1(a[7]), .A2(b[3]), .ZN(y[115]) );
  OR2_X1 U239bar ( .A1(abar[7]), .A2(bbar[3]), .ZN(ybar[115]) );
  AND2_X1 U240 ( .A1(a[7]), .A2(b[2]), .ZN(y[114]) );
  OR2_X1 U240bar ( .A1(abar[7]), .A2(bbar[2]), .ZN(ybar[114]) );
  AND2_X1 U241 ( .A1(a[7]), .A2(b[1]), .ZN(y[113]) );
  OR2_X1 U241bar ( .A1(abar[7]), .A2(bbar[1]), .ZN(ybar[113]) );
  AND2_X1 U242 ( .A1(a[7]), .A2(b[0]), .ZN(y[112]) );
  OR2_X1 U242bar ( .A1(abar[7]), .A2(bbar[0]), .ZN(ybar[112]) );
  AND2_X1 U243 ( .A1(b[15]), .A2(a[6]), .ZN(y[111]) );
  OR2_X1 U243bar ( .A1(bbar[15]), .A2(abar[6]), .ZN(ybar[111]) );
  AND2_X1 U244 ( .A1(b[14]), .A2(a[6]), .ZN(y[110]) );
  OR2_X1 U244bar ( .A1(bbar[14]), .A2(abar[6]), .ZN(ybar[110]) );
  AND2_X1 U245 ( .A1(b[10]), .A2(a[0]), .ZN(y[10]) );
  OR2_X1 U245bar ( .A1(bbar[10]), .A2(abar[0]), .ZN(ybar[10]) );
  AND2_X1 U246 ( .A1(b[13]), .A2(a[6]), .ZN(y[109]) );
  OR2_X1 U246bar ( .A1(bbar[13]), .A2(abar[6]), .ZN(ybar[109]) );
  AND2_X1 U247 ( .A1(b[12]), .A2(a[6]), .ZN(y[108]) );
  OR2_X1 U247bar ( .A1(bbar[12]), .A2(abar[6]), .ZN(ybar[108]) );
  AND2_X1 U248 ( .A1(b[11]), .A2(a[6]), .ZN(y[107]) );
  OR2_X1 U248bar ( .A1(bbar[11]), .A2(abar[6]), .ZN(ybar[107]) );
  AND2_X1 U249 ( .A1(b[10]), .A2(a[6]), .ZN(y[106]) );
  OR2_X1 U249bar ( .A1(bbar[10]), .A2(abar[6]), .ZN(ybar[106]) );
  AND2_X1 U250 ( .A1(a[6]), .A2(b[9]), .ZN(y[105]) );
  OR2_X1 U250bar ( .A1(abar[6]), .A2(bbar[9]), .ZN(ybar[105]) );
  AND2_X1 U251 ( .A1(b[8]), .A2(a[6]), .ZN(y[104]) );
  OR2_X1 U251bar ( .A1(bbar[8]), .A2(abar[6]), .ZN(ybar[104]) );
  AND2_X1 U252 ( .A1(b[7]), .A2(a[6]), .ZN(y[103]) );
  OR2_X1 U252bar ( .A1(bbar[7]), .A2(abar[6]), .ZN(ybar[103]) );
  AND2_X1 U253 ( .A1(b[6]), .A2(a[6]), .ZN(y[102]) );
  OR2_X1 U253bar ( .A1(bbar[6]), .A2(abar[6]), .ZN(ybar[102]) );
  AND2_X1 U254 ( .A1(b[5]), .A2(a[6]), .ZN(y[101]) );
  OR2_X1 U254bar ( .A1(bbar[5]), .A2(abar[6]), .ZN(ybar[101]) );
  AND2_X1 U255 ( .A1(b[4]), .A2(a[6]), .ZN(y[100]) );
  OR2_X1 U255bar ( .A1(bbar[4]), .A2(abar[6]), .ZN(ybar[100]) );
  AND2_X1 U256 ( .A1(b[0]), .A2(a[0]), .ZN(y[0]) );
  OR2_X1 U256bar ( .A1(bbar[0]), .A2(abar[0]), .ZN(ybar[0]) );
endmodule

module decode_13 ( in, inbar, out, outbar );

  input wire [7:0] in;
  input wire [7:0] inbar;
//input_done

  output wire [255:0] out;
  output wire [255:0] outbar;
//output_done

  wire [15:0] level1;
  wire [31:0] level2;
  wire [15:0] level1bar;
  wire [31:0] level2bar;
//wire_done

  CD2_52 cd_l1_1 ( .a(in[1]), .abar(inbar[1]), .b(in[0]), .bbar(inbar[0]), .y(level1[3:0]), .ybar(level1bar[3:0]) );
  CD2_51 cd_l1_2 ( .a(in[3]), .abar(inbar[3]), .b(in[2]), .bbar(inbar[2]), .y(level1[7:4]), .ybar(level1bar[7:4]) );
  CD2_50 cd_l1_3 ( .a(in[5]), .abar(inbar[5]), .b(in[4]), .bbar(inbar[4]), .y(level1[11:8]), .ybar(level1bar[11:8]) );
  CD2_49 cd_l1_4 ( .a(in[7]), .abar(inbar[7]), .b(in[6]), .bbar(inbar[6]), .y(level1[15:12]), .ybar(level1bar[15:12]) );

  CD4_26 cd_l2_1 ( .a(level1[7:4]), .abar(level1bar[7:4]), .b(level1[3:0]), .bbar(level1bar[3:0]), 
        .y(level2[15:0]), .ybar(level2bar[15:0]) );
  CD4_25 cd_l2_2 ( .a(level1[15:12]), .abar(level1bar[15:12]), .b(level1[11:8]), .bbar(level1bar[11:8]), 
        .y(level2[31:16]), .ybar(level2bar[31:16]) );
  CD16_13 cd_l3 ( .a(level2[31:16]), .abar(level2bar[31:16]), .b(level2[15:0]), .bbar(level2bar[15:0]), 
        .y(out), .ybar(outbar) );
endmodule

module encode_13 ( in, inbar, out, outbar );

  input wire [255:0] in;
  input wire [255:0] inbar;
//input_done

  output wire [7:0] out;
  output wire [7:0] outbar;
//output_done

  wire in_81;
  wire in_80;
  wire in_79;
  wire in_78;
  wire in_77;
  wire in_76;
  wire in_75;
  wire in_74;
  wire in_73;
  wire in_72;
  wire in_71;
  wire in_70;
  wire in_69;
  wire in_68;
  wire in_67;
  wire in_66;
  wire in_65;
  wire in_64;
  wire in_63;
  wire in_62;
  wire in_61;
  wire in_60;
  wire in_59;
  wire in_58;
  wire in_57;
  wire in_56;
  wire in_55;
  wire in_54;
  wire in_53;
  wire in_52;
  wire in_51;
  wire in_50;
  wire in_49;
  wire in_48;
  wire in_47;
  wire in_46;
  wire in_45;
  wire in_44;
  wire in_43;
  wire in_42;
  wire in_41;
  wire in_40;
  wire in_39;
  wire in_38;
  wire in_37;
  wire in_36;
  wire in_35;
  wire in_34;
  wire in_33;
  wire in_32;
  wire in_31;
  wire in_30;
  wire in_29;
  wire in_28;
  wire in_27;
  wire in_26;
  wire in_25;
  wire in_24;
  wire in_23;
  wire in_22;
  wire in_21;
  wire in_20;
  wire in_19;
  wire in_18;
  wire in_17;
  wire in_16;
  wire in_15;
  wire in_14;
  wire in_13;
  wire in_12;
  wire in_11;
  wire in_10;
  wire in_9;
  wire in_8;
  wire in_7;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_3;
  wire in_2;
  wire in_1;
  wire in_0;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire in_81bar;
  wire in_80bar;
  wire in_79bar;
  wire in_78bar;
  wire in_77bar;
  wire in_76bar;
  wire in_75bar;
  wire in_74bar;
  wire in_73bar;
  wire in_72bar;
  wire in_71bar;
  wire in_70bar;
  wire in_69bar;
  wire in_68bar;
  wire in_67bar;
  wire in_66bar;
  wire in_65bar;
  wire in_64bar;
  wire in_63bar;
  wire in_62bar;
  wire in_61bar;
  wire in_60bar;
  wire in_59bar;
  wire in_58bar;
  wire in_57bar;
  wire in_56bar;
  wire in_55bar;
  wire in_54bar;
  wire in_53bar;
  wire in_52bar;
  wire in_51bar;
  wire in_50bar;
  wire in_49bar;
  wire in_48bar;
  wire in_47bar;
  wire in_46bar;
  wire in_45bar;
  wire in_44bar;
  wire in_43bar;
  wire in_42bar;
  wire in_41bar;
  wire in_40bar;
  wire in_39bar;
  wire in_38bar;
  wire in_37bar;
  wire in_36bar;
  wire in_35bar;
  wire in_34bar;
  wire in_33bar;
  wire in_32bar;
  wire in_31bar;
  wire in_30bar;
  wire in_29bar;
  wire in_28bar;
  wire in_27bar;
  wire in_26bar;
  wire in_25bar;
  wire in_24bar;
  wire in_23bar;
  wire in_22bar;
  wire in_21bar;
  wire in_20bar;
  wire in_19bar;
  wire in_18bar;
  wire in_17bar;
  wire in_16bar;
  wire in_15bar;
  wire in_14bar;
  wire in_13bar;
  wire in_12bar;
  wire in_11bar;
  wire in_10bar;
  wire in_9bar;
  wire in_8bar;
  wire in_7bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_3bar;
  wire in_2bar;
  wire in_1bar;
  wire in_0bar;
  wire n487bar;
  wire n488bar;
  wire n489bar;
  wire n490bar;
  wire n491bar;
  wire n492bar;
  wire n493bar;
  wire n494bar;
  wire n495bar;
  wire n496bar;
  wire n497bar;
  wire n498bar;
  wire n499bar;
  wire n500bar;
  wire n501bar;
  wire n502bar;
  wire n503bar;
  wire n504bar;
  wire n505bar;
  wire n506bar;
  wire n507bar;
  wire n508bar;
  wire n509bar;
  wire n510bar;
  wire n511bar;
  wire n512bar;
  wire n513bar;
  wire n514bar;
  wire n515bar;
  wire n516bar;
  wire n517bar;
  wire n518bar;
  wire n519bar;
  wire n520bar;
  wire n521bar;
  wire n522bar;
  wire n523bar;
  wire n524bar;
  wire n525bar;
  wire n526bar;
  wire n527bar;
  wire n528bar;
  wire n529bar;
  wire n530bar;
  wire n531bar;
  wire n532bar;
  wire n533bar;
  wire n534bar;
  wire n535bar;
  wire n536bar;
  wire n537bar;
  wire n538bar;
  wire n539bar;
  wire n540bar;
  wire n541bar;
  wire n542bar;
  wire n543bar;
  wire n544bar;
  wire n545bar;
  wire n546bar;
  wire n547bar;
  wire n548bar;
  wire n549bar;
  wire n550bar;
  wire n551bar;
  wire n552bar;
  wire n553bar;
  wire n554bar;
  wire n555bar;
  wire n556bar;
  wire n557bar;
  wire n558bar;
  wire n559bar;
  wire n560bar;
  wire n561bar;
  wire n562bar;
  wire n563bar;
  wire n564bar;
  wire n565bar;
  wire n566bar;
  wire n567bar;
  wire n568bar;
  wire n569bar;
  wire n570bar;
  wire n571bar;
  wire n572bar;
  wire n573bar;
  wire n574bar;
  wire n575bar;
  wire n576bar;
  wire n577bar;
  wire n578bar;
  wire n579bar;
  wire n580bar;
  wire n581bar;
  wire n582bar;
  wire n583bar;
  wire n584bar;
  wire n585bar;
  wire n586bar;
  wire n587bar;
  wire n588bar;
  wire n589bar;
  wire n590bar;
  wire n591bar;
  wire n592bar;
  wire n593bar;
  wire n594bar;
  wire n595bar;
  wire n596bar;
  wire n597bar;
  wire n598bar;
  wire n599bar;
  wire n600bar;
  wire n601bar;
  wire n602bar;
  wire n603bar;
  wire n604bar;
  wire n605bar;
  wire n606bar;
  wire n607bar;
  wire n608bar;
  wire n609bar;
  wire n610bar;
  wire n611bar;
  wire n612bar;
  wire n613bar;
  wire n614bar;
  wire n615bar;
  wire n616bar;
  wire n617bar;
  wire n618bar;
  wire n619bar;
  wire n620bar;
  wire n621bar;
  wire n622bar;
  wire n623bar;
  wire n624bar;
  wire n625bar;
  wire n626bar;
  wire n627bar;
  wire n628bar;
  wire n629bar;
  wire n630bar;
  wire n631bar;
  wire n632bar;
  wire n633bar;
  wire n634bar;
  wire n635bar;
  wire n636bar;
  wire n637bar;
  wire n638bar;
  wire n639bar;
  wire n640bar;
  wire n641bar;
  wire n642bar;
  wire n643bar;
  wire n644bar;
  wire n645bar;
  wire n646bar;
  wire n647bar;
  wire n648bar;
  wire n649bar;
  wire n650bar;
  wire n651bar;
  wire n652bar;
  wire n653bar;
  wire n654bar;
  wire n655bar;
  wire n656bar;
  wire n657bar;
  wire n658bar;
  wire n659bar;
  wire n660bar;
  wire n661bar;
  wire n662bar;
  wire n663bar;
  wire n664bar;
  wire n665bar;
  wire n666bar;
  wire n667bar;
  wire n668bar;
  wire n669bar;
  wire n670bar;
  wire n671bar;
  wire n672bar;
  wire n673bar;
  wire n674bar;
  wire n675bar;
  wire n676bar;
  wire n677bar;
  wire n678bar;
  wire n679bar;
  wire n680bar;
  wire n681bar;
  wire n682bar;
  wire n683bar;
  wire n684bar;
  wire n685bar;
  wire n686bar;
  wire n687bar;
  wire n688bar;
  wire n689bar;
  wire n690bar;
  wire n691bar;
  wire n692bar;
  wire n693bar;
  wire n694bar;
  wire n695bar;
  wire n696bar;
  wire n697bar;
  wire n698bar;
  wire n699bar;
  wire n700bar;
  wire n701bar;
  wire n702bar;
  wire n703bar;
  wire n704bar;
  wire n705bar;
  wire n706bar;
  wire n707bar;
  wire n708bar;
  wire n709bar;
  wire n710bar;
  wire n711bar;
  wire n712bar;
  wire n713bar;
  wire n714bar;
  wire n715bar;
  wire n716bar;
  wire n717bar;
  wire n718bar;
  wire n719bar;
  wire n720bar;
  wire n721bar;
  wire n722bar;
  wire n723bar;
  wire n724bar;
  wire n725bar;
  wire n726bar;
  wire n727bar;
  wire n728bar;
  wire n729bar;
  wire n730bar;
  wire n731bar;
  wire n732bar;
  wire n733bar;
  wire n734bar;
  wire n735bar;
  wire n736bar;
  wire n737bar;
  wire n738bar;
  wire n739bar;
  wire n740bar;
  wire n741bar;
  wire n742bar;
  wire n743bar;
  wire n744bar;
  wire n745bar;
  wire n746bar;
  wire n747bar;
  wire n748bar;
  wire n749bar;
  wire n750bar;
  wire n751bar;
  wire n752bar;
  wire n753bar;
  wire n754bar;
  wire n755bar;
  wire n756bar;
  wire n757bar;
  wire n758bar;
  wire n759bar;
  wire n760bar;
  wire n761bar;
  wire n762bar;
  wire n763bar;
  wire n764bar;
  wire n765bar;
  wire n766bar;
  wire n767bar;
  wire n768bar;
  wire n769bar;
  wire n770bar;
  wire n771bar;
  wire n772bar;
  wire n773bar;
  wire n774bar;
  wire n775bar;
  wire n776bar;
  wire n777bar;
  wire n778bar;
  wire n779bar;
  wire n780bar;
  wire n781bar;
  wire n782bar;
  wire n783bar;
  wire n784bar;
  wire n785bar;
  wire n786bar;
  wire n787bar;
  wire n788bar;
  wire n789bar;
  wire n790bar;
  wire n791bar;
  wire n792bar;
  wire n793bar;
  wire n794bar;
  wire n795bar;
  wire n796bar;
  wire n797bar;
  wire n798bar;
  wire n799bar;
  wire n800bar;
  wire n801bar;
  wire n802bar;
  wire n803bar;
  wire n804bar;
  wire n805bar;
  wire n806bar;
  wire n807bar;
  wire n808bar;
  wire n809bar;
  wire n810bar;
  wire n811bar;
  wire n812bar;
  wire n813bar;
  wire n814bar;
  wire n815bar;
  wire n816bar;
  wire n817bar;
  wire n818bar;
  wire n819bar;
  wire n820bar;
  wire n821bar;
  wire n822bar;
  wire n823bar;
  wire n824bar;
  wire n825bar;
  wire n826bar;
  wire n827bar;
  wire n828bar;
  wire n829bar;
  wire n830bar;
  wire n831bar;
  wire n832bar;
  wire n833bar;
  wire n834bar;
  wire n835bar;
  wire n836bar;
  wire n837bar;
  wire n838bar;
  wire n839bar;
  wire n840bar;
  wire n841bar;
  wire n842bar;
  wire n843bar;
  wire n844bar;
  wire n845bar;
  wire n846bar;
  wire n847bar;
  wire n848bar;
  wire n849bar;
  wire n850bar;
  wire n851bar;
  wire n852bar;
  wire n853bar;
  wire n854bar;
  wire n855bar;
  wire n856bar;
  wire n857bar;
  wire n858bar;
  wire n859bar;
  wire n860bar;
  wire n861bar;
  wire n862bar;
  wire n863bar;
  wire n864bar;
  wire n865bar;
  wire n866bar;
  wire n867bar;
  wire n868bar;
  wire n869bar;
  wire n870bar;
  wire n871bar;
  wire n872bar;
  wire n873bar;
  wire n874bar;
  wire n875bar;
  wire n876bar;
  wire n877bar;
  wire n878bar;
  wire n879bar;
  wire n880bar;
  wire n881bar;
  wire n882bar;
  wire n883bar;
  wire n884bar;
  wire n885bar;
  wire n886bar;
  wire n887bar;
  wire n888bar;
  wire n889bar;
  wire n890bar;
  wire n891bar;
  wire n892bar;
  wire n893bar;
  wire n894bar;
  wire n895bar;
  wire n896bar;
  wire n897bar;
  wire n898bar;
  wire n899bar;
  wire n900bar;
  wire n901bar;
  wire n902bar;
  wire n903bar;
  wire n904bar;
  wire n905bar;
  wire n906bar;
  wire n907bar;
  wire n908bar;
  wire n909bar;
  wire n910bar;
  wire n911bar;
  wire n912bar;
  wire n913bar;
  wire n914bar;
  wire n915bar;
  wire n916bar;
  wire n917bar;
  wire n918bar;
  wire n919bar;
  wire n920bar;
  wire n921bar;
  wire n922bar;
  wire n923bar;
  wire n924bar;
  wire n925bar;
  wire n926bar;
  wire n927bar;
  wire n928bar;
  wire n929bar;
  wire n930bar;
  wire n931bar;
  wire n932bar;
  wire n933bar;
  wire n934bar;
  wire n935bar;
  wire n936bar;
  wire n937bar;
  wire n938bar;
  wire n939bar;
  wire n940bar;
  wire n941bar;
  wire n942bar;
  wire n943bar;
  wire n944bar;
  wire n945bar;
  wire n946bar;
  wire n947bar;
  wire n948bar;
  wire n949bar;
  wire n950bar;
  wire n951bar;
  wire n952bar;
  wire n953bar;
  wire n954bar;
  wire n955bar;
  wire n956bar;
  wire n957bar;
  wire n958bar;
  wire n959bar;
  wire n960bar;
  wire n961bar;
  wire n962bar;
  wire n963bar;
  wire n964bar;
  wire n965bar;
  wire n966bar;
  wire n967bar;
  wire n968bar;
  wire n969bar;
  wire n970bar;
  wire n971bar;
  wire n972bar;
//wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];
  assign in_81bar = inbar[81];
  assign in_80bar = inbar[80];
  assign in_79bar = inbar[79];
  assign in_78bar = inbar[78];
  assign in_77bar = inbar[77];
  assign in_76bar = inbar[76];
  assign in_75bar = inbar[75];
  assign in_74bar = inbar[74];
  assign in_73bar = inbar[73];
  assign in_72bar = inbar[72];
  assign in_71bar = inbar[71];
  assign in_70bar = inbar[70];
  assign in_69bar = inbar[69];
  assign in_68bar = inbar[68];
  assign in_67bar = inbar[67];
  assign in_66bar = inbar[66];
  assign in_65bar = inbar[65];
  assign in_64bar = inbar[64];
  assign in_63bar = inbar[63];
  assign in_62bar = inbar[62];
  assign in_61bar = inbar[61];
  assign in_60bar = inbar[60];
  assign in_59bar = inbar[59];
  assign in_58bar = inbar[58];
  assign in_57bar = inbar[57];
  assign in_56bar = inbar[56];
  assign in_55bar = inbar[55];
  assign in_54bar = inbar[54];
  assign in_53bar = inbar[53];
  assign in_52bar = inbar[52];
  assign in_51bar = inbar[51];
  assign in_50bar = inbar[50];
  assign in_49bar = inbar[49];
  assign in_48bar = inbar[48];
  assign in_47bar = inbar[47];
  assign in_46bar = inbar[46];
  assign in_45bar = inbar[45];
  assign in_44bar = inbar[44];
  assign in_43bar = inbar[43];
  assign in_42bar = inbar[42];
  assign in_41bar = inbar[41];
  assign in_40bar = inbar[40];
  assign in_39bar = inbar[39];
  assign in_38bar = inbar[38];
  assign in_37bar = inbar[37];
  assign in_36bar = inbar[36];
  assign in_35bar = inbar[35];
  assign in_34bar = inbar[34];
  assign in_33bar = inbar[33];
  assign in_32bar = inbar[32];
  assign in_31bar = inbar[31];
  assign in_30bar = inbar[30];
  assign in_29bar = inbar[29];
  assign in_28bar = inbar[28];
  assign in_27bar = inbar[27];
  assign in_26bar = inbar[26];
  assign in_25bar = inbar[25];
  assign in_24bar = inbar[24];
  assign in_23bar = inbar[23];
  assign in_22bar = inbar[22];
  assign in_21bar = inbar[21];
  assign in_20bar = inbar[20];
  assign in_19bar = inbar[19];
  assign in_18bar = inbar[18];
  assign in_17bar = inbar[17];
  assign in_16bar = inbar[16];
  assign in_15bar = inbar[15];
  assign in_14bar = inbar[14];
  assign in_13bar = inbar[13];
  assign in_12bar = inbar[12];
  assign in_11bar = inbar[11];
  assign in_10bar = inbar[10];
  assign in_9bar = inbar[9];
  assign in_8bar = inbar[8];
  assign in_7bar = inbar[7];
  assign in_6bar = inbar[6];
  assign in_5bar = inbar[5];
  assign in_4bar = inbar[4];
  assign in_3bar = inbar[3];
  assign in_2bar = inbar[2];
  assign in_1bar = inbar[1];
  assign in_0bar = inbar[0];
//assign_done

  OR2_X1 U1 ( .A1(n972), .A2(n971), .ZN(out[7]) );
  AND2_X1 U1bar ( .A1(n972bar), .A2(n971bar), .ZN(outbar[7]) );
  OR2_X1 U2 ( .A1(n970), .A2(n969), .ZN(n971) );
  AND2_X1 U2bar ( .A1(n970bar), .A2(n969bar), .ZN(n971bar) );
  OR2_X1 U3 ( .A1(n968), .A2(n967), .ZN(n969) );
  AND2_X1 U3bar ( .A1(n968bar), .A2(n967bar), .ZN(n969bar) );
  OR2_X1 U4 ( .A1(n966), .A2(n965), .ZN(n967) );
  AND2_X1 U4bar ( .A1(n966bar), .A2(n965bar), .ZN(n967bar) );
  OR2_X1 U5 ( .A1(n964), .A2(n963), .ZN(n968) );
  AND2_X1 U5bar ( .A1(n964bar), .A2(n963bar), .ZN(n968bar) );
  OR2_X1 U6 ( .A1(in[116]), .A2(n962), .ZN(n963) );
  AND2_X1 U6bar ( .A1(inbar[116]), .A2(n962bar), .ZN(n963bar) );
  OR2_X1 U7 ( .A1(n961), .A2(n960), .ZN(n970) );
  AND2_X1 U7bar ( .A1(n961bar), .A2(n960bar), .ZN(n970bar) );
  OR2_X1 U8 ( .A1(in[150]), .A2(in[127]), .ZN(n960) );
  AND2_X1 U8bar ( .A1(inbar[150]), .A2(inbar[127]), .ZN(n960bar) );
  OR2_X1 U9 ( .A1(in[160]), .A2(n959), .ZN(n961) );
  AND2_X1 U9bar ( .A1(inbar[160]), .A2(n959bar), .ZN(n961bar) );
  OR2_X1 U10 ( .A1(in[252]), .A2(in[168]), .ZN(n959) );
  AND2_X1 U10bar ( .A1(inbar[252]), .A2(inbar[168]), .ZN(n959bar) );
  OR2_X1 U11 ( .A1(n958), .A2(n957), .ZN(n972) );
  AND2_X1 U11bar ( .A1(n958bar), .A2(n957bar), .ZN(n972bar) );
  OR2_X1 U12 ( .A1(n956), .A2(n955), .ZN(n957) );
  AND2_X1 U12bar ( .A1(n956bar), .A2(n955bar), .ZN(n957bar) );
  OR2_X1 U13 ( .A1(in_17), .A2(in[96]), .ZN(n955) );
  AND2_X1 U13bar ( .A1(in_17bar), .A2(inbar[96]), .ZN(n955bar) );
  OR2_X1 U14 ( .A1(in_23), .A2(n954), .ZN(n956) );
  AND2_X1 U14bar ( .A1(in_23bar), .A2(n954bar), .ZN(n956bar) );
  OR2_X1 U15 ( .A1(in_31), .A2(in_26), .ZN(n954) );
  AND2_X1 U15bar ( .A1(in_31bar), .A2(in_26bar), .ZN(n954bar) );
  OR2_X1 U16 ( .A1(n953), .A2(n952), .ZN(n958) );
  AND2_X1 U16bar ( .A1(n953bar), .A2(n952bar), .ZN(n958bar) );
  OR2_X1 U17 ( .A1(in_58), .A2(in_4), .ZN(n952) );
  AND2_X1 U17bar ( .A1(in_58bar), .A2(in_4bar), .ZN(n952bar) );
  OR2_X1 U18 ( .A1(in_59), .A2(n951), .ZN(n953) );
  AND2_X1 U18bar ( .A1(in_59bar), .A2(n951bar), .ZN(n953bar) );
  OR2_X1 U19 ( .A1(in_71), .A2(in_62), .ZN(n951) );
  AND2_X1 U19bar ( .A1(in_71bar), .A2(in_62bar), .ZN(n951bar) );
  OR2_X1 U20 ( .A1(n950), .A2(n949), .ZN(out[6]) );
  AND2_X1 U20bar ( .A1(n950bar), .A2(n949bar), .ZN(outbar[6]) );
  OR2_X1 U21 ( .A1(n948), .A2(n947), .ZN(n949) );
  AND2_X1 U21bar ( .A1(n948bar), .A2(n947bar), .ZN(n949bar) );
  OR2_X1 U22 ( .A1(n946), .A2(n945), .ZN(n947) );
  AND2_X1 U22bar ( .A1(n946bar), .A2(n945bar), .ZN(n947bar) );
  OR2_X1 U23 ( .A1(n944), .A2(n943), .ZN(n945) );
  AND2_X1 U23bar ( .A1(n944bar), .A2(n943bar), .ZN(n945bar) );
  OR2_X1 U24 ( .A1(n942), .A2(n941), .ZN(n946) );
  AND2_X1 U24bar ( .A1(n942bar), .A2(n941bar), .ZN(n946bar) );
  OR2_X1 U25 ( .A1(in[101]), .A2(n940), .ZN(n941) );
  AND2_X1 U25bar ( .A1(inbar[101]), .A2(n940bar), .ZN(n941bar) );
  OR2_X1 U26 ( .A1(n939), .A2(n938), .ZN(n948) );
  AND2_X1 U26bar ( .A1(n939bar), .A2(n938bar), .ZN(n948bar) );
  OR2_X1 U27 ( .A1(in[114]), .A2(in[104]), .ZN(n938) );
  AND2_X1 U27bar ( .A1(inbar[114]), .A2(inbar[104]), .ZN(n938bar) );
  OR2_X1 U28 ( .A1(in[128]), .A2(n937), .ZN(n939) );
  AND2_X1 U28bar ( .A1(inbar[128]), .A2(n937bar), .ZN(n939bar) );
  OR2_X1 U29 ( .A1(in[136]), .A2(in[134]), .ZN(n937) );
  AND2_X1 U29bar ( .A1(inbar[136]), .A2(inbar[134]), .ZN(n937bar) );
  OR2_X1 U30 ( .A1(n936), .A2(n935), .ZN(n950) );
  AND2_X1 U30bar ( .A1(n936bar), .A2(n935bar), .ZN(n950bar) );
  OR2_X1 U31 ( .A1(n934), .A2(n933), .ZN(n935) );
  AND2_X1 U31bar ( .A1(n934bar), .A2(n933bar), .ZN(n935bar) );
  OR2_X1 U32 ( .A1(in[177]), .A2(in[164]), .ZN(n933) );
  AND2_X1 U32bar ( .A1(inbar[177]), .A2(inbar[164]), .ZN(n933bar) );
  OR2_X1 U33 ( .A1(in[212]), .A2(n932), .ZN(n934) );
  AND2_X1 U33bar ( .A1(inbar[212]), .A2(n932bar), .ZN(n934bar) );
  OR2_X1 U34 ( .A1(in[248]), .A2(in[221]), .ZN(n932) );
  AND2_X1 U34bar ( .A1(inbar[248]), .A2(inbar[221]), .ZN(n932bar) );
  OR2_X1 U35 ( .A1(n931), .A2(n930), .ZN(n936) );
  AND2_X1 U35bar ( .A1(n931bar), .A2(n930bar), .ZN(n936bar) );
  OR2_X1 U36 ( .A1(in_18), .A2(in[93]), .ZN(n930) );
  AND2_X1 U36bar ( .A1(in_18bar), .A2(inbar[93]), .ZN(n930bar) );
  OR2_X1 U37 ( .A1(in_31), .A2(n929), .ZN(n931) );
  AND2_X1 U37bar ( .A1(in_31bar), .A2(n929bar), .ZN(n931bar) );
  OR2_X1 U38 ( .A1(in_7), .A2(in_39), .ZN(n929) );
  AND2_X1 U38bar ( .A1(in_7bar), .A2(in_39bar), .ZN(n929bar) );
  OR2_X1 U39 ( .A1(n928), .A2(n927), .ZN(out[5]) );
  AND2_X1 U39bar ( .A1(n928bar), .A2(n927bar), .ZN(outbar[5]) );
  OR2_X1 U40 ( .A1(n926), .A2(n925), .ZN(n927) );
  AND2_X1 U40bar ( .A1(n926bar), .A2(n925bar), .ZN(n927bar) );
  OR2_X1 U41 ( .A1(n924), .A2(n923), .ZN(n925) );
  AND2_X1 U41bar ( .A1(n924bar), .A2(n923bar), .ZN(n925bar) );
  OR2_X1 U42 ( .A1(n922), .A2(n921), .ZN(n923) );
  AND2_X1 U42bar ( .A1(n922bar), .A2(n921bar), .ZN(n923bar) );
  OR2_X1 U43 ( .A1(n940), .A2(n920), .ZN(n924) );
  AND2_X1 U43bar ( .A1(n940bar), .A2(n920bar), .ZN(n924bar) );
  OR2_X1 U44 ( .A1(in[111]), .A2(n919), .ZN(n920) );
  AND2_X1 U44bar ( .A1(inbar[111]), .A2(n919bar), .ZN(n920bar) );
  OR2_X1 U45 ( .A1(n918), .A2(n917), .ZN(n940) );
  AND2_X1 U45bar ( .A1(n918bar), .A2(n917bar), .ZN(n940bar) );
  OR2_X1 U46 ( .A1(n916), .A2(n915), .ZN(n917) );
  AND2_X1 U46bar ( .A1(n916bar), .A2(n915bar), .ZN(n917bar) );
  OR2_X1 U47 ( .A1(n914), .A2(n913), .ZN(n915) );
  AND2_X1 U47bar ( .A1(n914bar), .A2(n913bar), .ZN(n915bar) );
  OR2_X1 U48 ( .A1(in[140]), .A2(in[131]), .ZN(n913) );
  AND2_X1 U48bar ( .A1(inbar[140]), .A2(inbar[131]), .ZN(n913bar) );
  OR2_X1 U49 ( .A1(in[160]), .A2(in[144]), .ZN(n914) );
  AND2_X1 U49bar ( .A1(inbar[160]), .A2(inbar[144]), .ZN(n914bar) );
  OR2_X1 U50 ( .A1(n912), .A2(n911), .ZN(n916) );
  AND2_X1 U50bar ( .A1(n912bar), .A2(n911bar), .ZN(n916bar) );
  OR2_X1 U51 ( .A1(in[179]), .A2(in[174]), .ZN(n911) );
  AND2_X1 U51bar ( .A1(inbar[179]), .A2(inbar[174]), .ZN(n911bar) );
  OR2_X1 U52 ( .A1(in[188]), .A2(in[184]), .ZN(n912) );
  AND2_X1 U52bar ( .A1(inbar[188]), .A2(inbar[184]), .ZN(n912bar) );
  OR2_X1 U53 ( .A1(n910), .A2(n909), .ZN(n918) );
  AND2_X1 U53bar ( .A1(n910bar), .A2(n909bar), .ZN(n918bar) );
  OR2_X1 U54 ( .A1(n908), .A2(n907), .ZN(n909) );
  AND2_X1 U54bar ( .A1(n908bar), .A2(n907bar), .ZN(n909bar) );
  OR2_X1 U55 ( .A1(in[216]), .A2(in[200]), .ZN(n907) );
  AND2_X1 U55bar ( .A1(inbar[216]), .A2(inbar[200]), .ZN(n907bar) );
  OR2_X1 U56 ( .A1(in[228]), .A2(in[224]), .ZN(n908) );
  AND2_X1 U56bar ( .A1(inbar[228]), .A2(inbar[224]), .ZN(n908bar) );
  OR2_X1 U57 ( .A1(n906), .A2(n905), .ZN(n910) );
  AND2_X1 U57bar ( .A1(n906bar), .A2(n905bar), .ZN(n910bar) );
  OR2_X1 U58 ( .A1(in[247]), .A2(in[235]), .ZN(n905) );
  AND2_X1 U58bar ( .A1(inbar[247]), .A2(inbar[235]), .ZN(n905bar) );
  OR2_X1 U59 ( .A1(in_42), .A2(in[83]), .ZN(n906) );
  AND2_X1 U59bar ( .A1(in_42bar), .A2(inbar[83]), .ZN(n906bar) );
  OR2_X1 U60 ( .A1(n904), .A2(n903), .ZN(n926) );
  AND2_X1 U60bar ( .A1(n904bar), .A2(n903bar), .ZN(n926bar) );
  OR2_X1 U61 ( .A1(in[166]), .A2(in[123]), .ZN(n903) );
  AND2_X1 U61bar ( .A1(inbar[166]), .A2(inbar[123]), .ZN(n903bar) );
  OR2_X1 U62 ( .A1(in[170]), .A2(n902), .ZN(n904) );
  AND2_X1 U62bar ( .A1(inbar[170]), .A2(n902bar), .ZN(n904bar) );
  OR2_X1 U63 ( .A1(in[194]), .A2(in[183]), .ZN(n902) );
  AND2_X1 U63bar ( .A1(inbar[194]), .A2(inbar[183]), .ZN(n902bar) );
  OR2_X1 U64 ( .A1(n901), .A2(n900), .ZN(n928) );
  AND2_X1 U64bar ( .A1(n901bar), .A2(n900bar), .ZN(n928bar) );
  OR2_X1 U65 ( .A1(n899), .A2(n898), .ZN(n900) );
  AND2_X1 U65bar ( .A1(n899bar), .A2(n898bar), .ZN(n900bar) );
  OR2_X1 U66 ( .A1(in[241]), .A2(in[238]), .ZN(n898) );
  AND2_X1 U66bar ( .A1(inbar[241]), .A2(inbar[238]), .ZN(n898bar) );
  OR2_X1 U67 ( .A1(in[250]), .A2(n897), .ZN(n899) );
  AND2_X1 U67bar ( .A1(inbar[250]), .A2(n897bar), .ZN(n899bar) );
  OR2_X1 U68 ( .A1(in_24), .A2(in[84]), .ZN(n897) );
  AND2_X1 U68bar ( .A1(in_24bar), .A2(inbar[84]), .ZN(n897bar) );
  OR2_X1 U69 ( .A1(n896), .A2(n895), .ZN(n901) );
  AND2_X1 U69bar ( .A1(n896bar), .A2(n895bar), .ZN(n901bar) );
  OR2_X1 U70 ( .A1(in_41), .A2(in_29), .ZN(n895) );
  AND2_X1 U70bar ( .A1(in_41bar), .A2(in_29bar), .ZN(n895bar) );
  OR2_X1 U71 ( .A1(in_66), .A2(n894), .ZN(n896) );
  AND2_X1 U71bar ( .A1(in_66bar), .A2(n894bar), .ZN(n896bar) );
  OR2_X1 U72 ( .A1(in_76), .A2(in_71), .ZN(n894) );
  AND2_X1 U72bar ( .A1(in_76bar), .A2(in_71bar), .ZN(n894bar) );
  OR2_X1 U73 ( .A1(n893), .A2(n892), .ZN(out[4]) );
  AND2_X1 U73bar ( .A1(n893bar), .A2(n892bar), .ZN(outbar[4]) );
  OR2_X1 U74 ( .A1(n891), .A2(n890), .ZN(n892) );
  AND2_X1 U74bar ( .A1(n891bar), .A2(n890bar), .ZN(n892bar) );
  OR2_X1 U75 ( .A1(n889), .A2(n888), .ZN(n890) );
  AND2_X1 U75bar ( .A1(n889bar), .A2(n888bar), .ZN(n890bar) );
  OR2_X1 U76 ( .A1(n922), .A2(n887), .ZN(n888) );
  AND2_X1 U76bar ( .A1(n922bar), .A2(n887bar), .ZN(n888bar) );
  OR2_X1 U77 ( .A1(n886), .A2(n885), .ZN(n922) );
  AND2_X1 U77bar ( .A1(n886bar), .A2(n885bar), .ZN(n922bar) );
  OR2_X1 U78 ( .A1(n884), .A2(n883), .ZN(n885) );
  AND2_X1 U78bar ( .A1(n884bar), .A2(n883bar), .ZN(n885bar) );
  OR2_X1 U79 ( .A1(n882), .A2(n881), .ZN(n883) );
  AND2_X1 U79bar ( .A1(n882bar), .A2(n881bar), .ZN(n883bar) );
  OR2_X1 U80 ( .A1(in[118]), .A2(in[109]), .ZN(n881) );
  AND2_X1 U80bar ( .A1(inbar[118]), .A2(inbar[109]), .ZN(n881bar) );
  OR2_X1 U81 ( .A1(in[139]), .A2(in[120]), .ZN(n882) );
  AND2_X1 U81bar ( .A1(inbar[139]), .A2(inbar[120]), .ZN(n882bar) );
  OR2_X1 U82 ( .A1(n880), .A2(n879), .ZN(n884) );
  AND2_X1 U82bar ( .A1(n880bar), .A2(n879bar), .ZN(n884bar) );
  OR2_X1 U83 ( .A1(in[198]), .A2(in[154]), .ZN(n879) );
  AND2_X1 U83bar ( .A1(inbar[198]), .A2(inbar[154]), .ZN(n879bar) );
  OR2_X1 U84 ( .A1(in[210]), .A2(in[205]), .ZN(n880) );
  AND2_X1 U84bar ( .A1(inbar[210]), .A2(inbar[205]), .ZN(n880bar) );
  OR2_X1 U85 ( .A1(n878), .A2(n877), .ZN(n886) );
  AND2_X1 U85bar ( .A1(n878bar), .A2(n877bar), .ZN(n886bar) );
  OR2_X1 U86 ( .A1(n876), .A2(n875), .ZN(n877) );
  AND2_X1 U86bar ( .A1(n876bar), .A2(n875bar), .ZN(n877bar) );
  OR2_X1 U87 ( .A1(in[219]), .A2(in[217]), .ZN(n875) );
  AND2_X1 U87bar ( .A1(inbar[219]), .A2(inbar[217]), .ZN(n875bar) );
  OR2_X1 U88 ( .A1(in[86]), .A2(in[252]), .ZN(n876) );
  AND2_X1 U88bar ( .A1(inbar[86]), .A2(inbar[252]), .ZN(n876bar) );
  OR2_X1 U89 ( .A1(n874), .A2(n873), .ZN(n878) );
  AND2_X1 U89bar ( .A1(n874bar), .A2(n873bar), .ZN(n878bar) );
  OR2_X1 U90 ( .A1(in_40), .A2(in[91]), .ZN(n873) );
  AND2_X1 U90bar ( .A1(in_40bar), .A2(inbar[91]), .ZN(n873bar) );
  OR2_X1 U91 ( .A1(in_8), .A2(in_46), .ZN(n874) );
  AND2_X1 U91bar ( .A1(in_8bar), .A2(in_46bar), .ZN(n874bar) );
  OR2_X1 U92 ( .A1(n872), .A2(n871), .ZN(n889) );
  AND2_X1 U92bar ( .A1(n872bar), .A2(n871bar), .ZN(n889bar) );
  OR2_X1 U93 ( .A1(in[117]), .A2(n943), .ZN(n871) );
  AND2_X1 U93bar ( .A1(inbar[117]), .A2(n943bar), .ZN(n871bar) );
  OR2_X1 U94 ( .A1(n870), .A2(n869), .ZN(n943) );
  AND2_X1 U94bar ( .A1(n870bar), .A2(n869bar), .ZN(n943bar) );
  OR2_X1 U95 ( .A1(n868), .A2(n867), .ZN(n869) );
  AND2_X1 U95bar ( .A1(n868bar), .A2(n867bar), .ZN(n869bar) );
  OR2_X1 U96 ( .A1(n866), .A2(n865), .ZN(n867) );
  AND2_X1 U96bar ( .A1(n866bar), .A2(n865bar), .ZN(n867bar) );
  OR2_X1 U97 ( .A1(n864), .A2(n863), .ZN(n865) );
  AND2_X1 U97bar ( .A1(n864bar), .A2(n863bar), .ZN(n865bar) );
  OR2_X1 U98 ( .A1(in[108]), .A2(n919), .ZN(n866) );
  AND2_X1 U98bar ( .A1(inbar[108]), .A2(n919bar), .ZN(n866bar) );
  OR2_X1 U99 ( .A1(n862), .A2(n861), .ZN(n919) );
  AND2_X1 U99bar ( .A1(n862bar), .A2(n861bar), .ZN(n919bar) );
  OR2_X1 U100 ( .A1(n860), .A2(n859), .ZN(n861) );
  AND2_X1 U100bar ( .A1(n860bar), .A2(n859bar), .ZN(n861bar) );
  OR2_X1 U101 ( .A1(n858), .A2(n857), .ZN(n859) );
  AND2_X1 U101bar ( .A1(n858bar), .A2(n857bar), .ZN(n859bar) );
  OR2_X1 U102 ( .A1(in[119]), .A2(in[105]), .ZN(n857) );
  AND2_X1 U102bar ( .A1(inbar[119]), .A2(inbar[105]), .ZN(n857bar) );
  OR2_X1 U103 ( .A1(in[186]), .A2(in[175]), .ZN(n858) );
  AND2_X1 U103bar ( .A1(inbar[186]), .A2(inbar[175]), .ZN(n858bar) );
  OR2_X1 U104 ( .A1(n856), .A2(n855), .ZN(n860) );
  AND2_X1 U104bar ( .A1(n856bar), .A2(n855bar), .ZN(n860bar) );
  OR2_X1 U105 ( .A1(in[202]), .A2(in[193]), .ZN(n855) );
  AND2_X1 U105bar ( .A1(inbar[202]), .A2(inbar[193]), .ZN(n855bar) );
  OR2_X1 U106 ( .A1(in[225]), .A2(in[208]), .ZN(n856) );
  AND2_X1 U106bar ( .A1(inbar[225]), .A2(inbar[208]), .ZN(n856bar) );
  OR2_X1 U107 ( .A1(n854), .A2(n853), .ZN(n862) );
  AND2_X1 U107bar ( .A1(n854bar), .A2(n853bar), .ZN(n862bar) );
  OR2_X1 U108 ( .A1(n852), .A2(n851), .ZN(n853) );
  AND2_X1 U108bar ( .A1(n852bar), .A2(n851bar), .ZN(n853bar) );
  OR2_X1 U109 ( .A1(in_1), .A2(in[85]), .ZN(n851) );
  AND2_X1 U109bar ( .A1(in_1bar), .A2(inbar[85]), .ZN(n851bar) );
  OR2_X1 U110 ( .A1(in_23), .A2(in_19), .ZN(n852) );
  AND2_X1 U110bar ( .A1(in_23bar), .A2(in_19bar), .ZN(n852bar) );
  OR2_X1 U111 ( .A1(n850), .A2(n849), .ZN(n854) );
  AND2_X1 U111bar ( .A1(n850bar), .A2(n849bar), .ZN(n854bar) );
  OR2_X1 U112 ( .A1(in_43), .A2(in_33), .ZN(n849) );
  AND2_X1 U112bar ( .A1(in_43bar), .A2(in_33bar), .ZN(n849bar) );
  OR2_X1 U113 ( .A1(in_63), .A2(in_44), .ZN(n850) );
  AND2_X1 U113bar ( .A1(in_63bar), .A2(in_44bar), .ZN(n850bar) );
  OR2_X1 U114 ( .A1(n848), .A2(n847), .ZN(n868) );
  AND2_X1 U114bar ( .A1(n848bar), .A2(n847bar), .ZN(n868bar) );
  OR2_X1 U115 ( .A1(in[141]), .A2(in[112]), .ZN(n847) );
  AND2_X1 U115bar ( .A1(inbar[141]), .A2(inbar[112]), .ZN(n847bar) );
  OR2_X1 U116 ( .A1(in[147]), .A2(n846), .ZN(n848) );
  AND2_X1 U116bar ( .A1(inbar[147]), .A2(n846bar), .ZN(n848bar) );
  OR2_X1 U117 ( .A1(in[181]), .A2(in[167]), .ZN(n846) );
  AND2_X1 U117bar ( .A1(inbar[181]), .A2(inbar[167]), .ZN(n846bar) );
  OR2_X1 U118 ( .A1(n845), .A2(n844), .ZN(n870) );
  AND2_X1 U118bar ( .A1(n845bar), .A2(n844bar), .ZN(n870bar) );
  OR2_X1 U119 ( .A1(n843), .A2(n842), .ZN(n844) );
  AND2_X1 U119bar ( .A1(n843bar), .A2(n842bar), .ZN(n844bar) );
  OR2_X1 U120 ( .A1(in[229]), .A2(in[201]), .ZN(n842) );
  AND2_X1 U120bar ( .A1(inbar[229]), .A2(inbar[201]), .ZN(n842bar) );
  OR2_X1 U121 ( .A1(in[237]), .A2(n841), .ZN(n843) );
  AND2_X1 U121bar ( .A1(inbar[237]), .A2(n841bar), .ZN(n843bar) );
  OR2_X1 U122 ( .A1(in[94]), .A2(in[253]), .ZN(n841) );
  AND2_X1 U122bar ( .A1(inbar[94]), .A2(inbar[253]), .ZN(n841bar) );
  OR2_X1 U123 ( .A1(n840), .A2(n839), .ZN(n845) );
  AND2_X1 U123bar ( .A1(n840bar), .A2(n839bar), .ZN(n845bar) );
  OR2_X1 U124 ( .A1(in_21), .A2(in[96]), .ZN(n839) );
  AND2_X1 U124bar ( .A1(in_21bar), .A2(inbar[96]), .ZN(n839bar) );
  OR2_X1 U125 ( .A1(in_25), .A2(n838), .ZN(n840) );
  AND2_X1 U125bar ( .A1(in_25bar), .A2(n838bar), .ZN(n840bar) );
  OR2_X1 U126 ( .A1(in_81), .A2(in_45), .ZN(n838) );
  AND2_X1 U126bar ( .A1(in_81bar), .A2(in_45bar), .ZN(n838bar) );
  OR2_X1 U127 ( .A1(n837), .A2(n836), .ZN(n891) );
  AND2_X1 U127bar ( .A1(n837bar), .A2(n836bar), .ZN(n891bar) );
  OR2_X1 U128 ( .A1(in[142]), .A2(in[124]), .ZN(n836) );
  AND2_X1 U128bar ( .A1(inbar[142]), .A2(inbar[124]), .ZN(n836bar) );
  OR2_X1 U129 ( .A1(in[150]), .A2(n835), .ZN(n837) );
  AND2_X1 U129bar ( .A1(inbar[150]), .A2(n835bar), .ZN(n837bar) );
  OR2_X1 U130 ( .A1(in[172]), .A2(in[155]), .ZN(n835) );
  AND2_X1 U130bar ( .A1(inbar[172]), .A2(inbar[155]), .ZN(n835bar) );
  OR2_X1 U131 ( .A1(n834), .A2(n833), .ZN(n893) );
  AND2_X1 U131bar ( .A1(n834bar), .A2(n833bar), .ZN(n893bar) );
  OR2_X1 U132 ( .A1(n832), .A2(n831), .ZN(n833) );
  AND2_X1 U132bar ( .A1(n832bar), .A2(n831bar), .ZN(n833bar) );
  OR2_X1 U133 ( .A1(in[196]), .A2(in[173]), .ZN(n831) );
  AND2_X1 U133bar ( .A1(inbar[196]), .A2(inbar[173]), .ZN(n831bar) );
  OR2_X1 U134 ( .A1(in[222]), .A2(n830), .ZN(n832) );
  AND2_X1 U134bar ( .A1(inbar[222]), .A2(n830bar), .ZN(n832bar) );
  OR2_X1 U135 ( .A1(in[227]), .A2(in[226]), .ZN(n830) );
  AND2_X1 U135bar ( .A1(inbar[227]), .A2(inbar[226]), .ZN(n830bar) );
  OR2_X1 U136 ( .A1(n829), .A2(n828), .ZN(n834) );
  AND2_X1 U136bar ( .A1(n829bar), .A2(n828bar), .ZN(n834bar) );
  OR2_X1 U137 ( .A1(in[249]), .A2(in[231]), .ZN(n828) );
  AND2_X1 U137bar ( .A1(inbar[249]), .A2(inbar[231]), .ZN(n828bar) );
  OR2_X1 U138 ( .A1(in_28), .A2(n827), .ZN(n829) );
  AND2_X1 U138bar ( .A1(in_28bar), .A2(n827bar), .ZN(n829bar) );
  OR2_X1 U139 ( .A1(in_52), .A2(in_47), .ZN(n827) );
  AND2_X1 U139bar ( .A1(in_52bar), .A2(in_47bar), .ZN(n827bar) );
  OR2_X1 U140 ( .A1(n826), .A2(n825), .ZN(out[3]) );
  AND2_X1 U140bar ( .A1(n826bar), .A2(n825bar), .ZN(outbar[3]) );
  OR2_X1 U141 ( .A1(n824), .A2(n823), .ZN(n825) );
  AND2_X1 U141bar ( .A1(n824bar), .A2(n823bar), .ZN(n825bar) );
  OR2_X1 U142 ( .A1(n822), .A2(n821), .ZN(n823) );
  AND2_X1 U142bar ( .A1(n822bar), .A2(n821bar), .ZN(n823bar) );
  OR2_X1 U143 ( .A1(n820), .A2(n819), .ZN(n821) );
  AND2_X1 U143bar ( .A1(n820bar), .A2(n819bar), .ZN(n821bar) );
  OR2_X1 U144 ( .A1(n964), .A2(n818), .ZN(n822) );
  AND2_X1 U144bar ( .A1(n964bar), .A2(n818bar), .ZN(n822bar) );
  OR2_X1 U145 ( .A1(in[118]), .A2(n817), .ZN(n818) );
  AND2_X1 U145bar ( .A1(inbar[118]), .A2(n817bar), .ZN(n818bar) );
  OR2_X1 U146 ( .A1(n816), .A2(n815), .ZN(n964) );
  AND2_X1 U146bar ( .A1(n816bar), .A2(n815bar), .ZN(n964bar) );
  OR2_X1 U147 ( .A1(n814), .A2(n813), .ZN(n815) );
  AND2_X1 U147bar ( .A1(n814bar), .A2(n813bar), .ZN(n815bar) );
  OR2_X1 U148 ( .A1(n812), .A2(n811), .ZN(n813) );
  AND2_X1 U148bar ( .A1(n812bar), .A2(n811bar), .ZN(n813bar) );
  OR2_X1 U149 ( .A1(in[122]), .A2(in[111]), .ZN(n811) );
  AND2_X1 U149bar ( .A1(inbar[122]), .A2(inbar[111]), .ZN(n811bar) );
  OR2_X1 U150 ( .A1(in[154]), .A2(in[151]), .ZN(n812) );
  AND2_X1 U150bar ( .A1(inbar[154]), .A2(inbar[151]), .ZN(n812bar) );
  OR2_X1 U151 ( .A1(n810), .A2(n809), .ZN(n814) );
  AND2_X1 U151bar ( .A1(n810bar), .A2(n809bar), .ZN(n814bar) );
  OR2_X1 U152 ( .A1(in[187]), .A2(in[177]), .ZN(n809) );
  AND2_X1 U152bar ( .A1(inbar[187]), .A2(inbar[177]), .ZN(n809bar) );
  OR2_X1 U153 ( .A1(in[200]), .A2(in[192]), .ZN(n810) );
  AND2_X1 U153bar ( .A1(inbar[200]), .A2(inbar[192]), .ZN(n810bar) );
  OR2_X1 U154 ( .A1(n808), .A2(n807), .ZN(n816) );
  AND2_X1 U154bar ( .A1(n808bar), .A2(n807bar), .ZN(n816bar) );
  OR2_X1 U155 ( .A1(n806), .A2(n805), .ZN(n807) );
  AND2_X1 U155bar ( .A1(n806bar), .A2(n805bar), .ZN(n807bar) );
  OR2_X1 U156 ( .A1(in[225]), .A2(in[207]), .ZN(n805) );
  AND2_X1 U156bar ( .A1(inbar[225]), .A2(inbar[207]), .ZN(n805bar) );
  OR2_X1 U157 ( .A1(in[98]), .A2(in[226]), .ZN(n806) );
  AND2_X1 U157bar ( .A1(inbar[98]), .A2(inbar[226]), .ZN(n806bar) );
  OR2_X1 U158 ( .A1(n804), .A2(n803), .ZN(n808) );
  AND2_X1 U158bar ( .A1(n804bar), .A2(n803bar), .ZN(n808bar) );
  OR2_X1 U159 ( .A1(in_20), .A2(in_16), .ZN(n803) );
  AND2_X1 U159bar ( .A1(in_20bar), .A2(in_16bar), .ZN(n803bar) );
  OR2_X1 U160 ( .A1(in_55), .A2(in_45), .ZN(n804) );
  AND2_X1 U160bar ( .A1(in_55bar), .A2(in_45bar), .ZN(n804bar) );
  OR2_X1 U161 ( .A1(n802), .A2(n801), .ZN(n824) );
  AND2_X1 U161bar ( .A1(n802bar), .A2(n801bar), .ZN(n824bar) );
  OR2_X1 U162 ( .A1(in[162]), .A2(in[149]), .ZN(n801) );
  AND2_X1 U162bar ( .A1(inbar[162]), .A2(inbar[149]), .ZN(n801bar) );
  OR2_X1 U163 ( .A1(in[163]), .A2(n800), .ZN(n802) );
  AND2_X1 U163bar ( .A1(inbar[163]), .A2(n800bar), .ZN(n802bar) );
  OR2_X1 U164 ( .A1(in[191]), .A2(in[189]), .ZN(n800) );
  AND2_X1 U164bar ( .A1(inbar[191]), .A2(inbar[189]), .ZN(n800bar) );
  OR2_X1 U165 ( .A1(n799), .A2(n798), .ZN(n826) );
  AND2_X1 U165bar ( .A1(n799bar), .A2(n798bar), .ZN(n826bar) );
  OR2_X1 U166 ( .A1(n797), .A2(n796), .ZN(n798) );
  AND2_X1 U166bar ( .A1(n797bar), .A2(n796bar), .ZN(n798bar) );
  OR2_X1 U167 ( .A1(in[212]), .A2(in[193]), .ZN(n796) );
  AND2_X1 U167bar ( .A1(inbar[212]), .A2(inbar[193]), .ZN(n796bar) );
  OR2_X1 U168 ( .A1(in[238]), .A2(n795), .ZN(n797) );
  AND2_X1 U168bar ( .A1(inbar[238]), .A2(n795bar), .ZN(n797bar) );
  OR2_X1 U169 ( .A1(in[88]), .A2(in[247]), .ZN(n795) );
  AND2_X1 U169bar ( .A1(inbar[88]), .A2(inbar[247]), .ZN(n795bar) );
  OR2_X1 U170 ( .A1(n794), .A2(n793), .ZN(n799) );
  AND2_X1 U170bar ( .A1(n794bar), .A2(n793bar), .ZN(n799bar) );
  OR2_X1 U171 ( .A1(in[94]), .A2(in[92]), .ZN(n793) );
  AND2_X1 U171bar ( .A1(inbar[94]), .A2(inbar[92]), .ZN(n793bar) );
  OR2_X1 U172 ( .A1(in_52), .A2(n792), .ZN(n794) );
  AND2_X1 U172bar ( .A1(in_52bar), .A2(n792bar), .ZN(n794bar) );
  OR2_X1 U173 ( .A1(in_70), .A2(in_67), .ZN(n792) );
  AND2_X1 U173bar ( .A1(in_70bar), .A2(in_67bar), .ZN(n792bar) );
  OR2_X1 U174 ( .A1(n791), .A2(n790), .ZN(out[2]) );
  AND2_X1 U174bar ( .A1(n791bar), .A2(n790bar), .ZN(outbar[2]) );
  OR2_X1 U175 ( .A1(n789), .A2(n788), .ZN(n790) );
  AND2_X1 U175bar ( .A1(n789bar), .A2(n788bar), .ZN(n790bar) );
  OR2_X1 U176 ( .A1(n787), .A2(n786), .ZN(n788) );
  AND2_X1 U176bar ( .A1(n787bar), .A2(n786bar), .ZN(n788bar) );
  OR2_X1 U177 ( .A1(n819), .A2(n785), .ZN(n786) );
  AND2_X1 U177bar ( .A1(n819bar), .A2(n785bar), .ZN(n786bar) );
  OR2_X1 U178 ( .A1(n784), .A2(n783), .ZN(n819) );
  AND2_X1 U178bar ( .A1(n784bar), .A2(n783bar), .ZN(n819bar) );
  OR2_X1 U179 ( .A1(n782), .A2(n781), .ZN(n783) );
  AND2_X1 U179bar ( .A1(n782bar), .A2(n781bar), .ZN(n783bar) );
  OR2_X1 U180 ( .A1(n780), .A2(n779), .ZN(n781) );
  AND2_X1 U180bar ( .A1(n780bar), .A2(n779bar), .ZN(n781bar) );
  OR2_X1 U181 ( .A1(n962), .A2(n778), .ZN(n779) );
  AND2_X1 U181bar ( .A1(n962bar), .A2(n778bar), .ZN(n779bar) );
  OR2_X1 U182 ( .A1(n777), .A2(n776), .ZN(n962) );
  AND2_X1 U182bar ( .A1(n777bar), .A2(n776bar), .ZN(n962bar) );
  OR2_X1 U183 ( .A1(n775), .A2(n774), .ZN(n776) );
  AND2_X1 U183bar ( .A1(n775bar), .A2(n774bar), .ZN(n776bar) );
  OR2_X1 U184 ( .A1(n773), .A2(n772), .ZN(n774) );
  AND2_X1 U184bar ( .A1(n773bar), .A2(n772bar), .ZN(n774bar) );
  OR2_X1 U185 ( .A1(in[131]), .A2(in[120]), .ZN(n772) );
  AND2_X1 U185bar ( .A1(inbar[131]), .A2(inbar[120]), .ZN(n772bar) );
  OR2_X1 U186 ( .A1(in[153]), .A2(in[147]), .ZN(n773) );
  AND2_X1 U186bar ( .A1(inbar[153]), .A2(inbar[147]), .ZN(n773bar) );
  OR2_X1 U187 ( .A1(n771), .A2(n770), .ZN(n775) );
  AND2_X1 U187bar ( .A1(n771bar), .A2(n770bar), .ZN(n775bar) );
  OR2_X1 U188 ( .A1(in[170]), .A2(in[156]), .ZN(n770) );
  AND2_X1 U188bar ( .A1(inbar[170]), .A2(inbar[156]), .ZN(n770bar) );
  OR2_X1 U189 ( .A1(in[223]), .A2(in[190]), .ZN(n771) );
  AND2_X1 U189bar ( .A1(inbar[223]), .A2(inbar[190]), .ZN(n771bar) );
  OR2_X1 U190 ( .A1(n769), .A2(n768), .ZN(n777) );
  AND2_X1 U190bar ( .A1(n769bar), .A2(n768bar), .ZN(n777bar) );
  OR2_X1 U191 ( .A1(n767), .A2(n766), .ZN(n768) );
  AND2_X1 U191bar ( .A1(n767bar), .A2(n766bar), .ZN(n768bar) );
  OR2_X1 U192 ( .A1(in[236]), .A2(in[230]), .ZN(n766) );
  AND2_X1 U192bar ( .A1(inbar[236]), .A2(inbar[230]), .ZN(n766bar) );
  OR2_X1 U193 ( .A1(in[85]), .A2(in[240]), .ZN(n767) );
  AND2_X1 U193bar ( .A1(inbar[85]), .A2(inbar[240]), .ZN(n767bar) );
  OR2_X1 U194 ( .A1(n765), .A2(n764), .ZN(n769) );
  AND2_X1 U194bar ( .A1(n765bar), .A2(n764bar), .ZN(n769bar) );
  OR2_X1 U195 ( .A1(in_12), .A2(in[90]), .ZN(n764) );
  AND2_X1 U195bar ( .A1(in_12bar), .A2(inbar[90]), .ZN(n764bar) );
  OR2_X1 U196 ( .A1(in_39), .A2(in_28), .ZN(n765) );
  AND2_X1 U196bar ( .A1(in_39bar), .A2(in_28bar), .ZN(n765bar) );
  OR2_X1 U197 ( .A1(in[109]), .A2(n763), .ZN(n780) );
  AND2_X1 U197bar ( .A1(inbar[109]), .A2(n763bar), .ZN(n780bar) );
  OR2_X1 U198 ( .A1(n762), .A2(n761), .ZN(n782) );
  AND2_X1 U198bar ( .A1(n762bar), .A2(n761bar), .ZN(n782bar) );
  OR2_X1 U199 ( .A1(in[138]), .A2(in[129]), .ZN(n761) );
  AND2_X1 U199bar ( .A1(inbar[138]), .A2(inbar[129]), .ZN(n761bar) );
  OR2_X1 U200 ( .A1(in[157]), .A2(n760), .ZN(n762) );
  AND2_X1 U200bar ( .A1(inbar[157]), .A2(n760bar), .ZN(n762bar) );
  OR2_X1 U201 ( .A1(in[182]), .A2(in[167]), .ZN(n760) );
  AND2_X1 U201bar ( .A1(inbar[182]), .A2(inbar[167]), .ZN(n760bar) );
  OR2_X1 U202 ( .A1(n759), .A2(n758), .ZN(n784) );
  AND2_X1 U202bar ( .A1(n759bar), .A2(n758bar), .ZN(n784bar) );
  OR2_X1 U203 ( .A1(n757), .A2(n756), .ZN(n758) );
  AND2_X1 U203bar ( .A1(n757bar), .A2(n756bar), .ZN(n758bar) );
  OR2_X1 U204 ( .A1(in[195]), .A2(in[184]), .ZN(n756) );
  AND2_X1 U204bar ( .A1(inbar[195]), .A2(inbar[184]), .ZN(n756bar) );
  OR2_X1 U205 ( .A1(in[196]), .A2(n755), .ZN(n757) );
  AND2_X1 U205bar ( .A1(inbar[196]), .A2(n755bar), .ZN(n757bar) );
  OR2_X1 U206 ( .A1(in[215]), .A2(in[209]), .ZN(n755) );
  AND2_X1 U206bar ( .A1(inbar[215]), .A2(inbar[209]), .ZN(n755bar) );
  OR2_X1 U207 ( .A1(n754), .A2(n753), .ZN(n759) );
  AND2_X1 U207bar ( .A1(n754bar), .A2(n753bar), .ZN(n759bar) );
  OR2_X1 U208 ( .A1(in[93]), .A2(in[233]), .ZN(n753) );
  AND2_X1 U208bar ( .A1(inbar[93]), .A2(inbar[233]), .ZN(n753bar) );
  OR2_X1 U209 ( .A1(in_1), .A2(n752), .ZN(n754) );
  AND2_X1 U209bar ( .A1(in_1bar), .A2(n752bar), .ZN(n754bar) );
  OR2_X1 U210 ( .A1(in_69), .A2(in_66), .ZN(n752) );
  AND2_X1 U210bar ( .A1(in_69bar), .A2(in_66bar), .ZN(n752bar) );
  OR2_X1 U211 ( .A1(n966), .A2(n751), .ZN(n787) );
  AND2_X1 U211bar ( .A1(n966bar), .A2(n751bar), .ZN(n787bar) );
  OR2_X1 U212 ( .A1(in[134]), .A2(n750), .ZN(n751) );
  AND2_X1 U212bar ( .A1(inbar[134]), .A2(n750bar), .ZN(n751bar) );
  OR2_X1 U213 ( .A1(n749), .A2(n748), .ZN(n966) );
  AND2_X1 U213bar ( .A1(n749bar), .A2(n748bar), .ZN(n966bar) );
  OR2_X1 U214 ( .A1(n747), .A2(n746), .ZN(n748) );
  AND2_X1 U214bar ( .A1(n747bar), .A2(n746bar), .ZN(n748bar) );
  OR2_X1 U215 ( .A1(n745), .A2(n744), .ZN(n746) );
  AND2_X1 U215bar ( .A1(n745bar), .A2(n744bar), .ZN(n746bar) );
  OR2_X1 U216 ( .A1(in[136]), .A2(in[121]), .ZN(n744) );
  AND2_X1 U216bar ( .A1(inbar[136]), .A2(inbar[121]), .ZN(n744bar) );
  OR2_X1 U217 ( .A1(in[186]), .A2(in[174]), .ZN(n745) );
  AND2_X1 U217bar ( .A1(inbar[186]), .A2(inbar[174]), .ZN(n745bar) );
  OR2_X1 U218 ( .A1(n743), .A2(n742), .ZN(n747) );
  AND2_X1 U218bar ( .A1(n743bar), .A2(n742bar), .ZN(n747bar) );
  OR2_X1 U219 ( .A1(in[198]), .A2(in[197]), .ZN(n742) );
  AND2_X1 U219bar ( .A1(inbar[198]), .A2(inbar[197]), .ZN(n742bar) );
  OR2_X1 U220 ( .A1(in[214]), .A2(in[199]), .ZN(n743) );
  AND2_X1 U220bar ( .A1(inbar[214]), .A2(inbar[199]), .ZN(n743bar) );
  OR2_X1 U221 ( .A1(n741), .A2(n740), .ZN(n749) );
  AND2_X1 U221bar ( .A1(n741bar), .A2(n740bar), .ZN(n749bar) );
  OR2_X1 U222 ( .A1(n739), .A2(n738), .ZN(n740) );
  AND2_X1 U222bar ( .A1(n739bar), .A2(n738bar), .ZN(n740bar) );
  OR2_X1 U223 ( .A1(in[231]), .A2(in[220]), .ZN(n738) );
  AND2_X1 U223bar ( .A1(inbar[231]), .A2(inbar[220]), .ZN(n738bar) );
  OR2_X1 U224 ( .A1(in_25), .A2(in[245]), .ZN(n739) );
  AND2_X1 U224bar ( .A1(in_25bar), .A2(inbar[245]), .ZN(n739bar) );
  OR2_X1 U225 ( .A1(n737), .A2(n736), .ZN(n741) );
  AND2_X1 U225bar ( .A1(n737bar), .A2(n736bar), .ZN(n741bar) );
  OR2_X1 U226 ( .A1(in_53), .A2(in_29), .ZN(n736) );
  AND2_X1 U226bar ( .A1(in_53bar), .A2(in_29bar), .ZN(n736bar) );
  OR2_X1 U227 ( .A1(in_79), .A2(in_74), .ZN(n737) );
  AND2_X1 U227bar ( .A1(in_79bar), .A2(in_74bar), .ZN(n737bar) );
  OR2_X1 U228 ( .A1(n735), .A2(n734), .ZN(n789) );
  AND2_X1 U228bar ( .A1(n735bar), .A2(n734bar), .ZN(n789bar) );
  OR2_X1 U229 ( .A1(in[152]), .A2(in[140]), .ZN(n734) );
  AND2_X1 U229bar ( .A1(inbar[152]), .A2(inbar[140]), .ZN(n734bar) );
  OR2_X1 U230 ( .A1(in[155]), .A2(n733), .ZN(n735) );
  AND2_X1 U230bar ( .A1(inbar[155]), .A2(n733bar), .ZN(n735bar) );
  OR2_X1 U231 ( .A1(in[166]), .A2(in[165]), .ZN(n733) );
  AND2_X1 U231bar ( .A1(inbar[166]), .A2(inbar[165]), .ZN(n733bar) );
  OR2_X1 U232 ( .A1(n732), .A2(n731), .ZN(n791) );
  AND2_X1 U232bar ( .A1(n732bar), .A2(n731bar), .ZN(n791bar) );
  OR2_X1 U233 ( .A1(n730), .A2(n729), .ZN(n731) );
  AND2_X1 U233bar ( .A1(n730bar), .A2(n729bar), .ZN(n731bar) );
  OR2_X1 U234 ( .A1(in[202]), .A2(in[185]), .ZN(n729) );
  AND2_X1 U234bar ( .A1(inbar[202]), .A2(inbar[185]), .ZN(n729bar) );
  OR2_X1 U235 ( .A1(in[211]), .A2(n728), .ZN(n730) );
  AND2_X1 U235bar ( .A1(inbar[211]), .A2(n728bar), .ZN(n730bar) );
  OR2_X1 U236 ( .A1(in[255]), .A2(in[253]), .ZN(n728) );
  AND2_X1 U236bar ( .A1(inbar[255]), .A2(inbar[253]), .ZN(n728bar) );
  OR2_X1 U237 ( .A1(n727), .A2(n726), .ZN(n732) );
  AND2_X1 U237bar ( .A1(n727bar), .A2(n726bar), .ZN(n732bar) );
  OR2_X1 U238 ( .A1(in_35), .A2(in_15), .ZN(n726) );
  AND2_X1 U238bar ( .A1(in_35bar), .A2(in_15bar), .ZN(n726bar) );
  OR2_X1 U239 ( .A1(in_36), .A2(n725), .ZN(n727) );
  AND2_X1 U239bar ( .A1(in_36bar), .A2(n725bar), .ZN(n727bar) );
  OR2_X1 U240 ( .A1(in_48), .A2(in_40), .ZN(n725) );
  AND2_X1 U240bar ( .A1(in_48bar), .A2(in_40bar), .ZN(n725bar) );
  OR2_X1 U241 ( .A1(n724), .A2(n723), .ZN(out[1]) );
  AND2_X1 U241bar ( .A1(n724bar), .A2(n723bar), .ZN(outbar[1]) );
  OR2_X1 U242 ( .A1(n722), .A2(n721), .ZN(n723) );
  AND2_X1 U242bar ( .A1(n722bar), .A2(n721bar), .ZN(n723bar) );
  OR2_X1 U243 ( .A1(n720), .A2(n719), .ZN(n721) );
  AND2_X1 U243bar ( .A1(n720bar), .A2(n719bar), .ZN(n721bar) );
  OR2_X1 U244 ( .A1(n921), .A2(n887), .ZN(n719) );
  AND2_X1 U244bar ( .A1(n921bar), .A2(n887bar), .ZN(n719bar) );
  OR2_X1 U245 ( .A1(n718), .A2(n717), .ZN(n887) );
  AND2_X1 U245bar ( .A1(n718bar), .A2(n717bar), .ZN(n887bar) );
  OR2_X1 U246 ( .A1(n716), .A2(n715), .ZN(n717) );
  AND2_X1 U246bar ( .A1(n716bar), .A2(n715bar), .ZN(n717bar) );
  OR2_X1 U247 ( .A1(n714), .A2(n713), .ZN(n715) );
  AND2_X1 U247bar ( .A1(n714bar), .A2(n713bar), .ZN(n715bar) );
  OR2_X1 U248 ( .A1(in[116]), .A2(in[110]), .ZN(n713) );
  AND2_X1 U248bar ( .A1(inbar[116]), .A2(inbar[110]), .ZN(n713bar) );
  OR2_X1 U249 ( .A1(in[133]), .A2(in[130]), .ZN(n714) );
  AND2_X1 U249bar ( .A1(inbar[133]), .A2(inbar[130]), .ZN(n714bar) );
  OR2_X1 U250 ( .A1(n712), .A2(n711), .ZN(n716) );
  AND2_X1 U250bar ( .A1(n712bar), .A2(n711bar), .ZN(n716bar) );
  OR2_X1 U251 ( .A1(in[203]), .A2(in[135]), .ZN(n711) );
  AND2_X1 U251bar ( .A1(inbar[203]), .A2(inbar[135]), .ZN(n711bar) );
  OR2_X1 U252 ( .A1(in[232]), .A2(in[223]), .ZN(n712) );
  AND2_X1 U252bar ( .A1(inbar[232]), .A2(inbar[223]), .ZN(n712bar) );
  OR2_X1 U253 ( .A1(n710), .A2(n709), .ZN(n718) );
  AND2_X1 U253bar ( .A1(n710bar), .A2(n709bar), .ZN(n718bar) );
  OR2_X1 U254 ( .A1(n708), .A2(n707), .ZN(n709) );
  AND2_X1 U254bar ( .A1(n708bar), .A2(n707bar), .ZN(n709bar) );
  OR2_X1 U255 ( .A1(in[255]), .A2(in[233]), .ZN(n707) );
  AND2_X1 U255bar ( .A1(inbar[255]), .A2(inbar[233]), .ZN(n707bar) );
  OR2_X1 U256 ( .A1(in_53), .A2(in_34), .ZN(n708) );
  AND2_X1 U256bar ( .A1(in_53bar), .A2(in_34bar), .ZN(n708bar) );
  OR2_X1 U257 ( .A1(n706), .A2(n705), .ZN(n710) );
  AND2_X1 U257bar ( .A1(n706bar), .A2(n705bar), .ZN(n710bar) );
  OR2_X1 U258 ( .A1(in_57), .A2(in_55), .ZN(n705) );
  AND2_X1 U258bar ( .A1(in_57bar), .A2(in_55bar), .ZN(n705bar) );
  OR2_X1 U259 ( .A1(in_68), .A2(in_67), .ZN(n706) );
  AND2_X1 U259bar ( .A1(in_68bar), .A2(in_67bar), .ZN(n706bar) );
  OR2_X1 U260 ( .A1(n704), .A2(n703), .ZN(n921) );
  AND2_X1 U260bar ( .A1(n704bar), .A2(n703bar), .ZN(n921bar) );
  OR2_X1 U261 ( .A1(n702), .A2(n701), .ZN(n703) );
  AND2_X1 U261bar ( .A1(n702bar), .A2(n701bar), .ZN(n703bar) );
  OR2_X1 U262 ( .A1(n700), .A2(n699), .ZN(n701) );
  AND2_X1 U262bar ( .A1(n700bar), .A2(n699bar), .ZN(n701bar) );
  OR2_X1 U263 ( .A1(n944), .A2(n872), .ZN(n699) );
  AND2_X1 U263bar ( .A1(n944bar), .A2(n872bar), .ZN(n699bar) );
  OR2_X1 U264 ( .A1(n698), .A2(n697), .ZN(n872) );
  AND2_X1 U264bar ( .A1(n698bar), .A2(n697bar), .ZN(n872bar) );
  OR2_X1 U265 ( .A1(n696), .A2(n695), .ZN(n697) );
  AND2_X1 U265bar ( .A1(n696bar), .A2(n695bar), .ZN(n697bar) );
  OR2_X1 U266 ( .A1(n694), .A2(n693), .ZN(n695) );
  AND2_X1 U266bar ( .A1(n694bar), .A2(n693bar), .ZN(n695bar) );
  OR2_X1 U267 ( .A1(in[121]), .A2(in[102]), .ZN(n693) );
  AND2_X1 U267bar ( .A1(inbar[121]), .A2(inbar[102]), .ZN(n693bar) );
  OR2_X1 U268 ( .A1(in[162]), .A2(in[161]), .ZN(n694) );
  AND2_X1 U268bar ( .A1(inbar[162]), .A2(inbar[161]), .ZN(n694bar) );
  OR2_X1 U269 ( .A1(n692), .A2(n691), .ZN(n696) );
  AND2_X1 U269bar ( .A1(n692bar), .A2(n691bar), .ZN(n696bar) );
  OR2_X1 U270 ( .A1(in[192]), .A2(in[178]), .ZN(n691) );
  AND2_X1 U270bar ( .A1(inbar[192]), .A2(inbar[178]), .ZN(n691bar) );
  OR2_X1 U271 ( .A1(in[244]), .A2(in[209]), .ZN(n692) );
  AND2_X1 U271bar ( .A1(inbar[244]), .A2(inbar[209]), .ZN(n692bar) );
  OR2_X1 U272 ( .A1(n690), .A2(n689), .ZN(n698) );
  AND2_X1 U272bar ( .A1(n690bar), .A2(n689bar), .ZN(n698bar) );
  OR2_X1 U273 ( .A1(n688), .A2(n687), .ZN(n689) );
  AND2_X1 U273bar ( .A1(n688bar), .A2(n687bar), .ZN(n689bar) );
  OR2_X1 U274 ( .A1(in[90]), .A2(in[254]), .ZN(n687) );
  AND2_X1 U274bar ( .A1(inbar[90]), .A2(inbar[254]), .ZN(n687bar) );
  OR2_X1 U275 ( .A1(in_36), .A2(in_32), .ZN(n688) );
  AND2_X1 U275bar ( .A1(in_36bar), .A2(in_32bar), .ZN(n688bar) );
  OR2_X1 U276 ( .A1(n686), .A2(n685), .ZN(n690) );
  AND2_X1 U276bar ( .A1(n686bar), .A2(n685bar), .ZN(n690bar) );
  OR2_X1 U277 ( .A1(in_62), .A2(in_37), .ZN(n685) );
  AND2_X1 U277bar ( .A1(in_62bar), .A2(in_37bar), .ZN(n685bar) );
  OR2_X1 U278 ( .A1(in_75), .A2(in_73), .ZN(n686) );
  AND2_X1 U278bar ( .A1(in_75bar), .A2(in_73bar), .ZN(n686bar) );
  OR2_X1 U279 ( .A1(n684), .A2(n683), .ZN(n944) );
  AND2_X1 U279bar ( .A1(n684bar), .A2(n683bar), .ZN(n944bar) );
  OR2_X1 U280 ( .A1(n682), .A2(n681), .ZN(n683) );
  AND2_X1 U280bar ( .A1(n682bar), .A2(n681bar), .ZN(n683bar) );
  OR2_X1 U281 ( .A1(n680), .A2(n679), .ZN(n681) );
  AND2_X1 U281bar ( .A1(n680bar), .A2(n679bar), .ZN(n681bar) );
  OR2_X1 U282 ( .A1(in[171]), .A2(in[153]), .ZN(n679) );
  AND2_X1 U282bar ( .A1(inbar[171]), .A2(inbar[153]), .ZN(n679bar) );
  OR2_X1 U283 ( .A1(in[187]), .A2(in[176]), .ZN(n680) );
  AND2_X1 U283bar ( .A1(inbar[187]), .A2(inbar[176]), .ZN(n680bar) );
  OR2_X1 U284 ( .A1(n678), .A2(n677), .ZN(n682) );
  AND2_X1 U284bar ( .A1(n678bar), .A2(n677bar), .ZN(n682bar) );
  OR2_X1 U285 ( .A1(in[245]), .A2(in[211]), .ZN(n677) );
  AND2_X1 U285bar ( .A1(inbar[245]), .A2(inbar[211]), .ZN(n677bar) );
  OR2_X1 U286 ( .A1(in[97]), .A2(in[88]), .ZN(n678) );
  AND2_X1 U286bar ( .A1(inbar[97]), .A2(inbar[88]), .ZN(n678bar) );
  OR2_X1 U287 ( .A1(n676), .A2(n675), .ZN(n684) );
  AND2_X1 U287bar ( .A1(n676bar), .A2(n675bar), .ZN(n684bar) );
  OR2_X1 U288 ( .A1(n674), .A2(n673), .ZN(n675) );
  AND2_X1 U288bar ( .A1(n674bar), .A2(n673bar), .ZN(n675bar) );
  OR2_X1 U289 ( .A1(in_10), .A2(in_0), .ZN(n673) );
  AND2_X1 U289bar ( .A1(in_10bar), .A2(in_0bar), .ZN(n673bar) );
  OR2_X1 U290 ( .A1(in_59), .A2(in_5), .ZN(n674) );
  AND2_X1 U290bar ( .A1(in_59bar), .A2(in_5bar), .ZN(n674bar) );
  OR2_X1 U291 ( .A1(n672), .A2(n671), .ZN(n676) );
  AND2_X1 U291bar ( .A1(n672bar), .A2(n671bar), .ZN(n676bar) );
  OR2_X1 U292 ( .A1(in_60), .A2(in_6), .ZN(n671) );
  AND2_X1 U292bar ( .A1(in_60bar), .A2(in_6bar), .ZN(n671bar) );
  OR2_X1 U293 ( .A1(in_77), .A2(in_69), .ZN(n672) );
  AND2_X1 U293bar ( .A1(in_77bar), .A2(in_69bar), .ZN(n672bar) );
  OR2_X1 U294 ( .A1(in[113]), .A2(n864), .ZN(n700) );
  AND2_X1 U294bar ( .A1(inbar[113]), .A2(n864bar), .ZN(n700bar) );
  OR2_X1 U295 ( .A1(n670), .A2(n669), .ZN(n864) );
  AND2_X1 U295bar ( .A1(n670bar), .A2(n669bar), .ZN(n864bar) );
  OR2_X1 U296 ( .A1(n668), .A2(n667), .ZN(n669) );
  AND2_X1 U296bar ( .A1(n668bar), .A2(n667bar), .ZN(n669bar) );
  OR2_X1 U297 ( .A1(n666), .A2(n665), .ZN(n667) );
  AND2_X1 U297bar ( .A1(n666bar), .A2(n665bar), .ZN(n667bar) );
  OR2_X1 U298 ( .A1(in[125]), .A2(in[107]), .ZN(n665) );
  AND2_X1 U298bar ( .A1(inbar[125]), .A2(inbar[107]), .ZN(n665bar) );
  OR2_X1 U299 ( .A1(in[138]), .A2(in[126]), .ZN(n666) );
  AND2_X1 U299bar ( .A1(inbar[138]), .A2(inbar[126]), .ZN(n666bar) );
  OR2_X1 U300 ( .A1(n664), .A2(n663), .ZN(n668) );
  AND2_X1 U300bar ( .A1(n664bar), .A2(n663bar), .ZN(n668bar) );
  OR2_X1 U301 ( .A1(in[189]), .A2(in[143]), .ZN(n663) );
  AND2_X1 U301bar ( .A1(inbar[189]), .A2(inbar[143]), .ZN(n663bar) );
  OR2_X1 U302 ( .A1(in[99]), .A2(in[214]), .ZN(n664) );
  AND2_X1 U302bar ( .A1(inbar[99]), .A2(inbar[214]), .ZN(n664bar) );
  OR2_X1 U303 ( .A1(n662), .A2(n661), .ZN(n670) );
  AND2_X1 U303bar ( .A1(n662bar), .A2(n661bar), .ZN(n670bar) );
  OR2_X1 U304 ( .A1(n660), .A2(n659), .ZN(n661) );
  AND2_X1 U304bar ( .A1(n660bar), .A2(n659bar), .ZN(n661bar) );
  OR2_X1 U305 ( .A1(in_15), .A2(in_12), .ZN(n659) );
  AND2_X1 U305bar ( .A1(in_15bar), .A2(in_12bar), .ZN(n659bar) );
  OR2_X1 U306 ( .A1(in_20), .A2(in_2), .ZN(n660) );
  AND2_X1 U306bar ( .A1(in_20bar), .A2(in_2bar), .ZN(n660bar) );
  OR2_X1 U307 ( .A1(n658), .A2(n657), .ZN(n662) );
  AND2_X1 U307bar ( .A1(n658bar), .A2(n657bar), .ZN(n662bar) );
  OR2_X1 U308 ( .A1(in_30), .A2(in_3), .ZN(n657) );
  AND2_X1 U308bar ( .A1(in_30bar), .A2(in_3bar), .ZN(n657bar) );
  OR2_X1 U309 ( .A1(in_4), .A2(in_38), .ZN(n658) );
  AND2_X1 U309bar ( .A1(in_4bar), .A2(in_38bar), .ZN(n658bar) );
  OR2_X1 U310 ( .A1(n656), .A2(n655), .ZN(n702) );
  AND2_X1 U310bar ( .A1(n656bar), .A2(n655bar), .ZN(n702bar) );
  OR2_X1 U311 ( .A1(in[148]), .A2(in[137]), .ZN(n655) );
  AND2_X1 U311bar ( .A1(inbar[148]), .A2(inbar[137]), .ZN(n655bar) );
  OR2_X1 U312 ( .A1(in[149]), .A2(n654), .ZN(n656) );
  AND2_X1 U312bar ( .A1(inbar[149]), .A2(n654bar), .ZN(n656bar) );
  OR2_X1 U313 ( .A1(in[195]), .A2(in[190]), .ZN(n654) );
  AND2_X1 U313bar ( .A1(inbar[195]), .A2(inbar[190]), .ZN(n654bar) );
  OR2_X1 U314 ( .A1(n653), .A2(n652), .ZN(n704) );
  AND2_X1 U314bar ( .A1(n653bar), .A2(n652bar), .ZN(n704bar) );
  OR2_X1 U315 ( .A1(n651), .A2(n650), .ZN(n652) );
  AND2_X1 U315bar ( .A1(n651bar), .A2(n650bar), .ZN(n652bar) );
  OR2_X1 U316 ( .A1(in[98]), .A2(in[197]), .ZN(n650) );
  AND2_X1 U316bar ( .A1(inbar[98]), .A2(inbar[197]), .ZN(n650bar) );
  OR2_X1 U317 ( .A1(in_11), .A2(n649), .ZN(n651) );
  AND2_X1 U317bar ( .A1(in_11bar), .A2(n649bar), .ZN(n651bar) );
  OR2_X1 U318 ( .A1(in_26), .A2(in_14), .ZN(n649) );
  AND2_X1 U318bar ( .A1(in_26bar), .A2(in_14bar), .ZN(n649bar) );
  OR2_X1 U319 ( .A1(n648), .A2(n647), .ZN(n653) );
  AND2_X1 U319bar ( .A1(n648bar), .A2(n647bar), .ZN(n653bar) );
  OR2_X1 U320 ( .A1(in_35), .A2(in_27), .ZN(n647) );
  AND2_X1 U320bar ( .A1(in_35bar), .A2(in_27bar), .ZN(n647bar) );
  OR2_X1 U321 ( .A1(in_50), .A2(n646), .ZN(n648) );
  AND2_X1 U321bar ( .A1(in_50bar), .A2(n646bar), .ZN(n648bar) );
  OR2_X1 U322 ( .A1(in_78), .A2(in_61), .ZN(n646) );
  AND2_X1 U322bar ( .A1(in_78bar), .A2(in_61bar), .ZN(n646bar) );
  OR2_X1 U323 ( .A1(n942), .A2(n645), .ZN(n720) );
  AND2_X1 U323bar ( .A1(n942bar), .A2(n645bar), .ZN(n720bar) );
  OR2_X1 U324 ( .A1(in[106]), .A2(n863), .ZN(n645) );
  AND2_X1 U324bar ( .A1(inbar[106]), .A2(n863bar), .ZN(n645bar) );
  OR2_X1 U325 ( .A1(n644), .A2(n643), .ZN(n863) );
  AND2_X1 U325bar ( .A1(n644bar), .A2(n643bar), .ZN(n863bar) );
  OR2_X1 U326 ( .A1(n642), .A2(n641), .ZN(n643) );
  AND2_X1 U326bar ( .A1(n642bar), .A2(n641bar), .ZN(n643bar) );
  OR2_X1 U327 ( .A1(n640), .A2(n639), .ZN(n641) );
  AND2_X1 U327bar ( .A1(n640bar), .A2(n639bar), .ZN(n641bar) );
  OR2_X1 U328 ( .A1(in[127]), .A2(in[122]), .ZN(n639) );
  AND2_X1 U328bar ( .A1(inbar[127]), .A2(inbar[122]), .ZN(n639bar) );
  OR2_X1 U329 ( .A1(in[156]), .A2(in[132]), .ZN(n640) );
  AND2_X1 U329bar ( .A1(inbar[156]), .A2(inbar[132]), .ZN(n640bar) );
  OR2_X1 U330 ( .A1(n638), .A2(n637), .ZN(n642) );
  AND2_X1 U330bar ( .A1(n638bar), .A2(n637bar), .ZN(n642bar) );
  OR2_X1 U331 ( .A1(in[159]), .A2(in[157]), .ZN(n637) );
  AND2_X1 U331bar ( .A1(inbar[159]), .A2(inbar[157]), .ZN(n637bar) );
  OR2_X1 U332 ( .A1(in[185]), .A2(in[169]), .ZN(n638) );
  AND2_X1 U332bar ( .A1(inbar[185]), .A2(inbar[169]), .ZN(n638bar) );
  OR2_X1 U333 ( .A1(n636), .A2(n635), .ZN(n644) );
  AND2_X1 U333bar ( .A1(n636bar), .A2(n635bar), .ZN(n644bar) );
  OR2_X1 U334 ( .A1(n634), .A2(n633), .ZN(n635) );
  AND2_X1 U334bar ( .A1(n634bar), .A2(n633bar), .ZN(n635bar) );
  OR2_X1 U335 ( .A1(in[239]), .A2(in[218]), .ZN(n633) );
  AND2_X1 U335bar ( .A1(inbar[239]), .A2(inbar[218]), .ZN(n633bar) );
  OR2_X1 U336 ( .A1(in_13), .A2(in[87]), .ZN(n634) );
  AND2_X1 U336bar ( .A1(in_13bar), .A2(inbar[87]), .ZN(n634bar) );
  OR2_X1 U337 ( .A1(n632), .A2(n631), .ZN(n636) );
  AND2_X1 U337bar ( .A1(n632bar), .A2(n631bar), .ZN(n636bar) );
  OR2_X1 U338 ( .A1(in_72), .A2(in_70), .ZN(n631) );
  AND2_X1 U338bar ( .A1(in_72bar), .A2(in_70bar), .ZN(n631bar) );
  OR2_X1 U339 ( .A1(in_80), .A2(in_74), .ZN(n632) );
  AND2_X1 U339bar ( .A1(in_80bar), .A2(in_74bar), .ZN(n632bar) );
  OR2_X1 U340 ( .A1(n630), .A2(n629), .ZN(n942) );
  AND2_X1 U340bar ( .A1(n630bar), .A2(n629bar), .ZN(n942bar) );
  OR2_X1 U341 ( .A1(n628), .A2(n627), .ZN(n629) );
  AND2_X1 U341bar ( .A1(n628bar), .A2(n627bar), .ZN(n629bar) );
  OR2_X1 U342 ( .A1(n626), .A2(n625), .ZN(n627) );
  AND2_X1 U342bar ( .A1(n626bar), .A2(n625bar), .ZN(n627bar) );
  OR2_X1 U343 ( .A1(in[146]), .A2(in[100]), .ZN(n625) );
  AND2_X1 U343bar ( .A1(inbar[146]), .A2(inbar[100]), .ZN(n625bar) );
  OR2_X1 U344 ( .A1(in[168]), .A2(in[152]), .ZN(n626) );
  AND2_X1 U344bar ( .A1(inbar[168]), .A2(inbar[152]), .ZN(n626bar) );
  OR2_X1 U345 ( .A1(n624), .A2(n623), .ZN(n628) );
  AND2_X1 U345bar ( .A1(n624bar), .A2(n623bar), .ZN(n628bar) );
  OR2_X1 U346 ( .A1(in[199]), .A2(in[182]), .ZN(n623) );
  AND2_X1 U346bar ( .A1(inbar[199]), .A2(inbar[182]), .ZN(n623bar) );
  OR2_X1 U347 ( .A1(in[236]), .A2(in[204]), .ZN(n624) );
  AND2_X1 U347bar ( .A1(inbar[236]), .A2(inbar[204]), .ZN(n624bar) );
  OR2_X1 U348 ( .A1(n622), .A2(n621), .ZN(n630) );
  AND2_X1 U348bar ( .A1(n622bar), .A2(n621bar), .ZN(n630bar) );
  OR2_X1 U349 ( .A1(n620), .A2(n619), .ZN(n621) );
  AND2_X1 U349bar ( .A1(n620bar), .A2(n619bar), .ZN(n621bar) );
  OR2_X1 U350 ( .A1(in[89]), .A2(in[246]), .ZN(n619) );
  AND2_X1 U350bar ( .A1(inbar[89]), .A2(inbar[246]), .ZN(n619bar) );
  OR2_X1 U351 ( .A1(in[95]), .A2(in[92]), .ZN(n620) );
  AND2_X1 U351bar ( .A1(inbar[95]), .A2(inbar[92]), .ZN(n620bar) );
  OR2_X1 U352 ( .A1(n618), .A2(n617), .ZN(n622) );
  AND2_X1 U352bar ( .A1(n618bar), .A2(n617bar), .ZN(n622bar) );
  OR2_X1 U353 ( .A1(in_22), .A2(in_16), .ZN(n617) );
  AND2_X1 U353bar ( .A1(in_22bar), .A2(in_16bar), .ZN(n617bar) );
  OR2_X1 U354 ( .A1(in_51), .A2(in_49), .ZN(n618) );
  AND2_X1 U354bar ( .A1(in_51bar), .A2(in_49bar), .ZN(n618bar) );
  OR2_X1 U355 ( .A1(n616), .A2(n615), .ZN(n722) );
  AND2_X1 U355bar ( .A1(n616bar), .A2(n615bar), .ZN(n722bar) );
  OR2_X1 U356 ( .A1(in[158]), .A2(in[115]), .ZN(n615) );
  AND2_X1 U356bar ( .A1(inbar[158]), .A2(inbar[115]), .ZN(n615bar) );
  OR2_X1 U357 ( .A1(in[163]), .A2(n614), .ZN(n616) );
  AND2_X1 U357bar ( .A1(inbar[163]), .A2(n614bar), .ZN(n616bar) );
  OR2_X1 U358 ( .A1(in[206]), .A2(in[165]), .ZN(n614) );
  AND2_X1 U358bar ( .A1(inbar[206]), .A2(inbar[165]), .ZN(n614bar) );
  OR2_X1 U359 ( .A1(n613), .A2(n612), .ZN(n724) );
  AND2_X1 U359bar ( .A1(n613bar), .A2(n612bar), .ZN(n724bar) );
  OR2_X1 U360 ( .A1(n611), .A2(n610), .ZN(n612) );
  AND2_X1 U360bar ( .A1(n611bar), .A2(n610bar), .ZN(n612bar) );
  OR2_X1 U361 ( .A1(in[213]), .A2(in[207]), .ZN(n610) );
  AND2_X1 U361bar ( .A1(inbar[213]), .A2(inbar[207]), .ZN(n610bar) );
  OR2_X1 U362 ( .A1(in[215]), .A2(n609), .ZN(n611) );
  AND2_X1 U362bar ( .A1(inbar[215]), .A2(n609bar), .ZN(n611bar) );
  OR2_X1 U363 ( .A1(in[230]), .A2(in[220]), .ZN(n609) );
  AND2_X1 U363bar ( .A1(inbar[230]), .A2(inbar[220]), .ZN(n609bar) );
  OR2_X1 U364 ( .A1(n608), .A2(n607), .ZN(n613) );
  AND2_X1 U364bar ( .A1(n608bar), .A2(n607bar), .ZN(n613bar) );
  OR2_X1 U365 ( .A1(in[251]), .A2(in[234]), .ZN(n607) );
  AND2_X1 U365bar ( .A1(inbar[251]), .A2(inbar[234]), .ZN(n607bar) );
  OR2_X1 U366 ( .A1(in_17), .A2(n606), .ZN(n608) );
  AND2_X1 U366bar ( .A1(in_17bar), .A2(n606bar), .ZN(n608bar) );
  OR2_X1 U367 ( .A1(in_65), .A2(in_56), .ZN(n606) );
  AND2_X1 U367bar ( .A1(in_65bar), .A2(in_56bar), .ZN(n606bar) );
  OR2_X1 U368 ( .A1(n605), .A2(n604), .ZN(out[0]) );
  AND2_X1 U368bar ( .A1(n605bar), .A2(n604bar), .ZN(outbar[0]) );
  OR2_X1 U369 ( .A1(n603), .A2(n602), .ZN(n604) );
  AND2_X1 U369bar ( .A1(n603bar), .A2(n602bar), .ZN(n604bar) );
  OR2_X1 U370 ( .A1(n601), .A2(n600), .ZN(n602) );
  AND2_X1 U370bar ( .A1(n601bar), .A2(n600bar), .ZN(n602bar) );
  OR2_X1 U371 ( .A1(n820), .A2(n785), .ZN(n600) );
  AND2_X1 U371bar ( .A1(n820bar), .A2(n785bar), .ZN(n600bar) );
  OR2_X1 U372 ( .A1(n599), .A2(n598), .ZN(n785) );
  AND2_X1 U372bar ( .A1(n599bar), .A2(n598bar), .ZN(n785bar) );
  OR2_X1 U373 ( .A1(n597), .A2(n596), .ZN(n598) );
  AND2_X1 U373bar ( .A1(n597bar), .A2(n596bar), .ZN(n598bar) );
  OR2_X1 U374 ( .A1(n595), .A2(n594), .ZN(n596) );
  AND2_X1 U374bar ( .A1(n595bar), .A2(n594bar), .ZN(n596bar) );
  OR2_X1 U375 ( .A1(in[135]), .A2(in[104]), .ZN(n594) );
  AND2_X1 U375bar ( .A1(inbar[135]), .A2(inbar[104]), .ZN(n594bar) );
  OR2_X1 U376 ( .A1(in[188]), .A2(in[178]), .ZN(n595) );
  AND2_X1 U376bar ( .A1(inbar[188]), .A2(inbar[178]), .ZN(n595bar) );
  OR2_X1 U377 ( .A1(n593), .A2(n592), .ZN(n597) );
  AND2_X1 U377bar ( .A1(n593bar), .A2(n592bar), .ZN(n597bar) );
  OR2_X1 U378 ( .A1(in[217]), .A2(in[194]), .ZN(n592) );
  AND2_X1 U378bar ( .A1(inbar[217]), .A2(inbar[194]), .ZN(n592bar) );
  OR2_X1 U379 ( .A1(in[237]), .A2(in[218]), .ZN(n593) );
  AND2_X1 U379bar ( .A1(inbar[237]), .A2(inbar[218]), .ZN(n593bar) );
  OR2_X1 U380 ( .A1(n591), .A2(n590), .ZN(n599) );
  AND2_X1 U380bar ( .A1(n591bar), .A2(n590bar), .ZN(n599bar) );
  OR2_X1 U381 ( .A1(n589), .A2(n588), .ZN(n590) );
  AND2_X1 U381bar ( .A1(n589bar), .A2(n588bar), .ZN(n590bar) );
  OR2_X1 U382 ( .A1(in_2), .A2(in_10), .ZN(n588) );
  AND2_X1 U382bar ( .A1(in_2bar), .A2(in_10bar), .ZN(n588bar) );
  OR2_X1 U383 ( .A1(in_47), .A2(in_22), .ZN(n589) );
  AND2_X1 U383bar ( .A1(in_47bar), .A2(in_22bar), .ZN(n589bar) );
  OR2_X1 U384 ( .A1(n587), .A2(n586), .ZN(n591) );
  AND2_X1 U384bar ( .A1(n587bar), .A2(n586bar), .ZN(n591bar) );
  OR2_X1 U385 ( .A1(in_56), .A2(in_54), .ZN(n586) );
  AND2_X1 U385bar ( .A1(in_56bar), .A2(in_54bar), .ZN(n586bar) );
  OR2_X1 U386 ( .A1(in_63), .A2(in_61), .ZN(n587) );
  AND2_X1 U386bar ( .A1(in_63bar), .A2(in_61bar), .ZN(n587bar) );
  OR2_X1 U387 ( .A1(n585), .A2(n584), .ZN(n820) );
  AND2_X1 U387bar ( .A1(n585bar), .A2(n584bar), .ZN(n820bar) );
  OR2_X1 U388 ( .A1(n583), .A2(n582), .ZN(n584) );
  AND2_X1 U388bar ( .A1(n583bar), .A2(n582bar), .ZN(n584bar) );
  OR2_X1 U389 ( .A1(n581), .A2(n580), .ZN(n582) );
  AND2_X1 U389bar ( .A1(n581bar), .A2(n580bar), .ZN(n582bar) );
  OR2_X1 U390 ( .A1(in[158]), .A2(in[142]), .ZN(n580) );
  AND2_X1 U390bar ( .A1(inbar[158]), .A2(inbar[142]), .ZN(n580bar) );
  OR2_X1 U391 ( .A1(in[175]), .A2(in[164]), .ZN(n581) );
  AND2_X1 U391bar ( .A1(inbar[175]), .A2(inbar[164]), .ZN(n581bar) );
  OR2_X1 U392 ( .A1(n579), .A2(n578), .ZN(n583) );
  AND2_X1 U392bar ( .A1(n579bar), .A2(n578bar), .ZN(n583bar) );
  OR2_X1 U393 ( .A1(in[228]), .A2(in[204]), .ZN(n578) );
  AND2_X1 U393bar ( .A1(inbar[228]), .A2(inbar[204]), .ZN(n578bar) );
  OR2_X1 U394 ( .A1(in[91]), .A2(in[87]), .ZN(n579) );
  AND2_X1 U394bar ( .A1(inbar[91]), .A2(inbar[87]), .ZN(n579bar) );
  OR2_X1 U395 ( .A1(n577), .A2(n576), .ZN(n585) );
  AND2_X1 U395bar ( .A1(n577bar), .A2(n576bar), .ZN(n585bar) );
  OR2_X1 U396 ( .A1(n575), .A2(n574), .ZN(n576) );
  AND2_X1 U396bar ( .A1(n575bar), .A2(n574bar), .ZN(n576bar) );
  OR2_X1 U397 ( .A1(in_21), .A2(in_11), .ZN(n574) );
  AND2_X1 U397bar ( .A1(in_21bar), .A2(in_11bar), .ZN(n574bar) );
  OR2_X1 U398 ( .A1(in_5), .A2(in_3), .ZN(n575) );
  AND2_X1 U398bar ( .A1(in_5bar), .A2(in_3bar), .ZN(n575bar) );
  OR2_X1 U399 ( .A1(n573), .A2(n572), .ZN(n577) );
  AND2_X1 U399bar ( .A1(n573bar), .A2(n572bar), .ZN(n577bar) );
  OR2_X1 U400 ( .A1(in_68), .A2(in_64), .ZN(n572) );
  AND2_X1 U400bar ( .A1(in_68bar), .A2(in_64bar), .ZN(n572bar) );
  OR2_X1 U401 ( .A1(in_76), .A2(in_73), .ZN(n573) );
  AND2_X1 U401bar ( .A1(in_76bar), .A2(in_73bar), .ZN(n573bar) );
  OR2_X1 U402 ( .A1(n778), .A2(n571), .ZN(n601) );
  AND2_X1 U402bar ( .A1(n778bar), .A2(n571bar), .ZN(n601bar) );
  OR2_X1 U403 ( .A1(in[100]), .A2(n965), .ZN(n571) );
  AND2_X1 U403bar ( .A1(inbar[100]), .A2(n965bar), .ZN(n571bar) );
  OR2_X1 U404 ( .A1(n570), .A2(n569), .ZN(n965) );
  AND2_X1 U404bar ( .A1(n570bar), .A2(n569bar), .ZN(n965bar) );
  OR2_X1 U405 ( .A1(n568), .A2(n567), .ZN(n569) );
  AND2_X1 U405bar ( .A1(n568bar), .A2(n567bar), .ZN(n569bar) );
  OR2_X1 U406 ( .A1(n566), .A2(n565), .ZN(n567) );
  AND2_X1 U406bar ( .A1(n566bar), .A2(n565bar), .ZN(n567bar) );
  OR2_X1 U407 ( .A1(n817), .A2(n750), .ZN(n565) );
  AND2_X1 U407bar ( .A1(n817bar), .A2(n750bar), .ZN(n565bar) );
  OR2_X1 U408 ( .A1(n564), .A2(n563), .ZN(n750) );
  AND2_X1 U408bar ( .A1(n564bar), .A2(n563bar), .ZN(n750bar) );
  OR2_X1 U409 ( .A1(n562), .A2(n561), .ZN(n563) );
  AND2_X1 U409bar ( .A1(n562bar), .A2(n561bar), .ZN(n563bar) );
  OR2_X1 U410 ( .A1(n560), .A2(n559), .ZN(n561) );
  AND2_X1 U410bar ( .A1(n560bar), .A2(n559bar), .ZN(n561bar) );
  OR2_X1 U411 ( .A1(in[119]), .A2(in[103]), .ZN(n559) );
  AND2_X1 U411bar ( .A1(inbar[119]), .A2(inbar[103]), .ZN(n559bar) );
  OR2_X1 U412 ( .A1(in[137]), .A2(in[133]), .ZN(n560) );
  AND2_X1 U412bar ( .A1(inbar[137]), .A2(inbar[133]), .ZN(n560bar) );
  OR2_X1 U413 ( .A1(n558), .A2(n557), .ZN(n562) );
  AND2_X1 U413bar ( .A1(n558bar), .A2(n557bar), .ZN(n562bar) );
  OR2_X1 U414 ( .A1(in[176]), .A2(in[173]), .ZN(n557) );
  AND2_X1 U414bar ( .A1(inbar[176]), .A2(inbar[173]), .ZN(n557bar) );
  OR2_X1 U415 ( .A1(in[210]), .A2(in[181]), .ZN(n558) );
  AND2_X1 U415bar ( .A1(inbar[210]), .A2(inbar[181]), .ZN(n558bar) );
  OR2_X1 U416 ( .A1(n556), .A2(n555), .ZN(n564) );
  AND2_X1 U416bar ( .A1(n556bar), .A2(n555bar), .ZN(n564bar) );
  OR2_X1 U417 ( .A1(n554), .A2(n553), .ZN(n555) );
  AND2_X1 U417bar ( .A1(n554bar), .A2(n553bar), .ZN(n555bar) );
  OR2_X1 U418 ( .A1(in_13), .A2(in[234]), .ZN(n553) );
  AND2_X1 U418bar ( .A1(in_13bar), .A2(inbar[234]), .ZN(n553bar) );
  OR2_X1 U419 ( .A1(in_38), .A2(in_32), .ZN(n554) );
  AND2_X1 U419bar ( .A1(in_38bar), .A2(in_32bar), .ZN(n554bar) );
  OR2_X1 U420 ( .A1(n552), .A2(n551), .ZN(n556) );
  AND2_X1 U420bar ( .A1(n552bar), .A2(n551bar), .ZN(n556bar) );
  OR2_X1 U421 ( .A1(in_42), .A2(in_41), .ZN(n551) );
  AND2_X1 U421bar ( .A1(in_42bar), .A2(in_41bar), .ZN(n551bar) );
  OR2_X1 U422 ( .A1(in_7), .A2(in_49), .ZN(n552) );
  AND2_X1 U422bar ( .A1(in_7bar), .A2(in_49bar), .ZN(n552bar) );
  OR2_X1 U423 ( .A1(n550), .A2(n549), .ZN(n817) );
  AND2_X1 U423bar ( .A1(n550bar), .A2(n549bar), .ZN(n817bar) );
  OR2_X1 U424 ( .A1(n548), .A2(n547), .ZN(n549) );
  AND2_X1 U424bar ( .A1(n548bar), .A2(n547bar), .ZN(n549bar) );
  OR2_X1 U425 ( .A1(n546), .A2(n545), .ZN(n547) );
  AND2_X1 U425bar ( .A1(n546bar), .A2(n545bar), .ZN(n547bar) );
  OR2_X1 U426 ( .A1(in[159]), .A2(in[105]), .ZN(n545) );
  AND2_X1 U426bar ( .A1(inbar[159]), .A2(inbar[105]), .ZN(n545bar) );
  OR2_X1 U427 ( .A1(in[206]), .A2(in[183]), .ZN(n546) );
  AND2_X1 U427bar ( .A1(inbar[206]), .A2(inbar[183]), .ZN(n546bar) );
  OR2_X1 U428 ( .A1(n544), .A2(n543), .ZN(n548) );
  AND2_X1 U428bar ( .A1(n544bar), .A2(n543bar), .ZN(n548bar) );
  OR2_X1 U429 ( .A1(in[229]), .A2(in[219]), .ZN(n543) );
  AND2_X1 U429bar ( .A1(inbar[229]), .A2(inbar[219]), .ZN(n543bar) );
  OR2_X1 U430 ( .A1(in[235]), .A2(in[232]), .ZN(n544) );
  AND2_X1 U430bar ( .A1(inbar[235]), .A2(inbar[232]), .ZN(n544bar) );
  OR2_X1 U431 ( .A1(n542), .A2(n541), .ZN(n550) );
  AND2_X1 U431bar ( .A1(n542bar), .A2(n541bar), .ZN(n550bar) );
  OR2_X1 U432 ( .A1(n540), .A2(n539), .ZN(n541) );
  AND2_X1 U432bar ( .A1(n540bar), .A2(n539bar), .ZN(n541bar) );
  OR2_X1 U433 ( .A1(in[249]), .A2(in[242]), .ZN(n539) );
  AND2_X1 U433bar ( .A1(inbar[249]), .A2(inbar[242]), .ZN(n539bar) );
  OR2_X1 U434 ( .A1(in[89]), .A2(in[254]), .ZN(n540) );
  AND2_X1 U434bar ( .A1(inbar[89]), .A2(inbar[254]), .ZN(n540bar) );
  OR2_X1 U435 ( .A1(n538), .A2(n537), .ZN(n542) );
  AND2_X1 U435bar ( .A1(n538bar), .A2(n537bar), .ZN(n542bar) );
  OR2_X1 U436 ( .A1(in_14), .A2(in[99]), .ZN(n537) );
  AND2_X1 U436bar ( .A1(in_14bar), .A2(inbar[99]), .ZN(n537bar) );
  OR2_X1 U437 ( .A1(in_60), .A2(in_18), .ZN(n538) );
  AND2_X1 U437bar ( .A1(in_60bar), .A2(in_18bar), .ZN(n538bar) );
  OR2_X1 U438 ( .A1(in[113]), .A2(n763), .ZN(n566) );
  AND2_X1 U438bar ( .A1(inbar[113]), .A2(n763bar), .ZN(n566bar) );
  OR2_X1 U439 ( .A1(n536), .A2(n535), .ZN(n763) );
  AND2_X1 U439bar ( .A1(n536bar), .A2(n535bar), .ZN(n763bar) );
  OR2_X1 U440 ( .A1(n534), .A2(n533), .ZN(n535) );
  AND2_X1 U440bar ( .A1(n534bar), .A2(n533bar), .ZN(n535bar) );
  OR2_X1 U441 ( .A1(n532), .A2(n531), .ZN(n533) );
  AND2_X1 U441bar ( .A1(n532bar), .A2(n531bar), .ZN(n533bar) );
  OR2_X1 U442 ( .A1(in[115]), .A2(in[110]), .ZN(n531) );
  AND2_X1 U442bar ( .A1(inbar[115]), .A2(inbar[110]), .ZN(n531bar) );
  OR2_X1 U443 ( .A1(in[125]), .A2(in[117]), .ZN(n532) );
  AND2_X1 U443bar ( .A1(inbar[125]), .A2(inbar[117]), .ZN(n532bar) );
  OR2_X1 U444 ( .A1(n530), .A2(n529), .ZN(n534) );
  AND2_X1 U444bar ( .A1(n530bar), .A2(n529bar), .ZN(n534bar) );
  OR2_X1 U445 ( .A1(in[180]), .A2(in[128]), .ZN(n529) );
  AND2_X1 U445bar ( .A1(inbar[180]), .A2(inbar[128]), .ZN(n529bar) );
  OR2_X1 U446 ( .A1(in[205]), .A2(in[201]), .ZN(n530) );
  AND2_X1 U446bar ( .A1(inbar[205]), .A2(inbar[201]), .ZN(n530bar) );
  OR2_X1 U447 ( .A1(n528), .A2(n527), .ZN(n536) );
  AND2_X1 U447bar ( .A1(n528bar), .A2(n527bar), .ZN(n536bar) );
  OR2_X1 U448 ( .A1(n526), .A2(n525), .ZN(n527) );
  AND2_X1 U448bar ( .A1(n526bar), .A2(n525bar), .ZN(n527bar) );
  OR2_X1 U449 ( .A1(in[244]), .A2(in[239]), .ZN(n525) );
  AND2_X1 U449bar ( .A1(inbar[244]), .A2(inbar[239]), .ZN(n525bar) );
  OR2_X1 U450 ( .A1(in[95]), .A2(in[83]), .ZN(n526) );
  AND2_X1 U450bar ( .A1(inbar[95]), .A2(inbar[83]), .ZN(n526bar) );
  OR2_X1 U451 ( .A1(n524), .A2(n523), .ZN(n528) );
  AND2_X1 U451bar ( .A1(n524bar), .A2(n523bar), .ZN(n528bar) );
  OR2_X1 U452 ( .A1(in_24), .A2(in[97]), .ZN(n523) );
  AND2_X1 U452bar ( .A1(in_24bar), .A2(inbar[97]), .ZN(n523bar) );
  OR2_X1 U453 ( .A1(in_33), .A2(in_27), .ZN(n524) );
  AND2_X1 U453bar ( .A1(in_33bar), .A2(in_27bar), .ZN(n524bar) );
  OR2_X1 U454 ( .A1(n522), .A2(n521), .ZN(n568) );
  AND2_X1 U454bar ( .A1(n522bar), .A2(n521bar), .ZN(n568bar) );
  OR2_X1 U455 ( .A1(in[145]), .A2(in[126]), .ZN(n521) );
  AND2_X1 U455bar ( .A1(inbar[145]), .A2(inbar[126]), .ZN(n521bar) );
  OR2_X1 U456 ( .A1(in[169]), .A2(n520), .ZN(n522) );
  AND2_X1 U456bar ( .A1(inbar[169]), .A2(n520bar), .ZN(n522bar) );
  OR2_X1 U457 ( .A1(in[221]), .A2(in[172]), .ZN(n520) );
  AND2_X1 U457bar ( .A1(inbar[221]), .A2(inbar[172]), .ZN(n520bar) );
  OR2_X1 U458 ( .A1(n519), .A2(n518), .ZN(n570) );
  AND2_X1 U458bar ( .A1(n519bar), .A2(n518bar), .ZN(n570bar) );
  OR2_X1 U459 ( .A1(n517), .A2(n516), .ZN(n518) );
  AND2_X1 U459bar ( .A1(n517bar), .A2(n516bar), .ZN(n518bar) );
  OR2_X1 U460 ( .A1(in[241]), .A2(in[224]), .ZN(n516) );
  AND2_X1 U460bar ( .A1(inbar[241]), .A2(inbar[224]), .ZN(n516bar) );
  OR2_X1 U461 ( .A1(in[86]), .A2(n515), .ZN(n517) );
  AND2_X1 U461bar ( .A1(inbar[86]), .A2(n515bar), .ZN(n517bar) );
  OR2_X1 U462 ( .A1(in_43), .A2(in_34), .ZN(n515) );
  AND2_X1 U462bar ( .A1(in_43bar), .A2(in_34bar), .ZN(n515bar) );
  OR2_X1 U463 ( .A1(n514), .A2(n513), .ZN(n519) );
  AND2_X1 U463bar ( .A1(n514bar), .A2(n513bar), .ZN(n519bar) );
  OR2_X1 U464 ( .A1(in_65), .A2(in_51), .ZN(n513) );
  AND2_X1 U464bar ( .A1(in_65bar), .A2(in_51bar), .ZN(n513bar) );
  OR2_X1 U465 ( .A1(in_75), .A2(n512), .ZN(n514) );
  AND2_X1 U465bar ( .A1(in_75bar), .A2(n512bar), .ZN(n514bar) );
  OR2_X1 U466 ( .A1(in_81), .A2(in_77), .ZN(n512) );
  AND2_X1 U466bar ( .A1(in_81bar), .A2(in_77bar), .ZN(n512bar) );
  OR2_X1 U467 ( .A1(n511), .A2(n510), .ZN(n778) );
  AND2_X1 U467bar ( .A1(n511bar), .A2(n510bar), .ZN(n778bar) );
  OR2_X1 U468 ( .A1(n509), .A2(n508), .ZN(n510) );
  AND2_X1 U468bar ( .A1(n509bar), .A2(n508bar), .ZN(n510bar) );
  OR2_X1 U469 ( .A1(n507), .A2(n506), .ZN(n508) );
  AND2_X1 U469bar ( .A1(n507bar), .A2(n506bar), .ZN(n508bar) );
  OR2_X1 U470 ( .A1(in[107]), .A2(in[101]), .ZN(n506) );
  AND2_X1 U470bar ( .A1(inbar[107]), .A2(inbar[101]), .ZN(n506bar) );
  OR2_X1 U471 ( .A1(in[139]), .A2(in[132]), .ZN(n507) );
  AND2_X1 U471bar ( .A1(inbar[139]), .A2(inbar[132]), .ZN(n507bar) );
  OR2_X1 U472 ( .A1(n505), .A2(n504), .ZN(n509) );
  AND2_X1 U472bar ( .A1(n505bar), .A2(n504bar), .ZN(n509bar) );
  OR2_X1 U473 ( .A1(in[146]), .A2(in[141]), .ZN(n504) );
  AND2_X1 U473bar ( .A1(inbar[146]), .A2(inbar[141]), .ZN(n504bar) );
  OR2_X1 U474 ( .A1(in[203]), .A2(in[179]), .ZN(n505) );
  AND2_X1 U474bar ( .A1(inbar[203]), .A2(inbar[179]), .ZN(n505bar) );
  OR2_X1 U475 ( .A1(n503), .A2(n502), .ZN(n511) );
  AND2_X1 U475bar ( .A1(n503bar), .A2(n502bar), .ZN(n511bar) );
  OR2_X1 U476 ( .A1(n501), .A2(n500), .ZN(n502) );
  AND2_X1 U476bar ( .A1(n501bar), .A2(n500bar), .ZN(n502bar) );
  OR2_X1 U477 ( .A1(in[243]), .A2(in[222]), .ZN(n500) );
  AND2_X1 U477bar ( .A1(inbar[243]), .A2(inbar[222]), .ZN(n500bar) );
  OR2_X1 U478 ( .A1(in[251]), .A2(in[250]), .ZN(n501) );
  AND2_X1 U478bar ( .A1(inbar[251]), .A2(inbar[250]), .ZN(n501bar) );
  OR2_X1 U479 ( .A1(n499), .A2(n498), .ZN(n503) );
  AND2_X1 U479bar ( .A1(n499bar), .A2(n498bar), .ZN(n503bar) );
  OR2_X1 U480 ( .A1(in_37), .A2(in_19), .ZN(n498) );
  AND2_X1 U480bar ( .A1(in_37bar), .A2(in_19bar), .ZN(n498bar) );
  OR2_X1 U481 ( .A1(in_78), .A2(in_6), .ZN(n499) );
  AND2_X1 U481bar ( .A1(in_78bar), .A2(in_6bar), .ZN(n499bar) );
  OR2_X1 U482 ( .A1(n497), .A2(n496), .ZN(n603) );
  AND2_X1 U482bar ( .A1(n497bar), .A2(n496bar), .ZN(n603bar) );
  OR2_X1 U483 ( .A1(in[112]), .A2(in[102]), .ZN(n496) );
  AND2_X1 U483bar ( .A1(inbar[112]), .A2(inbar[102]), .ZN(n496bar) );
  OR2_X1 U484 ( .A1(in[123]), .A2(n495), .ZN(n497) );
  AND2_X1 U484bar ( .A1(inbar[123]), .A2(n495bar), .ZN(n497bar) );
  OR2_X1 U485 ( .A1(in[143]), .A2(in[130]), .ZN(n495) );
  AND2_X1 U485bar ( .A1(inbar[143]), .A2(inbar[130]), .ZN(n495bar) );
  OR2_X1 U486 ( .A1(n494), .A2(n493), .ZN(n605) );
  AND2_X1 U486bar ( .A1(n494bar), .A2(n493bar), .ZN(n605bar) );
  OR2_X1 U487 ( .A1(n492), .A2(n491), .ZN(n493) );
  AND2_X1 U487bar ( .A1(n492bar), .A2(n491bar), .ZN(n493bar) );
  OR2_X1 U488 ( .A1(in[216]), .A2(in[213]), .ZN(n491) );
  AND2_X1 U488bar ( .A1(inbar[216]), .A2(inbar[213]), .ZN(n491bar) );
  OR2_X1 U489 ( .A1(in[227]), .A2(n490), .ZN(n492) );
  AND2_X1 U489bar ( .A1(inbar[227]), .A2(n490bar), .ZN(n492bar) );
  OR2_X1 U490 ( .A1(in_0), .A2(in[248]), .ZN(n490) );
  AND2_X1 U490bar ( .A1(in_0bar), .A2(inbar[248]), .ZN(n490bar) );
  OR2_X1 U491 ( .A1(n489), .A2(n488), .ZN(n494) );
  AND2_X1 U491bar ( .A1(n489bar), .A2(n488bar), .ZN(n494bar) );
  OR2_X1 U492 ( .A1(in_46), .A2(in_44), .ZN(n488) );
  AND2_X1 U492bar ( .A1(in_46bar), .A2(in_44bar), .ZN(n488bar) );
  OR2_X1 U493 ( .A1(in_50), .A2(n487), .ZN(n489) );
  AND2_X1 U493bar ( .A1(in_50bar), .A2(n487bar), .ZN(n489bar) );
  OR2_X1 U494 ( .A1(in_9), .A2(in_80), .ZN(n487) );
  AND2_X1 U494bar ( .A1(in_9bar), .A2(in_80bar), .ZN(n487bar) );
endmodule

module sBox_13 ( in, inbar, out, outbar );

  input wire [7:0] in;
  input wire [7:0] inbar;
//input_done

  output wire [7:0] out;
  output wire [7:0] outbar;
//output_done

  wire [255:0] decodeOut;
  wire [255:0] decodeOutbar;
//wire_done

  decode_13 dec ( .in(in), .inbar(inbar), .out(decodeOut), .outbar(decodeOutbar) );
  encode_13 enc ( .in(decodeOut), .inbar(decodeOutbar), .out(out), .outbar(outbar) );
endmodule

module CD2_53 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD2_54 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD2_55 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD2_56 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD4_27 ( a, abar, b, bbar, y, ybar );

  input wire [3:0] a;
  input wire [3:0] b;
  input wire [3:0] abar;
  input wire [3:0] bbar;
//input_done

  output wire [15:0] y;
  output wire [15:0] ybar;
//output_done

//wire_done

  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]) );
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]) );
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]) );
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]) );
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]) );
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]) );
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]) );
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]) );
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]) );
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]) );
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]) );
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]) );
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]) );
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]) );
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]) );
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]) );
endmodule

module CD4_28 ( a, abar, b, bbar, y, ybar );

  input wire [3:0] a;
  input wire [3:0] b;
  input wire [3:0] abar;
  input wire [3:0] bbar;
//input_done

  output wire [15:0] y;
  output wire [15:0] ybar;
//output_done

//wire_done

  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]) );
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]) );
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]) );
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]) );
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]) );
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]) );
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]) );
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]) );
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]) );
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]) );
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]) );
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]) );
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]) );
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]) );
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]) );
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]) );
endmodule

module CD16_14 ( a, abar, b, bbar, y, ybar );

  input wire [15:0] a;
  input wire [15:0] b;
  input wire [15:0] abar;
  input wire [15:0] bbar;
//input_done

  output wire [255:0] y;
  output wire [255:0] ybar;
//output_done

//wire_done

  AND2_X1 U1 ( .A1(b[9]), .A2(a[0]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[9]), .A2(abar[0]), .ZN(ybar[9]) );
  AND2_X1 U2 ( .A1(b[3]), .A2(a[6]), .ZN(y[99]) );
  OR2_X1 U2bar ( .A1(bbar[3]), .A2(abar[6]), .ZN(ybar[99]) );
  AND2_X1 U3 ( .A1(b[2]), .A2(a[6]), .ZN(y[98]) );
  OR2_X1 U3bar ( .A1(bbar[2]), .A2(abar[6]), .ZN(ybar[98]) );
  AND2_X1 U4 ( .A1(b[1]), .A2(a[6]), .ZN(y[97]) );
  OR2_X1 U4bar ( .A1(bbar[1]), .A2(abar[6]), .ZN(ybar[97]) );
  AND2_X1 U5 ( .A1(b[0]), .A2(a[6]), .ZN(y[96]) );
  OR2_X1 U5bar ( .A1(bbar[0]), .A2(abar[6]), .ZN(ybar[96]) );
  AND2_X1 U6 ( .A1(b[15]), .A2(a[5]), .ZN(y[95]) );
  OR2_X1 U6bar ( .A1(bbar[15]), .A2(abar[5]), .ZN(ybar[95]) );
  AND2_X1 U7 ( .A1(b[14]), .A2(a[5]), .ZN(y[94]) );
  OR2_X1 U7bar ( .A1(bbar[14]), .A2(abar[5]), .ZN(ybar[94]) );
  AND2_X1 U8 ( .A1(b[13]), .A2(a[5]), .ZN(y[93]) );
  OR2_X1 U8bar ( .A1(bbar[13]), .A2(abar[5]), .ZN(ybar[93]) );
  AND2_X1 U9 ( .A1(b[12]), .A2(a[5]), .ZN(y[92]) );
  OR2_X1 U9bar ( .A1(bbar[12]), .A2(abar[5]), .ZN(ybar[92]) );
  AND2_X1 U10 ( .A1(b[11]), .A2(a[5]), .ZN(y[91]) );
  OR2_X1 U10bar ( .A1(bbar[11]), .A2(abar[5]), .ZN(ybar[91]) );
  AND2_X1 U11 ( .A1(b[10]), .A2(a[5]), .ZN(y[90]) );
  OR2_X1 U11bar ( .A1(bbar[10]), .A2(abar[5]), .ZN(ybar[90]) );
  AND2_X1 U12 ( .A1(b[8]), .A2(a[0]), .ZN(y[8]) );
  OR2_X1 U12bar ( .A1(bbar[8]), .A2(abar[0]), .ZN(ybar[8]) );
  AND2_X1 U13 ( .A1(a[5]), .A2(b[9]), .ZN(y[89]) );
  OR2_X1 U13bar ( .A1(abar[5]), .A2(bbar[9]), .ZN(ybar[89]) );
  AND2_X1 U14 ( .A1(b[8]), .A2(a[5]), .ZN(y[88]) );
  OR2_X1 U14bar ( .A1(bbar[8]), .A2(abar[5]), .ZN(ybar[88]) );
  AND2_X1 U15 ( .A1(b[7]), .A2(a[5]), .ZN(y[87]) );
  OR2_X1 U15bar ( .A1(bbar[7]), .A2(abar[5]), .ZN(ybar[87]) );
  AND2_X1 U16 ( .A1(b[6]), .A2(a[5]), .ZN(y[86]) );
  OR2_X1 U16bar ( .A1(bbar[6]), .A2(abar[5]), .ZN(ybar[86]) );
  AND2_X1 U17 ( .A1(b[5]), .A2(a[5]), .ZN(y[85]) );
  OR2_X1 U17bar ( .A1(bbar[5]), .A2(abar[5]), .ZN(ybar[85]) );
  AND2_X1 U18 ( .A1(b[4]), .A2(a[5]), .ZN(y[84]) );
  OR2_X1 U18bar ( .A1(bbar[4]), .A2(abar[5]), .ZN(ybar[84]) );
  AND2_X1 U19 ( .A1(a[5]), .A2(b[3]), .ZN(y[83]) );
  OR2_X1 U19bar ( .A1(abar[5]), .A2(bbar[3]), .ZN(ybar[83]) );
  AND2_X1 U20 ( .A1(a[5]), .A2(b[2]), .ZN(y[82]) );
  OR2_X1 U20bar ( .A1(abar[5]), .A2(bbar[2]), .ZN(ybar[82]) );
  AND2_X1 U21 ( .A1(a[5]), .A2(b[1]), .ZN(y[81]) );
  OR2_X1 U21bar ( .A1(abar[5]), .A2(bbar[1]), .ZN(ybar[81]) );
  AND2_X1 U22 ( .A1(a[5]), .A2(b[0]), .ZN(y[80]) );
  OR2_X1 U22bar ( .A1(abar[5]), .A2(bbar[0]), .ZN(ybar[80]) );
  AND2_X1 U23 ( .A1(b[7]), .A2(a[0]), .ZN(y[7]) );
  OR2_X1 U23bar ( .A1(bbar[7]), .A2(abar[0]), .ZN(ybar[7]) );
  AND2_X1 U24 ( .A1(a[4]), .A2(b[15]), .ZN(y[79]) );
  OR2_X1 U24bar ( .A1(abar[4]), .A2(bbar[15]), .ZN(ybar[79]) );
  AND2_X1 U25 ( .A1(a[4]), .A2(b[14]), .ZN(y[78]) );
  OR2_X1 U25bar ( .A1(abar[4]), .A2(bbar[14]), .ZN(ybar[78]) );
  AND2_X1 U26 ( .A1(a[4]), .A2(b[13]), .ZN(y[77]) );
  OR2_X1 U26bar ( .A1(abar[4]), .A2(bbar[13]), .ZN(ybar[77]) );
  AND2_X1 U27 ( .A1(a[4]), .A2(b[12]), .ZN(y[76]) );
  OR2_X1 U27bar ( .A1(abar[4]), .A2(bbar[12]), .ZN(ybar[76]) );
  AND2_X1 U28 ( .A1(a[4]), .A2(b[11]), .ZN(y[75]) );
  OR2_X1 U28bar ( .A1(abar[4]), .A2(bbar[11]), .ZN(ybar[75]) );
  AND2_X1 U29 ( .A1(a[4]), .A2(b[10]), .ZN(y[74]) );
  OR2_X1 U29bar ( .A1(abar[4]), .A2(bbar[10]), .ZN(ybar[74]) );
  AND2_X1 U30 ( .A1(a[4]), .A2(b[9]), .ZN(y[73]) );
  OR2_X1 U30bar ( .A1(abar[4]), .A2(bbar[9]), .ZN(ybar[73]) );
  AND2_X1 U31 ( .A1(a[4]), .A2(b[8]), .ZN(y[72]) );
  OR2_X1 U31bar ( .A1(abar[4]), .A2(bbar[8]), .ZN(ybar[72]) );
  AND2_X1 U32 ( .A1(a[4]), .A2(b[7]), .ZN(y[71]) );
  OR2_X1 U32bar ( .A1(abar[4]), .A2(bbar[7]), .ZN(ybar[71]) );
  AND2_X1 U33 ( .A1(a[4]), .A2(b[6]), .ZN(y[70]) );
  OR2_X1 U33bar ( .A1(abar[4]), .A2(bbar[6]), .ZN(ybar[70]) );
  AND2_X1 U34 ( .A1(b[6]), .A2(a[0]), .ZN(y[6]) );
  OR2_X1 U34bar ( .A1(bbar[6]), .A2(abar[0]), .ZN(ybar[6]) );
  AND2_X1 U35 ( .A1(a[4]), .A2(b[5]), .ZN(y[69]) );
  OR2_X1 U35bar ( .A1(abar[4]), .A2(bbar[5]), .ZN(ybar[69]) );
  AND2_X1 U36 ( .A1(a[4]), .A2(b[4]), .ZN(y[68]) );
  OR2_X1 U36bar ( .A1(abar[4]), .A2(bbar[4]), .ZN(ybar[68]) );
  AND2_X1 U37 ( .A1(a[4]), .A2(b[3]), .ZN(y[67]) );
  OR2_X1 U37bar ( .A1(abar[4]), .A2(bbar[3]), .ZN(ybar[67]) );
  AND2_X1 U38 ( .A1(a[4]), .A2(b[2]), .ZN(y[66]) );
  OR2_X1 U38bar ( .A1(abar[4]), .A2(bbar[2]), .ZN(ybar[66]) );
  AND2_X1 U39 ( .A1(a[4]), .A2(b[1]), .ZN(y[65]) );
  OR2_X1 U39bar ( .A1(abar[4]), .A2(bbar[1]), .ZN(ybar[65]) );
  AND2_X1 U40 ( .A1(a[4]), .A2(b[0]), .ZN(y[64]) );
  OR2_X1 U40bar ( .A1(abar[4]), .A2(bbar[0]), .ZN(ybar[64]) );
  AND2_X1 U41 ( .A1(a[3]), .A2(b[15]), .ZN(y[63]) );
  OR2_X1 U41bar ( .A1(abar[3]), .A2(bbar[15]), .ZN(ybar[63]) );
  AND2_X1 U42 ( .A1(a[3]), .A2(b[14]), .ZN(y[62]) );
  OR2_X1 U42bar ( .A1(abar[3]), .A2(bbar[14]), .ZN(ybar[62]) );
  AND2_X1 U43 ( .A1(a[3]), .A2(b[13]), .ZN(y[61]) );
  OR2_X1 U43bar ( .A1(abar[3]), .A2(bbar[13]), .ZN(ybar[61]) );
  AND2_X1 U44 ( .A1(a[3]), .A2(b[12]), .ZN(y[60]) );
  OR2_X1 U44bar ( .A1(abar[3]), .A2(bbar[12]), .ZN(ybar[60]) );
  AND2_X1 U45 ( .A1(b[5]), .A2(a[0]), .ZN(y[5]) );
  OR2_X1 U45bar ( .A1(bbar[5]), .A2(abar[0]), .ZN(ybar[5]) );
  AND2_X1 U46 ( .A1(a[3]), .A2(b[11]), .ZN(y[59]) );
  OR2_X1 U46bar ( .A1(abar[3]), .A2(bbar[11]), .ZN(ybar[59]) );
  AND2_X1 U47 ( .A1(a[3]), .A2(b[10]), .ZN(y[58]) );
  OR2_X1 U47bar ( .A1(abar[3]), .A2(bbar[10]), .ZN(ybar[58]) );
  AND2_X1 U48 ( .A1(a[3]), .A2(b[9]), .ZN(y[57]) );
  OR2_X1 U48bar ( .A1(abar[3]), .A2(bbar[9]), .ZN(ybar[57]) );
  AND2_X1 U49 ( .A1(a[3]), .A2(b[8]), .ZN(y[56]) );
  OR2_X1 U49bar ( .A1(abar[3]), .A2(bbar[8]), .ZN(ybar[56]) );
  AND2_X1 U50 ( .A1(a[3]), .A2(b[7]), .ZN(y[55]) );
  OR2_X1 U50bar ( .A1(abar[3]), .A2(bbar[7]), .ZN(ybar[55]) );
  AND2_X1 U51 ( .A1(a[3]), .A2(b[6]), .ZN(y[54]) );
  OR2_X1 U51bar ( .A1(abar[3]), .A2(bbar[6]), .ZN(ybar[54]) );
  AND2_X1 U52 ( .A1(a[3]), .A2(b[5]), .ZN(y[53]) );
  OR2_X1 U52bar ( .A1(abar[3]), .A2(bbar[5]), .ZN(ybar[53]) );
  AND2_X1 U53 ( .A1(a[3]), .A2(b[4]), .ZN(y[52]) );
  OR2_X1 U53bar ( .A1(abar[3]), .A2(bbar[4]), .ZN(ybar[52]) );
  AND2_X1 U54 ( .A1(a[3]), .A2(b[3]), .ZN(y[51]) );
  OR2_X1 U54bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[51]) );
  AND2_X1 U55 ( .A1(a[3]), .A2(b[2]), .ZN(y[50]) );
  OR2_X1 U55bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[50]) );
  AND2_X1 U56 ( .A1(b[4]), .A2(a[0]), .ZN(y[4]) );
  OR2_X1 U56bar ( .A1(bbar[4]), .A2(abar[0]), .ZN(ybar[4]) );
  AND2_X1 U57 ( .A1(a[3]), .A2(b[1]), .ZN(y[49]) );
  OR2_X1 U57bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[49]) );
  AND2_X1 U58 ( .A1(a[3]), .A2(b[0]), .ZN(y[48]) );
  OR2_X1 U58bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[48]) );
  AND2_X1 U59 ( .A1(a[2]), .A2(b[15]), .ZN(y[47]) );
  OR2_X1 U59bar ( .A1(abar[2]), .A2(bbar[15]), .ZN(ybar[47]) );
  AND2_X1 U60 ( .A1(a[2]), .A2(b[14]), .ZN(y[46]) );
  OR2_X1 U60bar ( .A1(abar[2]), .A2(bbar[14]), .ZN(ybar[46]) );
  AND2_X1 U61 ( .A1(a[2]), .A2(b[13]), .ZN(y[45]) );
  OR2_X1 U61bar ( .A1(abar[2]), .A2(bbar[13]), .ZN(ybar[45]) );
  AND2_X1 U62 ( .A1(a[2]), .A2(b[12]), .ZN(y[44]) );
  OR2_X1 U62bar ( .A1(abar[2]), .A2(bbar[12]), .ZN(ybar[44]) );
  AND2_X1 U63 ( .A1(a[2]), .A2(b[11]), .ZN(y[43]) );
  OR2_X1 U63bar ( .A1(abar[2]), .A2(bbar[11]), .ZN(ybar[43]) );
  AND2_X1 U64 ( .A1(a[2]), .A2(b[10]), .ZN(y[42]) );
  OR2_X1 U64bar ( .A1(abar[2]), .A2(bbar[10]), .ZN(ybar[42]) );
  AND2_X1 U65 ( .A1(a[2]), .A2(b[9]), .ZN(y[41]) );
  OR2_X1 U65bar ( .A1(abar[2]), .A2(bbar[9]), .ZN(ybar[41]) );
  AND2_X1 U66 ( .A1(a[2]), .A2(b[8]), .ZN(y[40]) );
  OR2_X1 U66bar ( .A1(abar[2]), .A2(bbar[8]), .ZN(ybar[40]) );
  AND2_X1 U67 ( .A1(b[3]), .A2(a[0]), .ZN(y[3]) );
  OR2_X1 U67bar ( .A1(bbar[3]), .A2(abar[0]), .ZN(ybar[3]) );
  AND2_X1 U68 ( .A1(a[2]), .A2(b[7]), .ZN(y[39]) );
  OR2_X1 U68bar ( .A1(abar[2]), .A2(bbar[7]), .ZN(ybar[39]) );
  AND2_X1 U69 ( .A1(a[2]), .A2(b[6]), .ZN(y[38]) );
  OR2_X1 U69bar ( .A1(abar[2]), .A2(bbar[6]), .ZN(ybar[38]) );
  AND2_X1 U70 ( .A1(a[2]), .A2(b[5]), .ZN(y[37]) );
  OR2_X1 U70bar ( .A1(abar[2]), .A2(bbar[5]), .ZN(ybar[37]) );
  AND2_X1 U71 ( .A1(a[2]), .A2(b[4]), .ZN(y[36]) );
  OR2_X1 U71bar ( .A1(abar[2]), .A2(bbar[4]), .ZN(ybar[36]) );
  AND2_X1 U72 ( .A1(a[2]), .A2(b[3]), .ZN(y[35]) );
  OR2_X1 U72bar ( .A1(abar[2]), .A2(bbar[3]), .ZN(ybar[35]) );
  AND2_X1 U73 ( .A1(a[2]), .A2(b[2]), .ZN(y[34]) );
  OR2_X1 U73bar ( .A1(abar[2]), .A2(bbar[2]), .ZN(ybar[34]) );
  AND2_X1 U74 ( .A1(a[2]), .A2(b[1]), .ZN(y[33]) );
  OR2_X1 U74bar ( .A1(abar[2]), .A2(bbar[1]), .ZN(ybar[33]) );
  AND2_X1 U75 ( .A1(a[2]), .A2(b[0]), .ZN(y[32]) );
  OR2_X1 U75bar ( .A1(abar[2]), .A2(bbar[0]), .ZN(ybar[32]) );
  AND2_X1 U76 ( .A1(a[1]), .A2(b[15]), .ZN(y[31]) );
  OR2_X1 U76bar ( .A1(abar[1]), .A2(bbar[15]), .ZN(ybar[31]) );
  AND2_X1 U77 ( .A1(a[1]), .A2(b[14]), .ZN(y[30]) );
  OR2_X1 U77bar ( .A1(abar[1]), .A2(bbar[14]), .ZN(ybar[30]) );
  AND2_X1 U78 ( .A1(b[2]), .A2(a[0]), .ZN(y[2]) );
  OR2_X1 U78bar ( .A1(bbar[2]), .A2(abar[0]), .ZN(ybar[2]) );
  AND2_X1 U79 ( .A1(a[1]), .A2(b[13]), .ZN(y[29]) );
  OR2_X1 U79bar ( .A1(abar[1]), .A2(bbar[13]), .ZN(ybar[29]) );
  AND2_X1 U80 ( .A1(a[1]), .A2(b[12]), .ZN(y[28]) );
  OR2_X1 U80bar ( .A1(abar[1]), .A2(bbar[12]), .ZN(ybar[28]) );
  AND2_X1 U81 ( .A1(a[1]), .A2(b[11]), .ZN(y[27]) );
  OR2_X1 U81bar ( .A1(abar[1]), .A2(bbar[11]), .ZN(ybar[27]) );
  AND2_X1 U82 ( .A1(a[1]), .A2(b[10]), .ZN(y[26]) );
  OR2_X1 U82bar ( .A1(abar[1]), .A2(bbar[10]), .ZN(ybar[26]) );
  AND2_X1 U83 ( .A1(a[1]), .A2(b[9]), .ZN(y[25]) );
  OR2_X1 U83bar ( .A1(abar[1]), .A2(bbar[9]), .ZN(ybar[25]) );
  AND2_X1 U84 ( .A1(a[15]), .A2(b[15]), .ZN(y[255]) );
  OR2_X1 U84bar ( .A1(abar[15]), .A2(bbar[15]), .ZN(ybar[255]) );
  AND2_X1 U85 ( .A1(a[15]), .A2(b[14]), .ZN(y[254]) );
  OR2_X1 U85bar ( .A1(abar[15]), .A2(bbar[14]), .ZN(ybar[254]) );
  AND2_X1 U86 ( .A1(a[15]), .A2(b[13]), .ZN(y[253]) );
  OR2_X1 U86bar ( .A1(abar[15]), .A2(bbar[13]), .ZN(ybar[253]) );
  AND2_X1 U87 ( .A1(a[15]), .A2(b[12]), .ZN(y[252]) );
  OR2_X1 U87bar ( .A1(abar[15]), .A2(bbar[12]), .ZN(ybar[252]) );
  AND2_X1 U88 ( .A1(a[15]), .A2(b[11]), .ZN(y[251]) );
  OR2_X1 U88bar ( .A1(abar[15]), .A2(bbar[11]), .ZN(ybar[251]) );
  AND2_X1 U89 ( .A1(a[15]), .A2(b[10]), .ZN(y[250]) );
  OR2_X1 U89bar ( .A1(abar[15]), .A2(bbar[10]), .ZN(ybar[250]) );
  AND2_X1 U90 ( .A1(a[1]), .A2(b[8]), .ZN(y[24]) );
  OR2_X1 U90bar ( .A1(abar[1]), .A2(bbar[8]), .ZN(ybar[24]) );
  AND2_X1 U91 ( .A1(a[15]), .A2(b[9]), .ZN(y[249]) );
  OR2_X1 U91bar ( .A1(abar[15]), .A2(bbar[9]), .ZN(ybar[249]) );
  AND2_X1 U92 ( .A1(a[15]), .A2(b[8]), .ZN(y[248]) );
  OR2_X1 U92bar ( .A1(abar[15]), .A2(bbar[8]), .ZN(ybar[248]) );
  AND2_X1 U93 ( .A1(a[15]), .A2(b[7]), .ZN(y[247]) );
  OR2_X1 U93bar ( .A1(abar[15]), .A2(bbar[7]), .ZN(ybar[247]) );
  AND2_X1 U94 ( .A1(a[15]), .A2(b[6]), .ZN(y[246]) );
  OR2_X1 U94bar ( .A1(abar[15]), .A2(bbar[6]), .ZN(ybar[246]) );
  AND2_X1 U95 ( .A1(a[15]), .A2(b[5]), .ZN(y[245]) );
  OR2_X1 U95bar ( .A1(abar[15]), .A2(bbar[5]), .ZN(ybar[245]) );
  AND2_X1 U96 ( .A1(a[15]), .A2(b[4]), .ZN(y[244]) );
  OR2_X1 U96bar ( .A1(abar[15]), .A2(bbar[4]), .ZN(ybar[244]) );
  AND2_X1 U97 ( .A1(a[15]), .A2(b[3]), .ZN(y[243]) );
  OR2_X1 U97bar ( .A1(abar[15]), .A2(bbar[3]), .ZN(ybar[243]) );
  AND2_X1 U98 ( .A1(a[15]), .A2(b[2]), .ZN(y[242]) );
  OR2_X1 U98bar ( .A1(abar[15]), .A2(bbar[2]), .ZN(ybar[242]) );
  AND2_X1 U99 ( .A1(a[15]), .A2(b[1]), .ZN(y[241]) );
  OR2_X1 U99bar ( .A1(abar[15]), .A2(bbar[1]), .ZN(ybar[241]) );
  AND2_X1 U100 ( .A1(a[15]), .A2(b[0]), .ZN(y[240]) );
  OR2_X1 U100bar ( .A1(abar[15]), .A2(bbar[0]), .ZN(ybar[240]) );
  AND2_X1 U101 ( .A1(a[1]), .A2(b[7]), .ZN(y[23]) );
  OR2_X1 U101bar ( .A1(abar[1]), .A2(bbar[7]), .ZN(ybar[23]) );
  AND2_X1 U102 ( .A1(a[14]), .A2(b[15]), .ZN(y[239]) );
  OR2_X1 U102bar ( .A1(abar[14]), .A2(bbar[15]), .ZN(ybar[239]) );
  AND2_X1 U103 ( .A1(a[14]), .A2(b[14]), .ZN(y[238]) );
  OR2_X1 U103bar ( .A1(abar[14]), .A2(bbar[14]), .ZN(ybar[238]) );
  AND2_X1 U104 ( .A1(a[14]), .A2(b[13]), .ZN(y[237]) );
  OR2_X1 U104bar ( .A1(abar[14]), .A2(bbar[13]), .ZN(ybar[237]) );
  AND2_X1 U105 ( .A1(a[14]), .A2(b[12]), .ZN(y[236]) );
  OR2_X1 U105bar ( .A1(abar[14]), .A2(bbar[12]), .ZN(ybar[236]) );
  AND2_X1 U106 ( .A1(a[14]), .A2(b[11]), .ZN(y[235]) );
  OR2_X1 U106bar ( .A1(abar[14]), .A2(bbar[11]), .ZN(ybar[235]) );
  AND2_X1 U107 ( .A1(a[14]), .A2(b[10]), .ZN(y[234]) );
  OR2_X1 U107bar ( .A1(abar[14]), .A2(bbar[10]), .ZN(ybar[234]) );
  AND2_X1 U108 ( .A1(a[14]), .A2(b[9]), .ZN(y[233]) );
  OR2_X1 U108bar ( .A1(abar[14]), .A2(bbar[9]), .ZN(ybar[233]) );
  AND2_X1 U109 ( .A1(a[14]), .A2(b[8]), .ZN(y[232]) );
  OR2_X1 U109bar ( .A1(abar[14]), .A2(bbar[8]), .ZN(ybar[232]) );
  AND2_X1 U110 ( .A1(a[14]), .A2(b[7]), .ZN(y[231]) );
  OR2_X1 U110bar ( .A1(abar[14]), .A2(bbar[7]), .ZN(ybar[231]) );
  AND2_X1 U111 ( .A1(a[14]), .A2(b[6]), .ZN(y[230]) );
  OR2_X1 U111bar ( .A1(abar[14]), .A2(bbar[6]), .ZN(ybar[230]) );
  AND2_X1 U112 ( .A1(a[1]), .A2(b[6]), .ZN(y[22]) );
  OR2_X1 U112bar ( .A1(abar[1]), .A2(bbar[6]), .ZN(ybar[22]) );
  AND2_X1 U113 ( .A1(a[14]), .A2(b[5]), .ZN(y[229]) );
  OR2_X1 U113bar ( .A1(abar[14]), .A2(bbar[5]), .ZN(ybar[229]) );
  AND2_X1 U114 ( .A1(a[14]), .A2(b[4]), .ZN(y[228]) );
  OR2_X1 U114bar ( .A1(abar[14]), .A2(bbar[4]), .ZN(ybar[228]) );
  AND2_X1 U115 ( .A1(a[14]), .A2(b[3]), .ZN(y[227]) );
  OR2_X1 U115bar ( .A1(abar[14]), .A2(bbar[3]), .ZN(ybar[227]) );
  AND2_X1 U116 ( .A1(a[14]), .A2(b[2]), .ZN(y[226]) );
  OR2_X1 U116bar ( .A1(abar[14]), .A2(bbar[2]), .ZN(ybar[226]) );
  AND2_X1 U117 ( .A1(a[14]), .A2(b[1]), .ZN(y[225]) );
  OR2_X1 U117bar ( .A1(abar[14]), .A2(bbar[1]), .ZN(ybar[225]) );
  AND2_X1 U118 ( .A1(a[14]), .A2(b[0]), .ZN(y[224]) );
  OR2_X1 U118bar ( .A1(abar[14]), .A2(bbar[0]), .ZN(ybar[224]) );
  AND2_X1 U119 ( .A1(a[13]), .A2(b[15]), .ZN(y[223]) );
  OR2_X1 U119bar ( .A1(abar[13]), .A2(bbar[15]), .ZN(ybar[223]) );
  AND2_X1 U120 ( .A1(a[13]), .A2(b[14]), .ZN(y[222]) );
  OR2_X1 U120bar ( .A1(abar[13]), .A2(bbar[14]), .ZN(ybar[222]) );
  AND2_X1 U121 ( .A1(a[13]), .A2(b[13]), .ZN(y[221]) );
  OR2_X1 U121bar ( .A1(abar[13]), .A2(bbar[13]), .ZN(ybar[221]) );
  AND2_X1 U122 ( .A1(a[13]), .A2(b[12]), .ZN(y[220]) );
  OR2_X1 U122bar ( .A1(abar[13]), .A2(bbar[12]), .ZN(ybar[220]) );
  AND2_X1 U123 ( .A1(a[1]), .A2(b[5]), .ZN(y[21]) );
  OR2_X1 U123bar ( .A1(abar[1]), .A2(bbar[5]), .ZN(ybar[21]) );
  AND2_X1 U124 ( .A1(a[13]), .A2(b[11]), .ZN(y[219]) );
  OR2_X1 U124bar ( .A1(abar[13]), .A2(bbar[11]), .ZN(ybar[219]) );
  AND2_X1 U125 ( .A1(a[13]), .A2(b[10]), .ZN(y[218]) );
  OR2_X1 U125bar ( .A1(abar[13]), .A2(bbar[10]), .ZN(ybar[218]) );
  AND2_X1 U126 ( .A1(a[13]), .A2(b[9]), .ZN(y[217]) );
  OR2_X1 U126bar ( .A1(abar[13]), .A2(bbar[9]), .ZN(ybar[217]) );
  AND2_X1 U127 ( .A1(a[13]), .A2(b[8]), .ZN(y[216]) );
  OR2_X1 U127bar ( .A1(abar[13]), .A2(bbar[8]), .ZN(ybar[216]) );
  AND2_X1 U128 ( .A1(a[13]), .A2(b[7]), .ZN(y[215]) );
  OR2_X1 U128bar ( .A1(abar[13]), .A2(bbar[7]), .ZN(ybar[215]) );
  AND2_X1 U129 ( .A1(a[13]), .A2(b[6]), .ZN(y[214]) );
  OR2_X1 U129bar ( .A1(abar[13]), .A2(bbar[6]), .ZN(ybar[214]) );
  AND2_X1 U130 ( .A1(a[13]), .A2(b[5]), .ZN(y[213]) );
  OR2_X1 U130bar ( .A1(abar[13]), .A2(bbar[5]), .ZN(ybar[213]) );
  AND2_X1 U131 ( .A1(a[13]), .A2(b[4]), .ZN(y[212]) );
  OR2_X1 U131bar ( .A1(abar[13]), .A2(bbar[4]), .ZN(ybar[212]) );
  AND2_X1 U132 ( .A1(a[13]), .A2(b[3]), .ZN(y[211]) );
  OR2_X1 U132bar ( .A1(abar[13]), .A2(bbar[3]), .ZN(ybar[211]) );
  AND2_X1 U133 ( .A1(a[13]), .A2(b[2]), .ZN(y[210]) );
  OR2_X1 U133bar ( .A1(abar[13]), .A2(bbar[2]), .ZN(ybar[210]) );
  AND2_X1 U134 ( .A1(a[1]), .A2(b[4]), .ZN(y[20]) );
  OR2_X1 U134bar ( .A1(abar[1]), .A2(bbar[4]), .ZN(ybar[20]) );
  AND2_X1 U135 ( .A1(a[13]), .A2(b[1]), .ZN(y[209]) );
  OR2_X1 U135bar ( .A1(abar[13]), .A2(bbar[1]), .ZN(ybar[209]) );
  AND2_X1 U136 ( .A1(a[13]), .A2(b[0]), .ZN(y[208]) );
  OR2_X1 U136bar ( .A1(abar[13]), .A2(bbar[0]), .ZN(ybar[208]) );
  AND2_X1 U137 ( .A1(a[12]), .A2(b[15]), .ZN(y[207]) );
  OR2_X1 U137bar ( .A1(abar[12]), .A2(bbar[15]), .ZN(ybar[207]) );
  AND2_X1 U138 ( .A1(a[12]), .A2(b[14]), .ZN(y[206]) );
  OR2_X1 U138bar ( .A1(abar[12]), .A2(bbar[14]), .ZN(ybar[206]) );
  AND2_X1 U139 ( .A1(a[12]), .A2(b[13]), .ZN(y[205]) );
  OR2_X1 U139bar ( .A1(abar[12]), .A2(bbar[13]), .ZN(ybar[205]) );
  AND2_X1 U140 ( .A1(a[12]), .A2(b[12]), .ZN(y[204]) );
  OR2_X1 U140bar ( .A1(abar[12]), .A2(bbar[12]), .ZN(ybar[204]) );
  AND2_X1 U141 ( .A1(a[12]), .A2(b[11]), .ZN(y[203]) );
  OR2_X1 U141bar ( .A1(abar[12]), .A2(bbar[11]), .ZN(ybar[203]) );
  AND2_X1 U142 ( .A1(a[12]), .A2(b[10]), .ZN(y[202]) );
  OR2_X1 U142bar ( .A1(abar[12]), .A2(bbar[10]), .ZN(ybar[202]) );
  AND2_X1 U143 ( .A1(a[12]), .A2(b[9]), .ZN(y[201]) );
  OR2_X1 U143bar ( .A1(abar[12]), .A2(bbar[9]), .ZN(ybar[201]) );
  AND2_X1 U144 ( .A1(a[12]), .A2(b[8]), .ZN(y[200]) );
  OR2_X1 U144bar ( .A1(abar[12]), .A2(bbar[8]), .ZN(ybar[200]) );
  AND2_X1 U145 ( .A1(b[1]), .A2(a[0]), .ZN(y[1]) );
  OR2_X1 U145bar ( .A1(bbar[1]), .A2(abar[0]), .ZN(ybar[1]) );
  AND2_X1 U146 ( .A1(a[1]), .A2(b[3]), .ZN(y[19]) );
  OR2_X1 U146bar ( .A1(abar[1]), .A2(bbar[3]), .ZN(ybar[19]) );
  AND2_X1 U147 ( .A1(a[12]), .A2(b[7]), .ZN(y[199]) );
  OR2_X1 U147bar ( .A1(abar[12]), .A2(bbar[7]), .ZN(ybar[199]) );
  AND2_X1 U148 ( .A1(a[12]), .A2(b[6]), .ZN(y[198]) );
  OR2_X1 U148bar ( .A1(abar[12]), .A2(bbar[6]), .ZN(ybar[198]) );
  AND2_X1 U149 ( .A1(a[12]), .A2(b[5]), .ZN(y[197]) );
  OR2_X1 U149bar ( .A1(abar[12]), .A2(bbar[5]), .ZN(ybar[197]) );
  AND2_X1 U150 ( .A1(a[12]), .A2(b[4]), .ZN(y[196]) );
  OR2_X1 U150bar ( .A1(abar[12]), .A2(bbar[4]), .ZN(ybar[196]) );
  AND2_X1 U151 ( .A1(a[12]), .A2(b[3]), .ZN(y[195]) );
  OR2_X1 U151bar ( .A1(abar[12]), .A2(bbar[3]), .ZN(ybar[195]) );
  AND2_X1 U152 ( .A1(a[12]), .A2(b[2]), .ZN(y[194]) );
  OR2_X1 U152bar ( .A1(abar[12]), .A2(bbar[2]), .ZN(ybar[194]) );
  AND2_X1 U153 ( .A1(a[12]), .A2(b[1]), .ZN(y[193]) );
  OR2_X1 U153bar ( .A1(abar[12]), .A2(bbar[1]), .ZN(ybar[193]) );
  AND2_X1 U154 ( .A1(a[12]), .A2(b[0]), .ZN(y[192]) );
  OR2_X1 U154bar ( .A1(abar[12]), .A2(bbar[0]), .ZN(ybar[192]) );
  AND2_X1 U155 ( .A1(a[11]), .A2(b[15]), .ZN(y[191]) );
  OR2_X1 U155bar ( .A1(abar[11]), .A2(bbar[15]), .ZN(ybar[191]) );
  AND2_X1 U156 ( .A1(a[11]), .A2(b[14]), .ZN(y[190]) );
  OR2_X1 U156bar ( .A1(abar[11]), .A2(bbar[14]), .ZN(ybar[190]) );
  AND2_X1 U157 ( .A1(a[1]), .A2(b[2]), .ZN(y[18]) );
  OR2_X1 U157bar ( .A1(abar[1]), .A2(bbar[2]), .ZN(ybar[18]) );
  AND2_X1 U158 ( .A1(a[11]), .A2(b[13]), .ZN(y[189]) );
  OR2_X1 U158bar ( .A1(abar[11]), .A2(bbar[13]), .ZN(ybar[189]) );
  AND2_X1 U159 ( .A1(a[11]), .A2(b[12]), .ZN(y[188]) );
  OR2_X1 U159bar ( .A1(abar[11]), .A2(bbar[12]), .ZN(ybar[188]) );
  AND2_X1 U160 ( .A1(a[11]), .A2(b[11]), .ZN(y[187]) );
  OR2_X1 U160bar ( .A1(abar[11]), .A2(bbar[11]), .ZN(ybar[187]) );
  AND2_X1 U161 ( .A1(a[11]), .A2(b[10]), .ZN(y[186]) );
  OR2_X1 U161bar ( .A1(abar[11]), .A2(bbar[10]), .ZN(ybar[186]) );
  AND2_X1 U162 ( .A1(a[11]), .A2(b[9]), .ZN(y[185]) );
  OR2_X1 U162bar ( .A1(abar[11]), .A2(bbar[9]), .ZN(ybar[185]) );
  AND2_X1 U163 ( .A1(a[11]), .A2(b[8]), .ZN(y[184]) );
  OR2_X1 U163bar ( .A1(abar[11]), .A2(bbar[8]), .ZN(ybar[184]) );
  AND2_X1 U164 ( .A1(a[11]), .A2(b[7]), .ZN(y[183]) );
  OR2_X1 U164bar ( .A1(abar[11]), .A2(bbar[7]), .ZN(ybar[183]) );
  AND2_X1 U165 ( .A1(a[11]), .A2(b[6]), .ZN(y[182]) );
  OR2_X1 U165bar ( .A1(abar[11]), .A2(bbar[6]), .ZN(ybar[182]) );
  AND2_X1 U166 ( .A1(a[11]), .A2(b[5]), .ZN(y[181]) );
  OR2_X1 U166bar ( .A1(abar[11]), .A2(bbar[5]), .ZN(ybar[181]) );
  AND2_X1 U167 ( .A1(a[11]), .A2(b[4]), .ZN(y[180]) );
  OR2_X1 U167bar ( .A1(abar[11]), .A2(bbar[4]), .ZN(ybar[180]) );
  AND2_X1 U168 ( .A1(a[1]), .A2(b[1]), .ZN(y[17]) );
  OR2_X1 U168bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[17]) );
  AND2_X1 U169 ( .A1(a[11]), .A2(b[3]), .ZN(y[179]) );
  OR2_X1 U169bar ( .A1(abar[11]), .A2(bbar[3]), .ZN(ybar[179]) );
  AND2_X1 U170 ( .A1(a[11]), .A2(b[2]), .ZN(y[178]) );
  OR2_X1 U170bar ( .A1(abar[11]), .A2(bbar[2]), .ZN(ybar[178]) );
  AND2_X1 U171 ( .A1(a[11]), .A2(b[1]), .ZN(y[177]) );
  OR2_X1 U171bar ( .A1(abar[11]), .A2(bbar[1]), .ZN(ybar[177]) );
  AND2_X1 U172 ( .A1(a[11]), .A2(b[0]), .ZN(y[176]) );
  OR2_X1 U172bar ( .A1(abar[11]), .A2(bbar[0]), .ZN(ybar[176]) );
  AND2_X1 U173 ( .A1(a[10]), .A2(b[15]), .ZN(y[175]) );
  OR2_X1 U173bar ( .A1(abar[10]), .A2(bbar[15]), .ZN(ybar[175]) );
  AND2_X1 U174 ( .A1(a[10]), .A2(b[14]), .ZN(y[174]) );
  OR2_X1 U174bar ( .A1(abar[10]), .A2(bbar[14]), .ZN(ybar[174]) );
  AND2_X1 U175 ( .A1(a[10]), .A2(b[13]), .ZN(y[173]) );
  OR2_X1 U175bar ( .A1(abar[10]), .A2(bbar[13]), .ZN(ybar[173]) );
  AND2_X1 U176 ( .A1(a[10]), .A2(b[12]), .ZN(y[172]) );
  OR2_X1 U176bar ( .A1(abar[10]), .A2(bbar[12]), .ZN(ybar[172]) );
  AND2_X1 U177 ( .A1(a[10]), .A2(b[11]), .ZN(y[171]) );
  OR2_X1 U177bar ( .A1(abar[10]), .A2(bbar[11]), .ZN(ybar[171]) );
  AND2_X1 U178 ( .A1(a[10]), .A2(b[10]), .ZN(y[170]) );
  OR2_X1 U178bar ( .A1(abar[10]), .A2(bbar[10]), .ZN(ybar[170]) );
  AND2_X1 U179 ( .A1(a[1]), .A2(b[0]), .ZN(y[16]) );
  OR2_X1 U179bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[16]) );
  AND2_X1 U180 ( .A1(a[10]), .A2(b[9]), .ZN(y[169]) );
  OR2_X1 U180bar ( .A1(abar[10]), .A2(bbar[9]), .ZN(ybar[169]) );
  AND2_X1 U181 ( .A1(a[10]), .A2(b[8]), .ZN(y[168]) );
  OR2_X1 U181bar ( .A1(abar[10]), .A2(bbar[8]), .ZN(ybar[168]) );
  AND2_X1 U182 ( .A1(a[10]), .A2(b[7]), .ZN(y[167]) );
  OR2_X1 U182bar ( .A1(abar[10]), .A2(bbar[7]), .ZN(ybar[167]) );
  AND2_X1 U183 ( .A1(a[10]), .A2(b[6]), .ZN(y[166]) );
  OR2_X1 U183bar ( .A1(abar[10]), .A2(bbar[6]), .ZN(ybar[166]) );
  AND2_X1 U184 ( .A1(a[10]), .A2(b[5]), .ZN(y[165]) );
  OR2_X1 U184bar ( .A1(abar[10]), .A2(bbar[5]), .ZN(ybar[165]) );
  AND2_X1 U185 ( .A1(a[10]), .A2(b[4]), .ZN(y[164]) );
  OR2_X1 U185bar ( .A1(abar[10]), .A2(bbar[4]), .ZN(ybar[164]) );
  AND2_X1 U186 ( .A1(a[10]), .A2(b[3]), .ZN(y[163]) );
  OR2_X1 U186bar ( .A1(abar[10]), .A2(bbar[3]), .ZN(ybar[163]) );
  AND2_X1 U187 ( .A1(a[10]), .A2(b[2]), .ZN(y[162]) );
  OR2_X1 U187bar ( .A1(abar[10]), .A2(bbar[2]), .ZN(ybar[162]) );
  AND2_X1 U188 ( .A1(a[10]), .A2(b[1]), .ZN(y[161]) );
  OR2_X1 U188bar ( .A1(abar[10]), .A2(bbar[1]), .ZN(ybar[161]) );
  AND2_X1 U189 ( .A1(a[10]), .A2(b[0]), .ZN(y[160]) );
  OR2_X1 U189bar ( .A1(abar[10]), .A2(bbar[0]), .ZN(ybar[160]) );
  AND2_X1 U190 ( .A1(b[15]), .A2(a[0]), .ZN(y[15]) );
  OR2_X1 U190bar ( .A1(bbar[15]), .A2(abar[0]), .ZN(ybar[15]) );
  AND2_X1 U191 ( .A1(a[9]), .A2(b[15]), .ZN(y[159]) );
  OR2_X1 U191bar ( .A1(abar[9]), .A2(bbar[15]), .ZN(ybar[159]) );
  AND2_X1 U192 ( .A1(a[9]), .A2(b[14]), .ZN(y[158]) );
  OR2_X1 U192bar ( .A1(abar[9]), .A2(bbar[14]), .ZN(ybar[158]) );
  AND2_X1 U193 ( .A1(a[9]), .A2(b[13]), .ZN(y[157]) );
  OR2_X1 U193bar ( .A1(abar[9]), .A2(bbar[13]), .ZN(ybar[157]) );
  AND2_X1 U194 ( .A1(a[9]), .A2(b[12]), .ZN(y[156]) );
  OR2_X1 U194bar ( .A1(abar[9]), .A2(bbar[12]), .ZN(ybar[156]) );
  AND2_X1 U195 ( .A1(a[9]), .A2(b[11]), .ZN(y[155]) );
  OR2_X1 U195bar ( .A1(abar[9]), .A2(bbar[11]), .ZN(ybar[155]) );
  AND2_X1 U196 ( .A1(a[9]), .A2(b[10]), .ZN(y[154]) );
  OR2_X1 U196bar ( .A1(abar[9]), .A2(bbar[10]), .ZN(ybar[154]) );
  AND2_X1 U197 ( .A1(a[9]), .A2(b[9]), .ZN(y[153]) );
  OR2_X1 U197bar ( .A1(abar[9]), .A2(bbar[9]), .ZN(ybar[153]) );
  AND2_X1 U198 ( .A1(a[9]), .A2(b[8]), .ZN(y[152]) );
  OR2_X1 U198bar ( .A1(abar[9]), .A2(bbar[8]), .ZN(ybar[152]) );
  AND2_X1 U199 ( .A1(a[9]), .A2(b[7]), .ZN(y[151]) );
  OR2_X1 U199bar ( .A1(abar[9]), .A2(bbar[7]), .ZN(ybar[151]) );
  AND2_X1 U200 ( .A1(a[9]), .A2(b[6]), .ZN(y[150]) );
  OR2_X1 U200bar ( .A1(abar[9]), .A2(bbar[6]), .ZN(ybar[150]) );
  AND2_X1 U201 ( .A1(b[14]), .A2(a[0]), .ZN(y[14]) );
  OR2_X1 U201bar ( .A1(bbar[14]), .A2(abar[0]), .ZN(ybar[14]) );
  AND2_X1 U202 ( .A1(a[9]), .A2(b[5]), .ZN(y[149]) );
  OR2_X1 U202bar ( .A1(abar[9]), .A2(bbar[5]), .ZN(ybar[149]) );
  AND2_X1 U203 ( .A1(a[9]), .A2(b[4]), .ZN(y[148]) );
  OR2_X1 U203bar ( .A1(abar[9]), .A2(bbar[4]), .ZN(ybar[148]) );
  AND2_X1 U204 ( .A1(a[9]), .A2(b[3]), .ZN(y[147]) );
  OR2_X1 U204bar ( .A1(abar[9]), .A2(bbar[3]), .ZN(ybar[147]) );
  AND2_X1 U205 ( .A1(a[9]), .A2(b[2]), .ZN(y[146]) );
  OR2_X1 U205bar ( .A1(abar[9]), .A2(bbar[2]), .ZN(ybar[146]) );
  AND2_X1 U206 ( .A1(a[9]), .A2(b[1]), .ZN(y[145]) );
  OR2_X1 U206bar ( .A1(abar[9]), .A2(bbar[1]), .ZN(ybar[145]) );
  AND2_X1 U207 ( .A1(a[9]), .A2(b[0]), .ZN(y[144]) );
  OR2_X1 U207bar ( .A1(abar[9]), .A2(bbar[0]), .ZN(ybar[144]) );
  AND2_X1 U208 ( .A1(a[8]), .A2(b[15]), .ZN(y[143]) );
  OR2_X1 U208bar ( .A1(abar[8]), .A2(bbar[15]), .ZN(ybar[143]) );
  AND2_X1 U209 ( .A1(a[8]), .A2(b[14]), .ZN(y[142]) );
  OR2_X1 U209bar ( .A1(abar[8]), .A2(bbar[14]), .ZN(ybar[142]) );
  AND2_X1 U210 ( .A1(a[8]), .A2(b[13]), .ZN(y[141]) );
  OR2_X1 U210bar ( .A1(abar[8]), .A2(bbar[13]), .ZN(ybar[141]) );
  AND2_X1 U211 ( .A1(a[8]), .A2(b[12]), .ZN(y[140]) );
  OR2_X1 U211bar ( .A1(abar[8]), .A2(bbar[12]), .ZN(ybar[140]) );
  AND2_X1 U212 ( .A1(b[13]), .A2(a[0]), .ZN(y[13]) );
  OR2_X1 U212bar ( .A1(bbar[13]), .A2(abar[0]), .ZN(ybar[13]) );
  AND2_X1 U213 ( .A1(a[8]), .A2(b[11]), .ZN(y[139]) );
  OR2_X1 U213bar ( .A1(abar[8]), .A2(bbar[11]), .ZN(ybar[139]) );
  AND2_X1 U214 ( .A1(a[8]), .A2(b[10]), .ZN(y[138]) );
  OR2_X1 U214bar ( .A1(abar[8]), .A2(bbar[10]), .ZN(ybar[138]) );
  AND2_X1 U215 ( .A1(a[8]), .A2(b[9]), .ZN(y[137]) );
  OR2_X1 U215bar ( .A1(abar[8]), .A2(bbar[9]), .ZN(ybar[137]) );
  AND2_X1 U216 ( .A1(a[8]), .A2(b[8]), .ZN(y[136]) );
  OR2_X1 U216bar ( .A1(abar[8]), .A2(bbar[8]), .ZN(ybar[136]) );
  AND2_X1 U217 ( .A1(a[8]), .A2(b[7]), .ZN(y[135]) );
  OR2_X1 U217bar ( .A1(abar[8]), .A2(bbar[7]), .ZN(ybar[135]) );
  AND2_X1 U218 ( .A1(a[8]), .A2(b[6]), .ZN(y[134]) );
  OR2_X1 U218bar ( .A1(abar[8]), .A2(bbar[6]), .ZN(ybar[134]) );
  AND2_X1 U219 ( .A1(a[8]), .A2(b[5]), .ZN(y[133]) );
  OR2_X1 U219bar ( .A1(abar[8]), .A2(bbar[5]), .ZN(ybar[133]) );
  AND2_X1 U220 ( .A1(a[8]), .A2(b[4]), .ZN(y[132]) );
  OR2_X1 U220bar ( .A1(abar[8]), .A2(bbar[4]), .ZN(ybar[132]) );
  AND2_X1 U221 ( .A1(a[8]), .A2(b[3]), .ZN(y[131]) );
  OR2_X1 U221bar ( .A1(abar[8]), .A2(bbar[3]), .ZN(ybar[131]) );
  AND2_X1 U222 ( .A1(a[8]), .A2(b[2]), .ZN(y[130]) );
  OR2_X1 U222bar ( .A1(abar[8]), .A2(bbar[2]), .ZN(ybar[130]) );
  AND2_X1 U223 ( .A1(b[12]), .A2(a[0]), .ZN(y[12]) );
  OR2_X1 U223bar ( .A1(bbar[12]), .A2(abar[0]), .ZN(ybar[12]) );
  AND2_X1 U224 ( .A1(a[8]), .A2(b[1]), .ZN(y[129]) );
  OR2_X1 U224bar ( .A1(abar[8]), .A2(bbar[1]), .ZN(ybar[129]) );
  AND2_X1 U225 ( .A1(a[8]), .A2(b[0]), .ZN(y[128]) );
  OR2_X1 U225bar ( .A1(abar[8]), .A2(bbar[0]), .ZN(ybar[128]) );
  AND2_X1 U226 ( .A1(a[7]), .A2(b[15]), .ZN(y[127]) );
  OR2_X1 U226bar ( .A1(abar[7]), .A2(bbar[15]), .ZN(ybar[127]) );
  AND2_X1 U227 ( .A1(a[7]), .A2(b[14]), .ZN(y[126]) );
  OR2_X1 U227bar ( .A1(abar[7]), .A2(bbar[14]), .ZN(ybar[126]) );
  AND2_X1 U228 ( .A1(a[7]), .A2(b[13]), .ZN(y[125]) );
  OR2_X1 U228bar ( .A1(abar[7]), .A2(bbar[13]), .ZN(ybar[125]) );
  AND2_X1 U229 ( .A1(a[7]), .A2(b[12]), .ZN(y[124]) );
  OR2_X1 U229bar ( .A1(abar[7]), .A2(bbar[12]), .ZN(ybar[124]) );
  AND2_X1 U230 ( .A1(a[7]), .A2(b[11]), .ZN(y[123]) );
  OR2_X1 U230bar ( .A1(abar[7]), .A2(bbar[11]), .ZN(ybar[123]) );
  AND2_X1 U231 ( .A1(a[7]), .A2(b[10]), .ZN(y[122]) );
  OR2_X1 U231bar ( .A1(abar[7]), .A2(bbar[10]), .ZN(ybar[122]) );
  AND2_X1 U232 ( .A1(a[7]), .A2(b[9]), .ZN(y[121]) );
  OR2_X1 U232bar ( .A1(abar[7]), .A2(bbar[9]), .ZN(ybar[121]) );
  AND2_X1 U233 ( .A1(a[7]), .A2(b[8]), .ZN(y[120]) );
  OR2_X1 U233bar ( .A1(abar[7]), .A2(bbar[8]), .ZN(ybar[120]) );
  AND2_X1 U234 ( .A1(b[11]), .A2(a[0]), .ZN(y[11]) );
  OR2_X1 U234bar ( .A1(bbar[11]), .A2(abar[0]), .ZN(ybar[11]) );
  AND2_X1 U235 ( .A1(a[7]), .A2(b[7]), .ZN(y[119]) );
  OR2_X1 U235bar ( .A1(abar[7]), .A2(bbar[7]), .ZN(ybar[119]) );
  AND2_X1 U236 ( .A1(a[7]), .A2(b[6]), .ZN(y[118]) );
  OR2_X1 U236bar ( .A1(abar[7]), .A2(bbar[6]), .ZN(ybar[118]) );
  AND2_X1 U237 ( .A1(a[7]), .A2(b[5]), .ZN(y[117]) );
  OR2_X1 U237bar ( .A1(abar[7]), .A2(bbar[5]), .ZN(ybar[117]) );
  AND2_X1 U238 ( .A1(a[7]), .A2(b[4]), .ZN(y[116]) );
  OR2_X1 U238bar ( .A1(abar[7]), .A2(bbar[4]), .ZN(ybar[116]) );
  AND2_X1 U239 ( .A1(a[7]), .A2(b[3]), .ZN(y[115]) );
  OR2_X1 U239bar ( .A1(abar[7]), .A2(bbar[3]), .ZN(ybar[115]) );
  AND2_X1 U240 ( .A1(a[7]), .A2(b[2]), .ZN(y[114]) );
  OR2_X1 U240bar ( .A1(abar[7]), .A2(bbar[2]), .ZN(ybar[114]) );
  AND2_X1 U241 ( .A1(a[7]), .A2(b[1]), .ZN(y[113]) );
  OR2_X1 U241bar ( .A1(abar[7]), .A2(bbar[1]), .ZN(ybar[113]) );
  AND2_X1 U242 ( .A1(a[7]), .A2(b[0]), .ZN(y[112]) );
  OR2_X1 U242bar ( .A1(abar[7]), .A2(bbar[0]), .ZN(ybar[112]) );
  AND2_X1 U243 ( .A1(b[15]), .A2(a[6]), .ZN(y[111]) );
  OR2_X1 U243bar ( .A1(bbar[15]), .A2(abar[6]), .ZN(ybar[111]) );
  AND2_X1 U244 ( .A1(b[14]), .A2(a[6]), .ZN(y[110]) );
  OR2_X1 U244bar ( .A1(bbar[14]), .A2(abar[6]), .ZN(ybar[110]) );
  AND2_X1 U245 ( .A1(b[10]), .A2(a[0]), .ZN(y[10]) );
  OR2_X1 U245bar ( .A1(bbar[10]), .A2(abar[0]), .ZN(ybar[10]) );
  AND2_X1 U246 ( .A1(b[13]), .A2(a[6]), .ZN(y[109]) );
  OR2_X1 U246bar ( .A1(bbar[13]), .A2(abar[6]), .ZN(ybar[109]) );
  AND2_X1 U247 ( .A1(b[12]), .A2(a[6]), .ZN(y[108]) );
  OR2_X1 U247bar ( .A1(bbar[12]), .A2(abar[6]), .ZN(ybar[108]) );
  AND2_X1 U248 ( .A1(b[11]), .A2(a[6]), .ZN(y[107]) );
  OR2_X1 U248bar ( .A1(bbar[11]), .A2(abar[6]), .ZN(ybar[107]) );
  AND2_X1 U249 ( .A1(b[10]), .A2(a[6]), .ZN(y[106]) );
  OR2_X1 U249bar ( .A1(bbar[10]), .A2(abar[6]), .ZN(ybar[106]) );
  AND2_X1 U250 ( .A1(a[6]), .A2(b[9]), .ZN(y[105]) );
  OR2_X1 U250bar ( .A1(abar[6]), .A2(bbar[9]), .ZN(ybar[105]) );
  AND2_X1 U251 ( .A1(b[8]), .A2(a[6]), .ZN(y[104]) );
  OR2_X1 U251bar ( .A1(bbar[8]), .A2(abar[6]), .ZN(ybar[104]) );
  AND2_X1 U252 ( .A1(b[7]), .A2(a[6]), .ZN(y[103]) );
  OR2_X1 U252bar ( .A1(bbar[7]), .A2(abar[6]), .ZN(ybar[103]) );
  AND2_X1 U253 ( .A1(b[6]), .A2(a[6]), .ZN(y[102]) );
  OR2_X1 U253bar ( .A1(bbar[6]), .A2(abar[6]), .ZN(ybar[102]) );
  AND2_X1 U254 ( .A1(b[5]), .A2(a[6]), .ZN(y[101]) );
  OR2_X1 U254bar ( .A1(bbar[5]), .A2(abar[6]), .ZN(ybar[101]) );
  AND2_X1 U255 ( .A1(b[4]), .A2(a[6]), .ZN(y[100]) );
  OR2_X1 U255bar ( .A1(bbar[4]), .A2(abar[6]), .ZN(ybar[100]) );
  AND2_X1 U256 ( .A1(b[0]), .A2(a[0]), .ZN(y[0]) );
  OR2_X1 U256bar ( .A1(bbar[0]), .A2(abar[0]), .ZN(ybar[0]) );
endmodule

module decode_14 ( in, inbar, out, outbar );

  input wire [7:0] in;
  input wire [7:0] inbar;
//input_done

  output wire [255:0] out;
  output wire [255:0] outbar;
//output_done

  wire [15:0] level1;
  wire [31:0] level2;
  wire [15:0] level1bar;
  wire [31:0] level2bar;
//wire_done

  CD2_56 cd_l1_1 ( .a(in[1]), .abar(inbar[1]), .b(in[0]), .bbar(inbar[0]), .y(level1[3:0]), .ybar(level1bar[3:0]) );
  CD2_55 cd_l1_2 ( .a(in[3]), .abar(inbar[3]), .b(in[2]), .bbar(inbar[2]), .y(level1[7:4]), .ybar(level1bar[7:4]) );
  CD2_54 cd_l1_3 ( .a(in[5]), .abar(inbar[5]), .b(in[4]), .bbar(inbar[4]), .y(level1[11:8]), .ybar(level1bar[11:8]) );
  CD2_53 cd_l1_4 ( .a(in[7]), .abar(inbar[7]), .b(in[6]), .bbar(inbar[6]), .y(level1[15:12]), .ybar(level1bar[15:12]) );

  CD4_28 cd_l2_1 ( .a(level1[7:4]), .abar(level1bar[7:4]), .b(level1[3:0]), .bbar(level1bar[3:0]), 
        .y(level2[15:0]), .ybar(level2bar[15:0]) );
  CD4_27 cd_l2_2 ( .a(level1[15:12]), .abar(level1bar[15:12]), .b(level1[11:8]), .bbar(level1bar[11:8]), 
        .y(level2[31:16]), .ybar(level2bar[31:16]) );
  CD16_14 cd_l3 ( .a(level2[31:16]), .abar(level2bar[31:16]), .b(level2[15:0]), .bbar(level2bar[15:0]), 
        .y(out), .ybar(outbar) );
endmodule

module encode_14 ( in, inbar, out, outbar );

  input wire [255:0] in;
  input wire [255:0] inbar;
//input_done

  output wire [7:0] out;
  output wire [7:0] outbar;
//output_done

  wire in_81;
  wire in_80;
  wire in_79;
  wire in_78;
  wire in_77;
  wire in_76;
  wire in_75;
  wire in_74;
  wire in_73;
  wire in_72;
  wire in_71;
  wire in_70;
  wire in_69;
  wire in_68;
  wire in_67;
  wire in_66;
  wire in_65;
  wire in_64;
  wire in_63;
  wire in_62;
  wire in_61;
  wire in_60;
  wire in_59;
  wire in_58;
  wire in_57;
  wire in_56;
  wire in_55;
  wire in_54;
  wire in_53;
  wire in_52;
  wire in_51;
  wire in_50;
  wire in_49;
  wire in_48;
  wire in_47;
  wire in_46;
  wire in_45;
  wire in_44;
  wire in_43;
  wire in_42;
  wire in_41;
  wire in_40;
  wire in_39;
  wire in_38;
  wire in_37;
  wire in_36;
  wire in_35;
  wire in_34;
  wire in_33;
  wire in_32;
  wire in_31;
  wire in_30;
  wire in_29;
  wire in_28;
  wire in_27;
  wire in_26;
  wire in_25;
  wire in_24;
  wire in_23;
  wire in_22;
  wire in_21;
  wire in_20;
  wire in_19;
  wire in_18;
  wire in_17;
  wire in_16;
  wire in_15;
  wire in_14;
  wire in_13;
  wire in_12;
  wire in_11;
  wire in_10;
  wire in_9;
  wire in_8;
  wire in_7;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_3;
  wire in_2;
  wire in_1;
  wire in_0;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire in_81bar;
  wire in_80bar;
  wire in_79bar;
  wire in_78bar;
  wire in_77bar;
  wire in_76bar;
  wire in_75bar;
  wire in_74bar;
  wire in_73bar;
  wire in_72bar;
  wire in_71bar;
  wire in_70bar;
  wire in_69bar;
  wire in_68bar;
  wire in_67bar;
  wire in_66bar;
  wire in_65bar;
  wire in_64bar;
  wire in_63bar;
  wire in_62bar;
  wire in_61bar;
  wire in_60bar;
  wire in_59bar;
  wire in_58bar;
  wire in_57bar;
  wire in_56bar;
  wire in_55bar;
  wire in_54bar;
  wire in_53bar;
  wire in_52bar;
  wire in_51bar;
  wire in_50bar;
  wire in_49bar;
  wire in_48bar;
  wire in_47bar;
  wire in_46bar;
  wire in_45bar;
  wire in_44bar;
  wire in_43bar;
  wire in_42bar;
  wire in_41bar;
  wire in_40bar;
  wire in_39bar;
  wire in_38bar;
  wire in_37bar;
  wire in_36bar;
  wire in_35bar;
  wire in_34bar;
  wire in_33bar;
  wire in_32bar;
  wire in_31bar;
  wire in_30bar;
  wire in_29bar;
  wire in_28bar;
  wire in_27bar;
  wire in_26bar;
  wire in_25bar;
  wire in_24bar;
  wire in_23bar;
  wire in_22bar;
  wire in_21bar;
  wire in_20bar;
  wire in_19bar;
  wire in_18bar;
  wire in_17bar;
  wire in_16bar;
  wire in_15bar;
  wire in_14bar;
  wire in_13bar;
  wire in_12bar;
  wire in_11bar;
  wire in_10bar;
  wire in_9bar;
  wire in_8bar;
  wire in_7bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_3bar;
  wire in_2bar;
  wire in_1bar;
  wire in_0bar;
  wire n487bar;
  wire n488bar;
  wire n489bar;
  wire n490bar;
  wire n491bar;
  wire n492bar;
  wire n493bar;
  wire n494bar;
  wire n495bar;
  wire n496bar;
  wire n497bar;
  wire n498bar;
  wire n499bar;
  wire n500bar;
  wire n501bar;
  wire n502bar;
  wire n503bar;
  wire n504bar;
  wire n505bar;
  wire n506bar;
  wire n507bar;
  wire n508bar;
  wire n509bar;
  wire n510bar;
  wire n511bar;
  wire n512bar;
  wire n513bar;
  wire n514bar;
  wire n515bar;
  wire n516bar;
  wire n517bar;
  wire n518bar;
  wire n519bar;
  wire n520bar;
  wire n521bar;
  wire n522bar;
  wire n523bar;
  wire n524bar;
  wire n525bar;
  wire n526bar;
  wire n527bar;
  wire n528bar;
  wire n529bar;
  wire n530bar;
  wire n531bar;
  wire n532bar;
  wire n533bar;
  wire n534bar;
  wire n535bar;
  wire n536bar;
  wire n537bar;
  wire n538bar;
  wire n539bar;
  wire n540bar;
  wire n541bar;
  wire n542bar;
  wire n543bar;
  wire n544bar;
  wire n545bar;
  wire n546bar;
  wire n547bar;
  wire n548bar;
  wire n549bar;
  wire n550bar;
  wire n551bar;
  wire n552bar;
  wire n553bar;
  wire n554bar;
  wire n555bar;
  wire n556bar;
  wire n557bar;
  wire n558bar;
  wire n559bar;
  wire n560bar;
  wire n561bar;
  wire n562bar;
  wire n563bar;
  wire n564bar;
  wire n565bar;
  wire n566bar;
  wire n567bar;
  wire n568bar;
  wire n569bar;
  wire n570bar;
  wire n571bar;
  wire n572bar;
  wire n573bar;
  wire n574bar;
  wire n575bar;
  wire n576bar;
  wire n577bar;
  wire n578bar;
  wire n579bar;
  wire n580bar;
  wire n581bar;
  wire n582bar;
  wire n583bar;
  wire n584bar;
  wire n585bar;
  wire n586bar;
  wire n587bar;
  wire n588bar;
  wire n589bar;
  wire n590bar;
  wire n591bar;
  wire n592bar;
  wire n593bar;
  wire n594bar;
  wire n595bar;
  wire n596bar;
  wire n597bar;
  wire n598bar;
  wire n599bar;
  wire n600bar;
  wire n601bar;
  wire n602bar;
  wire n603bar;
  wire n604bar;
  wire n605bar;
  wire n606bar;
  wire n607bar;
  wire n608bar;
  wire n609bar;
  wire n610bar;
  wire n611bar;
  wire n612bar;
  wire n613bar;
  wire n614bar;
  wire n615bar;
  wire n616bar;
  wire n617bar;
  wire n618bar;
  wire n619bar;
  wire n620bar;
  wire n621bar;
  wire n622bar;
  wire n623bar;
  wire n624bar;
  wire n625bar;
  wire n626bar;
  wire n627bar;
  wire n628bar;
  wire n629bar;
  wire n630bar;
  wire n631bar;
  wire n632bar;
  wire n633bar;
  wire n634bar;
  wire n635bar;
  wire n636bar;
  wire n637bar;
  wire n638bar;
  wire n639bar;
  wire n640bar;
  wire n641bar;
  wire n642bar;
  wire n643bar;
  wire n644bar;
  wire n645bar;
  wire n646bar;
  wire n647bar;
  wire n648bar;
  wire n649bar;
  wire n650bar;
  wire n651bar;
  wire n652bar;
  wire n653bar;
  wire n654bar;
  wire n655bar;
  wire n656bar;
  wire n657bar;
  wire n658bar;
  wire n659bar;
  wire n660bar;
  wire n661bar;
  wire n662bar;
  wire n663bar;
  wire n664bar;
  wire n665bar;
  wire n666bar;
  wire n667bar;
  wire n668bar;
  wire n669bar;
  wire n670bar;
  wire n671bar;
  wire n672bar;
  wire n673bar;
  wire n674bar;
  wire n675bar;
  wire n676bar;
  wire n677bar;
  wire n678bar;
  wire n679bar;
  wire n680bar;
  wire n681bar;
  wire n682bar;
  wire n683bar;
  wire n684bar;
  wire n685bar;
  wire n686bar;
  wire n687bar;
  wire n688bar;
  wire n689bar;
  wire n690bar;
  wire n691bar;
  wire n692bar;
  wire n693bar;
  wire n694bar;
  wire n695bar;
  wire n696bar;
  wire n697bar;
  wire n698bar;
  wire n699bar;
  wire n700bar;
  wire n701bar;
  wire n702bar;
  wire n703bar;
  wire n704bar;
  wire n705bar;
  wire n706bar;
  wire n707bar;
  wire n708bar;
  wire n709bar;
  wire n710bar;
  wire n711bar;
  wire n712bar;
  wire n713bar;
  wire n714bar;
  wire n715bar;
  wire n716bar;
  wire n717bar;
  wire n718bar;
  wire n719bar;
  wire n720bar;
  wire n721bar;
  wire n722bar;
  wire n723bar;
  wire n724bar;
  wire n725bar;
  wire n726bar;
  wire n727bar;
  wire n728bar;
  wire n729bar;
  wire n730bar;
  wire n731bar;
  wire n732bar;
  wire n733bar;
  wire n734bar;
  wire n735bar;
  wire n736bar;
  wire n737bar;
  wire n738bar;
  wire n739bar;
  wire n740bar;
  wire n741bar;
  wire n742bar;
  wire n743bar;
  wire n744bar;
  wire n745bar;
  wire n746bar;
  wire n747bar;
  wire n748bar;
  wire n749bar;
  wire n750bar;
  wire n751bar;
  wire n752bar;
  wire n753bar;
  wire n754bar;
  wire n755bar;
  wire n756bar;
  wire n757bar;
  wire n758bar;
  wire n759bar;
  wire n760bar;
  wire n761bar;
  wire n762bar;
  wire n763bar;
  wire n764bar;
  wire n765bar;
  wire n766bar;
  wire n767bar;
  wire n768bar;
  wire n769bar;
  wire n770bar;
  wire n771bar;
  wire n772bar;
  wire n773bar;
  wire n774bar;
  wire n775bar;
  wire n776bar;
  wire n777bar;
  wire n778bar;
  wire n779bar;
  wire n780bar;
  wire n781bar;
  wire n782bar;
  wire n783bar;
  wire n784bar;
  wire n785bar;
  wire n786bar;
  wire n787bar;
  wire n788bar;
  wire n789bar;
  wire n790bar;
  wire n791bar;
  wire n792bar;
  wire n793bar;
  wire n794bar;
  wire n795bar;
  wire n796bar;
  wire n797bar;
  wire n798bar;
  wire n799bar;
  wire n800bar;
  wire n801bar;
  wire n802bar;
  wire n803bar;
  wire n804bar;
  wire n805bar;
  wire n806bar;
  wire n807bar;
  wire n808bar;
  wire n809bar;
  wire n810bar;
  wire n811bar;
  wire n812bar;
  wire n813bar;
  wire n814bar;
  wire n815bar;
  wire n816bar;
  wire n817bar;
  wire n818bar;
  wire n819bar;
  wire n820bar;
  wire n821bar;
  wire n822bar;
  wire n823bar;
  wire n824bar;
  wire n825bar;
  wire n826bar;
  wire n827bar;
  wire n828bar;
  wire n829bar;
  wire n830bar;
  wire n831bar;
  wire n832bar;
  wire n833bar;
  wire n834bar;
  wire n835bar;
  wire n836bar;
  wire n837bar;
  wire n838bar;
  wire n839bar;
  wire n840bar;
  wire n841bar;
  wire n842bar;
  wire n843bar;
  wire n844bar;
  wire n845bar;
  wire n846bar;
  wire n847bar;
  wire n848bar;
  wire n849bar;
  wire n850bar;
  wire n851bar;
  wire n852bar;
  wire n853bar;
  wire n854bar;
  wire n855bar;
  wire n856bar;
  wire n857bar;
  wire n858bar;
  wire n859bar;
  wire n860bar;
  wire n861bar;
  wire n862bar;
  wire n863bar;
  wire n864bar;
  wire n865bar;
  wire n866bar;
  wire n867bar;
  wire n868bar;
  wire n869bar;
  wire n870bar;
  wire n871bar;
  wire n872bar;
  wire n873bar;
  wire n874bar;
  wire n875bar;
  wire n876bar;
  wire n877bar;
  wire n878bar;
  wire n879bar;
  wire n880bar;
  wire n881bar;
  wire n882bar;
  wire n883bar;
  wire n884bar;
  wire n885bar;
  wire n886bar;
  wire n887bar;
  wire n888bar;
  wire n889bar;
  wire n890bar;
  wire n891bar;
  wire n892bar;
  wire n893bar;
  wire n894bar;
  wire n895bar;
  wire n896bar;
  wire n897bar;
  wire n898bar;
  wire n899bar;
  wire n900bar;
  wire n901bar;
  wire n902bar;
  wire n903bar;
  wire n904bar;
  wire n905bar;
  wire n906bar;
  wire n907bar;
  wire n908bar;
  wire n909bar;
  wire n910bar;
  wire n911bar;
  wire n912bar;
  wire n913bar;
  wire n914bar;
  wire n915bar;
  wire n916bar;
  wire n917bar;
  wire n918bar;
  wire n919bar;
  wire n920bar;
  wire n921bar;
  wire n922bar;
  wire n923bar;
  wire n924bar;
  wire n925bar;
  wire n926bar;
  wire n927bar;
  wire n928bar;
  wire n929bar;
  wire n930bar;
  wire n931bar;
  wire n932bar;
  wire n933bar;
  wire n934bar;
  wire n935bar;
  wire n936bar;
  wire n937bar;
  wire n938bar;
  wire n939bar;
  wire n940bar;
  wire n941bar;
  wire n942bar;
  wire n943bar;
  wire n944bar;
  wire n945bar;
  wire n946bar;
  wire n947bar;
  wire n948bar;
  wire n949bar;
  wire n950bar;
  wire n951bar;
  wire n952bar;
  wire n953bar;
  wire n954bar;
  wire n955bar;
  wire n956bar;
  wire n957bar;
  wire n958bar;
  wire n959bar;
  wire n960bar;
  wire n961bar;
  wire n962bar;
  wire n963bar;
  wire n964bar;
  wire n965bar;
  wire n966bar;
  wire n967bar;
  wire n968bar;
  wire n969bar;
  wire n970bar;
  wire n971bar;
  wire n972bar;
//wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];
  assign in_81bar = inbar[81];
  assign in_80bar = inbar[80];
  assign in_79bar = inbar[79];
  assign in_78bar = inbar[78];
  assign in_77bar = inbar[77];
  assign in_76bar = inbar[76];
  assign in_75bar = inbar[75];
  assign in_74bar = inbar[74];
  assign in_73bar = inbar[73];
  assign in_72bar = inbar[72];
  assign in_71bar = inbar[71];
  assign in_70bar = inbar[70];
  assign in_69bar = inbar[69];
  assign in_68bar = inbar[68];
  assign in_67bar = inbar[67];
  assign in_66bar = inbar[66];
  assign in_65bar = inbar[65];
  assign in_64bar = inbar[64];
  assign in_63bar = inbar[63];
  assign in_62bar = inbar[62];
  assign in_61bar = inbar[61];
  assign in_60bar = inbar[60];
  assign in_59bar = inbar[59];
  assign in_58bar = inbar[58];
  assign in_57bar = inbar[57];
  assign in_56bar = inbar[56];
  assign in_55bar = inbar[55];
  assign in_54bar = inbar[54];
  assign in_53bar = inbar[53];
  assign in_52bar = inbar[52];
  assign in_51bar = inbar[51];
  assign in_50bar = inbar[50];
  assign in_49bar = inbar[49];
  assign in_48bar = inbar[48];
  assign in_47bar = inbar[47];
  assign in_46bar = inbar[46];
  assign in_45bar = inbar[45];
  assign in_44bar = inbar[44];
  assign in_43bar = inbar[43];
  assign in_42bar = inbar[42];
  assign in_41bar = inbar[41];
  assign in_40bar = inbar[40];
  assign in_39bar = inbar[39];
  assign in_38bar = inbar[38];
  assign in_37bar = inbar[37];
  assign in_36bar = inbar[36];
  assign in_35bar = inbar[35];
  assign in_34bar = inbar[34];
  assign in_33bar = inbar[33];
  assign in_32bar = inbar[32];
  assign in_31bar = inbar[31];
  assign in_30bar = inbar[30];
  assign in_29bar = inbar[29];
  assign in_28bar = inbar[28];
  assign in_27bar = inbar[27];
  assign in_26bar = inbar[26];
  assign in_25bar = inbar[25];
  assign in_24bar = inbar[24];
  assign in_23bar = inbar[23];
  assign in_22bar = inbar[22];
  assign in_21bar = inbar[21];
  assign in_20bar = inbar[20];
  assign in_19bar = inbar[19];
  assign in_18bar = inbar[18];
  assign in_17bar = inbar[17];
  assign in_16bar = inbar[16];
  assign in_15bar = inbar[15];
  assign in_14bar = inbar[14];
  assign in_13bar = inbar[13];
  assign in_12bar = inbar[12];
  assign in_11bar = inbar[11];
  assign in_10bar = inbar[10];
  assign in_9bar = inbar[9];
  assign in_8bar = inbar[8];
  assign in_7bar = inbar[7];
  assign in_6bar = inbar[6];
  assign in_5bar = inbar[5];
  assign in_4bar = inbar[4];
  assign in_3bar = inbar[3];
  assign in_2bar = inbar[2];
  assign in_1bar = inbar[1];
  assign in_0bar = inbar[0];
//assign_done

  OR2_X1 U1 ( .A1(n972), .A2(n971), .ZN(out[7]) );
  AND2_X1 U1bar ( .A1(n972bar), .A2(n971bar), .ZN(outbar[7]) );
  OR2_X1 U2 ( .A1(n970), .A2(n969), .ZN(n971) );
  AND2_X1 U2bar ( .A1(n970bar), .A2(n969bar), .ZN(n971bar) );
  OR2_X1 U3 ( .A1(n968), .A2(n967), .ZN(n969) );
  AND2_X1 U3bar ( .A1(n968bar), .A2(n967bar), .ZN(n969bar) );
  OR2_X1 U4 ( .A1(n966), .A2(n965), .ZN(n967) );
  AND2_X1 U4bar ( .A1(n966bar), .A2(n965bar), .ZN(n967bar) );
  OR2_X1 U5 ( .A1(n964), .A2(n963), .ZN(n968) );
  AND2_X1 U5bar ( .A1(n964bar), .A2(n963bar), .ZN(n968bar) );
  OR2_X1 U6 ( .A1(in[116]), .A2(n962), .ZN(n963) );
  AND2_X1 U6bar ( .A1(inbar[116]), .A2(n962bar), .ZN(n963bar) );
  OR2_X1 U7 ( .A1(n961), .A2(n960), .ZN(n970) );
  AND2_X1 U7bar ( .A1(n961bar), .A2(n960bar), .ZN(n970bar) );
  OR2_X1 U8 ( .A1(in[150]), .A2(in[127]), .ZN(n960) );
  AND2_X1 U8bar ( .A1(inbar[150]), .A2(inbar[127]), .ZN(n960bar) );
  OR2_X1 U9 ( .A1(in[160]), .A2(n959), .ZN(n961) );
  AND2_X1 U9bar ( .A1(inbar[160]), .A2(n959bar), .ZN(n961bar) );
  OR2_X1 U10 ( .A1(in[252]), .A2(in[168]), .ZN(n959) );
  AND2_X1 U10bar ( .A1(inbar[252]), .A2(inbar[168]), .ZN(n959bar) );
  OR2_X1 U11 ( .A1(n958), .A2(n957), .ZN(n972) );
  AND2_X1 U11bar ( .A1(n958bar), .A2(n957bar), .ZN(n972bar) );
  OR2_X1 U12 ( .A1(n956), .A2(n955), .ZN(n957) );
  AND2_X1 U12bar ( .A1(n956bar), .A2(n955bar), .ZN(n957bar) );
  OR2_X1 U13 ( .A1(in_17), .A2(in[96]), .ZN(n955) );
  AND2_X1 U13bar ( .A1(in_17bar), .A2(inbar[96]), .ZN(n955bar) );
  OR2_X1 U14 ( .A1(in_23), .A2(n954), .ZN(n956) );
  AND2_X1 U14bar ( .A1(in_23bar), .A2(n954bar), .ZN(n956bar) );
  OR2_X1 U15 ( .A1(in_31), .A2(in_26), .ZN(n954) );
  AND2_X1 U15bar ( .A1(in_31bar), .A2(in_26bar), .ZN(n954bar) );
  OR2_X1 U16 ( .A1(n953), .A2(n952), .ZN(n958) );
  AND2_X1 U16bar ( .A1(n953bar), .A2(n952bar), .ZN(n958bar) );
  OR2_X1 U17 ( .A1(in_58), .A2(in_4), .ZN(n952) );
  AND2_X1 U17bar ( .A1(in_58bar), .A2(in_4bar), .ZN(n952bar) );
  OR2_X1 U18 ( .A1(in_59), .A2(n951), .ZN(n953) );
  AND2_X1 U18bar ( .A1(in_59bar), .A2(n951bar), .ZN(n953bar) );
  OR2_X1 U19 ( .A1(in_71), .A2(in_62), .ZN(n951) );
  AND2_X1 U19bar ( .A1(in_71bar), .A2(in_62bar), .ZN(n951bar) );
  OR2_X1 U20 ( .A1(n950), .A2(n949), .ZN(out[6]) );
  AND2_X1 U20bar ( .A1(n950bar), .A2(n949bar), .ZN(outbar[6]) );
  OR2_X1 U21 ( .A1(n948), .A2(n947), .ZN(n949) );
  AND2_X1 U21bar ( .A1(n948bar), .A2(n947bar), .ZN(n949bar) );
  OR2_X1 U22 ( .A1(n946), .A2(n945), .ZN(n947) );
  AND2_X1 U22bar ( .A1(n946bar), .A2(n945bar), .ZN(n947bar) );
  OR2_X1 U23 ( .A1(n944), .A2(n943), .ZN(n945) );
  AND2_X1 U23bar ( .A1(n944bar), .A2(n943bar), .ZN(n945bar) );
  OR2_X1 U24 ( .A1(n942), .A2(n941), .ZN(n946) );
  AND2_X1 U24bar ( .A1(n942bar), .A2(n941bar), .ZN(n946bar) );
  OR2_X1 U25 ( .A1(in[101]), .A2(n940), .ZN(n941) );
  AND2_X1 U25bar ( .A1(inbar[101]), .A2(n940bar), .ZN(n941bar) );
  OR2_X1 U26 ( .A1(n939), .A2(n938), .ZN(n948) );
  AND2_X1 U26bar ( .A1(n939bar), .A2(n938bar), .ZN(n948bar) );
  OR2_X1 U27 ( .A1(in[114]), .A2(in[104]), .ZN(n938) );
  AND2_X1 U27bar ( .A1(inbar[114]), .A2(inbar[104]), .ZN(n938bar) );
  OR2_X1 U28 ( .A1(in[128]), .A2(n937), .ZN(n939) );
  AND2_X1 U28bar ( .A1(inbar[128]), .A2(n937bar), .ZN(n939bar) );
  OR2_X1 U29 ( .A1(in[136]), .A2(in[134]), .ZN(n937) );
  AND2_X1 U29bar ( .A1(inbar[136]), .A2(inbar[134]), .ZN(n937bar) );
  OR2_X1 U30 ( .A1(n936), .A2(n935), .ZN(n950) );
  AND2_X1 U30bar ( .A1(n936bar), .A2(n935bar), .ZN(n950bar) );
  OR2_X1 U31 ( .A1(n934), .A2(n933), .ZN(n935) );
  AND2_X1 U31bar ( .A1(n934bar), .A2(n933bar), .ZN(n935bar) );
  OR2_X1 U32 ( .A1(in[177]), .A2(in[164]), .ZN(n933) );
  AND2_X1 U32bar ( .A1(inbar[177]), .A2(inbar[164]), .ZN(n933bar) );
  OR2_X1 U33 ( .A1(in[212]), .A2(n932), .ZN(n934) );
  AND2_X1 U33bar ( .A1(inbar[212]), .A2(n932bar), .ZN(n934bar) );
  OR2_X1 U34 ( .A1(in[248]), .A2(in[221]), .ZN(n932) );
  AND2_X1 U34bar ( .A1(inbar[248]), .A2(inbar[221]), .ZN(n932bar) );
  OR2_X1 U35 ( .A1(n931), .A2(n930), .ZN(n936) );
  AND2_X1 U35bar ( .A1(n931bar), .A2(n930bar), .ZN(n936bar) );
  OR2_X1 U36 ( .A1(in_18), .A2(in[93]), .ZN(n930) );
  AND2_X1 U36bar ( .A1(in_18bar), .A2(inbar[93]), .ZN(n930bar) );
  OR2_X1 U37 ( .A1(in_31), .A2(n929), .ZN(n931) );
  AND2_X1 U37bar ( .A1(in_31bar), .A2(n929bar), .ZN(n931bar) );
  OR2_X1 U38 ( .A1(in_7), .A2(in_39), .ZN(n929) );
  AND2_X1 U38bar ( .A1(in_7bar), .A2(in_39bar), .ZN(n929bar) );
  OR2_X1 U39 ( .A1(n928), .A2(n927), .ZN(out[5]) );
  AND2_X1 U39bar ( .A1(n928bar), .A2(n927bar), .ZN(outbar[5]) );
  OR2_X1 U40 ( .A1(n926), .A2(n925), .ZN(n927) );
  AND2_X1 U40bar ( .A1(n926bar), .A2(n925bar), .ZN(n927bar) );
  OR2_X1 U41 ( .A1(n924), .A2(n923), .ZN(n925) );
  AND2_X1 U41bar ( .A1(n924bar), .A2(n923bar), .ZN(n925bar) );
  OR2_X1 U42 ( .A1(n922), .A2(n921), .ZN(n923) );
  AND2_X1 U42bar ( .A1(n922bar), .A2(n921bar), .ZN(n923bar) );
  OR2_X1 U43 ( .A1(n940), .A2(n920), .ZN(n924) );
  AND2_X1 U43bar ( .A1(n940bar), .A2(n920bar), .ZN(n924bar) );
  OR2_X1 U44 ( .A1(in[111]), .A2(n919), .ZN(n920) );
  AND2_X1 U44bar ( .A1(inbar[111]), .A2(n919bar), .ZN(n920bar) );
  OR2_X1 U45 ( .A1(n918), .A2(n917), .ZN(n940) );
  AND2_X1 U45bar ( .A1(n918bar), .A2(n917bar), .ZN(n940bar) );
  OR2_X1 U46 ( .A1(n916), .A2(n915), .ZN(n917) );
  AND2_X1 U46bar ( .A1(n916bar), .A2(n915bar), .ZN(n917bar) );
  OR2_X1 U47 ( .A1(n914), .A2(n913), .ZN(n915) );
  AND2_X1 U47bar ( .A1(n914bar), .A2(n913bar), .ZN(n915bar) );
  OR2_X1 U48 ( .A1(in[140]), .A2(in[131]), .ZN(n913) );
  AND2_X1 U48bar ( .A1(inbar[140]), .A2(inbar[131]), .ZN(n913bar) );
  OR2_X1 U49 ( .A1(in[160]), .A2(in[144]), .ZN(n914) );
  AND2_X1 U49bar ( .A1(inbar[160]), .A2(inbar[144]), .ZN(n914bar) );
  OR2_X1 U50 ( .A1(n912), .A2(n911), .ZN(n916) );
  AND2_X1 U50bar ( .A1(n912bar), .A2(n911bar), .ZN(n916bar) );
  OR2_X1 U51 ( .A1(in[179]), .A2(in[174]), .ZN(n911) );
  AND2_X1 U51bar ( .A1(inbar[179]), .A2(inbar[174]), .ZN(n911bar) );
  OR2_X1 U52 ( .A1(in[188]), .A2(in[184]), .ZN(n912) );
  AND2_X1 U52bar ( .A1(inbar[188]), .A2(inbar[184]), .ZN(n912bar) );
  OR2_X1 U53 ( .A1(n910), .A2(n909), .ZN(n918) );
  AND2_X1 U53bar ( .A1(n910bar), .A2(n909bar), .ZN(n918bar) );
  OR2_X1 U54 ( .A1(n908), .A2(n907), .ZN(n909) );
  AND2_X1 U54bar ( .A1(n908bar), .A2(n907bar), .ZN(n909bar) );
  OR2_X1 U55 ( .A1(in[216]), .A2(in[200]), .ZN(n907) );
  AND2_X1 U55bar ( .A1(inbar[216]), .A2(inbar[200]), .ZN(n907bar) );
  OR2_X1 U56 ( .A1(in[228]), .A2(in[224]), .ZN(n908) );
  AND2_X1 U56bar ( .A1(inbar[228]), .A2(inbar[224]), .ZN(n908bar) );
  OR2_X1 U57 ( .A1(n906), .A2(n905), .ZN(n910) );
  AND2_X1 U57bar ( .A1(n906bar), .A2(n905bar), .ZN(n910bar) );
  OR2_X1 U58 ( .A1(in[247]), .A2(in[235]), .ZN(n905) );
  AND2_X1 U58bar ( .A1(inbar[247]), .A2(inbar[235]), .ZN(n905bar) );
  OR2_X1 U59 ( .A1(in_42), .A2(in[83]), .ZN(n906) );
  AND2_X1 U59bar ( .A1(in_42bar), .A2(inbar[83]), .ZN(n906bar) );
  OR2_X1 U60 ( .A1(n904), .A2(n903), .ZN(n926) );
  AND2_X1 U60bar ( .A1(n904bar), .A2(n903bar), .ZN(n926bar) );
  OR2_X1 U61 ( .A1(in[166]), .A2(in[123]), .ZN(n903) );
  AND2_X1 U61bar ( .A1(inbar[166]), .A2(inbar[123]), .ZN(n903bar) );
  OR2_X1 U62 ( .A1(in[170]), .A2(n902), .ZN(n904) );
  AND2_X1 U62bar ( .A1(inbar[170]), .A2(n902bar), .ZN(n904bar) );
  OR2_X1 U63 ( .A1(in[194]), .A2(in[183]), .ZN(n902) );
  AND2_X1 U63bar ( .A1(inbar[194]), .A2(inbar[183]), .ZN(n902bar) );
  OR2_X1 U64 ( .A1(n901), .A2(n900), .ZN(n928) );
  AND2_X1 U64bar ( .A1(n901bar), .A2(n900bar), .ZN(n928bar) );
  OR2_X1 U65 ( .A1(n899), .A2(n898), .ZN(n900) );
  AND2_X1 U65bar ( .A1(n899bar), .A2(n898bar), .ZN(n900bar) );
  OR2_X1 U66 ( .A1(in[241]), .A2(in[238]), .ZN(n898) );
  AND2_X1 U66bar ( .A1(inbar[241]), .A2(inbar[238]), .ZN(n898bar) );
  OR2_X1 U67 ( .A1(in[250]), .A2(n897), .ZN(n899) );
  AND2_X1 U67bar ( .A1(inbar[250]), .A2(n897bar), .ZN(n899bar) );
  OR2_X1 U68 ( .A1(in_24), .A2(in[84]), .ZN(n897) );
  AND2_X1 U68bar ( .A1(in_24bar), .A2(inbar[84]), .ZN(n897bar) );
  OR2_X1 U69 ( .A1(n896), .A2(n895), .ZN(n901) );
  AND2_X1 U69bar ( .A1(n896bar), .A2(n895bar), .ZN(n901bar) );
  OR2_X1 U70 ( .A1(in_41), .A2(in_29), .ZN(n895) );
  AND2_X1 U70bar ( .A1(in_41bar), .A2(in_29bar), .ZN(n895bar) );
  OR2_X1 U71 ( .A1(in_66), .A2(n894), .ZN(n896) );
  AND2_X1 U71bar ( .A1(in_66bar), .A2(n894bar), .ZN(n896bar) );
  OR2_X1 U72 ( .A1(in_76), .A2(in_71), .ZN(n894) );
  AND2_X1 U72bar ( .A1(in_76bar), .A2(in_71bar), .ZN(n894bar) );
  OR2_X1 U73 ( .A1(n893), .A2(n892), .ZN(out[4]) );
  AND2_X1 U73bar ( .A1(n893bar), .A2(n892bar), .ZN(outbar[4]) );
  OR2_X1 U74 ( .A1(n891), .A2(n890), .ZN(n892) );
  AND2_X1 U74bar ( .A1(n891bar), .A2(n890bar), .ZN(n892bar) );
  OR2_X1 U75 ( .A1(n889), .A2(n888), .ZN(n890) );
  AND2_X1 U75bar ( .A1(n889bar), .A2(n888bar), .ZN(n890bar) );
  OR2_X1 U76 ( .A1(n922), .A2(n887), .ZN(n888) );
  AND2_X1 U76bar ( .A1(n922bar), .A2(n887bar), .ZN(n888bar) );
  OR2_X1 U77 ( .A1(n886), .A2(n885), .ZN(n922) );
  AND2_X1 U77bar ( .A1(n886bar), .A2(n885bar), .ZN(n922bar) );
  OR2_X1 U78 ( .A1(n884), .A2(n883), .ZN(n885) );
  AND2_X1 U78bar ( .A1(n884bar), .A2(n883bar), .ZN(n885bar) );
  OR2_X1 U79 ( .A1(n882), .A2(n881), .ZN(n883) );
  AND2_X1 U79bar ( .A1(n882bar), .A2(n881bar), .ZN(n883bar) );
  OR2_X1 U80 ( .A1(in[118]), .A2(in[109]), .ZN(n881) );
  AND2_X1 U80bar ( .A1(inbar[118]), .A2(inbar[109]), .ZN(n881bar) );
  OR2_X1 U81 ( .A1(in[139]), .A2(in[120]), .ZN(n882) );
  AND2_X1 U81bar ( .A1(inbar[139]), .A2(inbar[120]), .ZN(n882bar) );
  OR2_X1 U82 ( .A1(n880), .A2(n879), .ZN(n884) );
  AND2_X1 U82bar ( .A1(n880bar), .A2(n879bar), .ZN(n884bar) );
  OR2_X1 U83 ( .A1(in[198]), .A2(in[154]), .ZN(n879) );
  AND2_X1 U83bar ( .A1(inbar[198]), .A2(inbar[154]), .ZN(n879bar) );
  OR2_X1 U84 ( .A1(in[210]), .A2(in[205]), .ZN(n880) );
  AND2_X1 U84bar ( .A1(inbar[210]), .A2(inbar[205]), .ZN(n880bar) );
  OR2_X1 U85 ( .A1(n878), .A2(n877), .ZN(n886) );
  AND2_X1 U85bar ( .A1(n878bar), .A2(n877bar), .ZN(n886bar) );
  OR2_X1 U86 ( .A1(n876), .A2(n875), .ZN(n877) );
  AND2_X1 U86bar ( .A1(n876bar), .A2(n875bar), .ZN(n877bar) );
  OR2_X1 U87 ( .A1(in[219]), .A2(in[217]), .ZN(n875) );
  AND2_X1 U87bar ( .A1(inbar[219]), .A2(inbar[217]), .ZN(n875bar) );
  OR2_X1 U88 ( .A1(in[86]), .A2(in[252]), .ZN(n876) );
  AND2_X1 U88bar ( .A1(inbar[86]), .A2(inbar[252]), .ZN(n876bar) );
  OR2_X1 U89 ( .A1(n874), .A2(n873), .ZN(n878) );
  AND2_X1 U89bar ( .A1(n874bar), .A2(n873bar), .ZN(n878bar) );
  OR2_X1 U90 ( .A1(in_40), .A2(in[91]), .ZN(n873) );
  AND2_X1 U90bar ( .A1(in_40bar), .A2(inbar[91]), .ZN(n873bar) );
  OR2_X1 U91 ( .A1(in_8), .A2(in_46), .ZN(n874) );
  AND2_X1 U91bar ( .A1(in_8bar), .A2(in_46bar), .ZN(n874bar) );
  OR2_X1 U92 ( .A1(n872), .A2(n871), .ZN(n889) );
  AND2_X1 U92bar ( .A1(n872bar), .A2(n871bar), .ZN(n889bar) );
  OR2_X1 U93 ( .A1(in[117]), .A2(n943), .ZN(n871) );
  AND2_X1 U93bar ( .A1(inbar[117]), .A2(n943bar), .ZN(n871bar) );
  OR2_X1 U94 ( .A1(n870), .A2(n869), .ZN(n943) );
  AND2_X1 U94bar ( .A1(n870bar), .A2(n869bar), .ZN(n943bar) );
  OR2_X1 U95 ( .A1(n868), .A2(n867), .ZN(n869) );
  AND2_X1 U95bar ( .A1(n868bar), .A2(n867bar), .ZN(n869bar) );
  OR2_X1 U96 ( .A1(n866), .A2(n865), .ZN(n867) );
  AND2_X1 U96bar ( .A1(n866bar), .A2(n865bar), .ZN(n867bar) );
  OR2_X1 U97 ( .A1(n864), .A2(n863), .ZN(n865) );
  AND2_X1 U97bar ( .A1(n864bar), .A2(n863bar), .ZN(n865bar) );
  OR2_X1 U98 ( .A1(in[108]), .A2(n919), .ZN(n866) );
  AND2_X1 U98bar ( .A1(inbar[108]), .A2(n919bar), .ZN(n866bar) );
  OR2_X1 U99 ( .A1(n862), .A2(n861), .ZN(n919) );
  AND2_X1 U99bar ( .A1(n862bar), .A2(n861bar), .ZN(n919bar) );
  OR2_X1 U100 ( .A1(n860), .A2(n859), .ZN(n861) );
  AND2_X1 U100bar ( .A1(n860bar), .A2(n859bar), .ZN(n861bar) );
  OR2_X1 U101 ( .A1(n858), .A2(n857), .ZN(n859) );
  AND2_X1 U101bar ( .A1(n858bar), .A2(n857bar), .ZN(n859bar) );
  OR2_X1 U102 ( .A1(in[119]), .A2(in[105]), .ZN(n857) );
  AND2_X1 U102bar ( .A1(inbar[119]), .A2(inbar[105]), .ZN(n857bar) );
  OR2_X1 U103 ( .A1(in[186]), .A2(in[175]), .ZN(n858) );
  AND2_X1 U103bar ( .A1(inbar[186]), .A2(inbar[175]), .ZN(n858bar) );
  OR2_X1 U104 ( .A1(n856), .A2(n855), .ZN(n860) );
  AND2_X1 U104bar ( .A1(n856bar), .A2(n855bar), .ZN(n860bar) );
  OR2_X1 U105 ( .A1(in[202]), .A2(in[193]), .ZN(n855) );
  AND2_X1 U105bar ( .A1(inbar[202]), .A2(inbar[193]), .ZN(n855bar) );
  OR2_X1 U106 ( .A1(in[225]), .A2(in[208]), .ZN(n856) );
  AND2_X1 U106bar ( .A1(inbar[225]), .A2(inbar[208]), .ZN(n856bar) );
  OR2_X1 U107 ( .A1(n854), .A2(n853), .ZN(n862) );
  AND2_X1 U107bar ( .A1(n854bar), .A2(n853bar), .ZN(n862bar) );
  OR2_X1 U108 ( .A1(n852), .A2(n851), .ZN(n853) );
  AND2_X1 U108bar ( .A1(n852bar), .A2(n851bar), .ZN(n853bar) );
  OR2_X1 U109 ( .A1(in_1), .A2(in[85]), .ZN(n851) );
  AND2_X1 U109bar ( .A1(in_1bar), .A2(inbar[85]), .ZN(n851bar) );
  OR2_X1 U110 ( .A1(in_23), .A2(in_19), .ZN(n852) );
  AND2_X1 U110bar ( .A1(in_23bar), .A2(in_19bar), .ZN(n852bar) );
  OR2_X1 U111 ( .A1(n850), .A2(n849), .ZN(n854) );
  AND2_X1 U111bar ( .A1(n850bar), .A2(n849bar), .ZN(n854bar) );
  OR2_X1 U112 ( .A1(in_43), .A2(in_33), .ZN(n849) );
  AND2_X1 U112bar ( .A1(in_43bar), .A2(in_33bar), .ZN(n849bar) );
  OR2_X1 U113 ( .A1(in_63), .A2(in_44), .ZN(n850) );
  AND2_X1 U113bar ( .A1(in_63bar), .A2(in_44bar), .ZN(n850bar) );
  OR2_X1 U114 ( .A1(n848), .A2(n847), .ZN(n868) );
  AND2_X1 U114bar ( .A1(n848bar), .A2(n847bar), .ZN(n868bar) );
  OR2_X1 U115 ( .A1(in[141]), .A2(in[112]), .ZN(n847) );
  AND2_X1 U115bar ( .A1(inbar[141]), .A2(inbar[112]), .ZN(n847bar) );
  OR2_X1 U116 ( .A1(in[147]), .A2(n846), .ZN(n848) );
  AND2_X1 U116bar ( .A1(inbar[147]), .A2(n846bar), .ZN(n848bar) );
  OR2_X1 U117 ( .A1(in[181]), .A2(in[167]), .ZN(n846) );
  AND2_X1 U117bar ( .A1(inbar[181]), .A2(inbar[167]), .ZN(n846bar) );
  OR2_X1 U118 ( .A1(n845), .A2(n844), .ZN(n870) );
  AND2_X1 U118bar ( .A1(n845bar), .A2(n844bar), .ZN(n870bar) );
  OR2_X1 U119 ( .A1(n843), .A2(n842), .ZN(n844) );
  AND2_X1 U119bar ( .A1(n843bar), .A2(n842bar), .ZN(n844bar) );
  OR2_X1 U120 ( .A1(in[229]), .A2(in[201]), .ZN(n842) );
  AND2_X1 U120bar ( .A1(inbar[229]), .A2(inbar[201]), .ZN(n842bar) );
  OR2_X1 U121 ( .A1(in[237]), .A2(n841), .ZN(n843) );
  AND2_X1 U121bar ( .A1(inbar[237]), .A2(n841bar), .ZN(n843bar) );
  OR2_X1 U122 ( .A1(in[94]), .A2(in[253]), .ZN(n841) );
  AND2_X1 U122bar ( .A1(inbar[94]), .A2(inbar[253]), .ZN(n841bar) );
  OR2_X1 U123 ( .A1(n840), .A2(n839), .ZN(n845) );
  AND2_X1 U123bar ( .A1(n840bar), .A2(n839bar), .ZN(n845bar) );
  OR2_X1 U124 ( .A1(in_21), .A2(in[96]), .ZN(n839) );
  AND2_X1 U124bar ( .A1(in_21bar), .A2(inbar[96]), .ZN(n839bar) );
  OR2_X1 U125 ( .A1(in_25), .A2(n838), .ZN(n840) );
  AND2_X1 U125bar ( .A1(in_25bar), .A2(n838bar), .ZN(n840bar) );
  OR2_X1 U126 ( .A1(in_81), .A2(in_45), .ZN(n838) );
  AND2_X1 U126bar ( .A1(in_81bar), .A2(in_45bar), .ZN(n838bar) );
  OR2_X1 U127 ( .A1(n837), .A2(n836), .ZN(n891) );
  AND2_X1 U127bar ( .A1(n837bar), .A2(n836bar), .ZN(n891bar) );
  OR2_X1 U128 ( .A1(in[142]), .A2(in[124]), .ZN(n836) );
  AND2_X1 U128bar ( .A1(inbar[142]), .A2(inbar[124]), .ZN(n836bar) );
  OR2_X1 U129 ( .A1(in[150]), .A2(n835), .ZN(n837) );
  AND2_X1 U129bar ( .A1(inbar[150]), .A2(n835bar), .ZN(n837bar) );
  OR2_X1 U130 ( .A1(in[172]), .A2(in[155]), .ZN(n835) );
  AND2_X1 U130bar ( .A1(inbar[172]), .A2(inbar[155]), .ZN(n835bar) );
  OR2_X1 U131 ( .A1(n834), .A2(n833), .ZN(n893) );
  AND2_X1 U131bar ( .A1(n834bar), .A2(n833bar), .ZN(n893bar) );
  OR2_X1 U132 ( .A1(n832), .A2(n831), .ZN(n833) );
  AND2_X1 U132bar ( .A1(n832bar), .A2(n831bar), .ZN(n833bar) );
  OR2_X1 U133 ( .A1(in[196]), .A2(in[173]), .ZN(n831) );
  AND2_X1 U133bar ( .A1(inbar[196]), .A2(inbar[173]), .ZN(n831bar) );
  OR2_X1 U134 ( .A1(in[222]), .A2(n830), .ZN(n832) );
  AND2_X1 U134bar ( .A1(inbar[222]), .A2(n830bar), .ZN(n832bar) );
  OR2_X1 U135 ( .A1(in[227]), .A2(in[226]), .ZN(n830) );
  AND2_X1 U135bar ( .A1(inbar[227]), .A2(inbar[226]), .ZN(n830bar) );
  OR2_X1 U136 ( .A1(n829), .A2(n828), .ZN(n834) );
  AND2_X1 U136bar ( .A1(n829bar), .A2(n828bar), .ZN(n834bar) );
  OR2_X1 U137 ( .A1(in[249]), .A2(in[231]), .ZN(n828) );
  AND2_X1 U137bar ( .A1(inbar[249]), .A2(inbar[231]), .ZN(n828bar) );
  OR2_X1 U138 ( .A1(in_28), .A2(n827), .ZN(n829) );
  AND2_X1 U138bar ( .A1(in_28bar), .A2(n827bar), .ZN(n829bar) );
  OR2_X1 U139 ( .A1(in_52), .A2(in_47), .ZN(n827) );
  AND2_X1 U139bar ( .A1(in_52bar), .A2(in_47bar), .ZN(n827bar) );
  OR2_X1 U140 ( .A1(n826), .A2(n825), .ZN(out[3]) );
  AND2_X1 U140bar ( .A1(n826bar), .A2(n825bar), .ZN(outbar[3]) );
  OR2_X1 U141 ( .A1(n824), .A2(n823), .ZN(n825) );
  AND2_X1 U141bar ( .A1(n824bar), .A2(n823bar), .ZN(n825bar) );
  OR2_X1 U142 ( .A1(n822), .A2(n821), .ZN(n823) );
  AND2_X1 U142bar ( .A1(n822bar), .A2(n821bar), .ZN(n823bar) );
  OR2_X1 U143 ( .A1(n820), .A2(n819), .ZN(n821) );
  AND2_X1 U143bar ( .A1(n820bar), .A2(n819bar), .ZN(n821bar) );
  OR2_X1 U144 ( .A1(n964), .A2(n818), .ZN(n822) );
  AND2_X1 U144bar ( .A1(n964bar), .A2(n818bar), .ZN(n822bar) );
  OR2_X1 U145 ( .A1(in[118]), .A2(n817), .ZN(n818) );
  AND2_X1 U145bar ( .A1(inbar[118]), .A2(n817bar), .ZN(n818bar) );
  OR2_X1 U146 ( .A1(n816), .A2(n815), .ZN(n964) );
  AND2_X1 U146bar ( .A1(n816bar), .A2(n815bar), .ZN(n964bar) );
  OR2_X1 U147 ( .A1(n814), .A2(n813), .ZN(n815) );
  AND2_X1 U147bar ( .A1(n814bar), .A2(n813bar), .ZN(n815bar) );
  OR2_X1 U148 ( .A1(n812), .A2(n811), .ZN(n813) );
  AND2_X1 U148bar ( .A1(n812bar), .A2(n811bar), .ZN(n813bar) );
  OR2_X1 U149 ( .A1(in[122]), .A2(in[111]), .ZN(n811) );
  AND2_X1 U149bar ( .A1(inbar[122]), .A2(inbar[111]), .ZN(n811bar) );
  OR2_X1 U150 ( .A1(in[154]), .A2(in[151]), .ZN(n812) );
  AND2_X1 U150bar ( .A1(inbar[154]), .A2(inbar[151]), .ZN(n812bar) );
  OR2_X1 U151 ( .A1(n810), .A2(n809), .ZN(n814) );
  AND2_X1 U151bar ( .A1(n810bar), .A2(n809bar), .ZN(n814bar) );
  OR2_X1 U152 ( .A1(in[187]), .A2(in[177]), .ZN(n809) );
  AND2_X1 U152bar ( .A1(inbar[187]), .A2(inbar[177]), .ZN(n809bar) );
  OR2_X1 U153 ( .A1(in[200]), .A2(in[192]), .ZN(n810) );
  AND2_X1 U153bar ( .A1(inbar[200]), .A2(inbar[192]), .ZN(n810bar) );
  OR2_X1 U154 ( .A1(n808), .A2(n807), .ZN(n816) );
  AND2_X1 U154bar ( .A1(n808bar), .A2(n807bar), .ZN(n816bar) );
  OR2_X1 U155 ( .A1(n806), .A2(n805), .ZN(n807) );
  AND2_X1 U155bar ( .A1(n806bar), .A2(n805bar), .ZN(n807bar) );
  OR2_X1 U156 ( .A1(in[225]), .A2(in[207]), .ZN(n805) );
  AND2_X1 U156bar ( .A1(inbar[225]), .A2(inbar[207]), .ZN(n805bar) );
  OR2_X1 U157 ( .A1(in[98]), .A2(in[226]), .ZN(n806) );
  AND2_X1 U157bar ( .A1(inbar[98]), .A2(inbar[226]), .ZN(n806bar) );
  OR2_X1 U158 ( .A1(n804), .A2(n803), .ZN(n808) );
  AND2_X1 U158bar ( .A1(n804bar), .A2(n803bar), .ZN(n808bar) );
  OR2_X1 U159 ( .A1(in_20), .A2(in_16), .ZN(n803) );
  AND2_X1 U159bar ( .A1(in_20bar), .A2(in_16bar), .ZN(n803bar) );
  OR2_X1 U160 ( .A1(in_55), .A2(in_45), .ZN(n804) );
  AND2_X1 U160bar ( .A1(in_55bar), .A2(in_45bar), .ZN(n804bar) );
  OR2_X1 U161 ( .A1(n802), .A2(n801), .ZN(n824) );
  AND2_X1 U161bar ( .A1(n802bar), .A2(n801bar), .ZN(n824bar) );
  OR2_X1 U162 ( .A1(in[162]), .A2(in[149]), .ZN(n801) );
  AND2_X1 U162bar ( .A1(inbar[162]), .A2(inbar[149]), .ZN(n801bar) );
  OR2_X1 U163 ( .A1(in[163]), .A2(n800), .ZN(n802) );
  AND2_X1 U163bar ( .A1(inbar[163]), .A2(n800bar), .ZN(n802bar) );
  OR2_X1 U164 ( .A1(in[191]), .A2(in[189]), .ZN(n800) );
  AND2_X1 U164bar ( .A1(inbar[191]), .A2(inbar[189]), .ZN(n800bar) );
  OR2_X1 U165 ( .A1(n799), .A2(n798), .ZN(n826) );
  AND2_X1 U165bar ( .A1(n799bar), .A2(n798bar), .ZN(n826bar) );
  OR2_X1 U166 ( .A1(n797), .A2(n796), .ZN(n798) );
  AND2_X1 U166bar ( .A1(n797bar), .A2(n796bar), .ZN(n798bar) );
  OR2_X1 U167 ( .A1(in[212]), .A2(in[193]), .ZN(n796) );
  AND2_X1 U167bar ( .A1(inbar[212]), .A2(inbar[193]), .ZN(n796bar) );
  OR2_X1 U168 ( .A1(in[238]), .A2(n795), .ZN(n797) );
  AND2_X1 U168bar ( .A1(inbar[238]), .A2(n795bar), .ZN(n797bar) );
  OR2_X1 U169 ( .A1(in[88]), .A2(in[247]), .ZN(n795) );
  AND2_X1 U169bar ( .A1(inbar[88]), .A2(inbar[247]), .ZN(n795bar) );
  OR2_X1 U170 ( .A1(n794), .A2(n793), .ZN(n799) );
  AND2_X1 U170bar ( .A1(n794bar), .A2(n793bar), .ZN(n799bar) );
  OR2_X1 U171 ( .A1(in[94]), .A2(in[92]), .ZN(n793) );
  AND2_X1 U171bar ( .A1(inbar[94]), .A2(inbar[92]), .ZN(n793bar) );
  OR2_X1 U172 ( .A1(in_52), .A2(n792), .ZN(n794) );
  AND2_X1 U172bar ( .A1(in_52bar), .A2(n792bar), .ZN(n794bar) );
  OR2_X1 U173 ( .A1(in_70), .A2(in_67), .ZN(n792) );
  AND2_X1 U173bar ( .A1(in_70bar), .A2(in_67bar), .ZN(n792bar) );
  OR2_X1 U174 ( .A1(n791), .A2(n790), .ZN(out[2]) );
  AND2_X1 U174bar ( .A1(n791bar), .A2(n790bar), .ZN(outbar[2]) );
  OR2_X1 U175 ( .A1(n789), .A2(n788), .ZN(n790) );
  AND2_X1 U175bar ( .A1(n789bar), .A2(n788bar), .ZN(n790bar) );
  OR2_X1 U176 ( .A1(n787), .A2(n786), .ZN(n788) );
  AND2_X1 U176bar ( .A1(n787bar), .A2(n786bar), .ZN(n788bar) );
  OR2_X1 U177 ( .A1(n819), .A2(n785), .ZN(n786) );
  AND2_X1 U177bar ( .A1(n819bar), .A2(n785bar), .ZN(n786bar) );
  OR2_X1 U178 ( .A1(n784), .A2(n783), .ZN(n819) );
  AND2_X1 U178bar ( .A1(n784bar), .A2(n783bar), .ZN(n819bar) );
  OR2_X1 U179 ( .A1(n782), .A2(n781), .ZN(n783) );
  AND2_X1 U179bar ( .A1(n782bar), .A2(n781bar), .ZN(n783bar) );
  OR2_X1 U180 ( .A1(n780), .A2(n779), .ZN(n781) );
  AND2_X1 U180bar ( .A1(n780bar), .A2(n779bar), .ZN(n781bar) );
  OR2_X1 U181 ( .A1(n962), .A2(n778), .ZN(n779) );
  AND2_X1 U181bar ( .A1(n962bar), .A2(n778bar), .ZN(n779bar) );
  OR2_X1 U182 ( .A1(n777), .A2(n776), .ZN(n962) );
  AND2_X1 U182bar ( .A1(n777bar), .A2(n776bar), .ZN(n962bar) );
  OR2_X1 U183 ( .A1(n775), .A2(n774), .ZN(n776) );
  AND2_X1 U183bar ( .A1(n775bar), .A2(n774bar), .ZN(n776bar) );
  OR2_X1 U184 ( .A1(n773), .A2(n772), .ZN(n774) );
  AND2_X1 U184bar ( .A1(n773bar), .A2(n772bar), .ZN(n774bar) );
  OR2_X1 U185 ( .A1(in[131]), .A2(in[120]), .ZN(n772) );
  AND2_X1 U185bar ( .A1(inbar[131]), .A2(inbar[120]), .ZN(n772bar) );
  OR2_X1 U186 ( .A1(in[153]), .A2(in[147]), .ZN(n773) );
  AND2_X1 U186bar ( .A1(inbar[153]), .A2(inbar[147]), .ZN(n773bar) );
  OR2_X1 U187 ( .A1(n771), .A2(n770), .ZN(n775) );
  AND2_X1 U187bar ( .A1(n771bar), .A2(n770bar), .ZN(n775bar) );
  OR2_X1 U188 ( .A1(in[170]), .A2(in[156]), .ZN(n770) );
  AND2_X1 U188bar ( .A1(inbar[170]), .A2(inbar[156]), .ZN(n770bar) );
  OR2_X1 U189 ( .A1(in[223]), .A2(in[190]), .ZN(n771) );
  AND2_X1 U189bar ( .A1(inbar[223]), .A2(inbar[190]), .ZN(n771bar) );
  OR2_X1 U190 ( .A1(n769), .A2(n768), .ZN(n777) );
  AND2_X1 U190bar ( .A1(n769bar), .A2(n768bar), .ZN(n777bar) );
  OR2_X1 U191 ( .A1(n767), .A2(n766), .ZN(n768) );
  AND2_X1 U191bar ( .A1(n767bar), .A2(n766bar), .ZN(n768bar) );
  OR2_X1 U192 ( .A1(in[236]), .A2(in[230]), .ZN(n766) );
  AND2_X1 U192bar ( .A1(inbar[236]), .A2(inbar[230]), .ZN(n766bar) );
  OR2_X1 U193 ( .A1(in[85]), .A2(in[240]), .ZN(n767) );
  AND2_X1 U193bar ( .A1(inbar[85]), .A2(inbar[240]), .ZN(n767bar) );
  OR2_X1 U194 ( .A1(n765), .A2(n764), .ZN(n769) );
  AND2_X1 U194bar ( .A1(n765bar), .A2(n764bar), .ZN(n769bar) );
  OR2_X1 U195 ( .A1(in_12), .A2(in[90]), .ZN(n764) );
  AND2_X1 U195bar ( .A1(in_12bar), .A2(inbar[90]), .ZN(n764bar) );
  OR2_X1 U196 ( .A1(in_39), .A2(in_28), .ZN(n765) );
  AND2_X1 U196bar ( .A1(in_39bar), .A2(in_28bar), .ZN(n765bar) );
  OR2_X1 U197 ( .A1(in[109]), .A2(n763), .ZN(n780) );
  AND2_X1 U197bar ( .A1(inbar[109]), .A2(n763bar), .ZN(n780bar) );
  OR2_X1 U198 ( .A1(n762), .A2(n761), .ZN(n782) );
  AND2_X1 U198bar ( .A1(n762bar), .A2(n761bar), .ZN(n782bar) );
  OR2_X1 U199 ( .A1(in[138]), .A2(in[129]), .ZN(n761) );
  AND2_X1 U199bar ( .A1(inbar[138]), .A2(inbar[129]), .ZN(n761bar) );
  OR2_X1 U200 ( .A1(in[157]), .A2(n760), .ZN(n762) );
  AND2_X1 U200bar ( .A1(inbar[157]), .A2(n760bar), .ZN(n762bar) );
  OR2_X1 U201 ( .A1(in[182]), .A2(in[167]), .ZN(n760) );
  AND2_X1 U201bar ( .A1(inbar[182]), .A2(inbar[167]), .ZN(n760bar) );
  OR2_X1 U202 ( .A1(n759), .A2(n758), .ZN(n784) );
  AND2_X1 U202bar ( .A1(n759bar), .A2(n758bar), .ZN(n784bar) );
  OR2_X1 U203 ( .A1(n757), .A2(n756), .ZN(n758) );
  AND2_X1 U203bar ( .A1(n757bar), .A2(n756bar), .ZN(n758bar) );
  OR2_X1 U204 ( .A1(in[195]), .A2(in[184]), .ZN(n756) );
  AND2_X1 U204bar ( .A1(inbar[195]), .A2(inbar[184]), .ZN(n756bar) );
  OR2_X1 U205 ( .A1(in[196]), .A2(n755), .ZN(n757) );
  AND2_X1 U205bar ( .A1(inbar[196]), .A2(n755bar), .ZN(n757bar) );
  OR2_X1 U206 ( .A1(in[215]), .A2(in[209]), .ZN(n755) );
  AND2_X1 U206bar ( .A1(inbar[215]), .A2(inbar[209]), .ZN(n755bar) );
  OR2_X1 U207 ( .A1(n754), .A2(n753), .ZN(n759) );
  AND2_X1 U207bar ( .A1(n754bar), .A2(n753bar), .ZN(n759bar) );
  OR2_X1 U208 ( .A1(in[93]), .A2(in[233]), .ZN(n753) );
  AND2_X1 U208bar ( .A1(inbar[93]), .A2(inbar[233]), .ZN(n753bar) );
  OR2_X1 U209 ( .A1(in_1), .A2(n752), .ZN(n754) );
  AND2_X1 U209bar ( .A1(in_1bar), .A2(n752bar), .ZN(n754bar) );
  OR2_X1 U210 ( .A1(in_69), .A2(in_66), .ZN(n752) );
  AND2_X1 U210bar ( .A1(in_69bar), .A2(in_66bar), .ZN(n752bar) );
  OR2_X1 U211 ( .A1(n966), .A2(n751), .ZN(n787) );
  AND2_X1 U211bar ( .A1(n966bar), .A2(n751bar), .ZN(n787bar) );
  OR2_X1 U212 ( .A1(in[134]), .A2(n750), .ZN(n751) );
  AND2_X1 U212bar ( .A1(inbar[134]), .A2(n750bar), .ZN(n751bar) );
  OR2_X1 U213 ( .A1(n749), .A2(n748), .ZN(n966) );
  AND2_X1 U213bar ( .A1(n749bar), .A2(n748bar), .ZN(n966bar) );
  OR2_X1 U214 ( .A1(n747), .A2(n746), .ZN(n748) );
  AND2_X1 U214bar ( .A1(n747bar), .A2(n746bar), .ZN(n748bar) );
  OR2_X1 U215 ( .A1(n745), .A2(n744), .ZN(n746) );
  AND2_X1 U215bar ( .A1(n745bar), .A2(n744bar), .ZN(n746bar) );
  OR2_X1 U216 ( .A1(in[136]), .A2(in[121]), .ZN(n744) );
  AND2_X1 U216bar ( .A1(inbar[136]), .A2(inbar[121]), .ZN(n744bar) );
  OR2_X1 U217 ( .A1(in[186]), .A2(in[174]), .ZN(n745) );
  AND2_X1 U217bar ( .A1(inbar[186]), .A2(inbar[174]), .ZN(n745bar) );
  OR2_X1 U218 ( .A1(n743), .A2(n742), .ZN(n747) );
  AND2_X1 U218bar ( .A1(n743bar), .A2(n742bar), .ZN(n747bar) );
  OR2_X1 U219 ( .A1(in[198]), .A2(in[197]), .ZN(n742) );
  AND2_X1 U219bar ( .A1(inbar[198]), .A2(inbar[197]), .ZN(n742bar) );
  OR2_X1 U220 ( .A1(in[214]), .A2(in[199]), .ZN(n743) );
  AND2_X1 U220bar ( .A1(inbar[214]), .A2(inbar[199]), .ZN(n743bar) );
  OR2_X1 U221 ( .A1(n741), .A2(n740), .ZN(n749) );
  AND2_X1 U221bar ( .A1(n741bar), .A2(n740bar), .ZN(n749bar) );
  OR2_X1 U222 ( .A1(n739), .A2(n738), .ZN(n740) );
  AND2_X1 U222bar ( .A1(n739bar), .A2(n738bar), .ZN(n740bar) );
  OR2_X1 U223 ( .A1(in[231]), .A2(in[220]), .ZN(n738) );
  AND2_X1 U223bar ( .A1(inbar[231]), .A2(inbar[220]), .ZN(n738bar) );
  OR2_X1 U224 ( .A1(in_25), .A2(in[245]), .ZN(n739) );
  AND2_X1 U224bar ( .A1(in_25bar), .A2(inbar[245]), .ZN(n739bar) );
  OR2_X1 U225 ( .A1(n737), .A2(n736), .ZN(n741) );
  AND2_X1 U225bar ( .A1(n737bar), .A2(n736bar), .ZN(n741bar) );
  OR2_X1 U226 ( .A1(in_53), .A2(in_29), .ZN(n736) );
  AND2_X1 U226bar ( .A1(in_53bar), .A2(in_29bar), .ZN(n736bar) );
  OR2_X1 U227 ( .A1(in_79), .A2(in_74), .ZN(n737) );
  AND2_X1 U227bar ( .A1(in_79bar), .A2(in_74bar), .ZN(n737bar) );
  OR2_X1 U228 ( .A1(n735), .A2(n734), .ZN(n789) );
  AND2_X1 U228bar ( .A1(n735bar), .A2(n734bar), .ZN(n789bar) );
  OR2_X1 U229 ( .A1(in[152]), .A2(in[140]), .ZN(n734) );
  AND2_X1 U229bar ( .A1(inbar[152]), .A2(inbar[140]), .ZN(n734bar) );
  OR2_X1 U230 ( .A1(in[155]), .A2(n733), .ZN(n735) );
  AND2_X1 U230bar ( .A1(inbar[155]), .A2(n733bar), .ZN(n735bar) );
  OR2_X1 U231 ( .A1(in[166]), .A2(in[165]), .ZN(n733) );
  AND2_X1 U231bar ( .A1(inbar[166]), .A2(inbar[165]), .ZN(n733bar) );
  OR2_X1 U232 ( .A1(n732), .A2(n731), .ZN(n791) );
  AND2_X1 U232bar ( .A1(n732bar), .A2(n731bar), .ZN(n791bar) );
  OR2_X1 U233 ( .A1(n730), .A2(n729), .ZN(n731) );
  AND2_X1 U233bar ( .A1(n730bar), .A2(n729bar), .ZN(n731bar) );
  OR2_X1 U234 ( .A1(in[202]), .A2(in[185]), .ZN(n729) );
  AND2_X1 U234bar ( .A1(inbar[202]), .A2(inbar[185]), .ZN(n729bar) );
  OR2_X1 U235 ( .A1(in[211]), .A2(n728), .ZN(n730) );
  AND2_X1 U235bar ( .A1(inbar[211]), .A2(n728bar), .ZN(n730bar) );
  OR2_X1 U236 ( .A1(in[255]), .A2(in[253]), .ZN(n728) );
  AND2_X1 U236bar ( .A1(inbar[255]), .A2(inbar[253]), .ZN(n728bar) );
  OR2_X1 U237 ( .A1(n727), .A2(n726), .ZN(n732) );
  AND2_X1 U237bar ( .A1(n727bar), .A2(n726bar), .ZN(n732bar) );
  OR2_X1 U238 ( .A1(in_35), .A2(in_15), .ZN(n726) );
  AND2_X1 U238bar ( .A1(in_35bar), .A2(in_15bar), .ZN(n726bar) );
  OR2_X1 U239 ( .A1(in_36), .A2(n725), .ZN(n727) );
  AND2_X1 U239bar ( .A1(in_36bar), .A2(n725bar), .ZN(n727bar) );
  OR2_X1 U240 ( .A1(in_48), .A2(in_40), .ZN(n725) );
  AND2_X1 U240bar ( .A1(in_48bar), .A2(in_40bar), .ZN(n725bar) );
  OR2_X1 U241 ( .A1(n724), .A2(n723), .ZN(out[1]) );
  AND2_X1 U241bar ( .A1(n724bar), .A2(n723bar), .ZN(outbar[1]) );
  OR2_X1 U242 ( .A1(n722), .A2(n721), .ZN(n723) );
  AND2_X1 U242bar ( .A1(n722bar), .A2(n721bar), .ZN(n723bar) );
  OR2_X1 U243 ( .A1(n720), .A2(n719), .ZN(n721) );
  AND2_X1 U243bar ( .A1(n720bar), .A2(n719bar), .ZN(n721bar) );
  OR2_X1 U244 ( .A1(n921), .A2(n887), .ZN(n719) );
  AND2_X1 U244bar ( .A1(n921bar), .A2(n887bar), .ZN(n719bar) );
  OR2_X1 U245 ( .A1(n718), .A2(n717), .ZN(n887) );
  AND2_X1 U245bar ( .A1(n718bar), .A2(n717bar), .ZN(n887bar) );
  OR2_X1 U246 ( .A1(n716), .A2(n715), .ZN(n717) );
  AND2_X1 U246bar ( .A1(n716bar), .A2(n715bar), .ZN(n717bar) );
  OR2_X1 U247 ( .A1(n714), .A2(n713), .ZN(n715) );
  AND2_X1 U247bar ( .A1(n714bar), .A2(n713bar), .ZN(n715bar) );
  OR2_X1 U248 ( .A1(in[116]), .A2(in[110]), .ZN(n713) );
  AND2_X1 U248bar ( .A1(inbar[116]), .A2(inbar[110]), .ZN(n713bar) );
  OR2_X1 U249 ( .A1(in[133]), .A2(in[130]), .ZN(n714) );
  AND2_X1 U249bar ( .A1(inbar[133]), .A2(inbar[130]), .ZN(n714bar) );
  OR2_X1 U250 ( .A1(n712), .A2(n711), .ZN(n716) );
  AND2_X1 U250bar ( .A1(n712bar), .A2(n711bar), .ZN(n716bar) );
  OR2_X1 U251 ( .A1(in[203]), .A2(in[135]), .ZN(n711) );
  AND2_X1 U251bar ( .A1(inbar[203]), .A2(inbar[135]), .ZN(n711bar) );
  OR2_X1 U252 ( .A1(in[232]), .A2(in[223]), .ZN(n712) );
  AND2_X1 U252bar ( .A1(inbar[232]), .A2(inbar[223]), .ZN(n712bar) );
  OR2_X1 U253 ( .A1(n710), .A2(n709), .ZN(n718) );
  AND2_X1 U253bar ( .A1(n710bar), .A2(n709bar), .ZN(n718bar) );
  OR2_X1 U254 ( .A1(n708), .A2(n707), .ZN(n709) );
  AND2_X1 U254bar ( .A1(n708bar), .A2(n707bar), .ZN(n709bar) );
  OR2_X1 U255 ( .A1(in[255]), .A2(in[233]), .ZN(n707) );
  AND2_X1 U255bar ( .A1(inbar[255]), .A2(inbar[233]), .ZN(n707bar) );
  OR2_X1 U256 ( .A1(in_53), .A2(in_34), .ZN(n708) );
  AND2_X1 U256bar ( .A1(in_53bar), .A2(in_34bar), .ZN(n708bar) );
  OR2_X1 U257 ( .A1(n706), .A2(n705), .ZN(n710) );
  AND2_X1 U257bar ( .A1(n706bar), .A2(n705bar), .ZN(n710bar) );
  OR2_X1 U258 ( .A1(in_57), .A2(in_55), .ZN(n705) );
  AND2_X1 U258bar ( .A1(in_57bar), .A2(in_55bar), .ZN(n705bar) );
  OR2_X1 U259 ( .A1(in_68), .A2(in_67), .ZN(n706) );
  AND2_X1 U259bar ( .A1(in_68bar), .A2(in_67bar), .ZN(n706bar) );
  OR2_X1 U260 ( .A1(n704), .A2(n703), .ZN(n921) );
  AND2_X1 U260bar ( .A1(n704bar), .A2(n703bar), .ZN(n921bar) );
  OR2_X1 U261 ( .A1(n702), .A2(n701), .ZN(n703) );
  AND2_X1 U261bar ( .A1(n702bar), .A2(n701bar), .ZN(n703bar) );
  OR2_X1 U262 ( .A1(n700), .A2(n699), .ZN(n701) );
  AND2_X1 U262bar ( .A1(n700bar), .A2(n699bar), .ZN(n701bar) );
  OR2_X1 U263 ( .A1(n944), .A2(n872), .ZN(n699) );
  AND2_X1 U263bar ( .A1(n944bar), .A2(n872bar), .ZN(n699bar) );
  OR2_X1 U264 ( .A1(n698), .A2(n697), .ZN(n872) );
  AND2_X1 U264bar ( .A1(n698bar), .A2(n697bar), .ZN(n872bar) );
  OR2_X1 U265 ( .A1(n696), .A2(n695), .ZN(n697) );
  AND2_X1 U265bar ( .A1(n696bar), .A2(n695bar), .ZN(n697bar) );
  OR2_X1 U266 ( .A1(n694), .A2(n693), .ZN(n695) );
  AND2_X1 U266bar ( .A1(n694bar), .A2(n693bar), .ZN(n695bar) );
  OR2_X1 U267 ( .A1(in[121]), .A2(in[102]), .ZN(n693) );
  AND2_X1 U267bar ( .A1(inbar[121]), .A2(inbar[102]), .ZN(n693bar) );
  OR2_X1 U268 ( .A1(in[162]), .A2(in[161]), .ZN(n694) );
  AND2_X1 U268bar ( .A1(inbar[162]), .A2(inbar[161]), .ZN(n694bar) );
  OR2_X1 U269 ( .A1(n692), .A2(n691), .ZN(n696) );
  AND2_X1 U269bar ( .A1(n692bar), .A2(n691bar), .ZN(n696bar) );
  OR2_X1 U270 ( .A1(in[192]), .A2(in[178]), .ZN(n691) );
  AND2_X1 U270bar ( .A1(inbar[192]), .A2(inbar[178]), .ZN(n691bar) );
  OR2_X1 U271 ( .A1(in[244]), .A2(in[209]), .ZN(n692) );
  AND2_X1 U271bar ( .A1(inbar[244]), .A2(inbar[209]), .ZN(n692bar) );
  OR2_X1 U272 ( .A1(n690), .A2(n689), .ZN(n698) );
  AND2_X1 U272bar ( .A1(n690bar), .A2(n689bar), .ZN(n698bar) );
  OR2_X1 U273 ( .A1(n688), .A2(n687), .ZN(n689) );
  AND2_X1 U273bar ( .A1(n688bar), .A2(n687bar), .ZN(n689bar) );
  OR2_X1 U274 ( .A1(in[90]), .A2(in[254]), .ZN(n687) );
  AND2_X1 U274bar ( .A1(inbar[90]), .A2(inbar[254]), .ZN(n687bar) );
  OR2_X1 U275 ( .A1(in_36), .A2(in_32), .ZN(n688) );
  AND2_X1 U275bar ( .A1(in_36bar), .A2(in_32bar), .ZN(n688bar) );
  OR2_X1 U276 ( .A1(n686), .A2(n685), .ZN(n690) );
  AND2_X1 U276bar ( .A1(n686bar), .A2(n685bar), .ZN(n690bar) );
  OR2_X1 U277 ( .A1(in_62), .A2(in_37), .ZN(n685) );
  AND2_X1 U277bar ( .A1(in_62bar), .A2(in_37bar), .ZN(n685bar) );
  OR2_X1 U278 ( .A1(in_75), .A2(in_73), .ZN(n686) );
  AND2_X1 U278bar ( .A1(in_75bar), .A2(in_73bar), .ZN(n686bar) );
  OR2_X1 U279 ( .A1(n684), .A2(n683), .ZN(n944) );
  AND2_X1 U279bar ( .A1(n684bar), .A2(n683bar), .ZN(n944bar) );
  OR2_X1 U280 ( .A1(n682), .A2(n681), .ZN(n683) );
  AND2_X1 U280bar ( .A1(n682bar), .A2(n681bar), .ZN(n683bar) );
  OR2_X1 U281 ( .A1(n680), .A2(n679), .ZN(n681) );
  AND2_X1 U281bar ( .A1(n680bar), .A2(n679bar), .ZN(n681bar) );
  OR2_X1 U282 ( .A1(in[171]), .A2(in[153]), .ZN(n679) );
  AND2_X1 U282bar ( .A1(inbar[171]), .A2(inbar[153]), .ZN(n679bar) );
  OR2_X1 U283 ( .A1(in[187]), .A2(in[176]), .ZN(n680) );
  AND2_X1 U283bar ( .A1(inbar[187]), .A2(inbar[176]), .ZN(n680bar) );
  OR2_X1 U284 ( .A1(n678), .A2(n677), .ZN(n682) );
  AND2_X1 U284bar ( .A1(n678bar), .A2(n677bar), .ZN(n682bar) );
  OR2_X1 U285 ( .A1(in[245]), .A2(in[211]), .ZN(n677) );
  AND2_X1 U285bar ( .A1(inbar[245]), .A2(inbar[211]), .ZN(n677bar) );
  OR2_X1 U286 ( .A1(in[97]), .A2(in[88]), .ZN(n678) );
  AND2_X1 U286bar ( .A1(inbar[97]), .A2(inbar[88]), .ZN(n678bar) );
  OR2_X1 U287 ( .A1(n676), .A2(n675), .ZN(n684) );
  AND2_X1 U287bar ( .A1(n676bar), .A2(n675bar), .ZN(n684bar) );
  OR2_X1 U288 ( .A1(n674), .A2(n673), .ZN(n675) );
  AND2_X1 U288bar ( .A1(n674bar), .A2(n673bar), .ZN(n675bar) );
  OR2_X1 U289 ( .A1(in_10), .A2(in_0), .ZN(n673) );
  AND2_X1 U289bar ( .A1(in_10bar), .A2(in_0bar), .ZN(n673bar) );
  OR2_X1 U290 ( .A1(in_59), .A2(in_5), .ZN(n674) );
  AND2_X1 U290bar ( .A1(in_59bar), .A2(in_5bar), .ZN(n674bar) );
  OR2_X1 U291 ( .A1(n672), .A2(n671), .ZN(n676) );
  AND2_X1 U291bar ( .A1(n672bar), .A2(n671bar), .ZN(n676bar) );
  OR2_X1 U292 ( .A1(in_60), .A2(in_6), .ZN(n671) );
  AND2_X1 U292bar ( .A1(in_60bar), .A2(in_6bar), .ZN(n671bar) );
  OR2_X1 U293 ( .A1(in_77), .A2(in_69), .ZN(n672) );
  AND2_X1 U293bar ( .A1(in_77bar), .A2(in_69bar), .ZN(n672bar) );
  OR2_X1 U294 ( .A1(in[113]), .A2(n864), .ZN(n700) );
  AND2_X1 U294bar ( .A1(inbar[113]), .A2(n864bar), .ZN(n700bar) );
  OR2_X1 U295 ( .A1(n670), .A2(n669), .ZN(n864) );
  AND2_X1 U295bar ( .A1(n670bar), .A2(n669bar), .ZN(n864bar) );
  OR2_X1 U296 ( .A1(n668), .A2(n667), .ZN(n669) );
  AND2_X1 U296bar ( .A1(n668bar), .A2(n667bar), .ZN(n669bar) );
  OR2_X1 U297 ( .A1(n666), .A2(n665), .ZN(n667) );
  AND2_X1 U297bar ( .A1(n666bar), .A2(n665bar), .ZN(n667bar) );
  OR2_X1 U298 ( .A1(in[125]), .A2(in[107]), .ZN(n665) );
  AND2_X1 U298bar ( .A1(inbar[125]), .A2(inbar[107]), .ZN(n665bar) );
  OR2_X1 U299 ( .A1(in[138]), .A2(in[126]), .ZN(n666) );
  AND2_X1 U299bar ( .A1(inbar[138]), .A2(inbar[126]), .ZN(n666bar) );
  OR2_X1 U300 ( .A1(n664), .A2(n663), .ZN(n668) );
  AND2_X1 U300bar ( .A1(n664bar), .A2(n663bar), .ZN(n668bar) );
  OR2_X1 U301 ( .A1(in[189]), .A2(in[143]), .ZN(n663) );
  AND2_X1 U301bar ( .A1(inbar[189]), .A2(inbar[143]), .ZN(n663bar) );
  OR2_X1 U302 ( .A1(in[99]), .A2(in[214]), .ZN(n664) );
  AND2_X1 U302bar ( .A1(inbar[99]), .A2(inbar[214]), .ZN(n664bar) );
  OR2_X1 U303 ( .A1(n662), .A2(n661), .ZN(n670) );
  AND2_X1 U303bar ( .A1(n662bar), .A2(n661bar), .ZN(n670bar) );
  OR2_X1 U304 ( .A1(n660), .A2(n659), .ZN(n661) );
  AND2_X1 U304bar ( .A1(n660bar), .A2(n659bar), .ZN(n661bar) );
  OR2_X1 U305 ( .A1(in_15), .A2(in_12), .ZN(n659) );
  AND2_X1 U305bar ( .A1(in_15bar), .A2(in_12bar), .ZN(n659bar) );
  OR2_X1 U306 ( .A1(in_20), .A2(in_2), .ZN(n660) );
  AND2_X1 U306bar ( .A1(in_20bar), .A2(in_2bar), .ZN(n660bar) );
  OR2_X1 U307 ( .A1(n658), .A2(n657), .ZN(n662) );
  AND2_X1 U307bar ( .A1(n658bar), .A2(n657bar), .ZN(n662bar) );
  OR2_X1 U308 ( .A1(in_30), .A2(in_3), .ZN(n657) );
  AND2_X1 U308bar ( .A1(in_30bar), .A2(in_3bar), .ZN(n657bar) );
  OR2_X1 U309 ( .A1(in_4), .A2(in_38), .ZN(n658) );
  AND2_X1 U309bar ( .A1(in_4bar), .A2(in_38bar), .ZN(n658bar) );
  OR2_X1 U310 ( .A1(n656), .A2(n655), .ZN(n702) );
  AND2_X1 U310bar ( .A1(n656bar), .A2(n655bar), .ZN(n702bar) );
  OR2_X1 U311 ( .A1(in[148]), .A2(in[137]), .ZN(n655) );
  AND2_X1 U311bar ( .A1(inbar[148]), .A2(inbar[137]), .ZN(n655bar) );
  OR2_X1 U312 ( .A1(in[149]), .A2(n654), .ZN(n656) );
  AND2_X1 U312bar ( .A1(inbar[149]), .A2(n654bar), .ZN(n656bar) );
  OR2_X1 U313 ( .A1(in[195]), .A2(in[190]), .ZN(n654) );
  AND2_X1 U313bar ( .A1(inbar[195]), .A2(inbar[190]), .ZN(n654bar) );
  OR2_X1 U314 ( .A1(n653), .A2(n652), .ZN(n704) );
  AND2_X1 U314bar ( .A1(n653bar), .A2(n652bar), .ZN(n704bar) );
  OR2_X1 U315 ( .A1(n651), .A2(n650), .ZN(n652) );
  AND2_X1 U315bar ( .A1(n651bar), .A2(n650bar), .ZN(n652bar) );
  OR2_X1 U316 ( .A1(in[98]), .A2(in[197]), .ZN(n650) );
  AND2_X1 U316bar ( .A1(inbar[98]), .A2(inbar[197]), .ZN(n650bar) );
  OR2_X1 U317 ( .A1(in_11), .A2(n649), .ZN(n651) );
  AND2_X1 U317bar ( .A1(in_11bar), .A2(n649bar), .ZN(n651bar) );
  OR2_X1 U318 ( .A1(in_26), .A2(in_14), .ZN(n649) );
  AND2_X1 U318bar ( .A1(in_26bar), .A2(in_14bar), .ZN(n649bar) );
  OR2_X1 U319 ( .A1(n648), .A2(n647), .ZN(n653) );
  AND2_X1 U319bar ( .A1(n648bar), .A2(n647bar), .ZN(n653bar) );
  OR2_X1 U320 ( .A1(in_35), .A2(in_27), .ZN(n647) );
  AND2_X1 U320bar ( .A1(in_35bar), .A2(in_27bar), .ZN(n647bar) );
  OR2_X1 U321 ( .A1(in_50), .A2(n646), .ZN(n648) );
  AND2_X1 U321bar ( .A1(in_50bar), .A2(n646bar), .ZN(n648bar) );
  OR2_X1 U322 ( .A1(in_78), .A2(in_61), .ZN(n646) );
  AND2_X1 U322bar ( .A1(in_78bar), .A2(in_61bar), .ZN(n646bar) );
  OR2_X1 U323 ( .A1(n942), .A2(n645), .ZN(n720) );
  AND2_X1 U323bar ( .A1(n942bar), .A2(n645bar), .ZN(n720bar) );
  OR2_X1 U324 ( .A1(in[106]), .A2(n863), .ZN(n645) );
  AND2_X1 U324bar ( .A1(inbar[106]), .A2(n863bar), .ZN(n645bar) );
  OR2_X1 U325 ( .A1(n644), .A2(n643), .ZN(n863) );
  AND2_X1 U325bar ( .A1(n644bar), .A2(n643bar), .ZN(n863bar) );
  OR2_X1 U326 ( .A1(n642), .A2(n641), .ZN(n643) );
  AND2_X1 U326bar ( .A1(n642bar), .A2(n641bar), .ZN(n643bar) );
  OR2_X1 U327 ( .A1(n640), .A2(n639), .ZN(n641) );
  AND2_X1 U327bar ( .A1(n640bar), .A2(n639bar), .ZN(n641bar) );
  OR2_X1 U328 ( .A1(in[127]), .A2(in[122]), .ZN(n639) );
  AND2_X1 U328bar ( .A1(inbar[127]), .A2(inbar[122]), .ZN(n639bar) );
  OR2_X1 U329 ( .A1(in[156]), .A2(in[132]), .ZN(n640) );
  AND2_X1 U329bar ( .A1(inbar[156]), .A2(inbar[132]), .ZN(n640bar) );
  OR2_X1 U330 ( .A1(n638), .A2(n637), .ZN(n642) );
  AND2_X1 U330bar ( .A1(n638bar), .A2(n637bar), .ZN(n642bar) );
  OR2_X1 U331 ( .A1(in[159]), .A2(in[157]), .ZN(n637) );
  AND2_X1 U331bar ( .A1(inbar[159]), .A2(inbar[157]), .ZN(n637bar) );
  OR2_X1 U332 ( .A1(in[185]), .A2(in[169]), .ZN(n638) );
  AND2_X1 U332bar ( .A1(inbar[185]), .A2(inbar[169]), .ZN(n638bar) );
  OR2_X1 U333 ( .A1(n636), .A2(n635), .ZN(n644) );
  AND2_X1 U333bar ( .A1(n636bar), .A2(n635bar), .ZN(n644bar) );
  OR2_X1 U334 ( .A1(n634), .A2(n633), .ZN(n635) );
  AND2_X1 U334bar ( .A1(n634bar), .A2(n633bar), .ZN(n635bar) );
  OR2_X1 U335 ( .A1(in[239]), .A2(in[218]), .ZN(n633) );
  AND2_X1 U335bar ( .A1(inbar[239]), .A2(inbar[218]), .ZN(n633bar) );
  OR2_X1 U336 ( .A1(in_13), .A2(in[87]), .ZN(n634) );
  AND2_X1 U336bar ( .A1(in_13bar), .A2(inbar[87]), .ZN(n634bar) );
  OR2_X1 U337 ( .A1(n632), .A2(n631), .ZN(n636) );
  AND2_X1 U337bar ( .A1(n632bar), .A2(n631bar), .ZN(n636bar) );
  OR2_X1 U338 ( .A1(in_72), .A2(in_70), .ZN(n631) );
  AND2_X1 U338bar ( .A1(in_72bar), .A2(in_70bar), .ZN(n631bar) );
  OR2_X1 U339 ( .A1(in_80), .A2(in_74), .ZN(n632) );
  AND2_X1 U339bar ( .A1(in_80bar), .A2(in_74bar), .ZN(n632bar) );
  OR2_X1 U340 ( .A1(n630), .A2(n629), .ZN(n942) );
  AND2_X1 U340bar ( .A1(n630bar), .A2(n629bar), .ZN(n942bar) );
  OR2_X1 U341 ( .A1(n628), .A2(n627), .ZN(n629) );
  AND2_X1 U341bar ( .A1(n628bar), .A2(n627bar), .ZN(n629bar) );
  OR2_X1 U342 ( .A1(n626), .A2(n625), .ZN(n627) );
  AND2_X1 U342bar ( .A1(n626bar), .A2(n625bar), .ZN(n627bar) );
  OR2_X1 U343 ( .A1(in[146]), .A2(in[100]), .ZN(n625) );
  AND2_X1 U343bar ( .A1(inbar[146]), .A2(inbar[100]), .ZN(n625bar) );
  OR2_X1 U344 ( .A1(in[168]), .A2(in[152]), .ZN(n626) );
  AND2_X1 U344bar ( .A1(inbar[168]), .A2(inbar[152]), .ZN(n626bar) );
  OR2_X1 U345 ( .A1(n624), .A2(n623), .ZN(n628) );
  AND2_X1 U345bar ( .A1(n624bar), .A2(n623bar), .ZN(n628bar) );
  OR2_X1 U346 ( .A1(in[199]), .A2(in[182]), .ZN(n623) );
  AND2_X1 U346bar ( .A1(inbar[199]), .A2(inbar[182]), .ZN(n623bar) );
  OR2_X1 U347 ( .A1(in[236]), .A2(in[204]), .ZN(n624) );
  AND2_X1 U347bar ( .A1(inbar[236]), .A2(inbar[204]), .ZN(n624bar) );
  OR2_X1 U348 ( .A1(n622), .A2(n621), .ZN(n630) );
  AND2_X1 U348bar ( .A1(n622bar), .A2(n621bar), .ZN(n630bar) );
  OR2_X1 U349 ( .A1(n620), .A2(n619), .ZN(n621) );
  AND2_X1 U349bar ( .A1(n620bar), .A2(n619bar), .ZN(n621bar) );
  OR2_X1 U350 ( .A1(in[89]), .A2(in[246]), .ZN(n619) );
  AND2_X1 U350bar ( .A1(inbar[89]), .A2(inbar[246]), .ZN(n619bar) );
  OR2_X1 U351 ( .A1(in[95]), .A2(in[92]), .ZN(n620) );
  AND2_X1 U351bar ( .A1(inbar[95]), .A2(inbar[92]), .ZN(n620bar) );
  OR2_X1 U352 ( .A1(n618), .A2(n617), .ZN(n622) );
  AND2_X1 U352bar ( .A1(n618bar), .A2(n617bar), .ZN(n622bar) );
  OR2_X1 U353 ( .A1(in_22), .A2(in_16), .ZN(n617) );
  AND2_X1 U353bar ( .A1(in_22bar), .A2(in_16bar), .ZN(n617bar) );
  OR2_X1 U354 ( .A1(in_51), .A2(in_49), .ZN(n618) );
  AND2_X1 U354bar ( .A1(in_51bar), .A2(in_49bar), .ZN(n618bar) );
  OR2_X1 U355 ( .A1(n616), .A2(n615), .ZN(n722) );
  AND2_X1 U355bar ( .A1(n616bar), .A2(n615bar), .ZN(n722bar) );
  OR2_X1 U356 ( .A1(in[158]), .A2(in[115]), .ZN(n615) );
  AND2_X1 U356bar ( .A1(inbar[158]), .A2(inbar[115]), .ZN(n615bar) );
  OR2_X1 U357 ( .A1(in[163]), .A2(n614), .ZN(n616) );
  AND2_X1 U357bar ( .A1(inbar[163]), .A2(n614bar), .ZN(n616bar) );
  OR2_X1 U358 ( .A1(in[206]), .A2(in[165]), .ZN(n614) );
  AND2_X1 U358bar ( .A1(inbar[206]), .A2(inbar[165]), .ZN(n614bar) );
  OR2_X1 U359 ( .A1(n613), .A2(n612), .ZN(n724) );
  AND2_X1 U359bar ( .A1(n613bar), .A2(n612bar), .ZN(n724bar) );
  OR2_X1 U360 ( .A1(n611), .A2(n610), .ZN(n612) );
  AND2_X1 U360bar ( .A1(n611bar), .A2(n610bar), .ZN(n612bar) );
  OR2_X1 U361 ( .A1(in[213]), .A2(in[207]), .ZN(n610) );
  AND2_X1 U361bar ( .A1(inbar[213]), .A2(inbar[207]), .ZN(n610bar) );
  OR2_X1 U362 ( .A1(in[215]), .A2(n609), .ZN(n611) );
  AND2_X1 U362bar ( .A1(inbar[215]), .A2(n609bar), .ZN(n611bar) );
  OR2_X1 U363 ( .A1(in[230]), .A2(in[220]), .ZN(n609) );
  AND2_X1 U363bar ( .A1(inbar[230]), .A2(inbar[220]), .ZN(n609bar) );
  OR2_X1 U364 ( .A1(n608), .A2(n607), .ZN(n613) );
  AND2_X1 U364bar ( .A1(n608bar), .A2(n607bar), .ZN(n613bar) );
  OR2_X1 U365 ( .A1(in[251]), .A2(in[234]), .ZN(n607) );
  AND2_X1 U365bar ( .A1(inbar[251]), .A2(inbar[234]), .ZN(n607bar) );
  OR2_X1 U366 ( .A1(in_17), .A2(n606), .ZN(n608) );
  AND2_X1 U366bar ( .A1(in_17bar), .A2(n606bar), .ZN(n608bar) );
  OR2_X1 U367 ( .A1(in_65), .A2(in_56), .ZN(n606) );
  AND2_X1 U367bar ( .A1(in_65bar), .A2(in_56bar), .ZN(n606bar) );
  OR2_X1 U368 ( .A1(n605), .A2(n604), .ZN(out[0]) );
  AND2_X1 U368bar ( .A1(n605bar), .A2(n604bar), .ZN(outbar[0]) );
  OR2_X1 U369 ( .A1(n603), .A2(n602), .ZN(n604) );
  AND2_X1 U369bar ( .A1(n603bar), .A2(n602bar), .ZN(n604bar) );
  OR2_X1 U370 ( .A1(n601), .A2(n600), .ZN(n602) );
  AND2_X1 U370bar ( .A1(n601bar), .A2(n600bar), .ZN(n602bar) );
  OR2_X1 U371 ( .A1(n820), .A2(n785), .ZN(n600) );
  AND2_X1 U371bar ( .A1(n820bar), .A2(n785bar), .ZN(n600bar) );
  OR2_X1 U372 ( .A1(n599), .A2(n598), .ZN(n785) );
  AND2_X1 U372bar ( .A1(n599bar), .A2(n598bar), .ZN(n785bar) );
  OR2_X1 U373 ( .A1(n597), .A2(n596), .ZN(n598) );
  AND2_X1 U373bar ( .A1(n597bar), .A2(n596bar), .ZN(n598bar) );
  OR2_X1 U374 ( .A1(n595), .A2(n594), .ZN(n596) );
  AND2_X1 U374bar ( .A1(n595bar), .A2(n594bar), .ZN(n596bar) );
  OR2_X1 U375 ( .A1(in[135]), .A2(in[104]), .ZN(n594) );
  AND2_X1 U375bar ( .A1(inbar[135]), .A2(inbar[104]), .ZN(n594bar) );
  OR2_X1 U376 ( .A1(in[188]), .A2(in[178]), .ZN(n595) );
  AND2_X1 U376bar ( .A1(inbar[188]), .A2(inbar[178]), .ZN(n595bar) );
  OR2_X1 U377 ( .A1(n593), .A2(n592), .ZN(n597) );
  AND2_X1 U377bar ( .A1(n593bar), .A2(n592bar), .ZN(n597bar) );
  OR2_X1 U378 ( .A1(in[217]), .A2(in[194]), .ZN(n592) );
  AND2_X1 U378bar ( .A1(inbar[217]), .A2(inbar[194]), .ZN(n592bar) );
  OR2_X1 U379 ( .A1(in[237]), .A2(in[218]), .ZN(n593) );
  AND2_X1 U379bar ( .A1(inbar[237]), .A2(inbar[218]), .ZN(n593bar) );
  OR2_X1 U380 ( .A1(n591), .A2(n590), .ZN(n599) );
  AND2_X1 U380bar ( .A1(n591bar), .A2(n590bar), .ZN(n599bar) );
  OR2_X1 U381 ( .A1(n589), .A2(n588), .ZN(n590) );
  AND2_X1 U381bar ( .A1(n589bar), .A2(n588bar), .ZN(n590bar) );
  OR2_X1 U382 ( .A1(in_2), .A2(in_10), .ZN(n588) );
  AND2_X1 U382bar ( .A1(in_2bar), .A2(in_10bar), .ZN(n588bar) );
  OR2_X1 U383 ( .A1(in_47), .A2(in_22), .ZN(n589) );
  AND2_X1 U383bar ( .A1(in_47bar), .A2(in_22bar), .ZN(n589bar) );
  OR2_X1 U384 ( .A1(n587), .A2(n586), .ZN(n591) );
  AND2_X1 U384bar ( .A1(n587bar), .A2(n586bar), .ZN(n591bar) );
  OR2_X1 U385 ( .A1(in_56), .A2(in_54), .ZN(n586) );
  AND2_X1 U385bar ( .A1(in_56bar), .A2(in_54bar), .ZN(n586bar) );
  OR2_X1 U386 ( .A1(in_63), .A2(in_61), .ZN(n587) );
  AND2_X1 U386bar ( .A1(in_63bar), .A2(in_61bar), .ZN(n587bar) );
  OR2_X1 U387 ( .A1(n585), .A2(n584), .ZN(n820) );
  AND2_X1 U387bar ( .A1(n585bar), .A2(n584bar), .ZN(n820bar) );
  OR2_X1 U388 ( .A1(n583), .A2(n582), .ZN(n584) );
  AND2_X1 U388bar ( .A1(n583bar), .A2(n582bar), .ZN(n584bar) );
  OR2_X1 U389 ( .A1(n581), .A2(n580), .ZN(n582) );
  AND2_X1 U389bar ( .A1(n581bar), .A2(n580bar), .ZN(n582bar) );
  OR2_X1 U390 ( .A1(in[158]), .A2(in[142]), .ZN(n580) );
  AND2_X1 U390bar ( .A1(inbar[158]), .A2(inbar[142]), .ZN(n580bar) );
  OR2_X1 U391 ( .A1(in[175]), .A2(in[164]), .ZN(n581) );
  AND2_X1 U391bar ( .A1(inbar[175]), .A2(inbar[164]), .ZN(n581bar) );
  OR2_X1 U392 ( .A1(n579), .A2(n578), .ZN(n583) );
  AND2_X1 U392bar ( .A1(n579bar), .A2(n578bar), .ZN(n583bar) );
  OR2_X1 U393 ( .A1(in[228]), .A2(in[204]), .ZN(n578) );
  AND2_X1 U393bar ( .A1(inbar[228]), .A2(inbar[204]), .ZN(n578bar) );
  OR2_X1 U394 ( .A1(in[91]), .A2(in[87]), .ZN(n579) );
  AND2_X1 U394bar ( .A1(inbar[91]), .A2(inbar[87]), .ZN(n579bar) );
  OR2_X1 U395 ( .A1(n577), .A2(n576), .ZN(n585) );
  AND2_X1 U395bar ( .A1(n577bar), .A2(n576bar), .ZN(n585bar) );
  OR2_X1 U396 ( .A1(n575), .A2(n574), .ZN(n576) );
  AND2_X1 U396bar ( .A1(n575bar), .A2(n574bar), .ZN(n576bar) );
  OR2_X1 U397 ( .A1(in_21), .A2(in_11), .ZN(n574) );
  AND2_X1 U397bar ( .A1(in_21bar), .A2(in_11bar), .ZN(n574bar) );
  OR2_X1 U398 ( .A1(in_5), .A2(in_3), .ZN(n575) );
  AND2_X1 U398bar ( .A1(in_5bar), .A2(in_3bar), .ZN(n575bar) );
  OR2_X1 U399 ( .A1(n573), .A2(n572), .ZN(n577) );
  AND2_X1 U399bar ( .A1(n573bar), .A2(n572bar), .ZN(n577bar) );
  OR2_X1 U400 ( .A1(in_68), .A2(in_64), .ZN(n572) );
  AND2_X1 U400bar ( .A1(in_68bar), .A2(in_64bar), .ZN(n572bar) );
  OR2_X1 U401 ( .A1(in_76), .A2(in_73), .ZN(n573) );
  AND2_X1 U401bar ( .A1(in_76bar), .A2(in_73bar), .ZN(n573bar) );
  OR2_X1 U402 ( .A1(n778), .A2(n571), .ZN(n601) );
  AND2_X1 U402bar ( .A1(n778bar), .A2(n571bar), .ZN(n601bar) );
  OR2_X1 U403 ( .A1(in[100]), .A2(n965), .ZN(n571) );
  AND2_X1 U403bar ( .A1(inbar[100]), .A2(n965bar), .ZN(n571bar) );
  OR2_X1 U404 ( .A1(n570), .A2(n569), .ZN(n965) );
  AND2_X1 U404bar ( .A1(n570bar), .A2(n569bar), .ZN(n965bar) );
  OR2_X1 U405 ( .A1(n568), .A2(n567), .ZN(n569) );
  AND2_X1 U405bar ( .A1(n568bar), .A2(n567bar), .ZN(n569bar) );
  OR2_X1 U406 ( .A1(n566), .A2(n565), .ZN(n567) );
  AND2_X1 U406bar ( .A1(n566bar), .A2(n565bar), .ZN(n567bar) );
  OR2_X1 U407 ( .A1(n817), .A2(n750), .ZN(n565) );
  AND2_X1 U407bar ( .A1(n817bar), .A2(n750bar), .ZN(n565bar) );
  OR2_X1 U408 ( .A1(n564), .A2(n563), .ZN(n750) );
  AND2_X1 U408bar ( .A1(n564bar), .A2(n563bar), .ZN(n750bar) );
  OR2_X1 U409 ( .A1(n562), .A2(n561), .ZN(n563) );
  AND2_X1 U409bar ( .A1(n562bar), .A2(n561bar), .ZN(n563bar) );
  OR2_X1 U410 ( .A1(n560), .A2(n559), .ZN(n561) );
  AND2_X1 U410bar ( .A1(n560bar), .A2(n559bar), .ZN(n561bar) );
  OR2_X1 U411 ( .A1(in[119]), .A2(in[103]), .ZN(n559) );
  AND2_X1 U411bar ( .A1(inbar[119]), .A2(inbar[103]), .ZN(n559bar) );
  OR2_X1 U412 ( .A1(in[137]), .A2(in[133]), .ZN(n560) );
  AND2_X1 U412bar ( .A1(inbar[137]), .A2(inbar[133]), .ZN(n560bar) );
  OR2_X1 U413 ( .A1(n558), .A2(n557), .ZN(n562) );
  AND2_X1 U413bar ( .A1(n558bar), .A2(n557bar), .ZN(n562bar) );
  OR2_X1 U414 ( .A1(in[176]), .A2(in[173]), .ZN(n557) );
  AND2_X1 U414bar ( .A1(inbar[176]), .A2(inbar[173]), .ZN(n557bar) );
  OR2_X1 U415 ( .A1(in[210]), .A2(in[181]), .ZN(n558) );
  AND2_X1 U415bar ( .A1(inbar[210]), .A2(inbar[181]), .ZN(n558bar) );
  OR2_X1 U416 ( .A1(n556), .A2(n555), .ZN(n564) );
  AND2_X1 U416bar ( .A1(n556bar), .A2(n555bar), .ZN(n564bar) );
  OR2_X1 U417 ( .A1(n554), .A2(n553), .ZN(n555) );
  AND2_X1 U417bar ( .A1(n554bar), .A2(n553bar), .ZN(n555bar) );
  OR2_X1 U418 ( .A1(in_13), .A2(in[234]), .ZN(n553) );
  AND2_X1 U418bar ( .A1(in_13bar), .A2(inbar[234]), .ZN(n553bar) );
  OR2_X1 U419 ( .A1(in_38), .A2(in_32), .ZN(n554) );
  AND2_X1 U419bar ( .A1(in_38bar), .A2(in_32bar), .ZN(n554bar) );
  OR2_X1 U420 ( .A1(n552), .A2(n551), .ZN(n556) );
  AND2_X1 U420bar ( .A1(n552bar), .A2(n551bar), .ZN(n556bar) );
  OR2_X1 U421 ( .A1(in_42), .A2(in_41), .ZN(n551) );
  AND2_X1 U421bar ( .A1(in_42bar), .A2(in_41bar), .ZN(n551bar) );
  OR2_X1 U422 ( .A1(in_7), .A2(in_49), .ZN(n552) );
  AND2_X1 U422bar ( .A1(in_7bar), .A2(in_49bar), .ZN(n552bar) );
  OR2_X1 U423 ( .A1(n550), .A2(n549), .ZN(n817) );
  AND2_X1 U423bar ( .A1(n550bar), .A2(n549bar), .ZN(n817bar) );
  OR2_X1 U424 ( .A1(n548), .A2(n547), .ZN(n549) );
  AND2_X1 U424bar ( .A1(n548bar), .A2(n547bar), .ZN(n549bar) );
  OR2_X1 U425 ( .A1(n546), .A2(n545), .ZN(n547) );
  AND2_X1 U425bar ( .A1(n546bar), .A2(n545bar), .ZN(n547bar) );
  OR2_X1 U426 ( .A1(in[159]), .A2(in[105]), .ZN(n545) );
  AND2_X1 U426bar ( .A1(inbar[159]), .A2(inbar[105]), .ZN(n545bar) );
  OR2_X1 U427 ( .A1(in[206]), .A2(in[183]), .ZN(n546) );
  AND2_X1 U427bar ( .A1(inbar[206]), .A2(inbar[183]), .ZN(n546bar) );
  OR2_X1 U428 ( .A1(n544), .A2(n543), .ZN(n548) );
  AND2_X1 U428bar ( .A1(n544bar), .A2(n543bar), .ZN(n548bar) );
  OR2_X1 U429 ( .A1(in[229]), .A2(in[219]), .ZN(n543) );
  AND2_X1 U429bar ( .A1(inbar[229]), .A2(inbar[219]), .ZN(n543bar) );
  OR2_X1 U430 ( .A1(in[235]), .A2(in[232]), .ZN(n544) );
  AND2_X1 U430bar ( .A1(inbar[235]), .A2(inbar[232]), .ZN(n544bar) );
  OR2_X1 U431 ( .A1(n542), .A2(n541), .ZN(n550) );
  AND2_X1 U431bar ( .A1(n542bar), .A2(n541bar), .ZN(n550bar) );
  OR2_X1 U432 ( .A1(n540), .A2(n539), .ZN(n541) );
  AND2_X1 U432bar ( .A1(n540bar), .A2(n539bar), .ZN(n541bar) );
  OR2_X1 U433 ( .A1(in[249]), .A2(in[242]), .ZN(n539) );
  AND2_X1 U433bar ( .A1(inbar[249]), .A2(inbar[242]), .ZN(n539bar) );
  OR2_X1 U434 ( .A1(in[89]), .A2(in[254]), .ZN(n540) );
  AND2_X1 U434bar ( .A1(inbar[89]), .A2(inbar[254]), .ZN(n540bar) );
  OR2_X1 U435 ( .A1(n538), .A2(n537), .ZN(n542) );
  AND2_X1 U435bar ( .A1(n538bar), .A2(n537bar), .ZN(n542bar) );
  OR2_X1 U436 ( .A1(in_14), .A2(in[99]), .ZN(n537) );
  AND2_X1 U436bar ( .A1(in_14bar), .A2(inbar[99]), .ZN(n537bar) );
  OR2_X1 U437 ( .A1(in_60), .A2(in_18), .ZN(n538) );
  AND2_X1 U437bar ( .A1(in_60bar), .A2(in_18bar), .ZN(n538bar) );
  OR2_X1 U438 ( .A1(in[113]), .A2(n763), .ZN(n566) );
  AND2_X1 U438bar ( .A1(inbar[113]), .A2(n763bar), .ZN(n566bar) );
  OR2_X1 U439 ( .A1(n536), .A2(n535), .ZN(n763) );
  AND2_X1 U439bar ( .A1(n536bar), .A2(n535bar), .ZN(n763bar) );
  OR2_X1 U440 ( .A1(n534), .A2(n533), .ZN(n535) );
  AND2_X1 U440bar ( .A1(n534bar), .A2(n533bar), .ZN(n535bar) );
  OR2_X1 U441 ( .A1(n532), .A2(n531), .ZN(n533) );
  AND2_X1 U441bar ( .A1(n532bar), .A2(n531bar), .ZN(n533bar) );
  OR2_X1 U442 ( .A1(in[115]), .A2(in[110]), .ZN(n531) );
  AND2_X1 U442bar ( .A1(inbar[115]), .A2(inbar[110]), .ZN(n531bar) );
  OR2_X1 U443 ( .A1(in[125]), .A2(in[117]), .ZN(n532) );
  AND2_X1 U443bar ( .A1(inbar[125]), .A2(inbar[117]), .ZN(n532bar) );
  OR2_X1 U444 ( .A1(n530), .A2(n529), .ZN(n534) );
  AND2_X1 U444bar ( .A1(n530bar), .A2(n529bar), .ZN(n534bar) );
  OR2_X1 U445 ( .A1(in[180]), .A2(in[128]), .ZN(n529) );
  AND2_X1 U445bar ( .A1(inbar[180]), .A2(inbar[128]), .ZN(n529bar) );
  OR2_X1 U446 ( .A1(in[205]), .A2(in[201]), .ZN(n530) );
  AND2_X1 U446bar ( .A1(inbar[205]), .A2(inbar[201]), .ZN(n530bar) );
  OR2_X1 U447 ( .A1(n528), .A2(n527), .ZN(n536) );
  AND2_X1 U447bar ( .A1(n528bar), .A2(n527bar), .ZN(n536bar) );
  OR2_X1 U448 ( .A1(n526), .A2(n525), .ZN(n527) );
  AND2_X1 U448bar ( .A1(n526bar), .A2(n525bar), .ZN(n527bar) );
  OR2_X1 U449 ( .A1(in[244]), .A2(in[239]), .ZN(n525) );
  AND2_X1 U449bar ( .A1(inbar[244]), .A2(inbar[239]), .ZN(n525bar) );
  OR2_X1 U450 ( .A1(in[95]), .A2(in[83]), .ZN(n526) );
  AND2_X1 U450bar ( .A1(inbar[95]), .A2(inbar[83]), .ZN(n526bar) );
  OR2_X1 U451 ( .A1(n524), .A2(n523), .ZN(n528) );
  AND2_X1 U451bar ( .A1(n524bar), .A2(n523bar), .ZN(n528bar) );
  OR2_X1 U452 ( .A1(in_24), .A2(in[97]), .ZN(n523) );
  AND2_X1 U452bar ( .A1(in_24bar), .A2(inbar[97]), .ZN(n523bar) );
  OR2_X1 U453 ( .A1(in_33), .A2(in_27), .ZN(n524) );
  AND2_X1 U453bar ( .A1(in_33bar), .A2(in_27bar), .ZN(n524bar) );
  OR2_X1 U454 ( .A1(n522), .A2(n521), .ZN(n568) );
  AND2_X1 U454bar ( .A1(n522bar), .A2(n521bar), .ZN(n568bar) );
  OR2_X1 U455 ( .A1(in[145]), .A2(in[126]), .ZN(n521) );
  AND2_X1 U455bar ( .A1(inbar[145]), .A2(inbar[126]), .ZN(n521bar) );
  OR2_X1 U456 ( .A1(in[169]), .A2(n520), .ZN(n522) );
  AND2_X1 U456bar ( .A1(inbar[169]), .A2(n520bar), .ZN(n522bar) );
  OR2_X1 U457 ( .A1(in[221]), .A2(in[172]), .ZN(n520) );
  AND2_X1 U457bar ( .A1(inbar[221]), .A2(inbar[172]), .ZN(n520bar) );
  OR2_X1 U458 ( .A1(n519), .A2(n518), .ZN(n570) );
  AND2_X1 U458bar ( .A1(n519bar), .A2(n518bar), .ZN(n570bar) );
  OR2_X1 U459 ( .A1(n517), .A2(n516), .ZN(n518) );
  AND2_X1 U459bar ( .A1(n517bar), .A2(n516bar), .ZN(n518bar) );
  OR2_X1 U460 ( .A1(in[241]), .A2(in[224]), .ZN(n516) );
  AND2_X1 U460bar ( .A1(inbar[241]), .A2(inbar[224]), .ZN(n516bar) );
  OR2_X1 U461 ( .A1(in[86]), .A2(n515), .ZN(n517) );
  AND2_X1 U461bar ( .A1(inbar[86]), .A2(n515bar), .ZN(n517bar) );
  OR2_X1 U462 ( .A1(in_43), .A2(in_34), .ZN(n515) );
  AND2_X1 U462bar ( .A1(in_43bar), .A2(in_34bar), .ZN(n515bar) );
  OR2_X1 U463 ( .A1(n514), .A2(n513), .ZN(n519) );
  AND2_X1 U463bar ( .A1(n514bar), .A2(n513bar), .ZN(n519bar) );
  OR2_X1 U464 ( .A1(in_65), .A2(in_51), .ZN(n513) );
  AND2_X1 U464bar ( .A1(in_65bar), .A2(in_51bar), .ZN(n513bar) );
  OR2_X1 U465 ( .A1(in_75), .A2(n512), .ZN(n514) );
  AND2_X1 U465bar ( .A1(in_75bar), .A2(n512bar), .ZN(n514bar) );
  OR2_X1 U466 ( .A1(in_81), .A2(in_77), .ZN(n512) );
  AND2_X1 U466bar ( .A1(in_81bar), .A2(in_77bar), .ZN(n512bar) );
  OR2_X1 U467 ( .A1(n511), .A2(n510), .ZN(n778) );
  AND2_X1 U467bar ( .A1(n511bar), .A2(n510bar), .ZN(n778bar) );
  OR2_X1 U468 ( .A1(n509), .A2(n508), .ZN(n510) );
  AND2_X1 U468bar ( .A1(n509bar), .A2(n508bar), .ZN(n510bar) );
  OR2_X1 U469 ( .A1(n507), .A2(n506), .ZN(n508) );
  AND2_X1 U469bar ( .A1(n507bar), .A2(n506bar), .ZN(n508bar) );
  OR2_X1 U470 ( .A1(in[107]), .A2(in[101]), .ZN(n506) );
  AND2_X1 U470bar ( .A1(inbar[107]), .A2(inbar[101]), .ZN(n506bar) );
  OR2_X1 U471 ( .A1(in[139]), .A2(in[132]), .ZN(n507) );
  AND2_X1 U471bar ( .A1(inbar[139]), .A2(inbar[132]), .ZN(n507bar) );
  OR2_X1 U472 ( .A1(n505), .A2(n504), .ZN(n509) );
  AND2_X1 U472bar ( .A1(n505bar), .A2(n504bar), .ZN(n509bar) );
  OR2_X1 U473 ( .A1(in[146]), .A2(in[141]), .ZN(n504) );
  AND2_X1 U473bar ( .A1(inbar[146]), .A2(inbar[141]), .ZN(n504bar) );
  OR2_X1 U474 ( .A1(in[203]), .A2(in[179]), .ZN(n505) );
  AND2_X1 U474bar ( .A1(inbar[203]), .A2(inbar[179]), .ZN(n505bar) );
  OR2_X1 U475 ( .A1(n503), .A2(n502), .ZN(n511) );
  AND2_X1 U475bar ( .A1(n503bar), .A2(n502bar), .ZN(n511bar) );
  OR2_X1 U476 ( .A1(n501), .A2(n500), .ZN(n502) );
  AND2_X1 U476bar ( .A1(n501bar), .A2(n500bar), .ZN(n502bar) );
  OR2_X1 U477 ( .A1(in[243]), .A2(in[222]), .ZN(n500) );
  AND2_X1 U477bar ( .A1(inbar[243]), .A2(inbar[222]), .ZN(n500bar) );
  OR2_X1 U478 ( .A1(in[251]), .A2(in[250]), .ZN(n501) );
  AND2_X1 U478bar ( .A1(inbar[251]), .A2(inbar[250]), .ZN(n501bar) );
  OR2_X1 U479 ( .A1(n499), .A2(n498), .ZN(n503) );
  AND2_X1 U479bar ( .A1(n499bar), .A2(n498bar), .ZN(n503bar) );
  OR2_X1 U480 ( .A1(in_37), .A2(in_19), .ZN(n498) );
  AND2_X1 U480bar ( .A1(in_37bar), .A2(in_19bar), .ZN(n498bar) );
  OR2_X1 U481 ( .A1(in_78), .A2(in_6), .ZN(n499) );
  AND2_X1 U481bar ( .A1(in_78bar), .A2(in_6bar), .ZN(n499bar) );
  OR2_X1 U482 ( .A1(n497), .A2(n496), .ZN(n603) );
  AND2_X1 U482bar ( .A1(n497bar), .A2(n496bar), .ZN(n603bar) );
  OR2_X1 U483 ( .A1(in[112]), .A2(in[102]), .ZN(n496) );
  AND2_X1 U483bar ( .A1(inbar[112]), .A2(inbar[102]), .ZN(n496bar) );
  OR2_X1 U484 ( .A1(in[123]), .A2(n495), .ZN(n497) );
  AND2_X1 U484bar ( .A1(inbar[123]), .A2(n495bar), .ZN(n497bar) );
  OR2_X1 U485 ( .A1(in[143]), .A2(in[130]), .ZN(n495) );
  AND2_X1 U485bar ( .A1(inbar[143]), .A2(inbar[130]), .ZN(n495bar) );
  OR2_X1 U486 ( .A1(n494), .A2(n493), .ZN(n605) );
  AND2_X1 U486bar ( .A1(n494bar), .A2(n493bar), .ZN(n605bar) );
  OR2_X1 U487 ( .A1(n492), .A2(n491), .ZN(n493) );
  AND2_X1 U487bar ( .A1(n492bar), .A2(n491bar), .ZN(n493bar) );
  OR2_X1 U488 ( .A1(in[216]), .A2(in[213]), .ZN(n491) );
  AND2_X1 U488bar ( .A1(inbar[216]), .A2(inbar[213]), .ZN(n491bar) );
  OR2_X1 U489 ( .A1(in[227]), .A2(n490), .ZN(n492) );
  AND2_X1 U489bar ( .A1(inbar[227]), .A2(n490bar), .ZN(n492bar) );
  OR2_X1 U490 ( .A1(in_0), .A2(in[248]), .ZN(n490) );
  AND2_X1 U490bar ( .A1(in_0bar), .A2(inbar[248]), .ZN(n490bar) );
  OR2_X1 U491 ( .A1(n489), .A2(n488), .ZN(n494) );
  AND2_X1 U491bar ( .A1(n489bar), .A2(n488bar), .ZN(n494bar) );
  OR2_X1 U492 ( .A1(in_46), .A2(in_44), .ZN(n488) );
  AND2_X1 U492bar ( .A1(in_46bar), .A2(in_44bar), .ZN(n488bar) );
  OR2_X1 U493 ( .A1(in_50), .A2(n487), .ZN(n489) );
  AND2_X1 U493bar ( .A1(in_50bar), .A2(n487bar), .ZN(n489bar) );
  OR2_X1 U494 ( .A1(in_9), .A2(in_80), .ZN(n487) );
  AND2_X1 U494bar ( .A1(in_9bar), .A2(in_80bar), .ZN(n487bar) );
endmodule

module sBox_14 ( in, inbar, out, outbar );

  input wire [7:0] in;
  input wire [7:0] inbar;
//input_done

  output wire [7:0] out;
  output wire [7:0] outbar;
//output_done

  wire [255:0] decodeOut;
  wire [255:0] decodeOutbar;
//wire_done

  decode_14 dec ( .in(in), .inbar(inbar), .out(decodeOut), .outbar(decodeOutbar) );
  encode_14 enc ( .in(decodeOut), .inbar(decodeOutbar), .out(out), .outbar(outbar) );
endmodule

module CD2_57 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD2_58 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD2_59 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD2_60 ( a, abar, b, bbar, y, ybar );

  input wire a;
  input wire b;
  input wire abar;
  input wire bbar;
//input_done

  output wire [3:0] y;
  output wire [3:0] ybar;
//output_done

  wire n1;
  wire n2;
  wire n1bar;
  wire n2bar;
//wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]) );
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]) );
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]) );
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]) );
endmodule

module CD4_29 ( a, abar, b, bbar, y, ybar );

  input wire [3:0] a;
  input wire [3:0] b;
  input wire [3:0] abar;
  input wire [3:0] bbar;
//input_done

  output wire [15:0] y;
  output wire [15:0] ybar;
//output_done

//wire_done

  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]) );
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]) );
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]) );
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]) );
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]) );
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]) );
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]) );
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]) );
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]) );
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]) );
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]) );
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]) );
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]) );
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]) );
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]) );
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]) );
endmodule

module CD4_30 ( a, abar, b, bbar, y, ybar );

  input wire [3:0] a;
  input wire [3:0] b;
  input wire [3:0] abar;
  input wire [3:0] bbar;
//input_done

  output wire [15:0] y;
  output wire [15:0] ybar;
//output_done

//wire_done

  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]) );
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]) );
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]) );
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]) );
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]) );
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]) );
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]) );
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]) );
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]) );
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]) );
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]) );
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]) );
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]) );
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]) );
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]) );
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]) );
endmodule

module CD16_15 ( a, abar, b, bbar, y, ybar );

  input wire [15:0] a;
  input wire [15:0] b;
  input wire [15:0] abar;
  input wire [15:0] bbar;
//input_done

  output wire [255:0] y;
  output wire [255:0] ybar;
//output_done

//wire_done

  AND2_X1 U1 ( .A1(b[9]), .A2(a[0]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[9]), .A2(abar[0]), .ZN(ybar[9]) );
  AND2_X1 U2 ( .A1(b[3]), .A2(a[6]), .ZN(y[99]) );
  OR2_X1 U2bar ( .A1(bbar[3]), .A2(abar[6]), .ZN(ybar[99]) );
  AND2_X1 U3 ( .A1(b[2]), .A2(a[6]), .ZN(y[98]) );
  OR2_X1 U3bar ( .A1(bbar[2]), .A2(abar[6]), .ZN(ybar[98]) );
  AND2_X1 U4 ( .A1(b[1]), .A2(a[6]), .ZN(y[97]) );
  OR2_X1 U4bar ( .A1(bbar[1]), .A2(abar[6]), .ZN(ybar[97]) );
  AND2_X1 U5 ( .A1(b[0]), .A2(a[6]), .ZN(y[96]) );
  OR2_X1 U5bar ( .A1(bbar[0]), .A2(abar[6]), .ZN(ybar[96]) );
  AND2_X1 U6 ( .A1(b[15]), .A2(a[5]), .ZN(y[95]) );
  OR2_X1 U6bar ( .A1(bbar[15]), .A2(abar[5]), .ZN(ybar[95]) );
  AND2_X1 U7 ( .A1(b[14]), .A2(a[5]), .ZN(y[94]) );
  OR2_X1 U7bar ( .A1(bbar[14]), .A2(abar[5]), .ZN(ybar[94]) );
  AND2_X1 U8 ( .A1(b[13]), .A2(a[5]), .ZN(y[93]) );
  OR2_X1 U8bar ( .A1(bbar[13]), .A2(abar[5]), .ZN(ybar[93]) );
  AND2_X1 U9 ( .A1(b[12]), .A2(a[5]), .ZN(y[92]) );
  OR2_X1 U9bar ( .A1(bbar[12]), .A2(abar[5]), .ZN(ybar[92]) );
  AND2_X1 U10 ( .A1(b[11]), .A2(a[5]), .ZN(y[91]) );
  OR2_X1 U10bar ( .A1(bbar[11]), .A2(abar[5]), .ZN(ybar[91]) );
  AND2_X1 U11 ( .A1(b[10]), .A2(a[5]), .ZN(y[90]) );
  OR2_X1 U11bar ( .A1(bbar[10]), .A2(abar[5]), .ZN(ybar[90]) );
  AND2_X1 U12 ( .A1(b[8]), .A2(a[0]), .ZN(y[8]) );
  OR2_X1 U12bar ( .A1(bbar[8]), .A2(abar[0]), .ZN(ybar[8]) );
  AND2_X1 U13 ( .A1(a[5]), .A2(b[9]), .ZN(y[89]) );
  OR2_X1 U13bar ( .A1(abar[5]), .A2(bbar[9]), .ZN(ybar[89]) );
  AND2_X1 U14 ( .A1(b[8]), .A2(a[5]), .ZN(y[88]) );
  OR2_X1 U14bar ( .A1(bbar[8]), .A2(abar[5]), .ZN(ybar[88]) );
  AND2_X1 U15 ( .A1(b[7]), .A2(a[5]), .ZN(y[87]) );
  OR2_X1 U15bar ( .A1(bbar[7]), .A2(abar[5]), .ZN(ybar[87]) );
  AND2_X1 U16 ( .A1(b[6]), .A2(a[5]), .ZN(y[86]) );
  OR2_X1 U16bar ( .A1(bbar[6]), .A2(abar[5]), .ZN(ybar[86]) );
  AND2_X1 U17 ( .A1(b[5]), .A2(a[5]), .ZN(y[85]) );
  OR2_X1 U17bar ( .A1(bbar[5]), .A2(abar[5]), .ZN(ybar[85]) );
  AND2_X1 U18 ( .A1(b[4]), .A2(a[5]), .ZN(y[84]) );
  OR2_X1 U18bar ( .A1(bbar[4]), .A2(abar[5]), .ZN(ybar[84]) );
  AND2_X1 U19 ( .A1(a[5]), .A2(b[3]), .ZN(y[83]) );
  OR2_X1 U19bar ( .A1(abar[5]), .A2(bbar[3]), .ZN(ybar[83]) );
  AND2_X1 U20 ( .A1(a[5]), .A2(b[2]), .ZN(y[82]) );
  OR2_X1 U20bar ( .A1(abar[5]), .A2(bbar[2]), .ZN(ybar[82]) );
  AND2_X1 U21 ( .A1(a[5]), .A2(b[1]), .ZN(y[81]) );
  OR2_X1 U21bar ( .A1(abar[5]), .A2(bbar[1]), .ZN(ybar[81]) );
  AND2_X1 U22 ( .A1(a[5]), .A2(b[0]), .ZN(y[80]) );
  OR2_X1 U22bar ( .A1(abar[5]), .A2(bbar[0]), .ZN(ybar[80]) );
  AND2_X1 U23 ( .A1(b[7]), .A2(a[0]), .ZN(y[7]) );
  OR2_X1 U23bar ( .A1(bbar[7]), .A2(abar[0]), .ZN(ybar[7]) );
  AND2_X1 U24 ( .A1(a[4]), .A2(b[15]), .ZN(y[79]) );
  OR2_X1 U24bar ( .A1(abar[4]), .A2(bbar[15]), .ZN(ybar[79]) );
  AND2_X1 U25 ( .A1(a[4]), .A2(b[14]), .ZN(y[78]) );
  OR2_X1 U25bar ( .A1(abar[4]), .A2(bbar[14]), .ZN(ybar[78]) );
  AND2_X1 U26 ( .A1(a[4]), .A2(b[13]), .ZN(y[77]) );
  OR2_X1 U26bar ( .A1(abar[4]), .A2(bbar[13]), .ZN(ybar[77]) );
  AND2_X1 U27 ( .A1(a[4]), .A2(b[12]), .ZN(y[76]) );
  OR2_X1 U27bar ( .A1(abar[4]), .A2(bbar[12]), .ZN(ybar[76]) );
  AND2_X1 U28 ( .A1(a[4]), .A2(b[11]), .ZN(y[75]) );
  OR2_X1 U28bar ( .A1(abar[4]), .A2(bbar[11]), .ZN(ybar[75]) );
  AND2_X1 U29 ( .A1(a[4]), .A2(b[10]), .ZN(y[74]) );
  OR2_X1 U29bar ( .A1(abar[4]), .A2(bbar[10]), .ZN(ybar[74]) );
  AND2_X1 U30 ( .A1(a[4]), .A2(b[9]), .ZN(y[73]) );
  OR2_X1 U30bar ( .A1(abar[4]), .A2(bbar[9]), .ZN(ybar[73]) );
  AND2_X1 U31 ( .A1(a[4]), .A2(b[8]), .ZN(y[72]) );
  OR2_X1 U31bar ( .A1(abar[4]), .A2(bbar[8]), .ZN(ybar[72]) );
  AND2_X1 U32 ( .A1(a[4]), .A2(b[7]), .ZN(y[71]) );
  OR2_X1 U32bar ( .A1(abar[4]), .A2(bbar[7]), .ZN(ybar[71]) );
  AND2_X1 U33 ( .A1(a[4]), .A2(b[6]), .ZN(y[70]) );
  OR2_X1 U33bar ( .A1(abar[4]), .A2(bbar[6]), .ZN(ybar[70]) );
  AND2_X1 U34 ( .A1(b[6]), .A2(a[0]), .ZN(y[6]) );
  OR2_X1 U34bar ( .A1(bbar[6]), .A2(abar[0]), .ZN(ybar[6]) );
  AND2_X1 U35 ( .A1(a[4]), .A2(b[5]), .ZN(y[69]) );
  OR2_X1 U35bar ( .A1(abar[4]), .A2(bbar[5]), .ZN(ybar[69]) );
  AND2_X1 U36 ( .A1(a[4]), .A2(b[4]), .ZN(y[68]) );
  OR2_X1 U36bar ( .A1(abar[4]), .A2(bbar[4]), .ZN(ybar[68]) );
  AND2_X1 U37 ( .A1(a[4]), .A2(b[3]), .ZN(y[67]) );
  OR2_X1 U37bar ( .A1(abar[4]), .A2(bbar[3]), .ZN(ybar[67]) );
  AND2_X1 U38 ( .A1(a[4]), .A2(b[2]), .ZN(y[66]) );
  OR2_X1 U38bar ( .A1(abar[4]), .A2(bbar[2]), .ZN(ybar[66]) );
  AND2_X1 U39 ( .A1(a[4]), .A2(b[1]), .ZN(y[65]) );
  OR2_X1 U39bar ( .A1(abar[4]), .A2(bbar[1]), .ZN(ybar[65]) );
  AND2_X1 U40 ( .A1(a[4]), .A2(b[0]), .ZN(y[64]) );
  OR2_X1 U40bar ( .A1(abar[4]), .A2(bbar[0]), .ZN(ybar[64]) );
  AND2_X1 U41 ( .A1(a[3]), .A2(b[15]), .ZN(y[63]) );
  OR2_X1 U41bar ( .A1(abar[3]), .A2(bbar[15]), .ZN(ybar[63]) );
  AND2_X1 U42 ( .A1(a[3]), .A2(b[14]), .ZN(y[62]) );
  OR2_X1 U42bar ( .A1(abar[3]), .A2(bbar[14]), .ZN(ybar[62]) );
  AND2_X1 U43 ( .A1(a[3]), .A2(b[13]), .ZN(y[61]) );
  OR2_X1 U43bar ( .A1(abar[3]), .A2(bbar[13]), .ZN(ybar[61]) );
  AND2_X1 U44 ( .A1(a[3]), .A2(b[12]), .ZN(y[60]) );
  OR2_X1 U44bar ( .A1(abar[3]), .A2(bbar[12]), .ZN(ybar[60]) );
  AND2_X1 U45 ( .A1(b[5]), .A2(a[0]), .ZN(y[5]) );
  OR2_X1 U45bar ( .A1(bbar[5]), .A2(abar[0]), .ZN(ybar[5]) );
  AND2_X1 U46 ( .A1(a[3]), .A2(b[11]), .ZN(y[59]) );
  OR2_X1 U46bar ( .A1(abar[3]), .A2(bbar[11]), .ZN(ybar[59]) );
  AND2_X1 U47 ( .A1(a[3]), .A2(b[10]), .ZN(y[58]) );
  OR2_X1 U47bar ( .A1(abar[3]), .A2(bbar[10]), .ZN(ybar[58]) );
  AND2_X1 U48 ( .A1(a[3]), .A2(b[9]), .ZN(y[57]) );
  OR2_X1 U48bar ( .A1(abar[3]), .A2(bbar[9]), .ZN(ybar[57]) );
  AND2_X1 U49 ( .A1(a[3]), .A2(b[8]), .ZN(y[56]) );
  OR2_X1 U49bar ( .A1(abar[3]), .A2(bbar[8]), .ZN(ybar[56]) );
  AND2_X1 U50 ( .A1(a[3]), .A2(b[7]), .ZN(y[55]) );
  OR2_X1 U50bar ( .A1(abar[3]), .A2(bbar[7]), .ZN(ybar[55]) );
  AND2_X1 U51 ( .A1(a[3]), .A2(b[6]), .ZN(y[54]) );
  OR2_X1 U51bar ( .A1(abar[3]), .A2(bbar[6]), .ZN(ybar[54]) );
  AND2_X1 U52 ( .A1(a[3]), .A2(b[5]), .ZN(y[53]) );
  OR2_X1 U52bar ( .A1(abar[3]), .A2(bbar[5]), .ZN(ybar[53]) );
  AND2_X1 U53 ( .A1(a[3]), .A2(b[4]), .ZN(y[52]) );
  OR2_X1 U53bar ( .A1(abar[3]), .A2(bbar[4]), .ZN(ybar[52]) );
  AND2_X1 U54 ( .A1(a[3]), .A2(b[3]), .ZN(y[51]) );
  OR2_X1 U54bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[51]) );
  AND2_X1 U55 ( .A1(a[3]), .A2(b[2]), .ZN(y[50]) );
  OR2_X1 U55bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[50]) );
  AND2_X1 U56 ( .A1(b[4]), .A2(a[0]), .ZN(y[4]) );
  OR2_X1 U56bar ( .A1(bbar[4]), .A2(abar[0]), .ZN(ybar[4]) );
  AND2_X1 U57 ( .A1(a[3]), .A2(b[1]), .ZN(y[49]) );
  OR2_X1 U57bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[49]) );
  AND2_X1 U58 ( .A1(a[3]), .A2(b[0]), .ZN(y[48]) );
  OR2_X1 U58bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[48]) );
  AND2_X1 U59 ( .A1(a[2]), .A2(b[15]), .ZN(y[47]) );
  OR2_X1 U59bar ( .A1(abar[2]), .A2(bbar[15]), .ZN(ybar[47]) );
  AND2_X1 U60 ( .A1(a[2]), .A2(b[14]), .ZN(y[46]) );
  OR2_X1 U60bar ( .A1(abar[2]), .A2(bbar[14]), .ZN(ybar[46]) );
  AND2_X1 U61 ( .A1(a[2]), .A2(b[13]), .ZN(y[45]) );
  OR2_X1 U61bar ( .A1(abar[2]), .A2(bbar[13]), .ZN(ybar[45]) );
  AND2_X1 U62 ( .A1(a[2]), .A2(b[12]), .ZN(y[44]) );
  OR2_X1 U62bar ( .A1(abar[2]), .A2(bbar[12]), .ZN(ybar[44]) );
  AND2_X1 U63 ( .A1(a[2]), .A2(b[11]), .ZN(y[43]) );
  OR2_X1 U63bar ( .A1(abar[2]), .A2(bbar[11]), .ZN(ybar[43]) );
  AND2_X1 U64 ( .A1(a[2]), .A2(b[10]), .ZN(y[42]) );
  OR2_X1 U64bar ( .A1(abar[2]), .A2(bbar[10]), .ZN(ybar[42]) );
  AND2_X1 U65 ( .A1(a[2]), .A2(b[9]), .ZN(y[41]) );
  OR2_X1 U65bar ( .A1(abar[2]), .A2(bbar[9]), .ZN(ybar[41]) );
  AND2_X1 U66 ( .A1(a[2]), .A2(b[8]), .ZN(y[40]) );
  OR2_X1 U66bar ( .A1(abar[2]), .A2(bbar[8]), .ZN(ybar[40]) );
  AND2_X1 U67 ( .A1(b[3]), .A2(a[0]), .ZN(y[3]) );
  OR2_X1 U67bar ( .A1(bbar[3]), .A2(abar[0]), .ZN(ybar[3]) );
  AND2_X1 U68 ( .A1(a[2]), .A2(b[7]), .ZN(y[39]) );
  OR2_X1 U68bar ( .A1(abar[2]), .A2(bbar[7]), .ZN(ybar[39]) );
  AND2_X1 U69 ( .A1(a[2]), .A2(b[6]), .ZN(y[38]) );
  OR2_X1 U69bar ( .A1(abar[2]), .A2(bbar[6]), .ZN(ybar[38]) );
  AND2_X1 U70 ( .A1(a[2]), .A2(b[5]), .ZN(y[37]) );
  OR2_X1 U70bar ( .A1(abar[2]), .A2(bbar[5]), .ZN(ybar[37]) );
  AND2_X1 U71 ( .A1(a[2]), .A2(b[4]), .ZN(y[36]) );
  OR2_X1 U71bar ( .A1(abar[2]), .A2(bbar[4]), .ZN(ybar[36]) );
  AND2_X1 U72 ( .A1(a[2]), .A2(b[3]), .ZN(y[35]) );
  OR2_X1 U72bar ( .A1(abar[2]), .A2(bbar[3]), .ZN(ybar[35]) );
  AND2_X1 U73 ( .A1(a[2]), .A2(b[2]), .ZN(y[34]) );
  OR2_X1 U73bar ( .A1(abar[2]), .A2(bbar[2]), .ZN(ybar[34]) );
  AND2_X1 U74 ( .A1(a[2]), .A2(b[1]), .ZN(y[33]) );
  OR2_X1 U74bar ( .A1(abar[2]), .A2(bbar[1]), .ZN(ybar[33]) );
  AND2_X1 U75 ( .A1(a[2]), .A2(b[0]), .ZN(y[32]) );
  OR2_X1 U75bar ( .A1(abar[2]), .A2(bbar[0]), .ZN(ybar[32]) );
  AND2_X1 U76 ( .A1(a[1]), .A2(b[15]), .ZN(y[31]) );
  OR2_X1 U76bar ( .A1(abar[1]), .A2(bbar[15]), .ZN(ybar[31]) );
  AND2_X1 U77 ( .A1(a[1]), .A2(b[14]), .ZN(y[30]) );
  OR2_X1 U77bar ( .A1(abar[1]), .A2(bbar[14]), .ZN(ybar[30]) );
  AND2_X1 U78 ( .A1(b[2]), .A2(a[0]), .ZN(y[2]) );
  OR2_X1 U78bar ( .A1(bbar[2]), .A2(abar[0]), .ZN(ybar[2]) );
  AND2_X1 U79 ( .A1(a[1]), .A2(b[13]), .ZN(y[29]) );
  OR2_X1 U79bar ( .A1(abar[1]), .A2(bbar[13]), .ZN(ybar[29]) );
  AND2_X1 U80 ( .A1(a[1]), .A2(b[12]), .ZN(y[28]) );
  OR2_X1 U80bar ( .A1(abar[1]), .A2(bbar[12]), .ZN(ybar[28]) );
  AND2_X1 U81 ( .A1(a[1]), .A2(b[11]), .ZN(y[27]) );
  OR2_X1 U81bar ( .A1(abar[1]), .A2(bbar[11]), .ZN(ybar[27]) );
  AND2_X1 U82 ( .A1(a[1]), .A2(b[10]), .ZN(y[26]) );
  OR2_X1 U82bar ( .A1(abar[1]), .A2(bbar[10]), .ZN(ybar[26]) );
  AND2_X1 U83 ( .A1(a[1]), .A2(b[9]), .ZN(y[25]) );
  OR2_X1 U83bar ( .A1(abar[1]), .A2(bbar[9]), .ZN(ybar[25]) );
  AND2_X1 U84 ( .A1(a[15]), .A2(b[15]), .ZN(y[255]) );
  OR2_X1 U84bar ( .A1(abar[15]), .A2(bbar[15]), .ZN(ybar[255]) );
  AND2_X1 U85 ( .A1(a[15]), .A2(b[14]), .ZN(y[254]) );
  OR2_X1 U85bar ( .A1(abar[15]), .A2(bbar[14]), .ZN(ybar[254]) );
  AND2_X1 U86 ( .A1(a[15]), .A2(b[13]), .ZN(y[253]) );
  OR2_X1 U86bar ( .A1(abar[15]), .A2(bbar[13]), .ZN(ybar[253]) );
  AND2_X1 U87 ( .A1(a[15]), .A2(b[12]), .ZN(y[252]) );
  OR2_X1 U87bar ( .A1(abar[15]), .A2(bbar[12]), .ZN(ybar[252]) );
  AND2_X1 U88 ( .A1(a[15]), .A2(b[11]), .ZN(y[251]) );
  OR2_X1 U88bar ( .A1(abar[15]), .A2(bbar[11]), .ZN(ybar[251]) );
  AND2_X1 U89 ( .A1(a[15]), .A2(b[10]), .ZN(y[250]) );
  OR2_X1 U89bar ( .A1(abar[15]), .A2(bbar[10]), .ZN(ybar[250]) );
  AND2_X1 U90 ( .A1(a[1]), .A2(b[8]), .ZN(y[24]) );
  OR2_X1 U90bar ( .A1(abar[1]), .A2(bbar[8]), .ZN(ybar[24]) );
  AND2_X1 U91 ( .A1(a[15]), .A2(b[9]), .ZN(y[249]) );
  OR2_X1 U91bar ( .A1(abar[15]), .A2(bbar[9]), .ZN(ybar[249]) );
  AND2_X1 U92 ( .A1(a[15]), .A2(b[8]), .ZN(y[248]) );
  OR2_X1 U92bar ( .A1(abar[15]), .A2(bbar[8]), .ZN(ybar[248]) );
  AND2_X1 U93 ( .A1(a[15]), .A2(b[7]), .ZN(y[247]) );
  OR2_X1 U93bar ( .A1(abar[15]), .A2(bbar[7]), .ZN(ybar[247]) );
  AND2_X1 U94 ( .A1(a[15]), .A2(b[6]), .ZN(y[246]) );
  OR2_X1 U94bar ( .A1(abar[15]), .A2(bbar[6]), .ZN(ybar[246]) );
  AND2_X1 U95 ( .A1(a[15]), .A2(b[5]), .ZN(y[245]) );
  OR2_X1 U95bar ( .A1(abar[15]), .A2(bbar[5]), .ZN(ybar[245]) );
  AND2_X1 U96 ( .A1(a[15]), .A2(b[4]), .ZN(y[244]) );
  OR2_X1 U96bar ( .A1(abar[15]), .A2(bbar[4]), .ZN(ybar[244]) );
  AND2_X1 U97 ( .A1(a[15]), .A2(b[3]), .ZN(y[243]) );
  OR2_X1 U97bar ( .A1(abar[15]), .A2(bbar[3]), .ZN(ybar[243]) );
  AND2_X1 U98 ( .A1(a[15]), .A2(b[2]), .ZN(y[242]) );
  OR2_X1 U98bar ( .A1(abar[15]), .A2(bbar[2]), .ZN(ybar[242]) );
  AND2_X1 U99 ( .A1(a[15]), .A2(b[1]), .ZN(y[241]) );
  OR2_X1 U99bar ( .A1(abar[15]), .A2(bbar[1]), .ZN(ybar[241]) );
  AND2_X1 U100 ( .A1(a[15]), .A2(b[0]), .ZN(y[240]) );
  OR2_X1 U100bar ( .A1(abar[15]), .A2(bbar[0]), .ZN(ybar[240]) );
  AND2_X1 U101 ( .A1(a[1]), .A2(b[7]), .ZN(y[23]) );
  OR2_X1 U101bar ( .A1(abar[1]), .A2(bbar[7]), .ZN(ybar[23]) );
  AND2_X1 U102 ( .A1(a[14]), .A2(b[15]), .ZN(y[239]) );
  OR2_X1 U102bar ( .A1(abar[14]), .A2(bbar[15]), .ZN(ybar[239]) );
  AND2_X1 U103 ( .A1(a[14]), .A2(b[14]), .ZN(y[238]) );
  OR2_X1 U103bar ( .A1(abar[14]), .A2(bbar[14]), .ZN(ybar[238]) );
  AND2_X1 U104 ( .A1(a[14]), .A2(b[13]), .ZN(y[237]) );
  OR2_X1 U104bar ( .A1(abar[14]), .A2(bbar[13]), .ZN(ybar[237]) );
  AND2_X1 U105 ( .A1(a[14]), .A2(b[12]), .ZN(y[236]) );
  OR2_X1 U105bar ( .A1(abar[14]), .A2(bbar[12]), .ZN(ybar[236]) );
  AND2_X1 U106 ( .A1(a[14]), .A2(b[11]), .ZN(y[235]) );
  OR2_X1 U106bar ( .A1(abar[14]), .A2(bbar[11]), .ZN(ybar[235]) );
  AND2_X1 U107 ( .A1(a[14]), .A2(b[10]), .ZN(y[234]) );
  OR2_X1 U107bar ( .A1(abar[14]), .A2(bbar[10]), .ZN(ybar[234]) );
  AND2_X1 U108 ( .A1(a[14]), .A2(b[9]), .ZN(y[233]) );
  OR2_X1 U108bar ( .A1(abar[14]), .A2(bbar[9]), .ZN(ybar[233]) );
  AND2_X1 U109 ( .A1(a[14]), .A2(b[8]), .ZN(y[232]) );
  OR2_X1 U109bar ( .A1(abar[14]), .A2(bbar[8]), .ZN(ybar[232]) );
  AND2_X1 U110 ( .A1(a[14]), .A2(b[7]), .ZN(y[231]) );
  OR2_X1 U110bar ( .A1(abar[14]), .A2(bbar[7]), .ZN(ybar[231]) );
  AND2_X1 U111 ( .A1(a[14]), .A2(b[6]), .ZN(y[230]) );
  OR2_X1 U111bar ( .A1(abar[14]), .A2(bbar[6]), .ZN(ybar[230]) );
  AND2_X1 U112 ( .A1(a[1]), .A2(b[6]), .ZN(y[22]) );
  OR2_X1 U112bar ( .A1(abar[1]), .A2(bbar[6]), .ZN(ybar[22]) );
  AND2_X1 U113 ( .A1(a[14]), .A2(b[5]), .ZN(y[229]) );
  OR2_X1 U113bar ( .A1(abar[14]), .A2(bbar[5]), .ZN(ybar[229]) );
  AND2_X1 U114 ( .A1(a[14]), .A2(b[4]), .ZN(y[228]) );
  OR2_X1 U114bar ( .A1(abar[14]), .A2(bbar[4]), .ZN(ybar[228]) );
  AND2_X1 U115 ( .A1(a[14]), .A2(b[3]), .ZN(y[227]) );
  OR2_X1 U115bar ( .A1(abar[14]), .A2(bbar[3]), .ZN(ybar[227]) );
  AND2_X1 U116 ( .A1(a[14]), .A2(b[2]), .ZN(y[226]) );
  OR2_X1 U116bar ( .A1(abar[14]), .A2(bbar[2]), .ZN(ybar[226]) );
  AND2_X1 U117 ( .A1(a[14]), .A2(b[1]), .ZN(y[225]) );
  OR2_X1 U117bar ( .A1(abar[14]), .A2(bbar[1]), .ZN(ybar[225]) );
  AND2_X1 U118 ( .A1(a[14]), .A2(b[0]), .ZN(y[224]) );
  OR2_X1 U118bar ( .A1(abar[14]), .A2(bbar[0]), .ZN(ybar[224]) );
  AND2_X1 U119 ( .A1(a[13]), .A2(b[15]), .ZN(y[223]) );
  OR2_X1 U119bar ( .A1(abar[13]), .A2(bbar[15]), .ZN(ybar[223]) );
  AND2_X1 U120 ( .A1(a[13]), .A2(b[14]), .ZN(y[222]) );
  OR2_X1 U120bar ( .A1(abar[13]), .A2(bbar[14]), .ZN(ybar[222]) );
  AND2_X1 U121 ( .A1(a[13]), .A2(b[13]), .ZN(y[221]) );
  OR2_X1 U121bar ( .A1(abar[13]), .A2(bbar[13]), .ZN(ybar[221]) );
  AND2_X1 U122 ( .A1(a[13]), .A2(b[12]), .ZN(y[220]) );
  OR2_X1 U122bar ( .A1(abar[13]), .A2(bbar[12]), .ZN(ybar[220]) );
  AND2_X1 U123 ( .A1(a[1]), .A2(b[5]), .ZN(y[21]) );
  OR2_X1 U123bar ( .A1(abar[1]), .A2(bbar[5]), .ZN(ybar[21]) );
  AND2_X1 U124 ( .A1(a[13]), .A2(b[11]), .ZN(y[219]) );
  OR2_X1 U124bar ( .A1(abar[13]), .A2(bbar[11]), .ZN(ybar[219]) );
  AND2_X1 U125 ( .A1(a[13]), .A2(b[10]), .ZN(y[218]) );
  OR2_X1 U125bar ( .A1(abar[13]), .A2(bbar[10]), .ZN(ybar[218]) );
  AND2_X1 U126 ( .A1(a[13]), .A2(b[9]), .ZN(y[217]) );
  OR2_X1 U126bar ( .A1(abar[13]), .A2(bbar[9]), .ZN(ybar[217]) );
  AND2_X1 U127 ( .A1(a[13]), .A2(b[8]), .ZN(y[216]) );
  OR2_X1 U127bar ( .A1(abar[13]), .A2(bbar[8]), .ZN(ybar[216]) );
  AND2_X1 U128 ( .A1(a[13]), .A2(b[7]), .ZN(y[215]) );
  OR2_X1 U128bar ( .A1(abar[13]), .A2(bbar[7]), .ZN(ybar[215]) );
  AND2_X1 U129 ( .A1(a[13]), .A2(b[6]), .ZN(y[214]) );
  OR2_X1 U129bar ( .A1(abar[13]), .A2(bbar[6]), .ZN(ybar[214]) );
  AND2_X1 U130 ( .A1(a[13]), .A2(b[5]), .ZN(y[213]) );
  OR2_X1 U130bar ( .A1(abar[13]), .A2(bbar[5]), .ZN(ybar[213]) );
  AND2_X1 U131 ( .A1(a[13]), .A2(b[4]), .ZN(y[212]) );
  OR2_X1 U131bar ( .A1(abar[13]), .A2(bbar[4]), .ZN(ybar[212]) );
  AND2_X1 U132 ( .A1(a[13]), .A2(b[3]), .ZN(y[211]) );
  OR2_X1 U132bar ( .A1(abar[13]), .A2(bbar[3]), .ZN(ybar[211]) );
  AND2_X1 U133 ( .A1(a[13]), .A2(b[2]), .ZN(y[210]) );
  OR2_X1 U133bar ( .A1(abar[13]), .A2(bbar[2]), .ZN(ybar[210]) );
  AND2_X1 U134 ( .A1(a[1]), .A2(b[4]), .ZN(y[20]) );
  OR2_X1 U134bar ( .A1(abar[1]), .A2(bbar[4]), .ZN(ybar[20]) );
  AND2_X1 U135 ( .A1(a[13]), .A2(b[1]), .ZN(y[209]) );
  OR2_X1 U135bar ( .A1(abar[13]), .A2(bbar[1]), .ZN(ybar[209]) );
  AND2_X1 U136 ( .A1(a[13]), .A2(b[0]), .ZN(y[208]) );
  OR2_X1 U136bar ( .A1(abar[13]), .A2(bbar[0]), .ZN(ybar[208]) );
  AND2_X1 U137 ( .A1(a[12]), .A2(b[15]), .ZN(y[207]) );
  OR2_X1 U137bar ( .A1(abar[12]), .A2(bbar[15]), .ZN(ybar[207]) );
  AND2_X1 U138 ( .A1(a[12]), .A2(b[14]), .ZN(y[206]) );
  OR2_X1 U138bar ( .A1(abar[12]), .A2(bbar[14]), .ZN(ybar[206]) );
  AND2_X1 U139 ( .A1(a[12]), .A2(b[13]), .ZN(y[205]) );
  OR2_X1 U139bar ( .A1(abar[12]), .A2(bbar[13]), .ZN(ybar[205]) );
  AND2_X1 U140 ( .A1(a[12]), .A2(b[12]), .ZN(y[204]) );
  OR2_X1 U140bar ( .A1(abar[12]), .A2(bbar[12]), .ZN(ybar[204]) );
  AND2_X1 U141 ( .A1(a[12]), .A2(b[11]), .ZN(y[203]) );
  OR2_X1 U141bar ( .A1(abar[12]), .A2(bbar[11]), .ZN(ybar[203]) );
  AND2_X1 U142 ( .A1(a[12]), .A2(b[10]), .ZN(y[202]) );
  OR2_X1 U142bar ( .A1(abar[12]), .A2(bbar[10]), .ZN(ybar[202]) );
  AND2_X1 U143 ( .A1(a[12]), .A2(b[9]), .ZN(y[201]) );
  OR2_X1 U143bar ( .A1(abar[12]), .A2(bbar[9]), .ZN(ybar[201]) );
  AND2_X1 U144 ( .A1(a[12]), .A2(b[8]), .ZN(y[200]) );
  OR2_X1 U144bar ( .A1(abar[12]), .A2(bbar[8]), .ZN(ybar[200]) );
  AND2_X1 U145 ( .A1(b[1]), .A2(a[0]), .ZN(y[1]) );
  OR2_X1 U145bar ( .A1(bbar[1]), .A2(abar[0]), .ZN(ybar[1]) );
  AND2_X1 U146 ( .A1(a[1]), .A2(b[3]), .ZN(y[19]) );
  OR2_X1 U146bar ( .A1(abar[1]), .A2(bbar[3]), .ZN(ybar[19]) );
  AND2_X1 U147 ( .A1(a[12]), .A2(b[7]), .ZN(y[199]) );
  OR2_X1 U147bar ( .A1(abar[12]), .A2(bbar[7]), .ZN(ybar[199]) );
  AND2_X1 U148 ( .A1(a[12]), .A2(b[6]), .ZN(y[198]) );
  OR2_X1 U148bar ( .A1(abar[12]), .A2(bbar[6]), .ZN(ybar[198]) );
  AND2_X1 U149 ( .A1(a[12]), .A2(b[5]), .ZN(y[197]) );
  OR2_X1 U149bar ( .A1(abar[12]), .A2(bbar[5]), .ZN(ybar[197]) );
  AND2_X1 U150 ( .A1(a[12]), .A2(b[4]), .ZN(y[196]) );
  OR2_X1 U150bar ( .A1(abar[12]), .A2(bbar[4]), .ZN(ybar[196]) );
  AND2_X1 U151 ( .A1(a[12]), .A2(b[3]), .ZN(y[195]) );
  OR2_X1 U151bar ( .A1(abar[12]), .A2(bbar[3]), .ZN(ybar[195]) );
  AND2_X1 U152 ( .A1(a[12]), .A2(b[2]), .ZN(y[194]) );
  OR2_X1 U152bar ( .A1(abar[12]), .A2(bbar[2]), .ZN(ybar[194]) );
  AND2_X1 U153 ( .A1(a[12]), .A2(b[1]), .ZN(y[193]) );
  OR2_X1 U153bar ( .A1(abar[12]), .A2(bbar[1]), .ZN(ybar[193]) );
  AND2_X1 U154 ( .A1(a[12]), .A2(b[0]), .ZN(y[192]) );
  OR2_X1 U154bar ( .A1(abar[12]), .A2(bbar[0]), .ZN(ybar[192]) );
  AND2_X1 U155 ( .A1(a[11]), .A2(b[15]), .ZN(y[191]) );
  OR2_X1 U155bar ( .A1(abar[11]), .A2(bbar[15]), .ZN(ybar[191]) );
  AND2_X1 U156 ( .A1(a[11]), .A2(b[14]), .ZN(y[190]) );
  OR2_X1 U156bar ( .A1(abar[11]), .A2(bbar[14]), .ZN(ybar[190]) );
  AND2_X1 U157 ( .A1(a[1]), .A2(b[2]), .ZN(y[18]) );
  OR2_X1 U157bar ( .A1(abar[1]), .A2(bbar[2]), .ZN(ybar[18]) );
  AND2_X1 U158 ( .A1(a[11]), .A2(b[13]), .ZN(y[189]) );
  OR2_X1 U158bar ( .A1(abar[11]), .A2(bbar[13]), .ZN(ybar[189]) );
  AND2_X1 U159 ( .A1(a[11]), .A2(b[12]), .ZN(y[188]) );
  OR2_X1 U159bar ( .A1(abar[11]), .A2(bbar[12]), .ZN(ybar[188]) );
  AND2_X1 U160 ( .A1(a[11]), .A2(b[11]), .ZN(y[187]) );
  OR2_X1 U160bar ( .A1(abar[11]), .A2(bbar[11]), .ZN(ybar[187]) );
  AND2_X1 U161 ( .A1(a[11]), .A2(b[10]), .ZN(y[186]) );
  OR2_X1 U161bar ( .A1(abar[11]), .A2(bbar[10]), .ZN(ybar[186]) );
  AND2_X1 U162 ( .A1(a[11]), .A2(b[9]), .ZN(y[185]) );
  OR2_X1 U162bar ( .A1(abar[11]), .A2(bbar[9]), .ZN(ybar[185]) );
  AND2_X1 U163 ( .A1(a[11]), .A2(b[8]), .ZN(y[184]) );
  OR2_X1 U163bar ( .A1(abar[11]), .A2(bbar[8]), .ZN(ybar[184]) );
  AND2_X1 U164 ( .A1(a[11]), .A2(b[7]), .ZN(y[183]) );
  OR2_X1 U164bar ( .A1(abar[11]), .A2(bbar[7]), .ZN(ybar[183]) );
  AND2_X1 U165 ( .A1(a[11]), .A2(b[6]), .ZN(y[182]) );
  OR2_X1 U165bar ( .A1(abar[11]), .A2(bbar[6]), .ZN(ybar[182]) );
  AND2_X1 U166 ( .A1(a[11]), .A2(b[5]), .ZN(y[181]) );
  OR2_X1 U166bar ( .A1(abar[11]), .A2(bbar[5]), .ZN(ybar[181]) );
  AND2_X1 U167 ( .A1(a[11]), .A2(b[4]), .ZN(y[180]) );
  OR2_X1 U167bar ( .A1(abar[11]), .A2(bbar[4]), .ZN(ybar[180]) );
  AND2_X1 U168 ( .A1(a[1]), .A2(b[1]), .ZN(y[17]) );
  OR2_X1 U168bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[17]) );
  AND2_X1 U169 ( .A1(a[11]), .A2(b[3]), .ZN(y[179]) );
  OR2_X1 U169bar ( .A1(abar[11]), .A2(bbar[3]), .ZN(ybar[179]) );
  AND2_X1 U170 ( .A1(a[11]), .A2(b[2]), .ZN(y[178]) );
  OR2_X1 U170bar ( .A1(abar[11]), .A2(bbar[2]), .ZN(ybar[178]) );
  AND2_X1 U171 ( .A1(a[11]), .A2(b[1]), .ZN(y[177]) );
  OR2_X1 U171bar ( .A1(abar[11]), .A2(bbar[1]), .ZN(ybar[177]) );
  AND2_X1 U172 ( .A1(a[11]), .A2(b[0]), .ZN(y[176]) );
  OR2_X1 U172bar ( .A1(abar[11]), .A2(bbar[0]), .ZN(ybar[176]) );
  AND2_X1 U173 ( .A1(a[10]), .A2(b[15]), .ZN(y[175]) );
  OR2_X1 U173bar ( .A1(abar[10]), .A2(bbar[15]), .ZN(ybar[175]) );
  AND2_X1 U174 ( .A1(a[10]), .A2(b[14]), .ZN(y[174]) );
  OR2_X1 U174bar ( .A1(abar[10]), .A2(bbar[14]), .ZN(ybar[174]) );
  AND2_X1 U175 ( .A1(a[10]), .A2(b[13]), .ZN(y[173]) );
  OR2_X1 U175bar ( .A1(abar[10]), .A2(bbar[13]), .ZN(ybar[173]) );
  AND2_X1 U176 ( .A1(a[10]), .A2(b[12]), .ZN(y[172]) );
  OR2_X1 U176bar ( .A1(abar[10]), .A2(bbar[12]), .ZN(ybar[172]) );
  AND2_X1 U177 ( .A1(a[10]), .A2(b[11]), .ZN(y[171]) );
  OR2_X1 U177bar ( .A1(abar[10]), .A2(bbar[11]), .ZN(ybar[171]) );
  AND2_X1 U178 ( .A1(a[10]), .A2(b[10]), .ZN(y[170]) );
  OR2_X1 U178bar ( .A1(abar[10]), .A2(bbar[10]), .ZN(ybar[170]) );
  AND2_X1 U179 ( .A1(a[1]), .A2(b[0]), .ZN(y[16]) );
  OR2_X1 U179bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[16]) );
  AND2_X1 U180 ( .A1(a[10]), .A2(b[9]), .ZN(y[169]) );
  OR2_X1 U180bar ( .A1(abar[10]), .A2(bbar[9]), .ZN(ybar[169]) );
  AND2_X1 U181 ( .A1(a[10]), .A2(b[8]), .ZN(y[168]) );
  OR2_X1 U181bar ( .A1(abar[10]), .A2(bbar[8]), .ZN(ybar[168]) );
  AND2_X1 U182 ( .A1(a[10]), .A2(b[7]), .ZN(y[167]) );
  OR2_X1 U182bar ( .A1(abar[10]), .A2(bbar[7]), .ZN(ybar[167]) );
  AND2_X1 U183 ( .A1(a[10]), .A2(b[6]), .ZN(y[166]) );
  OR2_X1 U183bar ( .A1(abar[10]), .A2(bbar[6]), .ZN(ybar[166]) );
  AND2_X1 U184 ( .A1(a[10]), .A2(b[5]), .ZN(y[165]) );
  OR2_X1 U184bar ( .A1(abar[10]), .A2(bbar[5]), .ZN(ybar[165]) );
  AND2_X1 U185 ( .A1(a[10]), .A2(b[4]), .ZN(y[164]) );
  OR2_X1 U185bar ( .A1(abar[10]), .A2(bbar[4]), .ZN(ybar[164]) );
  AND2_X1 U186 ( .A1(a[10]), .A2(b[3]), .ZN(y[163]) );
  OR2_X1 U186bar ( .A1(abar[10]), .A2(bbar[3]), .ZN(ybar[163]) );
  AND2_X1 U187 ( .A1(a[10]), .A2(b[2]), .ZN(y[162]) );
  OR2_X1 U187bar ( .A1(abar[10]), .A2(bbar[2]), .ZN(ybar[162]) );
  AND2_X1 U188 ( .A1(a[10]), .A2(b[1]), .ZN(y[161]) );
  OR2_X1 U188bar ( .A1(abar[10]), .A2(bbar[1]), .ZN(ybar[161]) );
  AND2_X1 U189 ( .A1(a[10]), .A2(b[0]), .ZN(y[160]) );
  OR2_X1 U189bar ( .A1(abar[10]), .A2(bbar[0]), .ZN(ybar[160]) );
  AND2_X1 U190 ( .A1(b[15]), .A2(a[0]), .ZN(y[15]) );
  OR2_X1 U190bar ( .A1(bbar[15]), .A2(abar[0]), .ZN(ybar[15]) );
  AND2_X1 U191 ( .A1(a[9]), .A2(b[15]), .ZN(y[159]) );
  OR2_X1 U191bar ( .A1(abar[9]), .A2(bbar[15]), .ZN(ybar[159]) );
  AND2_X1 U192 ( .A1(a[9]), .A2(b[14]), .ZN(y[158]) );
  OR2_X1 U192bar ( .A1(abar[9]), .A2(bbar[14]), .ZN(ybar[158]) );
  AND2_X1 U193 ( .A1(a[9]), .A2(b[13]), .ZN(y[157]) );
  OR2_X1 U193bar ( .A1(abar[9]), .A2(bbar[13]), .ZN(ybar[157]) );
  AND2_X1 U194 ( .A1(a[9]), .A2(b[12]), .ZN(y[156]) );
  OR2_X1 U194bar ( .A1(abar[9]), .A2(bbar[12]), .ZN(ybar[156]) );
  AND2_X1 U195 ( .A1(a[9]), .A2(b[11]), .ZN(y[155]) );
  OR2_X1 U195bar ( .A1(abar[9]), .A2(bbar[11]), .ZN(ybar[155]) );
  AND2_X1 U196 ( .A1(a[9]), .A2(b[10]), .ZN(y[154]) );
  OR2_X1 U196bar ( .A1(abar[9]), .A2(bbar[10]), .ZN(ybar[154]) );
  AND2_X1 U197 ( .A1(a[9]), .A2(b[9]), .ZN(y[153]) );
  OR2_X1 U197bar ( .A1(abar[9]), .A2(bbar[9]), .ZN(ybar[153]) );
  AND2_X1 U198 ( .A1(a[9]), .A2(b[8]), .ZN(y[152]) );
  OR2_X1 U198bar ( .A1(abar[9]), .A2(bbar[8]), .ZN(ybar[152]) );
  AND2_X1 U199 ( .A1(a[9]), .A2(b[7]), .ZN(y[151]) );
  OR2_X1 U199bar ( .A1(abar[9]), .A2(bbar[7]), .ZN(ybar[151]) );
  AND2_X1 U200 ( .A1(a[9]), .A2(b[6]), .ZN(y[150]) );
  OR2_X1 U200bar ( .A1(abar[9]), .A2(bbar[6]), .ZN(ybar[150]) );
  AND2_X1 U201 ( .A1(b[14]), .A2(a[0]), .ZN(y[14]) );
  OR2_X1 U201bar ( .A1(bbar[14]), .A2(abar[0]), .ZN(ybar[14]) );
  AND2_X1 U202 ( .A1(a[9]), .A2(b[5]), .ZN(y[149]) );
  OR2_X1 U202bar ( .A1(abar[9]), .A2(bbar[5]), .ZN(ybar[149]) );
  AND2_X1 U203 ( .A1(a[9]), .A2(b[4]), .ZN(y[148]) );
  OR2_X1 U203bar ( .A1(abar[9]), .A2(bbar[4]), .ZN(ybar[148]) );
  AND2_X1 U204 ( .A1(a[9]), .A2(b[3]), .ZN(y[147]) );
  OR2_X1 U204bar ( .A1(abar[9]), .A2(bbar[3]), .ZN(ybar[147]) );
  AND2_X1 U205 ( .A1(a[9]), .A2(b[2]), .ZN(y[146]) );
  OR2_X1 U205bar ( .A1(abar[9]), .A2(bbar[2]), .ZN(ybar[146]) );
  AND2_X1 U206 ( .A1(a[9]), .A2(b[1]), .ZN(y[145]) );
  OR2_X1 U206bar ( .A1(abar[9]), .A2(bbar[1]), .ZN(ybar[145]) );
  AND2_X1 U207 ( .A1(a[9]), .A2(b[0]), .ZN(y[144]) );
  OR2_X1 U207bar ( .A1(abar[9]), .A2(bbar[0]), .ZN(ybar[144]) );
  AND2_X1 U208 ( .A1(a[8]), .A2(b[15]), .ZN(y[143]) );
  OR2_X1 U208bar ( .A1(abar[8]), .A2(bbar[15]), .ZN(ybar[143]) );
  AND2_X1 U209 ( .A1(a[8]), .A2(b[14]), .ZN(y[142]) );
  OR2_X1 U209bar ( .A1(abar[8]), .A2(bbar[14]), .ZN(ybar[142]) );
  AND2_X1 U210 ( .A1(a[8]), .A2(b[13]), .ZN(y[141]) );
  OR2_X1 U210bar ( .A1(abar[8]), .A2(bbar[13]), .ZN(ybar[141]) );
  AND2_X1 U211 ( .A1(a[8]), .A2(b[12]), .ZN(y[140]) );
  OR2_X1 U211bar ( .A1(abar[8]), .A2(bbar[12]), .ZN(ybar[140]) );
  AND2_X1 U212 ( .A1(b[13]), .A2(a[0]), .ZN(y[13]) );
  OR2_X1 U212bar ( .A1(bbar[13]), .A2(abar[0]), .ZN(ybar[13]) );
  AND2_X1 U213 ( .A1(a[8]), .A2(b[11]), .ZN(y[139]) );
  OR2_X1 U213bar ( .A1(abar[8]), .A2(bbar[11]), .ZN(ybar[139]) );
  AND2_X1 U214 ( .A1(a[8]), .A2(b[10]), .ZN(y[138]) );
  OR2_X1 U214bar ( .A1(abar[8]), .A2(bbar[10]), .ZN(ybar[138]) );
  AND2_X1 U215 ( .A1(a[8]), .A2(b[9]), .ZN(y[137]) );
  OR2_X1 U215bar ( .A1(abar[8]), .A2(bbar[9]), .ZN(ybar[137]) );
  AND2_X1 U216 ( .A1(a[8]), .A2(b[8]), .ZN(y[136]) );
  OR2_X1 U216bar ( .A1(abar[8]), .A2(bbar[8]), .ZN(ybar[136]) );
  AND2_X1 U217 ( .A1(a[8]), .A2(b[7]), .ZN(y[135]) );
  OR2_X1 U217bar ( .A1(abar[8]), .A2(bbar[7]), .ZN(ybar[135]) );
  AND2_X1 U218 ( .A1(a[8]), .A2(b[6]), .ZN(y[134]) );
  OR2_X1 U218bar ( .A1(abar[8]), .A2(bbar[6]), .ZN(ybar[134]) );
  AND2_X1 U219 ( .A1(a[8]), .A2(b[5]), .ZN(y[133]) );
  OR2_X1 U219bar ( .A1(abar[8]), .A2(bbar[5]), .ZN(ybar[133]) );
  AND2_X1 U220 ( .A1(a[8]), .A2(b[4]), .ZN(y[132]) );
  OR2_X1 U220bar ( .A1(abar[8]), .A2(bbar[4]), .ZN(ybar[132]) );
  AND2_X1 U221 ( .A1(a[8]), .A2(b[3]), .ZN(y[131]) );
  OR2_X1 U221bar ( .A1(abar[8]), .A2(bbar[3]), .ZN(ybar[131]) );
  AND2_X1 U222 ( .A1(a[8]), .A2(b[2]), .ZN(y[130]) );
  OR2_X1 U222bar ( .A1(abar[8]), .A2(bbar[2]), .ZN(ybar[130]) );
  AND2_X1 U223 ( .A1(b[12]), .A2(a[0]), .ZN(y[12]) );
  OR2_X1 U223bar ( .A1(bbar[12]), .A2(abar[0]), .ZN(ybar[12]) );
  AND2_X1 U224 ( .A1(a[8]), .A2(b[1]), .ZN(y[129]) );
  OR2_X1 U224bar ( .A1(abar[8]), .A2(bbar[1]), .ZN(ybar[129]) );
  AND2_X1 U225 ( .A1(a[8]), .A2(b[0]), .ZN(y[128]) );
  OR2_X1 U225bar ( .A1(abar[8]), .A2(bbar[0]), .ZN(ybar[128]) );
  AND2_X1 U226 ( .A1(a[7]), .A2(b[15]), .ZN(y[127]) );
  OR2_X1 U226bar ( .A1(abar[7]), .A2(bbar[15]), .ZN(ybar[127]) );
  AND2_X1 U227 ( .A1(a[7]), .A2(b[14]), .ZN(y[126]) );
  OR2_X1 U227bar ( .A1(abar[7]), .A2(bbar[14]), .ZN(ybar[126]) );
  AND2_X1 U228 ( .A1(a[7]), .A2(b[13]), .ZN(y[125]) );
  OR2_X1 U228bar ( .A1(abar[7]), .A2(bbar[13]), .ZN(ybar[125]) );
  AND2_X1 U229 ( .A1(a[7]), .A2(b[12]), .ZN(y[124]) );
  OR2_X1 U229bar ( .A1(abar[7]), .A2(bbar[12]), .ZN(ybar[124]) );
  AND2_X1 U230 ( .A1(a[7]), .A2(b[11]), .ZN(y[123]) );
  OR2_X1 U230bar ( .A1(abar[7]), .A2(bbar[11]), .ZN(ybar[123]) );
  AND2_X1 U231 ( .A1(a[7]), .A2(b[10]), .ZN(y[122]) );
  OR2_X1 U231bar ( .A1(abar[7]), .A2(bbar[10]), .ZN(ybar[122]) );
  AND2_X1 U232 ( .A1(a[7]), .A2(b[9]), .ZN(y[121]) );
  OR2_X1 U232bar ( .A1(abar[7]), .A2(bbar[9]), .ZN(ybar[121]) );
  AND2_X1 U233 ( .A1(a[7]), .A2(b[8]), .ZN(y[120]) );
  OR2_X1 U233bar ( .A1(abar[7]), .A2(bbar[8]), .ZN(ybar[120]) );
  AND2_X1 U234 ( .A1(b[11]), .A2(a[0]), .ZN(y[11]) );
  OR2_X1 U234bar ( .A1(bbar[11]), .A2(abar[0]), .ZN(ybar[11]) );
  AND2_X1 U235 ( .A1(a[7]), .A2(b[7]), .ZN(y[119]) );
  OR2_X1 U235bar ( .A1(abar[7]), .A2(bbar[7]), .ZN(ybar[119]) );
  AND2_X1 U236 ( .A1(a[7]), .A2(b[6]), .ZN(y[118]) );
  OR2_X1 U236bar ( .A1(abar[7]), .A2(bbar[6]), .ZN(ybar[118]) );
  AND2_X1 U237 ( .A1(a[7]), .A2(b[5]), .ZN(y[117]) );
  OR2_X1 U237bar ( .A1(abar[7]), .A2(bbar[5]), .ZN(ybar[117]) );
  AND2_X1 U238 ( .A1(a[7]), .A2(b[4]), .ZN(y[116]) );
  OR2_X1 U238bar ( .A1(abar[7]), .A2(bbar[4]), .ZN(ybar[116]) );
  AND2_X1 U239 ( .A1(a[7]), .A2(b[3]), .ZN(y[115]) );
  OR2_X1 U239bar ( .A1(abar[7]), .A2(bbar[3]), .ZN(ybar[115]) );
  AND2_X1 U240 ( .A1(a[7]), .A2(b[2]), .ZN(y[114]) );
  OR2_X1 U240bar ( .A1(abar[7]), .A2(bbar[2]), .ZN(ybar[114]) );
  AND2_X1 U241 ( .A1(a[7]), .A2(b[1]), .ZN(y[113]) );
  OR2_X1 U241bar ( .A1(abar[7]), .A2(bbar[1]), .ZN(ybar[113]) );
  AND2_X1 U242 ( .A1(a[7]), .A2(b[0]), .ZN(y[112]) );
  OR2_X1 U242bar ( .A1(abar[7]), .A2(bbar[0]), .ZN(ybar[112]) );
  AND2_X1 U243 ( .A1(b[15]), .A2(a[6]), .ZN(y[111]) );
  OR2_X1 U243bar ( .A1(bbar[15]), .A2(abar[6]), .ZN(ybar[111]) );
  AND2_X1 U244 ( .A1(b[14]), .A2(a[6]), .ZN(y[110]) );
  OR2_X1 U244bar ( .A1(bbar[14]), .A2(abar[6]), .ZN(ybar[110]) );
  AND2_X1 U245 ( .A1(b[10]), .A2(a[0]), .ZN(y[10]) );
  OR2_X1 U245bar ( .A1(bbar[10]), .A2(abar[0]), .ZN(ybar[10]) );
  AND2_X1 U246 ( .A1(b[13]), .A2(a[6]), .ZN(y[109]) );
  OR2_X1 U246bar ( .A1(bbar[13]), .A2(abar[6]), .ZN(ybar[109]) );
  AND2_X1 U247 ( .A1(b[12]), .A2(a[6]), .ZN(y[108]) );
  OR2_X1 U247bar ( .A1(bbar[12]), .A2(abar[6]), .ZN(ybar[108]) );
  AND2_X1 U248 ( .A1(b[11]), .A2(a[6]), .ZN(y[107]) );
  OR2_X1 U248bar ( .A1(bbar[11]), .A2(abar[6]), .ZN(ybar[107]) );
  AND2_X1 U249 ( .A1(b[10]), .A2(a[6]), .ZN(y[106]) );
  OR2_X1 U249bar ( .A1(bbar[10]), .A2(abar[6]), .ZN(ybar[106]) );
  AND2_X1 U250 ( .A1(a[6]), .A2(b[9]), .ZN(y[105]) );
  OR2_X1 U250bar ( .A1(abar[6]), .A2(bbar[9]), .ZN(ybar[105]) );
  AND2_X1 U251 ( .A1(b[8]), .A2(a[6]), .ZN(y[104]) );
  OR2_X1 U251bar ( .A1(bbar[8]), .A2(abar[6]), .ZN(ybar[104]) );
  AND2_X1 U252 ( .A1(b[7]), .A2(a[6]), .ZN(y[103]) );
  OR2_X1 U252bar ( .A1(bbar[7]), .A2(abar[6]), .ZN(ybar[103]) );
  AND2_X1 U253 ( .A1(b[6]), .A2(a[6]), .ZN(y[102]) );
  OR2_X1 U253bar ( .A1(bbar[6]), .A2(abar[6]), .ZN(ybar[102]) );
  AND2_X1 U254 ( .A1(b[5]), .A2(a[6]), .ZN(y[101]) );
  OR2_X1 U254bar ( .A1(bbar[5]), .A2(abar[6]), .ZN(ybar[101]) );
  AND2_X1 U255 ( .A1(b[4]), .A2(a[6]), .ZN(y[100]) );
  OR2_X1 U255bar ( .A1(bbar[4]), .A2(abar[6]), .ZN(ybar[100]) );
  AND2_X1 U256 ( .A1(b[0]), .A2(a[0]), .ZN(y[0]) );
  OR2_X1 U256bar ( .A1(bbar[0]), .A2(abar[0]), .ZN(ybar[0]) );
endmodule

module decode_15 ( in, inbar, out, outbar );

  input wire [7:0] in;
  input wire [7:0] inbar;
//input_done

  output wire [255:0] out;
  output wire [255:0] outbar;
//output_done

  wire [15:0] level1;
  wire [31:0] level2;
  wire [15:0] level1bar;
  wire [31:0] level2bar;
//wire_done

  CD2_60 cd_l1_1 ( .a(in[1]), .abar(inbar[1]), .b(in[0]), .bbar(inbar[0]), .y(level1[3:0]), .ybar(level1bar[3:0]) );
  CD2_59 cd_l1_2 ( .a(in[3]), .abar(inbar[3]), .b(in[2]), .bbar(inbar[2]), .y(level1[7:4]), .ybar(level1bar[7:4]) );
  CD2_58 cd_l1_3 ( .a(in[5]), .abar(inbar[5]), .b(in[4]), .bbar(inbar[4]), .y(level1[11:8]), .ybar(level1bar[11:8]) );
  CD2_57 cd_l1_4 ( .a(in[7]), .abar(inbar[7]), .b(in[6]), .bbar(inbar[6]), .y(level1[15:12]), .ybar(level1bar[15:12]) );

  CD4_30 cd_l2_1 ( .a(level1[7:4]), .abar(level1bar[7:4]), .b(level1[3:0]), .bbar(level1bar[3:0]), 
        .y(level2[15:0]), .ybar(level2bar[15:0]) );
  CD4_29 cd_l2_2 ( .a(level1[15:12]), .abar(level1bar[15:12]), .b(level1[11:8]), .bbar(level1bar[11:8]), 
        .y(level2[31:16]), .ybar(level2bar[31:16]) );
  CD16_15 cd_l3 ( .a(level2[31:16]), .abar(level2bar[31:16]), .b(level2[15:0]), .bbar(level2bar[15:0]), 
        .y(out), .ybar(outbar) );
endmodule

module encode_15 ( in, inbar, out, outbar );

  input wire [255:0] in;
  input wire [255:0] inbar;
//input_done

  output wire [7:0] out;
  output wire [7:0] outbar;
//output_done

  wire in_81;
  wire in_80;
  wire in_79;
  wire in_78;
  wire in_77;
  wire in_76;
  wire in_75;
  wire in_74;
  wire in_73;
  wire in_72;
  wire in_71;
  wire in_70;
  wire in_69;
  wire in_68;
  wire in_67;
  wire in_66;
  wire in_65;
  wire in_64;
  wire in_63;
  wire in_62;
  wire in_61;
  wire in_60;
  wire in_59;
  wire in_58;
  wire in_57;
  wire in_56;
  wire in_55;
  wire in_54;
  wire in_53;
  wire in_52;
  wire in_51;
  wire in_50;
  wire in_49;
  wire in_48;
  wire in_47;
  wire in_46;
  wire in_45;
  wire in_44;
  wire in_43;
  wire in_42;
  wire in_41;
  wire in_40;
  wire in_39;
  wire in_38;
  wire in_37;
  wire in_36;
  wire in_35;
  wire in_34;
  wire in_33;
  wire in_32;
  wire in_31;
  wire in_30;
  wire in_29;
  wire in_28;
  wire in_27;
  wire in_26;
  wire in_25;
  wire in_24;
  wire in_23;
  wire in_22;
  wire in_21;
  wire in_20;
  wire in_19;
  wire in_18;
  wire in_17;
  wire in_16;
  wire in_15;
  wire in_14;
  wire in_13;
  wire in_12;
  wire in_11;
  wire in_10;
  wire in_9;
  wire in_8;
  wire in_7;
  wire in_6;
  wire in_5;
  wire in_4;
  wire in_3;
  wire in_2;
  wire in_1;
  wire in_0;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire in_81bar;
  wire in_80bar;
  wire in_79bar;
  wire in_78bar;
  wire in_77bar;
  wire in_76bar;
  wire in_75bar;
  wire in_74bar;
  wire in_73bar;
  wire in_72bar;
  wire in_71bar;
  wire in_70bar;
  wire in_69bar;
  wire in_68bar;
  wire in_67bar;
  wire in_66bar;
  wire in_65bar;
  wire in_64bar;
  wire in_63bar;
  wire in_62bar;
  wire in_61bar;
  wire in_60bar;
  wire in_59bar;
  wire in_58bar;
  wire in_57bar;
  wire in_56bar;
  wire in_55bar;
  wire in_54bar;
  wire in_53bar;
  wire in_52bar;
  wire in_51bar;
  wire in_50bar;
  wire in_49bar;
  wire in_48bar;
  wire in_47bar;
  wire in_46bar;
  wire in_45bar;
  wire in_44bar;
  wire in_43bar;
  wire in_42bar;
  wire in_41bar;
  wire in_40bar;
  wire in_39bar;
  wire in_38bar;
  wire in_37bar;
  wire in_36bar;
  wire in_35bar;
  wire in_34bar;
  wire in_33bar;
  wire in_32bar;
  wire in_31bar;
  wire in_30bar;
  wire in_29bar;
  wire in_28bar;
  wire in_27bar;
  wire in_26bar;
  wire in_25bar;
  wire in_24bar;
  wire in_23bar;
  wire in_22bar;
  wire in_21bar;
  wire in_20bar;
  wire in_19bar;
  wire in_18bar;
  wire in_17bar;
  wire in_16bar;
  wire in_15bar;
  wire in_14bar;
  wire in_13bar;
  wire in_12bar;
  wire in_11bar;
  wire in_10bar;
  wire in_9bar;
  wire in_8bar;
  wire in_7bar;
  wire in_6bar;
  wire in_5bar;
  wire in_4bar;
  wire in_3bar;
  wire in_2bar;
  wire in_1bar;
  wire in_0bar;
  wire n487bar;
  wire n488bar;
  wire n489bar;
  wire n490bar;
  wire n491bar;
  wire n492bar;
  wire n493bar;
  wire n494bar;
  wire n495bar;
  wire n496bar;
  wire n497bar;
  wire n498bar;
  wire n499bar;
  wire n500bar;
  wire n501bar;
  wire n502bar;
  wire n503bar;
  wire n504bar;
  wire n505bar;
  wire n506bar;
  wire n507bar;
  wire n508bar;
  wire n509bar;
  wire n510bar;
  wire n511bar;
  wire n512bar;
  wire n513bar;
  wire n514bar;
  wire n515bar;
  wire n516bar;
  wire n517bar;
  wire n518bar;
  wire n519bar;
  wire n520bar;
  wire n521bar;
  wire n522bar;
  wire n523bar;
  wire n524bar;
  wire n525bar;
  wire n526bar;
  wire n527bar;
  wire n528bar;
  wire n529bar;
  wire n530bar;
  wire n531bar;
  wire n532bar;
  wire n533bar;
  wire n534bar;
  wire n535bar;
  wire n536bar;
  wire n537bar;
  wire n538bar;
  wire n539bar;
  wire n540bar;
  wire n541bar;
  wire n542bar;
  wire n543bar;
  wire n544bar;
  wire n545bar;
  wire n546bar;
  wire n547bar;
  wire n548bar;
  wire n549bar;
  wire n550bar;
  wire n551bar;
  wire n552bar;
  wire n553bar;
  wire n554bar;
  wire n555bar;
  wire n556bar;
  wire n557bar;
  wire n558bar;
  wire n559bar;
  wire n560bar;
  wire n561bar;
  wire n562bar;
  wire n563bar;
  wire n564bar;
  wire n565bar;
  wire n566bar;
  wire n567bar;
  wire n568bar;
  wire n569bar;
  wire n570bar;
  wire n571bar;
  wire n572bar;
  wire n573bar;
  wire n574bar;
  wire n575bar;
  wire n576bar;
  wire n577bar;
  wire n578bar;
  wire n579bar;
  wire n580bar;
  wire n581bar;
  wire n582bar;
  wire n583bar;
  wire n584bar;
  wire n585bar;
  wire n586bar;
  wire n587bar;
  wire n588bar;
  wire n589bar;
  wire n590bar;
  wire n591bar;
  wire n592bar;
  wire n593bar;
  wire n594bar;
  wire n595bar;
  wire n596bar;
  wire n597bar;
  wire n598bar;
  wire n599bar;
  wire n600bar;
  wire n601bar;
  wire n602bar;
  wire n603bar;
  wire n604bar;
  wire n605bar;
  wire n606bar;
  wire n607bar;
  wire n608bar;
  wire n609bar;
  wire n610bar;
  wire n611bar;
  wire n612bar;
  wire n613bar;
  wire n614bar;
  wire n615bar;
  wire n616bar;
  wire n617bar;
  wire n618bar;
  wire n619bar;
  wire n620bar;
  wire n621bar;
  wire n622bar;
  wire n623bar;
  wire n624bar;
  wire n625bar;
  wire n626bar;
  wire n627bar;
  wire n628bar;
  wire n629bar;
  wire n630bar;
  wire n631bar;
  wire n632bar;
  wire n633bar;
  wire n634bar;
  wire n635bar;
  wire n636bar;
  wire n637bar;
  wire n638bar;
  wire n639bar;
  wire n640bar;
  wire n641bar;
  wire n642bar;
  wire n643bar;
  wire n644bar;
  wire n645bar;
  wire n646bar;
  wire n647bar;
  wire n648bar;
  wire n649bar;
  wire n650bar;
  wire n651bar;
  wire n652bar;
  wire n653bar;
  wire n654bar;
  wire n655bar;
  wire n656bar;
  wire n657bar;
  wire n658bar;
  wire n659bar;
  wire n660bar;
  wire n661bar;
  wire n662bar;
  wire n663bar;
  wire n664bar;
  wire n665bar;
  wire n666bar;
  wire n667bar;
  wire n668bar;
  wire n669bar;
  wire n670bar;
  wire n671bar;
  wire n672bar;
  wire n673bar;
  wire n674bar;
  wire n675bar;
  wire n676bar;
  wire n677bar;
  wire n678bar;
  wire n679bar;
  wire n680bar;
  wire n681bar;
  wire n682bar;
  wire n683bar;
  wire n684bar;
  wire n685bar;
  wire n686bar;
  wire n687bar;
  wire n688bar;
  wire n689bar;
  wire n690bar;
  wire n691bar;
  wire n692bar;
  wire n693bar;
  wire n694bar;
  wire n695bar;
  wire n696bar;
  wire n697bar;
  wire n698bar;
  wire n699bar;
  wire n700bar;
  wire n701bar;
  wire n702bar;
  wire n703bar;
  wire n704bar;
  wire n705bar;
  wire n706bar;
  wire n707bar;
  wire n708bar;
  wire n709bar;
  wire n710bar;
  wire n711bar;
  wire n712bar;
  wire n713bar;
  wire n714bar;
  wire n715bar;
  wire n716bar;
  wire n717bar;
  wire n718bar;
  wire n719bar;
  wire n720bar;
  wire n721bar;
  wire n722bar;
  wire n723bar;
  wire n724bar;
  wire n725bar;
  wire n726bar;
  wire n727bar;
  wire n728bar;
  wire n729bar;
  wire n730bar;
  wire n731bar;
  wire n732bar;
  wire n733bar;
  wire n734bar;
  wire n735bar;
  wire n736bar;
  wire n737bar;
  wire n738bar;
  wire n739bar;
  wire n740bar;
  wire n741bar;
  wire n742bar;
  wire n743bar;
  wire n744bar;
  wire n745bar;
  wire n746bar;
  wire n747bar;
  wire n748bar;
  wire n749bar;
  wire n750bar;
  wire n751bar;
  wire n752bar;
  wire n753bar;
  wire n754bar;
  wire n755bar;
  wire n756bar;
  wire n757bar;
  wire n758bar;
  wire n759bar;
  wire n760bar;
  wire n761bar;
  wire n762bar;
  wire n763bar;
  wire n764bar;
  wire n765bar;
  wire n766bar;
  wire n767bar;
  wire n768bar;
  wire n769bar;
  wire n770bar;
  wire n771bar;
  wire n772bar;
  wire n773bar;
  wire n774bar;
  wire n775bar;
  wire n776bar;
  wire n777bar;
  wire n778bar;
  wire n779bar;
  wire n780bar;
  wire n781bar;
  wire n782bar;
  wire n783bar;
  wire n784bar;
  wire n785bar;
  wire n786bar;
  wire n787bar;
  wire n788bar;
  wire n789bar;
  wire n790bar;
  wire n791bar;
  wire n792bar;
  wire n793bar;
  wire n794bar;
  wire n795bar;
  wire n796bar;
  wire n797bar;
  wire n798bar;
  wire n799bar;
  wire n800bar;
  wire n801bar;
  wire n802bar;
  wire n803bar;
  wire n804bar;
  wire n805bar;
  wire n806bar;
  wire n807bar;
  wire n808bar;
  wire n809bar;
  wire n810bar;
  wire n811bar;
  wire n812bar;
  wire n813bar;
  wire n814bar;
  wire n815bar;
  wire n816bar;
  wire n817bar;
  wire n818bar;
  wire n819bar;
  wire n820bar;
  wire n821bar;
  wire n822bar;
  wire n823bar;
  wire n824bar;
  wire n825bar;
  wire n826bar;
  wire n827bar;
  wire n828bar;
  wire n829bar;
  wire n830bar;
  wire n831bar;
  wire n832bar;
  wire n833bar;
  wire n834bar;
  wire n835bar;
  wire n836bar;
  wire n837bar;
  wire n838bar;
  wire n839bar;
  wire n840bar;
  wire n841bar;
  wire n842bar;
  wire n843bar;
  wire n844bar;
  wire n845bar;
  wire n846bar;
  wire n847bar;
  wire n848bar;
  wire n849bar;
  wire n850bar;
  wire n851bar;
  wire n852bar;
  wire n853bar;
  wire n854bar;
  wire n855bar;
  wire n856bar;
  wire n857bar;
  wire n858bar;
  wire n859bar;
  wire n860bar;
  wire n861bar;
  wire n862bar;
  wire n863bar;
  wire n864bar;
  wire n865bar;
  wire n866bar;
  wire n867bar;
  wire n868bar;
  wire n869bar;
  wire n870bar;
  wire n871bar;
  wire n872bar;
  wire n873bar;
  wire n874bar;
  wire n875bar;
  wire n876bar;
  wire n877bar;
  wire n878bar;
  wire n879bar;
  wire n880bar;
  wire n881bar;
  wire n882bar;
  wire n883bar;
  wire n884bar;
  wire n885bar;
  wire n886bar;
  wire n887bar;
  wire n888bar;
  wire n889bar;
  wire n890bar;
  wire n891bar;
  wire n892bar;
  wire n893bar;
  wire n894bar;
  wire n895bar;
  wire n896bar;
  wire n897bar;
  wire n898bar;
  wire n899bar;
  wire n900bar;
  wire n901bar;
  wire n902bar;
  wire n903bar;
  wire n904bar;
  wire n905bar;
  wire n906bar;
  wire n907bar;
  wire n908bar;
  wire n909bar;
  wire n910bar;
  wire n911bar;
  wire n912bar;
  wire n913bar;
  wire n914bar;
  wire n915bar;
  wire n916bar;
  wire n917bar;
  wire n918bar;
  wire n919bar;
  wire n920bar;
  wire n921bar;
  wire n922bar;
  wire n923bar;
  wire n924bar;
  wire n925bar;
  wire n926bar;
  wire n927bar;
  wire n928bar;
  wire n929bar;
  wire n930bar;
  wire n931bar;
  wire n932bar;
  wire n933bar;
  wire n934bar;
  wire n935bar;
  wire n936bar;
  wire n937bar;
  wire n938bar;
  wire n939bar;
  wire n940bar;
  wire n941bar;
  wire n942bar;
  wire n943bar;
  wire n944bar;
  wire n945bar;
  wire n946bar;
  wire n947bar;
  wire n948bar;
  wire n949bar;
  wire n950bar;
  wire n951bar;
  wire n952bar;
  wire n953bar;
  wire n954bar;
  wire n955bar;
  wire n956bar;
  wire n957bar;
  wire n958bar;
  wire n959bar;
  wire n960bar;
  wire n961bar;
  wire n962bar;
  wire n963bar;
  wire n964bar;
  wire n965bar;
  wire n966bar;
  wire n967bar;
  wire n968bar;
  wire n969bar;
  wire n970bar;
  wire n971bar;
  wire n972bar;
//wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];
  assign in_81bar = inbar[81];
  assign in_80bar = inbar[80];
  assign in_79bar = inbar[79];
  assign in_78bar = inbar[78];
  assign in_77bar = inbar[77];
  assign in_76bar = inbar[76];
  assign in_75bar = inbar[75];
  assign in_74bar = inbar[74];
  assign in_73bar = inbar[73];
  assign in_72bar = inbar[72];
  assign in_71bar = inbar[71];
  assign in_70bar = inbar[70];
  assign in_69bar = inbar[69];
  assign in_68bar = inbar[68];
  assign in_67bar = inbar[67];
  assign in_66bar = inbar[66];
  assign in_65bar = inbar[65];
  assign in_64bar = inbar[64];
  assign in_63bar = inbar[63];
  assign in_62bar = inbar[62];
  assign in_61bar = inbar[61];
  assign in_60bar = inbar[60];
  assign in_59bar = inbar[59];
  assign in_58bar = inbar[58];
  assign in_57bar = inbar[57];
  assign in_56bar = inbar[56];
  assign in_55bar = inbar[55];
  assign in_54bar = inbar[54];
  assign in_53bar = inbar[53];
  assign in_52bar = inbar[52];
  assign in_51bar = inbar[51];
  assign in_50bar = inbar[50];
  assign in_49bar = inbar[49];
  assign in_48bar = inbar[48];
  assign in_47bar = inbar[47];
  assign in_46bar = inbar[46];
  assign in_45bar = inbar[45];
  assign in_44bar = inbar[44];
  assign in_43bar = inbar[43];
  assign in_42bar = inbar[42];
  assign in_41bar = inbar[41];
  assign in_40bar = inbar[40];
  assign in_39bar = inbar[39];
  assign in_38bar = inbar[38];
  assign in_37bar = inbar[37];
  assign in_36bar = inbar[36];
  assign in_35bar = inbar[35];
  assign in_34bar = inbar[34];
  assign in_33bar = inbar[33];
  assign in_32bar = inbar[32];
  assign in_31bar = inbar[31];
  assign in_30bar = inbar[30];
  assign in_29bar = inbar[29];
  assign in_28bar = inbar[28];
  assign in_27bar = inbar[27];
  assign in_26bar = inbar[26];
  assign in_25bar = inbar[25];
  assign in_24bar = inbar[24];
  assign in_23bar = inbar[23];
  assign in_22bar = inbar[22];
  assign in_21bar = inbar[21];
  assign in_20bar = inbar[20];
  assign in_19bar = inbar[19];
  assign in_18bar = inbar[18];
  assign in_17bar = inbar[17];
  assign in_16bar = inbar[16];
  assign in_15bar = inbar[15];
  assign in_14bar = inbar[14];
  assign in_13bar = inbar[13];
  assign in_12bar = inbar[12];
  assign in_11bar = inbar[11];
  assign in_10bar = inbar[10];
  assign in_9bar = inbar[9];
  assign in_8bar = inbar[8];
  assign in_7bar = inbar[7];
  assign in_6bar = inbar[6];
  assign in_5bar = inbar[5];
  assign in_4bar = inbar[4];
  assign in_3bar = inbar[3];
  assign in_2bar = inbar[2];
  assign in_1bar = inbar[1];
  assign in_0bar = inbar[0];
//assign_done

  OR2_X1 U1 ( .A1(n972), .A2(n971), .ZN(out[7]) );
  AND2_X1 U1bar ( .A1(n972bar), .A2(n971bar), .ZN(outbar[7]) );
  OR2_X1 U2 ( .A1(n970), .A2(n969), .ZN(n971) );
  AND2_X1 U2bar ( .A1(n970bar), .A2(n969bar), .ZN(n971bar) );
  OR2_X1 U3 ( .A1(n968), .A2(n967), .ZN(n969) );
  AND2_X1 U3bar ( .A1(n968bar), .A2(n967bar), .ZN(n969bar) );
  OR2_X1 U4 ( .A1(n966), .A2(n965), .ZN(n967) );
  AND2_X1 U4bar ( .A1(n966bar), .A2(n965bar), .ZN(n967bar) );
  OR2_X1 U5 ( .A1(n964), .A2(n963), .ZN(n968) );
  AND2_X1 U5bar ( .A1(n964bar), .A2(n963bar), .ZN(n968bar) );
  OR2_X1 U6 ( .A1(in[116]), .A2(n962), .ZN(n963) );
  AND2_X1 U6bar ( .A1(inbar[116]), .A2(n962bar), .ZN(n963bar) );
  OR2_X1 U7 ( .A1(n961), .A2(n960), .ZN(n970) );
  AND2_X1 U7bar ( .A1(n961bar), .A2(n960bar), .ZN(n970bar) );
  OR2_X1 U8 ( .A1(in[150]), .A2(in[127]), .ZN(n960) );
  AND2_X1 U8bar ( .A1(inbar[150]), .A2(inbar[127]), .ZN(n960bar) );
  OR2_X1 U9 ( .A1(in[160]), .A2(n959), .ZN(n961) );
  AND2_X1 U9bar ( .A1(inbar[160]), .A2(n959bar), .ZN(n961bar) );
  OR2_X1 U10 ( .A1(in[252]), .A2(in[168]), .ZN(n959) );
  AND2_X1 U10bar ( .A1(inbar[252]), .A2(inbar[168]), .ZN(n959bar) );
  OR2_X1 U11 ( .A1(n958), .A2(n957), .ZN(n972) );
  AND2_X1 U11bar ( .A1(n958bar), .A2(n957bar), .ZN(n972bar) );
  OR2_X1 U12 ( .A1(n956), .A2(n955), .ZN(n957) );
  AND2_X1 U12bar ( .A1(n956bar), .A2(n955bar), .ZN(n957bar) );
  OR2_X1 U13 ( .A1(in_17), .A2(in[96]), .ZN(n955) );
  AND2_X1 U13bar ( .A1(in_17bar), .A2(inbar[96]), .ZN(n955bar) );
  OR2_X1 U14 ( .A1(in_23), .A2(n954), .ZN(n956) );
  AND2_X1 U14bar ( .A1(in_23bar), .A2(n954bar), .ZN(n956bar) );
  OR2_X1 U15 ( .A1(in_31), .A2(in_26), .ZN(n954) );
  AND2_X1 U15bar ( .A1(in_31bar), .A2(in_26bar), .ZN(n954bar) );
  OR2_X1 U16 ( .A1(n953), .A2(n952), .ZN(n958) );
  AND2_X1 U16bar ( .A1(n953bar), .A2(n952bar), .ZN(n958bar) );
  OR2_X1 U17 ( .A1(in_58), .A2(in_4), .ZN(n952) );
  AND2_X1 U17bar ( .A1(in_58bar), .A2(in_4bar), .ZN(n952bar) );
  OR2_X1 U18 ( .A1(in_59), .A2(n951), .ZN(n953) );
  AND2_X1 U18bar ( .A1(in_59bar), .A2(n951bar), .ZN(n953bar) );
  OR2_X1 U19 ( .A1(in_71), .A2(in_62), .ZN(n951) );
  AND2_X1 U19bar ( .A1(in_71bar), .A2(in_62bar), .ZN(n951bar) );
  OR2_X1 U20 ( .A1(n950), .A2(n949), .ZN(out[6]) );
  AND2_X1 U20bar ( .A1(n950bar), .A2(n949bar), .ZN(outbar[6]) );
  OR2_X1 U21 ( .A1(n948), .A2(n947), .ZN(n949) );
  AND2_X1 U21bar ( .A1(n948bar), .A2(n947bar), .ZN(n949bar) );
  OR2_X1 U22 ( .A1(n946), .A2(n945), .ZN(n947) );
  AND2_X1 U22bar ( .A1(n946bar), .A2(n945bar), .ZN(n947bar) );
  OR2_X1 U23 ( .A1(n944), .A2(n943), .ZN(n945) );
  AND2_X1 U23bar ( .A1(n944bar), .A2(n943bar), .ZN(n945bar) );
  OR2_X1 U24 ( .A1(n942), .A2(n941), .ZN(n946) );
  AND2_X1 U24bar ( .A1(n942bar), .A2(n941bar), .ZN(n946bar) );
  OR2_X1 U25 ( .A1(in[101]), .A2(n940), .ZN(n941) );
  AND2_X1 U25bar ( .A1(inbar[101]), .A2(n940bar), .ZN(n941bar) );
  OR2_X1 U26 ( .A1(n939), .A2(n938), .ZN(n948) );
  AND2_X1 U26bar ( .A1(n939bar), .A2(n938bar), .ZN(n948bar) );
  OR2_X1 U27 ( .A1(in[114]), .A2(in[104]), .ZN(n938) );
  AND2_X1 U27bar ( .A1(inbar[114]), .A2(inbar[104]), .ZN(n938bar) );
  OR2_X1 U28 ( .A1(in[128]), .A2(n937), .ZN(n939) );
  AND2_X1 U28bar ( .A1(inbar[128]), .A2(n937bar), .ZN(n939bar) );
  OR2_X1 U29 ( .A1(in[136]), .A2(in[134]), .ZN(n937) );
  AND2_X1 U29bar ( .A1(inbar[136]), .A2(inbar[134]), .ZN(n937bar) );
  OR2_X1 U30 ( .A1(n936), .A2(n935), .ZN(n950) );
  AND2_X1 U30bar ( .A1(n936bar), .A2(n935bar), .ZN(n950bar) );
  OR2_X1 U31 ( .A1(n934), .A2(n933), .ZN(n935) );
  AND2_X1 U31bar ( .A1(n934bar), .A2(n933bar), .ZN(n935bar) );
  OR2_X1 U32 ( .A1(in[177]), .A2(in[164]), .ZN(n933) );
  AND2_X1 U32bar ( .A1(inbar[177]), .A2(inbar[164]), .ZN(n933bar) );
  OR2_X1 U33 ( .A1(in[212]), .A2(n932), .ZN(n934) );
  AND2_X1 U33bar ( .A1(inbar[212]), .A2(n932bar), .ZN(n934bar) );
  OR2_X1 U34 ( .A1(in[248]), .A2(in[221]), .ZN(n932) );
  AND2_X1 U34bar ( .A1(inbar[248]), .A2(inbar[221]), .ZN(n932bar) );
  OR2_X1 U35 ( .A1(n931), .A2(n930), .ZN(n936) );
  AND2_X1 U35bar ( .A1(n931bar), .A2(n930bar), .ZN(n936bar) );
  OR2_X1 U36 ( .A1(in_18), .A2(in[93]), .ZN(n930) );
  AND2_X1 U36bar ( .A1(in_18bar), .A2(inbar[93]), .ZN(n930bar) );
  OR2_X1 U37 ( .A1(in_31), .A2(n929), .ZN(n931) );
  AND2_X1 U37bar ( .A1(in_31bar), .A2(n929bar), .ZN(n931bar) );
  OR2_X1 U38 ( .A1(in_7), .A2(in_39), .ZN(n929) );
  AND2_X1 U38bar ( .A1(in_7bar), .A2(in_39bar), .ZN(n929bar) );
  OR2_X1 U39 ( .A1(n928), .A2(n927), .ZN(out[5]) );
  AND2_X1 U39bar ( .A1(n928bar), .A2(n927bar), .ZN(outbar[5]) );
  OR2_X1 U40 ( .A1(n926), .A2(n925), .ZN(n927) );
  AND2_X1 U40bar ( .A1(n926bar), .A2(n925bar), .ZN(n927bar) );
  OR2_X1 U41 ( .A1(n924), .A2(n923), .ZN(n925) );
  AND2_X1 U41bar ( .A1(n924bar), .A2(n923bar), .ZN(n925bar) );
  OR2_X1 U42 ( .A1(n922), .A2(n921), .ZN(n923) );
  AND2_X1 U42bar ( .A1(n922bar), .A2(n921bar), .ZN(n923bar) );
  OR2_X1 U43 ( .A1(n940), .A2(n920), .ZN(n924) );
  AND2_X1 U43bar ( .A1(n940bar), .A2(n920bar), .ZN(n924bar) );
  OR2_X1 U44 ( .A1(in[111]), .A2(n919), .ZN(n920) );
  AND2_X1 U44bar ( .A1(inbar[111]), .A2(n919bar), .ZN(n920bar) );
  OR2_X1 U45 ( .A1(n918), .A2(n917), .ZN(n940) );
  AND2_X1 U45bar ( .A1(n918bar), .A2(n917bar), .ZN(n940bar) );
  OR2_X1 U46 ( .A1(n916), .A2(n915), .ZN(n917) );
  AND2_X1 U46bar ( .A1(n916bar), .A2(n915bar), .ZN(n917bar) );
  OR2_X1 U47 ( .A1(n914), .A2(n913), .ZN(n915) );
  AND2_X1 U47bar ( .A1(n914bar), .A2(n913bar), .ZN(n915bar) );
  OR2_X1 U48 ( .A1(in[140]), .A2(in[131]), .ZN(n913) );
  AND2_X1 U48bar ( .A1(inbar[140]), .A2(inbar[131]), .ZN(n913bar) );
  OR2_X1 U49 ( .A1(in[160]), .A2(in[144]), .ZN(n914) );
  AND2_X1 U49bar ( .A1(inbar[160]), .A2(inbar[144]), .ZN(n914bar) );
  OR2_X1 U50 ( .A1(n912), .A2(n911), .ZN(n916) );
  AND2_X1 U50bar ( .A1(n912bar), .A2(n911bar), .ZN(n916bar) );
  OR2_X1 U51 ( .A1(in[179]), .A2(in[174]), .ZN(n911) );
  AND2_X1 U51bar ( .A1(inbar[179]), .A2(inbar[174]), .ZN(n911bar) );
  OR2_X1 U52 ( .A1(in[188]), .A2(in[184]), .ZN(n912) );
  AND2_X1 U52bar ( .A1(inbar[188]), .A2(inbar[184]), .ZN(n912bar) );
  OR2_X1 U53 ( .A1(n910), .A2(n909), .ZN(n918) );
  AND2_X1 U53bar ( .A1(n910bar), .A2(n909bar), .ZN(n918bar) );
  OR2_X1 U54 ( .A1(n908), .A2(n907), .ZN(n909) );
  AND2_X1 U54bar ( .A1(n908bar), .A2(n907bar), .ZN(n909bar) );
  OR2_X1 U55 ( .A1(in[216]), .A2(in[200]), .ZN(n907) );
  AND2_X1 U55bar ( .A1(inbar[216]), .A2(inbar[200]), .ZN(n907bar) );
  OR2_X1 U56 ( .A1(in[228]), .A2(in[224]), .ZN(n908) );
  AND2_X1 U56bar ( .A1(inbar[228]), .A2(inbar[224]), .ZN(n908bar) );
  OR2_X1 U57 ( .A1(n906), .A2(n905), .ZN(n910) );
  AND2_X1 U57bar ( .A1(n906bar), .A2(n905bar), .ZN(n910bar) );
  OR2_X1 U58 ( .A1(in[247]), .A2(in[235]), .ZN(n905) );
  AND2_X1 U58bar ( .A1(inbar[247]), .A2(inbar[235]), .ZN(n905bar) );
  OR2_X1 U59 ( .A1(in_42), .A2(in[83]), .ZN(n906) );
  AND2_X1 U59bar ( .A1(in_42bar), .A2(inbar[83]), .ZN(n906bar) );
  OR2_X1 U60 ( .A1(n904), .A2(n903), .ZN(n926) );
  AND2_X1 U60bar ( .A1(n904bar), .A2(n903bar), .ZN(n926bar) );
  OR2_X1 U61 ( .A1(in[166]), .A2(in[123]), .ZN(n903) );
  AND2_X1 U61bar ( .A1(inbar[166]), .A2(inbar[123]), .ZN(n903bar) );
  OR2_X1 U62 ( .A1(in[170]), .A2(n902), .ZN(n904) );
  AND2_X1 U62bar ( .A1(inbar[170]), .A2(n902bar), .ZN(n904bar) );
  OR2_X1 U63 ( .A1(in[194]), .A2(in[183]), .ZN(n902) );
  AND2_X1 U63bar ( .A1(inbar[194]), .A2(inbar[183]), .ZN(n902bar) );
  OR2_X1 U64 ( .A1(n901), .A2(n900), .ZN(n928) );
  AND2_X1 U64bar ( .A1(n901bar), .A2(n900bar), .ZN(n928bar) );
  OR2_X1 U65 ( .A1(n899), .A2(n898), .ZN(n900) );
  AND2_X1 U65bar ( .A1(n899bar), .A2(n898bar), .ZN(n900bar) );
  OR2_X1 U66 ( .A1(in[241]), .A2(in[238]), .ZN(n898) );
  AND2_X1 U66bar ( .A1(inbar[241]), .A2(inbar[238]), .ZN(n898bar) );
  OR2_X1 U67 ( .A1(in[250]), .A2(n897), .ZN(n899) );
  AND2_X1 U67bar ( .A1(inbar[250]), .A2(n897bar), .ZN(n899bar) );
  OR2_X1 U68 ( .A1(in_24), .A2(in[84]), .ZN(n897) );
  AND2_X1 U68bar ( .A1(in_24bar), .A2(inbar[84]), .ZN(n897bar) );
  OR2_X1 U69 ( .A1(n896), .A2(n895), .ZN(n901) );
  AND2_X1 U69bar ( .A1(n896bar), .A2(n895bar), .ZN(n901bar) );
  OR2_X1 U70 ( .A1(in_41), .A2(in_29), .ZN(n895) );
  AND2_X1 U70bar ( .A1(in_41bar), .A2(in_29bar), .ZN(n895bar) );
  OR2_X1 U71 ( .A1(in_66), .A2(n894), .ZN(n896) );
  AND2_X1 U71bar ( .A1(in_66bar), .A2(n894bar), .ZN(n896bar) );
  OR2_X1 U72 ( .A1(in_76), .A2(in_71), .ZN(n894) );
  AND2_X1 U72bar ( .A1(in_76bar), .A2(in_71bar), .ZN(n894bar) );
  OR2_X1 U73 ( .A1(n893), .A2(n892), .ZN(out[4]) );
  AND2_X1 U73bar ( .A1(n893bar), .A2(n892bar), .ZN(outbar[4]) );
  OR2_X1 U74 ( .A1(n891), .A2(n890), .ZN(n892) );
  AND2_X1 U74bar ( .A1(n891bar), .A2(n890bar), .ZN(n892bar) );
  OR2_X1 U75 ( .A1(n889), .A2(n888), .ZN(n890) );
  AND2_X1 U75bar ( .A1(n889bar), .A2(n888bar), .ZN(n890bar) );
  OR2_X1 U76 ( .A1(n922), .A2(n887), .ZN(n888) );
  AND2_X1 U76bar ( .A1(n922bar), .A2(n887bar), .ZN(n888bar) );
  OR2_X1 U77 ( .A1(n886), .A2(n885), .ZN(n922) );
  AND2_X1 U77bar ( .A1(n886bar), .A2(n885bar), .ZN(n922bar) );
  OR2_X1 U78 ( .A1(n884), .A2(n883), .ZN(n885) );
  AND2_X1 U78bar ( .A1(n884bar), .A2(n883bar), .ZN(n885bar) );
  OR2_X1 U79 ( .A1(n882), .A2(n881), .ZN(n883) );
  AND2_X1 U79bar ( .A1(n882bar), .A2(n881bar), .ZN(n883bar) );
  OR2_X1 U80 ( .A1(in[118]), .A2(in[109]), .ZN(n881) );
  AND2_X1 U80bar ( .A1(inbar[118]), .A2(inbar[109]), .ZN(n881bar) );
  OR2_X1 U81 ( .A1(in[139]), .A2(in[120]), .ZN(n882) );
  AND2_X1 U81bar ( .A1(inbar[139]), .A2(inbar[120]), .ZN(n882bar) );
  OR2_X1 U82 ( .A1(n880), .A2(n879), .ZN(n884) );
  AND2_X1 U82bar ( .A1(n880bar), .A2(n879bar), .ZN(n884bar) );
  OR2_X1 U83 ( .A1(in[198]), .A2(in[154]), .ZN(n879) );
  AND2_X1 U83bar ( .A1(inbar[198]), .A2(inbar[154]), .ZN(n879bar) );
  OR2_X1 U84 ( .A1(in[210]), .A2(in[205]), .ZN(n880) );
  AND2_X1 U84bar ( .A1(inbar[210]), .A2(inbar[205]), .ZN(n880bar) );
  OR2_X1 U85 ( .A1(n878), .A2(n877), .ZN(n886) );
  AND2_X1 U85bar ( .A1(n878bar), .A2(n877bar), .ZN(n886bar) );
  OR2_X1 U86 ( .A1(n876), .A2(n875), .ZN(n877) );
  AND2_X1 U86bar ( .A1(n876bar), .A2(n875bar), .ZN(n877bar) );
  OR2_X1 U87 ( .A1(in[219]), .A2(in[217]), .ZN(n875) );
  AND2_X1 U87bar ( .A1(inbar[219]), .A2(inbar[217]), .ZN(n875bar) );
  OR2_X1 U88 ( .A1(in[86]), .A2(in[252]), .ZN(n876) );
  AND2_X1 U88bar ( .A1(inbar[86]), .A2(inbar[252]), .ZN(n876bar) );
  OR2_X1 U89 ( .A1(n874), .A2(n873), .ZN(n878) );
  AND2_X1 U89bar ( .A1(n874bar), .A2(n873bar), .ZN(n878bar) );
  OR2_X1 U90 ( .A1(in_40), .A2(in[91]), .ZN(n873) );
  AND2_X1 U90bar ( .A1(in_40bar), .A2(inbar[91]), .ZN(n873bar) );
  OR2_X1 U91 ( .A1(in_8), .A2(in_46), .ZN(n874) );
  AND2_X1 U91bar ( .A1(in_8bar), .A2(in_46bar), .ZN(n874bar) );
  OR2_X1 U92 ( .A1(n872), .A2(n871), .ZN(n889) );
  AND2_X1 U92bar ( .A1(n872bar), .A2(n871bar), .ZN(n889bar) );
  OR2_X1 U93 ( .A1(in[117]), .A2(n943), .ZN(n871) );
  AND2_X1 U93bar ( .A1(inbar[117]), .A2(n943bar), .ZN(n871bar) );
  OR2_X1 U94 ( .A1(n870), .A2(n869), .ZN(n943) );
  AND2_X1 U94bar ( .A1(n870bar), .A2(n869bar), .ZN(n943bar) );
  OR2_X1 U95 ( .A1(n868), .A2(n867), .ZN(n869) );
  AND2_X1 U95bar ( .A1(n868bar), .A2(n867bar), .ZN(n869bar) );
  OR2_X1 U96 ( .A1(n866), .A2(n865), .ZN(n867) );
  AND2_X1 U96bar ( .A1(n866bar), .A2(n865bar), .ZN(n867bar) );
  OR2_X1 U97 ( .A1(n864), .A2(n863), .ZN(n865) );
  AND2_X1 U97bar ( .A1(n864bar), .A2(n863bar), .ZN(n865bar) );
  OR2_X1 U98 ( .A1(in[108]), .A2(n919), .ZN(n866) );
  AND2_X1 U98bar ( .A1(inbar[108]), .A2(n919bar), .ZN(n866bar) );
  OR2_X1 U99 ( .A1(n862), .A2(n861), .ZN(n919) );
  AND2_X1 U99bar ( .A1(n862bar), .A2(n861bar), .ZN(n919bar) );
  OR2_X1 U100 ( .A1(n860), .A2(n859), .ZN(n861) );
  AND2_X1 U100bar ( .A1(n860bar), .A2(n859bar), .ZN(n861bar) );
  OR2_X1 U101 ( .A1(n858), .A2(n857), .ZN(n859) );
  AND2_X1 U101bar ( .A1(n858bar), .A2(n857bar), .ZN(n859bar) );
  OR2_X1 U102 ( .A1(in[119]), .A2(in[105]), .ZN(n857) );
  AND2_X1 U102bar ( .A1(inbar[119]), .A2(inbar[105]), .ZN(n857bar) );
  OR2_X1 U103 ( .A1(in[186]), .A2(in[175]), .ZN(n858) );
  AND2_X1 U103bar ( .A1(inbar[186]), .A2(inbar[175]), .ZN(n858bar) );
  OR2_X1 U104 ( .A1(n856), .A2(n855), .ZN(n860) );
  AND2_X1 U104bar ( .A1(n856bar), .A2(n855bar), .ZN(n860bar) );
  OR2_X1 U105 ( .A1(in[202]), .A2(in[193]), .ZN(n855) );
  AND2_X1 U105bar ( .A1(inbar[202]), .A2(inbar[193]), .ZN(n855bar) );
  OR2_X1 U106 ( .A1(in[225]), .A2(in[208]), .ZN(n856) );
  AND2_X1 U106bar ( .A1(inbar[225]), .A2(inbar[208]), .ZN(n856bar) );
  OR2_X1 U107 ( .A1(n854), .A2(n853), .ZN(n862) );
  AND2_X1 U107bar ( .A1(n854bar), .A2(n853bar), .ZN(n862bar) );
  OR2_X1 U108 ( .A1(n852), .A2(n851), .ZN(n853) );
  AND2_X1 U108bar ( .A1(n852bar), .A2(n851bar), .ZN(n853bar) );
  OR2_X1 U109 ( .A1(in_1), .A2(in[85]), .ZN(n851) );
  AND2_X1 U109bar ( .A1(in_1bar), .A2(inbar[85]), .ZN(n851bar) );
  OR2_X1 U110 ( .A1(in_23), .A2(in_19), .ZN(n852) );
  AND2_X1 U110bar ( .A1(in_23bar), .A2(in_19bar), .ZN(n852bar) );
  OR2_X1 U111 ( .A1(n850), .A2(n849), .ZN(n854) );
  AND2_X1 U111bar ( .A1(n850bar), .A2(n849bar), .ZN(n854bar) );
  OR2_X1 U112 ( .A1(in_43), .A2(in_33), .ZN(n849) );
  AND2_X1 U112bar ( .A1(in_43bar), .A2(in_33bar), .ZN(n849bar) );
  OR2_X1 U113 ( .A1(in_63), .A2(in_44), .ZN(n850) );
  AND2_X1 U113bar ( .A1(in_63bar), .A2(in_44bar), .ZN(n850bar) );
  OR2_X1 U114 ( .A1(n848), .A2(n847), .ZN(n868) );
  AND2_X1 U114bar ( .A1(n848bar), .A2(n847bar), .ZN(n868bar) );
  OR2_X1 U115 ( .A1(in[141]), .A2(in[112]), .ZN(n847) );
  AND2_X1 U115bar ( .A1(inbar[141]), .A2(inbar[112]), .ZN(n847bar) );
  OR2_X1 U116 ( .A1(in[147]), .A2(n846), .ZN(n848) );
  AND2_X1 U116bar ( .A1(inbar[147]), .A2(n846bar), .ZN(n848bar) );
  OR2_X1 U117 ( .A1(in[181]), .A2(in[167]), .ZN(n846) );
  AND2_X1 U117bar ( .A1(inbar[181]), .A2(inbar[167]), .ZN(n846bar) );
  OR2_X1 U118 ( .A1(n845), .A2(n844), .ZN(n870) );
  AND2_X1 U118bar ( .A1(n845bar), .A2(n844bar), .ZN(n870bar) );
  OR2_X1 U119 ( .A1(n843), .A2(n842), .ZN(n844) );
  AND2_X1 U119bar ( .A1(n843bar), .A2(n842bar), .ZN(n844bar) );
  OR2_X1 U120 ( .A1(in[229]), .A2(in[201]), .ZN(n842) );
  AND2_X1 U120bar ( .A1(inbar[229]), .A2(inbar[201]), .ZN(n842bar) );
  OR2_X1 U121 ( .A1(in[237]), .A2(n841), .ZN(n843) );
  AND2_X1 U121bar ( .A1(inbar[237]), .A2(n841bar), .ZN(n843bar) );
  OR2_X1 U122 ( .A1(in[94]), .A2(in[253]), .ZN(n841) );
  AND2_X1 U122bar ( .A1(inbar[94]), .A2(inbar[253]), .ZN(n841bar) );
  OR2_X1 U123 ( .A1(n840), .A2(n839), .ZN(n845) );
  AND2_X1 U123bar ( .A1(n840bar), .A2(n839bar), .ZN(n845bar) );
  OR2_X1 U124 ( .A1(in_21), .A2(in[96]), .ZN(n839) );
  AND2_X1 U124bar ( .A1(in_21bar), .A2(inbar[96]), .ZN(n839bar) );
  OR2_X1 U125 ( .A1(in_25), .A2(n838), .ZN(n840) );
  AND2_X1 U125bar ( .A1(in_25bar), .A2(n838bar), .ZN(n840bar) );
  OR2_X1 U126 ( .A1(in_81), .A2(in_45), .ZN(n838) );
  AND2_X1 U126bar ( .A1(in_81bar), .A2(in_45bar), .ZN(n838bar) );
  OR2_X1 U127 ( .A1(n837), .A2(n836), .ZN(n891) );
  AND2_X1 U127bar ( .A1(n837bar), .A2(n836bar), .ZN(n891bar) );
  OR2_X1 U128 ( .A1(in[142]), .A2(in[124]), .ZN(n836) );
  AND2_X1 U128bar ( .A1(inbar[142]), .A2(inbar[124]), .ZN(n836bar) );
  OR2_X1 U129 ( .A1(in[150]), .A2(n835), .ZN(n837) );
  AND2_X1 U129bar ( .A1(inbar[150]), .A2(n835bar), .ZN(n837bar) );
  OR2_X1 U130 ( .A1(in[172]), .A2(in[155]), .ZN(n835) );
  AND2_X1 U130bar ( .A1(inbar[172]), .A2(inbar[155]), .ZN(n835bar) );
  OR2_X1 U131 ( .A1(n834), .A2(n833), .ZN(n893) );
  AND2_X1 U131bar ( .A1(n834bar), .A2(n833bar), .ZN(n893bar) );
  OR2_X1 U132 ( .A1(n832), .A2(n831), .ZN(n833) );
  AND2_X1 U132bar ( .A1(n832bar), .A2(n831bar), .ZN(n833bar) );
  OR2_X1 U133 ( .A1(in[196]), .A2(in[173]), .ZN(n831) );
  AND2_X1 U133bar ( .A1(inbar[196]), .A2(inbar[173]), .ZN(n831bar) );
  OR2_X1 U134 ( .A1(in[222]), .A2(n830), .ZN(n832) );
  AND2_X1 U134bar ( .A1(inbar[222]), .A2(n830bar), .ZN(n832bar) );
  OR2_X1 U135 ( .A1(in[227]), .A2(in[226]), .ZN(n830) );
  AND2_X1 U135bar ( .A1(inbar[227]), .A2(inbar[226]), .ZN(n830bar) );
  OR2_X1 U136 ( .A1(n829), .A2(n828), .ZN(n834) );
  AND2_X1 U136bar ( .A1(n829bar), .A2(n828bar), .ZN(n834bar) );
  OR2_X1 U137 ( .A1(in[249]), .A2(in[231]), .ZN(n828) );
  AND2_X1 U137bar ( .A1(inbar[249]), .A2(inbar[231]), .ZN(n828bar) );
  OR2_X1 U138 ( .A1(in_28), .A2(n827), .ZN(n829) );
  AND2_X1 U138bar ( .A1(in_28bar), .A2(n827bar), .ZN(n829bar) );
  OR2_X1 U139 ( .A1(in_52), .A2(in_47), .ZN(n827) );
  AND2_X1 U139bar ( .A1(in_52bar), .A2(in_47bar), .ZN(n827bar) );
  OR2_X1 U140 ( .A1(n826), .A2(n825), .ZN(out[3]) );
  AND2_X1 U140bar ( .A1(n826bar), .A2(n825bar), .ZN(outbar[3]) );
  OR2_X1 U141 ( .A1(n824), .A2(n823), .ZN(n825) );
  AND2_X1 U141bar ( .A1(n824bar), .A2(n823bar), .ZN(n825bar) );
  OR2_X1 U142 ( .A1(n822), .A2(n821), .ZN(n823) );
  AND2_X1 U142bar ( .A1(n822bar), .A2(n821bar), .ZN(n823bar) );
  OR2_X1 U143 ( .A1(n820), .A2(n819), .ZN(n821) );
  AND2_X1 U143bar ( .A1(n820bar), .A2(n819bar), .ZN(n821bar) );
  OR2_X1 U144 ( .A1(n964), .A2(n818), .ZN(n822) );
  AND2_X1 U144bar ( .A1(n964bar), .A2(n818bar), .ZN(n822bar) );
  OR2_X1 U145 ( .A1(in[118]), .A2(n817), .ZN(n818) );
  AND2_X1 U145bar ( .A1(inbar[118]), .A2(n817bar), .ZN(n818bar) );
  OR2_X1 U146 ( .A1(n816), .A2(n815), .ZN(n964) );
  AND2_X1 U146bar ( .A1(n816bar), .A2(n815bar), .ZN(n964bar) );
  OR2_X1 U147 ( .A1(n814), .A2(n813), .ZN(n815) );
  AND2_X1 U147bar ( .A1(n814bar), .A2(n813bar), .ZN(n815bar) );
  OR2_X1 U148 ( .A1(n812), .A2(n811), .ZN(n813) );
  AND2_X1 U148bar ( .A1(n812bar), .A2(n811bar), .ZN(n813bar) );
  OR2_X1 U149 ( .A1(in[122]), .A2(in[111]), .ZN(n811) );
  AND2_X1 U149bar ( .A1(inbar[122]), .A2(inbar[111]), .ZN(n811bar) );
  OR2_X1 U150 ( .A1(in[154]), .A2(in[151]), .ZN(n812) );
  AND2_X1 U150bar ( .A1(inbar[154]), .A2(inbar[151]), .ZN(n812bar) );
  OR2_X1 U151 ( .A1(n810), .A2(n809), .ZN(n814) );
  AND2_X1 U151bar ( .A1(n810bar), .A2(n809bar), .ZN(n814bar) );
  OR2_X1 U152 ( .A1(in[187]), .A2(in[177]), .ZN(n809) );
  AND2_X1 U152bar ( .A1(inbar[187]), .A2(inbar[177]), .ZN(n809bar) );
  OR2_X1 U153 ( .A1(in[200]), .A2(in[192]), .ZN(n810) );
  AND2_X1 U153bar ( .A1(inbar[200]), .A2(inbar[192]), .ZN(n810bar) );
  OR2_X1 U154 ( .A1(n808), .A2(n807), .ZN(n816) );
  AND2_X1 U154bar ( .A1(n808bar), .A2(n807bar), .ZN(n816bar) );
  OR2_X1 U155 ( .A1(n806), .A2(n805), .ZN(n807) );
  AND2_X1 U155bar ( .A1(n806bar), .A2(n805bar), .ZN(n807bar) );
  OR2_X1 U156 ( .A1(in[225]), .A2(in[207]), .ZN(n805) );
  AND2_X1 U156bar ( .A1(inbar[225]), .A2(inbar[207]), .ZN(n805bar) );
  OR2_X1 U157 ( .A1(in[98]), .A2(in[226]), .ZN(n806) );
  AND2_X1 U157bar ( .A1(inbar[98]), .A2(inbar[226]), .ZN(n806bar) );
  OR2_X1 U158 ( .A1(n804), .A2(n803), .ZN(n808) );
  AND2_X1 U158bar ( .A1(n804bar), .A2(n803bar), .ZN(n808bar) );
  OR2_X1 U159 ( .A1(in_20), .A2(in_16), .ZN(n803) );
  AND2_X1 U159bar ( .A1(in_20bar), .A2(in_16bar), .ZN(n803bar) );
  OR2_X1 U160 ( .A1(in_55), .A2(in_45), .ZN(n804) );
  AND2_X1 U160bar ( .A1(in_55bar), .A2(in_45bar), .ZN(n804bar) );
  OR2_X1 U161 ( .A1(n802), .A2(n801), .ZN(n824) );
  AND2_X1 U161bar ( .A1(n802bar), .A2(n801bar), .ZN(n824bar) );
  OR2_X1 U162 ( .A1(in[162]), .A2(in[149]), .ZN(n801) );
  AND2_X1 U162bar ( .A1(inbar[162]), .A2(inbar[149]), .ZN(n801bar) );
  OR2_X1 U163 ( .A1(in[163]), .A2(n800), .ZN(n802) );
  AND2_X1 U163bar ( .A1(inbar[163]), .A2(n800bar), .ZN(n802bar) );
  OR2_X1 U164 ( .A1(in[191]), .A2(in[189]), .ZN(n800) );
  AND2_X1 U164bar ( .A1(inbar[191]), .A2(inbar[189]), .ZN(n800bar) );
  OR2_X1 U165 ( .A1(n799), .A2(n798), .ZN(n826) );
  AND2_X1 U165bar ( .A1(n799bar), .A2(n798bar), .ZN(n826bar) );
  OR2_X1 U166 ( .A1(n797), .A2(n796), .ZN(n798) );
  AND2_X1 U166bar ( .A1(n797bar), .A2(n796bar), .ZN(n798bar) );
  OR2_X1 U167 ( .A1(in[212]), .A2(in[193]), .ZN(n796) );
  AND2_X1 U167bar ( .A1(inbar[212]), .A2(inbar[193]), .ZN(n796bar) );
  OR2_X1 U168 ( .A1(in[238]), .A2(n795), .ZN(n797) );
  AND2_X1 U168bar ( .A1(inbar[238]), .A2(n795bar), .ZN(n797bar) );
  OR2_X1 U169 ( .A1(in[88]), .A2(in[247]), .ZN(n795) );
  AND2_X1 U169bar ( .A1(inbar[88]), .A2(inbar[247]), .ZN(n795bar) );
  OR2_X1 U170 ( .A1(n794), .A2(n793), .ZN(n799) );
  AND2_X1 U170bar ( .A1(n794bar), .A2(n793bar), .ZN(n799bar) );
  OR2_X1 U171 ( .A1(in[94]), .A2(in[92]), .ZN(n793) );
  AND2_X1 U171bar ( .A1(inbar[94]), .A2(inbar[92]), .ZN(n793bar) );
  OR2_X1 U172 ( .A1(in_52), .A2(n792), .ZN(n794) );
  AND2_X1 U172bar ( .A1(in_52bar), .A2(n792bar), .ZN(n794bar) );
  OR2_X1 U173 ( .A1(in_70), .A2(in_67), .ZN(n792) );
  AND2_X1 U173bar ( .A1(in_70bar), .A2(in_67bar), .ZN(n792bar) );
  OR2_X1 U174 ( .A1(n791), .A2(n790), .ZN(out[2]) );
  AND2_X1 U174bar ( .A1(n791bar), .A2(n790bar), .ZN(outbar[2]) );
  OR2_X1 U175 ( .A1(n789), .A2(n788), .ZN(n790) );
  AND2_X1 U175bar ( .A1(n789bar), .A2(n788bar), .ZN(n790bar) );
  OR2_X1 U176 ( .A1(n787), .A2(n786), .ZN(n788) );
  AND2_X1 U176bar ( .A1(n787bar), .A2(n786bar), .ZN(n788bar) );
  OR2_X1 U177 ( .A1(n819), .A2(n785), .ZN(n786) );
  AND2_X1 U177bar ( .A1(n819bar), .A2(n785bar), .ZN(n786bar) );
  OR2_X1 U178 ( .A1(n784), .A2(n783), .ZN(n819) );
  AND2_X1 U178bar ( .A1(n784bar), .A2(n783bar), .ZN(n819bar) );
  OR2_X1 U179 ( .A1(n782), .A2(n781), .ZN(n783) );
  AND2_X1 U179bar ( .A1(n782bar), .A2(n781bar), .ZN(n783bar) );
  OR2_X1 U180 ( .A1(n780), .A2(n779), .ZN(n781) );
  AND2_X1 U180bar ( .A1(n780bar), .A2(n779bar), .ZN(n781bar) );
  OR2_X1 U181 ( .A1(n962), .A2(n778), .ZN(n779) );
  AND2_X1 U181bar ( .A1(n962bar), .A2(n778bar), .ZN(n779bar) );
  OR2_X1 U182 ( .A1(n777), .A2(n776), .ZN(n962) );
  AND2_X1 U182bar ( .A1(n777bar), .A2(n776bar), .ZN(n962bar) );
  OR2_X1 U183 ( .A1(n775), .A2(n774), .ZN(n776) );
  AND2_X1 U183bar ( .A1(n775bar), .A2(n774bar), .ZN(n776bar) );
  OR2_X1 U184 ( .A1(n773), .A2(n772), .ZN(n774) );
  AND2_X1 U184bar ( .A1(n773bar), .A2(n772bar), .ZN(n774bar) );
  OR2_X1 U185 ( .A1(in[131]), .A2(in[120]), .ZN(n772) );
  AND2_X1 U185bar ( .A1(inbar[131]), .A2(inbar[120]), .ZN(n772bar) );
  OR2_X1 U186 ( .A1(in[153]), .A2(in[147]), .ZN(n773) );
  AND2_X1 U186bar ( .A1(inbar[153]), .A2(inbar[147]), .ZN(n773bar) );
  OR2_X1 U187 ( .A1(n771), .A2(n770), .ZN(n775) );
  AND2_X1 U187bar ( .A1(n771bar), .A2(n770bar), .ZN(n775bar) );
  OR2_X1 U188 ( .A1(in[170]), .A2(in[156]), .ZN(n770) );
  AND2_X1 U188bar ( .A1(inbar[170]), .A2(inbar[156]), .ZN(n770bar) );
  OR2_X1 U189 ( .A1(in[223]), .A2(in[190]), .ZN(n771) );
  AND2_X1 U189bar ( .A1(inbar[223]), .A2(inbar[190]), .ZN(n771bar) );
  OR2_X1 U190 ( .A1(n769), .A2(n768), .ZN(n777) );
  AND2_X1 U190bar ( .A1(n769bar), .A2(n768bar), .ZN(n777bar) );
  OR2_X1 U191 ( .A1(n767), .A2(n766), .ZN(n768) );
  AND2_X1 U191bar ( .A1(n767bar), .A2(n766bar), .ZN(n768bar) );
  OR2_X1 U192 ( .A1(in[236]), .A2(in[230]), .ZN(n766) );
  AND2_X1 U192bar ( .A1(inbar[236]), .A2(inbar[230]), .ZN(n766bar) );
  OR2_X1 U193 ( .A1(in[85]), .A2(in[240]), .ZN(n767) );
  AND2_X1 U193bar ( .A1(inbar[85]), .A2(inbar[240]), .ZN(n767bar) );
  OR2_X1 U194 ( .A1(n765), .A2(n764), .ZN(n769) );
  AND2_X1 U194bar ( .A1(n765bar), .A2(n764bar), .ZN(n769bar) );
  OR2_X1 U195 ( .A1(in_12), .A2(in[90]), .ZN(n764) );
  AND2_X1 U195bar ( .A1(in_12bar), .A2(inbar[90]), .ZN(n764bar) );
  OR2_X1 U196 ( .A1(in_39), .A2(in_28), .ZN(n765) );
  AND2_X1 U196bar ( .A1(in_39bar), .A2(in_28bar), .ZN(n765bar) );
  OR2_X1 U197 ( .A1(in[109]), .A2(n763), .ZN(n780) );
  AND2_X1 U197bar ( .A1(inbar[109]), .A2(n763bar), .ZN(n780bar) );
  OR2_X1 U198 ( .A1(n762), .A2(n761), .ZN(n782) );
  AND2_X1 U198bar ( .A1(n762bar), .A2(n761bar), .ZN(n782bar) );
  OR2_X1 U199 ( .A1(in[138]), .A2(in[129]), .ZN(n761) );
  AND2_X1 U199bar ( .A1(inbar[138]), .A2(inbar[129]), .ZN(n761bar) );
  OR2_X1 U200 ( .A1(in[157]), .A2(n760), .ZN(n762) );
  AND2_X1 U200bar ( .A1(inbar[157]), .A2(n760bar), .ZN(n762bar) );
  OR2_X1 U201 ( .A1(in[182]), .A2(in[167]), .ZN(n760) );
  AND2_X1 U201bar ( .A1(inbar[182]), .A2(inbar[167]), .ZN(n760bar) );
  OR2_X1 U202 ( .A1(n759), .A2(n758), .ZN(n784) );
  AND2_X1 U202bar ( .A1(n759bar), .A2(n758bar), .ZN(n784bar) );
  OR2_X1 U203 ( .A1(n757), .A2(n756), .ZN(n758) );
  AND2_X1 U203bar ( .A1(n757bar), .A2(n756bar), .ZN(n758bar) );
  OR2_X1 U204 ( .A1(in[195]), .A2(in[184]), .ZN(n756) );
  AND2_X1 U204bar ( .A1(inbar[195]), .A2(inbar[184]), .ZN(n756bar) );
  OR2_X1 U205 ( .A1(in[196]), .A2(n755), .ZN(n757) );
  AND2_X1 U205bar ( .A1(inbar[196]), .A2(n755bar), .ZN(n757bar) );
  OR2_X1 U206 ( .A1(in[215]), .A2(in[209]), .ZN(n755) );
  AND2_X1 U206bar ( .A1(inbar[215]), .A2(inbar[209]), .ZN(n755bar) );
  OR2_X1 U207 ( .A1(n754), .A2(n753), .ZN(n759) );
  AND2_X1 U207bar ( .A1(n754bar), .A2(n753bar), .ZN(n759bar) );
  OR2_X1 U208 ( .A1(in[93]), .A2(in[233]), .ZN(n753) );
  AND2_X1 U208bar ( .A1(inbar[93]), .A2(inbar[233]), .ZN(n753bar) );
  OR2_X1 U209 ( .A1(in_1), .A2(n752), .ZN(n754) );
  AND2_X1 U209bar ( .A1(in_1bar), .A2(n752bar), .ZN(n754bar) );
  OR2_X1 U210 ( .A1(in_69), .A2(in_66), .ZN(n752) );
  AND2_X1 U210bar ( .A1(in_69bar), .A2(in_66bar), .ZN(n752bar) );
  OR2_X1 U211 ( .A1(n966), .A2(n751), .ZN(n787) );
  AND2_X1 U211bar ( .A1(n966bar), .A2(n751bar), .ZN(n787bar) );
  OR2_X1 U212 ( .A1(in[134]), .A2(n750), .ZN(n751) );
  AND2_X1 U212bar ( .A1(inbar[134]), .A2(n750bar), .ZN(n751bar) );
  OR2_X1 U213 ( .A1(n749), .A2(n748), .ZN(n966) );
  AND2_X1 U213bar ( .A1(n749bar), .A2(n748bar), .ZN(n966bar) );
  OR2_X1 U214 ( .A1(n747), .A2(n746), .ZN(n748) );
  AND2_X1 U214bar ( .A1(n747bar), .A2(n746bar), .ZN(n748bar) );
  OR2_X1 U215 ( .A1(n745), .A2(n744), .ZN(n746) );
  AND2_X1 U215bar ( .A1(n745bar), .A2(n744bar), .ZN(n746bar) );
  OR2_X1 U216 ( .A1(in[136]), .A2(in[121]), .ZN(n744) );
  AND2_X1 U216bar ( .A1(inbar[136]), .A2(inbar[121]), .ZN(n744bar) );
  OR2_X1 U217 ( .A1(in[186]), .A2(in[174]), .ZN(n745) );
  AND2_X1 U217bar ( .A1(inbar[186]), .A2(inbar[174]), .ZN(n745bar) );
  OR2_X1 U218 ( .A1(n743), .A2(n742), .ZN(n747) );
  AND2_X1 U218bar ( .A1(n743bar), .A2(n742bar), .ZN(n747bar) );
  OR2_X1 U219 ( .A1(in[198]), .A2(in[197]), .ZN(n742) );
  AND2_X1 U219bar ( .A1(inbar[198]), .A2(inbar[197]), .ZN(n742bar) );
  OR2_X1 U220 ( .A1(in[214]), .A2(in[199]), .ZN(n743) );
  AND2_X1 U220bar ( .A1(inbar[214]), .A2(inbar[199]), .ZN(n743bar) );
  OR2_X1 U221 ( .A1(n741), .A2(n740), .ZN(n749) );
  AND2_X1 U221bar ( .A1(n741bar), .A2(n740bar), .ZN(n749bar) );
  OR2_X1 U222 ( .A1(n739), .A2(n738), .ZN(n740) );
  AND2_X1 U222bar ( .A1(n739bar), .A2(n738bar), .ZN(n740bar) );
  OR2_X1 U223 ( .A1(in[231]), .A2(in[220]), .ZN(n738) );
  AND2_X1 U223bar ( .A1(inbar[231]), .A2(inbar[220]), .ZN(n738bar) );
  OR2_X1 U224 ( .A1(in_25), .A2(in[245]), .ZN(n739) );
  AND2_X1 U224bar ( .A1(in_25bar), .A2(inbar[245]), .ZN(n739bar) );
  OR2_X1 U225 ( .A1(n737), .A2(n736), .ZN(n741) );
  AND2_X1 U225bar ( .A1(n737bar), .A2(n736bar), .ZN(n741bar) );
  OR2_X1 U226 ( .A1(in_53), .A2(in_29), .ZN(n736) );
  AND2_X1 U226bar ( .A1(in_53bar), .A2(in_29bar), .ZN(n736bar) );
  OR2_X1 U227 ( .A1(in_79), .A2(in_74), .ZN(n737) );
  AND2_X1 U227bar ( .A1(in_79bar), .A2(in_74bar), .ZN(n737bar) );
  OR2_X1 U228 ( .A1(n735), .A2(n734), .ZN(n789) );
  AND2_X1 U228bar ( .A1(n735bar), .A2(n734bar), .ZN(n789bar) );
  OR2_X1 U229 ( .A1(in[152]), .A2(in[140]), .ZN(n734) );
  AND2_X1 U229bar ( .A1(inbar[152]), .A2(inbar[140]), .ZN(n734bar) );
  OR2_X1 U230 ( .A1(in[155]), .A2(n733), .ZN(n735) );
  AND2_X1 U230bar ( .A1(inbar[155]), .A2(n733bar), .ZN(n735bar) );
  OR2_X1 U231 ( .A1(in[166]), .A2(in[165]), .ZN(n733) );
  AND2_X1 U231bar ( .A1(inbar[166]), .A2(inbar[165]), .ZN(n733bar) );
  OR2_X1 U232 ( .A1(n732), .A2(n731), .ZN(n791) );
  AND2_X1 U232bar ( .A1(n732bar), .A2(n731bar), .ZN(n791bar) );
  OR2_X1 U233 ( .A1(n730), .A2(n729), .ZN(n731) );
  AND2_X1 U233bar ( .A1(n730bar), .A2(n729bar), .ZN(n731bar) );
  OR2_X1 U234 ( .A1(in[202]), .A2(in[185]), .ZN(n729) );
  AND2_X1 U234bar ( .A1(inbar[202]), .A2(inbar[185]), .ZN(n729bar) );
  OR2_X1 U235 ( .A1(in[211]), .A2(n728), .ZN(n730) );
  AND2_X1 U235bar ( .A1(inbar[211]), .A2(n728bar), .ZN(n730bar) );
  OR2_X1 U236 ( .A1(in[255]), .A2(in[253]), .ZN(n728) );
  AND2_X1 U236bar ( .A1(inbar[255]), .A2(inbar[253]), .ZN(n728bar) );
  OR2_X1 U237 ( .A1(n727), .A2(n726), .ZN(n732) );
  AND2_X1 U237bar ( .A1(n727bar), .A2(n726bar), .ZN(n732bar) );
  OR2_X1 U238 ( .A1(in_35), .A2(in_15), .ZN(n726) );
  AND2_X1 U238bar ( .A1(in_35bar), .A2(in_15bar), .ZN(n726bar) );
  OR2_X1 U239 ( .A1(in_36), .A2(n725), .ZN(n727) );
  AND2_X1 U239bar ( .A1(in_36bar), .A2(n725bar), .ZN(n727bar) );
  OR2_X1 U240 ( .A1(in_48), .A2(in_40), .ZN(n725) );
  AND2_X1 U240bar ( .A1(in_48bar), .A2(in_40bar), .ZN(n725bar) );
  OR2_X1 U241 ( .A1(n724), .A2(n723), .ZN(out[1]) );
  AND2_X1 U241bar ( .A1(n724bar), .A2(n723bar), .ZN(outbar[1]) );
  OR2_X1 U242 ( .A1(n722), .A2(n721), .ZN(n723) );
  AND2_X1 U242bar ( .A1(n722bar), .A2(n721bar), .ZN(n723bar) );
  OR2_X1 U243 ( .A1(n720), .A2(n719), .ZN(n721) );
  AND2_X1 U243bar ( .A1(n720bar), .A2(n719bar), .ZN(n721bar) );
  OR2_X1 U244 ( .A1(n921), .A2(n887), .ZN(n719) );
  AND2_X1 U244bar ( .A1(n921bar), .A2(n887bar), .ZN(n719bar) );
  OR2_X1 U245 ( .A1(n718), .A2(n717), .ZN(n887) );
  AND2_X1 U245bar ( .A1(n718bar), .A2(n717bar), .ZN(n887bar) );
  OR2_X1 U246 ( .A1(n716), .A2(n715), .ZN(n717) );
  AND2_X1 U246bar ( .A1(n716bar), .A2(n715bar), .ZN(n717bar) );
  OR2_X1 U247 ( .A1(n714), .A2(n713), .ZN(n715) );
  AND2_X1 U247bar ( .A1(n714bar), .A2(n713bar), .ZN(n715bar) );
  OR2_X1 U248 ( .A1(in[116]), .A2(in[110]), .ZN(n713) );
  AND2_X1 U248bar ( .A1(inbar[116]), .A2(inbar[110]), .ZN(n713bar) );
  OR2_X1 U249 ( .A1(in[133]), .A2(in[130]), .ZN(n714) );
  AND2_X1 U249bar ( .A1(inbar[133]), .A2(inbar[130]), .ZN(n714bar) );
  OR2_X1 U250 ( .A1(n712), .A2(n711), .ZN(n716) );
  AND2_X1 U250bar ( .A1(n712bar), .A2(n711bar), .ZN(n716bar) );
  OR2_X1 U251 ( .A1(in[203]), .A2(in[135]), .ZN(n711) );
  AND2_X1 U251bar ( .A1(inbar[203]), .A2(inbar[135]), .ZN(n711bar) );
  OR2_X1 U252 ( .A1(in[232]), .A2(in[223]), .ZN(n712) );
  AND2_X1 U252bar ( .A1(inbar[232]), .A2(inbar[223]), .ZN(n712bar) );
  OR2_X1 U253 ( .A1(n710), .A2(n709), .ZN(n718) );
  AND2_X1 U253bar ( .A1(n710bar), .A2(n709bar), .ZN(n718bar) );
  OR2_X1 U254 ( .A1(n708), .A2(n707), .ZN(n709) );
  AND2_X1 U254bar ( .A1(n708bar), .A2(n707bar), .ZN(n709bar) );
  OR2_X1 U255 ( .A1(in[255]), .A2(in[233]), .ZN(n707) );
  AND2_X1 U255bar ( .A1(inbar[255]), .A2(inbar[233]), .ZN(n707bar) );
  OR2_X1 U256 ( .A1(in_53), .A2(in_34), .ZN(n708) );
  AND2_X1 U256bar ( .A1(in_53bar), .A2(in_34bar), .ZN(n708bar) );
  OR2_X1 U257 ( .A1(n706), .A2(n705), .ZN(n710) );
  AND2_X1 U257bar ( .A1(n706bar), .A2(n705bar), .ZN(n710bar) );
  OR2_X1 U258 ( .A1(in_57), .A2(in_55), .ZN(n705) );
  AND2_X1 U258bar ( .A1(in_57bar), .A2(in_55bar), .ZN(n705bar) );
  OR2_X1 U259 ( .A1(in_68), .A2(in_67), .ZN(n706) );
  AND2_X1 U259bar ( .A1(in_68bar), .A2(in_67bar), .ZN(n706bar) );
  OR2_X1 U260 ( .A1(n704), .A2(n703), .ZN(n921) );
  AND2_X1 U260bar ( .A1(n704bar), .A2(n703bar), .ZN(n921bar) );
  OR2_X1 U261 ( .A1(n702), .A2(n701), .ZN(n703) );
  AND2_X1 U261bar ( .A1(n702bar), .A2(n701bar), .ZN(n703bar) );
  OR2_X1 U262 ( .A1(n700), .A2(n699), .ZN(n701) );
  AND2_X1 U262bar ( .A1(n700bar), .A2(n699bar), .ZN(n701bar) );
  OR2_X1 U263 ( .A1(n944), .A2(n872), .ZN(n699) );
  AND2_X1 U263bar ( .A1(n944bar), .A2(n872bar), .ZN(n699bar) );
  OR2_X1 U264 ( .A1(n698), .A2(n697), .ZN(n872) );
  AND2_X1 U264bar ( .A1(n698bar), .A2(n697bar), .ZN(n872bar) );
  OR2_X1 U265 ( .A1(n696), .A2(n695), .ZN(n697) );
  AND2_X1 U265bar ( .A1(n696bar), .A2(n695bar), .ZN(n697bar) );
  OR2_X1 U266 ( .A1(n694), .A2(n693), .ZN(n695) );
  AND2_X1 U266bar ( .A1(n694bar), .A2(n693bar), .ZN(n695bar) );
  OR2_X1 U267 ( .A1(in[121]), .A2(in[102]), .ZN(n693) );
  AND2_X1 U267bar ( .A1(inbar[121]), .A2(inbar[102]), .ZN(n693bar) );
  OR2_X1 U268 ( .A1(in[162]), .A2(in[161]), .ZN(n694) );
  AND2_X1 U268bar ( .A1(inbar[162]), .A2(inbar[161]), .ZN(n694bar) );
  OR2_X1 U269 ( .A1(n692), .A2(n691), .ZN(n696) );
  AND2_X1 U269bar ( .A1(n692bar), .A2(n691bar), .ZN(n696bar) );
  OR2_X1 U270 ( .A1(in[192]), .A2(in[178]), .ZN(n691) );
  AND2_X1 U270bar ( .A1(inbar[192]), .A2(inbar[178]), .ZN(n691bar) );
  OR2_X1 U271 ( .A1(in[244]), .A2(in[209]), .ZN(n692) );
  AND2_X1 U271bar ( .A1(inbar[244]), .A2(inbar[209]), .ZN(n692bar) );
  OR2_X1 U272 ( .A1(n690), .A2(n689), .ZN(n698) );
  AND2_X1 U272bar ( .A1(n690bar), .A2(n689bar), .ZN(n698bar) );
  OR2_X1 U273 ( .A1(n688), .A2(n687), .ZN(n689) );
  AND2_X1 U273bar ( .A1(n688bar), .A2(n687bar), .ZN(n689bar) );
  OR2_X1 U274 ( .A1(in[90]), .A2(in[254]), .ZN(n687) );
  AND2_X1 U274bar ( .A1(inbar[90]), .A2(inbar[254]), .ZN(n687bar) );
  OR2_X1 U275 ( .A1(in_36), .A2(in_32), .ZN(n688) );
  AND2_X1 U275bar ( .A1(in_36bar), .A2(in_32bar), .ZN(n688bar) );
  OR2_X1 U276 ( .A1(n686), .A2(n685), .ZN(n690) );
  AND2_X1 U276bar ( .A1(n686bar), .A2(n685bar), .ZN(n690bar) );
  OR2_X1 U277 ( .A1(in_62), .A2(in_37), .ZN(n685) );
  AND2_X1 U277bar ( .A1(in_62bar), .A2(in_37bar), .ZN(n685bar) );
  OR2_X1 U278 ( .A1(in_75), .A2(in_73), .ZN(n686) );
  AND2_X1 U278bar ( .A1(in_75bar), .A2(in_73bar), .ZN(n686bar) );
  OR2_X1 U279 ( .A1(n684), .A2(n683), .ZN(n944) );
  AND2_X1 U279bar ( .A1(n684bar), .A2(n683bar), .ZN(n944bar) );
  OR2_X1 U280 ( .A1(n682), .A2(n681), .ZN(n683) );
  AND2_X1 U280bar ( .A1(n682bar), .A2(n681bar), .ZN(n683bar) );
  OR2_X1 U281 ( .A1(n680), .A2(n679), .ZN(n681) );
  AND2_X1 U281bar ( .A1(n680bar), .A2(n679bar), .ZN(n681bar) );
  OR2_X1 U282 ( .A1(in[171]), .A2(in[153]), .ZN(n679) );
  AND2_X1 U282bar ( .A1(inbar[171]), .A2(inbar[153]), .ZN(n679bar) );
  OR2_X1 U283 ( .A1(in[187]), .A2(in[176]), .ZN(n680) );
  AND2_X1 U283bar ( .A1(inbar[187]), .A2(inbar[176]), .ZN(n680bar) );
  OR2_X1 U284 ( .A1(n678), .A2(n677), .ZN(n682) );
  AND2_X1 U284bar ( .A1(n678bar), .A2(n677bar), .ZN(n682bar) );
  OR2_X1 U285 ( .A1(in[245]), .A2(in[211]), .ZN(n677) );
  AND2_X1 U285bar ( .A1(inbar[245]), .A2(inbar[211]), .ZN(n677bar) );
  OR2_X1 U286 ( .A1(in[97]), .A2(in[88]), .ZN(n678) );
  AND2_X1 U286bar ( .A1(inbar[97]), .A2(inbar[88]), .ZN(n678bar) );
  OR2_X1 U287 ( .A1(n676), .A2(n675), .ZN(n684) );
  AND2_X1 U287bar ( .A1(n676bar), .A2(n675bar), .ZN(n684bar) );
  OR2_X1 U288 ( .A1(n674), .A2(n673), .ZN(n675) );
  AND2_X1 U288bar ( .A1(n674bar), .A2(n673bar), .ZN(n675bar) );
  OR2_X1 U289 ( .A1(in_10), .A2(in_0), .ZN(n673) );
  AND2_X1 U289bar ( .A1(in_10bar), .A2(in_0bar), .ZN(n673bar) );
  OR2_X1 U290 ( .A1(in_59), .A2(in_5), .ZN(n674) );
  AND2_X1 U290bar ( .A1(in_59bar), .A2(in_5bar), .ZN(n674bar) );
  OR2_X1 U291 ( .A1(n672), .A2(n671), .ZN(n676) );
  AND2_X1 U291bar ( .A1(n672bar), .A2(n671bar), .ZN(n676bar) );
  OR2_X1 U292 ( .A1(in_60), .A2(in_6), .ZN(n671) );
  AND2_X1 U292bar ( .A1(in_60bar), .A2(in_6bar), .ZN(n671bar) );
  OR2_X1 U293 ( .A1(in_77), .A2(in_69), .ZN(n672) );
  AND2_X1 U293bar ( .A1(in_77bar), .A2(in_69bar), .ZN(n672bar) );
  OR2_X1 U294 ( .A1(in[113]), .A2(n864), .ZN(n700) );
  AND2_X1 U294bar ( .A1(inbar[113]), .A2(n864bar), .ZN(n700bar) );
  OR2_X1 U295 ( .A1(n670), .A2(n669), .ZN(n864) );
  AND2_X1 U295bar ( .A1(n670bar), .A2(n669bar), .ZN(n864bar) );
  OR2_X1 U296 ( .A1(n668), .A2(n667), .ZN(n669) );
  AND2_X1 U296bar ( .A1(n668bar), .A2(n667bar), .ZN(n669bar) );
  OR2_X1 U297 ( .A1(n666), .A2(n665), .ZN(n667) );
  AND2_X1 U297bar ( .A1(n666bar), .A2(n665bar), .ZN(n667bar) );
  OR2_X1 U298 ( .A1(in[125]), .A2(in[107]), .ZN(n665) );
  AND2_X1 U298bar ( .A1(inbar[125]), .A2(inbar[107]), .ZN(n665bar) );
  OR2_X1 U299 ( .A1(in[138]), .A2(in[126]), .ZN(n666) );
  AND2_X1 U299bar ( .A1(inbar[138]), .A2(inbar[126]), .ZN(n666bar) );
  OR2_X1 U300 ( .A1(n664), .A2(n663), .ZN(n668) );
  AND2_X1 U300bar ( .A1(n664bar), .A2(n663bar), .ZN(n668bar) );
  OR2_X1 U301 ( .A1(in[189]), .A2(in[143]), .ZN(n663) );
  AND2_X1 U301bar ( .A1(inbar[189]), .A2(inbar[143]), .ZN(n663bar) );
  OR2_X1 U302 ( .A1(in[99]), .A2(in[214]), .ZN(n664) );
  AND2_X1 U302bar ( .A1(inbar[99]), .A2(inbar[214]), .ZN(n664bar) );
  OR2_X1 U303 ( .A1(n662), .A2(n661), .ZN(n670) );
  AND2_X1 U303bar ( .A1(n662bar), .A2(n661bar), .ZN(n670bar) );
  OR2_X1 U304 ( .A1(n660), .A2(n659), .ZN(n661) );
  AND2_X1 U304bar ( .A1(n660bar), .A2(n659bar), .ZN(n661bar) );
  OR2_X1 U305 ( .A1(in_15), .A2(in_12), .ZN(n659) );
  AND2_X1 U305bar ( .A1(in_15bar), .A2(in_12bar), .ZN(n659bar) );
  OR2_X1 U306 ( .A1(in_20), .A2(in_2), .ZN(n660) );
  AND2_X1 U306bar ( .A1(in_20bar), .A2(in_2bar), .ZN(n660bar) );
  OR2_X1 U307 ( .A1(n658), .A2(n657), .ZN(n662) );
  AND2_X1 U307bar ( .A1(n658bar), .A2(n657bar), .ZN(n662bar) );
  OR2_X1 U308 ( .A1(in_30), .A2(in_3), .ZN(n657) );
  AND2_X1 U308bar ( .A1(in_30bar), .A2(in_3bar), .ZN(n657bar) );
  OR2_X1 U309 ( .A1(in_4), .A2(in_38), .ZN(n658) );
  AND2_X1 U309bar ( .A1(in_4bar), .A2(in_38bar), .ZN(n658bar) );
  OR2_X1 U310 ( .A1(n656), .A2(n655), .ZN(n702) );
  AND2_X1 U310bar ( .A1(n656bar), .A2(n655bar), .ZN(n702bar) );
  OR2_X1 U311 ( .A1(in[148]), .A2(in[137]), .ZN(n655) );
  AND2_X1 U311bar ( .A1(inbar[148]), .A2(inbar[137]), .ZN(n655bar) );
  OR2_X1 U312 ( .A1(in[149]), .A2(n654), .ZN(n656) );
  AND2_X1 U312bar ( .A1(inbar[149]), .A2(n654bar), .ZN(n656bar) );
  OR2_X1 U313 ( .A1(in[195]), .A2(in[190]), .ZN(n654) );
  AND2_X1 U313bar ( .A1(inbar[195]), .A2(inbar[190]), .ZN(n654bar) );
  OR2_X1 U314 ( .A1(n653), .A2(n652), .ZN(n704) );
  AND2_X1 U314bar ( .A1(n653bar), .A2(n652bar), .ZN(n704bar) );
  OR2_X1 U315 ( .A1(n651), .A2(n650), .ZN(n652) );
  AND2_X1 U315bar ( .A1(n651bar), .A2(n650bar), .ZN(n652bar) );
  OR2_X1 U316 ( .A1(in[98]), .A2(in[197]), .ZN(n650) );
  AND2_X1 U316bar ( .A1(inbar[98]), .A2(inbar[197]), .ZN(n650bar) );
  OR2_X1 U317 ( .A1(in_11), .A2(n649), .ZN(n651) );
  AND2_X1 U317bar ( .A1(in_11bar), .A2(n649bar), .ZN(n651bar) );
  OR2_X1 U318 ( .A1(in_26), .A2(in_14), .ZN(n649) );
  AND2_X1 U318bar ( .A1(in_26bar), .A2(in_14bar), .ZN(n649bar) );
  OR2_X1 U319 ( .A1(n648), .A2(n647), .ZN(n653) );
  AND2_X1 U319bar ( .A1(n648bar), .A2(n647bar), .ZN(n653bar) );
  OR2_X1 U320 ( .A1(in_35), .A2(in_27), .ZN(n647) );
  AND2_X1 U320bar ( .A1(in_35bar), .A2(in_27bar), .ZN(n647bar) );
  OR2_X1 U321 ( .A1(in_50), .A2(n646), .ZN(n648) );
  AND2_X1 U321bar ( .A1(in_50bar), .A2(n646bar), .ZN(n648bar) );
  OR2_X1 U322 ( .A1(in_78), .A2(in_61), .ZN(n646) );
  AND2_X1 U322bar ( .A1(in_78bar), .A2(in_61bar), .ZN(n646bar) );
  OR2_X1 U323 ( .A1(n942), .A2(n645), .ZN(n720) );
  AND2_X1 U323bar ( .A1(n942bar), .A2(n645bar), .ZN(n720bar) );
  OR2_X1 U324 ( .A1(in[106]), .A2(n863), .ZN(n645) );
  AND2_X1 U324bar ( .A1(inbar[106]), .A2(n863bar), .ZN(n645bar) );
  OR2_X1 U325 ( .A1(n644), .A2(n643), .ZN(n863) );
  AND2_X1 U325bar ( .A1(n644bar), .A2(n643bar), .ZN(n863bar) );
  OR2_X1 U326 ( .A1(n642), .A2(n641), .ZN(n643) );
  AND2_X1 U326bar ( .A1(n642bar), .A2(n641bar), .ZN(n643bar) );
  OR2_X1 U327 ( .A1(n640), .A2(n639), .ZN(n641) );
  AND2_X1 U327bar ( .A1(n640bar), .A2(n639bar), .ZN(n641bar) );
  OR2_X1 U328 ( .A1(in[127]), .A2(in[122]), .ZN(n639) );
  AND2_X1 U328bar ( .A1(inbar[127]), .A2(inbar[122]), .ZN(n639bar) );
  OR2_X1 U329 ( .A1(in[156]), .A2(in[132]), .ZN(n640) );
  AND2_X1 U329bar ( .A1(inbar[156]), .A2(inbar[132]), .ZN(n640bar) );
  OR2_X1 U330 ( .A1(n638), .A2(n637), .ZN(n642) );
  AND2_X1 U330bar ( .A1(n638bar), .A2(n637bar), .ZN(n642bar) );
  OR2_X1 U331 ( .A1(in[159]), .A2(in[157]), .ZN(n637) );
  AND2_X1 U331bar ( .A1(inbar[159]), .A2(inbar[157]), .ZN(n637bar) );
  OR2_X1 U332 ( .A1(in[185]), .A2(in[169]), .ZN(n638) );
  AND2_X1 U332bar ( .A1(inbar[185]), .A2(inbar[169]), .ZN(n638bar) );
  OR2_X1 U333 ( .A1(n636), .A2(n635), .ZN(n644) );
  AND2_X1 U333bar ( .A1(n636bar), .A2(n635bar), .ZN(n644bar) );
  OR2_X1 U334 ( .A1(n634), .A2(n633), .ZN(n635) );
  AND2_X1 U334bar ( .A1(n634bar), .A2(n633bar), .ZN(n635bar) );
  OR2_X1 U335 ( .A1(in[239]), .A2(in[218]), .ZN(n633) );
  AND2_X1 U335bar ( .A1(inbar[239]), .A2(inbar[218]), .ZN(n633bar) );
  OR2_X1 U336 ( .A1(in_13), .A2(in[87]), .ZN(n634) );
  AND2_X1 U336bar ( .A1(in_13bar), .A2(inbar[87]), .ZN(n634bar) );
  OR2_X1 U337 ( .A1(n632), .A2(n631), .ZN(n636) );
  AND2_X1 U337bar ( .A1(n632bar), .A2(n631bar), .ZN(n636bar) );
  OR2_X1 U338 ( .A1(in_72), .A2(in_70), .ZN(n631) );
  AND2_X1 U338bar ( .A1(in_72bar), .A2(in_70bar), .ZN(n631bar) );
  OR2_X1 U339 ( .A1(in_80), .A2(in_74), .ZN(n632) );
  AND2_X1 U339bar ( .A1(in_80bar), .A2(in_74bar), .ZN(n632bar) );
  OR2_X1 U340 ( .A1(n630), .A2(n629), .ZN(n942) );
  AND2_X1 U340bar ( .A1(n630bar), .A2(n629bar), .ZN(n942bar) );
  OR2_X1 U341 ( .A1(n628), .A2(n627), .ZN(n629) );
  AND2_X1 U341bar ( .A1(n628bar), .A2(n627bar), .ZN(n629bar) );
  OR2_X1 U342 ( .A1(n626), .A2(n625), .ZN(n627) );
  AND2_X1 U342bar ( .A1(n626bar), .A2(n625bar), .ZN(n627bar) );
  OR2_X1 U343 ( .A1(in[146]), .A2(in[100]), .ZN(n625) );
  AND2_X1 U343bar ( .A1(inbar[146]), .A2(inbar[100]), .ZN(n625bar) );
  OR2_X1 U344 ( .A1(in[168]), .A2(in[152]), .ZN(n626) );
  AND2_X1 U344bar ( .A1(inbar[168]), .A2(inbar[152]), .ZN(n626bar) );
  OR2_X1 U345 ( .A1(n624), .A2(n623), .ZN(n628) );
  AND2_X1 U345bar ( .A1(n624bar), .A2(n623bar), .ZN(n628bar) );
  OR2_X1 U346 ( .A1(in[199]), .A2(in[182]), .ZN(n623) );
  AND2_X1 U346bar ( .A1(inbar[199]), .A2(inbar[182]), .ZN(n623bar) );
  OR2_X1 U347 ( .A1(in[236]), .A2(in[204]), .ZN(n624) );
  AND2_X1 U347bar ( .A1(inbar[236]), .A2(inbar[204]), .ZN(n624bar) );
  OR2_X1 U348 ( .A1(n622), .A2(n621), .ZN(n630) );
  AND2_X1 U348bar ( .A1(n622bar), .A2(n621bar), .ZN(n630bar) );
  OR2_X1 U349 ( .A1(n620), .A2(n619), .ZN(n621) );
  AND2_X1 U349bar ( .A1(n620bar), .A2(n619bar), .ZN(n621bar) );
  OR2_X1 U350 ( .A1(in[89]), .A2(in[246]), .ZN(n619) );
  AND2_X1 U350bar ( .A1(inbar[89]), .A2(inbar[246]), .ZN(n619bar) );
  OR2_X1 U351 ( .A1(in[95]), .A2(in[92]), .ZN(n620) );
  AND2_X1 U351bar ( .A1(inbar[95]), .A2(inbar[92]), .ZN(n620bar) );
  OR2_X1 U352 ( .A1(n618), .A2(n617), .ZN(n622) );
  AND2_X1 U352bar ( .A1(n618bar), .A2(n617bar), .ZN(n622bar) );
  OR2_X1 U353 ( .A1(in_22), .A2(in_16), .ZN(n617) );
  AND2_X1 U353bar ( .A1(in_22bar), .A2(in_16bar), .ZN(n617bar) );
  OR2_X1 U354 ( .A1(in_51), .A2(in_49), .ZN(n618) );
  AND2_X1 U354bar ( .A1(in_51bar), .A2(in_49bar), .ZN(n618bar) );
  OR2_X1 U355 ( .A1(n616), .A2(n615), .ZN(n722) );
  AND2_X1 U355bar ( .A1(n616bar), .A2(n615bar), .ZN(n722bar) );
  OR2_X1 U356 ( .A1(in[158]), .A2(in[115]), .ZN(n615) );
  AND2_X1 U356bar ( .A1(inbar[158]), .A2(inbar[115]), .ZN(n615bar) );
  OR2_X1 U357 ( .A1(in[163]), .A2(n614), .ZN(n616) );
  AND2_X1 U357bar ( .A1(inbar[163]), .A2(n614bar), .ZN(n616bar) );
  OR2_X1 U358 ( .A1(in[206]), .A2(in[165]), .ZN(n614) );
  AND2_X1 U358bar ( .A1(inbar[206]), .A2(inbar[165]), .ZN(n614bar) );
  OR2_X1 U359 ( .A1(n613), .A2(n612), .ZN(n724) );
  AND2_X1 U359bar ( .A1(n613bar), .A2(n612bar), .ZN(n724bar) );
  OR2_X1 U360 ( .A1(n611), .A2(n610), .ZN(n612) );
  AND2_X1 U360bar ( .A1(n611bar), .A2(n610bar), .ZN(n612bar) );
  OR2_X1 U361 ( .A1(in[213]), .A2(in[207]), .ZN(n610) );
  AND2_X1 U361bar ( .A1(inbar[213]), .A2(inbar[207]), .ZN(n610bar) );
  OR2_X1 U362 ( .A1(in[215]), .A2(n609), .ZN(n611) );
  AND2_X1 U362bar ( .A1(inbar[215]), .A2(n609bar), .ZN(n611bar) );
  OR2_X1 U363 ( .A1(in[230]), .A2(in[220]), .ZN(n609) );
  AND2_X1 U363bar ( .A1(inbar[230]), .A2(inbar[220]), .ZN(n609bar) );
  OR2_X1 U364 ( .A1(n608), .A2(n607), .ZN(n613) );
  AND2_X1 U364bar ( .A1(n608bar), .A2(n607bar), .ZN(n613bar) );
  OR2_X1 U365 ( .A1(in[251]), .A2(in[234]), .ZN(n607) );
  AND2_X1 U365bar ( .A1(inbar[251]), .A2(inbar[234]), .ZN(n607bar) );
  OR2_X1 U366 ( .A1(in_17), .A2(n606), .ZN(n608) );
  AND2_X1 U366bar ( .A1(in_17bar), .A2(n606bar), .ZN(n608bar) );
  OR2_X1 U367 ( .A1(in_65), .A2(in_56), .ZN(n606) );
  AND2_X1 U367bar ( .A1(in_65bar), .A2(in_56bar), .ZN(n606bar) );
  OR2_X1 U368 ( .A1(n605), .A2(n604), .ZN(out[0]) );
  AND2_X1 U368bar ( .A1(n605bar), .A2(n604bar), .ZN(outbar[0]) );
  OR2_X1 U369 ( .A1(n603), .A2(n602), .ZN(n604) );
  AND2_X1 U369bar ( .A1(n603bar), .A2(n602bar), .ZN(n604bar) );
  OR2_X1 U370 ( .A1(n601), .A2(n600), .ZN(n602) );
  AND2_X1 U370bar ( .A1(n601bar), .A2(n600bar), .ZN(n602bar) );
  OR2_X1 U371 ( .A1(n820), .A2(n785), .ZN(n600) );
  AND2_X1 U371bar ( .A1(n820bar), .A2(n785bar), .ZN(n600bar) );
  OR2_X1 U372 ( .A1(n599), .A2(n598), .ZN(n785) );
  AND2_X1 U372bar ( .A1(n599bar), .A2(n598bar), .ZN(n785bar) );
  OR2_X1 U373 ( .A1(n597), .A2(n596), .ZN(n598) );
  AND2_X1 U373bar ( .A1(n597bar), .A2(n596bar), .ZN(n598bar) );
  OR2_X1 U374 ( .A1(n595), .A2(n594), .ZN(n596) );
  AND2_X1 U374bar ( .A1(n595bar), .A2(n594bar), .ZN(n596bar) );
  OR2_X1 U375 ( .A1(in[135]), .A2(in[104]), .ZN(n594) );
  AND2_X1 U375bar ( .A1(inbar[135]), .A2(inbar[104]), .ZN(n594bar) );
  OR2_X1 U376 ( .A1(in[188]), .A2(in[178]), .ZN(n595) );
  AND2_X1 U376bar ( .A1(inbar[188]), .A2(inbar[178]), .ZN(n595bar) );
  OR2_X1 U377 ( .A1(n593), .A2(n592), .ZN(n597) );
  AND2_X1 U377bar ( .A1(n593bar), .A2(n592bar), .ZN(n597bar) );
  OR2_X1 U378 ( .A1(in[217]), .A2(in[194]), .ZN(n592) );
  AND2_X1 U378bar ( .A1(inbar[217]), .A2(inbar[194]), .ZN(n592bar) );
  OR2_X1 U379 ( .A1(in[237]), .A2(in[218]), .ZN(n593) );
  AND2_X1 U379bar ( .A1(inbar[237]), .A2(inbar[218]), .ZN(n593bar) );
  OR2_X1 U380 ( .A1(n591), .A2(n590), .ZN(n599) );
  AND2_X1 U380bar ( .A1(n591bar), .A2(n590bar), .ZN(n599bar) );
  OR2_X1 U381 ( .A1(n589), .A2(n588), .ZN(n590) );
  AND2_X1 U381bar ( .A1(n589bar), .A2(n588bar), .ZN(n590bar) );
  OR2_X1 U382 ( .A1(in_2), .A2(in_10), .ZN(n588) );
  AND2_X1 U382bar ( .A1(in_2bar), .A2(in_10bar), .ZN(n588bar) );
  OR2_X1 U383 ( .A1(in_47), .A2(in_22), .ZN(n589) );
  AND2_X1 U383bar ( .A1(in_47bar), .A2(in_22bar), .ZN(n589bar) );
  OR2_X1 U384 ( .A1(n587), .A2(n586), .ZN(n591) );
  AND2_X1 U384bar ( .A1(n587bar), .A2(n586bar), .ZN(n591bar) );
  OR2_X1 U385 ( .A1(in_56), .A2(in_54), .ZN(n586) );
  AND2_X1 U385bar ( .A1(in_56bar), .A2(in_54bar), .ZN(n586bar) );
  OR2_X1 U386 ( .A1(in_63), .A2(in_61), .ZN(n587) );
  AND2_X1 U386bar ( .A1(in_63bar), .A2(in_61bar), .ZN(n587bar) );
  OR2_X1 U387 ( .A1(n585), .A2(n584), .ZN(n820) );
  AND2_X1 U387bar ( .A1(n585bar), .A2(n584bar), .ZN(n820bar) );
  OR2_X1 U388 ( .A1(n583), .A2(n582), .ZN(n584) );
  AND2_X1 U388bar ( .A1(n583bar), .A2(n582bar), .ZN(n584bar) );
  OR2_X1 U389 ( .A1(n581), .A2(n580), .ZN(n582) );
  AND2_X1 U389bar ( .A1(n581bar), .A2(n580bar), .ZN(n582bar) );
  OR2_X1 U390 ( .A1(in[158]), .A2(in[142]), .ZN(n580) );
  AND2_X1 U390bar ( .A1(inbar[158]), .A2(inbar[142]), .ZN(n580bar) );
  OR2_X1 U391 ( .A1(in[175]), .A2(in[164]), .ZN(n581) );
  AND2_X1 U391bar ( .A1(inbar[175]), .A2(inbar[164]), .ZN(n581bar) );
  OR2_X1 U392 ( .A1(n579), .A2(n578), .ZN(n583) );
  AND2_X1 U392bar ( .A1(n579bar), .A2(n578bar), .ZN(n583bar) );
  OR2_X1 U393 ( .A1(in[228]), .A2(in[204]), .ZN(n578) );
  AND2_X1 U393bar ( .A1(inbar[228]), .A2(inbar[204]), .ZN(n578bar) );
  OR2_X1 U394 ( .A1(in[91]), .A2(in[87]), .ZN(n579) );
  AND2_X1 U394bar ( .A1(inbar[91]), .A2(inbar[87]), .ZN(n579bar) );
  OR2_X1 U395 ( .A1(n577), .A2(n576), .ZN(n585) );
  AND2_X1 U395bar ( .A1(n577bar), .A2(n576bar), .ZN(n585bar) );
  OR2_X1 U396 ( .A1(n575), .A2(n574), .ZN(n576) );
  AND2_X1 U396bar ( .A1(n575bar), .A2(n574bar), .ZN(n576bar) );
  OR2_X1 U397 ( .A1(in_21), .A2(in_11), .ZN(n574) );
  AND2_X1 U397bar ( .A1(in_21bar), .A2(in_11bar), .ZN(n574bar) );
  OR2_X1 U398 ( .A1(in_5), .A2(in_3), .ZN(n575) );
  AND2_X1 U398bar ( .A1(in_5bar), .A2(in_3bar), .ZN(n575bar) );
  OR2_X1 U399 ( .A1(n573), .A2(n572), .ZN(n577) );
  AND2_X1 U399bar ( .A1(n573bar), .A2(n572bar), .ZN(n577bar) );
  OR2_X1 U400 ( .A1(in_68), .A2(in_64), .ZN(n572) );
  AND2_X1 U400bar ( .A1(in_68bar), .A2(in_64bar), .ZN(n572bar) );
  OR2_X1 U401 ( .A1(in_76), .A2(in_73), .ZN(n573) );
  AND2_X1 U401bar ( .A1(in_76bar), .A2(in_73bar), .ZN(n573bar) );
  OR2_X1 U402 ( .A1(n778), .A2(n571), .ZN(n601) );
  AND2_X1 U402bar ( .A1(n778bar), .A2(n571bar), .ZN(n601bar) );
  OR2_X1 U403 ( .A1(in[100]), .A2(n965), .ZN(n571) );
  AND2_X1 U403bar ( .A1(inbar[100]), .A2(n965bar), .ZN(n571bar) );
  OR2_X1 U404 ( .A1(n570), .A2(n569), .ZN(n965) );
  AND2_X1 U404bar ( .A1(n570bar), .A2(n569bar), .ZN(n965bar) );
  OR2_X1 U405 ( .A1(n568), .A2(n567), .ZN(n569) );
  AND2_X1 U405bar ( .A1(n568bar), .A2(n567bar), .ZN(n569bar) );
  OR2_X1 U406 ( .A1(n566), .A2(n565), .ZN(n567) );
  AND2_X1 U406bar ( .A1(n566bar), .A2(n565bar), .ZN(n567bar) );
  OR2_X1 U407 ( .A1(n817), .A2(n750), .ZN(n565) );
  AND2_X1 U407bar ( .A1(n817bar), .A2(n750bar), .ZN(n565bar) );
  OR2_X1 U408 ( .A1(n564), .A2(n563), .ZN(n750) );
  AND2_X1 U408bar ( .A1(n564bar), .A2(n563bar), .ZN(n750bar) );
  OR2_X1 U409 ( .A1(n562), .A2(n561), .ZN(n563) );
  AND2_X1 U409bar ( .A1(n562bar), .A2(n561bar), .ZN(n563bar) );
  OR2_X1 U410 ( .A1(n560), .A2(n559), .ZN(n561) );
  AND2_X1 U410bar ( .A1(n560bar), .A2(n559bar), .ZN(n561bar) );
  OR2_X1 U411 ( .A1(in[119]), .A2(in[103]), .ZN(n559) );
  AND2_X1 U411bar ( .A1(inbar[119]), .A2(inbar[103]), .ZN(n559bar) );
  OR2_X1 U412 ( .A1(in[137]), .A2(in[133]), .ZN(n560) );
  AND2_X1 U412bar ( .A1(inbar[137]), .A2(inbar[133]), .ZN(n560bar) );
  OR2_X1 U413 ( .A1(n558), .A2(n557), .ZN(n562) );
  AND2_X1 U413bar ( .A1(n558bar), .A2(n557bar), .ZN(n562bar) );
  OR2_X1 U414 ( .A1(in[176]), .A2(in[173]), .ZN(n557) );
  AND2_X1 U414bar ( .A1(inbar[176]), .A2(inbar[173]), .ZN(n557bar) );
  OR2_X1 U415 ( .A1(in[210]), .A2(in[181]), .ZN(n558) );
  AND2_X1 U415bar ( .A1(inbar[210]), .A2(inbar[181]), .ZN(n558bar) );
  OR2_X1 U416 ( .A1(n556), .A2(n555), .ZN(n564) );
  AND2_X1 U416bar ( .A1(n556bar), .A2(n555bar), .ZN(n564bar) );
  OR2_X1 U417 ( .A1(n554), .A2(n553), .ZN(n555) );
  AND2_X1 U417bar ( .A1(n554bar), .A2(n553bar), .ZN(n555bar) );
  OR2_X1 U418 ( .A1(in_13), .A2(in[234]), .ZN(n553) );
  AND2_X1 U418bar ( .A1(in_13bar), .A2(inbar[234]), .ZN(n553bar) );
  OR2_X1 U419 ( .A1(in_38), .A2(in_32), .ZN(n554) );
  AND2_X1 U419bar ( .A1(in_38bar), .A2(in_32bar), .ZN(n554bar) );
  OR2_X1 U420 ( .A1(n552), .A2(n551), .ZN(n556) );
  AND2_X1 U420bar ( .A1(n552bar), .A2(n551bar), .ZN(n556bar) );
  OR2_X1 U421 ( .A1(in_42), .A2(in_41), .ZN(n551) );
  AND2_X1 U421bar ( .A1(in_42bar), .A2(in_41bar), .ZN(n551bar) );
  OR2_X1 U422 ( .A1(in_7), .A2(in_49), .ZN(n552) );
  AND2_X1 U422bar ( .A1(in_7bar), .A2(in_49bar), .ZN(n552bar) );
  OR2_X1 U423 ( .A1(n550), .A2(n549), .ZN(n817) );
  AND2_X1 U423bar ( .A1(n550bar), .A2(n549bar), .ZN(n817bar) );
  OR2_X1 U424 ( .A1(n548), .A2(n547), .ZN(n549) );
  AND2_X1 U424bar ( .A1(n548bar), .A2(n547bar), .ZN(n549bar) );
  OR2_X1 U425 ( .A1(n546), .A2(n545), .ZN(n547) );
  AND2_X1 U425bar ( .A1(n546bar), .A2(n545bar), .ZN(n547bar) );
  OR2_X1 U426 ( .A1(in[159]), .A2(in[105]), .ZN(n545) );
  AND2_X1 U426bar ( .A1(inbar[159]), .A2(inbar[105]), .ZN(n545bar) );
  OR2_X1 U427 ( .A1(in[206]), .A2(in[183]), .ZN(n546) );
  AND2_X1 U427bar ( .A1(inbar[206]), .A2(inbar[183]), .ZN(n546bar) );
  OR2_X1 U428 ( .A1(n544), .A2(n543), .ZN(n548) );
  AND2_X1 U428bar ( .A1(n544bar), .A2(n543bar), .ZN(n548bar) );
  OR2_X1 U429 ( .A1(in[229]), .A2(in[219]), .ZN(n543) );
  AND2_X1 U429bar ( .A1(inbar[229]), .A2(inbar[219]), .ZN(n543bar) );
  OR2_X1 U430 ( .A1(in[235]), .A2(in[232]), .ZN(n544) );
  AND2_X1 U430bar ( .A1(inbar[235]), .A2(inbar[232]), .ZN(n544bar) );
  OR2_X1 U431 ( .A1(n542), .A2(n541), .ZN(n550) );
  AND2_X1 U431bar ( .A1(n542bar), .A2(n541bar), .ZN(n550bar) );
  OR2_X1 U432 ( .A1(n540), .A2(n539), .ZN(n541) );
  AND2_X1 U432bar ( .A1(n540bar), .A2(n539bar), .ZN(n541bar) );
  OR2_X1 U433 ( .A1(in[249]), .A2(in[242]), .ZN(n539) );
  AND2_X1 U433bar ( .A1(inbar[249]), .A2(inbar[242]), .ZN(n539bar) );
  OR2_X1 U434 ( .A1(in[89]), .A2(in[254]), .ZN(n540) );
  AND2_X1 U434bar ( .A1(inbar[89]), .A2(inbar[254]), .ZN(n540bar) );
  OR2_X1 U435 ( .A1(n538), .A2(n537), .ZN(n542) );
  AND2_X1 U435bar ( .A1(n538bar), .A2(n537bar), .ZN(n542bar) );
  OR2_X1 U436 ( .A1(in_14), .A2(in[99]), .ZN(n537) );
  AND2_X1 U436bar ( .A1(in_14bar), .A2(inbar[99]), .ZN(n537bar) );
  OR2_X1 U437 ( .A1(in_60), .A2(in_18), .ZN(n538) );
  AND2_X1 U437bar ( .A1(in_60bar), .A2(in_18bar), .ZN(n538bar) );
  OR2_X1 U438 ( .A1(in[113]), .A2(n763), .ZN(n566) );
  AND2_X1 U438bar ( .A1(inbar[113]), .A2(n763bar), .ZN(n566bar) );
  OR2_X1 U439 ( .A1(n536), .A2(n535), .ZN(n763) );
  AND2_X1 U439bar ( .A1(n536bar), .A2(n535bar), .ZN(n763bar) );
  OR2_X1 U440 ( .A1(n534), .A2(n533), .ZN(n535) );
  AND2_X1 U440bar ( .A1(n534bar), .A2(n533bar), .ZN(n535bar) );
  OR2_X1 U441 ( .A1(n532), .A2(n531), .ZN(n533) );
  AND2_X1 U441bar ( .A1(n532bar), .A2(n531bar), .ZN(n533bar) );
  OR2_X1 U442 ( .A1(in[115]), .A2(in[110]), .ZN(n531) );
  AND2_X1 U442bar ( .A1(inbar[115]), .A2(inbar[110]), .ZN(n531bar) );
  OR2_X1 U443 ( .A1(in[125]), .A2(in[117]), .ZN(n532) );
  AND2_X1 U443bar ( .A1(inbar[125]), .A2(inbar[117]), .ZN(n532bar) );
  OR2_X1 U444 ( .A1(n530), .A2(n529), .ZN(n534) );
  AND2_X1 U444bar ( .A1(n530bar), .A2(n529bar), .ZN(n534bar) );
  OR2_X1 U445 ( .A1(in[180]), .A2(in[128]), .ZN(n529) );
  AND2_X1 U445bar ( .A1(inbar[180]), .A2(inbar[128]), .ZN(n529bar) );
  OR2_X1 U446 ( .A1(in[205]), .A2(in[201]), .ZN(n530) );
  AND2_X1 U446bar ( .A1(inbar[205]), .A2(inbar[201]), .ZN(n530bar) );
  OR2_X1 U447 ( .A1(n528), .A2(n527), .ZN(n536) );
  AND2_X1 U447bar ( .A1(n528bar), .A2(n527bar), .ZN(n536bar) );
  OR2_X1 U448 ( .A1(n526), .A2(n525), .ZN(n527) );
  AND2_X1 U448bar ( .A1(n526bar), .A2(n525bar), .ZN(n527bar) );
  OR2_X1 U449 ( .A1(in[244]), .A2(in[239]), .ZN(n525) );
  AND2_X1 U449bar ( .A1(inbar[244]), .A2(inbar[239]), .ZN(n525bar) );
  OR2_X1 U450 ( .A1(in[95]), .A2(in[83]), .ZN(n526) );
  AND2_X1 U450bar ( .A1(inbar[95]), .A2(inbar[83]), .ZN(n526bar) );
  OR2_X1 U451 ( .A1(n524), .A2(n523), .ZN(n528) );
  AND2_X1 U451bar ( .A1(n524bar), .A2(n523bar), .ZN(n528bar) );
  OR2_X1 U452 ( .A1(in_24), .A2(in[97]), .ZN(n523) );
  AND2_X1 U452bar ( .A1(in_24bar), .A2(inbar[97]), .ZN(n523bar) );
  OR2_X1 U453 ( .A1(in_33), .A2(in_27), .ZN(n524) );
  AND2_X1 U453bar ( .A1(in_33bar), .A2(in_27bar), .ZN(n524bar) );
  OR2_X1 U454 ( .A1(n522), .A2(n521), .ZN(n568) );
  AND2_X1 U454bar ( .A1(n522bar), .A2(n521bar), .ZN(n568bar) );
  OR2_X1 U455 ( .A1(in[145]), .A2(in[126]), .ZN(n521) );
  AND2_X1 U455bar ( .A1(inbar[145]), .A2(inbar[126]), .ZN(n521bar) );
  OR2_X1 U456 ( .A1(in[169]), .A2(n520), .ZN(n522) );
  AND2_X1 U456bar ( .A1(inbar[169]), .A2(n520bar), .ZN(n522bar) );
  OR2_X1 U457 ( .A1(in[221]), .A2(in[172]), .ZN(n520) );
  AND2_X1 U457bar ( .A1(inbar[221]), .A2(inbar[172]), .ZN(n520bar) );
  OR2_X1 U458 ( .A1(n519), .A2(n518), .ZN(n570) );
  AND2_X1 U458bar ( .A1(n519bar), .A2(n518bar), .ZN(n570bar) );
  OR2_X1 U459 ( .A1(n517), .A2(n516), .ZN(n518) );
  AND2_X1 U459bar ( .A1(n517bar), .A2(n516bar), .ZN(n518bar) );
  OR2_X1 U460 ( .A1(in[241]), .A2(in[224]), .ZN(n516) );
  AND2_X1 U460bar ( .A1(inbar[241]), .A2(inbar[224]), .ZN(n516bar) );
  OR2_X1 U461 ( .A1(in[86]), .A2(n515), .ZN(n517) );
  AND2_X1 U461bar ( .A1(inbar[86]), .A2(n515bar), .ZN(n517bar) );
  OR2_X1 U462 ( .A1(in_43), .A2(in_34), .ZN(n515) );
  AND2_X1 U462bar ( .A1(in_43bar), .A2(in_34bar), .ZN(n515bar) );
  OR2_X1 U463 ( .A1(n514), .A2(n513), .ZN(n519) );
  AND2_X1 U463bar ( .A1(n514bar), .A2(n513bar), .ZN(n519bar) );
  OR2_X1 U464 ( .A1(in_65), .A2(in_51), .ZN(n513) );
  AND2_X1 U464bar ( .A1(in_65bar), .A2(in_51bar), .ZN(n513bar) );
  OR2_X1 U465 ( .A1(in_75), .A2(n512), .ZN(n514) );
  AND2_X1 U465bar ( .A1(in_75bar), .A2(n512bar), .ZN(n514bar) );
  OR2_X1 U466 ( .A1(in_81), .A2(in_77), .ZN(n512) );
  AND2_X1 U466bar ( .A1(in_81bar), .A2(in_77bar), .ZN(n512bar) );
  OR2_X1 U467 ( .A1(n511), .A2(n510), .ZN(n778) );
  AND2_X1 U467bar ( .A1(n511bar), .A2(n510bar), .ZN(n778bar) );
  OR2_X1 U468 ( .A1(n509), .A2(n508), .ZN(n510) );
  AND2_X1 U468bar ( .A1(n509bar), .A2(n508bar), .ZN(n510bar) );
  OR2_X1 U469 ( .A1(n507), .A2(n506), .ZN(n508) );
  AND2_X1 U469bar ( .A1(n507bar), .A2(n506bar), .ZN(n508bar) );
  OR2_X1 U470 ( .A1(in[107]), .A2(in[101]), .ZN(n506) );
  AND2_X1 U470bar ( .A1(inbar[107]), .A2(inbar[101]), .ZN(n506bar) );
  OR2_X1 U471 ( .A1(in[139]), .A2(in[132]), .ZN(n507) );
  AND2_X1 U471bar ( .A1(inbar[139]), .A2(inbar[132]), .ZN(n507bar) );
  OR2_X1 U472 ( .A1(n505), .A2(n504), .ZN(n509) );
  AND2_X1 U472bar ( .A1(n505bar), .A2(n504bar), .ZN(n509bar) );
  OR2_X1 U473 ( .A1(in[146]), .A2(in[141]), .ZN(n504) );
  AND2_X1 U473bar ( .A1(inbar[146]), .A2(inbar[141]), .ZN(n504bar) );
  OR2_X1 U474 ( .A1(in[203]), .A2(in[179]), .ZN(n505) );
  AND2_X1 U474bar ( .A1(inbar[203]), .A2(inbar[179]), .ZN(n505bar) );
  OR2_X1 U475 ( .A1(n503), .A2(n502), .ZN(n511) );
  AND2_X1 U475bar ( .A1(n503bar), .A2(n502bar), .ZN(n511bar) );
  OR2_X1 U476 ( .A1(n501), .A2(n500), .ZN(n502) );
  AND2_X1 U476bar ( .A1(n501bar), .A2(n500bar), .ZN(n502bar) );
  OR2_X1 U477 ( .A1(in[243]), .A2(in[222]), .ZN(n500) );
  AND2_X1 U477bar ( .A1(inbar[243]), .A2(inbar[222]), .ZN(n500bar) );
  OR2_X1 U478 ( .A1(in[251]), .A2(in[250]), .ZN(n501) );
  AND2_X1 U478bar ( .A1(inbar[251]), .A2(inbar[250]), .ZN(n501bar) );
  OR2_X1 U479 ( .A1(n499), .A2(n498), .ZN(n503) );
  AND2_X1 U479bar ( .A1(n499bar), .A2(n498bar), .ZN(n503bar) );
  OR2_X1 U480 ( .A1(in_37), .A2(in_19), .ZN(n498) );
  AND2_X1 U480bar ( .A1(in_37bar), .A2(in_19bar), .ZN(n498bar) );
  OR2_X1 U481 ( .A1(in_78), .A2(in_6), .ZN(n499) );
  AND2_X1 U481bar ( .A1(in_78bar), .A2(in_6bar), .ZN(n499bar) );
  OR2_X1 U482 ( .A1(n497), .A2(n496), .ZN(n603) );
  AND2_X1 U482bar ( .A1(n497bar), .A2(n496bar), .ZN(n603bar) );
  OR2_X1 U483 ( .A1(in[112]), .A2(in[102]), .ZN(n496) );
  AND2_X1 U483bar ( .A1(inbar[112]), .A2(inbar[102]), .ZN(n496bar) );
  OR2_X1 U484 ( .A1(in[123]), .A2(n495), .ZN(n497) );
  AND2_X1 U484bar ( .A1(inbar[123]), .A2(n495bar), .ZN(n497bar) );
  OR2_X1 U485 ( .A1(in[143]), .A2(in[130]), .ZN(n495) );
  AND2_X1 U485bar ( .A1(inbar[143]), .A2(inbar[130]), .ZN(n495bar) );
  OR2_X1 U486 ( .A1(n494), .A2(n493), .ZN(n605) );
  AND2_X1 U486bar ( .A1(n494bar), .A2(n493bar), .ZN(n605bar) );
  OR2_X1 U487 ( .A1(n492), .A2(n491), .ZN(n493) );
  AND2_X1 U487bar ( .A1(n492bar), .A2(n491bar), .ZN(n493bar) );
  OR2_X1 U488 ( .A1(in[216]), .A2(in[213]), .ZN(n491) );
  AND2_X1 U488bar ( .A1(inbar[216]), .A2(inbar[213]), .ZN(n491bar) );
  OR2_X1 U489 ( .A1(in[227]), .A2(n490), .ZN(n492) );
  AND2_X1 U489bar ( .A1(inbar[227]), .A2(n490bar), .ZN(n492bar) );
  OR2_X1 U490 ( .A1(in_0), .A2(in[248]), .ZN(n490) );
  AND2_X1 U490bar ( .A1(in_0bar), .A2(inbar[248]), .ZN(n490bar) );
  OR2_X1 U491 ( .A1(n489), .A2(n488), .ZN(n494) );
  AND2_X1 U491bar ( .A1(n489bar), .A2(n488bar), .ZN(n494bar) );
  OR2_X1 U492 ( .A1(in_46), .A2(in_44), .ZN(n488) );
  AND2_X1 U492bar ( .A1(in_46bar), .A2(in_44bar), .ZN(n488bar) );
  OR2_X1 U493 ( .A1(in_50), .A2(n487), .ZN(n489) );
  AND2_X1 U493bar ( .A1(in_50bar), .A2(n487bar), .ZN(n489bar) );
  OR2_X1 U494 ( .A1(in_9), .A2(in_80), .ZN(n487) );
  AND2_X1 U494bar ( .A1(in_9bar), .A2(in_80bar), .ZN(n487bar) );
endmodule

module sBox_15 ( in, inbar, out, outbar );

  input wire [7:0] in;
  input wire [7:0] inbar;
//input_done

  output wire [7:0] out;
  output wire [7:0] outbar;
//output_done

  wire [255:0] decodeOut;
  wire [255:0] decodeOutbar;
//wire_done

  decode_15 dec ( .in(in), .inbar(inbar), .out(decodeOut), .outbar(decodeOutbar) );
  encode_15 enc ( .in(decodeOut), .inbar(decodeOutbar), .out(out), .outbar(outbar) );
endmodule

module s_box_Precharge ( in, inbar, out, outbar );

  input wire [127:0] in;
  input wire [127:0] inbar;
//input_done

  output [127:0] out;
  output [127:0] outbar;
//output_done

//wire_done

  sBox_15 s0 ( .in(in[127:120]), .inbar(inbar[127:120]), .out(out[127:120]), .outbar(outbar[127:120]) );
  sBox_14 s1 ( .in(in[119:112]), .inbar(inbar[119:112]), .out(out[119:112]), .outbar(outbar[119:112]) );
  sBox_13 s2 ( .in(in[111:104]), .inbar(inbar[111:104]), .out(out[111:104]), .outbar(outbar[111:104]) );
  sBox_12 s3 ( .in(in[103:96]), .inbar(inbar[103:96]), .out(out[103:96]), .outbar(outbar[103:96]) );
  sBox_11 s4 ( .in(in[95:88]), .inbar(inbar[95:88]), .out(out[95:88]), .outbar(outbar[95:88]) );
  sBox_10 s5 ( .in(in[87:80]), .inbar(inbar[87:80]), .out(out[87:80]), .outbar(outbar[87:80]) );
  sBox_9 s6 ( .in(in[79:72]), .inbar(inbar[79:72]), .out(out[79:72]), .outbar(outbar[79:72]) );
  sBox_8 s7 ( .in(in[71:64]), .inbar(inbar[71:64]), .out(out[71:64]), .outbar(outbar[71:64]) );
  sBox_7 s8 ( .in(in[63:56]), .inbar(inbar[63:56]), .out(out[63:56]), .outbar(outbar[63:56]) );
  sBox_6 s9 ( .in(in[55:48]), .inbar(inbar[55:48]), .out(out[55:48]), .outbar(outbar[55:48]) );
  sBox_5 s10 ( .in(in[47:40]), .inbar(inbar[47:40]), .out(out[47:40]), .outbar(outbar[47:40]) );
  sBox_4 s11 ( .in(in[39:32]), .inbar(inbar[39:32]), .out(out[39:32]), .outbar(outbar[39:32]) );
  sBox_3 s12 ( .in(in[31:24]), .inbar(inbar[31:24]), .out(out[31:24]), .outbar(outbar[31:24]) );
  sBox_2 s13 ( .in(in[23:16]), .inbar(inbar[23:16]), .out(out[23:16]), .outbar(outbar[23:16]) );
  sBox_1 s14 ( .in(in[15:8]), .inbar(inbar[15:8]), .out(out[15:8]), .outbar(outbar[15:8]) );
  sBox_0 s15 ( .in(in[7:0]), .inbar(inbar[7:0]), .out(out[7:0]), .outbar(outbar[7:0]) );
endmodule

//done
