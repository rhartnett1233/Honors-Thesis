
module mux128_0 ( a, b, sel, y );
  input [127:0] a;
  input [127:0] b;
  input sel;
  //input_done

  output [127:0] y;
  //output_done

  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n1, n258, n259, n260;
  //wire_done

  OR2_X1 U2 ( .A1(n2), .A2(n3), .ZN(y[9]) );
  AND2_X1 U3 ( .A1(sel), .A2(b[9]), .ZN(n3) );
  AND2_X1 U4 ( .A1(a[9]), .A2(n258), .ZN(n2) );
  OR2_X1 U5 ( .A1(n4), .A2(n5), .ZN(y[99]) );
  AND2_X1 U6 ( .A1(b[99]), .A2(sel), .ZN(n5) );
  AND2_X1 U7 ( .A1(a[99]), .A2(n258), .ZN(n4) );
  OR2_X1 U8 ( .A1(n6), .A2(n7), .ZN(y[98]) );
  AND2_X1 U9 ( .A1(b[98]), .A2(sel), .ZN(n7) );
  AND2_X1 U10 ( .A1(a[98]), .A2(n258), .ZN(n6) );
  OR2_X1 U11 ( .A1(n8), .A2(n9), .ZN(y[97]) );
  AND2_X1 U12 ( .A1(b[97]), .A2(sel), .ZN(n9) );
  AND2_X1 U13 ( .A1(a[97]), .A2(n258), .ZN(n8) );
  OR2_X1 U14 ( .A1(n10), .A2(n11), .ZN(y[96]) );
  AND2_X1 U15 ( .A1(b[96]), .A2(sel), .ZN(n11) );
  AND2_X1 U16 ( .A1(a[96]), .A2(n258), .ZN(n10) );
  OR2_X1 U17 ( .A1(n12), .A2(n13), .ZN(y[95]) );
  AND2_X1 U18 ( .A1(b[95]), .A2(sel), .ZN(n13) );
  AND2_X1 U19 ( .A1(a[95]), .A2(n258), .ZN(n12) );
  OR2_X1 U20 ( .A1(n14), .A2(n15), .ZN(y[94]) );
  AND2_X1 U21 ( .A1(b[94]), .A2(sel), .ZN(n15) );
  AND2_X1 U22 ( .A1(a[94]), .A2(n258), .ZN(n14) );
  OR2_X1 U23 ( .A1(n16), .A2(n17), .ZN(y[93]) );
  AND2_X1 U24 ( .A1(b[93]), .A2(sel), .ZN(n17) );
  AND2_X1 U25 ( .A1(a[93]), .A2(n258), .ZN(n16) );
  OR2_X1 U26 ( .A1(n18), .A2(n19), .ZN(y[92]) );
  AND2_X1 U27 ( .A1(b[92]), .A2(sel), .ZN(n19) );
  AND2_X1 U28 ( .A1(a[92]), .A2(n258), .ZN(n18) );
  OR2_X1 U29 ( .A1(n20), .A2(n21), .ZN(y[91]) );
  AND2_X1 U30 ( .A1(b[91]), .A2(sel), .ZN(n21) );
  AND2_X1 U31 ( .A1(a[91]), .A2(n258), .ZN(n20) );
  OR2_X1 U32 ( .A1(n22), .A2(n23), .ZN(y[90]) );
  AND2_X1 U33 ( .A1(b[90]), .A2(sel), .ZN(n23) );
  AND2_X1 U34 ( .A1(a[90]), .A2(n258), .ZN(n22) );
  OR2_X1 U35 ( .A1(n24), .A2(n25), .ZN(y[8]) );
  AND2_X1 U36 ( .A1(b[8]), .A2(sel), .ZN(n25) );
  AND2_X1 U37 ( .A1(a[8]), .A2(n260), .ZN(n24) );
  OR2_X1 U38 ( .A1(n26), .A2(n27), .ZN(y[89]) );
  AND2_X1 U39 ( .A1(b[89]), .A2(sel), .ZN(n27) );
  AND2_X1 U40 ( .A1(a[89]), .A2(n258), .ZN(n26) );
  OR2_X1 U41 ( .A1(n28), .A2(n29), .ZN(y[88]) );
  AND2_X1 U42 ( .A1(b[88]), .A2(sel), .ZN(n29) );
  AND2_X1 U43 ( .A1(a[88]), .A2(n1), .ZN(n28) );
  OR2_X1 U44 ( .A1(n30), .A2(n31), .ZN(y[87]) );
  AND2_X1 U45 ( .A1(b[87]), .A2(sel), .ZN(n31) );
  AND2_X1 U46 ( .A1(a[87]), .A2(n259), .ZN(n30) );
  OR2_X1 U47 ( .A1(n32), .A2(n33), .ZN(y[86]) );
  AND2_X1 U48 ( .A1(b[86]), .A2(sel), .ZN(n33) );
  AND2_X1 U49 ( .A1(a[86]), .A2(n260), .ZN(n32) );
  OR2_X1 U50 ( .A1(n34), .A2(n35), .ZN(y[85]) );
  AND2_X1 U51 ( .A1(b[85]), .A2(sel), .ZN(n35) );
  AND2_X1 U52 ( .A1(a[85]), .A2(n1), .ZN(n34) );
  OR2_X1 U53 ( .A1(n36), .A2(n37), .ZN(y[84]) );
  AND2_X1 U54 ( .A1(b[84]), .A2(sel), .ZN(n37) );
  AND2_X1 U55 ( .A1(a[84]), .A2(n258), .ZN(n36) );
  OR2_X1 U56 ( .A1(n38), .A2(n39), .ZN(y[83]) );
  AND2_X1 U57 ( .A1(b[83]), .A2(sel), .ZN(n39) );
  AND2_X1 U58 ( .A1(a[83]), .A2(n1), .ZN(n38) );
  OR2_X1 U59 ( .A1(n40), .A2(n41), .ZN(y[82]) );
  AND2_X1 U60 ( .A1(b[82]), .A2(sel), .ZN(n41) );
  AND2_X1 U61 ( .A1(a[82]), .A2(n259), .ZN(n40) );
  OR2_X1 U62 ( .A1(n42), .A2(n43), .ZN(y[81]) );
  AND2_X1 U63 ( .A1(b[81]), .A2(sel), .ZN(n43) );
  AND2_X1 U64 ( .A1(a[81]), .A2(n260), .ZN(n42) );
  OR2_X1 U65 ( .A1(n44), .A2(n45), .ZN(y[80]) );
  AND2_X1 U66 ( .A1(b[80]), .A2(sel), .ZN(n45) );
  AND2_X1 U67 ( .A1(a[80]), .A2(n260), .ZN(n44) );
  OR2_X1 U68 ( .A1(n46), .A2(n47), .ZN(y[7]) );
  AND2_X1 U69 ( .A1(b[7]), .A2(sel), .ZN(n47) );
  AND2_X1 U70 ( .A1(a[7]), .A2(n258), .ZN(n46) );
  OR2_X1 U71 ( .A1(n48), .A2(n49), .ZN(y[79]) );
  AND2_X1 U72 ( .A1(b[79]), .A2(sel), .ZN(n49) );
  AND2_X1 U73 ( .A1(a[79]), .A2(n258), .ZN(n48) );
  OR2_X1 U74 ( .A1(n50), .A2(n51), .ZN(y[78]) );
  AND2_X1 U75 ( .A1(b[78]), .A2(sel), .ZN(n51) );
  AND2_X1 U76 ( .A1(a[78]), .A2(n259), .ZN(n50) );
  OR2_X1 U77 ( .A1(n52), .A2(n53), .ZN(y[77]) );
  AND2_X1 U78 ( .A1(b[77]), .A2(sel), .ZN(n53) );
  AND2_X1 U79 ( .A1(a[77]), .A2(n1), .ZN(n52) );
  OR2_X1 U80 ( .A1(n54), .A2(n55), .ZN(y[76]) );
  AND2_X1 U81 ( .A1(b[76]), .A2(sel), .ZN(n55) );
  AND2_X1 U82 ( .A1(a[76]), .A2(n1), .ZN(n54) );
  OR2_X1 U83 ( .A1(n56), .A2(n57), .ZN(y[75]) );
  AND2_X1 U84 ( .A1(b[75]), .A2(sel), .ZN(n57) );
  AND2_X1 U85 ( .A1(a[75]), .A2(n260), .ZN(n56) );
  OR2_X1 U86 ( .A1(n58), .A2(n59), .ZN(y[74]) );
  AND2_X1 U87 ( .A1(b[74]), .A2(sel), .ZN(n59) );
  AND2_X1 U88 ( .A1(a[74]), .A2(n1), .ZN(n58) );
  OR2_X1 U89 ( .A1(n60), .A2(n61), .ZN(y[73]) );
  AND2_X1 U90 ( .A1(b[73]), .A2(sel), .ZN(n61) );
  AND2_X1 U91 ( .A1(a[73]), .A2(n258), .ZN(n60) );
  OR2_X1 U92 ( .A1(n62), .A2(n63), .ZN(y[72]) );
  AND2_X1 U93 ( .A1(b[72]), .A2(sel), .ZN(n63) );
  AND2_X1 U94 ( .A1(a[72]), .A2(n259), .ZN(n62) );
  OR2_X1 U95 ( .A1(n64), .A2(n65), .ZN(y[71]) );
  AND2_X1 U96 ( .A1(b[71]), .A2(sel), .ZN(n65) );
  AND2_X1 U97 ( .A1(a[71]), .A2(n1), .ZN(n64) );
  OR2_X1 U98 ( .A1(n66), .A2(n67), .ZN(y[70]) );
  AND2_X1 U99 ( .A1(b[70]), .A2(sel), .ZN(n67) );
  AND2_X1 U100 ( .A1(a[70]), .A2(n260), .ZN(n66) );
  OR2_X1 U101 ( .A1(n68), .A2(n69), .ZN(y[6]) );
  AND2_X1 U102 ( .A1(b[6]), .A2(sel), .ZN(n69) );
  AND2_X1 U103 ( .A1(a[6]), .A2(n260), .ZN(n68) );
  OR2_X1 U104 ( .A1(n70), .A2(n71), .ZN(y[69]) );
  AND2_X1 U105 ( .A1(b[69]), .A2(sel), .ZN(n71) );
  AND2_X1 U106 ( .A1(a[69]), .A2(n260), .ZN(n70) );
  OR2_X1 U107 ( .A1(n72), .A2(n73), .ZN(y[68]) );
  AND2_X1 U108 ( .A1(b[68]), .A2(sel), .ZN(n73) );
  AND2_X1 U109 ( .A1(a[68]), .A2(n1), .ZN(n72) );
  OR2_X1 U110 ( .A1(n74), .A2(n75), .ZN(y[67]) );
  AND2_X1 U111 ( .A1(b[67]), .A2(sel), .ZN(n75) );
  AND2_X1 U112 ( .A1(a[67]), .A2(n260), .ZN(n74) );
  OR2_X1 U113 ( .A1(n76), .A2(n77), .ZN(y[66]) );
  AND2_X1 U114 ( .A1(b[66]), .A2(sel), .ZN(n77) );
  AND2_X1 U115 ( .A1(a[66]), .A2(n258), .ZN(n76) );
  OR2_X1 U116 ( .A1(n78), .A2(n79), .ZN(y[65]) );
  AND2_X1 U117 ( .A1(b[65]), .A2(sel), .ZN(n79) );
  AND2_X1 U118 ( .A1(a[65]), .A2(n1), .ZN(n78) );
  OR2_X1 U119 ( .A1(n80), .A2(n81), .ZN(y[64]) );
  AND2_X1 U120 ( .A1(b[64]), .A2(sel), .ZN(n81) );
  AND2_X1 U121 ( .A1(a[64]), .A2(n1), .ZN(n80) );
  OR2_X1 U122 ( .A1(n82), .A2(n83), .ZN(y[63]) );
  AND2_X1 U123 ( .A1(b[63]), .A2(sel), .ZN(n83) );
  AND2_X1 U124 ( .A1(a[63]), .A2(n259), .ZN(n82) );
  OR2_X1 U125 ( .A1(n84), .A2(n85), .ZN(y[62]) );
  AND2_X1 U126 ( .A1(b[62]), .A2(sel), .ZN(n85) );
  AND2_X1 U127 ( .A1(a[62]), .A2(n258), .ZN(n84) );
  OR2_X1 U128 ( .A1(n86), .A2(n87), .ZN(y[61]) );
  AND2_X1 U129 ( .A1(b[61]), .A2(sel), .ZN(n87) );
  AND2_X1 U130 ( .A1(a[61]), .A2(n260), .ZN(n86) );
  OR2_X1 U131 ( .A1(n88), .A2(n89), .ZN(y[60]) );
  AND2_X1 U132 ( .A1(b[60]), .A2(sel), .ZN(n89) );
  AND2_X1 U133 ( .A1(a[60]), .A2(n259), .ZN(n88) );
  OR2_X1 U134 ( .A1(n90), .A2(n91), .ZN(y[5]) );
  AND2_X1 U135 ( .A1(b[5]), .A2(sel), .ZN(n91) );
  AND2_X1 U136 ( .A1(a[5]), .A2(n1), .ZN(n90) );
  OR2_X1 U137 ( .A1(n92), .A2(n93), .ZN(y[59]) );
  AND2_X1 U138 ( .A1(b[59]), .A2(sel), .ZN(n93) );
  AND2_X1 U139 ( .A1(a[59]), .A2(n259), .ZN(n92) );
  OR2_X1 U140 ( .A1(n94), .A2(n95), .ZN(y[58]) );
  AND2_X1 U141 ( .A1(b[58]), .A2(sel), .ZN(n95) );
  AND2_X1 U142 ( .A1(a[58]), .A2(n258), .ZN(n94) );
  OR2_X1 U143 ( .A1(n96), .A2(n97), .ZN(y[57]) );
  AND2_X1 U144 ( .A1(b[57]), .A2(sel), .ZN(n97) );
  AND2_X1 U145 ( .A1(a[57]), .A2(n1), .ZN(n96) );
  OR2_X1 U146 ( .A1(n98), .A2(n99), .ZN(y[56]) );
  AND2_X1 U147 ( .A1(b[56]), .A2(sel), .ZN(n99) );
  AND2_X1 U148 ( .A1(a[56]), .A2(n259), .ZN(n98) );
  OR2_X1 U149 ( .A1(n100), .A2(n101), .ZN(y[55]) );
  AND2_X1 U150 ( .A1(b[55]), .A2(sel), .ZN(n101) );
  AND2_X1 U151 ( .A1(a[55]), .A2(n1), .ZN(n100) );
  OR2_X1 U152 ( .A1(n102), .A2(n103), .ZN(y[54]) );
  AND2_X1 U153 ( .A1(b[54]), .A2(sel), .ZN(n103) );
  AND2_X1 U154 ( .A1(a[54]), .A2(n259), .ZN(n102) );
  OR2_X1 U155 ( .A1(n104), .A2(n105), .ZN(y[53]) );
  AND2_X1 U156 ( .A1(b[53]), .A2(sel), .ZN(n105) );
  AND2_X1 U157 ( .A1(a[53]), .A2(n259), .ZN(n104) );
  OR2_X1 U158 ( .A1(n106), .A2(n107), .ZN(y[52]) );
  AND2_X1 U159 ( .A1(b[52]), .A2(sel), .ZN(n107) );
  AND2_X1 U160 ( .A1(a[52]), .A2(n260), .ZN(n106) );
  OR2_X1 U161 ( .A1(n108), .A2(n109), .ZN(y[51]) );
  AND2_X1 U162 ( .A1(b[51]), .A2(sel), .ZN(n109) );
  AND2_X1 U163 ( .A1(a[51]), .A2(n1), .ZN(n108) );
  OR2_X1 U164 ( .A1(n110), .A2(n111), .ZN(y[50]) );
  AND2_X1 U165 ( .A1(b[50]), .A2(sel), .ZN(n111) );
  AND2_X1 U166 ( .A1(a[50]), .A2(n259), .ZN(n110) );
  OR2_X1 U167 ( .A1(n112), .A2(n113), .ZN(y[4]) );
  AND2_X1 U168 ( .A1(b[4]), .A2(sel), .ZN(n113) );
  AND2_X1 U169 ( .A1(a[4]), .A2(n260), .ZN(n112) );
  OR2_X1 U170 ( .A1(n114), .A2(n115), .ZN(y[49]) );
  AND2_X1 U171 ( .A1(b[49]), .A2(sel), .ZN(n115) );
  AND2_X1 U172 ( .A1(a[49]), .A2(n1), .ZN(n114) );
  OR2_X1 U173 ( .A1(n116), .A2(n117), .ZN(y[48]) );
  AND2_X1 U174 ( .A1(b[48]), .A2(sel), .ZN(n117) );
  AND2_X1 U175 ( .A1(a[48]), .A2(n258), .ZN(n116) );
  OR2_X1 U176 ( .A1(n118), .A2(n119), .ZN(y[47]) );
  AND2_X1 U177 ( .A1(b[47]), .A2(sel), .ZN(n119) );
  AND2_X1 U178 ( .A1(a[47]), .A2(n260), .ZN(n118) );
  OR2_X1 U179 ( .A1(n120), .A2(n121), .ZN(y[46]) );
  AND2_X1 U180 ( .A1(b[46]), .A2(sel), .ZN(n121) );
  AND2_X1 U181 ( .A1(a[46]), .A2(n260), .ZN(n120) );
  OR2_X1 U182 ( .A1(n122), .A2(n123), .ZN(y[45]) );
  AND2_X1 U183 ( .A1(b[45]), .A2(sel), .ZN(n123) );
  AND2_X1 U184 ( .A1(a[45]), .A2(n258), .ZN(n122) );
  OR2_X1 U185 ( .A1(n124), .A2(n125), .ZN(y[44]) );
  AND2_X1 U186 ( .A1(b[44]), .A2(sel), .ZN(n125) );
  AND2_X1 U187 ( .A1(a[44]), .A2(n259), .ZN(n124) );
  OR2_X1 U188 ( .A1(n126), .A2(n127), .ZN(y[43]) );
  AND2_X1 U189 ( .A1(b[43]), .A2(sel), .ZN(n127) );
  AND2_X1 U190 ( .A1(a[43]), .A2(n258), .ZN(n126) );
  OR2_X1 U191 ( .A1(n128), .A2(n129), .ZN(y[42]) );
  AND2_X1 U192 ( .A1(b[42]), .A2(sel), .ZN(n129) );
  AND2_X1 U193 ( .A1(a[42]), .A2(n1), .ZN(n128) );
  OR2_X1 U194 ( .A1(n130), .A2(n131), .ZN(y[41]) );
  AND2_X1 U195 ( .A1(b[41]), .A2(sel), .ZN(n131) );
  AND2_X1 U196 ( .A1(a[41]), .A2(n260), .ZN(n130) );
  OR2_X1 U197 ( .A1(n132), .A2(n133), .ZN(y[40]) );
  AND2_X1 U198 ( .A1(b[40]), .A2(sel), .ZN(n133) );
  AND2_X1 U199 ( .A1(a[40]), .A2(n260), .ZN(n132) );
  OR2_X1 U200 ( .A1(n134), .A2(n135), .ZN(y[3]) );
  AND2_X1 U201 ( .A1(b[3]), .A2(sel), .ZN(n135) );
  AND2_X1 U202 ( .A1(a[3]), .A2(n258), .ZN(n134) );
  OR2_X1 U203 ( .A1(n136), .A2(n137), .ZN(y[39]) );
  AND2_X1 U204 ( .A1(b[39]), .A2(sel), .ZN(n137) );
  AND2_X1 U205 ( .A1(a[39]), .A2(n259), .ZN(n136) );
  OR2_X1 U206 ( .A1(n138), .A2(n139), .ZN(y[38]) );
  AND2_X1 U207 ( .A1(b[38]), .A2(sel), .ZN(n139) );
  AND2_X1 U208 ( .A1(a[38]), .A2(n259), .ZN(n138) );
  OR2_X1 U209 ( .A1(n140), .A2(n141), .ZN(y[37]) );
  AND2_X1 U210 ( .A1(b[37]), .A2(sel), .ZN(n141) );
  AND2_X1 U211 ( .A1(a[37]), .A2(n1), .ZN(n140) );
  OR2_X1 U212 ( .A1(n142), .A2(n143), .ZN(y[36]) );
  AND2_X1 U213 ( .A1(b[36]), .A2(sel), .ZN(n143) );
  AND2_X1 U214 ( .A1(a[36]), .A2(n260), .ZN(n142) );
  OR2_X1 U215 ( .A1(n144), .A2(n145), .ZN(y[35]) );
  AND2_X1 U216 ( .A1(b[35]), .A2(sel), .ZN(n145) );
  AND2_X1 U217 ( .A1(a[35]), .A2(n260), .ZN(n144) );
  OR2_X1 U218 ( .A1(n146), .A2(n147), .ZN(y[34]) );
  AND2_X1 U219 ( .A1(b[34]), .A2(sel), .ZN(n147) );
  AND2_X1 U220 ( .A1(a[34]), .A2(n1), .ZN(n146) );
  OR2_X1 U221 ( .A1(n148), .A2(n149), .ZN(y[33]) );
  AND2_X1 U222 ( .A1(b[33]), .A2(sel), .ZN(n149) );
  AND2_X1 U223 ( .A1(a[33]), .A2(n260), .ZN(n148) );
  OR2_X1 U224 ( .A1(n150), .A2(n151), .ZN(y[32]) );
  AND2_X1 U225 ( .A1(b[32]), .A2(sel), .ZN(n151) );
  AND2_X1 U226 ( .A1(a[32]), .A2(n258), .ZN(n150) );
  OR2_X1 U227 ( .A1(n152), .A2(n153), .ZN(y[31]) );
  AND2_X1 U228 ( .A1(b[31]), .A2(sel), .ZN(n153) );
  AND2_X1 U229 ( .A1(a[31]), .A2(n259), .ZN(n152) );
  OR2_X1 U230 ( .A1(n154), .A2(n155), .ZN(y[30]) );
  AND2_X1 U231 ( .A1(b[30]), .A2(sel), .ZN(n155) );
  AND2_X1 U232 ( .A1(a[30]), .A2(n260), .ZN(n154) );
  OR2_X1 U233 ( .A1(n156), .A2(n157), .ZN(y[2]) );
  AND2_X1 U234 ( .A1(b[2]), .A2(sel), .ZN(n157) );
  AND2_X1 U235 ( .A1(a[2]), .A2(n258), .ZN(n156) );
  OR2_X1 U236 ( .A1(n158), .A2(n159), .ZN(y[29]) );
  AND2_X1 U237 ( .A1(b[29]), .A2(sel), .ZN(n159) );
  AND2_X1 U238 ( .A1(a[29]), .A2(n259), .ZN(n158) );
  OR2_X1 U239 ( .A1(n160), .A2(n161), .ZN(y[28]) );
  AND2_X1 U240 ( .A1(b[28]), .A2(sel), .ZN(n161) );
  AND2_X1 U241 ( .A1(a[28]), .A2(n259), .ZN(n160) );
  OR2_X1 U242 ( .A1(n162), .A2(n163), .ZN(y[27]) );
  AND2_X1 U243 ( .A1(b[27]), .A2(sel), .ZN(n163) );
  AND2_X1 U244 ( .A1(a[27]), .A2(n260), .ZN(n162) );
  OR2_X1 U245 ( .A1(n164), .A2(n165), .ZN(y[26]) );
  AND2_X1 U246 ( .A1(b[26]), .A2(sel), .ZN(n165) );
  AND2_X1 U247 ( .A1(a[26]), .A2(n259), .ZN(n164) );
  OR2_X1 U248 ( .A1(n166), .A2(n167), .ZN(y[25]) );
  AND2_X1 U249 ( .A1(b[25]), .A2(sel), .ZN(n167) );
  AND2_X1 U250 ( .A1(a[25]), .A2(n259), .ZN(n166) );
  OR2_X1 U251 ( .A1(n168), .A2(n169), .ZN(y[24]) );
  AND2_X1 U252 ( .A1(b[24]), .A2(sel), .ZN(n169) );
  AND2_X1 U253 ( .A1(a[24]), .A2(n260), .ZN(n168) );
  OR2_X1 U254 ( .A1(n170), .A2(n171), .ZN(y[23]) );
  AND2_X1 U255 ( .A1(b[23]), .A2(sel), .ZN(n171) );
  AND2_X1 U256 ( .A1(a[23]), .A2(n1), .ZN(n170) );
  OR2_X1 U257 ( .A1(n172), .A2(n173), .ZN(y[22]) );
  AND2_X1 U258 ( .A1(b[22]), .A2(sel), .ZN(n173) );
  AND2_X1 U259 ( .A1(a[22]), .A2(n258), .ZN(n172) );
  OR2_X1 U260 ( .A1(n174), .A2(n175), .ZN(y[21]) );
  AND2_X1 U261 ( .A1(b[21]), .A2(sel), .ZN(n175) );
  AND2_X1 U262 ( .A1(a[21]), .A2(n259), .ZN(n174) );
  OR2_X1 U263 ( .A1(n176), .A2(n177), .ZN(y[20]) );
  AND2_X1 U264 ( .A1(b[20]), .A2(sel), .ZN(n177) );
  AND2_X1 U265 ( .A1(a[20]), .A2(n259), .ZN(n176) );
  OR2_X1 U266 ( .A1(n178), .A2(n179), .ZN(y[1]) );
  AND2_X1 U267 ( .A1(b[1]), .A2(sel), .ZN(n179) );
  AND2_X1 U268 ( .A1(a[1]), .A2(n1), .ZN(n178) );
  OR2_X1 U269 ( .A1(n180), .A2(n181), .ZN(y[19]) );
  AND2_X1 U270 ( .A1(b[19]), .A2(sel), .ZN(n181) );
  AND2_X1 U271 ( .A1(a[19]), .A2(n260), .ZN(n180) );
  OR2_X1 U272 ( .A1(n182), .A2(n183), .ZN(y[18]) );
  AND2_X1 U273 ( .A1(b[18]), .A2(sel), .ZN(n183) );
  AND2_X1 U274 ( .A1(a[18]), .A2(n258), .ZN(n182) );
  OR2_X1 U275 ( .A1(n184), .A2(n185), .ZN(y[17]) );
  AND2_X1 U276 ( .A1(b[17]), .A2(sel), .ZN(n185) );
  AND2_X1 U277 ( .A1(a[17]), .A2(n258), .ZN(n184) );
  OR2_X1 U278 ( .A1(n186), .A2(n187), .ZN(y[16]) );
  AND2_X1 U279 ( .A1(b[16]), .A2(sel), .ZN(n187) );
  AND2_X1 U280 ( .A1(a[16]), .A2(n260), .ZN(n186) );
  OR2_X1 U281 ( .A1(n188), .A2(n189), .ZN(y[15]) );
  AND2_X1 U282 ( .A1(b[15]), .A2(sel), .ZN(n189) );
  AND2_X1 U283 ( .A1(a[15]), .A2(n259), .ZN(n188) );
  OR2_X1 U284 ( .A1(n190), .A2(n191), .ZN(y[14]) );
  AND2_X1 U285 ( .A1(b[14]), .A2(sel), .ZN(n191) );
  AND2_X1 U286 ( .A1(a[14]), .A2(n1), .ZN(n190) );
  OR2_X1 U287 ( .A1(n192), .A2(n193), .ZN(y[13]) );
  AND2_X1 U288 ( .A1(b[13]), .A2(sel), .ZN(n193) );
  AND2_X1 U289 ( .A1(a[13]), .A2(n1), .ZN(n192) );
  OR2_X1 U290 ( .A1(n194), .A2(n195), .ZN(y[12]) );
  AND2_X1 U291 ( .A1(b[12]), .A2(sel), .ZN(n195) );
  AND2_X1 U292 ( .A1(a[12]), .A2(n260), .ZN(n194) );
  OR2_X1 U293 ( .A1(n196), .A2(n197), .ZN(y[127]) );
  AND2_X1 U294 ( .A1(b[127]), .A2(sel), .ZN(n197) );
  AND2_X1 U295 ( .A1(a[127]), .A2(n1), .ZN(n196) );
  OR2_X1 U296 ( .A1(n198), .A2(n199), .ZN(y[126]) );
  AND2_X1 U297 ( .A1(b[126]), .A2(sel), .ZN(n199) );
  AND2_X1 U298 ( .A1(a[126]), .A2(n259), .ZN(n198) );
  OR2_X1 U299 ( .A1(n200), .A2(n201), .ZN(y[125]) );
  AND2_X1 U300 ( .A1(b[125]), .A2(sel), .ZN(n201) );
  AND2_X1 U301 ( .A1(a[125]), .A2(n1), .ZN(n200) );
  OR2_X1 U302 ( .A1(n202), .A2(n203), .ZN(y[124]) );
  AND2_X1 U303 ( .A1(b[124]), .A2(sel), .ZN(n203) );
  AND2_X1 U304 ( .A1(a[124]), .A2(n259), .ZN(n202) );
  OR2_X1 U305 ( .A1(n204), .A2(n205), .ZN(y[123]) );
  AND2_X1 U306 ( .A1(b[123]), .A2(sel), .ZN(n205) );
  AND2_X1 U307 ( .A1(a[123]), .A2(n259), .ZN(n204) );
  OR2_X1 U308 ( .A1(n206), .A2(n207), .ZN(y[122]) );
  AND2_X1 U309 ( .A1(b[122]), .A2(sel), .ZN(n207) );
  AND2_X1 U310 ( .A1(a[122]), .A2(n1), .ZN(n206) );
  OR2_X1 U311 ( .A1(n208), .A2(n209), .ZN(y[121]) );
  AND2_X1 U312 ( .A1(b[121]), .A2(sel), .ZN(n209) );
  AND2_X1 U313 ( .A1(a[121]), .A2(n259), .ZN(n208) );
  OR2_X1 U314 ( .A1(n210), .A2(n211), .ZN(y[120]) );
  AND2_X1 U315 ( .A1(b[120]), .A2(sel), .ZN(n211) );
  AND2_X1 U316 ( .A1(a[120]), .A2(n259), .ZN(n210) );
  OR2_X1 U317 ( .A1(n212), .A2(n213), .ZN(y[11]) );
  AND2_X1 U318 ( .A1(b[11]), .A2(sel), .ZN(n213) );
  AND2_X1 U319 ( .A1(a[11]), .A2(n260), .ZN(n212) );
  OR2_X1 U320 ( .A1(n214), .A2(n215), .ZN(y[119]) );
  AND2_X1 U321 ( .A1(b[119]), .A2(sel), .ZN(n215) );
  AND2_X1 U322 ( .A1(a[119]), .A2(n260), .ZN(n214) );
  OR2_X1 U323 ( .A1(n216), .A2(n217), .ZN(y[118]) );
  AND2_X1 U324 ( .A1(b[118]), .A2(sel), .ZN(n217) );
  AND2_X1 U325 ( .A1(a[118]), .A2(n1), .ZN(n216) );
  OR2_X1 U326 ( .A1(n218), .A2(n219), .ZN(y[117]) );
  AND2_X1 U327 ( .A1(b[117]), .A2(sel), .ZN(n219) );
  AND2_X1 U328 ( .A1(a[117]), .A2(n259), .ZN(n218) );
  OR2_X1 U329 ( .A1(n220), .A2(n221), .ZN(y[116]) );
  AND2_X1 U330 ( .A1(b[116]), .A2(sel), .ZN(n221) );
  AND2_X1 U331 ( .A1(a[116]), .A2(n1), .ZN(n220) );
  OR2_X1 U332 ( .A1(n222), .A2(n223), .ZN(y[115]) );
  AND2_X1 U333 ( .A1(b[115]), .A2(sel), .ZN(n223) );
  AND2_X1 U334 ( .A1(a[115]), .A2(n258), .ZN(n222) );
  OR2_X1 U335 ( .A1(n224), .A2(n225), .ZN(y[114]) );
  AND2_X1 U336 ( .A1(b[114]), .A2(sel), .ZN(n225) );
  AND2_X1 U337 ( .A1(a[114]), .A2(n258), .ZN(n224) );
  OR2_X1 U338 ( .A1(n226), .A2(n227), .ZN(y[113]) );
  AND2_X1 U339 ( .A1(b[113]), .A2(sel), .ZN(n227) );
  AND2_X1 U340 ( .A1(a[113]), .A2(n259), .ZN(n226) );
  OR2_X1 U341 ( .A1(n228), .A2(n229), .ZN(y[112]) );
  AND2_X1 U342 ( .A1(b[112]), .A2(sel), .ZN(n229) );
  AND2_X1 U343 ( .A1(a[112]), .A2(n260), .ZN(n228) );
  OR2_X1 U344 ( .A1(n230), .A2(n231), .ZN(y[111]) );
  AND2_X1 U345 ( .A1(b[111]), .A2(sel), .ZN(n231) );
  AND2_X1 U346 ( .A1(a[111]), .A2(n1), .ZN(n230) );
  OR2_X1 U347 ( .A1(n232), .A2(n233), .ZN(y[110]) );
  AND2_X1 U348 ( .A1(b[110]), .A2(sel), .ZN(n233) );
  AND2_X1 U349 ( .A1(a[110]), .A2(n259), .ZN(n232) );
  OR2_X1 U350 ( .A1(n234), .A2(n235), .ZN(y[10]) );
  AND2_X1 U351 ( .A1(b[10]), .A2(sel), .ZN(n235) );
  AND2_X1 U352 ( .A1(a[10]), .A2(n1), .ZN(n234) );
  OR2_X1 U353 ( .A1(n236), .A2(n237), .ZN(y[109]) );
  AND2_X1 U354 ( .A1(b[109]), .A2(sel), .ZN(n237) );
  AND2_X1 U355 ( .A1(a[109]), .A2(n259), .ZN(n236) );
  OR2_X1 U356 ( .A1(n238), .A2(n239), .ZN(y[108]) );
  AND2_X1 U357 ( .A1(b[108]), .A2(sel), .ZN(n239) );
  AND2_X1 U358 ( .A1(a[108]), .A2(n1), .ZN(n238) );
  OR2_X1 U359 ( .A1(n240), .A2(n241), .ZN(y[107]) );
  AND2_X1 U360 ( .A1(b[107]), .A2(sel), .ZN(n241) );
  AND2_X1 U361 ( .A1(a[107]), .A2(n260), .ZN(n240) );
  OR2_X1 U362 ( .A1(n242), .A2(n243), .ZN(y[106]) );
  AND2_X1 U363 ( .A1(b[106]), .A2(sel), .ZN(n243) );
  AND2_X1 U364 ( .A1(a[106]), .A2(n1), .ZN(n242) );
  OR2_X1 U365 ( .A1(n244), .A2(n245), .ZN(y[105]) );
  AND2_X1 U366 ( .A1(b[105]), .A2(sel), .ZN(n245) );
  AND2_X1 U367 ( .A1(a[105]), .A2(n260), .ZN(n244) );
  OR2_X1 U368 ( .A1(n246), .A2(n247), .ZN(y[104]) );
  AND2_X1 U369 ( .A1(b[104]), .A2(sel), .ZN(n247) );
  AND2_X1 U370 ( .A1(a[104]), .A2(n258), .ZN(n246) );
  OR2_X1 U371 ( .A1(n248), .A2(n249), .ZN(y[103]) );
  AND2_X1 U372 ( .A1(b[103]), .A2(sel), .ZN(n249) );
  AND2_X1 U373 ( .A1(a[103]), .A2(n258), .ZN(n248) );
  OR2_X1 U374 ( .A1(n250), .A2(n251), .ZN(y[102]) );
  AND2_X1 U375 ( .A1(b[102]), .A2(sel), .ZN(n251) );
  AND2_X1 U376 ( .A1(a[102]), .A2(n260), .ZN(n250) );
  OR2_X1 U377 ( .A1(n252), .A2(n253), .ZN(y[101]) );
  AND2_X1 U378 ( .A1(b[101]), .A2(sel), .ZN(n253) );
  AND2_X1 U379 ( .A1(a[101]), .A2(n260), .ZN(n252) );
  OR2_X1 U380 ( .A1(n254), .A2(n255), .ZN(y[100]) );
  AND2_X1 U381 ( .A1(b[100]), .A2(sel), .ZN(n255) );
  AND2_X1 U382 ( .A1(a[100]), .A2(n259), .ZN(n254) );
  OR2_X1 U383 ( .A1(n256), .A2(n257), .ZN(y[0]) );
  AND2_X1 U384 ( .A1(b[0]), .A2(sel), .ZN(n257) );
  AND2_X1 U385 ( .A1(a[0]), .A2(n1), .ZN(n256) );
  INV_X1 U1 ( .A(sel), .ZN(n1) );
  INV_X1 U386 ( .A(sel), .ZN(n258) );
  INV_X1 U387 ( .A(sel), .ZN(n259) );
  INV_X1 U388 ( .A(sel), .ZN(n260) );
endmodule


module shiftRows ( in, out );
  input [127:0] in;
  //input_done

  output [127:0] out;
  //output_done

  //wire_done

  assign out[127] = in[127];
  assign out[126] = in[126];
  assign out[125] = in[125];
  assign out[124] = in[124];
  assign out[123] = in[123];
  assign out[122] = in[122];
  assign out[121] = in[121];
  assign out[120] = in[120];
  assign out[119] = in[87];
  assign out[118] = in[86];
  assign out[117] = in[85];
  assign out[116] = in[84];
  assign out[115] = in[83];
  assign out[114] = in[82];
  assign out[113] = in[81];
  assign out[112] = in[80];
  assign out[111] = in[47];
  assign out[110] = in[46];
  assign out[109] = in[45];
  assign out[108] = in[44];
  assign out[107] = in[43];
  assign out[106] = in[42];
  assign out[105] = in[41];
  assign out[104] = in[40];
  assign out[103] = in[7];
  assign out[102] = in[6];
  assign out[101] = in[5];
  assign out[100] = in[4];
  assign out[99] = in[3];
  assign out[98] = in[2];
  assign out[97] = in[1];
  assign out[96] = in[0];
  assign out[95] = in[95];
  assign out[94] = in[94];
  assign out[93] = in[93];
  assign out[92] = in[92];
  assign out[91] = in[91];
  assign out[90] = in[90];
  assign out[89] = in[89];
  assign out[88] = in[88];
  assign out[87] = in[55];
  assign out[86] = in[54];
  assign out[85] = in[53];
  assign out[84] = in[52];
  assign out[83] = in[51];
  assign out[82] = in[50];
  assign out[81] = in[49];
  assign out[80] = in[48];
  assign out[79] = in[15];
  assign out[78] = in[14];
  assign out[77] = in[13];
  assign out[76] = in[12];
  assign out[75] = in[11];
  assign out[74] = in[10];
  assign out[73] = in[9];
  assign out[72] = in[8];
  assign out[71] = in[103];
  assign out[70] = in[102];
  assign out[69] = in[101];
  assign out[68] = in[100];
  assign out[67] = in[99];
  assign out[66] = in[98];
  assign out[65] = in[97];
  assign out[64] = in[96];
  assign out[63] = in[63];
  assign out[62] = in[62];
  assign out[61] = in[61];
  assign out[60] = in[60];
  assign out[59] = in[59];
  assign out[58] = in[58];
  assign out[57] = in[57];
  assign out[56] = in[56];
  assign out[55] = in[23];
  assign out[54] = in[22];
  assign out[53] = in[21];
  assign out[52] = in[20];
  assign out[51] = in[19];
  assign out[50] = in[18];
  assign out[49] = in[17];
  assign out[48] = in[16];
  assign out[47] = in[111];
  assign out[46] = in[110];
  assign out[45] = in[109];
  assign out[44] = in[108];
  assign out[43] = in[107];
  assign out[42] = in[106];
  assign out[41] = in[105];
  assign out[40] = in[104];
  assign out[39] = in[71];
  assign out[38] = in[70];
  assign out[37] = in[69];
  assign out[36] = in[68];
  assign out[35] = in[67];
  assign out[34] = in[66];
  assign out[33] = in[65];
  assign out[32] = in[64];
  assign out[31] = in[31];
  assign out[30] = in[30];
  assign out[29] = in[29];
  assign out[28] = in[28];
  assign out[27] = in[27];
  assign out[26] = in[26];
  assign out[25] = in[25];
  assign out[24] = in[24];
  assign out[23] = in[119];
  assign out[22] = in[118];
  assign out[21] = in[117];
  assign out[20] = in[116];
  assign out[19] = in[115];
  assign out[18] = in[114];
  assign out[17] = in[113];
  assign out[16] = in[112];
  assign out[15] = in[79];
  assign out[14] = in[78];
  assign out[13] = in[77];
  assign out[12] = in[76];
  assign out[11] = in[75];
  assign out[10] = in[74];
  assign out[9] = in[73];
  assign out[8] = in[72];
  assign out[7] = in[39];
  assign out[6] = in[38];
  assign out[5] = in[37];
  assign out[4] = in[36];
  assign out[3] = in[35];
  assign out[2] = in[34];
  assign out[1] = in[33];
  assign out[0] = in[32];

endmodule


module CD2_0 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done

  wire   n1, n2;
  wire n1bar, n2bar;
  //wire_done

  assign n1bar = a;
  assign n1 = abar;
  assign n2bar = b;
  assign n2 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n2), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n2bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n1), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n1bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n1bar), .A2(n2bar), .ZN(ybar[0]);
endmodule




module CD4_0 ( a, b, y );
  input [3:0] a;
  input [3:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  //input_done

  output [15:0] y;
  reg [15:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]);
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]);
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]);
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]);
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]);
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]);
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]);
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]);
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]);
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]);
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]);
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]);
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]);
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]);
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]);
endmodule




module CD16_0 ( a, b, y );
  input [15:0] a;
  input [15:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign abar[8] = ~a[8];
  assign abar[9] = ~a[9];
  assign abar[10] = ~a[10];
  assign abar[11] = ~a[11];
  assign abar[12] = ~a[12];
  assign abar[13] = ~a[13];
  assign abar[14] = ~a[14];
  assign abar[15] = ~a[15];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign bbar[8] = ~b[8];
  assign bbar[9] = ~b[9];
  assign bbar[10] = ~b[10];
  assign bbar[11] = ~b[11];
  assign bbar[12] = ~b[12];
  assign bbar[13] = ~b[13];
  assign bbar[14] = ~b[14];
  assign bbar[15] = ~b[15];
  //input_done

  output [255:0] y;
  reg [255:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[9]), .A2(a[0]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[9]), .A2(abar[0]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[3]), .A2(a[6]), .ZN(y[99]) );
  OR2_X1 U2bar ( .A1(bbar[3]), .A2(abar[6]), .ZN(ybar[99]);
  AND2_X1 U3 ( .A1(b[2]), .A2(a[6]), .ZN(y[98]) );
  OR2_X1 U3bar ( .A1(bbar[2]), .A2(abar[6]), .ZN(ybar[98]);
  AND2_X1 U4 ( .A1(b[1]), .A2(a[6]), .ZN(y[97]) );
  OR2_X1 U4bar ( .A1(bbar[1]), .A2(abar[6]), .ZN(ybar[97]);
  AND2_X1 U5 ( .A1(b[0]), .A2(a[6]), .ZN(y[96]) );
  OR2_X1 U5bar ( .A1(bbar[0]), .A2(abar[6]), .ZN(ybar[96]);
  AND2_X1 U6 ( .A1(b[15]), .A2(a[5]), .ZN(y[95]) );
  OR2_X1 U6bar ( .A1(bbar[15]), .A2(abar[5]), .ZN(ybar[95]);
  AND2_X1 U7 ( .A1(b[14]), .A2(a[5]), .ZN(y[94]) );
  OR2_X1 U7bar ( .A1(bbar[14]), .A2(abar[5]), .ZN(ybar[94]);
  AND2_X1 U8 ( .A1(b[13]), .A2(a[5]), .ZN(y[93]) );
  OR2_X1 U8bar ( .A1(bbar[13]), .A2(abar[5]), .ZN(ybar[93]);
  AND2_X1 U9 ( .A1(b[12]), .A2(a[5]), .ZN(y[92]) );
  OR2_X1 U9bar ( .A1(bbar[12]), .A2(abar[5]), .ZN(ybar[92]);
  AND2_X1 U10 ( .A1(b[11]), .A2(a[5]), .ZN(y[91]) );
  OR2_X1 U10bar ( .A1(bbar[11]), .A2(abar[5]), .ZN(ybar[91]);
  AND2_X1 U11 ( .A1(b[10]), .A2(a[5]), .ZN(y[90]) );
  OR2_X1 U11bar ( .A1(bbar[10]), .A2(abar[5]), .ZN(ybar[90]);
  AND2_X1 U12 ( .A1(b[8]), .A2(a[0]), .ZN(y[8]) );
  OR2_X1 U12bar ( .A1(bbar[8]), .A2(abar[0]), .ZN(ybar[8]);
  AND2_X1 U13 ( .A1(a[5]), .A2(b[9]), .ZN(y[89]) );
  OR2_X1 U13bar ( .A1(abar[5]), .A2(bbar[9]), .ZN(ybar[89]);
  AND2_X1 U14 ( .A1(b[8]), .A2(a[5]), .ZN(y[88]) );
  OR2_X1 U14bar ( .A1(bbar[8]), .A2(abar[5]), .ZN(ybar[88]);
  AND2_X1 U15 ( .A1(b[7]), .A2(a[5]), .ZN(y[87]) );
  OR2_X1 U15bar ( .A1(bbar[7]), .A2(abar[5]), .ZN(ybar[87]);
  AND2_X1 U16 ( .A1(b[6]), .A2(a[5]), .ZN(y[86]) );
  OR2_X1 U16bar ( .A1(bbar[6]), .A2(abar[5]), .ZN(ybar[86]);
  AND2_X1 U17 ( .A1(b[5]), .A2(a[5]), .ZN(y[85]) );
  OR2_X1 U17bar ( .A1(bbar[5]), .A2(abar[5]), .ZN(ybar[85]);
  AND2_X1 U18 ( .A1(b[4]), .A2(a[5]), .ZN(y[84]) );
  OR2_X1 U18bar ( .A1(bbar[4]), .A2(abar[5]), .ZN(ybar[84]);
  AND2_X1 U19 ( .A1(a[5]), .A2(b[3]), .ZN(y[83]) );
  OR2_X1 U19bar ( .A1(abar[5]), .A2(bbar[3]), .ZN(ybar[83]);
  AND2_X1 U20 ( .A1(a[5]), .A2(b[2]), .ZN(y[82]) );
  OR2_X1 U20bar ( .A1(abar[5]), .A2(bbar[2]), .ZN(ybar[82]);
  AND2_X1 U21 ( .A1(a[5]), .A2(b[1]), .ZN(y[81]) );
  OR2_X1 U21bar ( .A1(abar[5]), .A2(bbar[1]), .ZN(ybar[81]);
  AND2_X1 U22 ( .A1(a[5]), .A2(b[0]), .ZN(y[80]) );
  OR2_X1 U22bar ( .A1(abar[5]), .A2(bbar[0]), .ZN(ybar[80]);
  AND2_X1 U23 ( .A1(b[7]), .A2(a[0]), .ZN(y[7]) );
  OR2_X1 U23bar ( .A1(bbar[7]), .A2(abar[0]), .ZN(ybar[7]);
  AND2_X1 U24 ( .A1(a[4]), .A2(b[15]), .ZN(y[79]) );
  OR2_X1 U24bar ( .A1(abar[4]), .A2(bbar[15]), .ZN(ybar[79]);
  AND2_X1 U25 ( .A1(a[4]), .A2(b[14]), .ZN(y[78]) );
  OR2_X1 U25bar ( .A1(abar[4]), .A2(bbar[14]), .ZN(ybar[78]);
  AND2_X1 U26 ( .A1(a[4]), .A2(b[13]), .ZN(y[77]) );
  OR2_X1 U26bar ( .A1(abar[4]), .A2(bbar[13]), .ZN(ybar[77]);
  AND2_X1 U27 ( .A1(a[4]), .A2(b[12]), .ZN(y[76]) );
  OR2_X1 U27bar ( .A1(abar[4]), .A2(bbar[12]), .ZN(ybar[76]);
  AND2_X1 U28 ( .A1(a[4]), .A2(b[11]), .ZN(y[75]) );
  OR2_X1 U28bar ( .A1(abar[4]), .A2(bbar[11]), .ZN(ybar[75]);
  AND2_X1 U29 ( .A1(a[4]), .A2(b[10]), .ZN(y[74]) );
  OR2_X1 U29bar ( .A1(abar[4]), .A2(bbar[10]), .ZN(ybar[74]);
  AND2_X1 U30 ( .A1(a[4]), .A2(b[9]), .ZN(y[73]) );
  OR2_X1 U30bar ( .A1(abar[4]), .A2(bbar[9]), .ZN(ybar[73]);
  AND2_X1 U31 ( .A1(a[4]), .A2(b[8]), .ZN(y[72]) );
  OR2_X1 U31bar ( .A1(abar[4]), .A2(bbar[8]), .ZN(ybar[72]);
  AND2_X1 U32 ( .A1(a[4]), .A2(b[7]), .ZN(y[71]) );
  OR2_X1 U32bar ( .A1(abar[4]), .A2(bbar[7]), .ZN(ybar[71]);
  AND2_X1 U33 ( .A1(a[4]), .A2(b[6]), .ZN(y[70]) );
  OR2_X1 U33bar ( .A1(abar[4]), .A2(bbar[6]), .ZN(ybar[70]);
  AND2_X1 U34 ( .A1(b[6]), .A2(a[0]), .ZN(y[6]) );
  OR2_X1 U34bar ( .A1(bbar[6]), .A2(abar[0]), .ZN(ybar[6]);
  AND2_X1 U35 ( .A1(a[4]), .A2(b[5]), .ZN(y[69]) );
  OR2_X1 U35bar ( .A1(abar[4]), .A2(bbar[5]), .ZN(ybar[69]);
  AND2_X1 U36 ( .A1(a[4]), .A2(b[4]), .ZN(y[68]) );
  OR2_X1 U36bar ( .A1(abar[4]), .A2(bbar[4]), .ZN(ybar[68]);
  AND2_X1 U37 ( .A1(a[4]), .A2(b[3]), .ZN(y[67]) );
  OR2_X1 U37bar ( .A1(abar[4]), .A2(bbar[3]), .ZN(ybar[67]);
  AND2_X1 U38 ( .A1(a[4]), .A2(b[2]), .ZN(y[66]) );
  OR2_X1 U38bar ( .A1(abar[4]), .A2(bbar[2]), .ZN(ybar[66]);
  AND2_X1 U39 ( .A1(a[4]), .A2(b[1]), .ZN(y[65]) );
  OR2_X1 U39bar ( .A1(abar[4]), .A2(bbar[1]), .ZN(ybar[65]);
  AND2_X1 U40 ( .A1(a[4]), .A2(b[0]), .ZN(y[64]) );
  OR2_X1 U40bar ( .A1(abar[4]), .A2(bbar[0]), .ZN(ybar[64]);
  AND2_X1 U41 ( .A1(a[3]), .A2(b[15]), .ZN(y[63]) );
  OR2_X1 U41bar ( .A1(abar[3]), .A2(bbar[15]), .ZN(ybar[63]);
  AND2_X1 U42 ( .A1(a[3]), .A2(b[14]), .ZN(y[62]) );
  OR2_X1 U42bar ( .A1(abar[3]), .A2(bbar[14]), .ZN(ybar[62]);
  AND2_X1 U43 ( .A1(a[3]), .A2(b[13]), .ZN(y[61]) );
  OR2_X1 U43bar ( .A1(abar[3]), .A2(bbar[13]), .ZN(ybar[61]);
  AND2_X1 U44 ( .A1(a[3]), .A2(b[12]), .ZN(y[60]) );
  OR2_X1 U44bar ( .A1(abar[3]), .A2(bbar[12]), .ZN(ybar[60]);
  AND2_X1 U45 ( .A1(b[5]), .A2(a[0]), .ZN(y[5]) );
  OR2_X1 U45bar ( .A1(bbar[5]), .A2(abar[0]), .ZN(ybar[5]);
  AND2_X1 U46 ( .A1(a[3]), .A2(b[11]), .ZN(y[59]) );
  OR2_X1 U46bar ( .A1(abar[3]), .A2(bbar[11]), .ZN(ybar[59]);
  AND2_X1 U47 ( .A1(a[3]), .A2(b[10]), .ZN(y[58]) );
  OR2_X1 U47bar ( .A1(abar[3]), .A2(bbar[10]), .ZN(ybar[58]);
  AND2_X1 U48 ( .A1(a[3]), .A2(b[9]), .ZN(y[57]) );
  OR2_X1 U48bar ( .A1(abar[3]), .A2(bbar[9]), .ZN(ybar[57]);
  AND2_X1 U49 ( .A1(a[3]), .A2(b[8]), .ZN(y[56]) );
  OR2_X1 U49bar ( .A1(abar[3]), .A2(bbar[8]), .ZN(ybar[56]);
  AND2_X1 U50 ( .A1(a[3]), .A2(b[7]), .ZN(y[55]) );
  OR2_X1 U50bar ( .A1(abar[3]), .A2(bbar[7]), .ZN(ybar[55]);
  AND2_X1 U51 ( .A1(a[3]), .A2(b[6]), .ZN(y[54]) );
  OR2_X1 U51bar ( .A1(abar[3]), .A2(bbar[6]), .ZN(ybar[54]);
  AND2_X1 U52 ( .A1(a[3]), .A2(b[5]), .ZN(y[53]) );
  OR2_X1 U52bar ( .A1(abar[3]), .A2(bbar[5]), .ZN(ybar[53]);
  AND2_X1 U53 ( .A1(a[3]), .A2(b[4]), .ZN(y[52]) );
  OR2_X1 U53bar ( .A1(abar[3]), .A2(bbar[4]), .ZN(ybar[52]);
  AND2_X1 U54 ( .A1(a[3]), .A2(b[3]), .ZN(y[51]) );
  OR2_X1 U54bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[51]);
  AND2_X1 U55 ( .A1(a[3]), .A2(b[2]), .ZN(y[50]) );
  OR2_X1 U55bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[50]);
  AND2_X1 U56 ( .A1(b[4]), .A2(a[0]), .ZN(y[4]) );
  OR2_X1 U56bar ( .A1(bbar[4]), .A2(abar[0]), .ZN(ybar[4]);
  AND2_X1 U57 ( .A1(a[3]), .A2(b[1]), .ZN(y[49]) );
  OR2_X1 U57bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[49]);
  AND2_X1 U58 ( .A1(a[3]), .A2(b[0]), .ZN(y[48]) );
  OR2_X1 U58bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[48]);
  AND2_X1 U59 ( .A1(a[2]), .A2(b[15]), .ZN(y[47]) );
  OR2_X1 U59bar ( .A1(abar[2]), .A2(bbar[15]), .ZN(ybar[47]);
  AND2_X1 U60 ( .A1(a[2]), .A2(b[14]), .ZN(y[46]) );
  OR2_X1 U60bar ( .A1(abar[2]), .A2(bbar[14]), .ZN(ybar[46]);
  AND2_X1 U61 ( .A1(a[2]), .A2(b[13]), .ZN(y[45]) );
  OR2_X1 U61bar ( .A1(abar[2]), .A2(bbar[13]), .ZN(ybar[45]);
  AND2_X1 U62 ( .A1(a[2]), .A2(b[12]), .ZN(y[44]) );
  OR2_X1 U62bar ( .A1(abar[2]), .A2(bbar[12]), .ZN(ybar[44]);
  AND2_X1 U63 ( .A1(a[2]), .A2(b[11]), .ZN(y[43]) );
  OR2_X1 U63bar ( .A1(abar[2]), .A2(bbar[11]), .ZN(ybar[43]);
  AND2_X1 U64 ( .A1(a[2]), .A2(b[10]), .ZN(y[42]) );
  OR2_X1 U64bar ( .A1(abar[2]), .A2(bbar[10]), .ZN(ybar[42]);
  AND2_X1 U65 ( .A1(a[2]), .A2(b[9]), .ZN(y[41]) );
  OR2_X1 U65bar ( .A1(abar[2]), .A2(bbar[9]), .ZN(ybar[41]);
  AND2_X1 U66 ( .A1(a[2]), .A2(b[8]), .ZN(y[40]) );
  OR2_X1 U66bar ( .A1(abar[2]), .A2(bbar[8]), .ZN(ybar[40]);
  AND2_X1 U67 ( .A1(b[3]), .A2(a[0]), .ZN(y[3]) );
  OR2_X1 U67bar ( .A1(bbar[3]), .A2(abar[0]), .ZN(ybar[3]);
  AND2_X1 U68 ( .A1(a[2]), .A2(b[7]), .ZN(y[39]) );
  OR2_X1 U68bar ( .A1(abar[2]), .A2(bbar[7]), .ZN(ybar[39]);
  AND2_X1 U69 ( .A1(a[2]), .A2(b[6]), .ZN(y[38]) );
  OR2_X1 U69bar ( .A1(abar[2]), .A2(bbar[6]), .ZN(ybar[38]);
  AND2_X1 U70 ( .A1(a[2]), .A2(b[5]), .ZN(y[37]) );
  OR2_X1 U70bar ( .A1(abar[2]), .A2(bbar[5]), .ZN(ybar[37]);
  AND2_X1 U71 ( .A1(a[2]), .A2(b[4]), .ZN(y[36]) );
  OR2_X1 U71bar ( .A1(abar[2]), .A2(bbar[4]), .ZN(ybar[36]);
  AND2_X1 U72 ( .A1(a[2]), .A2(b[3]), .ZN(y[35]) );
  OR2_X1 U72bar ( .A1(abar[2]), .A2(bbar[3]), .ZN(ybar[35]);
  AND2_X1 U73 ( .A1(a[2]), .A2(b[2]), .ZN(y[34]) );
  OR2_X1 U73bar ( .A1(abar[2]), .A2(bbar[2]), .ZN(ybar[34]);
  AND2_X1 U74 ( .A1(a[2]), .A2(b[1]), .ZN(y[33]) );
  OR2_X1 U74bar ( .A1(abar[2]), .A2(bbar[1]), .ZN(ybar[33]);
  AND2_X1 U75 ( .A1(a[2]), .A2(b[0]), .ZN(y[32]) );
  OR2_X1 U75bar ( .A1(abar[2]), .A2(bbar[0]), .ZN(ybar[32]);
  AND2_X1 U76 ( .A1(a[1]), .A2(b[15]), .ZN(y[31]) );
  OR2_X1 U76bar ( .A1(abar[1]), .A2(bbar[15]), .ZN(ybar[31]);
  AND2_X1 U77 ( .A1(a[1]), .A2(b[14]), .ZN(y[30]) );
  OR2_X1 U77bar ( .A1(abar[1]), .A2(bbar[14]), .ZN(ybar[30]);
  AND2_X1 U78 ( .A1(b[2]), .A2(a[0]), .ZN(y[2]) );
  OR2_X1 U78bar ( .A1(bbar[2]), .A2(abar[0]), .ZN(ybar[2]);
  AND2_X1 U79 ( .A1(a[1]), .A2(b[13]), .ZN(y[29]) );
  OR2_X1 U79bar ( .A1(abar[1]), .A2(bbar[13]), .ZN(ybar[29]);
  AND2_X1 U80 ( .A1(a[1]), .A2(b[12]), .ZN(y[28]) );
  OR2_X1 U80bar ( .A1(abar[1]), .A2(bbar[12]), .ZN(ybar[28]);
  AND2_X1 U81 ( .A1(a[1]), .A2(b[11]), .ZN(y[27]) );
  OR2_X1 U81bar ( .A1(abar[1]), .A2(bbar[11]), .ZN(ybar[27]);
  AND2_X1 U82 ( .A1(a[1]), .A2(b[10]), .ZN(y[26]) );
  OR2_X1 U82bar ( .A1(abar[1]), .A2(bbar[10]), .ZN(ybar[26]);
  AND2_X1 U83 ( .A1(a[1]), .A2(b[9]), .ZN(y[25]) );
  OR2_X1 U83bar ( .A1(abar[1]), .A2(bbar[9]), .ZN(ybar[25]);
  AND2_X1 U84 ( .A1(a[15]), .A2(b[15]), .ZN(y[255]) );
  OR2_X1 U84bar ( .A1(abar[15]), .A2(bbar[15]), .ZN(ybar[255]);
  AND2_X1 U85 ( .A1(a[15]), .A2(b[14]), .ZN(y[254]) );
  OR2_X1 U85bar ( .A1(abar[15]), .A2(bbar[14]), .ZN(ybar[254]);
  AND2_X1 U86 ( .A1(a[15]), .A2(b[13]), .ZN(y[253]) );
  OR2_X1 U86bar ( .A1(abar[15]), .A2(bbar[13]), .ZN(ybar[253]);
  AND2_X1 U87 ( .A1(a[15]), .A2(b[12]), .ZN(y[252]) );
  OR2_X1 U87bar ( .A1(abar[15]), .A2(bbar[12]), .ZN(ybar[252]);
  AND2_X1 U88 ( .A1(a[15]), .A2(b[11]), .ZN(y[251]) );
  OR2_X1 U88bar ( .A1(abar[15]), .A2(bbar[11]), .ZN(ybar[251]);
  AND2_X1 U89 ( .A1(a[15]), .A2(b[10]), .ZN(y[250]) );
  OR2_X1 U89bar ( .A1(abar[15]), .A2(bbar[10]), .ZN(ybar[250]);
  AND2_X1 U90 ( .A1(a[1]), .A2(b[8]), .ZN(y[24]) );
  OR2_X1 U90bar ( .A1(abar[1]), .A2(bbar[8]), .ZN(ybar[24]);
  AND2_X1 U91 ( .A1(a[15]), .A2(b[9]), .ZN(y[249]) );
  OR2_X1 U91bar ( .A1(abar[15]), .A2(bbar[9]), .ZN(ybar[249]);
  AND2_X1 U92 ( .A1(a[15]), .A2(b[8]), .ZN(y[248]) );
  OR2_X1 U92bar ( .A1(abar[15]), .A2(bbar[8]), .ZN(ybar[248]);
  AND2_X1 U93 ( .A1(a[15]), .A2(b[7]), .ZN(y[247]) );
  OR2_X1 U93bar ( .A1(abar[15]), .A2(bbar[7]), .ZN(ybar[247]);
  AND2_X1 U94 ( .A1(a[15]), .A2(b[6]), .ZN(y[246]) );
  OR2_X1 U94bar ( .A1(abar[15]), .A2(bbar[6]), .ZN(ybar[246]);
  AND2_X1 U95 ( .A1(a[15]), .A2(b[5]), .ZN(y[245]) );
  OR2_X1 U95bar ( .A1(abar[15]), .A2(bbar[5]), .ZN(ybar[245]);
  AND2_X1 U96 ( .A1(a[15]), .A2(b[4]), .ZN(y[244]) );
  OR2_X1 U96bar ( .A1(abar[15]), .A2(bbar[4]), .ZN(ybar[244]);
  AND2_X1 U97 ( .A1(a[15]), .A2(b[3]), .ZN(y[243]) );
  OR2_X1 U97bar ( .A1(abar[15]), .A2(bbar[3]), .ZN(ybar[243]);
  AND2_X1 U98 ( .A1(a[15]), .A2(b[2]), .ZN(y[242]) );
  OR2_X1 U98bar ( .A1(abar[15]), .A2(bbar[2]), .ZN(ybar[242]);
  AND2_X1 U99 ( .A1(a[15]), .A2(b[1]), .ZN(y[241]) );
  OR2_X1 U99bar ( .A1(abar[15]), .A2(bbar[1]), .ZN(ybar[241]);
  AND2_X1 U100 ( .A1(a[15]), .A2(b[0]), .ZN(y[240]) );
  OR2_X1 U100bar ( .A1(abar[15]), .A2(bbar[0]), .ZN(ybar[240]);
  AND2_X1 U101 ( .A1(a[1]), .A2(b[7]), .ZN(y[23]) );
  OR2_X1 U101bar ( .A1(abar[1]), .A2(bbar[7]), .ZN(ybar[23]);
  AND2_X1 U102 ( .A1(a[14]), .A2(b[15]), .ZN(y[239]) );
  OR2_X1 U102bar ( .A1(abar[14]), .A2(bbar[15]), .ZN(ybar[239]);
  AND2_X1 U103 ( .A1(a[14]), .A2(b[14]), .ZN(y[238]) );
  OR2_X1 U103bar ( .A1(abar[14]), .A2(bbar[14]), .ZN(ybar[238]);
  AND2_X1 U104 ( .A1(a[14]), .A2(b[13]), .ZN(y[237]) );
  OR2_X1 U104bar ( .A1(abar[14]), .A2(bbar[13]), .ZN(ybar[237]);
  AND2_X1 U105 ( .A1(a[14]), .A2(b[12]), .ZN(y[236]) );
  OR2_X1 U105bar ( .A1(abar[14]), .A2(bbar[12]), .ZN(ybar[236]);
  AND2_X1 U106 ( .A1(a[14]), .A2(b[11]), .ZN(y[235]) );
  OR2_X1 U106bar ( .A1(abar[14]), .A2(bbar[11]), .ZN(ybar[235]);
  AND2_X1 U107 ( .A1(a[14]), .A2(b[10]), .ZN(y[234]) );
  OR2_X1 U107bar ( .A1(abar[14]), .A2(bbar[10]), .ZN(ybar[234]);
  AND2_X1 U108 ( .A1(a[14]), .A2(b[9]), .ZN(y[233]) );
  OR2_X1 U108bar ( .A1(abar[14]), .A2(bbar[9]), .ZN(ybar[233]);
  AND2_X1 U109 ( .A1(a[14]), .A2(b[8]), .ZN(y[232]) );
  OR2_X1 U109bar ( .A1(abar[14]), .A2(bbar[8]), .ZN(ybar[232]);
  AND2_X1 U110 ( .A1(a[14]), .A2(b[7]), .ZN(y[231]) );
  OR2_X1 U110bar ( .A1(abar[14]), .A2(bbar[7]), .ZN(ybar[231]);
  AND2_X1 U111 ( .A1(a[14]), .A2(b[6]), .ZN(y[230]) );
  OR2_X1 U111bar ( .A1(abar[14]), .A2(bbar[6]), .ZN(ybar[230]);
  AND2_X1 U112 ( .A1(a[1]), .A2(b[6]), .ZN(y[22]) );
  OR2_X1 U112bar ( .A1(abar[1]), .A2(bbar[6]), .ZN(ybar[22]);
  AND2_X1 U113 ( .A1(a[14]), .A2(b[5]), .ZN(y[229]) );
  OR2_X1 U113bar ( .A1(abar[14]), .A2(bbar[5]), .ZN(ybar[229]);
  AND2_X1 U114 ( .A1(a[14]), .A2(b[4]), .ZN(y[228]) );
  OR2_X1 U114bar ( .A1(abar[14]), .A2(bbar[4]), .ZN(ybar[228]);
  AND2_X1 U115 ( .A1(a[14]), .A2(b[3]), .ZN(y[227]) );
  OR2_X1 U115bar ( .A1(abar[14]), .A2(bbar[3]), .ZN(ybar[227]);
  AND2_X1 U116 ( .A1(a[14]), .A2(b[2]), .ZN(y[226]) );
  OR2_X1 U116bar ( .A1(abar[14]), .A2(bbar[2]), .ZN(ybar[226]);
  AND2_X1 U117 ( .A1(a[14]), .A2(b[1]), .ZN(y[225]) );
  OR2_X1 U117bar ( .A1(abar[14]), .A2(bbar[1]), .ZN(ybar[225]);
  AND2_X1 U118 ( .A1(a[14]), .A2(b[0]), .ZN(y[224]) );
  OR2_X1 U118bar ( .A1(abar[14]), .A2(bbar[0]), .ZN(ybar[224]);
  AND2_X1 U119 ( .A1(a[13]), .A2(b[15]), .ZN(y[223]) );
  OR2_X1 U119bar ( .A1(abar[13]), .A2(bbar[15]), .ZN(ybar[223]);
  AND2_X1 U120 ( .A1(a[13]), .A2(b[14]), .ZN(y[222]) );
  OR2_X1 U120bar ( .A1(abar[13]), .A2(bbar[14]), .ZN(ybar[222]);
  AND2_X1 U121 ( .A1(a[13]), .A2(b[13]), .ZN(y[221]) );
  OR2_X1 U121bar ( .A1(abar[13]), .A2(bbar[13]), .ZN(ybar[221]);
  AND2_X1 U122 ( .A1(a[13]), .A2(b[12]), .ZN(y[220]) );
  OR2_X1 U122bar ( .A1(abar[13]), .A2(bbar[12]), .ZN(ybar[220]);
  AND2_X1 U123 ( .A1(a[1]), .A2(b[5]), .ZN(y[21]) );
  OR2_X1 U123bar ( .A1(abar[1]), .A2(bbar[5]), .ZN(ybar[21]);
  AND2_X1 U124 ( .A1(a[13]), .A2(b[11]), .ZN(y[219]) );
  OR2_X1 U124bar ( .A1(abar[13]), .A2(bbar[11]), .ZN(ybar[219]);
  AND2_X1 U125 ( .A1(a[13]), .A2(b[10]), .ZN(y[218]) );
  OR2_X1 U125bar ( .A1(abar[13]), .A2(bbar[10]), .ZN(ybar[218]);
  AND2_X1 U126 ( .A1(a[13]), .A2(b[9]), .ZN(y[217]) );
  OR2_X1 U126bar ( .A1(abar[13]), .A2(bbar[9]), .ZN(ybar[217]);
  AND2_X1 U127 ( .A1(a[13]), .A2(b[8]), .ZN(y[216]) );
  OR2_X1 U127bar ( .A1(abar[13]), .A2(bbar[8]), .ZN(ybar[216]);
  AND2_X1 U128 ( .A1(a[13]), .A2(b[7]), .ZN(y[215]) );
  OR2_X1 U128bar ( .A1(abar[13]), .A2(bbar[7]), .ZN(ybar[215]);
  AND2_X1 U129 ( .A1(a[13]), .A2(b[6]), .ZN(y[214]) );
  OR2_X1 U129bar ( .A1(abar[13]), .A2(bbar[6]), .ZN(ybar[214]);
  AND2_X1 U130 ( .A1(a[13]), .A2(b[5]), .ZN(y[213]) );
  OR2_X1 U130bar ( .A1(abar[13]), .A2(bbar[5]), .ZN(ybar[213]);
  AND2_X1 U131 ( .A1(a[13]), .A2(b[4]), .ZN(y[212]) );
  OR2_X1 U131bar ( .A1(abar[13]), .A2(bbar[4]), .ZN(ybar[212]);
  AND2_X1 U132 ( .A1(a[13]), .A2(b[3]), .ZN(y[211]) );
  OR2_X1 U132bar ( .A1(abar[13]), .A2(bbar[3]), .ZN(ybar[211]);
  AND2_X1 U133 ( .A1(a[13]), .A2(b[2]), .ZN(y[210]) );
  OR2_X1 U133bar ( .A1(abar[13]), .A2(bbar[2]), .ZN(ybar[210]);
  AND2_X1 U134 ( .A1(a[1]), .A2(b[4]), .ZN(y[20]) );
  OR2_X1 U134bar ( .A1(abar[1]), .A2(bbar[4]), .ZN(ybar[20]);
  AND2_X1 U135 ( .A1(a[13]), .A2(b[1]), .ZN(y[209]) );
  OR2_X1 U135bar ( .A1(abar[13]), .A2(bbar[1]), .ZN(ybar[209]);
  AND2_X1 U136 ( .A1(a[13]), .A2(b[0]), .ZN(y[208]) );
  OR2_X1 U136bar ( .A1(abar[13]), .A2(bbar[0]), .ZN(ybar[208]);
  AND2_X1 U137 ( .A1(a[12]), .A2(b[15]), .ZN(y[207]) );
  OR2_X1 U137bar ( .A1(abar[12]), .A2(bbar[15]), .ZN(ybar[207]);
  AND2_X1 U138 ( .A1(a[12]), .A2(b[14]), .ZN(y[206]) );
  OR2_X1 U138bar ( .A1(abar[12]), .A2(bbar[14]), .ZN(ybar[206]);
  AND2_X1 U139 ( .A1(a[12]), .A2(b[13]), .ZN(y[205]) );
  OR2_X1 U139bar ( .A1(abar[12]), .A2(bbar[13]), .ZN(ybar[205]);
  AND2_X1 U140 ( .A1(a[12]), .A2(b[12]), .ZN(y[204]) );
  OR2_X1 U140bar ( .A1(abar[12]), .A2(bbar[12]), .ZN(ybar[204]);
  AND2_X1 U141 ( .A1(a[12]), .A2(b[11]), .ZN(y[203]) );
  OR2_X1 U141bar ( .A1(abar[12]), .A2(bbar[11]), .ZN(ybar[203]);
  AND2_X1 U142 ( .A1(a[12]), .A2(b[10]), .ZN(y[202]) );
  OR2_X1 U142bar ( .A1(abar[12]), .A2(bbar[10]), .ZN(ybar[202]);
  AND2_X1 U143 ( .A1(a[12]), .A2(b[9]), .ZN(y[201]) );
  OR2_X1 U143bar ( .A1(abar[12]), .A2(bbar[9]), .ZN(ybar[201]);
  AND2_X1 U144 ( .A1(a[12]), .A2(b[8]), .ZN(y[200]) );
  OR2_X1 U144bar ( .A1(abar[12]), .A2(bbar[8]), .ZN(ybar[200]);
  AND2_X1 U145 ( .A1(b[1]), .A2(a[0]), .ZN(y[1]) );
  OR2_X1 U145bar ( .A1(bbar[1]), .A2(abar[0]), .ZN(ybar[1]);
  AND2_X1 U146 ( .A1(a[1]), .A2(b[3]), .ZN(y[19]) );
  OR2_X1 U146bar ( .A1(abar[1]), .A2(bbar[3]), .ZN(ybar[19]);
  AND2_X1 U147 ( .A1(a[12]), .A2(b[7]), .ZN(y[199]) );
  OR2_X1 U147bar ( .A1(abar[12]), .A2(bbar[7]), .ZN(ybar[199]);
  AND2_X1 U148 ( .A1(a[12]), .A2(b[6]), .ZN(y[198]) );
  OR2_X1 U148bar ( .A1(abar[12]), .A2(bbar[6]), .ZN(ybar[198]);
  AND2_X1 U149 ( .A1(a[12]), .A2(b[5]), .ZN(y[197]) );
  OR2_X1 U149bar ( .A1(abar[12]), .A2(bbar[5]), .ZN(ybar[197]);
  AND2_X1 U150 ( .A1(a[12]), .A2(b[4]), .ZN(y[196]) );
  OR2_X1 U150bar ( .A1(abar[12]), .A2(bbar[4]), .ZN(ybar[196]);
  AND2_X1 U151 ( .A1(a[12]), .A2(b[3]), .ZN(y[195]) );
  OR2_X1 U151bar ( .A1(abar[12]), .A2(bbar[3]), .ZN(ybar[195]);
  AND2_X1 U152 ( .A1(a[12]), .A2(b[2]), .ZN(y[194]) );
  OR2_X1 U152bar ( .A1(abar[12]), .A2(bbar[2]), .ZN(ybar[194]);
  AND2_X1 U153 ( .A1(a[12]), .A2(b[1]), .ZN(y[193]) );
  OR2_X1 U153bar ( .A1(abar[12]), .A2(bbar[1]), .ZN(ybar[193]);
  AND2_X1 U154 ( .A1(a[12]), .A2(b[0]), .ZN(y[192]) );
  OR2_X1 U154bar ( .A1(abar[12]), .A2(bbar[0]), .ZN(ybar[192]);
  AND2_X1 U155 ( .A1(a[11]), .A2(b[15]), .ZN(y[191]) );
  OR2_X1 U155bar ( .A1(abar[11]), .A2(bbar[15]), .ZN(ybar[191]);
  AND2_X1 U156 ( .A1(a[11]), .A2(b[14]), .ZN(y[190]) );
  OR2_X1 U156bar ( .A1(abar[11]), .A2(bbar[14]), .ZN(ybar[190]);
  AND2_X1 U157 ( .A1(a[1]), .A2(b[2]), .ZN(y[18]) );
  OR2_X1 U157bar ( .A1(abar[1]), .A2(bbar[2]), .ZN(ybar[18]);
  AND2_X1 U158 ( .A1(a[11]), .A2(b[13]), .ZN(y[189]) );
  OR2_X1 U158bar ( .A1(abar[11]), .A2(bbar[13]), .ZN(ybar[189]);
  AND2_X1 U159 ( .A1(a[11]), .A2(b[12]), .ZN(y[188]) );
  OR2_X1 U159bar ( .A1(abar[11]), .A2(bbar[12]), .ZN(ybar[188]);
  AND2_X1 U160 ( .A1(a[11]), .A2(b[11]), .ZN(y[187]) );
  OR2_X1 U160bar ( .A1(abar[11]), .A2(bbar[11]), .ZN(ybar[187]);
  AND2_X1 U161 ( .A1(a[11]), .A2(b[10]), .ZN(y[186]) );
  OR2_X1 U161bar ( .A1(abar[11]), .A2(bbar[10]), .ZN(ybar[186]);
  AND2_X1 U162 ( .A1(a[11]), .A2(b[9]), .ZN(y[185]) );
  OR2_X1 U162bar ( .A1(abar[11]), .A2(bbar[9]), .ZN(ybar[185]);
  AND2_X1 U163 ( .A1(a[11]), .A2(b[8]), .ZN(y[184]) );
  OR2_X1 U163bar ( .A1(abar[11]), .A2(bbar[8]), .ZN(ybar[184]);
  AND2_X1 U164 ( .A1(a[11]), .A2(b[7]), .ZN(y[183]) );
  OR2_X1 U164bar ( .A1(abar[11]), .A2(bbar[7]), .ZN(ybar[183]);
  AND2_X1 U165 ( .A1(a[11]), .A2(b[6]), .ZN(y[182]) );
  OR2_X1 U165bar ( .A1(abar[11]), .A2(bbar[6]), .ZN(ybar[182]);
  AND2_X1 U166 ( .A1(a[11]), .A2(b[5]), .ZN(y[181]) );
  OR2_X1 U166bar ( .A1(abar[11]), .A2(bbar[5]), .ZN(ybar[181]);
  AND2_X1 U167 ( .A1(a[11]), .A2(b[4]), .ZN(y[180]) );
  OR2_X1 U167bar ( .A1(abar[11]), .A2(bbar[4]), .ZN(ybar[180]);
  AND2_X1 U168 ( .A1(a[1]), .A2(b[1]), .ZN(y[17]) );
  OR2_X1 U168bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[17]);
  AND2_X1 U169 ( .A1(a[11]), .A2(b[3]), .ZN(y[179]) );
  OR2_X1 U169bar ( .A1(abar[11]), .A2(bbar[3]), .ZN(ybar[179]);
  AND2_X1 U170 ( .A1(a[11]), .A2(b[2]), .ZN(y[178]) );
  OR2_X1 U170bar ( .A1(abar[11]), .A2(bbar[2]), .ZN(ybar[178]);
  AND2_X1 U171 ( .A1(a[11]), .A2(b[1]), .ZN(y[177]) );
  OR2_X1 U171bar ( .A1(abar[11]), .A2(bbar[1]), .ZN(ybar[177]);
  AND2_X1 U172 ( .A1(a[11]), .A2(b[0]), .ZN(y[176]) );
  OR2_X1 U172bar ( .A1(abar[11]), .A2(bbar[0]), .ZN(ybar[176]);
  AND2_X1 U173 ( .A1(a[10]), .A2(b[15]), .ZN(y[175]) );
  OR2_X1 U173bar ( .A1(abar[10]), .A2(bbar[15]), .ZN(ybar[175]);
  AND2_X1 U174 ( .A1(a[10]), .A2(b[14]), .ZN(y[174]) );
  OR2_X1 U174bar ( .A1(abar[10]), .A2(bbar[14]), .ZN(ybar[174]);
  AND2_X1 U175 ( .A1(a[10]), .A2(b[13]), .ZN(y[173]) );
  OR2_X1 U175bar ( .A1(abar[10]), .A2(bbar[13]), .ZN(ybar[173]);
  AND2_X1 U176 ( .A1(a[10]), .A2(b[12]), .ZN(y[172]) );
  OR2_X1 U176bar ( .A1(abar[10]), .A2(bbar[12]), .ZN(ybar[172]);
  AND2_X1 U177 ( .A1(a[10]), .A2(b[11]), .ZN(y[171]) );
  OR2_X1 U177bar ( .A1(abar[10]), .A2(bbar[11]), .ZN(ybar[171]);
  AND2_X1 U178 ( .A1(a[10]), .A2(b[10]), .ZN(y[170]) );
  OR2_X1 U178bar ( .A1(abar[10]), .A2(bbar[10]), .ZN(ybar[170]);
  AND2_X1 U179 ( .A1(a[1]), .A2(b[0]), .ZN(y[16]) );
  OR2_X1 U179bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[16]);
  AND2_X1 U180 ( .A1(a[10]), .A2(b[9]), .ZN(y[169]) );
  OR2_X1 U180bar ( .A1(abar[10]), .A2(bbar[9]), .ZN(ybar[169]);
  AND2_X1 U181 ( .A1(a[10]), .A2(b[8]), .ZN(y[168]) );
  OR2_X1 U181bar ( .A1(abar[10]), .A2(bbar[8]), .ZN(ybar[168]);
  AND2_X1 U182 ( .A1(a[10]), .A2(b[7]), .ZN(y[167]) );
  OR2_X1 U182bar ( .A1(abar[10]), .A2(bbar[7]), .ZN(ybar[167]);
  AND2_X1 U183 ( .A1(a[10]), .A2(b[6]), .ZN(y[166]) );
  OR2_X1 U183bar ( .A1(abar[10]), .A2(bbar[6]), .ZN(ybar[166]);
  AND2_X1 U184 ( .A1(a[10]), .A2(b[5]), .ZN(y[165]) );
  OR2_X1 U184bar ( .A1(abar[10]), .A2(bbar[5]), .ZN(ybar[165]);
  AND2_X1 U185 ( .A1(a[10]), .A2(b[4]), .ZN(y[164]) );
  OR2_X1 U185bar ( .A1(abar[10]), .A2(bbar[4]), .ZN(ybar[164]);
  AND2_X1 U186 ( .A1(a[10]), .A2(b[3]), .ZN(y[163]) );
  OR2_X1 U186bar ( .A1(abar[10]), .A2(bbar[3]), .ZN(ybar[163]);
  AND2_X1 U187 ( .A1(a[10]), .A2(b[2]), .ZN(y[162]) );
  OR2_X1 U187bar ( .A1(abar[10]), .A2(bbar[2]), .ZN(ybar[162]);
  AND2_X1 U188 ( .A1(a[10]), .A2(b[1]), .ZN(y[161]) );
  OR2_X1 U188bar ( .A1(abar[10]), .A2(bbar[1]), .ZN(ybar[161]);
  AND2_X1 U189 ( .A1(a[10]), .A2(b[0]), .ZN(y[160]) );
  OR2_X1 U189bar ( .A1(abar[10]), .A2(bbar[0]), .ZN(ybar[160]);
  AND2_X1 U190 ( .A1(b[15]), .A2(a[0]), .ZN(y[15]) );
  OR2_X1 U190bar ( .A1(bbar[15]), .A2(abar[0]), .ZN(ybar[15]);
  AND2_X1 U191 ( .A1(a[9]), .A2(b[15]), .ZN(y[159]) );
  OR2_X1 U191bar ( .A1(abar[9]), .A2(bbar[15]), .ZN(ybar[159]);
  AND2_X1 U192 ( .A1(a[9]), .A2(b[14]), .ZN(y[158]) );
  OR2_X1 U192bar ( .A1(abar[9]), .A2(bbar[14]), .ZN(ybar[158]);
  AND2_X1 U193 ( .A1(a[9]), .A2(b[13]), .ZN(y[157]) );
  OR2_X1 U193bar ( .A1(abar[9]), .A2(bbar[13]), .ZN(ybar[157]);
  AND2_X1 U194 ( .A1(a[9]), .A2(b[12]), .ZN(y[156]) );
  OR2_X1 U194bar ( .A1(abar[9]), .A2(bbar[12]), .ZN(ybar[156]);
  AND2_X1 U195 ( .A1(a[9]), .A2(b[11]), .ZN(y[155]) );
  OR2_X1 U195bar ( .A1(abar[9]), .A2(bbar[11]), .ZN(ybar[155]);
  AND2_X1 U196 ( .A1(a[9]), .A2(b[10]), .ZN(y[154]) );
  OR2_X1 U196bar ( .A1(abar[9]), .A2(bbar[10]), .ZN(ybar[154]);
  AND2_X1 U197 ( .A1(a[9]), .A2(b[9]), .ZN(y[153]) );
  OR2_X1 U197bar ( .A1(abar[9]), .A2(bbar[9]), .ZN(ybar[153]);
  AND2_X1 U198 ( .A1(a[9]), .A2(b[8]), .ZN(y[152]) );
  OR2_X1 U198bar ( .A1(abar[9]), .A2(bbar[8]), .ZN(ybar[152]);
  AND2_X1 U199 ( .A1(a[9]), .A2(b[7]), .ZN(y[151]) );
  OR2_X1 U199bar ( .A1(abar[9]), .A2(bbar[7]), .ZN(ybar[151]);
  AND2_X1 U200 ( .A1(a[9]), .A2(b[6]), .ZN(y[150]) );
  OR2_X1 U200bar ( .A1(abar[9]), .A2(bbar[6]), .ZN(ybar[150]);
  AND2_X1 U201 ( .A1(b[14]), .A2(a[0]), .ZN(y[14]) );
  OR2_X1 U201bar ( .A1(bbar[14]), .A2(abar[0]), .ZN(ybar[14]);
  AND2_X1 U202 ( .A1(a[9]), .A2(b[5]), .ZN(y[149]) );
  OR2_X1 U202bar ( .A1(abar[9]), .A2(bbar[5]), .ZN(ybar[149]);
  AND2_X1 U203 ( .A1(a[9]), .A2(b[4]), .ZN(y[148]) );
  OR2_X1 U203bar ( .A1(abar[9]), .A2(bbar[4]), .ZN(ybar[148]);
  AND2_X1 U204 ( .A1(a[9]), .A2(b[3]), .ZN(y[147]) );
  OR2_X1 U204bar ( .A1(abar[9]), .A2(bbar[3]), .ZN(ybar[147]);
  AND2_X1 U205 ( .A1(a[9]), .A2(b[2]), .ZN(y[146]) );
  OR2_X1 U205bar ( .A1(abar[9]), .A2(bbar[2]), .ZN(ybar[146]);
  AND2_X1 U206 ( .A1(a[9]), .A2(b[1]), .ZN(y[145]) );
  OR2_X1 U206bar ( .A1(abar[9]), .A2(bbar[1]), .ZN(ybar[145]);
  AND2_X1 U207 ( .A1(a[9]), .A2(b[0]), .ZN(y[144]) );
  OR2_X1 U207bar ( .A1(abar[9]), .A2(bbar[0]), .ZN(ybar[144]);
  AND2_X1 U208 ( .A1(a[8]), .A2(b[15]), .ZN(y[143]) );
  OR2_X1 U208bar ( .A1(abar[8]), .A2(bbar[15]), .ZN(ybar[143]);
  AND2_X1 U209 ( .A1(a[8]), .A2(b[14]), .ZN(y[142]) );
  OR2_X1 U209bar ( .A1(abar[8]), .A2(bbar[14]), .ZN(ybar[142]);
  AND2_X1 U210 ( .A1(a[8]), .A2(b[13]), .ZN(y[141]) );
  OR2_X1 U210bar ( .A1(abar[8]), .A2(bbar[13]), .ZN(ybar[141]);
  AND2_X1 U211 ( .A1(a[8]), .A2(b[12]), .ZN(y[140]) );
  OR2_X1 U211bar ( .A1(abar[8]), .A2(bbar[12]), .ZN(ybar[140]);
  AND2_X1 U212 ( .A1(b[13]), .A2(a[0]), .ZN(y[13]) );
  OR2_X1 U212bar ( .A1(bbar[13]), .A2(abar[0]), .ZN(ybar[13]);
  AND2_X1 U213 ( .A1(a[8]), .A2(b[11]), .ZN(y[139]) );
  OR2_X1 U213bar ( .A1(abar[8]), .A2(bbar[11]), .ZN(ybar[139]);
  AND2_X1 U214 ( .A1(a[8]), .A2(b[10]), .ZN(y[138]) );
  OR2_X1 U214bar ( .A1(abar[8]), .A2(bbar[10]), .ZN(ybar[138]);
  AND2_X1 U215 ( .A1(a[8]), .A2(b[9]), .ZN(y[137]) );
  OR2_X1 U215bar ( .A1(abar[8]), .A2(bbar[9]), .ZN(ybar[137]);
  AND2_X1 U216 ( .A1(a[8]), .A2(b[8]), .ZN(y[136]) );
  OR2_X1 U216bar ( .A1(abar[8]), .A2(bbar[8]), .ZN(ybar[136]);
  AND2_X1 U217 ( .A1(a[8]), .A2(b[7]), .ZN(y[135]) );
  OR2_X1 U217bar ( .A1(abar[8]), .A2(bbar[7]), .ZN(ybar[135]);
  AND2_X1 U218 ( .A1(a[8]), .A2(b[6]), .ZN(y[134]) );
  OR2_X1 U218bar ( .A1(abar[8]), .A2(bbar[6]), .ZN(ybar[134]);
  AND2_X1 U219 ( .A1(a[8]), .A2(b[5]), .ZN(y[133]) );
  OR2_X1 U219bar ( .A1(abar[8]), .A2(bbar[5]), .ZN(ybar[133]);
  AND2_X1 U220 ( .A1(a[8]), .A2(b[4]), .ZN(y[132]) );
  OR2_X1 U220bar ( .A1(abar[8]), .A2(bbar[4]), .ZN(ybar[132]);
  AND2_X1 U221 ( .A1(a[8]), .A2(b[3]), .ZN(y[131]) );
  OR2_X1 U221bar ( .A1(abar[8]), .A2(bbar[3]), .ZN(ybar[131]);
  AND2_X1 U222 ( .A1(a[8]), .A2(b[2]), .ZN(y[130]) );
  OR2_X1 U222bar ( .A1(abar[8]), .A2(bbar[2]), .ZN(ybar[130]);
  AND2_X1 U223 ( .A1(b[12]), .A2(a[0]), .ZN(y[12]) );
  OR2_X1 U223bar ( .A1(bbar[12]), .A2(abar[0]), .ZN(ybar[12]);
  AND2_X1 U224 ( .A1(a[8]), .A2(b[1]), .ZN(y[129]) );
  OR2_X1 U224bar ( .A1(abar[8]), .A2(bbar[1]), .ZN(ybar[129]);
  AND2_X1 U225 ( .A1(a[8]), .A2(b[0]), .ZN(y[128]) );
  OR2_X1 U225bar ( .A1(abar[8]), .A2(bbar[0]), .ZN(ybar[128]);
  AND2_X1 U226 ( .A1(a[7]), .A2(b[15]), .ZN(y[127]) );
  OR2_X1 U226bar ( .A1(abar[7]), .A2(bbar[15]), .ZN(ybar[127]);
  AND2_X1 U227 ( .A1(a[7]), .A2(b[14]), .ZN(y[126]) );
  OR2_X1 U227bar ( .A1(abar[7]), .A2(bbar[14]), .ZN(ybar[126]);
  AND2_X1 U228 ( .A1(a[7]), .A2(b[13]), .ZN(y[125]) );
  OR2_X1 U228bar ( .A1(abar[7]), .A2(bbar[13]), .ZN(ybar[125]);
  AND2_X1 U229 ( .A1(a[7]), .A2(b[12]), .ZN(y[124]) );
  OR2_X1 U229bar ( .A1(abar[7]), .A2(bbar[12]), .ZN(ybar[124]);
  AND2_X1 U230 ( .A1(a[7]), .A2(b[11]), .ZN(y[123]) );
  OR2_X1 U230bar ( .A1(abar[7]), .A2(bbar[11]), .ZN(ybar[123]);
  AND2_X1 U231 ( .A1(a[7]), .A2(b[10]), .ZN(y[122]) );
  OR2_X1 U231bar ( .A1(abar[7]), .A2(bbar[10]), .ZN(ybar[122]);
  AND2_X1 U232 ( .A1(a[7]), .A2(b[9]), .ZN(y[121]) );
  OR2_X1 U232bar ( .A1(abar[7]), .A2(bbar[9]), .ZN(ybar[121]);
  AND2_X1 U233 ( .A1(a[7]), .A2(b[8]), .ZN(y[120]) );
  OR2_X1 U233bar ( .A1(abar[7]), .A2(bbar[8]), .ZN(ybar[120]);
  AND2_X1 U234 ( .A1(b[11]), .A2(a[0]), .ZN(y[11]) );
  OR2_X1 U234bar ( .A1(bbar[11]), .A2(abar[0]), .ZN(ybar[11]);
  AND2_X1 U235 ( .A1(a[7]), .A2(b[7]), .ZN(y[119]) );
  OR2_X1 U235bar ( .A1(abar[7]), .A2(bbar[7]), .ZN(ybar[119]);
  AND2_X1 U236 ( .A1(a[7]), .A2(b[6]), .ZN(y[118]) );
  OR2_X1 U236bar ( .A1(abar[7]), .A2(bbar[6]), .ZN(ybar[118]);
  AND2_X1 U237 ( .A1(a[7]), .A2(b[5]), .ZN(y[117]) );
  OR2_X1 U237bar ( .A1(abar[7]), .A2(bbar[5]), .ZN(ybar[117]);
  AND2_X1 U238 ( .A1(a[7]), .A2(b[4]), .ZN(y[116]) );
  OR2_X1 U238bar ( .A1(abar[7]), .A2(bbar[4]), .ZN(ybar[116]);
  AND2_X1 U239 ( .A1(a[7]), .A2(b[3]), .ZN(y[115]) );
  OR2_X1 U239bar ( .A1(abar[7]), .A2(bbar[3]), .ZN(ybar[115]);
  AND2_X1 U240 ( .A1(a[7]), .A2(b[2]), .ZN(y[114]) );
  OR2_X1 U240bar ( .A1(abar[7]), .A2(bbar[2]), .ZN(ybar[114]);
  AND2_X1 U241 ( .A1(a[7]), .A2(b[1]), .ZN(y[113]) );
  OR2_X1 U241bar ( .A1(abar[7]), .A2(bbar[1]), .ZN(ybar[113]);
  AND2_X1 U242 ( .A1(a[7]), .A2(b[0]), .ZN(y[112]) );
  OR2_X1 U242bar ( .A1(abar[7]), .A2(bbar[0]), .ZN(ybar[112]);
  AND2_X1 U243 ( .A1(b[15]), .A2(a[6]), .ZN(y[111]) );
  OR2_X1 U243bar ( .A1(bbar[15]), .A2(abar[6]), .ZN(ybar[111]);
  AND2_X1 U244 ( .A1(b[14]), .A2(a[6]), .ZN(y[110]) );
  OR2_X1 U244bar ( .A1(bbar[14]), .A2(abar[6]), .ZN(ybar[110]);
  AND2_X1 U245 ( .A1(b[10]), .A2(a[0]), .ZN(y[10]) );
  OR2_X1 U245bar ( .A1(bbar[10]), .A2(abar[0]), .ZN(ybar[10]);
  AND2_X1 U246 ( .A1(b[13]), .A2(a[6]), .ZN(y[109]) );
  OR2_X1 U246bar ( .A1(bbar[13]), .A2(abar[6]), .ZN(ybar[109]);
  AND2_X1 U247 ( .A1(b[12]), .A2(a[6]), .ZN(y[108]) );
  OR2_X1 U247bar ( .A1(bbar[12]), .A2(abar[6]), .ZN(ybar[108]);
  AND2_X1 U248 ( .A1(b[11]), .A2(a[6]), .ZN(y[107]) );
  OR2_X1 U248bar ( .A1(bbar[11]), .A2(abar[6]), .ZN(ybar[107]);
  AND2_X1 U249 ( .A1(b[10]), .A2(a[6]), .ZN(y[106]) );
  OR2_X1 U249bar ( .A1(bbar[10]), .A2(abar[6]), .ZN(ybar[106]);
  AND2_X1 U250 ( .A1(a[6]), .A2(b[9]), .ZN(y[105]) );
  OR2_X1 U250bar ( .A1(abar[6]), .A2(bbar[9]), .ZN(ybar[105]);
  AND2_X1 U251 ( .A1(b[8]), .A2(a[6]), .ZN(y[104]) );
  OR2_X1 U251bar ( .A1(bbar[8]), .A2(abar[6]), .ZN(ybar[104]);
  AND2_X1 U252 ( .A1(b[7]), .A2(a[6]), .ZN(y[103]) );
  OR2_X1 U252bar ( .A1(bbar[7]), .A2(abar[6]), .ZN(ybar[103]);
  AND2_X1 U253 ( .A1(b[6]), .A2(a[6]), .ZN(y[102]) );
  OR2_X1 U253bar ( .A1(bbar[6]), .A2(abar[6]), .ZN(ybar[102]);
  AND2_X1 U254 ( .A1(b[5]), .A2(a[6]), .ZN(y[101]) );
  OR2_X1 U254bar ( .A1(bbar[5]), .A2(abar[6]), .ZN(ybar[101]);
  AND2_X1 U255 ( .A1(b[4]), .A2(a[6]), .ZN(y[100]) );
  OR2_X1 U255bar ( .A1(bbar[4]), .A2(abar[6]), .ZN(ybar[100]);
  AND2_X1 U256 ( .A1(b[0]), .A2(a[0]), .ZN(y[0]) );
  OR2_X1 U256bar ( .A1(bbar[0]), .A2(abar[0]), .ZN(ybar[0]);
endmodule




module CD2_77 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done

  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_78 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_79 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD4_39 ( a, b, y );
  input [3:0] a;
  input [3:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  //input_done

  output [15:0] y;
  reg [15:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]);
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]);
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]);
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]);
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]);
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]);
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]);
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]);
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]);
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]);
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]);
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]);
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]);
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]);
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]);
endmodule




module decode_0 ( in, out );
  input [7:0] in;
  //input_done

  output [255:0] out;
  //output_done

  wire   [15:0] level1;
  wire   [31:0] level2;
  //wire_done

  CD2_0 cd_l1_1 ( .a(in[1]), .b(in[0]), .y(level1[3:0]) );
  CD2_79 cd_l1_2 ( .a(in[3]), .b(in[2]), .y(level1[7:4]) );
  CD2_78 cd_l1_3 ( .a(in[5]), .b(in[4]), .y(level1[11:8]) );
  CD2_77 cd_l1_4 ( .a(in[7]), .b(in[6]), .y(level1[15:12]) );
  CD4_0 cd_l2_1 ( .a(level1[7:4]), .b(level1[3:0]), .y(level2[15:0]) );
  CD4_39 cd_l2_2 ( .a(level1[15:12]), .b(level1[11:8]), .y(level2[31:16]) );
  CD16_0 cd_l3 ( .a(level2[31:16]), .b(level2[15:0]), .y(out) );
endmodule


module encode_0 ( in, out );
  input [255:0] in;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
  assign inbar[8] = ~in[8];
  assign inbar[9] = ~in[9];
  assign inbar[10] = ~in[10];
  assign inbar[11] = ~in[11];
  assign inbar[12] = ~in[12];
  assign inbar[13] = ~in[13];
  assign inbar[14] = ~in[14];
  assign inbar[15] = ~in[15];
  assign inbar[16] = ~in[16];
  assign inbar[17] = ~in[17];
  assign inbar[18] = ~in[18];
  assign inbar[19] = ~in[19];
  assign inbar[20] = ~in[20];
  assign inbar[21] = ~in[21];
  assign inbar[22] = ~in[22];
  assign inbar[23] = ~in[23];
  assign inbar[24] = ~in[24];
  assign inbar[25] = ~in[25];
  assign inbar[26] = ~in[26];
  assign inbar[27] = ~in[27];
  assign inbar[28] = ~in[28];
  assign inbar[29] = ~in[29];
  assign inbar[30] = ~in[30];
  assign inbar[31] = ~in[31];
  assign inbar[32] = ~in[32];
  assign inbar[33] = ~in[33];
  assign inbar[34] = ~in[34];
  assign inbar[35] = ~in[35];
  assign inbar[36] = ~in[36];
  assign inbar[37] = ~in[37];
  assign inbar[38] = ~in[38];
  assign inbar[39] = ~in[39];
  assign inbar[40] = ~in[40];
  assign inbar[41] = ~in[41];
  assign inbar[42] = ~in[42];
  assign inbar[43] = ~in[43];
  assign inbar[44] = ~in[44];
  assign inbar[45] = ~in[45];
  assign inbar[46] = ~in[46];
  assign inbar[47] = ~in[47];
  assign inbar[48] = ~in[48];
  assign inbar[49] = ~in[49];
  assign inbar[50] = ~in[50];
  assign inbar[51] = ~in[51];
  assign inbar[52] = ~in[52];
  assign inbar[53] = ~in[53];
  assign inbar[54] = ~in[54];
  assign inbar[55] = ~in[55];
  assign inbar[56] = ~in[56];
  assign inbar[57] = ~in[57];
  assign inbar[58] = ~in[58];
  assign inbar[59] = ~in[59];
  assign inbar[60] = ~in[60];
  assign inbar[61] = ~in[61];
  assign inbar[62] = ~in[62];
  assign inbar[63] = ~in[63];
  assign inbar[64] = ~in[64];
  assign inbar[65] = ~in[65];
  assign inbar[66] = ~in[66];
  assign inbar[67] = ~in[67];
  assign inbar[68] = ~in[68];
  assign inbar[69] = ~in[69];
  assign inbar[70] = ~in[70];
  assign inbar[71] = ~in[71];
  assign inbar[72] = ~in[72];
  assign inbar[73] = ~in[73];
  assign inbar[74] = ~in[74];
  assign inbar[75] = ~in[75];
  assign inbar[76] = ~in[76];
  assign inbar[77] = ~in[77];
  assign inbar[78] = ~in[78];
  assign inbar[79] = ~in[79];
  assign inbar[80] = ~in[80];
  assign inbar[81] = ~in[81];
  assign inbar[82] = ~in[82];
  assign inbar[83] = ~in[83];
  assign inbar[84] = ~in[84];
  assign inbar[85] = ~in[85];
  assign inbar[86] = ~in[86];
  assign inbar[87] = ~in[87];
  assign inbar[88] = ~in[88];
  assign inbar[89] = ~in[89];
  assign inbar[90] = ~in[90];
  assign inbar[91] = ~in[91];
  assign inbar[92] = ~in[92];
  assign inbar[93] = ~in[93];
  assign inbar[94] = ~in[94];
  assign inbar[95] = ~in[95];
  assign inbar[96] = ~in[96];
  assign inbar[97] = ~in[97];
  assign inbar[98] = ~in[98];
  assign inbar[99] = ~in[99];
  assign inbar[100] = ~in[100];
  assign inbar[101] = ~in[101];
  assign inbar[102] = ~in[102];
  assign inbar[103] = ~in[103];
  assign inbar[104] = ~in[104];
  assign inbar[105] = ~in[105];
  assign inbar[106] = ~in[106];
  assign inbar[107] = ~in[107];
  assign inbar[108] = ~in[108];
  assign inbar[109] = ~in[109];
  assign inbar[110] = ~in[110];
  assign inbar[111] = ~in[111];
  assign inbar[112] = ~in[112];
  assign inbar[113] = ~in[113];
  assign inbar[114] = ~in[114];
  assign inbar[115] = ~in[115];
  assign inbar[116] = ~in[116];
  assign inbar[117] = ~in[117];
  assign inbar[118] = ~in[118];
  assign inbar[119] = ~in[119];
  assign inbar[120] = ~in[120];
  assign inbar[121] = ~in[121];
  assign inbar[122] = ~in[122];
  assign inbar[123] = ~in[123];
  assign inbar[124] = ~in[124];
  assign inbar[125] = ~in[125];
  assign inbar[126] = ~in[126];
  assign inbar[127] = ~in[127];
  assign inbar[128] = ~in[128];
  assign inbar[129] = ~in[129];
  assign inbar[130] = ~in[130];
  assign inbar[131] = ~in[131];
  assign inbar[132] = ~in[132];
  assign inbar[133] = ~in[133];
  assign inbar[134] = ~in[134];
  assign inbar[135] = ~in[135];
  assign inbar[136] = ~in[136];
  assign inbar[137] = ~in[137];
  assign inbar[138] = ~in[138];
  assign inbar[139] = ~in[139];
  assign inbar[140] = ~in[140];
  assign inbar[141] = ~in[141];
  assign inbar[142] = ~in[142];
  assign inbar[143] = ~in[143];
  assign inbar[144] = ~in[144];
  assign inbar[145] = ~in[145];
  assign inbar[146] = ~in[146];
  assign inbar[147] = ~in[147];
  assign inbar[148] = ~in[148];
  assign inbar[149] = ~in[149];
  assign inbar[150] = ~in[150];
  assign inbar[151] = ~in[151];
  assign inbar[152] = ~in[152];
  assign inbar[153] = ~in[153];
  assign inbar[154] = ~in[154];
  assign inbar[155] = ~in[155];
  assign inbar[156] = ~in[156];
  assign inbar[157] = ~in[157];
  assign inbar[158] = ~in[158];
  assign inbar[159] = ~in[159];
  assign inbar[160] = ~in[160];
  assign inbar[161] = ~in[161];
  assign inbar[162] = ~in[162];
  assign inbar[163] = ~in[163];
  assign inbar[164] = ~in[164];
  assign inbar[165] = ~in[165];
  assign inbar[166] = ~in[166];
  assign inbar[167] = ~in[167];
  assign inbar[168] = ~in[168];
  assign inbar[169] = ~in[169];
  assign inbar[170] = ~in[170];
  assign inbar[171] = ~in[171];
  assign inbar[172] = ~in[172];
  assign inbar[173] = ~in[173];
  assign inbar[174] = ~in[174];
  assign inbar[175] = ~in[175];
  assign inbar[176] = ~in[176];
  assign inbar[177] = ~in[177];
  assign inbar[178] = ~in[178];
  assign inbar[179] = ~in[179];
  assign inbar[180] = ~in[180];
  assign inbar[181] = ~in[181];
  assign inbar[182] = ~in[182];
  assign inbar[183] = ~in[183];
  assign inbar[184] = ~in[184];
  assign inbar[185] = ~in[185];
  assign inbar[186] = ~in[186];
  assign inbar[187] = ~in[187];
  assign inbar[188] = ~in[188];
  assign inbar[189] = ~in[189];
  assign inbar[190] = ~in[190];
  assign inbar[191] = ~in[191];
  assign inbar[192] = ~in[192];
  assign inbar[193] = ~in[193];
  assign inbar[194] = ~in[194];
  assign inbar[195] = ~in[195];
  assign inbar[196] = ~in[196];
  assign inbar[197] = ~in[197];
  assign inbar[198] = ~in[198];
  assign inbar[199] = ~in[199];
  assign inbar[200] = ~in[200];
  assign inbar[201] = ~in[201];
  assign inbar[202] = ~in[202];
  assign inbar[203] = ~in[203];
  assign inbar[204] = ~in[204];
  assign inbar[205] = ~in[205];
  assign inbar[206] = ~in[206];
  assign inbar[207] = ~in[207];
  assign inbar[208] = ~in[208];
  assign inbar[209] = ~in[209];
  assign inbar[210] = ~in[210];
  assign inbar[211] = ~in[211];
  assign inbar[212] = ~in[212];
  assign inbar[213] = ~in[213];
  assign inbar[214] = ~in[214];
  assign inbar[215] = ~in[215];
  assign inbar[216] = ~in[216];
  assign inbar[217] = ~in[217];
  assign inbar[218] = ~in[218];
  assign inbar[219] = ~in[219];
  assign inbar[220] = ~in[220];
  assign inbar[221] = ~in[221];
  assign inbar[222] = ~in[222];
  assign inbar[223] = ~in[223];
  assign inbar[224] = ~in[224];
  assign inbar[225] = ~in[225];
  assign inbar[226] = ~in[226];
  assign inbar[227] = ~in[227];
  assign inbar[228] = ~in[228];
  assign inbar[229] = ~in[229];
  assign inbar[230] = ~in[230];
  assign inbar[231] = ~in[231];
  assign inbar[232] = ~in[232];
  assign inbar[233] = ~in[233];
  assign inbar[234] = ~in[234];
  assign inbar[235] = ~in[235];
  assign inbar[236] = ~in[236];
  assign inbar[237] = ~in[237];
  assign inbar[238] = ~in[238];
  assign inbar[239] = ~in[239];
  assign inbar[240] = ~in[240];
  assign inbar[241] = ~in[241];
  assign inbar[242] = ~in[242];
  assign inbar[243] = ~in[243];
  assign inbar[244] = ~in[244];
  assign inbar[245] = ~in[245];
  assign inbar[246] = ~in[246];
  assign inbar[247] = ~in[247];
  assign inbar[248] = ~in[248];
  assign inbar[249] = ~in[249];
  assign inbar[250] = ~in[250];
  assign inbar[251] = ~in[251];
  assign inbar[252] = ~in[252];
  assign inbar[253] = ~in[253];
  assign inbar[254] = ~in[254];
  assign inbar[255] = ~in[255];
  //input_done

  output [7:0] out;
  reg [7:0] outbar;
  //output_done

  wire   in_81, in_80, in_79, in_78, in_77, in_76, in_75, in_74, in_73, in_72,
         in_71, in_70, in_69, in_68, in_67, in_66, in_65, in_64, in_63, in_62,
         in_61, in_60, in_59, in_58, in_57, in_56, in_55, in_54, in_53, in_52,
         in_51, in_50, in_49, in_48, in_47, in_46, in_45, in_44, in_43, in_42,
         in_41, in_40, in_39, in_38, in_37, in_36, in_35, in_34, in_33, in_32,
         in_31, in_30, in_29, in_28, in_27, in_26, in_25, in_24, in_23, in_22,
         in_21, in_20, in_19, in_18, in_17, in_16, in_15, in_14, in_13, in_12,
         in_11, in_10, in_9, in_8, in_7, in_6, in_5, in_4, in_3, in_2, in_1,
         in_0, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486;
  wire in_81bar, in_80bar, in_79bar, in_78bar, in_77bar, in_76bar, in_75bar, in_74bar, in_73bar, in_72bar, in_71bar, in_70bar, in_69bar, in_68bar, in_67bar, in_66bar, in_65bar, in_64bar, in_63bar, in_62bar, in_61bar, in_60bar, in_59bar, in_58bar, in_57bar, in_56bar, in_55bar, in_54bar, in_53bar, in_52bar, in_51bar, in_50bar, in_49bar, in_48bar, in_47bar, in_46bar, in_45bar, in_44bar, in_43bar, in_42bar, in_41bar, in_40bar, in_39bar, in_38bar, in_37bar, in_36bar, in_35bar, in_34bar, in_33bar, in_32bar, in_31bar, in_30bar, in_29bar, in_28bar, in_27bar, in_26bar, in_25bar, in_24bar, in_23bar, in_22bar, in_21bar, in_20bar, in_19bar, in_18bar, in_17bar, in_16bar, in_15bar, in_14bar, in_13bar, in_12bar, in_11bar, in_10bar, in_9bar, in_8bar, in_7bar, in_6bar, in_5bar, in_4bar, in_3bar, in_2bar, in_1bar, in_0bar, n1bar, n2bar, n3bar, n4bar, n5bar, n6bar, n7bar, n8bar, n9bar, n10bar, n11bar, n12bar, n13bar, n14bar, n15bar, n16bar, n17bar, n18bar, n19bar, n20bar, n21bar, n22bar, n23bar, n24bar, n25bar, n26bar, n27bar, n28bar, n29bar, n30bar, n31bar, n32bar, n33bar, n34bar, n35bar, n36bar, n37bar, n38bar, n39bar, n40bar, n41bar, n42bar, n43bar, n44bar, n45bar, n46bar, n47bar, n48bar, n49bar, n50bar, n51bar, n52bar, n53bar, n54bar, n55bar, n56bar, n57bar, n58bar, n59bar, n60bar, n61bar, n62bar, n63bar, n64bar, n65bar, n66bar, n67bar, n68bar, n69bar, n70bar, n71bar, n72bar, n73bar, n74bar, n75bar, n76bar, n77bar, n78bar, n79bar, n80bar, n81bar, n82bar, n83bar, n84bar, n85bar, n86bar, n87bar, n88bar, n89bar, n90bar, n91bar, n92bar, n93bar, n94bar, n95bar, n96bar, n97bar, n98bar, n99bar, n100bar, n101bar, n102bar, n103bar, n104bar, n105bar, n106bar, n107bar, n108bar, n109bar, n110bar, n111bar, n112bar, n113bar, n114bar, n115bar, n116bar, n117bar, n118bar, n119bar, n120bar, n121bar, n122bar, n123bar, n124bar, n125bar, n126bar, n127bar, n128bar, n129bar, n130bar, n131bar, n132bar, n133bar, n134bar, n135bar, n136bar, n137bar, n138bar, n139bar, n140bar, n141bar, n142bar, n143bar, n144bar, n145bar, n146bar, n147bar, n148bar, n149bar, n150bar, n151bar, n152bar, n153bar, n154bar, n155bar, n156bar, n157bar, n158bar, n159bar, n160bar, n161bar, n162bar, n163bar, n164bar, n165bar, n166bar, n167bar, n168bar, n169bar, n170bar, n171bar, n172bar, n173bar, n174bar, n175bar, n176bar, n177bar, n178bar, n179bar, n180bar, n181bar, n182bar, n183bar, n184bar, n185bar, n186bar, n187bar, n188bar, n189bar, n190bar, n191bar, n192bar, n193bar, n194bar, n195bar, n196bar, n197bar, n198bar, n199bar, n200bar, n201bar, n202bar, n203bar, n204bar, n205bar, n206bar, n207bar, n208bar, n209bar, n210bar, n211bar, n212bar, n213bar, n214bar, n215bar, n216bar, n217bar, n218bar, n219bar, n220bar, n221bar, n222bar, n223bar, n224bar, n225bar, n226bar, n227bar, n228bar, n229bar, n230bar, n231bar, n232bar, n233bar, n234bar, n235bar, n236bar, n237bar, n238bar, n239bar, n240bar, n241bar, n242bar, n243bar, n244bar, n245bar, n246bar, n247bar, n248bar, n249bar, n250bar, n251bar, n252bar, n253bar, n254bar, n255bar, n256bar, n257bar, n258bar, n259bar, n260bar, n261bar, n262bar, n263bar, n264bar, n265bar, n266bar, n267bar, n268bar, n269bar, n270bar, n271bar, n272bar, n273bar, n274bar, n275bar, n276bar, n277bar, n278bar, n279bar, n280bar, n281bar, n282bar, n283bar, n284bar, n285bar, n286bar, n287bar, n288bar, n289bar, n290bar, n291bar, n292bar, n293bar, n294bar, n295bar, n296bar, n297bar, n298bar, n299bar, n300bar, n301bar, n302bar, n303bar, n304bar, n305bar, n306bar, n307bar, n308bar, n309bar, n310bar, n311bar, n312bar, n313bar, n314bar, n315bar, n316bar, n317bar, n318bar, n319bar, n320bar, n321bar, n322bar, n323bar, n324bar, n325bar, n326bar, n327bar, n328bar, n329bar, n330bar, n331bar, n332bar, n333bar, n334bar, n335bar, n336bar, n337bar, n338bar, n339bar, n340bar, n341bar, n342bar, n343bar, n344bar, n345bar, n346bar, n347bar, n348bar, n349bar, n350bar, n351bar, n352bar, n353bar, n354bar, n355bar, n356bar, n357bar, n358bar, n359bar, n360bar, n361bar, n362bar, n363bar, n364bar, n365bar, n366bar, n367bar, n368bar, n369bar, n370bar, n371bar, n372bar, n373bar, n374bar, n375bar, n376bar, n377bar, n378bar, n379bar, n380bar, n381bar, n382bar, n383bar, n384bar, n385bar, n386bar, n387bar, n388bar, n389bar, n390bar, n391bar, n392bar, n393bar, n394bar, n395bar, n396bar, n397bar, n398bar, n399bar, n400bar, n401bar, n402bar, n403bar, n404bar, n405bar, n406bar, n407bar, n408bar, n409bar, n410bar, n411bar, n412bar, n413bar, n414bar, n415bar, n416bar, n417bar, n418bar, n419bar, n420bar, n421bar, n422bar, n423bar, n424bar, n425bar, n426bar, n427bar, n428bar, n429bar, n430bar, n431bar, n432bar, n433bar, n434bar, n435bar, n436bar, n437bar, n438bar, n439bar, n440bar, n441bar, n442bar, n443bar, n444bar, n445bar, n446bar, n447bar, n448bar, n449bar, n450bar, n451bar, n452bar, n453bar, n454bar, n455bar, n456bar, n457bar, n458bar, n459bar, n460bar, n461bar, n462bar, n463bar, n464bar, n465bar, n466bar, n467bar, n468bar, n469bar, n470bar, n471bar, n472bar, n473bar, n474bar, n475bar, n476bar, n477bar, n478bar, n479bar, n480bar, n481bar, n482bar, n483bar, n484bar, n485bar, n486bar;
  //wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];

  OR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(out[7]) );
  AND2_X1 U1bar ( .A1(n1bar), .A2(n2bar), .ZN(outbar[7]);
  OR2_X1 U2 ( .A1(n3), .A2(n4), .ZN(n2) );
  AND2_X1 U2bar ( .A1(n3bar), .A2(n4bar), .ZN(n2bar);
  OR2_X1 U3 ( .A1(n5), .A2(n6), .ZN(n4) );
  AND2_X1 U3bar ( .A1(n5bar), .A2(n6bar), .ZN(n4bar);
  OR2_X1 U4 ( .A1(n7), .A2(n8), .ZN(n6) );
  AND2_X1 U4bar ( .A1(n7bar), .A2(n8bar), .ZN(n6bar);
  OR2_X1 U5 ( .A1(n9), .A2(n10), .ZN(n5) );
  AND2_X1 U5bar ( .A1(n9bar), .A2(n10bar), .ZN(n5bar);
  OR2_X1 U6 ( .A1(in[116]), .A2(n11), .ZN(n10) );
  AND2_X1 U6bar ( .A1(inbar[116]), .A2(n11bar), .ZN(n10bar);
  OR2_X1 U7 ( .A1(n12), .A2(n13), .ZN(n3) );
  AND2_X1 U7bar ( .A1(n12bar), .A2(n13bar), .ZN(n3bar);
  OR2_X1 U8 ( .A1(in[150]), .A2(in[127]), .ZN(n13) );
  AND2_X1 U8bar ( .A1(inbar[150]), .A2(inbar[127]), .ZN(n13bar);
  OR2_X1 U9 ( .A1(in[160]), .A2(n14), .ZN(n12) );
  AND2_X1 U9bar ( .A1(inbar[160]), .A2(n14bar), .ZN(n12bar);
  OR2_X1 U10 ( .A1(in[252]), .A2(in[168]), .ZN(n14) );
  AND2_X1 U10bar ( .A1(inbar[252]), .A2(inbar[168]), .ZN(n14bar);
  OR2_X1 U11 ( .A1(n15), .A2(n16), .ZN(n1) );
  AND2_X1 U11bar ( .A1(n15bar), .A2(n16bar), .ZN(n1bar);
  OR2_X1 U12 ( .A1(n17), .A2(n18), .ZN(n16) );
  AND2_X1 U12bar ( .A1(n17bar), .A2(n18bar), .ZN(n16bar);
  OR2_X1 U13 ( .A1(in_17), .A2(in[96]), .ZN(n18) );
  AND2_X1 U13bar ( .A1(in_17bar), .A2(inbar[96]), .ZN(n18bar);
  OR2_X1 U14 ( .A1(in_23), .A2(n19), .ZN(n17) );
  AND2_X1 U14bar ( .A1(in_23bar), .A2(n19bar), .ZN(n17bar);
  OR2_X1 U15 ( .A1(in_31), .A2(in_26), .ZN(n19) );
  AND2_X1 U15bar ( .A1(in_31bar), .A2(in_26bar), .ZN(n19bar);
  OR2_X1 U16 ( .A1(n20), .A2(n21), .ZN(n15) );
  AND2_X1 U16bar ( .A1(n20bar), .A2(n21bar), .ZN(n15bar);
  OR2_X1 U17 ( .A1(in_58), .A2(in_4), .ZN(n21) );
  AND2_X1 U17bar ( .A1(in_58bar), .A2(in_4bar), .ZN(n21bar);
  OR2_X1 U18 ( .A1(in_59), .A2(n22), .ZN(n20) );
  AND2_X1 U18bar ( .A1(in_59bar), .A2(n22bar), .ZN(n20bar);
  OR2_X1 U19 ( .A1(in_71), .A2(in_62), .ZN(n22) );
  AND2_X1 U19bar ( .A1(in_71bar), .A2(in_62bar), .ZN(n22bar);
  OR2_X1 U20 ( .A1(n23), .A2(n24), .ZN(out[6]) );
  AND2_X1 U20bar ( .A1(n23bar), .A2(n24bar), .ZN(outbar[6]);
  OR2_X1 U21 ( .A1(n25), .A2(n26), .ZN(n24) );
  AND2_X1 U21bar ( .A1(n25bar), .A2(n26bar), .ZN(n24bar);
  OR2_X1 U22 ( .A1(n27), .A2(n28), .ZN(n26) );
  AND2_X1 U22bar ( .A1(n27bar), .A2(n28bar), .ZN(n26bar);
  OR2_X1 U23 ( .A1(n29), .A2(n30), .ZN(n28) );
  AND2_X1 U23bar ( .A1(n29bar), .A2(n30bar), .ZN(n28bar);
  OR2_X1 U24 ( .A1(n31), .A2(n32), .ZN(n27) );
  AND2_X1 U24bar ( .A1(n31bar), .A2(n32bar), .ZN(n27bar);
  OR2_X1 U25 ( .A1(in[101]), .A2(n33), .ZN(n32) );
  AND2_X1 U25bar ( .A1(inbar[101]), .A2(n33bar), .ZN(n32bar);
  OR2_X1 U26 ( .A1(n34), .A2(n35), .ZN(n25) );
  AND2_X1 U26bar ( .A1(n34bar), .A2(n35bar), .ZN(n25bar);
  OR2_X1 U27 ( .A1(in[114]), .A2(in[104]), .ZN(n35) );
  AND2_X1 U27bar ( .A1(inbar[114]), .A2(inbar[104]), .ZN(n35bar);
  OR2_X1 U28 ( .A1(in[128]), .A2(n36), .ZN(n34) );
  AND2_X1 U28bar ( .A1(inbar[128]), .A2(n36bar), .ZN(n34bar);
  OR2_X1 U29 ( .A1(in[136]), .A2(in[134]), .ZN(n36) );
  AND2_X1 U29bar ( .A1(inbar[136]), .A2(inbar[134]), .ZN(n36bar);
  OR2_X1 U30 ( .A1(n37), .A2(n38), .ZN(n23) );
  AND2_X1 U30bar ( .A1(n37bar), .A2(n38bar), .ZN(n23bar);
  OR2_X1 U31 ( .A1(n39), .A2(n40), .ZN(n38) );
  AND2_X1 U31bar ( .A1(n39bar), .A2(n40bar), .ZN(n38bar);
  OR2_X1 U32 ( .A1(in[177]), .A2(in[164]), .ZN(n40) );
  AND2_X1 U32bar ( .A1(inbar[177]), .A2(inbar[164]), .ZN(n40bar);
  OR2_X1 U33 ( .A1(in[212]), .A2(n41), .ZN(n39) );
  AND2_X1 U33bar ( .A1(inbar[212]), .A2(n41bar), .ZN(n39bar);
  OR2_X1 U34 ( .A1(in[248]), .A2(in[221]), .ZN(n41) );
  AND2_X1 U34bar ( .A1(inbar[248]), .A2(inbar[221]), .ZN(n41bar);
  OR2_X1 U35 ( .A1(n42), .A2(n43), .ZN(n37) );
  AND2_X1 U35bar ( .A1(n42bar), .A2(n43bar), .ZN(n37bar);
  OR2_X1 U36 ( .A1(in_18), .A2(in[93]), .ZN(n43) );
  AND2_X1 U36bar ( .A1(in_18bar), .A2(inbar[93]), .ZN(n43bar);
  OR2_X1 U37 ( .A1(in_31), .A2(n44), .ZN(n42) );
  AND2_X1 U37bar ( .A1(in_31bar), .A2(n44bar), .ZN(n42bar);
  OR2_X1 U38 ( .A1(in_7), .A2(in_39), .ZN(n44) );
  AND2_X1 U38bar ( .A1(in_7bar), .A2(in_39bar), .ZN(n44bar);
  OR2_X1 U39 ( .A1(n45), .A2(n46), .ZN(out[5]) );
  AND2_X1 U39bar ( .A1(n45bar), .A2(n46bar), .ZN(outbar[5]);
  OR2_X1 U40 ( .A1(n47), .A2(n48), .ZN(n46) );
  AND2_X1 U40bar ( .A1(n47bar), .A2(n48bar), .ZN(n46bar);
  OR2_X1 U41 ( .A1(n49), .A2(n50), .ZN(n48) );
  AND2_X1 U41bar ( .A1(n49bar), .A2(n50bar), .ZN(n48bar);
  OR2_X1 U42 ( .A1(n51), .A2(n52), .ZN(n50) );
  AND2_X1 U42bar ( .A1(n51bar), .A2(n52bar), .ZN(n50bar);
  OR2_X1 U43 ( .A1(n33), .A2(n53), .ZN(n49) );
  AND2_X1 U43bar ( .A1(n33bar), .A2(n53bar), .ZN(n49bar);
  OR2_X1 U44 ( .A1(in[111]), .A2(n54), .ZN(n53) );
  AND2_X1 U44bar ( .A1(inbar[111]), .A2(n54bar), .ZN(n53bar);
  OR2_X1 U45 ( .A1(n55), .A2(n56), .ZN(n33) );
  AND2_X1 U45bar ( .A1(n55bar), .A2(n56bar), .ZN(n33bar);
  OR2_X1 U46 ( .A1(n57), .A2(n58), .ZN(n56) );
  AND2_X1 U46bar ( .A1(n57bar), .A2(n58bar), .ZN(n56bar);
  OR2_X1 U47 ( .A1(n59), .A2(n60), .ZN(n58) );
  AND2_X1 U47bar ( .A1(n59bar), .A2(n60bar), .ZN(n58bar);
  OR2_X1 U48 ( .A1(in[140]), .A2(in[131]), .ZN(n60) );
  AND2_X1 U48bar ( .A1(inbar[140]), .A2(inbar[131]), .ZN(n60bar);
  OR2_X1 U49 ( .A1(in[160]), .A2(in[144]), .ZN(n59) );
  AND2_X1 U49bar ( .A1(inbar[160]), .A2(inbar[144]), .ZN(n59bar);
  OR2_X1 U50 ( .A1(n61), .A2(n62), .ZN(n57) );
  AND2_X1 U50bar ( .A1(n61bar), .A2(n62bar), .ZN(n57bar);
  OR2_X1 U51 ( .A1(in[179]), .A2(in[174]), .ZN(n62) );
  AND2_X1 U51bar ( .A1(inbar[179]), .A2(inbar[174]), .ZN(n62bar);
  OR2_X1 U52 ( .A1(in[188]), .A2(in[184]), .ZN(n61) );
  AND2_X1 U52bar ( .A1(inbar[188]), .A2(inbar[184]), .ZN(n61bar);
  OR2_X1 U53 ( .A1(n63), .A2(n64), .ZN(n55) );
  AND2_X1 U53bar ( .A1(n63bar), .A2(n64bar), .ZN(n55bar);
  OR2_X1 U54 ( .A1(n65), .A2(n66), .ZN(n64) );
  AND2_X1 U54bar ( .A1(n65bar), .A2(n66bar), .ZN(n64bar);
  OR2_X1 U55 ( .A1(in[216]), .A2(in[200]), .ZN(n66) );
  AND2_X1 U55bar ( .A1(inbar[216]), .A2(inbar[200]), .ZN(n66bar);
  OR2_X1 U56 ( .A1(in[228]), .A2(in[224]), .ZN(n65) );
  AND2_X1 U56bar ( .A1(inbar[228]), .A2(inbar[224]), .ZN(n65bar);
  OR2_X1 U57 ( .A1(n67), .A2(n68), .ZN(n63) );
  AND2_X1 U57bar ( .A1(n67bar), .A2(n68bar), .ZN(n63bar);
  OR2_X1 U58 ( .A1(in[247]), .A2(in[235]), .ZN(n68) );
  AND2_X1 U58bar ( .A1(inbar[247]), .A2(inbar[235]), .ZN(n68bar);
  OR2_X1 U59 ( .A1(in_42), .A2(in[83]), .ZN(n67) );
  AND2_X1 U59bar ( .A1(in_42bar), .A2(inbar[83]), .ZN(n67bar);
  OR2_X1 U60 ( .A1(n69), .A2(n70), .ZN(n47) );
  AND2_X1 U60bar ( .A1(n69bar), .A2(n70bar), .ZN(n47bar);
  OR2_X1 U61 ( .A1(in[166]), .A2(in[123]), .ZN(n70) );
  AND2_X1 U61bar ( .A1(inbar[166]), .A2(inbar[123]), .ZN(n70bar);
  OR2_X1 U62 ( .A1(in[170]), .A2(n71), .ZN(n69) );
  AND2_X1 U62bar ( .A1(inbar[170]), .A2(n71bar), .ZN(n69bar);
  OR2_X1 U63 ( .A1(in[194]), .A2(in[183]), .ZN(n71) );
  AND2_X1 U63bar ( .A1(inbar[194]), .A2(inbar[183]), .ZN(n71bar);
  OR2_X1 U64 ( .A1(n72), .A2(n73), .ZN(n45) );
  AND2_X1 U64bar ( .A1(n72bar), .A2(n73bar), .ZN(n45bar);
  OR2_X1 U65 ( .A1(n74), .A2(n75), .ZN(n73) );
  AND2_X1 U65bar ( .A1(n74bar), .A2(n75bar), .ZN(n73bar);
  OR2_X1 U66 ( .A1(in[241]), .A2(in[238]), .ZN(n75) );
  AND2_X1 U66bar ( .A1(inbar[241]), .A2(inbar[238]), .ZN(n75bar);
  OR2_X1 U67 ( .A1(in[250]), .A2(n76), .ZN(n74) );
  AND2_X1 U67bar ( .A1(inbar[250]), .A2(n76bar), .ZN(n74bar);
  OR2_X1 U68 ( .A1(in_24), .A2(in[84]), .ZN(n76) );
  AND2_X1 U68bar ( .A1(in_24bar), .A2(inbar[84]), .ZN(n76bar);
  OR2_X1 U69 ( .A1(n77), .A2(n78), .ZN(n72) );
  AND2_X1 U69bar ( .A1(n77bar), .A2(n78bar), .ZN(n72bar);
  OR2_X1 U70 ( .A1(in_41), .A2(in_29), .ZN(n78) );
  AND2_X1 U70bar ( .A1(in_41bar), .A2(in_29bar), .ZN(n78bar);
  OR2_X1 U71 ( .A1(in_66), .A2(n79), .ZN(n77) );
  AND2_X1 U71bar ( .A1(in_66bar), .A2(n79bar), .ZN(n77bar);
  OR2_X1 U72 ( .A1(in_76), .A2(in_71), .ZN(n79) );
  AND2_X1 U72bar ( .A1(in_76bar), .A2(in_71bar), .ZN(n79bar);
  OR2_X1 U73 ( .A1(n80), .A2(n81), .ZN(out[4]) );
  AND2_X1 U73bar ( .A1(n80bar), .A2(n81bar), .ZN(outbar[4]);
  OR2_X1 U74 ( .A1(n82), .A2(n83), .ZN(n81) );
  AND2_X1 U74bar ( .A1(n82bar), .A2(n83bar), .ZN(n81bar);
  OR2_X1 U75 ( .A1(n84), .A2(n85), .ZN(n83) );
  AND2_X1 U75bar ( .A1(n84bar), .A2(n85bar), .ZN(n83bar);
  OR2_X1 U76 ( .A1(n51), .A2(n86), .ZN(n85) );
  AND2_X1 U76bar ( .A1(n51bar), .A2(n86bar), .ZN(n85bar);
  OR2_X1 U77 ( .A1(n87), .A2(n88), .ZN(n51) );
  AND2_X1 U77bar ( .A1(n87bar), .A2(n88bar), .ZN(n51bar);
  OR2_X1 U78 ( .A1(n89), .A2(n90), .ZN(n88) );
  AND2_X1 U78bar ( .A1(n89bar), .A2(n90bar), .ZN(n88bar);
  OR2_X1 U79 ( .A1(n91), .A2(n92), .ZN(n90) );
  AND2_X1 U79bar ( .A1(n91bar), .A2(n92bar), .ZN(n90bar);
  OR2_X1 U80 ( .A1(in[118]), .A2(in[109]), .ZN(n92) );
  AND2_X1 U80bar ( .A1(inbar[118]), .A2(inbar[109]), .ZN(n92bar);
  OR2_X1 U81 ( .A1(in[139]), .A2(in[120]), .ZN(n91) );
  AND2_X1 U81bar ( .A1(inbar[139]), .A2(inbar[120]), .ZN(n91bar);
  OR2_X1 U82 ( .A1(n93), .A2(n94), .ZN(n89) );
  AND2_X1 U82bar ( .A1(n93bar), .A2(n94bar), .ZN(n89bar);
  OR2_X1 U83 ( .A1(in[198]), .A2(in[154]), .ZN(n94) );
  AND2_X1 U83bar ( .A1(inbar[198]), .A2(inbar[154]), .ZN(n94bar);
  OR2_X1 U84 ( .A1(in[210]), .A2(in[205]), .ZN(n93) );
  AND2_X1 U84bar ( .A1(inbar[210]), .A2(inbar[205]), .ZN(n93bar);
  OR2_X1 U85 ( .A1(n95), .A2(n96), .ZN(n87) );
  AND2_X1 U85bar ( .A1(n95bar), .A2(n96bar), .ZN(n87bar);
  OR2_X1 U86 ( .A1(n97), .A2(n98), .ZN(n96) );
  AND2_X1 U86bar ( .A1(n97bar), .A2(n98bar), .ZN(n96bar);
  OR2_X1 U87 ( .A1(in[219]), .A2(in[217]), .ZN(n98) );
  AND2_X1 U87bar ( .A1(inbar[219]), .A2(inbar[217]), .ZN(n98bar);
  OR2_X1 U88 ( .A1(in[86]), .A2(in[252]), .ZN(n97) );
  AND2_X1 U88bar ( .A1(inbar[86]), .A2(inbar[252]), .ZN(n97bar);
  OR2_X1 U89 ( .A1(n99), .A2(n100), .ZN(n95) );
  AND2_X1 U89bar ( .A1(n99bar), .A2(n100bar), .ZN(n95bar);
  OR2_X1 U90 ( .A1(in_40), .A2(in[91]), .ZN(n100) );
  AND2_X1 U90bar ( .A1(in_40bar), .A2(inbar[91]), .ZN(n100bar);
  OR2_X1 U91 ( .A1(in_8), .A2(in_46), .ZN(n99) );
  AND2_X1 U91bar ( .A1(in_8bar), .A2(in_46bar), .ZN(n99bar);
  OR2_X1 U92 ( .A1(n101), .A2(n102), .ZN(n84) );
  AND2_X1 U92bar ( .A1(n101bar), .A2(n102bar), .ZN(n84bar);
  OR2_X1 U93 ( .A1(in[117]), .A2(n30), .ZN(n102) );
  AND2_X1 U93bar ( .A1(inbar[117]), .A2(n30bar), .ZN(n102bar);
  OR2_X1 U94 ( .A1(n103), .A2(n104), .ZN(n30) );
  AND2_X1 U94bar ( .A1(n103bar), .A2(n104bar), .ZN(n30bar);
  OR2_X1 U95 ( .A1(n105), .A2(n106), .ZN(n104) );
  AND2_X1 U95bar ( .A1(n105bar), .A2(n106bar), .ZN(n104bar);
  OR2_X1 U96 ( .A1(n107), .A2(n108), .ZN(n106) );
  AND2_X1 U96bar ( .A1(n107bar), .A2(n108bar), .ZN(n106bar);
  OR2_X1 U97 ( .A1(n109), .A2(n110), .ZN(n108) );
  AND2_X1 U97bar ( .A1(n109bar), .A2(n110bar), .ZN(n108bar);
  OR2_X1 U98 ( .A1(in[108]), .A2(n54), .ZN(n107) );
  AND2_X1 U98bar ( .A1(inbar[108]), .A2(n54bar), .ZN(n107bar);
  OR2_X1 U99 ( .A1(n111), .A2(n112), .ZN(n54) );
  AND2_X1 U99bar ( .A1(n111bar), .A2(n112bar), .ZN(n54bar);
  OR2_X1 U100 ( .A1(n113), .A2(n114), .ZN(n112) );
  AND2_X1 U100bar ( .A1(n113bar), .A2(n114bar), .ZN(n112bar);
  OR2_X1 U101 ( .A1(n115), .A2(n116), .ZN(n114) );
  AND2_X1 U101bar ( .A1(n115bar), .A2(n116bar), .ZN(n114bar);
  OR2_X1 U102 ( .A1(in[119]), .A2(in[105]), .ZN(n116) );
  AND2_X1 U102bar ( .A1(inbar[119]), .A2(inbar[105]), .ZN(n116bar);
  OR2_X1 U103 ( .A1(in[186]), .A2(in[175]), .ZN(n115) );
  AND2_X1 U103bar ( .A1(inbar[186]), .A2(inbar[175]), .ZN(n115bar);
  OR2_X1 U104 ( .A1(n117), .A2(n118), .ZN(n113) );
  AND2_X1 U104bar ( .A1(n117bar), .A2(n118bar), .ZN(n113bar);
  OR2_X1 U105 ( .A1(in[202]), .A2(in[193]), .ZN(n118) );
  AND2_X1 U105bar ( .A1(inbar[202]), .A2(inbar[193]), .ZN(n118bar);
  OR2_X1 U106 ( .A1(in[225]), .A2(in[208]), .ZN(n117) );
  AND2_X1 U106bar ( .A1(inbar[225]), .A2(inbar[208]), .ZN(n117bar);
  OR2_X1 U107 ( .A1(n119), .A2(n120), .ZN(n111) );
  AND2_X1 U107bar ( .A1(n119bar), .A2(n120bar), .ZN(n111bar);
  OR2_X1 U108 ( .A1(n121), .A2(n122), .ZN(n120) );
  AND2_X1 U108bar ( .A1(n121bar), .A2(n122bar), .ZN(n120bar);
  OR2_X1 U109 ( .A1(in_1), .A2(in[85]), .ZN(n122) );
  AND2_X1 U109bar ( .A1(in_1bar), .A2(inbar[85]), .ZN(n122bar);
  OR2_X1 U110 ( .A1(in_23), .A2(in_19), .ZN(n121) );
  AND2_X1 U110bar ( .A1(in_23bar), .A2(in_19bar), .ZN(n121bar);
  OR2_X1 U111 ( .A1(n123), .A2(n124), .ZN(n119) );
  AND2_X1 U111bar ( .A1(n123bar), .A2(n124bar), .ZN(n119bar);
  OR2_X1 U112 ( .A1(in_43), .A2(in_33), .ZN(n124) );
  AND2_X1 U112bar ( .A1(in_43bar), .A2(in_33bar), .ZN(n124bar);
  OR2_X1 U113 ( .A1(in_63), .A2(in_44), .ZN(n123) );
  AND2_X1 U113bar ( .A1(in_63bar), .A2(in_44bar), .ZN(n123bar);
  OR2_X1 U114 ( .A1(n125), .A2(n126), .ZN(n105) );
  AND2_X1 U114bar ( .A1(n125bar), .A2(n126bar), .ZN(n105bar);
  OR2_X1 U115 ( .A1(in[141]), .A2(in[112]), .ZN(n126) );
  AND2_X1 U115bar ( .A1(inbar[141]), .A2(inbar[112]), .ZN(n126bar);
  OR2_X1 U116 ( .A1(in[147]), .A2(n127), .ZN(n125) );
  AND2_X1 U116bar ( .A1(inbar[147]), .A2(n127bar), .ZN(n125bar);
  OR2_X1 U117 ( .A1(in[181]), .A2(in[167]), .ZN(n127) );
  AND2_X1 U117bar ( .A1(inbar[181]), .A2(inbar[167]), .ZN(n127bar);
  OR2_X1 U118 ( .A1(n128), .A2(n129), .ZN(n103) );
  AND2_X1 U118bar ( .A1(n128bar), .A2(n129bar), .ZN(n103bar);
  OR2_X1 U119 ( .A1(n130), .A2(n131), .ZN(n129) );
  AND2_X1 U119bar ( .A1(n130bar), .A2(n131bar), .ZN(n129bar);
  OR2_X1 U120 ( .A1(in[229]), .A2(in[201]), .ZN(n131) );
  AND2_X1 U120bar ( .A1(inbar[229]), .A2(inbar[201]), .ZN(n131bar);
  OR2_X1 U121 ( .A1(in[237]), .A2(n132), .ZN(n130) );
  AND2_X1 U121bar ( .A1(inbar[237]), .A2(n132bar), .ZN(n130bar);
  OR2_X1 U122 ( .A1(in[94]), .A2(in[253]), .ZN(n132) );
  AND2_X1 U122bar ( .A1(inbar[94]), .A2(inbar[253]), .ZN(n132bar);
  OR2_X1 U123 ( .A1(n133), .A2(n134), .ZN(n128) );
  AND2_X1 U123bar ( .A1(n133bar), .A2(n134bar), .ZN(n128bar);
  OR2_X1 U124 ( .A1(in_21), .A2(in[96]), .ZN(n134) );
  AND2_X1 U124bar ( .A1(in_21bar), .A2(inbar[96]), .ZN(n134bar);
  OR2_X1 U125 ( .A1(in_25), .A2(n135), .ZN(n133) );
  AND2_X1 U125bar ( .A1(in_25bar), .A2(n135bar), .ZN(n133bar);
  OR2_X1 U126 ( .A1(in_81), .A2(in_45), .ZN(n135) );
  AND2_X1 U126bar ( .A1(in_81bar), .A2(in_45bar), .ZN(n135bar);
  OR2_X1 U127 ( .A1(n136), .A2(n137), .ZN(n82) );
  AND2_X1 U127bar ( .A1(n136bar), .A2(n137bar), .ZN(n82bar);
  OR2_X1 U128 ( .A1(in[142]), .A2(in[124]), .ZN(n137) );
  AND2_X1 U128bar ( .A1(inbar[142]), .A2(inbar[124]), .ZN(n137bar);
  OR2_X1 U129 ( .A1(in[150]), .A2(n138), .ZN(n136) );
  AND2_X1 U129bar ( .A1(inbar[150]), .A2(n138bar), .ZN(n136bar);
  OR2_X1 U130 ( .A1(in[172]), .A2(in[155]), .ZN(n138) );
  AND2_X1 U130bar ( .A1(inbar[172]), .A2(inbar[155]), .ZN(n138bar);
  OR2_X1 U131 ( .A1(n139), .A2(n140), .ZN(n80) );
  AND2_X1 U131bar ( .A1(n139bar), .A2(n140bar), .ZN(n80bar);
  OR2_X1 U132 ( .A1(n141), .A2(n142), .ZN(n140) );
  AND2_X1 U132bar ( .A1(n141bar), .A2(n142bar), .ZN(n140bar);
  OR2_X1 U133 ( .A1(in[196]), .A2(in[173]), .ZN(n142) );
  AND2_X1 U133bar ( .A1(inbar[196]), .A2(inbar[173]), .ZN(n142bar);
  OR2_X1 U134 ( .A1(in[222]), .A2(n143), .ZN(n141) );
  AND2_X1 U134bar ( .A1(inbar[222]), .A2(n143bar), .ZN(n141bar);
  OR2_X1 U135 ( .A1(in[227]), .A2(in[226]), .ZN(n143) );
  AND2_X1 U135bar ( .A1(inbar[227]), .A2(inbar[226]), .ZN(n143bar);
  OR2_X1 U136 ( .A1(n144), .A2(n145), .ZN(n139) );
  AND2_X1 U136bar ( .A1(n144bar), .A2(n145bar), .ZN(n139bar);
  OR2_X1 U137 ( .A1(in[249]), .A2(in[231]), .ZN(n145) );
  AND2_X1 U137bar ( .A1(inbar[249]), .A2(inbar[231]), .ZN(n145bar);
  OR2_X1 U138 ( .A1(in_28), .A2(n146), .ZN(n144) );
  AND2_X1 U138bar ( .A1(in_28bar), .A2(n146bar), .ZN(n144bar);
  OR2_X1 U139 ( .A1(in_52), .A2(in_47), .ZN(n146) );
  AND2_X1 U139bar ( .A1(in_52bar), .A2(in_47bar), .ZN(n146bar);
  OR2_X1 U140 ( .A1(n147), .A2(n148), .ZN(out[3]) );
  AND2_X1 U140bar ( .A1(n147bar), .A2(n148bar), .ZN(outbar[3]);
  OR2_X1 U141 ( .A1(n149), .A2(n150), .ZN(n148) );
  AND2_X1 U141bar ( .A1(n149bar), .A2(n150bar), .ZN(n148bar);
  OR2_X1 U142 ( .A1(n151), .A2(n152), .ZN(n150) );
  AND2_X1 U142bar ( .A1(n151bar), .A2(n152bar), .ZN(n150bar);
  OR2_X1 U143 ( .A1(n153), .A2(n154), .ZN(n152) );
  AND2_X1 U143bar ( .A1(n153bar), .A2(n154bar), .ZN(n152bar);
  OR2_X1 U144 ( .A1(n9), .A2(n155), .ZN(n151) );
  AND2_X1 U144bar ( .A1(n9bar), .A2(n155bar), .ZN(n151bar);
  OR2_X1 U145 ( .A1(in[118]), .A2(n156), .ZN(n155) );
  AND2_X1 U145bar ( .A1(inbar[118]), .A2(n156bar), .ZN(n155bar);
  OR2_X1 U146 ( .A1(n157), .A2(n158), .ZN(n9) );
  AND2_X1 U146bar ( .A1(n157bar), .A2(n158bar), .ZN(n9bar);
  OR2_X1 U147 ( .A1(n159), .A2(n160), .ZN(n158) );
  AND2_X1 U147bar ( .A1(n159bar), .A2(n160bar), .ZN(n158bar);
  OR2_X1 U148 ( .A1(n161), .A2(n162), .ZN(n160) );
  AND2_X1 U148bar ( .A1(n161bar), .A2(n162bar), .ZN(n160bar);
  OR2_X1 U149 ( .A1(in[122]), .A2(in[111]), .ZN(n162) );
  AND2_X1 U149bar ( .A1(inbar[122]), .A2(inbar[111]), .ZN(n162bar);
  OR2_X1 U150 ( .A1(in[154]), .A2(in[151]), .ZN(n161) );
  AND2_X1 U150bar ( .A1(inbar[154]), .A2(inbar[151]), .ZN(n161bar);
  OR2_X1 U151 ( .A1(n163), .A2(n164), .ZN(n159) );
  AND2_X1 U151bar ( .A1(n163bar), .A2(n164bar), .ZN(n159bar);
  OR2_X1 U152 ( .A1(in[187]), .A2(in[177]), .ZN(n164) );
  AND2_X1 U152bar ( .A1(inbar[187]), .A2(inbar[177]), .ZN(n164bar);
  OR2_X1 U153 ( .A1(in[200]), .A2(in[192]), .ZN(n163) );
  AND2_X1 U153bar ( .A1(inbar[200]), .A2(inbar[192]), .ZN(n163bar);
  OR2_X1 U154 ( .A1(n165), .A2(n166), .ZN(n157) );
  AND2_X1 U154bar ( .A1(n165bar), .A2(n166bar), .ZN(n157bar);
  OR2_X1 U155 ( .A1(n167), .A2(n168), .ZN(n166) );
  AND2_X1 U155bar ( .A1(n167bar), .A2(n168bar), .ZN(n166bar);
  OR2_X1 U156 ( .A1(in[225]), .A2(in[207]), .ZN(n168) );
  AND2_X1 U156bar ( .A1(inbar[225]), .A2(inbar[207]), .ZN(n168bar);
  OR2_X1 U157 ( .A1(in[98]), .A2(in[226]), .ZN(n167) );
  AND2_X1 U157bar ( .A1(inbar[98]), .A2(inbar[226]), .ZN(n167bar);
  OR2_X1 U158 ( .A1(n169), .A2(n170), .ZN(n165) );
  AND2_X1 U158bar ( .A1(n169bar), .A2(n170bar), .ZN(n165bar);
  OR2_X1 U159 ( .A1(in_20), .A2(in_16), .ZN(n170) );
  AND2_X1 U159bar ( .A1(in_20bar), .A2(in_16bar), .ZN(n170bar);
  OR2_X1 U160 ( .A1(in_55), .A2(in_45), .ZN(n169) );
  AND2_X1 U160bar ( .A1(in_55bar), .A2(in_45bar), .ZN(n169bar);
  OR2_X1 U161 ( .A1(n171), .A2(n172), .ZN(n149) );
  AND2_X1 U161bar ( .A1(n171bar), .A2(n172bar), .ZN(n149bar);
  OR2_X1 U162 ( .A1(in[162]), .A2(in[149]), .ZN(n172) );
  AND2_X1 U162bar ( .A1(inbar[162]), .A2(inbar[149]), .ZN(n172bar);
  OR2_X1 U163 ( .A1(in[163]), .A2(n173), .ZN(n171) );
  AND2_X1 U163bar ( .A1(inbar[163]), .A2(n173bar), .ZN(n171bar);
  OR2_X1 U164 ( .A1(in[191]), .A2(in[189]), .ZN(n173) );
  AND2_X1 U164bar ( .A1(inbar[191]), .A2(inbar[189]), .ZN(n173bar);
  OR2_X1 U165 ( .A1(n174), .A2(n175), .ZN(n147) );
  AND2_X1 U165bar ( .A1(n174bar), .A2(n175bar), .ZN(n147bar);
  OR2_X1 U166 ( .A1(n176), .A2(n177), .ZN(n175) );
  AND2_X1 U166bar ( .A1(n176bar), .A2(n177bar), .ZN(n175bar);
  OR2_X1 U167 ( .A1(in[212]), .A2(in[193]), .ZN(n177) );
  AND2_X1 U167bar ( .A1(inbar[212]), .A2(inbar[193]), .ZN(n177bar);
  OR2_X1 U168 ( .A1(in[238]), .A2(n178), .ZN(n176) );
  AND2_X1 U168bar ( .A1(inbar[238]), .A2(n178bar), .ZN(n176bar);
  OR2_X1 U169 ( .A1(in[88]), .A2(in[247]), .ZN(n178) );
  AND2_X1 U169bar ( .A1(inbar[88]), .A2(inbar[247]), .ZN(n178bar);
  OR2_X1 U170 ( .A1(n179), .A2(n180), .ZN(n174) );
  AND2_X1 U170bar ( .A1(n179bar), .A2(n180bar), .ZN(n174bar);
  OR2_X1 U171 ( .A1(in[94]), .A2(in[92]), .ZN(n180) );
  AND2_X1 U171bar ( .A1(inbar[94]), .A2(inbar[92]), .ZN(n180bar);
  OR2_X1 U172 ( .A1(in_52), .A2(n181), .ZN(n179) );
  AND2_X1 U172bar ( .A1(in_52bar), .A2(n181bar), .ZN(n179bar);
  OR2_X1 U173 ( .A1(in_70), .A2(in_67), .ZN(n181) );
  AND2_X1 U173bar ( .A1(in_70bar), .A2(in_67bar), .ZN(n181bar);
  OR2_X1 U174 ( .A1(n182), .A2(n183), .ZN(out[2]) );
  AND2_X1 U174bar ( .A1(n182bar), .A2(n183bar), .ZN(outbar[2]);
  OR2_X1 U175 ( .A1(n184), .A2(n185), .ZN(n183) );
  AND2_X1 U175bar ( .A1(n184bar), .A2(n185bar), .ZN(n183bar);
  OR2_X1 U176 ( .A1(n186), .A2(n187), .ZN(n185) );
  AND2_X1 U176bar ( .A1(n186bar), .A2(n187bar), .ZN(n185bar);
  OR2_X1 U177 ( .A1(n154), .A2(n188), .ZN(n187) );
  AND2_X1 U177bar ( .A1(n154bar), .A2(n188bar), .ZN(n187bar);
  OR2_X1 U178 ( .A1(n189), .A2(n190), .ZN(n154) );
  AND2_X1 U178bar ( .A1(n189bar), .A2(n190bar), .ZN(n154bar);
  OR2_X1 U179 ( .A1(n191), .A2(n192), .ZN(n190) );
  AND2_X1 U179bar ( .A1(n191bar), .A2(n192bar), .ZN(n190bar);
  OR2_X1 U180 ( .A1(n193), .A2(n194), .ZN(n192) );
  AND2_X1 U180bar ( .A1(n193bar), .A2(n194bar), .ZN(n192bar);
  OR2_X1 U181 ( .A1(n11), .A2(n195), .ZN(n194) );
  AND2_X1 U181bar ( .A1(n11bar), .A2(n195bar), .ZN(n194bar);
  OR2_X1 U182 ( .A1(n196), .A2(n197), .ZN(n11) );
  AND2_X1 U182bar ( .A1(n196bar), .A2(n197bar), .ZN(n11bar);
  OR2_X1 U183 ( .A1(n198), .A2(n199), .ZN(n197) );
  AND2_X1 U183bar ( .A1(n198bar), .A2(n199bar), .ZN(n197bar);
  OR2_X1 U184 ( .A1(n200), .A2(n201), .ZN(n199) );
  AND2_X1 U184bar ( .A1(n200bar), .A2(n201bar), .ZN(n199bar);
  OR2_X1 U185 ( .A1(in[131]), .A2(in[120]), .ZN(n201) );
  AND2_X1 U185bar ( .A1(inbar[131]), .A2(inbar[120]), .ZN(n201bar);
  OR2_X1 U186 ( .A1(in[153]), .A2(in[147]), .ZN(n200) );
  AND2_X1 U186bar ( .A1(inbar[153]), .A2(inbar[147]), .ZN(n200bar);
  OR2_X1 U187 ( .A1(n202), .A2(n203), .ZN(n198) );
  AND2_X1 U187bar ( .A1(n202bar), .A2(n203bar), .ZN(n198bar);
  OR2_X1 U188 ( .A1(in[170]), .A2(in[156]), .ZN(n203) );
  AND2_X1 U188bar ( .A1(inbar[170]), .A2(inbar[156]), .ZN(n203bar);
  OR2_X1 U189 ( .A1(in[223]), .A2(in[190]), .ZN(n202) );
  AND2_X1 U189bar ( .A1(inbar[223]), .A2(inbar[190]), .ZN(n202bar);
  OR2_X1 U190 ( .A1(n204), .A2(n205), .ZN(n196) );
  AND2_X1 U190bar ( .A1(n204bar), .A2(n205bar), .ZN(n196bar);
  OR2_X1 U191 ( .A1(n206), .A2(n207), .ZN(n205) );
  AND2_X1 U191bar ( .A1(n206bar), .A2(n207bar), .ZN(n205bar);
  OR2_X1 U192 ( .A1(in[236]), .A2(in[230]), .ZN(n207) );
  AND2_X1 U192bar ( .A1(inbar[236]), .A2(inbar[230]), .ZN(n207bar);
  OR2_X1 U193 ( .A1(in[85]), .A2(in[240]), .ZN(n206) );
  AND2_X1 U193bar ( .A1(inbar[85]), .A2(inbar[240]), .ZN(n206bar);
  OR2_X1 U194 ( .A1(n208), .A2(n209), .ZN(n204) );
  AND2_X1 U194bar ( .A1(n208bar), .A2(n209bar), .ZN(n204bar);
  OR2_X1 U195 ( .A1(in_12), .A2(in[90]), .ZN(n209) );
  AND2_X1 U195bar ( .A1(in_12bar), .A2(inbar[90]), .ZN(n209bar);
  OR2_X1 U196 ( .A1(in_39), .A2(in_28), .ZN(n208) );
  AND2_X1 U196bar ( .A1(in_39bar), .A2(in_28bar), .ZN(n208bar);
  OR2_X1 U197 ( .A1(in[109]), .A2(n210), .ZN(n193) );
  AND2_X1 U197bar ( .A1(inbar[109]), .A2(n210bar), .ZN(n193bar);
  OR2_X1 U198 ( .A1(n211), .A2(n212), .ZN(n191) );
  AND2_X1 U198bar ( .A1(n211bar), .A2(n212bar), .ZN(n191bar);
  OR2_X1 U199 ( .A1(in[138]), .A2(in[129]), .ZN(n212) );
  AND2_X1 U199bar ( .A1(inbar[138]), .A2(inbar[129]), .ZN(n212bar);
  OR2_X1 U200 ( .A1(in[157]), .A2(n213), .ZN(n211) );
  AND2_X1 U200bar ( .A1(inbar[157]), .A2(n213bar), .ZN(n211bar);
  OR2_X1 U201 ( .A1(in[182]), .A2(in[167]), .ZN(n213) );
  AND2_X1 U201bar ( .A1(inbar[182]), .A2(inbar[167]), .ZN(n213bar);
  OR2_X1 U202 ( .A1(n214), .A2(n215), .ZN(n189) );
  AND2_X1 U202bar ( .A1(n214bar), .A2(n215bar), .ZN(n189bar);
  OR2_X1 U203 ( .A1(n216), .A2(n217), .ZN(n215) );
  AND2_X1 U203bar ( .A1(n216bar), .A2(n217bar), .ZN(n215bar);
  OR2_X1 U204 ( .A1(in[195]), .A2(in[184]), .ZN(n217) );
  AND2_X1 U204bar ( .A1(inbar[195]), .A2(inbar[184]), .ZN(n217bar);
  OR2_X1 U205 ( .A1(in[196]), .A2(n218), .ZN(n216) );
  AND2_X1 U205bar ( .A1(inbar[196]), .A2(n218bar), .ZN(n216bar);
  OR2_X1 U206 ( .A1(in[215]), .A2(in[209]), .ZN(n218) );
  AND2_X1 U206bar ( .A1(inbar[215]), .A2(inbar[209]), .ZN(n218bar);
  OR2_X1 U207 ( .A1(n219), .A2(n220), .ZN(n214) );
  AND2_X1 U207bar ( .A1(n219bar), .A2(n220bar), .ZN(n214bar);
  OR2_X1 U208 ( .A1(in[93]), .A2(in[233]), .ZN(n220) );
  AND2_X1 U208bar ( .A1(inbar[93]), .A2(inbar[233]), .ZN(n220bar);
  OR2_X1 U209 ( .A1(in_1), .A2(n221), .ZN(n219) );
  AND2_X1 U209bar ( .A1(in_1bar), .A2(n221bar), .ZN(n219bar);
  OR2_X1 U210 ( .A1(in_69), .A2(in_66), .ZN(n221) );
  AND2_X1 U210bar ( .A1(in_69bar), .A2(in_66bar), .ZN(n221bar);
  OR2_X1 U211 ( .A1(n7), .A2(n222), .ZN(n186) );
  AND2_X1 U211bar ( .A1(n7bar), .A2(n222bar), .ZN(n186bar);
  OR2_X1 U212 ( .A1(in[134]), .A2(n223), .ZN(n222) );
  AND2_X1 U212bar ( .A1(inbar[134]), .A2(n223bar), .ZN(n222bar);
  OR2_X1 U213 ( .A1(n224), .A2(n225), .ZN(n7) );
  AND2_X1 U213bar ( .A1(n224bar), .A2(n225bar), .ZN(n7bar);
  OR2_X1 U214 ( .A1(n226), .A2(n227), .ZN(n225) );
  AND2_X1 U214bar ( .A1(n226bar), .A2(n227bar), .ZN(n225bar);
  OR2_X1 U215 ( .A1(n228), .A2(n229), .ZN(n227) );
  AND2_X1 U215bar ( .A1(n228bar), .A2(n229bar), .ZN(n227bar);
  OR2_X1 U216 ( .A1(in[136]), .A2(in[121]), .ZN(n229) );
  AND2_X1 U216bar ( .A1(inbar[136]), .A2(inbar[121]), .ZN(n229bar);
  OR2_X1 U217 ( .A1(in[186]), .A2(in[174]), .ZN(n228) );
  AND2_X1 U217bar ( .A1(inbar[186]), .A2(inbar[174]), .ZN(n228bar);
  OR2_X1 U218 ( .A1(n230), .A2(n231), .ZN(n226) );
  AND2_X1 U218bar ( .A1(n230bar), .A2(n231bar), .ZN(n226bar);
  OR2_X1 U219 ( .A1(in[198]), .A2(in[197]), .ZN(n231) );
  AND2_X1 U219bar ( .A1(inbar[198]), .A2(inbar[197]), .ZN(n231bar);
  OR2_X1 U220 ( .A1(in[214]), .A2(in[199]), .ZN(n230) );
  AND2_X1 U220bar ( .A1(inbar[214]), .A2(inbar[199]), .ZN(n230bar);
  OR2_X1 U221 ( .A1(n232), .A2(n233), .ZN(n224) );
  AND2_X1 U221bar ( .A1(n232bar), .A2(n233bar), .ZN(n224bar);
  OR2_X1 U222 ( .A1(n234), .A2(n235), .ZN(n233) );
  AND2_X1 U222bar ( .A1(n234bar), .A2(n235bar), .ZN(n233bar);
  OR2_X1 U223 ( .A1(in[231]), .A2(in[220]), .ZN(n235) );
  AND2_X1 U223bar ( .A1(inbar[231]), .A2(inbar[220]), .ZN(n235bar);
  OR2_X1 U224 ( .A1(in_25), .A2(in[245]), .ZN(n234) );
  AND2_X1 U224bar ( .A1(in_25bar), .A2(inbar[245]), .ZN(n234bar);
  OR2_X1 U225 ( .A1(n236), .A2(n237), .ZN(n232) );
  AND2_X1 U225bar ( .A1(n236bar), .A2(n237bar), .ZN(n232bar);
  OR2_X1 U226 ( .A1(in_53), .A2(in_29), .ZN(n237) );
  AND2_X1 U226bar ( .A1(in_53bar), .A2(in_29bar), .ZN(n237bar);
  OR2_X1 U227 ( .A1(in_79), .A2(in_74), .ZN(n236) );
  AND2_X1 U227bar ( .A1(in_79bar), .A2(in_74bar), .ZN(n236bar);
  OR2_X1 U228 ( .A1(n238), .A2(n239), .ZN(n184) );
  AND2_X1 U228bar ( .A1(n238bar), .A2(n239bar), .ZN(n184bar);
  OR2_X1 U229 ( .A1(in[152]), .A2(in[140]), .ZN(n239) );
  AND2_X1 U229bar ( .A1(inbar[152]), .A2(inbar[140]), .ZN(n239bar);
  OR2_X1 U230 ( .A1(in[155]), .A2(n240), .ZN(n238) );
  AND2_X1 U230bar ( .A1(inbar[155]), .A2(n240bar), .ZN(n238bar);
  OR2_X1 U231 ( .A1(in[166]), .A2(in[165]), .ZN(n240) );
  AND2_X1 U231bar ( .A1(inbar[166]), .A2(inbar[165]), .ZN(n240bar);
  OR2_X1 U232 ( .A1(n241), .A2(n242), .ZN(n182) );
  AND2_X1 U232bar ( .A1(n241bar), .A2(n242bar), .ZN(n182bar);
  OR2_X1 U233 ( .A1(n243), .A2(n244), .ZN(n242) );
  AND2_X1 U233bar ( .A1(n243bar), .A2(n244bar), .ZN(n242bar);
  OR2_X1 U234 ( .A1(in[202]), .A2(in[185]), .ZN(n244) );
  AND2_X1 U234bar ( .A1(inbar[202]), .A2(inbar[185]), .ZN(n244bar);
  OR2_X1 U235 ( .A1(in[211]), .A2(n245), .ZN(n243) );
  AND2_X1 U235bar ( .A1(inbar[211]), .A2(n245bar), .ZN(n243bar);
  OR2_X1 U236 ( .A1(in[255]), .A2(in[253]), .ZN(n245) );
  AND2_X1 U236bar ( .A1(inbar[255]), .A2(inbar[253]), .ZN(n245bar);
  OR2_X1 U237 ( .A1(n246), .A2(n247), .ZN(n241) );
  AND2_X1 U237bar ( .A1(n246bar), .A2(n247bar), .ZN(n241bar);
  OR2_X1 U238 ( .A1(in_35), .A2(in_15), .ZN(n247) );
  AND2_X1 U238bar ( .A1(in_35bar), .A2(in_15bar), .ZN(n247bar);
  OR2_X1 U239 ( .A1(in_36), .A2(n248), .ZN(n246) );
  AND2_X1 U239bar ( .A1(in_36bar), .A2(n248bar), .ZN(n246bar);
  OR2_X1 U240 ( .A1(in_48), .A2(in_40), .ZN(n248) );
  AND2_X1 U240bar ( .A1(in_48bar), .A2(in_40bar), .ZN(n248bar);
  OR2_X1 U241 ( .A1(n249), .A2(n250), .ZN(out[1]) );
  AND2_X1 U241bar ( .A1(n249bar), .A2(n250bar), .ZN(outbar[1]);
  OR2_X1 U242 ( .A1(n251), .A2(n252), .ZN(n250) );
  AND2_X1 U242bar ( .A1(n251bar), .A2(n252bar), .ZN(n250bar);
  OR2_X1 U243 ( .A1(n253), .A2(n254), .ZN(n252) );
  AND2_X1 U243bar ( .A1(n253bar), .A2(n254bar), .ZN(n252bar);
  OR2_X1 U244 ( .A1(n52), .A2(n86), .ZN(n254) );
  AND2_X1 U244bar ( .A1(n52bar), .A2(n86bar), .ZN(n254bar);
  OR2_X1 U245 ( .A1(n255), .A2(n256), .ZN(n86) );
  AND2_X1 U245bar ( .A1(n255bar), .A2(n256bar), .ZN(n86bar);
  OR2_X1 U246 ( .A1(n257), .A2(n258), .ZN(n256) );
  AND2_X1 U246bar ( .A1(n257bar), .A2(n258bar), .ZN(n256bar);
  OR2_X1 U247 ( .A1(n259), .A2(n260), .ZN(n258) );
  AND2_X1 U247bar ( .A1(n259bar), .A2(n260bar), .ZN(n258bar);
  OR2_X1 U248 ( .A1(in[116]), .A2(in[110]), .ZN(n260) );
  AND2_X1 U248bar ( .A1(inbar[116]), .A2(inbar[110]), .ZN(n260bar);
  OR2_X1 U249 ( .A1(in[133]), .A2(in[130]), .ZN(n259) );
  AND2_X1 U249bar ( .A1(inbar[133]), .A2(inbar[130]), .ZN(n259bar);
  OR2_X1 U250 ( .A1(n261), .A2(n262), .ZN(n257) );
  AND2_X1 U250bar ( .A1(n261bar), .A2(n262bar), .ZN(n257bar);
  OR2_X1 U251 ( .A1(in[203]), .A2(in[135]), .ZN(n262) );
  AND2_X1 U251bar ( .A1(inbar[203]), .A2(inbar[135]), .ZN(n262bar);
  OR2_X1 U252 ( .A1(in[232]), .A2(in[223]), .ZN(n261) );
  AND2_X1 U252bar ( .A1(inbar[232]), .A2(inbar[223]), .ZN(n261bar);
  OR2_X1 U253 ( .A1(n263), .A2(n264), .ZN(n255) );
  AND2_X1 U253bar ( .A1(n263bar), .A2(n264bar), .ZN(n255bar);
  OR2_X1 U254 ( .A1(n265), .A2(n266), .ZN(n264) );
  AND2_X1 U254bar ( .A1(n265bar), .A2(n266bar), .ZN(n264bar);
  OR2_X1 U255 ( .A1(in[255]), .A2(in[233]), .ZN(n266) );
  AND2_X1 U255bar ( .A1(inbar[255]), .A2(inbar[233]), .ZN(n266bar);
  OR2_X1 U256 ( .A1(in_53), .A2(in_34), .ZN(n265) );
  AND2_X1 U256bar ( .A1(in_53bar), .A2(in_34bar), .ZN(n265bar);
  OR2_X1 U257 ( .A1(n267), .A2(n268), .ZN(n263) );
  AND2_X1 U257bar ( .A1(n267bar), .A2(n268bar), .ZN(n263bar);
  OR2_X1 U258 ( .A1(in_57), .A2(in_55), .ZN(n268) );
  AND2_X1 U258bar ( .A1(in_57bar), .A2(in_55bar), .ZN(n268bar);
  OR2_X1 U259 ( .A1(in_68), .A2(in_67), .ZN(n267) );
  AND2_X1 U259bar ( .A1(in_68bar), .A2(in_67bar), .ZN(n267bar);
  OR2_X1 U260 ( .A1(n269), .A2(n270), .ZN(n52) );
  AND2_X1 U260bar ( .A1(n269bar), .A2(n270bar), .ZN(n52bar);
  OR2_X1 U261 ( .A1(n271), .A2(n272), .ZN(n270) );
  AND2_X1 U261bar ( .A1(n271bar), .A2(n272bar), .ZN(n270bar);
  OR2_X1 U262 ( .A1(n273), .A2(n274), .ZN(n272) );
  AND2_X1 U262bar ( .A1(n273bar), .A2(n274bar), .ZN(n272bar);
  OR2_X1 U263 ( .A1(n29), .A2(n101), .ZN(n274) );
  AND2_X1 U263bar ( .A1(n29bar), .A2(n101bar), .ZN(n274bar);
  OR2_X1 U264 ( .A1(n275), .A2(n276), .ZN(n101) );
  AND2_X1 U264bar ( .A1(n275bar), .A2(n276bar), .ZN(n101bar);
  OR2_X1 U265 ( .A1(n277), .A2(n278), .ZN(n276) );
  AND2_X1 U265bar ( .A1(n277bar), .A2(n278bar), .ZN(n276bar);
  OR2_X1 U266 ( .A1(n279), .A2(n280), .ZN(n278) );
  AND2_X1 U266bar ( .A1(n279bar), .A2(n280bar), .ZN(n278bar);
  OR2_X1 U267 ( .A1(in[121]), .A2(in[102]), .ZN(n280) );
  AND2_X1 U267bar ( .A1(inbar[121]), .A2(inbar[102]), .ZN(n280bar);
  OR2_X1 U268 ( .A1(in[162]), .A2(in[161]), .ZN(n279) );
  AND2_X1 U268bar ( .A1(inbar[162]), .A2(inbar[161]), .ZN(n279bar);
  OR2_X1 U269 ( .A1(n281), .A2(n282), .ZN(n277) );
  AND2_X1 U269bar ( .A1(n281bar), .A2(n282bar), .ZN(n277bar);
  OR2_X1 U270 ( .A1(in[192]), .A2(in[178]), .ZN(n282) );
  AND2_X1 U270bar ( .A1(inbar[192]), .A2(inbar[178]), .ZN(n282bar);
  OR2_X1 U271 ( .A1(in[244]), .A2(in[209]), .ZN(n281) );
  AND2_X1 U271bar ( .A1(inbar[244]), .A2(inbar[209]), .ZN(n281bar);
  OR2_X1 U272 ( .A1(n283), .A2(n284), .ZN(n275) );
  AND2_X1 U272bar ( .A1(n283bar), .A2(n284bar), .ZN(n275bar);
  OR2_X1 U273 ( .A1(n285), .A2(n286), .ZN(n284) );
  AND2_X1 U273bar ( .A1(n285bar), .A2(n286bar), .ZN(n284bar);
  OR2_X1 U274 ( .A1(in[90]), .A2(in[254]), .ZN(n286) );
  AND2_X1 U274bar ( .A1(inbar[90]), .A2(inbar[254]), .ZN(n286bar);
  OR2_X1 U275 ( .A1(in_36), .A2(in_32), .ZN(n285) );
  AND2_X1 U275bar ( .A1(in_36bar), .A2(in_32bar), .ZN(n285bar);
  OR2_X1 U276 ( .A1(n287), .A2(n288), .ZN(n283) );
  AND2_X1 U276bar ( .A1(n287bar), .A2(n288bar), .ZN(n283bar);
  OR2_X1 U277 ( .A1(in_62), .A2(in_37), .ZN(n288) );
  AND2_X1 U277bar ( .A1(in_62bar), .A2(in_37bar), .ZN(n288bar);
  OR2_X1 U278 ( .A1(in_75), .A2(in_73), .ZN(n287) );
  AND2_X1 U278bar ( .A1(in_75bar), .A2(in_73bar), .ZN(n287bar);
  OR2_X1 U279 ( .A1(n289), .A2(n290), .ZN(n29) );
  AND2_X1 U279bar ( .A1(n289bar), .A2(n290bar), .ZN(n29bar);
  OR2_X1 U280 ( .A1(n291), .A2(n292), .ZN(n290) );
  AND2_X1 U280bar ( .A1(n291bar), .A2(n292bar), .ZN(n290bar);
  OR2_X1 U281 ( .A1(n293), .A2(n294), .ZN(n292) );
  AND2_X1 U281bar ( .A1(n293bar), .A2(n294bar), .ZN(n292bar);
  OR2_X1 U282 ( .A1(in[171]), .A2(in[153]), .ZN(n294) );
  AND2_X1 U282bar ( .A1(inbar[171]), .A2(inbar[153]), .ZN(n294bar);
  OR2_X1 U283 ( .A1(in[187]), .A2(in[176]), .ZN(n293) );
  AND2_X1 U283bar ( .A1(inbar[187]), .A2(inbar[176]), .ZN(n293bar);
  OR2_X1 U284 ( .A1(n295), .A2(n296), .ZN(n291) );
  AND2_X1 U284bar ( .A1(n295bar), .A2(n296bar), .ZN(n291bar);
  OR2_X1 U285 ( .A1(in[245]), .A2(in[211]), .ZN(n296) );
  AND2_X1 U285bar ( .A1(inbar[245]), .A2(inbar[211]), .ZN(n296bar);
  OR2_X1 U286 ( .A1(in[97]), .A2(in[88]), .ZN(n295) );
  AND2_X1 U286bar ( .A1(inbar[97]), .A2(inbar[88]), .ZN(n295bar);
  OR2_X1 U287 ( .A1(n297), .A2(n298), .ZN(n289) );
  AND2_X1 U287bar ( .A1(n297bar), .A2(n298bar), .ZN(n289bar);
  OR2_X1 U288 ( .A1(n299), .A2(n300), .ZN(n298) );
  AND2_X1 U288bar ( .A1(n299bar), .A2(n300bar), .ZN(n298bar);
  OR2_X1 U289 ( .A1(in_10), .A2(in_0), .ZN(n300) );
  AND2_X1 U289bar ( .A1(in_10bar), .A2(in_0bar), .ZN(n300bar);
  OR2_X1 U290 ( .A1(in_59), .A2(in_5), .ZN(n299) );
  AND2_X1 U290bar ( .A1(in_59bar), .A2(in_5bar), .ZN(n299bar);
  OR2_X1 U291 ( .A1(n301), .A2(n302), .ZN(n297) );
  AND2_X1 U291bar ( .A1(n301bar), .A2(n302bar), .ZN(n297bar);
  OR2_X1 U292 ( .A1(in_60), .A2(in_6), .ZN(n302) );
  AND2_X1 U292bar ( .A1(in_60bar), .A2(in_6bar), .ZN(n302bar);
  OR2_X1 U293 ( .A1(in_77), .A2(in_69), .ZN(n301) );
  AND2_X1 U293bar ( .A1(in_77bar), .A2(in_69bar), .ZN(n301bar);
  OR2_X1 U294 ( .A1(in[113]), .A2(n109), .ZN(n273) );
  AND2_X1 U294bar ( .A1(inbar[113]), .A2(n109bar), .ZN(n273bar);
  OR2_X1 U295 ( .A1(n303), .A2(n304), .ZN(n109) );
  AND2_X1 U295bar ( .A1(n303bar), .A2(n304bar), .ZN(n109bar);
  OR2_X1 U296 ( .A1(n305), .A2(n306), .ZN(n304) );
  AND2_X1 U296bar ( .A1(n305bar), .A2(n306bar), .ZN(n304bar);
  OR2_X1 U297 ( .A1(n307), .A2(n308), .ZN(n306) );
  AND2_X1 U297bar ( .A1(n307bar), .A2(n308bar), .ZN(n306bar);
  OR2_X1 U298 ( .A1(in[125]), .A2(in[107]), .ZN(n308) );
  AND2_X1 U298bar ( .A1(inbar[125]), .A2(inbar[107]), .ZN(n308bar);
  OR2_X1 U299 ( .A1(in[138]), .A2(in[126]), .ZN(n307) );
  AND2_X1 U299bar ( .A1(inbar[138]), .A2(inbar[126]), .ZN(n307bar);
  OR2_X1 U300 ( .A1(n309), .A2(n310), .ZN(n305) );
  AND2_X1 U300bar ( .A1(n309bar), .A2(n310bar), .ZN(n305bar);
  OR2_X1 U301 ( .A1(in[189]), .A2(in[143]), .ZN(n310) );
  AND2_X1 U301bar ( .A1(inbar[189]), .A2(inbar[143]), .ZN(n310bar);
  OR2_X1 U302 ( .A1(in[99]), .A2(in[214]), .ZN(n309) );
  AND2_X1 U302bar ( .A1(inbar[99]), .A2(inbar[214]), .ZN(n309bar);
  OR2_X1 U303 ( .A1(n311), .A2(n312), .ZN(n303) );
  AND2_X1 U303bar ( .A1(n311bar), .A2(n312bar), .ZN(n303bar);
  OR2_X1 U304 ( .A1(n313), .A2(n314), .ZN(n312) );
  AND2_X1 U304bar ( .A1(n313bar), .A2(n314bar), .ZN(n312bar);
  OR2_X1 U305 ( .A1(in_15), .A2(in_12), .ZN(n314) );
  AND2_X1 U305bar ( .A1(in_15bar), .A2(in_12bar), .ZN(n314bar);
  OR2_X1 U306 ( .A1(in_20), .A2(in_2), .ZN(n313) );
  AND2_X1 U306bar ( .A1(in_20bar), .A2(in_2bar), .ZN(n313bar);
  OR2_X1 U307 ( .A1(n315), .A2(n316), .ZN(n311) );
  AND2_X1 U307bar ( .A1(n315bar), .A2(n316bar), .ZN(n311bar);
  OR2_X1 U308 ( .A1(in_30), .A2(in_3), .ZN(n316) );
  AND2_X1 U308bar ( .A1(in_30bar), .A2(in_3bar), .ZN(n316bar);
  OR2_X1 U309 ( .A1(in_4), .A2(in_38), .ZN(n315) );
  AND2_X1 U309bar ( .A1(in_4bar), .A2(in_38bar), .ZN(n315bar);
  OR2_X1 U310 ( .A1(n317), .A2(n318), .ZN(n271) );
  AND2_X1 U310bar ( .A1(n317bar), .A2(n318bar), .ZN(n271bar);
  OR2_X1 U311 ( .A1(in[148]), .A2(in[137]), .ZN(n318) );
  AND2_X1 U311bar ( .A1(inbar[148]), .A2(inbar[137]), .ZN(n318bar);
  OR2_X1 U312 ( .A1(in[149]), .A2(n319), .ZN(n317) );
  AND2_X1 U312bar ( .A1(inbar[149]), .A2(n319bar), .ZN(n317bar);
  OR2_X1 U313 ( .A1(in[195]), .A2(in[190]), .ZN(n319) );
  AND2_X1 U313bar ( .A1(inbar[195]), .A2(inbar[190]), .ZN(n319bar);
  OR2_X1 U314 ( .A1(n320), .A2(n321), .ZN(n269) );
  AND2_X1 U314bar ( .A1(n320bar), .A2(n321bar), .ZN(n269bar);
  OR2_X1 U315 ( .A1(n322), .A2(n323), .ZN(n321) );
  AND2_X1 U315bar ( .A1(n322bar), .A2(n323bar), .ZN(n321bar);
  OR2_X1 U316 ( .A1(in[98]), .A2(in[197]), .ZN(n323) );
  AND2_X1 U316bar ( .A1(inbar[98]), .A2(inbar[197]), .ZN(n323bar);
  OR2_X1 U317 ( .A1(in_11), .A2(n324), .ZN(n322) );
  AND2_X1 U317bar ( .A1(in_11bar), .A2(n324bar), .ZN(n322bar);
  OR2_X1 U318 ( .A1(in_26), .A2(in_14), .ZN(n324) );
  AND2_X1 U318bar ( .A1(in_26bar), .A2(in_14bar), .ZN(n324bar);
  OR2_X1 U319 ( .A1(n325), .A2(n326), .ZN(n320) );
  AND2_X1 U319bar ( .A1(n325bar), .A2(n326bar), .ZN(n320bar);
  OR2_X1 U320 ( .A1(in_35), .A2(in_27), .ZN(n326) );
  AND2_X1 U320bar ( .A1(in_35bar), .A2(in_27bar), .ZN(n326bar);
  OR2_X1 U321 ( .A1(in_50), .A2(n327), .ZN(n325) );
  AND2_X1 U321bar ( .A1(in_50bar), .A2(n327bar), .ZN(n325bar);
  OR2_X1 U322 ( .A1(in_78), .A2(in_61), .ZN(n327) );
  AND2_X1 U322bar ( .A1(in_78bar), .A2(in_61bar), .ZN(n327bar);
  OR2_X1 U323 ( .A1(n31), .A2(n328), .ZN(n253) );
  AND2_X1 U323bar ( .A1(n31bar), .A2(n328bar), .ZN(n253bar);
  OR2_X1 U324 ( .A1(in[106]), .A2(n110), .ZN(n328) );
  AND2_X1 U324bar ( .A1(inbar[106]), .A2(n110bar), .ZN(n328bar);
  OR2_X1 U325 ( .A1(n329), .A2(n330), .ZN(n110) );
  AND2_X1 U325bar ( .A1(n329bar), .A2(n330bar), .ZN(n110bar);
  OR2_X1 U326 ( .A1(n331), .A2(n332), .ZN(n330) );
  AND2_X1 U326bar ( .A1(n331bar), .A2(n332bar), .ZN(n330bar);
  OR2_X1 U327 ( .A1(n333), .A2(n334), .ZN(n332) );
  AND2_X1 U327bar ( .A1(n333bar), .A2(n334bar), .ZN(n332bar);
  OR2_X1 U328 ( .A1(in[127]), .A2(in[122]), .ZN(n334) );
  AND2_X1 U328bar ( .A1(inbar[127]), .A2(inbar[122]), .ZN(n334bar);
  OR2_X1 U329 ( .A1(in[156]), .A2(in[132]), .ZN(n333) );
  AND2_X1 U329bar ( .A1(inbar[156]), .A2(inbar[132]), .ZN(n333bar);
  OR2_X1 U330 ( .A1(n335), .A2(n336), .ZN(n331) );
  AND2_X1 U330bar ( .A1(n335bar), .A2(n336bar), .ZN(n331bar);
  OR2_X1 U331 ( .A1(in[159]), .A2(in[157]), .ZN(n336) );
  AND2_X1 U331bar ( .A1(inbar[159]), .A2(inbar[157]), .ZN(n336bar);
  OR2_X1 U332 ( .A1(in[185]), .A2(in[169]), .ZN(n335) );
  AND2_X1 U332bar ( .A1(inbar[185]), .A2(inbar[169]), .ZN(n335bar);
  OR2_X1 U333 ( .A1(n337), .A2(n338), .ZN(n329) );
  AND2_X1 U333bar ( .A1(n337bar), .A2(n338bar), .ZN(n329bar);
  OR2_X1 U334 ( .A1(n339), .A2(n340), .ZN(n338) );
  AND2_X1 U334bar ( .A1(n339bar), .A2(n340bar), .ZN(n338bar);
  OR2_X1 U335 ( .A1(in[239]), .A2(in[218]), .ZN(n340) );
  AND2_X1 U335bar ( .A1(inbar[239]), .A2(inbar[218]), .ZN(n340bar);
  OR2_X1 U336 ( .A1(in_13), .A2(in[87]), .ZN(n339) );
  AND2_X1 U336bar ( .A1(in_13bar), .A2(inbar[87]), .ZN(n339bar);
  OR2_X1 U337 ( .A1(n341), .A2(n342), .ZN(n337) );
  AND2_X1 U337bar ( .A1(n341bar), .A2(n342bar), .ZN(n337bar);
  OR2_X1 U338 ( .A1(in_72), .A2(in_70), .ZN(n342) );
  AND2_X1 U338bar ( .A1(in_72bar), .A2(in_70bar), .ZN(n342bar);
  OR2_X1 U339 ( .A1(in_80), .A2(in_74), .ZN(n341) );
  AND2_X1 U339bar ( .A1(in_80bar), .A2(in_74bar), .ZN(n341bar);
  OR2_X1 U340 ( .A1(n343), .A2(n344), .ZN(n31) );
  AND2_X1 U340bar ( .A1(n343bar), .A2(n344bar), .ZN(n31bar);
  OR2_X1 U341 ( .A1(n345), .A2(n346), .ZN(n344) );
  AND2_X1 U341bar ( .A1(n345bar), .A2(n346bar), .ZN(n344bar);
  OR2_X1 U342 ( .A1(n347), .A2(n348), .ZN(n346) );
  AND2_X1 U342bar ( .A1(n347bar), .A2(n348bar), .ZN(n346bar);
  OR2_X1 U343 ( .A1(in[146]), .A2(in[100]), .ZN(n348) );
  AND2_X1 U343bar ( .A1(inbar[146]), .A2(inbar[100]), .ZN(n348bar);
  OR2_X1 U344 ( .A1(in[168]), .A2(in[152]), .ZN(n347) );
  AND2_X1 U344bar ( .A1(inbar[168]), .A2(inbar[152]), .ZN(n347bar);
  OR2_X1 U345 ( .A1(n349), .A2(n350), .ZN(n345) );
  AND2_X1 U345bar ( .A1(n349bar), .A2(n350bar), .ZN(n345bar);
  OR2_X1 U346 ( .A1(in[199]), .A2(in[182]), .ZN(n350) );
  AND2_X1 U346bar ( .A1(inbar[199]), .A2(inbar[182]), .ZN(n350bar);
  OR2_X1 U347 ( .A1(in[236]), .A2(in[204]), .ZN(n349) );
  AND2_X1 U347bar ( .A1(inbar[236]), .A2(inbar[204]), .ZN(n349bar);
  OR2_X1 U348 ( .A1(n351), .A2(n352), .ZN(n343) );
  AND2_X1 U348bar ( .A1(n351bar), .A2(n352bar), .ZN(n343bar);
  OR2_X1 U349 ( .A1(n353), .A2(n354), .ZN(n352) );
  AND2_X1 U349bar ( .A1(n353bar), .A2(n354bar), .ZN(n352bar);
  OR2_X1 U350 ( .A1(in[89]), .A2(in[246]), .ZN(n354) );
  AND2_X1 U350bar ( .A1(inbar[89]), .A2(inbar[246]), .ZN(n354bar);
  OR2_X1 U351 ( .A1(in[95]), .A2(in[92]), .ZN(n353) );
  AND2_X1 U351bar ( .A1(inbar[95]), .A2(inbar[92]), .ZN(n353bar);
  OR2_X1 U352 ( .A1(n355), .A2(n356), .ZN(n351) );
  AND2_X1 U352bar ( .A1(n355bar), .A2(n356bar), .ZN(n351bar);
  OR2_X1 U353 ( .A1(in_22), .A2(in_16), .ZN(n356) );
  AND2_X1 U353bar ( .A1(in_22bar), .A2(in_16bar), .ZN(n356bar);
  OR2_X1 U354 ( .A1(in_51), .A2(in_49), .ZN(n355) );
  AND2_X1 U354bar ( .A1(in_51bar), .A2(in_49bar), .ZN(n355bar);
  OR2_X1 U355 ( .A1(n357), .A2(n358), .ZN(n251) );
  AND2_X1 U355bar ( .A1(n357bar), .A2(n358bar), .ZN(n251bar);
  OR2_X1 U356 ( .A1(in[158]), .A2(in[115]), .ZN(n358) );
  AND2_X1 U356bar ( .A1(inbar[158]), .A2(inbar[115]), .ZN(n358bar);
  OR2_X1 U357 ( .A1(in[163]), .A2(n359), .ZN(n357) );
  AND2_X1 U357bar ( .A1(inbar[163]), .A2(n359bar), .ZN(n357bar);
  OR2_X1 U358 ( .A1(in[206]), .A2(in[165]), .ZN(n359) );
  AND2_X1 U358bar ( .A1(inbar[206]), .A2(inbar[165]), .ZN(n359bar);
  OR2_X1 U359 ( .A1(n360), .A2(n361), .ZN(n249) );
  AND2_X1 U359bar ( .A1(n360bar), .A2(n361bar), .ZN(n249bar);
  OR2_X1 U360 ( .A1(n362), .A2(n363), .ZN(n361) );
  AND2_X1 U360bar ( .A1(n362bar), .A2(n363bar), .ZN(n361bar);
  OR2_X1 U361 ( .A1(in[213]), .A2(in[207]), .ZN(n363) );
  AND2_X1 U361bar ( .A1(inbar[213]), .A2(inbar[207]), .ZN(n363bar);
  OR2_X1 U362 ( .A1(in[215]), .A2(n364), .ZN(n362) );
  AND2_X1 U362bar ( .A1(inbar[215]), .A2(n364bar), .ZN(n362bar);
  OR2_X1 U363 ( .A1(in[230]), .A2(in[220]), .ZN(n364) );
  AND2_X1 U363bar ( .A1(inbar[230]), .A2(inbar[220]), .ZN(n364bar);
  OR2_X1 U364 ( .A1(n365), .A2(n366), .ZN(n360) );
  AND2_X1 U364bar ( .A1(n365bar), .A2(n366bar), .ZN(n360bar);
  OR2_X1 U365 ( .A1(in[251]), .A2(in[234]), .ZN(n366) );
  AND2_X1 U365bar ( .A1(inbar[251]), .A2(inbar[234]), .ZN(n366bar);
  OR2_X1 U366 ( .A1(in_17), .A2(n367), .ZN(n365) );
  AND2_X1 U366bar ( .A1(in_17bar), .A2(n367bar), .ZN(n365bar);
  OR2_X1 U367 ( .A1(in_65), .A2(in_56), .ZN(n367) );
  AND2_X1 U367bar ( .A1(in_65bar), .A2(in_56bar), .ZN(n367bar);
  OR2_X1 U368 ( .A1(n368), .A2(n369), .ZN(out[0]) );
  AND2_X1 U368bar ( .A1(n368bar), .A2(n369bar), .ZN(outbar[0]);
  OR2_X1 U369 ( .A1(n370), .A2(n371), .ZN(n369) );
  AND2_X1 U369bar ( .A1(n370bar), .A2(n371bar), .ZN(n369bar);
  OR2_X1 U370 ( .A1(n372), .A2(n373), .ZN(n371) );
  AND2_X1 U370bar ( .A1(n372bar), .A2(n373bar), .ZN(n371bar);
  OR2_X1 U371 ( .A1(n153), .A2(n188), .ZN(n373) );
  AND2_X1 U371bar ( .A1(n153bar), .A2(n188bar), .ZN(n373bar);
  OR2_X1 U372 ( .A1(n374), .A2(n375), .ZN(n188) );
  AND2_X1 U372bar ( .A1(n374bar), .A2(n375bar), .ZN(n188bar);
  OR2_X1 U373 ( .A1(n376), .A2(n377), .ZN(n375) );
  AND2_X1 U373bar ( .A1(n376bar), .A2(n377bar), .ZN(n375bar);
  OR2_X1 U374 ( .A1(n378), .A2(n379), .ZN(n377) );
  AND2_X1 U374bar ( .A1(n378bar), .A2(n379bar), .ZN(n377bar);
  OR2_X1 U375 ( .A1(in[135]), .A2(in[104]), .ZN(n379) );
  AND2_X1 U375bar ( .A1(inbar[135]), .A2(inbar[104]), .ZN(n379bar);
  OR2_X1 U376 ( .A1(in[188]), .A2(in[178]), .ZN(n378) );
  AND2_X1 U376bar ( .A1(inbar[188]), .A2(inbar[178]), .ZN(n378bar);
  OR2_X1 U377 ( .A1(n380), .A2(n381), .ZN(n376) );
  AND2_X1 U377bar ( .A1(n380bar), .A2(n381bar), .ZN(n376bar);
  OR2_X1 U378 ( .A1(in[217]), .A2(in[194]), .ZN(n381) );
  AND2_X1 U378bar ( .A1(inbar[217]), .A2(inbar[194]), .ZN(n381bar);
  OR2_X1 U379 ( .A1(in[237]), .A2(in[218]), .ZN(n380) );
  AND2_X1 U379bar ( .A1(inbar[237]), .A2(inbar[218]), .ZN(n380bar);
  OR2_X1 U380 ( .A1(n382), .A2(n383), .ZN(n374) );
  AND2_X1 U380bar ( .A1(n382bar), .A2(n383bar), .ZN(n374bar);
  OR2_X1 U381 ( .A1(n384), .A2(n385), .ZN(n383) );
  AND2_X1 U381bar ( .A1(n384bar), .A2(n385bar), .ZN(n383bar);
  OR2_X1 U382 ( .A1(in_2), .A2(in_10), .ZN(n385) );
  AND2_X1 U382bar ( .A1(in_2bar), .A2(in_10bar), .ZN(n385bar);
  OR2_X1 U383 ( .A1(in_47), .A2(in_22), .ZN(n384) );
  AND2_X1 U383bar ( .A1(in_47bar), .A2(in_22bar), .ZN(n384bar);
  OR2_X1 U384 ( .A1(n386), .A2(n387), .ZN(n382) );
  AND2_X1 U384bar ( .A1(n386bar), .A2(n387bar), .ZN(n382bar);
  OR2_X1 U385 ( .A1(in_56), .A2(in_54), .ZN(n387) );
  AND2_X1 U385bar ( .A1(in_56bar), .A2(in_54bar), .ZN(n387bar);
  OR2_X1 U386 ( .A1(in_63), .A2(in_61), .ZN(n386) );
  AND2_X1 U386bar ( .A1(in_63bar), .A2(in_61bar), .ZN(n386bar);
  OR2_X1 U387 ( .A1(n388), .A2(n389), .ZN(n153) );
  AND2_X1 U387bar ( .A1(n388bar), .A2(n389bar), .ZN(n153bar);
  OR2_X1 U388 ( .A1(n390), .A2(n391), .ZN(n389) );
  AND2_X1 U388bar ( .A1(n390bar), .A2(n391bar), .ZN(n389bar);
  OR2_X1 U389 ( .A1(n392), .A2(n393), .ZN(n391) );
  AND2_X1 U389bar ( .A1(n392bar), .A2(n393bar), .ZN(n391bar);
  OR2_X1 U390 ( .A1(in[158]), .A2(in[142]), .ZN(n393) );
  AND2_X1 U390bar ( .A1(inbar[158]), .A2(inbar[142]), .ZN(n393bar);
  OR2_X1 U391 ( .A1(in[175]), .A2(in[164]), .ZN(n392) );
  AND2_X1 U391bar ( .A1(inbar[175]), .A2(inbar[164]), .ZN(n392bar);
  OR2_X1 U392 ( .A1(n394), .A2(n395), .ZN(n390) );
  AND2_X1 U392bar ( .A1(n394bar), .A2(n395bar), .ZN(n390bar);
  OR2_X1 U393 ( .A1(in[228]), .A2(in[204]), .ZN(n395) );
  AND2_X1 U393bar ( .A1(inbar[228]), .A2(inbar[204]), .ZN(n395bar);
  OR2_X1 U394 ( .A1(in[91]), .A2(in[87]), .ZN(n394) );
  AND2_X1 U394bar ( .A1(inbar[91]), .A2(inbar[87]), .ZN(n394bar);
  OR2_X1 U395 ( .A1(n396), .A2(n397), .ZN(n388) );
  AND2_X1 U395bar ( .A1(n396bar), .A2(n397bar), .ZN(n388bar);
  OR2_X1 U396 ( .A1(n398), .A2(n399), .ZN(n397) );
  AND2_X1 U396bar ( .A1(n398bar), .A2(n399bar), .ZN(n397bar);
  OR2_X1 U397 ( .A1(in_21), .A2(in_11), .ZN(n399) );
  AND2_X1 U397bar ( .A1(in_21bar), .A2(in_11bar), .ZN(n399bar);
  OR2_X1 U398 ( .A1(in_5), .A2(in_3), .ZN(n398) );
  AND2_X1 U398bar ( .A1(in_5bar), .A2(in_3bar), .ZN(n398bar);
  OR2_X1 U399 ( .A1(n400), .A2(n401), .ZN(n396) );
  AND2_X1 U399bar ( .A1(n400bar), .A2(n401bar), .ZN(n396bar);
  OR2_X1 U400 ( .A1(in_68), .A2(in_64), .ZN(n401) );
  AND2_X1 U400bar ( .A1(in_68bar), .A2(in_64bar), .ZN(n401bar);
  OR2_X1 U401 ( .A1(in_76), .A2(in_73), .ZN(n400) );
  AND2_X1 U401bar ( .A1(in_76bar), .A2(in_73bar), .ZN(n400bar);
  OR2_X1 U402 ( .A1(n195), .A2(n402), .ZN(n372) );
  AND2_X1 U402bar ( .A1(n195bar), .A2(n402bar), .ZN(n372bar);
  OR2_X1 U403 ( .A1(in[100]), .A2(n8), .ZN(n402) );
  AND2_X1 U403bar ( .A1(inbar[100]), .A2(n8bar), .ZN(n402bar);
  OR2_X1 U404 ( .A1(n403), .A2(n404), .ZN(n8) );
  AND2_X1 U404bar ( .A1(n403bar), .A2(n404bar), .ZN(n8bar);
  OR2_X1 U405 ( .A1(n405), .A2(n406), .ZN(n404) );
  AND2_X1 U405bar ( .A1(n405bar), .A2(n406bar), .ZN(n404bar);
  OR2_X1 U406 ( .A1(n407), .A2(n408), .ZN(n406) );
  AND2_X1 U406bar ( .A1(n407bar), .A2(n408bar), .ZN(n406bar);
  OR2_X1 U407 ( .A1(n156), .A2(n223), .ZN(n408) );
  AND2_X1 U407bar ( .A1(n156bar), .A2(n223bar), .ZN(n408bar);
  OR2_X1 U408 ( .A1(n409), .A2(n410), .ZN(n223) );
  AND2_X1 U408bar ( .A1(n409bar), .A2(n410bar), .ZN(n223bar);
  OR2_X1 U409 ( .A1(n411), .A2(n412), .ZN(n410) );
  AND2_X1 U409bar ( .A1(n411bar), .A2(n412bar), .ZN(n410bar);
  OR2_X1 U410 ( .A1(n413), .A2(n414), .ZN(n412) );
  AND2_X1 U410bar ( .A1(n413bar), .A2(n414bar), .ZN(n412bar);
  OR2_X1 U411 ( .A1(in[119]), .A2(in[103]), .ZN(n414) );
  AND2_X1 U411bar ( .A1(inbar[119]), .A2(inbar[103]), .ZN(n414bar);
  OR2_X1 U412 ( .A1(in[137]), .A2(in[133]), .ZN(n413) );
  AND2_X1 U412bar ( .A1(inbar[137]), .A2(inbar[133]), .ZN(n413bar);
  OR2_X1 U413 ( .A1(n415), .A2(n416), .ZN(n411) );
  AND2_X1 U413bar ( .A1(n415bar), .A2(n416bar), .ZN(n411bar);
  OR2_X1 U414 ( .A1(in[176]), .A2(in[173]), .ZN(n416) );
  AND2_X1 U414bar ( .A1(inbar[176]), .A2(inbar[173]), .ZN(n416bar);
  OR2_X1 U415 ( .A1(in[210]), .A2(in[181]), .ZN(n415) );
  AND2_X1 U415bar ( .A1(inbar[210]), .A2(inbar[181]), .ZN(n415bar);
  OR2_X1 U416 ( .A1(n417), .A2(n418), .ZN(n409) );
  AND2_X1 U416bar ( .A1(n417bar), .A2(n418bar), .ZN(n409bar);
  OR2_X1 U417 ( .A1(n419), .A2(n420), .ZN(n418) );
  AND2_X1 U417bar ( .A1(n419bar), .A2(n420bar), .ZN(n418bar);
  OR2_X1 U418 ( .A1(in_13), .A2(in[234]), .ZN(n420) );
  AND2_X1 U418bar ( .A1(in_13bar), .A2(inbar[234]), .ZN(n420bar);
  OR2_X1 U419 ( .A1(in_38), .A2(in_32), .ZN(n419) );
  AND2_X1 U419bar ( .A1(in_38bar), .A2(in_32bar), .ZN(n419bar);
  OR2_X1 U420 ( .A1(n421), .A2(n422), .ZN(n417) );
  AND2_X1 U420bar ( .A1(n421bar), .A2(n422bar), .ZN(n417bar);
  OR2_X1 U421 ( .A1(in_42), .A2(in_41), .ZN(n422) );
  AND2_X1 U421bar ( .A1(in_42bar), .A2(in_41bar), .ZN(n422bar);
  OR2_X1 U422 ( .A1(in_7), .A2(in_49), .ZN(n421) );
  AND2_X1 U422bar ( .A1(in_7bar), .A2(in_49bar), .ZN(n421bar);
  OR2_X1 U423 ( .A1(n423), .A2(n424), .ZN(n156) );
  AND2_X1 U423bar ( .A1(n423bar), .A2(n424bar), .ZN(n156bar);
  OR2_X1 U424 ( .A1(n425), .A2(n426), .ZN(n424) );
  AND2_X1 U424bar ( .A1(n425bar), .A2(n426bar), .ZN(n424bar);
  OR2_X1 U425 ( .A1(n427), .A2(n428), .ZN(n426) );
  AND2_X1 U425bar ( .A1(n427bar), .A2(n428bar), .ZN(n426bar);
  OR2_X1 U426 ( .A1(in[159]), .A2(in[105]), .ZN(n428) );
  AND2_X1 U426bar ( .A1(inbar[159]), .A2(inbar[105]), .ZN(n428bar);
  OR2_X1 U427 ( .A1(in[206]), .A2(in[183]), .ZN(n427) );
  AND2_X1 U427bar ( .A1(inbar[206]), .A2(inbar[183]), .ZN(n427bar);
  OR2_X1 U428 ( .A1(n429), .A2(n430), .ZN(n425) );
  AND2_X1 U428bar ( .A1(n429bar), .A2(n430bar), .ZN(n425bar);
  OR2_X1 U429 ( .A1(in[229]), .A2(in[219]), .ZN(n430) );
  AND2_X1 U429bar ( .A1(inbar[229]), .A2(inbar[219]), .ZN(n430bar);
  OR2_X1 U430 ( .A1(in[235]), .A2(in[232]), .ZN(n429) );
  AND2_X1 U430bar ( .A1(inbar[235]), .A2(inbar[232]), .ZN(n429bar);
  OR2_X1 U431 ( .A1(n431), .A2(n432), .ZN(n423) );
  AND2_X1 U431bar ( .A1(n431bar), .A2(n432bar), .ZN(n423bar);
  OR2_X1 U432 ( .A1(n433), .A2(n434), .ZN(n432) );
  AND2_X1 U432bar ( .A1(n433bar), .A2(n434bar), .ZN(n432bar);
  OR2_X1 U433 ( .A1(in[249]), .A2(in[242]), .ZN(n434) );
  AND2_X1 U433bar ( .A1(inbar[249]), .A2(inbar[242]), .ZN(n434bar);
  OR2_X1 U434 ( .A1(in[89]), .A2(in[254]), .ZN(n433) );
  AND2_X1 U434bar ( .A1(inbar[89]), .A2(inbar[254]), .ZN(n433bar);
  OR2_X1 U435 ( .A1(n435), .A2(n436), .ZN(n431) );
  AND2_X1 U435bar ( .A1(n435bar), .A2(n436bar), .ZN(n431bar);
  OR2_X1 U436 ( .A1(in_14), .A2(in[99]), .ZN(n436) );
  AND2_X1 U436bar ( .A1(in_14bar), .A2(inbar[99]), .ZN(n436bar);
  OR2_X1 U437 ( .A1(in_60), .A2(in_18), .ZN(n435) );
  AND2_X1 U437bar ( .A1(in_60bar), .A2(in_18bar), .ZN(n435bar);
  OR2_X1 U438 ( .A1(in[113]), .A2(n210), .ZN(n407) );
  AND2_X1 U438bar ( .A1(inbar[113]), .A2(n210bar), .ZN(n407bar);
  OR2_X1 U439 ( .A1(n437), .A2(n438), .ZN(n210) );
  AND2_X1 U439bar ( .A1(n437bar), .A2(n438bar), .ZN(n210bar);
  OR2_X1 U440 ( .A1(n439), .A2(n440), .ZN(n438) );
  AND2_X1 U440bar ( .A1(n439bar), .A2(n440bar), .ZN(n438bar);
  OR2_X1 U441 ( .A1(n441), .A2(n442), .ZN(n440) );
  AND2_X1 U441bar ( .A1(n441bar), .A2(n442bar), .ZN(n440bar);
  OR2_X1 U442 ( .A1(in[115]), .A2(in[110]), .ZN(n442) );
  AND2_X1 U442bar ( .A1(inbar[115]), .A2(inbar[110]), .ZN(n442bar);
  OR2_X1 U443 ( .A1(in[125]), .A2(in[117]), .ZN(n441) );
  AND2_X1 U443bar ( .A1(inbar[125]), .A2(inbar[117]), .ZN(n441bar);
  OR2_X1 U444 ( .A1(n443), .A2(n444), .ZN(n439) );
  AND2_X1 U444bar ( .A1(n443bar), .A2(n444bar), .ZN(n439bar);
  OR2_X1 U445 ( .A1(in[180]), .A2(in[128]), .ZN(n444) );
  AND2_X1 U445bar ( .A1(inbar[180]), .A2(inbar[128]), .ZN(n444bar);
  OR2_X1 U446 ( .A1(in[205]), .A2(in[201]), .ZN(n443) );
  AND2_X1 U446bar ( .A1(inbar[205]), .A2(inbar[201]), .ZN(n443bar);
  OR2_X1 U447 ( .A1(n445), .A2(n446), .ZN(n437) );
  AND2_X1 U447bar ( .A1(n445bar), .A2(n446bar), .ZN(n437bar);
  OR2_X1 U448 ( .A1(n447), .A2(n448), .ZN(n446) );
  AND2_X1 U448bar ( .A1(n447bar), .A2(n448bar), .ZN(n446bar);
  OR2_X1 U449 ( .A1(in[244]), .A2(in[239]), .ZN(n448) );
  AND2_X1 U449bar ( .A1(inbar[244]), .A2(inbar[239]), .ZN(n448bar);
  OR2_X1 U450 ( .A1(in[95]), .A2(in[83]), .ZN(n447) );
  AND2_X1 U450bar ( .A1(inbar[95]), .A2(inbar[83]), .ZN(n447bar);
  OR2_X1 U451 ( .A1(n449), .A2(n450), .ZN(n445) );
  AND2_X1 U451bar ( .A1(n449bar), .A2(n450bar), .ZN(n445bar);
  OR2_X1 U452 ( .A1(in_24), .A2(in[97]), .ZN(n450) );
  AND2_X1 U452bar ( .A1(in_24bar), .A2(inbar[97]), .ZN(n450bar);
  OR2_X1 U453 ( .A1(in_33), .A2(in_27), .ZN(n449) );
  AND2_X1 U453bar ( .A1(in_33bar), .A2(in_27bar), .ZN(n449bar);
  OR2_X1 U454 ( .A1(n451), .A2(n452), .ZN(n405) );
  AND2_X1 U454bar ( .A1(n451bar), .A2(n452bar), .ZN(n405bar);
  OR2_X1 U455 ( .A1(in[145]), .A2(in[126]), .ZN(n452) );
  AND2_X1 U455bar ( .A1(inbar[145]), .A2(inbar[126]), .ZN(n452bar);
  OR2_X1 U456 ( .A1(in[169]), .A2(n453), .ZN(n451) );
  AND2_X1 U456bar ( .A1(inbar[169]), .A2(n453bar), .ZN(n451bar);
  OR2_X1 U457 ( .A1(in[221]), .A2(in[172]), .ZN(n453) );
  AND2_X1 U457bar ( .A1(inbar[221]), .A2(inbar[172]), .ZN(n453bar);
  OR2_X1 U458 ( .A1(n454), .A2(n455), .ZN(n403) );
  AND2_X1 U458bar ( .A1(n454bar), .A2(n455bar), .ZN(n403bar);
  OR2_X1 U459 ( .A1(n456), .A2(n457), .ZN(n455) );
  AND2_X1 U459bar ( .A1(n456bar), .A2(n457bar), .ZN(n455bar);
  OR2_X1 U460 ( .A1(in[241]), .A2(in[224]), .ZN(n457) );
  AND2_X1 U460bar ( .A1(inbar[241]), .A2(inbar[224]), .ZN(n457bar);
  OR2_X1 U461 ( .A1(in[86]), .A2(n458), .ZN(n456) );
  AND2_X1 U461bar ( .A1(inbar[86]), .A2(n458bar), .ZN(n456bar);
  OR2_X1 U462 ( .A1(in_43), .A2(in_34), .ZN(n458) );
  AND2_X1 U462bar ( .A1(in_43bar), .A2(in_34bar), .ZN(n458bar);
  OR2_X1 U463 ( .A1(n459), .A2(n460), .ZN(n454) );
  AND2_X1 U463bar ( .A1(n459bar), .A2(n460bar), .ZN(n454bar);
  OR2_X1 U464 ( .A1(in_65), .A2(in_51), .ZN(n460) );
  AND2_X1 U464bar ( .A1(in_65bar), .A2(in_51bar), .ZN(n460bar);
  OR2_X1 U465 ( .A1(in_75), .A2(n461), .ZN(n459) );
  AND2_X1 U465bar ( .A1(in_75bar), .A2(n461bar), .ZN(n459bar);
  OR2_X1 U466 ( .A1(in_81), .A2(in_77), .ZN(n461) );
  AND2_X1 U466bar ( .A1(in_81bar), .A2(in_77bar), .ZN(n461bar);
  OR2_X1 U467 ( .A1(n462), .A2(n463), .ZN(n195) );
  AND2_X1 U467bar ( .A1(n462bar), .A2(n463bar), .ZN(n195bar);
  OR2_X1 U468 ( .A1(n464), .A2(n465), .ZN(n463) );
  AND2_X1 U468bar ( .A1(n464bar), .A2(n465bar), .ZN(n463bar);
  OR2_X1 U469 ( .A1(n466), .A2(n467), .ZN(n465) );
  AND2_X1 U469bar ( .A1(n466bar), .A2(n467bar), .ZN(n465bar);
  OR2_X1 U470 ( .A1(in[107]), .A2(in[101]), .ZN(n467) );
  AND2_X1 U470bar ( .A1(inbar[107]), .A2(inbar[101]), .ZN(n467bar);
  OR2_X1 U471 ( .A1(in[139]), .A2(in[132]), .ZN(n466) );
  AND2_X1 U471bar ( .A1(inbar[139]), .A2(inbar[132]), .ZN(n466bar);
  OR2_X1 U472 ( .A1(n468), .A2(n469), .ZN(n464) );
  AND2_X1 U472bar ( .A1(n468bar), .A2(n469bar), .ZN(n464bar);
  OR2_X1 U473 ( .A1(in[146]), .A2(in[141]), .ZN(n469) );
  AND2_X1 U473bar ( .A1(inbar[146]), .A2(inbar[141]), .ZN(n469bar);
  OR2_X1 U474 ( .A1(in[203]), .A2(in[179]), .ZN(n468) );
  AND2_X1 U474bar ( .A1(inbar[203]), .A2(inbar[179]), .ZN(n468bar);
  OR2_X1 U475 ( .A1(n470), .A2(n471), .ZN(n462) );
  AND2_X1 U475bar ( .A1(n470bar), .A2(n471bar), .ZN(n462bar);
  OR2_X1 U476 ( .A1(n472), .A2(n473), .ZN(n471) );
  AND2_X1 U476bar ( .A1(n472bar), .A2(n473bar), .ZN(n471bar);
  OR2_X1 U477 ( .A1(in[243]), .A2(in[222]), .ZN(n473) );
  AND2_X1 U477bar ( .A1(inbar[243]), .A2(inbar[222]), .ZN(n473bar);
  OR2_X1 U478 ( .A1(in[251]), .A2(in[250]), .ZN(n472) );
  AND2_X1 U478bar ( .A1(inbar[251]), .A2(inbar[250]), .ZN(n472bar);
  OR2_X1 U479 ( .A1(n474), .A2(n475), .ZN(n470) );
  AND2_X1 U479bar ( .A1(n474bar), .A2(n475bar), .ZN(n470bar);
  OR2_X1 U480 ( .A1(in_37), .A2(in_19), .ZN(n475) );
  AND2_X1 U480bar ( .A1(in_37bar), .A2(in_19bar), .ZN(n475bar);
  OR2_X1 U481 ( .A1(in_78), .A2(in_6), .ZN(n474) );
  AND2_X1 U481bar ( .A1(in_78bar), .A2(in_6bar), .ZN(n474bar);
  OR2_X1 U482 ( .A1(n476), .A2(n477), .ZN(n370) );
  AND2_X1 U482bar ( .A1(n476bar), .A2(n477bar), .ZN(n370bar);
  OR2_X1 U483 ( .A1(in[112]), .A2(in[102]), .ZN(n477) );
  AND2_X1 U483bar ( .A1(inbar[112]), .A2(inbar[102]), .ZN(n477bar);
  OR2_X1 U484 ( .A1(in[123]), .A2(n478), .ZN(n476) );
  AND2_X1 U484bar ( .A1(inbar[123]), .A2(n478bar), .ZN(n476bar);
  OR2_X1 U485 ( .A1(in[143]), .A2(in[130]), .ZN(n478) );
  AND2_X1 U485bar ( .A1(inbar[143]), .A2(inbar[130]), .ZN(n478bar);
  OR2_X1 U486 ( .A1(n479), .A2(n480), .ZN(n368) );
  AND2_X1 U486bar ( .A1(n479bar), .A2(n480bar), .ZN(n368bar);
  OR2_X1 U487 ( .A1(n481), .A2(n482), .ZN(n480) );
  AND2_X1 U487bar ( .A1(n481bar), .A2(n482bar), .ZN(n480bar);
  OR2_X1 U488 ( .A1(in[216]), .A2(in[213]), .ZN(n482) );
  AND2_X1 U488bar ( .A1(inbar[216]), .A2(inbar[213]), .ZN(n482bar);
  OR2_X1 U489 ( .A1(in[227]), .A2(n483), .ZN(n481) );
  AND2_X1 U489bar ( .A1(inbar[227]), .A2(n483bar), .ZN(n481bar);
  OR2_X1 U490 ( .A1(in_0), .A2(in[248]), .ZN(n483) );
  AND2_X1 U490bar ( .A1(in_0bar), .A2(inbar[248]), .ZN(n483bar);
  OR2_X1 U491 ( .A1(n484), .A2(n485), .ZN(n479) );
  AND2_X1 U491bar ( .A1(n484bar), .A2(n485bar), .ZN(n479bar);
  OR2_X1 U492 ( .A1(in_46), .A2(in_44), .ZN(n485) );
  AND2_X1 U492bar ( .A1(in_46bar), .A2(in_44bar), .ZN(n485bar);
  OR2_X1 U493 ( .A1(in_50), .A2(n486), .ZN(n484) );
  AND2_X1 U493bar ( .A1(in_50bar), .A2(n486bar), .ZN(n484bar);
  OR2_X1 U494 ( .A1(in_9), .A2(in_80), .ZN(n486) );
  AND2_X1 U494bar ( .A1(in_9bar), .A2(in_80bar), .ZN(n486bar);
endmodule




module sBox_0 ( in, out );
  input [7:0] in;
  //input_done

  output [7:0] out;
  //output_done

  wire   [255:0] decodeOut;
  //wire_done

  decode_0 dec ( .in(in), .out(decodeOut) );
  encode_0 enc ( .in(decodeOut), .out(out) );
endmodule


module scale2_0 ( in, out );
  input [7:0] in;
  //input_done

  output [7:0] out;
  //output_done

  wire   in_0, \in[6] , \in[5] , \in[4] , \in[1] , \in[7] , n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10;
  //wire_done

  assign in_0 = in[0];
  assign out[7] = \in[6] ;
  assign \in[6]  = in[6];
  assign out[6] = \in[5] ;
  assign \in[5]  = in[5];
  assign out[5] = \in[4] ;
  assign \in[4]  = in[4];
  assign out[2] = \in[1] ;
  assign \in[1]  = in[1];
  assign out[0] = \in[7] ;
  assign \in[7]  = in[7];

  INV_X1 U1 ( .A(\in[7]), .ZN(n1) );
  INV_X1 U2 ( .A(in[3]), .ZN(n2) );
  INV_X1 U3 ( .A(in[2]), .ZN(n3) );
  INV_X1 U4 ( .A(in_0), .ZN(n4) );
  OR2_X1 U5 ( .A1(n5), .A2(n6), .ZN(out[4]) );
  AND2_X1 U6 ( .A1(in[3]), .A2(n1), .ZN(n6) );
  AND2_X1 U7 ( .A1(\in[7]), .A2(n2), .ZN(n5) );
  OR2_X1 U8 ( .A1(n7), .A2(n8), .ZN(out[3]) );
  AND2_X1 U9 ( .A1(in[2]), .A2(n1), .ZN(n8) );
  AND2_X1 U10 ( .A1(\in[7]), .A2(n3), .ZN(n7) );
  OR2_X1 U11 ( .A1(n9), .A2(n10), .ZN(out[1]) );
  AND2_X1 U12 ( .A1(in_0), .A2(n1), .ZN(n10) );
  AND2_X1 U13 ( .A1(\in[7]), .A2(n4), .ZN(n9) );
endmodule


module byteXor_0 ( a, b, y );
  input [7:0] a;
  input [7:0] b;
  //input_done

  output [7:0] y;
  //output_done

  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32;
  //wire_done

  INV_X1 U1 ( .A(n18), .ZN(n1) );
  INV_X1 U2 ( .A(a[7]), .ZN(n2) );
  INV_X1 U3 ( .A(n20), .ZN(n3) );
  INV_X1 U4 ( .A(a[6]), .ZN(n4) );
  INV_X1 U5 ( .A(n22), .ZN(n5) );
  INV_X1 U6 ( .A(a[5]), .ZN(n6) );
  INV_X1 U7 ( .A(n24), .ZN(n7) );
  INV_X1 U8 ( .A(a[4]), .ZN(n8) );
  INV_X1 U9 ( .A(n26), .ZN(n9) );
  INV_X1 U10 ( .A(a[3]), .ZN(n10) );
  INV_X1 U11 ( .A(n28), .ZN(n11) );
  INV_X1 U12 ( .A(a[2]), .ZN(n12) );
  INV_X1 U13 ( .A(n30), .ZN(n13) );
  INV_X1 U14 ( .A(a[1]), .ZN(n14) );
  INV_X1 U15 ( .A(n32), .ZN(n15) );
  INV_X1 U16 ( .A(a[0]), .ZN(n16) );
  OR2_X1 U17 ( .A1(n17), .A2(n1), .ZN(y[7]) );
  OR2_X1 U18 ( .A1(n2), .A2(b[7]), .ZN(n18) );
  AND2_X1 U19 ( .A1(b[7]), .A2(n2), .ZN(n17) );
  OR2_X1 U20 ( .A1(n19), .A2(n3), .ZN(y[6]) );
  OR2_X1 U21 ( .A1(n4), .A2(b[6]), .ZN(n20) );
  AND2_X1 U22 ( .A1(b[6]), .A2(n4), .ZN(n19) );
  OR2_X1 U23 ( .A1(n21), .A2(n5), .ZN(y[5]) );
  OR2_X1 U24 ( .A1(n6), .A2(b[5]), .ZN(n22) );
  AND2_X1 U25 ( .A1(b[5]), .A2(n6), .ZN(n21) );
  OR2_X1 U26 ( .A1(n23), .A2(n7), .ZN(y[4]) );
  OR2_X1 U27 ( .A1(n8), .A2(b[4]), .ZN(n24) );
  AND2_X1 U28 ( .A1(b[4]), .A2(n8), .ZN(n23) );
  OR2_X1 U29 ( .A1(n25), .A2(n9), .ZN(y[3]) );
  OR2_X1 U30 ( .A1(n10), .A2(b[3]), .ZN(n26) );
  AND2_X1 U31 ( .A1(b[3]), .A2(n10), .ZN(n25) );
  OR2_X1 U32 ( .A1(n27), .A2(n11), .ZN(y[2]) );
  OR2_X1 U33 ( .A1(n12), .A2(b[2]), .ZN(n28) );
  AND2_X1 U34 ( .A1(b[2]), .A2(n12), .ZN(n27) );
  OR2_X1 U35 ( .A1(n29), .A2(n13), .ZN(y[1]) );
  OR2_X1 U36 ( .A1(n14), .A2(b[1]), .ZN(n30) );
  AND2_X1 U37 ( .A1(b[1]), .A2(n14), .ZN(n29) );
  OR2_X1 U38 ( .A1(n31), .A2(n15), .ZN(y[0]) );
  OR2_X1 U39 ( .A1(n16), .A2(b[0]), .ZN(n32) );
  AND2_X1 U40 ( .A1(b[0]), .A2(n16), .ZN(n31) );
endmodule


module byteXor4_0 ( a, b, c, d, y );
  input [7:0] a;
  input [7:0] b;
  input [7:0] c;
  input [7:0] d;
  //input_done

  output [7:0] y;
  //output_done

  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112;
  //wire_done

  INV_X1 U1 ( .A(n50), .ZN(n1) );
  INV_X1 U2 ( .A(a[7]), .ZN(n2) );
  INV_X1 U3 ( .A(n58), .ZN(n3) );
  INV_X1 U4 ( .A(a[6]), .ZN(n4) );
  INV_X1 U5 ( .A(n66), .ZN(n5) );
  INV_X1 U6 ( .A(a[5]), .ZN(n6) );
  INV_X1 U7 ( .A(n74), .ZN(n7) );
  INV_X1 U8 ( .A(a[4]), .ZN(n8) );
  INV_X1 U9 ( .A(n82), .ZN(n9) );
  INV_X1 U10 ( .A(a[3]), .ZN(n10) );
  INV_X1 U11 ( .A(n90), .ZN(n11) );
  INV_X1 U12 ( .A(a[2]), .ZN(n12) );
  INV_X1 U13 ( .A(n98), .ZN(n13) );
  INV_X1 U14 ( .A(a[1]), .ZN(n14) );
  INV_X1 U15 ( .A(n106), .ZN(n15) );
  INV_X1 U16 ( .A(a[0]), .ZN(n16) );
  INV_X1 U17 ( .A(b[7]), .ZN(n17) );
  INV_X1 U18 ( .A(b[6]), .ZN(n18) );
  INV_X1 U19 ( .A(b[5]), .ZN(n19) );
  INV_X1 U20 ( .A(b[4]), .ZN(n20) );
  INV_X1 U21 ( .A(b[3]), .ZN(n21) );
  INV_X1 U22 ( .A(b[2]), .ZN(n22) );
  INV_X1 U23 ( .A(b[1]), .ZN(n23) );
  INV_X1 U24 ( .A(b[0]), .ZN(n24) );
  INV_X1 U25 ( .A(n54), .ZN(n25) );
  INV_X1 U26 ( .A(c[7]), .ZN(n26) );
  INV_X1 U27 ( .A(n62), .ZN(n27) );
  INV_X1 U28 ( .A(c[6]), .ZN(n28) );
  INV_X1 U29 ( .A(n70), .ZN(n29) );
  INV_X1 U30 ( .A(c[5]), .ZN(n30) );
  INV_X1 U31 ( .A(n78), .ZN(n31) );
  INV_X1 U32 ( .A(c[4]), .ZN(n32) );
  INV_X1 U33 ( .A(n86), .ZN(n33) );
  INV_X1 U34 ( .A(c[3]), .ZN(n34) );
  INV_X1 U35 ( .A(n94), .ZN(n35) );
  INV_X1 U36 ( .A(c[2]), .ZN(n36) );
  INV_X1 U37 ( .A(n102), .ZN(n37) );
  INV_X1 U38 ( .A(c[1]), .ZN(n38) );
  INV_X1 U39 ( .A(n110), .ZN(n39) );
  INV_X1 U40 ( .A(c[0]), .ZN(n40) );
  INV_X1 U41 ( .A(d[7]), .ZN(n41) );
  INV_X1 U42 ( .A(d[6]), .ZN(n42) );
  INV_X1 U43 ( .A(d[5]), .ZN(n43) );
  INV_X1 U44 ( .A(d[4]), .ZN(n44) );
  INV_X1 U45 ( .A(d[3]), .ZN(n45) );
  INV_X1 U46 ( .A(d[2]), .ZN(n46) );
  INV_X1 U47 ( .A(d[1]), .ZN(n47) );
  INV_X1 U48 ( .A(d[0]), .ZN(n48) );
  OR2_X1 U49 ( .A1(n49), .A2(n1), .ZN(y[7]) );
  OR2_X1 U50 ( .A1(n51), .A2(n25), .ZN(n50) );
  AND2_X1 U51 ( .A1(n25), .A2(n51), .ZN(n49) );
  AND2_X1 U52 ( .A1(n52), .A2(n53), .ZN(n51) );
  OR2_X1 U53 ( .A1(n2), .A2(b[7]), .ZN(n53) );
  OR2_X1 U54 ( .A1(n17), .A2(a[7]), .ZN(n52) );
  AND2_X1 U55 ( .A1(n55), .A2(n56), .ZN(n54) );
  OR2_X1 U56 ( .A1(n26), .A2(d[7]), .ZN(n56) );
  OR2_X1 U57 ( .A1(n41), .A2(c[7]), .ZN(n55) );
  OR2_X1 U58 ( .A1(n57), .A2(n3), .ZN(y[6]) );
  OR2_X1 U59 ( .A1(n59), .A2(n27), .ZN(n58) );
  AND2_X1 U60 ( .A1(n27), .A2(n59), .ZN(n57) );
  AND2_X1 U61 ( .A1(n60), .A2(n61), .ZN(n59) );
  OR2_X1 U62 ( .A1(n4), .A2(b[6]), .ZN(n61) );
  OR2_X1 U63 ( .A1(n18), .A2(a[6]), .ZN(n60) );
  AND2_X1 U64 ( .A1(n63), .A2(n64), .ZN(n62) );
  OR2_X1 U65 ( .A1(n28), .A2(d[6]), .ZN(n64) );
  OR2_X1 U66 ( .A1(n42), .A2(c[6]), .ZN(n63) );
  OR2_X1 U67 ( .A1(n65), .A2(n5), .ZN(y[5]) );
  OR2_X1 U68 ( .A1(n67), .A2(n29), .ZN(n66) );
  AND2_X1 U69 ( .A1(n29), .A2(n67), .ZN(n65) );
  AND2_X1 U70 ( .A1(n68), .A2(n69), .ZN(n67) );
  OR2_X1 U71 ( .A1(n6), .A2(b[5]), .ZN(n69) );
  OR2_X1 U72 ( .A1(n19), .A2(a[5]), .ZN(n68) );
  AND2_X1 U73 ( .A1(n71), .A2(n72), .ZN(n70) );
  OR2_X1 U74 ( .A1(n30), .A2(d[5]), .ZN(n72) );
  OR2_X1 U75 ( .A1(n43), .A2(c[5]), .ZN(n71) );
  OR2_X1 U76 ( .A1(n73), .A2(n7), .ZN(y[4]) );
  OR2_X1 U77 ( .A1(n75), .A2(n31), .ZN(n74) );
  AND2_X1 U78 ( .A1(n31), .A2(n75), .ZN(n73) );
  AND2_X1 U79 ( .A1(n76), .A2(n77), .ZN(n75) );
  OR2_X1 U80 ( .A1(n8), .A2(b[4]), .ZN(n77) );
  OR2_X1 U81 ( .A1(n20), .A2(a[4]), .ZN(n76) );
  AND2_X1 U82 ( .A1(n79), .A2(n80), .ZN(n78) );
  OR2_X1 U83 ( .A1(n32), .A2(d[4]), .ZN(n80) );
  OR2_X1 U84 ( .A1(n44), .A2(c[4]), .ZN(n79) );
  OR2_X1 U85 ( .A1(n81), .A2(n9), .ZN(y[3]) );
  OR2_X1 U86 ( .A1(n83), .A2(n33), .ZN(n82) );
  AND2_X1 U87 ( .A1(n33), .A2(n83), .ZN(n81) );
  AND2_X1 U88 ( .A1(n84), .A2(n85), .ZN(n83) );
  OR2_X1 U89 ( .A1(n10), .A2(b[3]), .ZN(n85) );
  OR2_X1 U90 ( .A1(n21), .A2(a[3]), .ZN(n84) );
  AND2_X1 U91 ( .A1(n87), .A2(n88), .ZN(n86) );
  OR2_X1 U92 ( .A1(n34), .A2(d[3]), .ZN(n88) );
  OR2_X1 U93 ( .A1(n45), .A2(c[3]), .ZN(n87) );
  OR2_X1 U94 ( .A1(n89), .A2(n11), .ZN(y[2]) );
  OR2_X1 U95 ( .A1(n91), .A2(n35), .ZN(n90) );
  AND2_X1 U96 ( .A1(n35), .A2(n91), .ZN(n89) );
  AND2_X1 U97 ( .A1(n92), .A2(n93), .ZN(n91) );
  OR2_X1 U98 ( .A1(n12), .A2(b[2]), .ZN(n93) );
  OR2_X1 U99 ( .A1(n22), .A2(a[2]), .ZN(n92) );
  AND2_X1 U100 ( .A1(n95), .A2(n96), .ZN(n94) );
  OR2_X1 U101 ( .A1(n36), .A2(d[2]), .ZN(n96) );
  OR2_X1 U102 ( .A1(n46), .A2(c[2]), .ZN(n95) );
  OR2_X1 U103 ( .A1(n97), .A2(n13), .ZN(y[1]) );
  OR2_X1 U104 ( .A1(n99), .A2(n37), .ZN(n98) );
  AND2_X1 U105 ( .A1(n37), .A2(n99), .ZN(n97) );
  AND2_X1 U106 ( .A1(n100), .A2(n101), .ZN(n99) );
  OR2_X1 U107 ( .A1(n14), .A2(b[1]), .ZN(n101) );
  OR2_X1 U108 ( .A1(n23), .A2(a[1]), .ZN(n100) );
  AND2_X1 U109 ( .A1(n103), .A2(n104), .ZN(n102) );
  OR2_X1 U110 ( .A1(n38), .A2(d[1]), .ZN(n104) );
  OR2_X1 U111 ( .A1(n47), .A2(c[1]), .ZN(n103) );
  OR2_X1 U112 ( .A1(n105), .A2(n15), .ZN(y[0]) );
  OR2_X1 U113 ( .A1(n107), .A2(n39), .ZN(n106) );
  AND2_X1 U114 ( .A1(n39), .A2(n107), .ZN(n105) );
  AND2_X1 U115 ( .A1(n108), .A2(n109), .ZN(n107) );
  OR2_X1 U116 ( .A1(n16), .A2(b[0]), .ZN(n109) );
  OR2_X1 U117 ( .A1(n24), .A2(a[0]), .ZN(n108) );
  AND2_X1 U118 ( .A1(n111), .A2(n112), .ZN(n110) );
  OR2_X1 U119 ( .A1(n40), .A2(d[0]), .ZN(n112) );
  OR2_X1 U120 ( .A1(n48), .A2(c[0]), .ZN(n111) );
endmodule


module scale2_13 ( in, out );
  input [7:0] in;
  //input_done

  output [7:0] out;
  //output_done

  wire   in_0, \in[6] , \in[5] , \in[4] , \in[1] , \in[7] , n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20;
  //wire_done

  assign in_0 = in[0];
  assign out[7] = \in[6] ;
  assign \in[6]  = in[6];
  assign out[6] = \in[5] ;
  assign \in[5]  = in[5];
  assign out[5] = \in[4] ;
  assign \in[4]  = in[4];
  assign out[2] = \in[1] ;
  assign \in[1]  = in[1];
  assign out[0] = \in[7] ;
  assign \in[7]  = in[7];

  INV_X1 U1 ( .A(\in[7]), .ZN(n20) );
  INV_X1 U2 ( .A(in[3]), .ZN(n19) );
  INV_X1 U3 ( .A(in[2]), .ZN(n18) );
  INV_X1 U4 ( .A(in_0), .ZN(n17) );
  OR2_X1 U5 ( .A1(n16), .A2(n15), .ZN(out[4]) );
  AND2_X1 U6 ( .A1(in[3]), .A2(n20), .ZN(n15) );
  AND2_X1 U7 ( .A1(\in[7]), .A2(n19), .ZN(n16) );
  OR2_X1 U8 ( .A1(n14), .A2(n13), .ZN(out[3]) );
  AND2_X1 U9 ( .A1(in[2]), .A2(n20), .ZN(n13) );
  AND2_X1 U10 ( .A1(\in[7]), .A2(n18), .ZN(n14) );
  OR2_X1 U11 ( .A1(n12), .A2(n11), .ZN(out[1]) );
  AND2_X1 U12 ( .A1(in_0), .A2(n20), .ZN(n11) );
  AND2_X1 U13 ( .A1(\in[7]), .A2(n17), .ZN(n12) );
endmodule


module scale2_14 ( in, out );
  input [7:0] in;
  //input_done

  output [7:0] out;
  //output_done

  wire   in_0, \in[6] , \in[5] , \in[4] , \in[1] , \in[7] , n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20;
  //wire_done

  assign in_0 = in[0];
  assign out[7] = \in[6] ;
  assign \in[6]  = in[6];
  assign out[6] = \in[5] ;
  assign \in[5]  = in[5];
  assign out[5] = \in[4] ;
  assign \in[4]  = in[4];
  assign out[2] = \in[1] ;
  assign \in[1]  = in[1];
  assign out[0] = \in[7] ;
  assign \in[7]  = in[7];

  INV_X1 U1 ( .A(\in[7]), .ZN(n20) );
  INV_X1 U2 ( .A(in[3]), .ZN(n19) );
  INV_X1 U3 ( .A(in[2]), .ZN(n18) );
  INV_X1 U4 ( .A(in_0), .ZN(n17) );
  OR2_X1 U5 ( .A1(n16), .A2(n15), .ZN(out[4]) );
  AND2_X1 U6 ( .A1(in[3]), .A2(n20), .ZN(n15) );
  AND2_X1 U7 ( .A1(\in[7]), .A2(n19), .ZN(n16) );
  OR2_X1 U8 ( .A1(n14), .A2(n13), .ZN(out[3]) );
  AND2_X1 U9 ( .A1(in[2]), .A2(n20), .ZN(n13) );
  AND2_X1 U10 ( .A1(\in[7]), .A2(n18), .ZN(n14) );
  OR2_X1 U11 ( .A1(n12), .A2(n11), .ZN(out[1]) );
  AND2_X1 U12 ( .A1(in_0), .A2(n20), .ZN(n11) );
  AND2_X1 U13 ( .A1(\in[7]), .A2(n17), .ZN(n12) );
endmodule


module scale2_15 ( in, out );
  input [7:0] in;
  //input_done

  output [7:0] out;
  //output_done

  wire   in_0, \in[6] , \in[5] , \in[4] , \in[1] , \in[7] , n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20;
  //wire_done
         
  assign in_0 = in[0];
  assign out[7] = \in[6] ;
  assign \in[6]  = in[6];
  assign out[6] = \in[5] ;
  assign \in[5]  = in[5];
  assign out[5] = \in[4] ;
  assign \in[4]  = in[4];
  assign out[2] = \in[1] ;
  assign \in[1]  = in[1];
  assign out[0] = \in[7] ;
  assign \in[7]  = in[7];

  INV_X1 U1 ( .A(\in[7]), .ZN(n20) );
  INV_X1 U2 ( .A(in[3]), .ZN(n19) );
  INV_X1 U3 ( .A(in[2]), .ZN(n18) );
  INV_X1 U4 ( .A(in_0), .ZN(n17) );
  OR2_X1 U5 ( .A1(n16), .A2(n15), .ZN(out[4]) );
  AND2_X1 U6 ( .A1(in[3]), .A2(n20), .ZN(n15) );
  AND2_X1 U7 ( .A1(\in[7]), .A2(n19), .ZN(n16) );
  OR2_X1 U8 ( .A1(n14), .A2(n13), .ZN(out[3]) );
  AND2_X1 U9 ( .A1(in[2]), .A2(n20), .ZN(n13) );
  AND2_X1 U10 ( .A1(\in[7]), .A2(n18), .ZN(n14) );
  OR2_X1 U11 ( .A1(n12), .A2(n11), .ZN(out[1]) );
  AND2_X1 U12 ( .A1(in_0), .A2(n20), .ZN(n11) );
  AND2_X1 U13 ( .A1(\in[7]), .A2(n17), .ZN(n12) );
endmodule


module byteXor_14 ( a, b, y );
  input [7:0] a;
  input [7:0] b;
  //input_done

  output [7:0] y;
  //output_done

  wire   n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64;
  //wire_done

  INV_X1 U1 ( .A(n47), .ZN(n64) );
  INV_X1 U2 ( .A(a[7]), .ZN(n63) );
  INV_X1 U3 ( .A(n45), .ZN(n62) );
  INV_X1 U4 ( .A(a[6]), .ZN(n61) );
  INV_X1 U5 ( .A(n43), .ZN(n60) );
  INV_X1 U6 ( .A(a[5]), .ZN(n59) );
  INV_X1 U7 ( .A(n41), .ZN(n58) );
  INV_X1 U8 ( .A(a[4]), .ZN(n57) );
  INV_X1 U9 ( .A(n39), .ZN(n56) );
  INV_X1 U10 ( .A(a[3]), .ZN(n55) );
  INV_X1 U11 ( .A(n37), .ZN(n54) );
  INV_X1 U12 ( .A(a[2]), .ZN(n53) );
  INV_X1 U13 ( .A(n35), .ZN(n52) );
  INV_X1 U14 ( .A(a[1]), .ZN(n51) );
  INV_X1 U15 ( .A(n33), .ZN(n50) );
  INV_X1 U16 ( .A(a[0]), .ZN(n49) );
  OR2_X1 U17 ( .A1(n48), .A2(n64), .ZN(y[7]) );
  OR2_X1 U18 ( .A1(n63), .A2(b[7]), .ZN(n47) );
  AND2_X1 U19 ( .A1(b[7]), .A2(n63), .ZN(n48) );
  OR2_X1 U20 ( .A1(n46), .A2(n62), .ZN(y[6]) );
  OR2_X1 U21 ( .A1(n61), .A2(b[6]), .ZN(n45) );
  AND2_X1 U22 ( .A1(b[6]), .A2(n61), .ZN(n46) );
  OR2_X1 U23 ( .A1(n44), .A2(n60), .ZN(y[5]) );
  OR2_X1 U24 ( .A1(n59), .A2(b[5]), .ZN(n43) );
  AND2_X1 U25 ( .A1(b[5]), .A2(n59), .ZN(n44) );
  OR2_X1 U26 ( .A1(n42), .A2(n58), .ZN(y[4]) );
  OR2_X1 U27 ( .A1(n57), .A2(b[4]), .ZN(n41) );
  AND2_X1 U28 ( .A1(b[4]), .A2(n57), .ZN(n42) );
  OR2_X1 U29 ( .A1(n40), .A2(n56), .ZN(y[3]) );
  OR2_X1 U30 ( .A1(n55), .A2(b[3]), .ZN(n39) );
  AND2_X1 U31 ( .A1(b[3]), .A2(n55), .ZN(n40) );
  OR2_X1 U32 ( .A1(n38), .A2(n54), .ZN(y[2]) );
  OR2_X1 U33 ( .A1(n53), .A2(b[2]), .ZN(n37) );
  AND2_X1 U34 ( .A1(b[2]), .A2(n53), .ZN(n38) );
  OR2_X1 U35 ( .A1(n36), .A2(n52), .ZN(y[1]) );
  OR2_X1 U36 ( .A1(n51), .A2(b[1]), .ZN(n35) );
  AND2_X1 U37 ( .A1(b[1]), .A2(n51), .ZN(n36) );
  OR2_X1 U38 ( .A1(n34), .A2(n50), .ZN(y[0]) );
  OR2_X1 U39 ( .A1(n49), .A2(b[0]), .ZN(n33) );
  AND2_X1 U40 ( .A1(b[0]), .A2(n49), .ZN(n34) );
endmodule


module byteXor_15 ( a, b, y );
  input [7:0] a;
  input [7:0] b;
  //input_done

  output [7:0] y;
  //output_done

  wire   n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64;
  //wire_done

  INV_X1 U1 ( .A(n47), .ZN(n64) );
  INV_X1 U2 ( .A(a[7]), .ZN(n63) );
  INV_X1 U3 ( .A(n45), .ZN(n62) );
  INV_X1 U4 ( .A(a[6]), .ZN(n61) );
  INV_X1 U5 ( .A(n43), .ZN(n60) );
  INV_X1 U6 ( .A(a[5]), .ZN(n59) );
  INV_X1 U7 ( .A(n41), .ZN(n58) );
  INV_X1 U8 ( .A(a[4]), .ZN(n57) );
  INV_X1 U9 ( .A(n39), .ZN(n56) );
  INV_X1 U10 ( .A(a[3]), .ZN(n55) );
  INV_X1 U11 ( .A(n37), .ZN(n54) );
  INV_X1 U12 ( .A(a[2]), .ZN(n53) );
  INV_X1 U13 ( .A(n35), .ZN(n52) );
  INV_X1 U14 ( .A(a[1]), .ZN(n51) );
  INV_X1 U15 ( .A(n33), .ZN(n50) );
  INV_X1 U16 ( .A(a[0]), .ZN(n49) );
  OR2_X1 U17 ( .A1(n48), .A2(n64), .ZN(y[7]) );
  OR2_X1 U18 ( .A1(n63), .A2(b[7]), .ZN(n47) );
  AND2_X1 U19 ( .A1(b[7]), .A2(n63), .ZN(n48) );
  OR2_X1 U20 ( .A1(n46), .A2(n62), .ZN(y[6]) );
  OR2_X1 U21 ( .A1(n61), .A2(b[6]), .ZN(n45) );
  AND2_X1 U22 ( .A1(b[6]), .A2(n61), .ZN(n46) );
  OR2_X1 U23 ( .A1(n44), .A2(n60), .ZN(y[5]) );
  OR2_X1 U24 ( .A1(n59), .A2(b[5]), .ZN(n43) );
  AND2_X1 U25 ( .A1(b[5]), .A2(n59), .ZN(n44) );
  OR2_X1 U26 ( .A1(n42), .A2(n58), .ZN(y[4]) );
  OR2_X1 U27 ( .A1(n57), .A2(b[4]), .ZN(n41) );
  AND2_X1 U28 ( .A1(b[4]), .A2(n57), .ZN(n42) );
  OR2_X1 U29 ( .A1(n40), .A2(n56), .ZN(y[3]) );
  OR2_X1 U30 ( .A1(n55), .A2(b[3]), .ZN(n39) );
  AND2_X1 U31 ( .A1(b[3]), .A2(n55), .ZN(n40) );
  OR2_X1 U32 ( .A1(n38), .A2(n54), .ZN(y[2]) );
  OR2_X1 U33 ( .A1(n53), .A2(b[2]), .ZN(n37) );
  AND2_X1 U34 ( .A1(b[2]), .A2(n53), .ZN(n38) );
  OR2_X1 U35 ( .A1(n36), .A2(n52), .ZN(y[1]) );
  OR2_X1 U36 ( .A1(n51), .A2(b[1]), .ZN(n35) );
  AND2_X1 U37 ( .A1(b[1]), .A2(n51), .ZN(n36) );
  OR2_X1 U38 ( .A1(n34), .A2(n50), .ZN(y[0]) );
  OR2_X1 U39 ( .A1(n49), .A2(b[0]), .ZN(n33) );
  AND2_X1 U40 ( .A1(b[0]), .A2(n49), .ZN(n34) );
endmodule


module byteXor_16 ( a, b, y );
  input [7:0] a;
  input [7:0] b;
  //input_done

  output [7:0] y;
  //output_done

  wire   n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64;
  //wire_done

  INV_X1 U1 ( .A(n47), .ZN(n64) );
  INV_X1 U2 ( .A(a[7]), .ZN(n63) );
  INV_X1 U3 ( .A(n45), .ZN(n62) );
  INV_X1 U4 ( .A(a[6]), .ZN(n61) );
  INV_X1 U5 ( .A(n43), .ZN(n60) );
  INV_X1 U6 ( .A(a[5]), .ZN(n59) );
  INV_X1 U7 ( .A(n41), .ZN(n58) );
  INV_X1 U8 ( .A(a[4]), .ZN(n57) );
  INV_X1 U9 ( .A(n39), .ZN(n56) );
  INV_X1 U10 ( .A(a[3]), .ZN(n55) );
  INV_X1 U11 ( .A(n37), .ZN(n54) );
  INV_X1 U12 ( .A(a[2]), .ZN(n53) );
  INV_X1 U13 ( .A(n35), .ZN(n52) );
  INV_X1 U14 ( .A(a[1]), .ZN(n51) );
  INV_X1 U15 ( .A(n33), .ZN(n50) );
  INV_X1 U16 ( .A(a[0]), .ZN(n49) );
  OR2_X1 U17 ( .A1(n48), .A2(n64), .ZN(y[7]) );
  OR2_X1 U18 ( .A1(n63), .A2(b[7]), .ZN(n47) );
  AND2_X1 U19 ( .A1(b[7]), .A2(n63), .ZN(n48) );
  OR2_X1 U20 ( .A1(n46), .A2(n62), .ZN(y[6]) );
  OR2_X1 U21 ( .A1(n61), .A2(b[6]), .ZN(n45) );
  AND2_X1 U22 ( .A1(b[6]), .A2(n61), .ZN(n46) );
  OR2_X1 U23 ( .A1(n44), .A2(n60), .ZN(y[5]) );
  OR2_X1 U24 ( .A1(n59), .A2(b[5]), .ZN(n43) );
  AND2_X1 U25 ( .A1(b[5]), .A2(n59), .ZN(n44) );
  OR2_X1 U26 ( .A1(n42), .A2(n58), .ZN(y[4]) );
  OR2_X1 U27 ( .A1(n57), .A2(b[4]), .ZN(n41) );
  AND2_X1 U28 ( .A1(b[4]), .A2(n57), .ZN(n42) );
  OR2_X1 U29 ( .A1(n40), .A2(n56), .ZN(y[3]) );
  OR2_X1 U30 ( .A1(n55), .A2(b[3]), .ZN(n39) );
  AND2_X1 U31 ( .A1(b[3]), .A2(n55), .ZN(n40) );
  OR2_X1 U32 ( .A1(n38), .A2(n54), .ZN(y[2]) );
  OR2_X1 U33 ( .A1(n53), .A2(b[2]), .ZN(n37) );
  AND2_X1 U34 ( .A1(b[2]), .A2(n53), .ZN(n38) );
  OR2_X1 U35 ( .A1(n36), .A2(n52), .ZN(y[1]) );
  OR2_X1 U36 ( .A1(n51), .A2(b[1]), .ZN(n35) );
  AND2_X1 U37 ( .A1(b[1]), .A2(n51), .ZN(n36) );
  OR2_X1 U38 ( .A1(n34), .A2(n50), .ZN(y[0]) );
  OR2_X1 U39 ( .A1(n49), .A2(b[0]), .ZN(n33) );
  AND2_X1 U40 ( .A1(b[0]), .A2(n49), .ZN(n34) );
endmodule


module byteXor4_13 ( a, b, c, d, y );
  input [7:0] a;
  input [7:0] b;
  input [7:0] c;
  input [7:0] d;
  //input_done

  output [7:0] y;
  //output_done

  wire   n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224;
  //wire_done

  INV_X1 U1 ( .A(n175), .ZN(n224) );
  INV_X1 U2 ( .A(a[7]), .ZN(n223) );
  INV_X1 U3 ( .A(n167), .ZN(n222) );
  INV_X1 U4 ( .A(a[6]), .ZN(n221) );
  INV_X1 U5 ( .A(n159), .ZN(n220) );
  INV_X1 U6 ( .A(a[5]), .ZN(n219) );
  INV_X1 U7 ( .A(n151), .ZN(n218) );
  INV_X1 U8 ( .A(a[4]), .ZN(n217) );
  INV_X1 U9 ( .A(n143), .ZN(n216) );
  INV_X1 U10 ( .A(a[3]), .ZN(n215) );
  INV_X1 U11 ( .A(n135), .ZN(n214) );
  INV_X1 U12 ( .A(a[2]), .ZN(n213) );
  INV_X1 U13 ( .A(n127), .ZN(n212) );
  INV_X1 U14 ( .A(a[1]), .ZN(n211) );
  INV_X1 U15 ( .A(n119), .ZN(n210) );
  INV_X1 U16 ( .A(a[0]), .ZN(n209) );
  INV_X1 U17 ( .A(b[7]), .ZN(n208) );
  INV_X1 U18 ( .A(b[6]), .ZN(n207) );
  INV_X1 U19 ( .A(b[5]), .ZN(n206) );
  INV_X1 U20 ( .A(b[4]), .ZN(n205) );
  INV_X1 U21 ( .A(b[3]), .ZN(n204) );
  INV_X1 U22 ( .A(b[2]), .ZN(n203) );
  INV_X1 U23 ( .A(b[1]), .ZN(n202) );
  INV_X1 U24 ( .A(b[0]), .ZN(n201) );
  INV_X1 U25 ( .A(n171), .ZN(n200) );
  INV_X1 U26 ( .A(c[7]), .ZN(n199) );
  INV_X1 U27 ( .A(n163), .ZN(n198) );
  INV_X1 U28 ( .A(c[6]), .ZN(n197) );
  INV_X1 U29 ( .A(n155), .ZN(n196) );
  INV_X1 U30 ( .A(c[5]), .ZN(n195) );
  INV_X1 U31 ( .A(n147), .ZN(n194) );
  INV_X1 U32 ( .A(c[4]), .ZN(n193) );
  INV_X1 U33 ( .A(n139), .ZN(n192) );
  INV_X1 U34 ( .A(c[3]), .ZN(n191) );
  INV_X1 U35 ( .A(n131), .ZN(n190) );
  INV_X1 U36 ( .A(c[2]), .ZN(n189) );
  INV_X1 U37 ( .A(n123), .ZN(n188) );
  INV_X1 U38 ( .A(c[1]), .ZN(n187) );
  INV_X1 U39 ( .A(n115), .ZN(n186) );
  INV_X1 U40 ( .A(c[0]), .ZN(n185) );
  INV_X1 U41 ( .A(d[7]), .ZN(n184) );
  INV_X1 U42 ( .A(d[6]), .ZN(n183) );
  INV_X1 U43 ( .A(d[5]), .ZN(n182) );
  INV_X1 U44 ( .A(d[4]), .ZN(n181) );
  INV_X1 U45 ( .A(d[3]), .ZN(n180) );
  INV_X1 U46 ( .A(d[2]), .ZN(n179) );
  INV_X1 U47 ( .A(d[1]), .ZN(n178) );
  INV_X1 U48 ( .A(d[0]), .ZN(n177) );
  OR2_X1 U49 ( .A1(n176), .A2(n224), .ZN(y[7]) );
  OR2_X1 U50 ( .A1(n174), .A2(n200), .ZN(n175) );
  AND2_X1 U51 ( .A1(n200), .A2(n174), .ZN(n176) );
  AND2_X1 U52 ( .A1(n173), .A2(n172), .ZN(n174) );
  OR2_X1 U53 ( .A1(n223), .A2(b[7]), .ZN(n172) );
  OR2_X1 U54 ( .A1(n208), .A2(a[7]), .ZN(n173) );
  AND2_X1 U55 ( .A1(n170), .A2(n169), .ZN(n171) );
  OR2_X1 U56 ( .A1(n199), .A2(d[7]), .ZN(n169) );
  OR2_X1 U57 ( .A1(n184), .A2(c[7]), .ZN(n170) );
  OR2_X1 U58 ( .A1(n168), .A2(n222), .ZN(y[6]) );
  OR2_X1 U59 ( .A1(n166), .A2(n198), .ZN(n167) );
  AND2_X1 U60 ( .A1(n198), .A2(n166), .ZN(n168) );
  AND2_X1 U61 ( .A1(n165), .A2(n164), .ZN(n166) );
  OR2_X1 U62 ( .A1(n221), .A2(b[6]), .ZN(n164) );
  OR2_X1 U63 ( .A1(n207), .A2(a[6]), .ZN(n165) );
  AND2_X1 U64 ( .A1(n162), .A2(n161), .ZN(n163) );
  OR2_X1 U65 ( .A1(n197), .A2(d[6]), .ZN(n161) );
  OR2_X1 U66 ( .A1(n183), .A2(c[6]), .ZN(n162) );
  OR2_X1 U67 ( .A1(n160), .A2(n220), .ZN(y[5]) );
  OR2_X1 U68 ( .A1(n158), .A2(n196), .ZN(n159) );
  AND2_X1 U69 ( .A1(n196), .A2(n158), .ZN(n160) );
  AND2_X1 U70 ( .A1(n157), .A2(n156), .ZN(n158) );
  OR2_X1 U71 ( .A1(n219), .A2(b[5]), .ZN(n156) );
  OR2_X1 U72 ( .A1(n206), .A2(a[5]), .ZN(n157) );
  AND2_X1 U73 ( .A1(n154), .A2(n153), .ZN(n155) );
  OR2_X1 U74 ( .A1(n195), .A2(d[5]), .ZN(n153) );
  OR2_X1 U75 ( .A1(n182), .A2(c[5]), .ZN(n154) );
  OR2_X1 U76 ( .A1(n152), .A2(n218), .ZN(y[4]) );
  OR2_X1 U77 ( .A1(n150), .A2(n194), .ZN(n151) );
  AND2_X1 U78 ( .A1(n194), .A2(n150), .ZN(n152) );
  AND2_X1 U79 ( .A1(n149), .A2(n148), .ZN(n150) );
  OR2_X1 U80 ( .A1(n217), .A2(b[4]), .ZN(n148) );
  OR2_X1 U81 ( .A1(n205), .A2(a[4]), .ZN(n149) );
  AND2_X1 U82 ( .A1(n146), .A2(n145), .ZN(n147) );
  OR2_X1 U83 ( .A1(n193), .A2(d[4]), .ZN(n145) );
  OR2_X1 U84 ( .A1(n181), .A2(c[4]), .ZN(n146) );
  OR2_X1 U85 ( .A1(n144), .A2(n216), .ZN(y[3]) );
  OR2_X1 U86 ( .A1(n142), .A2(n192), .ZN(n143) );
  AND2_X1 U87 ( .A1(n192), .A2(n142), .ZN(n144) );
  AND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(n142) );
  OR2_X1 U89 ( .A1(n215), .A2(b[3]), .ZN(n140) );
  OR2_X1 U90 ( .A1(n204), .A2(a[3]), .ZN(n141) );
  AND2_X1 U91 ( .A1(n138), .A2(n137), .ZN(n139) );
  OR2_X1 U92 ( .A1(n191), .A2(d[3]), .ZN(n137) );
  OR2_X1 U93 ( .A1(n180), .A2(c[3]), .ZN(n138) );
  OR2_X1 U94 ( .A1(n136), .A2(n214), .ZN(y[2]) );
  OR2_X1 U95 ( .A1(n134), .A2(n190), .ZN(n135) );
  AND2_X1 U96 ( .A1(n190), .A2(n134), .ZN(n136) );
  AND2_X1 U97 ( .A1(n133), .A2(n132), .ZN(n134) );
  OR2_X1 U98 ( .A1(n213), .A2(b[2]), .ZN(n132) );
  OR2_X1 U99 ( .A1(n203), .A2(a[2]), .ZN(n133) );
  AND2_X1 U100 ( .A1(n130), .A2(n129), .ZN(n131) );
  OR2_X1 U101 ( .A1(n189), .A2(d[2]), .ZN(n129) );
  OR2_X1 U102 ( .A1(n179), .A2(c[2]), .ZN(n130) );
  OR2_X1 U103 ( .A1(n128), .A2(n212), .ZN(y[1]) );
  OR2_X1 U104 ( .A1(n126), .A2(n188), .ZN(n127) );
  AND2_X1 U105 ( .A1(n188), .A2(n126), .ZN(n128) );
  AND2_X1 U106 ( .A1(n125), .A2(n124), .ZN(n126) );
  OR2_X1 U107 ( .A1(n211), .A2(b[1]), .ZN(n124) );
  OR2_X1 U108 ( .A1(n202), .A2(a[1]), .ZN(n125) );
  AND2_X1 U109 ( .A1(n122), .A2(n121), .ZN(n123) );
  OR2_X1 U110 ( .A1(n187), .A2(d[1]), .ZN(n121) );
  OR2_X1 U111 ( .A1(n178), .A2(c[1]), .ZN(n122) );
  OR2_X1 U112 ( .A1(n120), .A2(n210), .ZN(y[0]) );
  OR2_X1 U113 ( .A1(n118), .A2(n186), .ZN(n119) );
  AND2_X1 U114 ( .A1(n186), .A2(n118), .ZN(n120) );
  AND2_X1 U115 ( .A1(n117), .A2(n116), .ZN(n118) );
  OR2_X1 U116 ( .A1(n209), .A2(b[0]), .ZN(n116) );
  OR2_X1 U117 ( .A1(n201), .A2(a[0]), .ZN(n117) );
  AND2_X1 U118 ( .A1(n114), .A2(n113), .ZN(n115) );
  OR2_X1 U119 ( .A1(n185), .A2(d[0]), .ZN(n113) );
  OR2_X1 U120 ( .A1(n177), .A2(c[0]), .ZN(n114) );
endmodule


module byteXor4_14 ( a, b, c, d, y );
  input [7:0] a;
  input [7:0] b;
  input [7:0] c;
  input [7:0] d;
  //input_done

  output [7:0] y;
  //output_done

  wire   n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224;
  //wire_done

  INV_X1 U1 ( .A(n175), .ZN(n224) );
  INV_X1 U2 ( .A(a[7]), .ZN(n223) );
  INV_X1 U3 ( .A(n167), .ZN(n222) );
  INV_X1 U4 ( .A(a[6]), .ZN(n221) );
  INV_X1 U5 ( .A(n159), .ZN(n220) );
  INV_X1 U6 ( .A(a[5]), .ZN(n219) );
  INV_X1 U7 ( .A(n151), .ZN(n218) );
  INV_X1 U8 ( .A(a[4]), .ZN(n217) );
  INV_X1 U9 ( .A(n143), .ZN(n216) );
  INV_X1 U10 ( .A(a[3]), .ZN(n215) );
  INV_X1 U11 ( .A(n135), .ZN(n214) );
  INV_X1 U12 ( .A(a[2]), .ZN(n213) );
  INV_X1 U13 ( .A(n127), .ZN(n212) );
  INV_X1 U14 ( .A(a[1]), .ZN(n211) );
  INV_X1 U15 ( .A(n119), .ZN(n210) );
  INV_X1 U16 ( .A(a[0]), .ZN(n209) );
  INV_X1 U17 ( .A(b[7]), .ZN(n208) );
  INV_X1 U18 ( .A(b[6]), .ZN(n207) );
  INV_X1 U19 ( .A(b[5]), .ZN(n206) );
  INV_X1 U20 ( .A(b[4]), .ZN(n205) );
  INV_X1 U21 ( .A(b[3]), .ZN(n204) );
  INV_X1 U22 ( .A(b[2]), .ZN(n203) );
  INV_X1 U23 ( .A(b[1]), .ZN(n202) );
  INV_X1 U24 ( .A(b[0]), .ZN(n201) );
  INV_X1 U25 ( .A(n171), .ZN(n200) );
  INV_X1 U26 ( .A(c[7]), .ZN(n199) );
  INV_X1 U27 ( .A(n163), .ZN(n198) );
  INV_X1 U28 ( .A(c[6]), .ZN(n197) );
  INV_X1 U29 ( .A(n155), .ZN(n196) );
  INV_X1 U30 ( .A(c[5]), .ZN(n195) );
  INV_X1 U31 ( .A(n147), .ZN(n194) );
  INV_X1 U32 ( .A(c[4]), .ZN(n193) );
  INV_X1 U33 ( .A(n139), .ZN(n192) );
  INV_X1 U34 ( .A(c[3]), .ZN(n191) );
  INV_X1 U35 ( .A(n131), .ZN(n190) );
  INV_X1 U36 ( .A(c[2]), .ZN(n189) );
  INV_X1 U37 ( .A(n123), .ZN(n188) );
  INV_X1 U38 ( .A(c[1]), .ZN(n187) );
  INV_X1 U39 ( .A(n115), .ZN(n186) );
  INV_X1 U40 ( .A(c[0]), .ZN(n185) );
  INV_X1 U41 ( .A(d[7]), .ZN(n184) );
  INV_X1 U42 ( .A(d[6]), .ZN(n183) );
  INV_X1 U43 ( .A(d[5]), .ZN(n182) );
  INV_X1 U44 ( .A(d[4]), .ZN(n181) );
  INV_X1 U45 ( .A(d[3]), .ZN(n180) );
  INV_X1 U46 ( .A(d[2]), .ZN(n179) );
  INV_X1 U47 ( .A(d[1]), .ZN(n178) );
  INV_X1 U48 ( .A(d[0]), .ZN(n177) );
  OR2_X1 U49 ( .A1(n176), .A2(n224), .ZN(y[7]) );
  OR2_X1 U50 ( .A1(n174), .A2(n200), .ZN(n175) );
  AND2_X1 U51 ( .A1(n200), .A2(n174), .ZN(n176) );
  AND2_X1 U52 ( .A1(n173), .A2(n172), .ZN(n174) );
  OR2_X1 U53 ( .A1(n223), .A2(b[7]), .ZN(n172) );
  OR2_X1 U54 ( .A1(n208), .A2(a[7]), .ZN(n173) );
  AND2_X1 U55 ( .A1(n170), .A2(n169), .ZN(n171) );
  OR2_X1 U56 ( .A1(n199), .A2(d[7]), .ZN(n169) );
  OR2_X1 U57 ( .A1(n184), .A2(c[7]), .ZN(n170) );
  OR2_X1 U58 ( .A1(n168), .A2(n222), .ZN(y[6]) );
  OR2_X1 U59 ( .A1(n166), .A2(n198), .ZN(n167) );
  AND2_X1 U60 ( .A1(n198), .A2(n166), .ZN(n168) );
  AND2_X1 U61 ( .A1(n165), .A2(n164), .ZN(n166) );
  OR2_X1 U62 ( .A1(n221), .A2(b[6]), .ZN(n164) );
  OR2_X1 U63 ( .A1(n207), .A2(a[6]), .ZN(n165) );
  AND2_X1 U64 ( .A1(n162), .A2(n161), .ZN(n163) );
  OR2_X1 U65 ( .A1(n197), .A2(d[6]), .ZN(n161) );
  OR2_X1 U66 ( .A1(n183), .A2(c[6]), .ZN(n162) );
  OR2_X1 U67 ( .A1(n160), .A2(n220), .ZN(y[5]) );
  OR2_X1 U68 ( .A1(n158), .A2(n196), .ZN(n159) );
  AND2_X1 U69 ( .A1(n196), .A2(n158), .ZN(n160) );
  AND2_X1 U70 ( .A1(n157), .A2(n156), .ZN(n158) );
  OR2_X1 U71 ( .A1(n219), .A2(b[5]), .ZN(n156) );
  OR2_X1 U72 ( .A1(n206), .A2(a[5]), .ZN(n157) );
  AND2_X1 U73 ( .A1(n154), .A2(n153), .ZN(n155) );
  OR2_X1 U74 ( .A1(n195), .A2(d[5]), .ZN(n153) );
  OR2_X1 U75 ( .A1(n182), .A2(c[5]), .ZN(n154) );
  OR2_X1 U76 ( .A1(n152), .A2(n218), .ZN(y[4]) );
  OR2_X1 U77 ( .A1(n150), .A2(n194), .ZN(n151) );
  AND2_X1 U78 ( .A1(n194), .A2(n150), .ZN(n152) );
  AND2_X1 U79 ( .A1(n149), .A2(n148), .ZN(n150) );
  OR2_X1 U80 ( .A1(n217), .A2(b[4]), .ZN(n148) );
  OR2_X1 U81 ( .A1(n205), .A2(a[4]), .ZN(n149) );
  AND2_X1 U82 ( .A1(n146), .A2(n145), .ZN(n147) );
  OR2_X1 U83 ( .A1(n193), .A2(d[4]), .ZN(n145) );
  OR2_X1 U84 ( .A1(n181), .A2(c[4]), .ZN(n146) );
  OR2_X1 U85 ( .A1(n144), .A2(n216), .ZN(y[3]) );
  OR2_X1 U86 ( .A1(n142), .A2(n192), .ZN(n143) );
  AND2_X1 U87 ( .A1(n192), .A2(n142), .ZN(n144) );
  AND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(n142) );
  OR2_X1 U89 ( .A1(n215), .A2(b[3]), .ZN(n140) );
  OR2_X1 U90 ( .A1(n204), .A2(a[3]), .ZN(n141) );
  AND2_X1 U91 ( .A1(n138), .A2(n137), .ZN(n139) );
  OR2_X1 U92 ( .A1(n191), .A2(d[3]), .ZN(n137) );
  OR2_X1 U93 ( .A1(n180), .A2(c[3]), .ZN(n138) );
  OR2_X1 U94 ( .A1(n136), .A2(n214), .ZN(y[2]) );
  OR2_X1 U95 ( .A1(n134), .A2(n190), .ZN(n135) );
  AND2_X1 U96 ( .A1(n190), .A2(n134), .ZN(n136) );
  AND2_X1 U97 ( .A1(n133), .A2(n132), .ZN(n134) );
  OR2_X1 U98 ( .A1(n213), .A2(b[2]), .ZN(n132) );
  OR2_X1 U99 ( .A1(n203), .A2(a[2]), .ZN(n133) );
  AND2_X1 U100 ( .A1(n130), .A2(n129), .ZN(n131) );
  OR2_X1 U101 ( .A1(n189), .A2(d[2]), .ZN(n129) );
  OR2_X1 U102 ( .A1(n179), .A2(c[2]), .ZN(n130) );
  OR2_X1 U103 ( .A1(n128), .A2(n212), .ZN(y[1]) );
  OR2_X1 U104 ( .A1(n126), .A2(n188), .ZN(n127) );
  AND2_X1 U105 ( .A1(n188), .A2(n126), .ZN(n128) );
  AND2_X1 U106 ( .A1(n125), .A2(n124), .ZN(n126) );
  OR2_X1 U107 ( .A1(n211), .A2(b[1]), .ZN(n124) );
  OR2_X1 U108 ( .A1(n202), .A2(a[1]), .ZN(n125) );
  AND2_X1 U109 ( .A1(n122), .A2(n121), .ZN(n123) );
  OR2_X1 U110 ( .A1(n187), .A2(d[1]), .ZN(n121) );
  OR2_X1 U111 ( .A1(n178), .A2(c[1]), .ZN(n122) );
  OR2_X1 U112 ( .A1(n120), .A2(n210), .ZN(y[0]) );
  OR2_X1 U113 ( .A1(n118), .A2(n186), .ZN(n119) );
  AND2_X1 U114 ( .A1(n186), .A2(n118), .ZN(n120) );
  AND2_X1 U115 ( .A1(n117), .A2(n116), .ZN(n118) );
  OR2_X1 U116 ( .A1(n209), .A2(b[0]), .ZN(n116) );
  OR2_X1 U117 ( .A1(n201), .A2(a[0]), .ZN(n117) );
  AND2_X1 U118 ( .A1(n114), .A2(n113), .ZN(n115) );
  OR2_X1 U119 ( .A1(n185), .A2(d[0]), .ZN(n113) );
  OR2_X1 U120 ( .A1(n177), .A2(c[0]), .ZN(n114) );
endmodule


module byteXor4_15 ( a, b, c, d, y );
  input [7:0] a;
  input [7:0] b;
  input [7:0] c;
  input [7:0] d;
  //input_done

  output [7:0] y;
  //output_done

  wire   n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224;
  //wire_done

  INV_X1 U1 ( .A(n175), .ZN(n224) );
  INV_X1 U2 ( .A(a[7]), .ZN(n223) );
  INV_X1 U3 ( .A(n167), .ZN(n222) );
  INV_X1 U4 ( .A(a[6]), .ZN(n221) );
  INV_X1 U5 ( .A(n159), .ZN(n220) );
  INV_X1 U6 ( .A(a[5]), .ZN(n219) );
  INV_X1 U7 ( .A(n151), .ZN(n218) );
  INV_X1 U8 ( .A(a[4]), .ZN(n217) );
  INV_X1 U9 ( .A(n143), .ZN(n216) );
  INV_X1 U10 ( .A(a[3]), .ZN(n215) );
  INV_X1 U11 ( .A(n135), .ZN(n214) );
  INV_X1 U12 ( .A(a[2]), .ZN(n213) );
  INV_X1 U13 ( .A(n127), .ZN(n212) );
  INV_X1 U14 ( .A(a[1]), .ZN(n211) );
  INV_X1 U15 ( .A(n119), .ZN(n210) );
  INV_X1 U16 ( .A(a[0]), .ZN(n209) );
  INV_X1 U17 ( .A(b[7]), .ZN(n208) );
  INV_X1 U18 ( .A(b[6]), .ZN(n207) );
  INV_X1 U19 ( .A(b[5]), .ZN(n206) );
  INV_X1 U20 ( .A(b[4]), .ZN(n205) );
  INV_X1 U21 ( .A(b[3]), .ZN(n204) );
  INV_X1 U22 ( .A(b[2]), .ZN(n203) );
  INV_X1 U23 ( .A(b[1]), .ZN(n202) );
  INV_X1 U24 ( .A(b[0]), .ZN(n201) );
  INV_X1 U25 ( .A(n171), .ZN(n200) );
  INV_X1 U26 ( .A(c[7]), .ZN(n199) );
  INV_X1 U27 ( .A(n163), .ZN(n198) );
  INV_X1 U28 ( .A(c[6]), .ZN(n197) );
  INV_X1 U29 ( .A(n155), .ZN(n196) );
  INV_X1 U30 ( .A(c[5]), .ZN(n195) );
  INV_X1 U31 ( .A(n147), .ZN(n194) );
  INV_X1 U32 ( .A(c[4]), .ZN(n193) );
  INV_X1 U33 ( .A(n139), .ZN(n192) );
  INV_X1 U34 ( .A(c[3]), .ZN(n191) );
  INV_X1 U35 ( .A(n131), .ZN(n190) );
  INV_X1 U36 ( .A(c[2]), .ZN(n189) );
  INV_X1 U37 ( .A(n123), .ZN(n188) );
  INV_X1 U38 ( .A(c[1]), .ZN(n187) );
  INV_X1 U39 ( .A(n115), .ZN(n186) );
  INV_X1 U40 ( .A(c[0]), .ZN(n185) );
  INV_X1 U41 ( .A(d[7]), .ZN(n184) );
  INV_X1 U42 ( .A(d[6]), .ZN(n183) );
  INV_X1 U43 ( .A(d[5]), .ZN(n182) );
  INV_X1 U44 ( .A(d[4]), .ZN(n181) );
  INV_X1 U45 ( .A(d[3]), .ZN(n180) );
  INV_X1 U46 ( .A(d[2]), .ZN(n179) );
  INV_X1 U47 ( .A(d[1]), .ZN(n178) );
  INV_X1 U48 ( .A(d[0]), .ZN(n177) );
  OR2_X1 U49 ( .A1(n176), .A2(n224), .ZN(y[7]) );
  OR2_X1 U50 ( .A1(n174), .A2(n200), .ZN(n175) );
  AND2_X1 U51 ( .A1(n200), .A2(n174), .ZN(n176) );
  AND2_X1 U52 ( .A1(n173), .A2(n172), .ZN(n174) );
  OR2_X1 U53 ( .A1(n223), .A2(b[7]), .ZN(n172) );
  OR2_X1 U54 ( .A1(n208), .A2(a[7]), .ZN(n173) );
  AND2_X1 U55 ( .A1(n170), .A2(n169), .ZN(n171) );
  OR2_X1 U56 ( .A1(n199), .A2(d[7]), .ZN(n169) );
  OR2_X1 U57 ( .A1(n184), .A2(c[7]), .ZN(n170) );
  OR2_X1 U58 ( .A1(n168), .A2(n222), .ZN(y[6]) );
  OR2_X1 U59 ( .A1(n166), .A2(n198), .ZN(n167) );
  AND2_X1 U60 ( .A1(n198), .A2(n166), .ZN(n168) );
  AND2_X1 U61 ( .A1(n165), .A2(n164), .ZN(n166) );
  OR2_X1 U62 ( .A1(n221), .A2(b[6]), .ZN(n164) );
  OR2_X1 U63 ( .A1(n207), .A2(a[6]), .ZN(n165) );
  AND2_X1 U64 ( .A1(n162), .A2(n161), .ZN(n163) );
  OR2_X1 U65 ( .A1(n197), .A2(d[6]), .ZN(n161) );
  OR2_X1 U66 ( .A1(n183), .A2(c[6]), .ZN(n162) );
  OR2_X1 U67 ( .A1(n160), .A2(n220), .ZN(y[5]) );
  OR2_X1 U68 ( .A1(n158), .A2(n196), .ZN(n159) );
  AND2_X1 U69 ( .A1(n196), .A2(n158), .ZN(n160) );
  AND2_X1 U70 ( .A1(n157), .A2(n156), .ZN(n158) );
  OR2_X1 U71 ( .A1(n219), .A2(b[5]), .ZN(n156) );
  OR2_X1 U72 ( .A1(n206), .A2(a[5]), .ZN(n157) );
  AND2_X1 U73 ( .A1(n154), .A2(n153), .ZN(n155) );
  OR2_X1 U74 ( .A1(n195), .A2(d[5]), .ZN(n153) );
  OR2_X1 U75 ( .A1(n182), .A2(c[5]), .ZN(n154) );
  OR2_X1 U76 ( .A1(n152), .A2(n218), .ZN(y[4]) );
  OR2_X1 U77 ( .A1(n150), .A2(n194), .ZN(n151) );
  AND2_X1 U78 ( .A1(n194), .A2(n150), .ZN(n152) );
  AND2_X1 U79 ( .A1(n149), .A2(n148), .ZN(n150) );
  OR2_X1 U80 ( .A1(n217), .A2(b[4]), .ZN(n148) );
  OR2_X1 U81 ( .A1(n205), .A2(a[4]), .ZN(n149) );
  AND2_X1 U82 ( .A1(n146), .A2(n145), .ZN(n147) );
  OR2_X1 U83 ( .A1(n193), .A2(d[4]), .ZN(n145) );
  OR2_X1 U84 ( .A1(n181), .A2(c[4]), .ZN(n146) );
  OR2_X1 U85 ( .A1(n144), .A2(n216), .ZN(y[3]) );
  OR2_X1 U86 ( .A1(n142), .A2(n192), .ZN(n143) );
  AND2_X1 U87 ( .A1(n192), .A2(n142), .ZN(n144) );
  AND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(n142) );
  OR2_X1 U89 ( .A1(n215), .A2(b[3]), .ZN(n140) );
  OR2_X1 U90 ( .A1(n204), .A2(a[3]), .ZN(n141) );
  AND2_X1 U91 ( .A1(n138), .A2(n137), .ZN(n139) );
  OR2_X1 U92 ( .A1(n191), .A2(d[3]), .ZN(n137) );
  OR2_X1 U93 ( .A1(n180), .A2(c[3]), .ZN(n138) );
  OR2_X1 U94 ( .A1(n136), .A2(n214), .ZN(y[2]) );
  OR2_X1 U95 ( .A1(n134), .A2(n190), .ZN(n135) );
  AND2_X1 U96 ( .A1(n190), .A2(n134), .ZN(n136) );
  AND2_X1 U97 ( .A1(n133), .A2(n132), .ZN(n134) );
  OR2_X1 U98 ( .A1(n213), .A2(b[2]), .ZN(n132) );
  OR2_X1 U99 ( .A1(n203), .A2(a[2]), .ZN(n133) );
  AND2_X1 U100 ( .A1(n130), .A2(n129), .ZN(n131) );
  OR2_X1 U101 ( .A1(n189), .A2(d[2]), .ZN(n129) );
  OR2_X1 U102 ( .A1(n179), .A2(c[2]), .ZN(n130) );
  OR2_X1 U103 ( .A1(n128), .A2(n212), .ZN(y[1]) );
  OR2_X1 U104 ( .A1(n126), .A2(n188), .ZN(n127) );
  AND2_X1 U105 ( .A1(n188), .A2(n126), .ZN(n128) );
  AND2_X1 U106 ( .A1(n125), .A2(n124), .ZN(n126) );
  OR2_X1 U107 ( .A1(n211), .A2(b[1]), .ZN(n124) );
  OR2_X1 U108 ( .A1(n202), .A2(a[1]), .ZN(n125) );
  AND2_X1 U109 ( .A1(n122), .A2(n121), .ZN(n123) );
  OR2_X1 U110 ( .A1(n187), .A2(d[1]), .ZN(n121) );
  OR2_X1 U111 ( .A1(n178), .A2(c[1]), .ZN(n122) );
  OR2_X1 U112 ( .A1(n120), .A2(n210), .ZN(y[0]) );
  OR2_X1 U113 ( .A1(n118), .A2(n186), .ZN(n119) );
  AND2_X1 U114 ( .A1(n186), .A2(n118), .ZN(n120) );
  AND2_X1 U115 ( .A1(n117), .A2(n116), .ZN(n118) );
  OR2_X1 U116 ( .A1(n209), .A2(b[0]), .ZN(n116) );
  OR2_X1 U117 ( .A1(n201), .A2(a[0]), .ZN(n117) );
  AND2_X1 U118 ( .A1(n114), .A2(n113), .ZN(n115) );
  OR2_X1 U119 ( .A1(n185), .A2(d[0]), .ZN(n113) );
  OR2_X1 U120 ( .A1(n177), .A2(c[0]), .ZN(n114) );
endmodule


module mixCol_0 ( in, out );
  input [31:0] in;
  //input_done

  output [31:0] out;
  //output_done

  wire   [7:0] b0_s2;
  wire   [7:0] b1_s2;
  wire   [7:0] b2_s2;
  wire   [7:0] b3_s2;
  wire   [7:0] b0_s3;
  wire   [7:0] b1_s3;
  wire   [7:0] b2_s3;
  wire   [7:0] b3_s3;
  //wire_done

  scale2_0 b0_scale2 ( .in(in[31:24]), .out(b0_s2) );
  scale2_15 b1_scale2 ( .in(in[23:16]), .out(b1_s2) );
  scale2_14 b2_scale2 ( .in(in[15:8]), .out(b2_s2) );
  scale2_13 b3_scale2 ( .in(in[7:0]), .out(b3_s2) );
  byteXor_0 b0_scale3 ( .a(in[31:24]), .b(b0_s2), .y(b0_s3) );
  byteXor_16 b1_scale3 ( .a(in[23:16]), .b(b1_s2), .y(b1_s3) );
  byteXor_15 b2_scale3 ( .a(in[15:8]), .b(b2_s2), .y(b2_s3) );
  byteXor_14 b3_scale3 ( .a(in[7:0]), .b(b3_s2), .y(b3_s3) );
  byteXor4_0 out0 ( .a(b0_s2), .b(b1_s3), .c(in[15:8]), .d(in[7:0]), .y(
        out[31:24]) );
  byteXor4_15 out1 ( .a(in[31:24]), .b(b1_s2), .c(b2_s3), .d(in[7:0]), .y(
        out[23:16]) );
  byteXor4_14 out2 ( .a(in[31:24]), .b(in[23:16]), .c(b2_s2), .d(b3_s3), .y(
        out[15:8]) );
  byteXor4_13 out3 ( .a(b0_s3), .b(in[23:16]), .c(in[15:8]), .d(b3_s2), .y(
        out[7:0]) );
endmodule


module CD2_1 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_2 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done

  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_3 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_4 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD4_1 ( a, b, y );
  input [3:0] a;
  input [3:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  //input_done

  output [15:0] y;
  reg [15:0] ybar;
  //output_done


  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
endmodule


module CD4_2 ( a, b, y );
  input [3:0] a;
  input [3:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  //input_done

  output [15:0] y;
  reg [15:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]);
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]);
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]);
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]);
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]);
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]);
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]);
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]);
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]);
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]);
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]);
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]);
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]);
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]);
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]);
endmodule




module CD4_2 ( a, b, y );
  input [3:0] a;
  input [3:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  //input_done

  output [15:0] y;
  reg [15:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]);
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]);
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]);
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]);
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]);
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]);
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]);
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]);
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]);
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]);
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]);
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]);
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]);
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]);
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]);
endmodule




module CD16_1 ( a, b, y );
  input [15:0] a;
  input [15:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign abar[8] = ~a[8];
  assign abar[9] = ~a[9];
  assign abar[10] = ~a[10];
  assign abar[11] = ~a[11];
  assign abar[12] = ~a[12];
  assign abar[13] = ~a[13];
  assign abar[14] = ~a[14];
  assign abar[15] = ~a[15];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign bbar[8] = ~b[8];
  assign bbar[9] = ~b[9];
  assign bbar[10] = ~b[10];
  assign bbar[11] = ~b[11];
  assign bbar[12] = ~b[12];
  assign bbar[13] = ~b[13];
  assign bbar[14] = ~b[14];
  assign bbar[15] = ~b[15];
  //input_done

  output [255:0] y;
  reg [255:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[9]), .A2(a[0]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[9]), .A2(abar[0]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[3]), .A2(a[6]), .ZN(y[99]) );
  OR2_X1 U2bar ( .A1(bbar[3]), .A2(abar[6]), .ZN(ybar[99]);
  AND2_X1 U3 ( .A1(b[2]), .A2(a[6]), .ZN(y[98]) );
  OR2_X1 U3bar ( .A1(bbar[2]), .A2(abar[6]), .ZN(ybar[98]);
  AND2_X1 U4 ( .A1(b[1]), .A2(a[6]), .ZN(y[97]) );
  OR2_X1 U4bar ( .A1(bbar[1]), .A2(abar[6]), .ZN(ybar[97]);
  AND2_X1 U5 ( .A1(b[0]), .A2(a[6]), .ZN(y[96]) );
  OR2_X1 U5bar ( .A1(bbar[0]), .A2(abar[6]), .ZN(ybar[96]);
  AND2_X1 U6 ( .A1(b[15]), .A2(a[5]), .ZN(y[95]) );
  OR2_X1 U6bar ( .A1(bbar[15]), .A2(abar[5]), .ZN(ybar[95]);
  AND2_X1 U7 ( .A1(b[14]), .A2(a[5]), .ZN(y[94]) );
  OR2_X1 U7bar ( .A1(bbar[14]), .A2(abar[5]), .ZN(ybar[94]);
  AND2_X1 U8 ( .A1(b[13]), .A2(a[5]), .ZN(y[93]) );
  OR2_X1 U8bar ( .A1(bbar[13]), .A2(abar[5]), .ZN(ybar[93]);
  AND2_X1 U9 ( .A1(b[12]), .A2(a[5]), .ZN(y[92]) );
  OR2_X1 U9bar ( .A1(bbar[12]), .A2(abar[5]), .ZN(ybar[92]);
  AND2_X1 U10 ( .A1(b[11]), .A2(a[5]), .ZN(y[91]) );
  OR2_X1 U10bar ( .A1(bbar[11]), .A2(abar[5]), .ZN(ybar[91]);
  AND2_X1 U11 ( .A1(b[10]), .A2(a[5]), .ZN(y[90]) );
  OR2_X1 U11bar ( .A1(bbar[10]), .A2(abar[5]), .ZN(ybar[90]);
  AND2_X1 U12 ( .A1(b[8]), .A2(a[0]), .ZN(y[8]) );
  OR2_X1 U12bar ( .A1(bbar[8]), .A2(abar[0]), .ZN(ybar[8]);
  AND2_X1 U13 ( .A1(a[5]), .A2(b[9]), .ZN(y[89]) );
  OR2_X1 U13bar ( .A1(abar[5]), .A2(bbar[9]), .ZN(ybar[89]);
  AND2_X1 U14 ( .A1(b[8]), .A2(a[5]), .ZN(y[88]) );
  OR2_X1 U14bar ( .A1(bbar[8]), .A2(abar[5]), .ZN(ybar[88]);
  AND2_X1 U15 ( .A1(b[7]), .A2(a[5]), .ZN(y[87]) );
  OR2_X1 U15bar ( .A1(bbar[7]), .A2(abar[5]), .ZN(ybar[87]);
  AND2_X1 U16 ( .A1(b[6]), .A2(a[5]), .ZN(y[86]) );
  OR2_X1 U16bar ( .A1(bbar[6]), .A2(abar[5]), .ZN(ybar[86]);
  AND2_X1 U17 ( .A1(b[5]), .A2(a[5]), .ZN(y[85]) );
  OR2_X1 U17bar ( .A1(bbar[5]), .A2(abar[5]), .ZN(ybar[85]);
  AND2_X1 U18 ( .A1(b[4]), .A2(a[5]), .ZN(y[84]) );
  OR2_X1 U18bar ( .A1(bbar[4]), .A2(abar[5]), .ZN(ybar[84]);
  AND2_X1 U19 ( .A1(a[5]), .A2(b[3]), .ZN(y[83]) );
  OR2_X1 U19bar ( .A1(abar[5]), .A2(bbar[3]), .ZN(ybar[83]);
  AND2_X1 U20 ( .A1(a[5]), .A2(b[2]), .ZN(y[82]) );
  OR2_X1 U20bar ( .A1(abar[5]), .A2(bbar[2]), .ZN(ybar[82]);
  AND2_X1 U21 ( .A1(a[5]), .A2(b[1]), .ZN(y[81]) );
  OR2_X1 U21bar ( .A1(abar[5]), .A2(bbar[1]), .ZN(ybar[81]);
  AND2_X1 U22 ( .A1(a[5]), .A2(b[0]), .ZN(y[80]) );
  OR2_X1 U22bar ( .A1(abar[5]), .A2(bbar[0]), .ZN(ybar[80]);
  AND2_X1 U23 ( .A1(b[7]), .A2(a[0]), .ZN(y[7]) );
  OR2_X1 U23bar ( .A1(bbar[7]), .A2(abar[0]), .ZN(ybar[7]);
  AND2_X1 U24 ( .A1(a[4]), .A2(b[15]), .ZN(y[79]) );
  OR2_X1 U24bar ( .A1(abar[4]), .A2(bbar[15]), .ZN(ybar[79]);
  AND2_X1 U25 ( .A1(a[4]), .A2(b[14]), .ZN(y[78]) );
  OR2_X1 U25bar ( .A1(abar[4]), .A2(bbar[14]), .ZN(ybar[78]);
  AND2_X1 U26 ( .A1(a[4]), .A2(b[13]), .ZN(y[77]) );
  OR2_X1 U26bar ( .A1(abar[4]), .A2(bbar[13]), .ZN(ybar[77]);
  AND2_X1 U27 ( .A1(a[4]), .A2(b[12]), .ZN(y[76]) );
  OR2_X1 U27bar ( .A1(abar[4]), .A2(bbar[12]), .ZN(ybar[76]);
  AND2_X1 U28 ( .A1(a[4]), .A2(b[11]), .ZN(y[75]) );
  OR2_X1 U28bar ( .A1(abar[4]), .A2(bbar[11]), .ZN(ybar[75]);
  AND2_X1 U29 ( .A1(a[4]), .A2(b[10]), .ZN(y[74]) );
  OR2_X1 U29bar ( .A1(abar[4]), .A2(bbar[10]), .ZN(ybar[74]);
  AND2_X1 U30 ( .A1(a[4]), .A2(b[9]), .ZN(y[73]) );
  OR2_X1 U30bar ( .A1(abar[4]), .A2(bbar[9]), .ZN(ybar[73]);
  AND2_X1 U31 ( .A1(a[4]), .A2(b[8]), .ZN(y[72]) );
  OR2_X1 U31bar ( .A1(abar[4]), .A2(bbar[8]), .ZN(ybar[72]);
  AND2_X1 U32 ( .A1(a[4]), .A2(b[7]), .ZN(y[71]) );
  OR2_X1 U32bar ( .A1(abar[4]), .A2(bbar[7]), .ZN(ybar[71]);
  AND2_X1 U33 ( .A1(a[4]), .A2(b[6]), .ZN(y[70]) );
  OR2_X1 U33bar ( .A1(abar[4]), .A2(bbar[6]), .ZN(ybar[70]);
  AND2_X1 U34 ( .A1(b[6]), .A2(a[0]), .ZN(y[6]) );
  OR2_X1 U34bar ( .A1(bbar[6]), .A2(abar[0]), .ZN(ybar[6]);
  AND2_X1 U35 ( .A1(a[4]), .A2(b[5]), .ZN(y[69]) );
  OR2_X1 U35bar ( .A1(abar[4]), .A2(bbar[5]), .ZN(ybar[69]);
  AND2_X1 U36 ( .A1(a[4]), .A2(b[4]), .ZN(y[68]) );
  OR2_X1 U36bar ( .A1(abar[4]), .A2(bbar[4]), .ZN(ybar[68]);
  AND2_X1 U37 ( .A1(a[4]), .A2(b[3]), .ZN(y[67]) );
  OR2_X1 U37bar ( .A1(abar[4]), .A2(bbar[3]), .ZN(ybar[67]);
  AND2_X1 U38 ( .A1(a[4]), .A2(b[2]), .ZN(y[66]) );
  OR2_X1 U38bar ( .A1(abar[4]), .A2(bbar[2]), .ZN(ybar[66]);
  AND2_X1 U39 ( .A1(a[4]), .A2(b[1]), .ZN(y[65]) );
  OR2_X1 U39bar ( .A1(abar[4]), .A2(bbar[1]), .ZN(ybar[65]);
  AND2_X1 U40 ( .A1(a[4]), .A2(b[0]), .ZN(y[64]) );
  OR2_X1 U40bar ( .A1(abar[4]), .A2(bbar[0]), .ZN(ybar[64]);
  AND2_X1 U41 ( .A1(a[3]), .A2(b[15]), .ZN(y[63]) );
  OR2_X1 U41bar ( .A1(abar[3]), .A2(bbar[15]), .ZN(ybar[63]);
  AND2_X1 U42 ( .A1(a[3]), .A2(b[14]), .ZN(y[62]) );
  OR2_X1 U42bar ( .A1(abar[3]), .A2(bbar[14]), .ZN(ybar[62]);
  AND2_X1 U43 ( .A1(a[3]), .A2(b[13]), .ZN(y[61]) );
  OR2_X1 U43bar ( .A1(abar[3]), .A2(bbar[13]), .ZN(ybar[61]);
  AND2_X1 U44 ( .A1(a[3]), .A2(b[12]), .ZN(y[60]) );
  OR2_X1 U44bar ( .A1(abar[3]), .A2(bbar[12]), .ZN(ybar[60]);
  AND2_X1 U45 ( .A1(b[5]), .A2(a[0]), .ZN(y[5]) );
  OR2_X1 U45bar ( .A1(bbar[5]), .A2(abar[0]), .ZN(ybar[5]);
  AND2_X1 U46 ( .A1(a[3]), .A2(b[11]), .ZN(y[59]) );
  OR2_X1 U46bar ( .A1(abar[3]), .A2(bbar[11]), .ZN(ybar[59]);
  AND2_X1 U47 ( .A1(a[3]), .A2(b[10]), .ZN(y[58]) );
  OR2_X1 U47bar ( .A1(abar[3]), .A2(bbar[10]), .ZN(ybar[58]);
  AND2_X1 U48 ( .A1(a[3]), .A2(b[9]), .ZN(y[57]) );
  OR2_X1 U48bar ( .A1(abar[3]), .A2(bbar[9]), .ZN(ybar[57]);
  AND2_X1 U49 ( .A1(a[3]), .A2(b[8]), .ZN(y[56]) );
  OR2_X1 U49bar ( .A1(abar[3]), .A2(bbar[8]), .ZN(ybar[56]);
  AND2_X1 U50 ( .A1(a[3]), .A2(b[7]), .ZN(y[55]) );
  OR2_X1 U50bar ( .A1(abar[3]), .A2(bbar[7]), .ZN(ybar[55]);
  AND2_X1 U51 ( .A1(a[3]), .A2(b[6]), .ZN(y[54]) );
  OR2_X1 U51bar ( .A1(abar[3]), .A2(bbar[6]), .ZN(ybar[54]);
  AND2_X1 U52 ( .A1(a[3]), .A2(b[5]), .ZN(y[53]) );
  OR2_X1 U52bar ( .A1(abar[3]), .A2(bbar[5]), .ZN(ybar[53]);
  AND2_X1 U53 ( .A1(a[3]), .A2(b[4]), .ZN(y[52]) );
  OR2_X1 U53bar ( .A1(abar[3]), .A2(bbar[4]), .ZN(ybar[52]);
  AND2_X1 U54 ( .A1(a[3]), .A2(b[3]), .ZN(y[51]) );
  OR2_X1 U54bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[51]);
  AND2_X1 U55 ( .A1(a[3]), .A2(b[2]), .ZN(y[50]) );
  OR2_X1 U55bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[50]);
  AND2_X1 U56 ( .A1(b[4]), .A2(a[0]), .ZN(y[4]) );
  OR2_X1 U56bar ( .A1(bbar[4]), .A2(abar[0]), .ZN(ybar[4]);
  AND2_X1 U57 ( .A1(a[3]), .A2(b[1]), .ZN(y[49]) );
  OR2_X1 U57bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[49]);
  AND2_X1 U58 ( .A1(a[3]), .A2(b[0]), .ZN(y[48]) );
  OR2_X1 U58bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[48]);
  AND2_X1 U59 ( .A1(a[2]), .A2(b[15]), .ZN(y[47]) );
  OR2_X1 U59bar ( .A1(abar[2]), .A2(bbar[15]), .ZN(ybar[47]);
  AND2_X1 U60 ( .A1(a[2]), .A2(b[14]), .ZN(y[46]) );
  OR2_X1 U60bar ( .A1(abar[2]), .A2(bbar[14]), .ZN(ybar[46]);
  AND2_X1 U61 ( .A1(a[2]), .A2(b[13]), .ZN(y[45]) );
  OR2_X1 U61bar ( .A1(abar[2]), .A2(bbar[13]), .ZN(ybar[45]);
  AND2_X1 U62 ( .A1(a[2]), .A2(b[12]), .ZN(y[44]) );
  OR2_X1 U62bar ( .A1(abar[2]), .A2(bbar[12]), .ZN(ybar[44]);
  AND2_X1 U63 ( .A1(a[2]), .A2(b[11]), .ZN(y[43]) );
  OR2_X1 U63bar ( .A1(abar[2]), .A2(bbar[11]), .ZN(ybar[43]);
  AND2_X1 U64 ( .A1(a[2]), .A2(b[10]), .ZN(y[42]) );
  OR2_X1 U64bar ( .A1(abar[2]), .A2(bbar[10]), .ZN(ybar[42]);
  AND2_X1 U65 ( .A1(a[2]), .A2(b[9]), .ZN(y[41]) );
  OR2_X1 U65bar ( .A1(abar[2]), .A2(bbar[9]), .ZN(ybar[41]);
  AND2_X1 U66 ( .A1(a[2]), .A2(b[8]), .ZN(y[40]) );
  OR2_X1 U66bar ( .A1(abar[2]), .A2(bbar[8]), .ZN(ybar[40]);
  AND2_X1 U67 ( .A1(b[3]), .A2(a[0]), .ZN(y[3]) );
  OR2_X1 U67bar ( .A1(bbar[3]), .A2(abar[0]), .ZN(ybar[3]);
  AND2_X1 U68 ( .A1(a[2]), .A2(b[7]), .ZN(y[39]) );
  OR2_X1 U68bar ( .A1(abar[2]), .A2(bbar[7]), .ZN(ybar[39]);
  AND2_X1 U69 ( .A1(a[2]), .A2(b[6]), .ZN(y[38]) );
  OR2_X1 U69bar ( .A1(abar[2]), .A2(bbar[6]), .ZN(ybar[38]);
  AND2_X1 U70 ( .A1(a[2]), .A2(b[5]), .ZN(y[37]) );
  OR2_X1 U70bar ( .A1(abar[2]), .A2(bbar[5]), .ZN(ybar[37]);
  AND2_X1 U71 ( .A1(a[2]), .A2(b[4]), .ZN(y[36]) );
  OR2_X1 U71bar ( .A1(abar[2]), .A2(bbar[4]), .ZN(ybar[36]);
  AND2_X1 U72 ( .A1(a[2]), .A2(b[3]), .ZN(y[35]) );
  OR2_X1 U72bar ( .A1(abar[2]), .A2(bbar[3]), .ZN(ybar[35]);
  AND2_X1 U73 ( .A1(a[2]), .A2(b[2]), .ZN(y[34]) );
  OR2_X1 U73bar ( .A1(abar[2]), .A2(bbar[2]), .ZN(ybar[34]);
  AND2_X1 U74 ( .A1(a[2]), .A2(b[1]), .ZN(y[33]) );
  OR2_X1 U74bar ( .A1(abar[2]), .A2(bbar[1]), .ZN(ybar[33]);
  AND2_X1 U75 ( .A1(a[2]), .A2(b[0]), .ZN(y[32]) );
  OR2_X1 U75bar ( .A1(abar[2]), .A2(bbar[0]), .ZN(ybar[32]);
  AND2_X1 U76 ( .A1(a[1]), .A2(b[15]), .ZN(y[31]) );
  OR2_X1 U76bar ( .A1(abar[1]), .A2(bbar[15]), .ZN(ybar[31]);
  AND2_X1 U77 ( .A1(a[1]), .A2(b[14]), .ZN(y[30]) );
  OR2_X1 U77bar ( .A1(abar[1]), .A2(bbar[14]), .ZN(ybar[30]);
  AND2_X1 U78 ( .A1(b[2]), .A2(a[0]), .ZN(y[2]) );
  OR2_X1 U78bar ( .A1(bbar[2]), .A2(abar[0]), .ZN(ybar[2]);
  AND2_X1 U79 ( .A1(a[1]), .A2(b[13]), .ZN(y[29]) );
  OR2_X1 U79bar ( .A1(abar[1]), .A2(bbar[13]), .ZN(ybar[29]);
  AND2_X1 U80 ( .A1(a[1]), .A2(b[12]), .ZN(y[28]) );
  OR2_X1 U80bar ( .A1(abar[1]), .A2(bbar[12]), .ZN(ybar[28]);
  AND2_X1 U81 ( .A1(a[1]), .A2(b[11]), .ZN(y[27]) );
  OR2_X1 U81bar ( .A1(abar[1]), .A2(bbar[11]), .ZN(ybar[27]);
  AND2_X1 U82 ( .A1(a[1]), .A2(b[10]), .ZN(y[26]) );
  OR2_X1 U82bar ( .A1(abar[1]), .A2(bbar[10]), .ZN(ybar[26]);
  AND2_X1 U83 ( .A1(a[1]), .A2(b[9]), .ZN(y[25]) );
  OR2_X1 U83bar ( .A1(abar[1]), .A2(bbar[9]), .ZN(ybar[25]);
  AND2_X1 U84 ( .A1(a[15]), .A2(b[15]), .ZN(y[255]) );
  OR2_X1 U84bar ( .A1(abar[15]), .A2(bbar[15]), .ZN(ybar[255]);
  AND2_X1 U85 ( .A1(a[15]), .A2(b[14]), .ZN(y[254]) );
  OR2_X1 U85bar ( .A1(abar[15]), .A2(bbar[14]), .ZN(ybar[254]);
  AND2_X1 U86 ( .A1(a[15]), .A2(b[13]), .ZN(y[253]) );
  OR2_X1 U86bar ( .A1(abar[15]), .A2(bbar[13]), .ZN(ybar[253]);
  AND2_X1 U87 ( .A1(a[15]), .A2(b[12]), .ZN(y[252]) );
  OR2_X1 U87bar ( .A1(abar[15]), .A2(bbar[12]), .ZN(ybar[252]);
  AND2_X1 U88 ( .A1(a[15]), .A2(b[11]), .ZN(y[251]) );
  OR2_X1 U88bar ( .A1(abar[15]), .A2(bbar[11]), .ZN(ybar[251]);
  AND2_X1 U89 ( .A1(a[15]), .A2(b[10]), .ZN(y[250]) );
  OR2_X1 U89bar ( .A1(abar[15]), .A2(bbar[10]), .ZN(ybar[250]);
  AND2_X1 U90 ( .A1(a[1]), .A2(b[8]), .ZN(y[24]) );
  OR2_X1 U90bar ( .A1(abar[1]), .A2(bbar[8]), .ZN(ybar[24]);
  AND2_X1 U91 ( .A1(a[15]), .A2(b[9]), .ZN(y[249]) );
  OR2_X1 U91bar ( .A1(abar[15]), .A2(bbar[9]), .ZN(ybar[249]);
  AND2_X1 U92 ( .A1(a[15]), .A2(b[8]), .ZN(y[248]) );
  OR2_X1 U92bar ( .A1(abar[15]), .A2(bbar[8]), .ZN(ybar[248]);
  AND2_X1 U93 ( .A1(a[15]), .A2(b[7]), .ZN(y[247]) );
  OR2_X1 U93bar ( .A1(abar[15]), .A2(bbar[7]), .ZN(ybar[247]);
  AND2_X1 U94 ( .A1(a[15]), .A2(b[6]), .ZN(y[246]) );
  OR2_X1 U94bar ( .A1(abar[15]), .A2(bbar[6]), .ZN(ybar[246]);
  AND2_X1 U95 ( .A1(a[15]), .A2(b[5]), .ZN(y[245]) );
  OR2_X1 U95bar ( .A1(abar[15]), .A2(bbar[5]), .ZN(ybar[245]);
  AND2_X1 U96 ( .A1(a[15]), .A2(b[4]), .ZN(y[244]) );
  OR2_X1 U96bar ( .A1(abar[15]), .A2(bbar[4]), .ZN(ybar[244]);
  AND2_X1 U97 ( .A1(a[15]), .A2(b[3]), .ZN(y[243]) );
  OR2_X1 U97bar ( .A1(abar[15]), .A2(bbar[3]), .ZN(ybar[243]);
  AND2_X1 U98 ( .A1(a[15]), .A2(b[2]), .ZN(y[242]) );
  OR2_X1 U98bar ( .A1(abar[15]), .A2(bbar[2]), .ZN(ybar[242]);
  AND2_X1 U99 ( .A1(a[15]), .A2(b[1]), .ZN(y[241]) );
  OR2_X1 U99bar ( .A1(abar[15]), .A2(bbar[1]), .ZN(ybar[241]);
  AND2_X1 U100 ( .A1(a[15]), .A2(b[0]), .ZN(y[240]) );
  OR2_X1 U100bar ( .A1(abar[15]), .A2(bbar[0]), .ZN(ybar[240]);
  AND2_X1 U101 ( .A1(a[1]), .A2(b[7]), .ZN(y[23]) );
  OR2_X1 U101bar ( .A1(abar[1]), .A2(bbar[7]), .ZN(ybar[23]);
  AND2_X1 U102 ( .A1(a[14]), .A2(b[15]), .ZN(y[239]) );
  OR2_X1 U102bar ( .A1(abar[14]), .A2(bbar[15]), .ZN(ybar[239]);
  AND2_X1 U103 ( .A1(a[14]), .A2(b[14]), .ZN(y[238]) );
  OR2_X1 U103bar ( .A1(abar[14]), .A2(bbar[14]), .ZN(ybar[238]);
  AND2_X1 U104 ( .A1(a[14]), .A2(b[13]), .ZN(y[237]) );
  OR2_X1 U104bar ( .A1(abar[14]), .A2(bbar[13]), .ZN(ybar[237]);
  AND2_X1 U105 ( .A1(a[14]), .A2(b[12]), .ZN(y[236]) );
  OR2_X1 U105bar ( .A1(abar[14]), .A2(bbar[12]), .ZN(ybar[236]);
  AND2_X1 U106 ( .A1(a[14]), .A2(b[11]), .ZN(y[235]) );
  OR2_X1 U106bar ( .A1(abar[14]), .A2(bbar[11]), .ZN(ybar[235]);
  AND2_X1 U107 ( .A1(a[14]), .A2(b[10]), .ZN(y[234]) );
  OR2_X1 U107bar ( .A1(abar[14]), .A2(bbar[10]), .ZN(ybar[234]);
  AND2_X1 U108 ( .A1(a[14]), .A2(b[9]), .ZN(y[233]) );
  OR2_X1 U108bar ( .A1(abar[14]), .A2(bbar[9]), .ZN(ybar[233]);
  AND2_X1 U109 ( .A1(a[14]), .A2(b[8]), .ZN(y[232]) );
  OR2_X1 U109bar ( .A1(abar[14]), .A2(bbar[8]), .ZN(ybar[232]);
  AND2_X1 U110 ( .A1(a[14]), .A2(b[7]), .ZN(y[231]) );
  OR2_X1 U110bar ( .A1(abar[14]), .A2(bbar[7]), .ZN(ybar[231]);
  AND2_X1 U111 ( .A1(a[14]), .A2(b[6]), .ZN(y[230]) );
  OR2_X1 U111bar ( .A1(abar[14]), .A2(bbar[6]), .ZN(ybar[230]);
  AND2_X1 U112 ( .A1(a[1]), .A2(b[6]), .ZN(y[22]) );
  OR2_X1 U112bar ( .A1(abar[1]), .A2(bbar[6]), .ZN(ybar[22]);
  AND2_X1 U113 ( .A1(a[14]), .A2(b[5]), .ZN(y[229]) );
  OR2_X1 U113bar ( .A1(abar[14]), .A2(bbar[5]), .ZN(ybar[229]);
  AND2_X1 U114 ( .A1(a[14]), .A2(b[4]), .ZN(y[228]) );
  OR2_X1 U114bar ( .A1(abar[14]), .A2(bbar[4]), .ZN(ybar[228]);
  AND2_X1 U115 ( .A1(a[14]), .A2(b[3]), .ZN(y[227]) );
  OR2_X1 U115bar ( .A1(abar[14]), .A2(bbar[3]), .ZN(ybar[227]);
  AND2_X1 U116 ( .A1(a[14]), .A2(b[2]), .ZN(y[226]) );
  OR2_X1 U116bar ( .A1(abar[14]), .A2(bbar[2]), .ZN(ybar[226]);
  AND2_X1 U117 ( .A1(a[14]), .A2(b[1]), .ZN(y[225]) );
  OR2_X1 U117bar ( .A1(abar[14]), .A2(bbar[1]), .ZN(ybar[225]);
  AND2_X1 U118 ( .A1(a[14]), .A2(b[0]), .ZN(y[224]) );
  OR2_X1 U118bar ( .A1(abar[14]), .A2(bbar[0]), .ZN(ybar[224]);
  AND2_X1 U119 ( .A1(a[13]), .A2(b[15]), .ZN(y[223]) );
  OR2_X1 U119bar ( .A1(abar[13]), .A2(bbar[15]), .ZN(ybar[223]);
  AND2_X1 U120 ( .A1(a[13]), .A2(b[14]), .ZN(y[222]) );
  OR2_X1 U120bar ( .A1(abar[13]), .A2(bbar[14]), .ZN(ybar[222]);
  AND2_X1 U121 ( .A1(a[13]), .A2(b[13]), .ZN(y[221]) );
  OR2_X1 U121bar ( .A1(abar[13]), .A2(bbar[13]), .ZN(ybar[221]);
  AND2_X1 U122 ( .A1(a[13]), .A2(b[12]), .ZN(y[220]) );
  OR2_X1 U122bar ( .A1(abar[13]), .A2(bbar[12]), .ZN(ybar[220]);
  AND2_X1 U123 ( .A1(a[1]), .A2(b[5]), .ZN(y[21]) );
  OR2_X1 U123bar ( .A1(abar[1]), .A2(bbar[5]), .ZN(ybar[21]);
  AND2_X1 U124 ( .A1(a[13]), .A2(b[11]), .ZN(y[219]) );
  OR2_X1 U124bar ( .A1(abar[13]), .A2(bbar[11]), .ZN(ybar[219]);
  AND2_X1 U125 ( .A1(a[13]), .A2(b[10]), .ZN(y[218]) );
  OR2_X1 U125bar ( .A1(abar[13]), .A2(bbar[10]), .ZN(ybar[218]);
  AND2_X1 U126 ( .A1(a[13]), .A2(b[9]), .ZN(y[217]) );
  OR2_X1 U126bar ( .A1(abar[13]), .A2(bbar[9]), .ZN(ybar[217]);
  AND2_X1 U127 ( .A1(a[13]), .A2(b[8]), .ZN(y[216]) );
  OR2_X1 U127bar ( .A1(abar[13]), .A2(bbar[8]), .ZN(ybar[216]);
  AND2_X1 U128 ( .A1(a[13]), .A2(b[7]), .ZN(y[215]) );
  OR2_X1 U128bar ( .A1(abar[13]), .A2(bbar[7]), .ZN(ybar[215]);
  AND2_X1 U129 ( .A1(a[13]), .A2(b[6]), .ZN(y[214]) );
  OR2_X1 U129bar ( .A1(abar[13]), .A2(bbar[6]), .ZN(ybar[214]);
  AND2_X1 U130 ( .A1(a[13]), .A2(b[5]), .ZN(y[213]) );
  OR2_X1 U130bar ( .A1(abar[13]), .A2(bbar[5]), .ZN(ybar[213]);
  AND2_X1 U131 ( .A1(a[13]), .A2(b[4]), .ZN(y[212]) );
  OR2_X1 U131bar ( .A1(abar[13]), .A2(bbar[4]), .ZN(ybar[212]);
  AND2_X1 U132 ( .A1(a[13]), .A2(b[3]), .ZN(y[211]) );
  OR2_X1 U132bar ( .A1(abar[13]), .A2(bbar[3]), .ZN(ybar[211]);
  AND2_X1 U133 ( .A1(a[13]), .A2(b[2]), .ZN(y[210]) );
  OR2_X1 U133bar ( .A1(abar[13]), .A2(bbar[2]), .ZN(ybar[210]);
  AND2_X1 U134 ( .A1(a[1]), .A2(b[4]), .ZN(y[20]) );
  OR2_X1 U134bar ( .A1(abar[1]), .A2(bbar[4]), .ZN(ybar[20]);
  AND2_X1 U135 ( .A1(a[13]), .A2(b[1]), .ZN(y[209]) );
  OR2_X1 U135bar ( .A1(abar[13]), .A2(bbar[1]), .ZN(ybar[209]);
  AND2_X1 U136 ( .A1(a[13]), .A2(b[0]), .ZN(y[208]) );
  OR2_X1 U136bar ( .A1(abar[13]), .A2(bbar[0]), .ZN(ybar[208]);
  AND2_X1 U137 ( .A1(a[12]), .A2(b[15]), .ZN(y[207]) );
  OR2_X1 U137bar ( .A1(abar[12]), .A2(bbar[15]), .ZN(ybar[207]);
  AND2_X1 U138 ( .A1(a[12]), .A2(b[14]), .ZN(y[206]) );
  OR2_X1 U138bar ( .A1(abar[12]), .A2(bbar[14]), .ZN(ybar[206]);
  AND2_X1 U139 ( .A1(a[12]), .A2(b[13]), .ZN(y[205]) );
  OR2_X1 U139bar ( .A1(abar[12]), .A2(bbar[13]), .ZN(ybar[205]);
  AND2_X1 U140 ( .A1(a[12]), .A2(b[12]), .ZN(y[204]) );
  OR2_X1 U140bar ( .A1(abar[12]), .A2(bbar[12]), .ZN(ybar[204]);
  AND2_X1 U141 ( .A1(a[12]), .A2(b[11]), .ZN(y[203]) );
  OR2_X1 U141bar ( .A1(abar[12]), .A2(bbar[11]), .ZN(ybar[203]);
  AND2_X1 U142 ( .A1(a[12]), .A2(b[10]), .ZN(y[202]) );
  OR2_X1 U142bar ( .A1(abar[12]), .A2(bbar[10]), .ZN(ybar[202]);
  AND2_X1 U143 ( .A1(a[12]), .A2(b[9]), .ZN(y[201]) );
  OR2_X1 U143bar ( .A1(abar[12]), .A2(bbar[9]), .ZN(ybar[201]);
  AND2_X1 U144 ( .A1(a[12]), .A2(b[8]), .ZN(y[200]) );
  OR2_X1 U144bar ( .A1(abar[12]), .A2(bbar[8]), .ZN(ybar[200]);
  AND2_X1 U145 ( .A1(b[1]), .A2(a[0]), .ZN(y[1]) );
  OR2_X1 U145bar ( .A1(bbar[1]), .A2(abar[0]), .ZN(ybar[1]);
  AND2_X1 U146 ( .A1(a[1]), .A2(b[3]), .ZN(y[19]) );
  OR2_X1 U146bar ( .A1(abar[1]), .A2(bbar[3]), .ZN(ybar[19]);
  AND2_X1 U147 ( .A1(a[12]), .A2(b[7]), .ZN(y[199]) );
  OR2_X1 U147bar ( .A1(abar[12]), .A2(bbar[7]), .ZN(ybar[199]);
  AND2_X1 U148 ( .A1(a[12]), .A2(b[6]), .ZN(y[198]) );
  OR2_X1 U148bar ( .A1(abar[12]), .A2(bbar[6]), .ZN(ybar[198]);
  AND2_X1 U149 ( .A1(a[12]), .A2(b[5]), .ZN(y[197]) );
  OR2_X1 U149bar ( .A1(abar[12]), .A2(bbar[5]), .ZN(ybar[197]);
  AND2_X1 U150 ( .A1(a[12]), .A2(b[4]), .ZN(y[196]) );
  OR2_X1 U150bar ( .A1(abar[12]), .A2(bbar[4]), .ZN(ybar[196]);
  AND2_X1 U151 ( .A1(a[12]), .A2(b[3]), .ZN(y[195]) );
  OR2_X1 U151bar ( .A1(abar[12]), .A2(bbar[3]), .ZN(ybar[195]);
  AND2_X1 U152 ( .A1(a[12]), .A2(b[2]), .ZN(y[194]) );
  OR2_X1 U152bar ( .A1(abar[12]), .A2(bbar[2]), .ZN(ybar[194]);
  AND2_X1 U153 ( .A1(a[12]), .A2(b[1]), .ZN(y[193]) );
  OR2_X1 U153bar ( .A1(abar[12]), .A2(bbar[1]), .ZN(ybar[193]);
  AND2_X1 U154 ( .A1(a[12]), .A2(b[0]), .ZN(y[192]) );
  OR2_X1 U154bar ( .A1(abar[12]), .A2(bbar[0]), .ZN(ybar[192]);
  AND2_X1 U155 ( .A1(a[11]), .A2(b[15]), .ZN(y[191]) );
  OR2_X1 U155bar ( .A1(abar[11]), .A2(bbar[15]), .ZN(ybar[191]);
  AND2_X1 U156 ( .A1(a[11]), .A2(b[14]), .ZN(y[190]) );
  OR2_X1 U156bar ( .A1(abar[11]), .A2(bbar[14]), .ZN(ybar[190]);
  AND2_X1 U157 ( .A1(a[1]), .A2(b[2]), .ZN(y[18]) );
  OR2_X1 U157bar ( .A1(abar[1]), .A2(bbar[2]), .ZN(ybar[18]);
  AND2_X1 U158 ( .A1(a[11]), .A2(b[13]), .ZN(y[189]) );
  OR2_X1 U158bar ( .A1(abar[11]), .A2(bbar[13]), .ZN(ybar[189]);
  AND2_X1 U159 ( .A1(a[11]), .A2(b[12]), .ZN(y[188]) );
  OR2_X1 U159bar ( .A1(abar[11]), .A2(bbar[12]), .ZN(ybar[188]);
  AND2_X1 U160 ( .A1(a[11]), .A2(b[11]), .ZN(y[187]) );
  OR2_X1 U160bar ( .A1(abar[11]), .A2(bbar[11]), .ZN(ybar[187]);
  AND2_X1 U161 ( .A1(a[11]), .A2(b[10]), .ZN(y[186]) );
  OR2_X1 U161bar ( .A1(abar[11]), .A2(bbar[10]), .ZN(ybar[186]);
  AND2_X1 U162 ( .A1(a[11]), .A2(b[9]), .ZN(y[185]) );
  OR2_X1 U162bar ( .A1(abar[11]), .A2(bbar[9]), .ZN(ybar[185]);
  AND2_X1 U163 ( .A1(a[11]), .A2(b[8]), .ZN(y[184]) );
  OR2_X1 U163bar ( .A1(abar[11]), .A2(bbar[8]), .ZN(ybar[184]);
  AND2_X1 U164 ( .A1(a[11]), .A2(b[7]), .ZN(y[183]) );
  OR2_X1 U164bar ( .A1(abar[11]), .A2(bbar[7]), .ZN(ybar[183]);
  AND2_X1 U165 ( .A1(a[11]), .A2(b[6]), .ZN(y[182]) );
  OR2_X1 U165bar ( .A1(abar[11]), .A2(bbar[6]), .ZN(ybar[182]);
  AND2_X1 U166 ( .A1(a[11]), .A2(b[5]), .ZN(y[181]) );
  OR2_X1 U166bar ( .A1(abar[11]), .A2(bbar[5]), .ZN(ybar[181]);
  AND2_X1 U167 ( .A1(a[11]), .A2(b[4]), .ZN(y[180]) );
  OR2_X1 U167bar ( .A1(abar[11]), .A2(bbar[4]), .ZN(ybar[180]);
  AND2_X1 U168 ( .A1(a[1]), .A2(b[1]), .ZN(y[17]) );
  OR2_X1 U168bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[17]);
  AND2_X1 U169 ( .A1(a[11]), .A2(b[3]), .ZN(y[179]) );
  OR2_X1 U169bar ( .A1(abar[11]), .A2(bbar[3]), .ZN(ybar[179]);
  AND2_X1 U170 ( .A1(a[11]), .A2(b[2]), .ZN(y[178]) );
  OR2_X1 U170bar ( .A1(abar[11]), .A2(bbar[2]), .ZN(ybar[178]);
  AND2_X1 U171 ( .A1(a[11]), .A2(b[1]), .ZN(y[177]) );
  OR2_X1 U171bar ( .A1(abar[11]), .A2(bbar[1]), .ZN(ybar[177]);
  AND2_X1 U172 ( .A1(a[11]), .A2(b[0]), .ZN(y[176]) );
  OR2_X1 U172bar ( .A1(abar[11]), .A2(bbar[0]), .ZN(ybar[176]);
  AND2_X1 U173 ( .A1(a[10]), .A2(b[15]), .ZN(y[175]) );
  OR2_X1 U173bar ( .A1(abar[10]), .A2(bbar[15]), .ZN(ybar[175]);
  AND2_X1 U174 ( .A1(a[10]), .A2(b[14]), .ZN(y[174]) );
  OR2_X1 U174bar ( .A1(abar[10]), .A2(bbar[14]), .ZN(ybar[174]);
  AND2_X1 U175 ( .A1(a[10]), .A2(b[13]), .ZN(y[173]) );
  OR2_X1 U175bar ( .A1(abar[10]), .A2(bbar[13]), .ZN(ybar[173]);
  AND2_X1 U176 ( .A1(a[10]), .A2(b[12]), .ZN(y[172]) );
  OR2_X1 U176bar ( .A1(abar[10]), .A2(bbar[12]), .ZN(ybar[172]);
  AND2_X1 U177 ( .A1(a[10]), .A2(b[11]), .ZN(y[171]) );
  OR2_X1 U177bar ( .A1(abar[10]), .A2(bbar[11]), .ZN(ybar[171]);
  AND2_X1 U178 ( .A1(a[10]), .A2(b[10]), .ZN(y[170]) );
  OR2_X1 U178bar ( .A1(abar[10]), .A2(bbar[10]), .ZN(ybar[170]);
  AND2_X1 U179 ( .A1(a[1]), .A2(b[0]), .ZN(y[16]) );
  OR2_X1 U179bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[16]);
  AND2_X1 U180 ( .A1(a[10]), .A2(b[9]), .ZN(y[169]) );
  OR2_X1 U180bar ( .A1(abar[10]), .A2(bbar[9]), .ZN(ybar[169]);
  AND2_X1 U181 ( .A1(a[10]), .A2(b[8]), .ZN(y[168]) );
  OR2_X1 U181bar ( .A1(abar[10]), .A2(bbar[8]), .ZN(ybar[168]);
  AND2_X1 U182 ( .A1(a[10]), .A2(b[7]), .ZN(y[167]) );
  OR2_X1 U182bar ( .A1(abar[10]), .A2(bbar[7]), .ZN(ybar[167]);
  AND2_X1 U183 ( .A1(a[10]), .A2(b[6]), .ZN(y[166]) );
  OR2_X1 U183bar ( .A1(abar[10]), .A2(bbar[6]), .ZN(ybar[166]);
  AND2_X1 U184 ( .A1(a[10]), .A2(b[5]), .ZN(y[165]) );
  OR2_X1 U184bar ( .A1(abar[10]), .A2(bbar[5]), .ZN(ybar[165]);
  AND2_X1 U185 ( .A1(a[10]), .A2(b[4]), .ZN(y[164]) );
  OR2_X1 U185bar ( .A1(abar[10]), .A2(bbar[4]), .ZN(ybar[164]);
  AND2_X1 U186 ( .A1(a[10]), .A2(b[3]), .ZN(y[163]) );
  OR2_X1 U186bar ( .A1(abar[10]), .A2(bbar[3]), .ZN(ybar[163]);
  AND2_X1 U187 ( .A1(a[10]), .A2(b[2]), .ZN(y[162]) );
  OR2_X1 U187bar ( .A1(abar[10]), .A2(bbar[2]), .ZN(ybar[162]);
  AND2_X1 U188 ( .A1(a[10]), .A2(b[1]), .ZN(y[161]) );
  OR2_X1 U188bar ( .A1(abar[10]), .A2(bbar[1]), .ZN(ybar[161]);
  AND2_X1 U189 ( .A1(a[10]), .A2(b[0]), .ZN(y[160]) );
  OR2_X1 U189bar ( .A1(abar[10]), .A2(bbar[0]), .ZN(ybar[160]);
  AND2_X1 U190 ( .A1(b[15]), .A2(a[0]), .ZN(y[15]) );
  OR2_X1 U190bar ( .A1(bbar[15]), .A2(abar[0]), .ZN(ybar[15]);
  AND2_X1 U191 ( .A1(a[9]), .A2(b[15]), .ZN(y[159]) );
  OR2_X1 U191bar ( .A1(abar[9]), .A2(bbar[15]), .ZN(ybar[159]);
  AND2_X1 U192 ( .A1(a[9]), .A2(b[14]), .ZN(y[158]) );
  OR2_X1 U192bar ( .A1(abar[9]), .A2(bbar[14]), .ZN(ybar[158]);
  AND2_X1 U193 ( .A1(a[9]), .A2(b[13]), .ZN(y[157]) );
  OR2_X1 U193bar ( .A1(abar[9]), .A2(bbar[13]), .ZN(ybar[157]);
  AND2_X1 U194 ( .A1(a[9]), .A2(b[12]), .ZN(y[156]) );
  OR2_X1 U194bar ( .A1(abar[9]), .A2(bbar[12]), .ZN(ybar[156]);
  AND2_X1 U195 ( .A1(a[9]), .A2(b[11]), .ZN(y[155]) );
  OR2_X1 U195bar ( .A1(abar[9]), .A2(bbar[11]), .ZN(ybar[155]);
  AND2_X1 U196 ( .A1(a[9]), .A2(b[10]), .ZN(y[154]) );
  OR2_X1 U196bar ( .A1(abar[9]), .A2(bbar[10]), .ZN(ybar[154]);
  AND2_X1 U197 ( .A1(a[9]), .A2(b[9]), .ZN(y[153]) );
  OR2_X1 U197bar ( .A1(abar[9]), .A2(bbar[9]), .ZN(ybar[153]);
  AND2_X1 U198 ( .A1(a[9]), .A2(b[8]), .ZN(y[152]) );
  OR2_X1 U198bar ( .A1(abar[9]), .A2(bbar[8]), .ZN(ybar[152]);
  AND2_X1 U199 ( .A1(a[9]), .A2(b[7]), .ZN(y[151]) );
  OR2_X1 U199bar ( .A1(abar[9]), .A2(bbar[7]), .ZN(ybar[151]);
  AND2_X1 U200 ( .A1(a[9]), .A2(b[6]), .ZN(y[150]) );
  OR2_X1 U200bar ( .A1(abar[9]), .A2(bbar[6]), .ZN(ybar[150]);
  AND2_X1 U201 ( .A1(b[14]), .A2(a[0]), .ZN(y[14]) );
  OR2_X1 U201bar ( .A1(bbar[14]), .A2(abar[0]), .ZN(ybar[14]);
  AND2_X1 U202 ( .A1(a[9]), .A2(b[5]), .ZN(y[149]) );
  OR2_X1 U202bar ( .A1(abar[9]), .A2(bbar[5]), .ZN(ybar[149]);
  AND2_X1 U203 ( .A1(a[9]), .A2(b[4]), .ZN(y[148]) );
  OR2_X1 U203bar ( .A1(abar[9]), .A2(bbar[4]), .ZN(ybar[148]);
  AND2_X1 U204 ( .A1(a[9]), .A2(b[3]), .ZN(y[147]) );
  OR2_X1 U204bar ( .A1(abar[9]), .A2(bbar[3]), .ZN(ybar[147]);
  AND2_X1 U205 ( .A1(a[9]), .A2(b[2]), .ZN(y[146]) );
  OR2_X1 U205bar ( .A1(abar[9]), .A2(bbar[2]), .ZN(ybar[146]);
  AND2_X1 U206 ( .A1(a[9]), .A2(b[1]), .ZN(y[145]) );
  OR2_X1 U206bar ( .A1(abar[9]), .A2(bbar[1]), .ZN(ybar[145]);
  AND2_X1 U207 ( .A1(a[9]), .A2(b[0]), .ZN(y[144]) );
  OR2_X1 U207bar ( .A1(abar[9]), .A2(bbar[0]), .ZN(ybar[144]);
  AND2_X1 U208 ( .A1(a[8]), .A2(b[15]), .ZN(y[143]) );
  OR2_X1 U208bar ( .A1(abar[8]), .A2(bbar[15]), .ZN(ybar[143]);
  AND2_X1 U209 ( .A1(a[8]), .A2(b[14]), .ZN(y[142]) );
  OR2_X1 U209bar ( .A1(abar[8]), .A2(bbar[14]), .ZN(ybar[142]);
  AND2_X1 U210 ( .A1(a[8]), .A2(b[13]), .ZN(y[141]) );
  OR2_X1 U210bar ( .A1(abar[8]), .A2(bbar[13]), .ZN(ybar[141]);
  AND2_X1 U211 ( .A1(a[8]), .A2(b[12]), .ZN(y[140]) );
  OR2_X1 U211bar ( .A1(abar[8]), .A2(bbar[12]), .ZN(ybar[140]);
  AND2_X1 U212 ( .A1(b[13]), .A2(a[0]), .ZN(y[13]) );
  OR2_X1 U212bar ( .A1(bbar[13]), .A2(abar[0]), .ZN(ybar[13]);
  AND2_X1 U213 ( .A1(a[8]), .A2(b[11]), .ZN(y[139]) );
  OR2_X1 U213bar ( .A1(abar[8]), .A2(bbar[11]), .ZN(ybar[139]);
  AND2_X1 U214 ( .A1(a[8]), .A2(b[10]), .ZN(y[138]) );
  OR2_X1 U214bar ( .A1(abar[8]), .A2(bbar[10]), .ZN(ybar[138]);
  AND2_X1 U215 ( .A1(a[8]), .A2(b[9]), .ZN(y[137]) );
  OR2_X1 U215bar ( .A1(abar[8]), .A2(bbar[9]), .ZN(ybar[137]);
  AND2_X1 U216 ( .A1(a[8]), .A2(b[8]), .ZN(y[136]) );
  OR2_X1 U216bar ( .A1(abar[8]), .A2(bbar[8]), .ZN(ybar[136]);
  AND2_X1 U217 ( .A1(a[8]), .A2(b[7]), .ZN(y[135]) );
  OR2_X1 U217bar ( .A1(abar[8]), .A2(bbar[7]), .ZN(ybar[135]);
  AND2_X1 U218 ( .A1(a[8]), .A2(b[6]), .ZN(y[134]) );
  OR2_X1 U218bar ( .A1(abar[8]), .A2(bbar[6]), .ZN(ybar[134]);
  AND2_X1 U219 ( .A1(a[8]), .A2(b[5]), .ZN(y[133]) );
  OR2_X1 U219bar ( .A1(abar[8]), .A2(bbar[5]), .ZN(ybar[133]);
  AND2_X1 U220 ( .A1(a[8]), .A2(b[4]), .ZN(y[132]) );
  OR2_X1 U220bar ( .A1(abar[8]), .A2(bbar[4]), .ZN(ybar[132]);
  AND2_X1 U221 ( .A1(a[8]), .A2(b[3]), .ZN(y[131]) );
  OR2_X1 U221bar ( .A1(abar[8]), .A2(bbar[3]), .ZN(ybar[131]);
  AND2_X1 U222 ( .A1(a[8]), .A2(b[2]), .ZN(y[130]) );
  OR2_X1 U222bar ( .A1(abar[8]), .A2(bbar[2]), .ZN(ybar[130]);
  AND2_X1 U223 ( .A1(b[12]), .A2(a[0]), .ZN(y[12]) );
  OR2_X1 U223bar ( .A1(bbar[12]), .A2(abar[0]), .ZN(ybar[12]);
  AND2_X1 U224 ( .A1(a[8]), .A2(b[1]), .ZN(y[129]) );
  OR2_X1 U224bar ( .A1(abar[8]), .A2(bbar[1]), .ZN(ybar[129]);
  AND2_X1 U225 ( .A1(a[8]), .A2(b[0]), .ZN(y[128]) );
  OR2_X1 U225bar ( .A1(abar[8]), .A2(bbar[0]), .ZN(ybar[128]);
  AND2_X1 U226 ( .A1(a[7]), .A2(b[15]), .ZN(y[127]) );
  OR2_X1 U226bar ( .A1(abar[7]), .A2(bbar[15]), .ZN(ybar[127]);
  AND2_X1 U227 ( .A1(a[7]), .A2(b[14]), .ZN(y[126]) );
  OR2_X1 U227bar ( .A1(abar[7]), .A2(bbar[14]), .ZN(ybar[126]);
  AND2_X1 U228 ( .A1(a[7]), .A2(b[13]), .ZN(y[125]) );
  OR2_X1 U228bar ( .A1(abar[7]), .A2(bbar[13]), .ZN(ybar[125]);
  AND2_X1 U229 ( .A1(a[7]), .A2(b[12]), .ZN(y[124]) );
  OR2_X1 U229bar ( .A1(abar[7]), .A2(bbar[12]), .ZN(ybar[124]);
  AND2_X1 U230 ( .A1(a[7]), .A2(b[11]), .ZN(y[123]) );
  OR2_X1 U230bar ( .A1(abar[7]), .A2(bbar[11]), .ZN(ybar[123]);
  AND2_X1 U231 ( .A1(a[7]), .A2(b[10]), .ZN(y[122]) );
  OR2_X1 U231bar ( .A1(abar[7]), .A2(bbar[10]), .ZN(ybar[122]);
  AND2_X1 U232 ( .A1(a[7]), .A2(b[9]), .ZN(y[121]) );
  OR2_X1 U232bar ( .A1(abar[7]), .A2(bbar[9]), .ZN(ybar[121]);
  AND2_X1 U233 ( .A1(a[7]), .A2(b[8]), .ZN(y[120]) );
  OR2_X1 U233bar ( .A1(abar[7]), .A2(bbar[8]), .ZN(ybar[120]);
  AND2_X1 U234 ( .A1(b[11]), .A2(a[0]), .ZN(y[11]) );
  OR2_X1 U234bar ( .A1(bbar[11]), .A2(abar[0]), .ZN(ybar[11]);
  AND2_X1 U235 ( .A1(a[7]), .A2(b[7]), .ZN(y[119]) );
  OR2_X1 U235bar ( .A1(abar[7]), .A2(bbar[7]), .ZN(ybar[119]);
  AND2_X1 U236 ( .A1(a[7]), .A2(b[6]), .ZN(y[118]) );
  OR2_X1 U236bar ( .A1(abar[7]), .A2(bbar[6]), .ZN(ybar[118]);
  AND2_X1 U237 ( .A1(a[7]), .A2(b[5]), .ZN(y[117]) );
  OR2_X1 U237bar ( .A1(abar[7]), .A2(bbar[5]), .ZN(ybar[117]);
  AND2_X1 U238 ( .A1(a[7]), .A2(b[4]), .ZN(y[116]) );
  OR2_X1 U238bar ( .A1(abar[7]), .A2(bbar[4]), .ZN(ybar[116]);
  AND2_X1 U239 ( .A1(a[7]), .A2(b[3]), .ZN(y[115]) );
  OR2_X1 U239bar ( .A1(abar[7]), .A2(bbar[3]), .ZN(ybar[115]);
  AND2_X1 U240 ( .A1(a[7]), .A2(b[2]), .ZN(y[114]) );
  OR2_X1 U240bar ( .A1(abar[7]), .A2(bbar[2]), .ZN(ybar[114]);
  AND2_X1 U241 ( .A1(a[7]), .A2(b[1]), .ZN(y[113]) );
  OR2_X1 U241bar ( .A1(abar[7]), .A2(bbar[1]), .ZN(ybar[113]);
  AND2_X1 U242 ( .A1(a[7]), .A2(b[0]), .ZN(y[112]) );
  OR2_X1 U242bar ( .A1(abar[7]), .A2(bbar[0]), .ZN(ybar[112]);
  AND2_X1 U243 ( .A1(b[15]), .A2(a[6]), .ZN(y[111]) );
  OR2_X1 U243bar ( .A1(bbar[15]), .A2(abar[6]), .ZN(ybar[111]);
  AND2_X1 U244 ( .A1(b[14]), .A2(a[6]), .ZN(y[110]) );
  OR2_X1 U244bar ( .A1(bbar[14]), .A2(abar[6]), .ZN(ybar[110]);
  AND2_X1 U245 ( .A1(b[10]), .A2(a[0]), .ZN(y[10]) );
  OR2_X1 U245bar ( .A1(bbar[10]), .A2(abar[0]), .ZN(ybar[10]);
  AND2_X1 U246 ( .A1(b[13]), .A2(a[6]), .ZN(y[109]) );
  OR2_X1 U246bar ( .A1(bbar[13]), .A2(abar[6]), .ZN(ybar[109]);
  AND2_X1 U247 ( .A1(b[12]), .A2(a[6]), .ZN(y[108]) );
  OR2_X1 U247bar ( .A1(bbar[12]), .A2(abar[6]), .ZN(ybar[108]);
  AND2_X1 U248 ( .A1(b[11]), .A2(a[6]), .ZN(y[107]) );
  OR2_X1 U248bar ( .A1(bbar[11]), .A2(abar[6]), .ZN(ybar[107]);
  AND2_X1 U249 ( .A1(b[10]), .A2(a[6]), .ZN(y[106]) );
  OR2_X1 U249bar ( .A1(bbar[10]), .A2(abar[6]), .ZN(ybar[106]);
  AND2_X1 U250 ( .A1(a[6]), .A2(b[9]), .ZN(y[105]) );
  OR2_X1 U250bar ( .A1(abar[6]), .A2(bbar[9]), .ZN(ybar[105]);
  AND2_X1 U251 ( .A1(b[8]), .A2(a[6]), .ZN(y[104]) );
  OR2_X1 U251bar ( .A1(bbar[8]), .A2(abar[6]), .ZN(ybar[104]);
  AND2_X1 U252 ( .A1(b[7]), .A2(a[6]), .ZN(y[103]) );
  OR2_X1 U252bar ( .A1(bbar[7]), .A2(abar[6]), .ZN(ybar[103]);
  AND2_X1 U253 ( .A1(b[6]), .A2(a[6]), .ZN(y[102]) );
  OR2_X1 U253bar ( .A1(bbar[6]), .A2(abar[6]), .ZN(ybar[102]);
  AND2_X1 U254 ( .A1(b[5]), .A2(a[6]), .ZN(y[101]) );
  OR2_X1 U254bar ( .A1(bbar[5]), .A2(abar[6]), .ZN(ybar[101]);
  AND2_X1 U255 ( .A1(b[4]), .A2(a[6]), .ZN(y[100]) );
  OR2_X1 U255bar ( .A1(bbar[4]), .A2(abar[6]), .ZN(ybar[100]);
  AND2_X1 U256 ( .A1(b[0]), .A2(a[0]), .ZN(y[0]) );
  OR2_X1 U256bar ( .A1(bbar[0]), .A2(abar[0]), .ZN(ybar[0]);
endmodule




module decode_1 ( in, out );
  input [7:0] in;
  //input_done

  output [255:0] out;
  //output_done

  wire   [15:0] level1;
  wire   [31:0] level2;
  //wire_done

  CD2_4 cd_l1_1 ( .a(in[1]), .b(in[0]), .y(level1[3:0]) );
  CD2_3 cd_l1_2 ( .a(in[3]), .b(in[2]), .y(level1[7:4]) );
  CD2_2 cd_l1_3 ( .a(in[5]), .b(in[4]), .y(level1[11:8]) );
  CD2_1 cd_l1_4 ( .a(in[7]), .b(in[6]), .y(level1[15:12]) );
  CD4_2 cd_l2_1 ( .a(level1[7:4]), .b(level1[3:0]), .y(level2[15:0]) );
  CD4_1 cd_l2_2 ( .a(level1[15:12]), .b(level1[11:8]), .y(level2[31:16]) );
  CD16_1 cd_l3 ( .a(level2[31:16]), .b(level2[15:0]), .y(out) );
endmodule


module encode_1 ( in, out );
  input [255:0] in;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
  assign inbar[8] = ~in[8];
  assign inbar[9] = ~in[9];
  assign inbar[10] = ~in[10];
  assign inbar[11] = ~in[11];
  assign inbar[12] = ~in[12];
  assign inbar[13] = ~in[13];
  assign inbar[14] = ~in[14];
  assign inbar[15] = ~in[15];
  assign inbar[16] = ~in[16];
  assign inbar[17] = ~in[17];
  assign inbar[18] = ~in[18];
  assign inbar[19] = ~in[19];
  assign inbar[20] = ~in[20];
  assign inbar[21] = ~in[21];
  assign inbar[22] = ~in[22];
  assign inbar[23] = ~in[23];
  assign inbar[24] = ~in[24];
  assign inbar[25] = ~in[25];
  assign inbar[26] = ~in[26];
  assign inbar[27] = ~in[27];
  assign inbar[28] = ~in[28];
  assign inbar[29] = ~in[29];
  assign inbar[30] = ~in[30];
  assign inbar[31] = ~in[31];
  assign inbar[32] = ~in[32];
  assign inbar[33] = ~in[33];
  assign inbar[34] = ~in[34];
  assign inbar[35] = ~in[35];
  assign inbar[36] = ~in[36];
  assign inbar[37] = ~in[37];
  assign inbar[38] = ~in[38];
  assign inbar[39] = ~in[39];
  assign inbar[40] = ~in[40];
  assign inbar[41] = ~in[41];
  assign inbar[42] = ~in[42];
  assign inbar[43] = ~in[43];
  assign inbar[44] = ~in[44];
  assign inbar[45] = ~in[45];
  assign inbar[46] = ~in[46];
  assign inbar[47] = ~in[47];
  assign inbar[48] = ~in[48];
  assign inbar[49] = ~in[49];
  assign inbar[50] = ~in[50];
  assign inbar[51] = ~in[51];
  assign inbar[52] = ~in[52];
  assign inbar[53] = ~in[53];
  assign inbar[54] = ~in[54];
  assign inbar[55] = ~in[55];
  assign inbar[56] = ~in[56];
  assign inbar[57] = ~in[57];
  assign inbar[58] = ~in[58];
  assign inbar[59] = ~in[59];
  assign inbar[60] = ~in[60];
  assign inbar[61] = ~in[61];
  assign inbar[62] = ~in[62];
  assign inbar[63] = ~in[63];
  assign inbar[64] = ~in[64];
  assign inbar[65] = ~in[65];
  assign inbar[66] = ~in[66];
  assign inbar[67] = ~in[67];
  assign inbar[68] = ~in[68];
  assign inbar[69] = ~in[69];
  assign inbar[70] = ~in[70];
  assign inbar[71] = ~in[71];
  assign inbar[72] = ~in[72];
  assign inbar[73] = ~in[73];
  assign inbar[74] = ~in[74];
  assign inbar[75] = ~in[75];
  assign inbar[76] = ~in[76];
  assign inbar[77] = ~in[77];
  assign inbar[78] = ~in[78];
  assign inbar[79] = ~in[79];
  assign inbar[80] = ~in[80];
  assign inbar[81] = ~in[81];
  assign inbar[82] = ~in[82];
  assign inbar[83] = ~in[83];
  assign inbar[84] = ~in[84];
  assign inbar[85] = ~in[85];
  assign inbar[86] = ~in[86];
  assign inbar[87] = ~in[87];
  assign inbar[88] = ~in[88];
  assign inbar[89] = ~in[89];
  assign inbar[90] = ~in[90];
  assign inbar[91] = ~in[91];
  assign inbar[92] = ~in[92];
  assign inbar[93] = ~in[93];
  assign inbar[94] = ~in[94];
  assign inbar[95] = ~in[95];
  assign inbar[96] = ~in[96];
  assign inbar[97] = ~in[97];
  assign inbar[98] = ~in[98];
  assign inbar[99] = ~in[99];
  assign inbar[100] = ~in[100];
  assign inbar[101] = ~in[101];
  assign inbar[102] = ~in[102];
  assign inbar[103] = ~in[103];
  assign inbar[104] = ~in[104];
  assign inbar[105] = ~in[105];
  assign inbar[106] = ~in[106];
  assign inbar[107] = ~in[107];
  assign inbar[108] = ~in[108];
  assign inbar[109] = ~in[109];
  assign inbar[110] = ~in[110];
  assign inbar[111] = ~in[111];
  assign inbar[112] = ~in[112];
  assign inbar[113] = ~in[113];
  assign inbar[114] = ~in[114];
  assign inbar[115] = ~in[115];
  assign inbar[116] = ~in[116];
  assign inbar[117] = ~in[117];
  assign inbar[118] = ~in[118];
  assign inbar[119] = ~in[119];
  assign inbar[120] = ~in[120];
  assign inbar[121] = ~in[121];
  assign inbar[122] = ~in[122];
  assign inbar[123] = ~in[123];
  assign inbar[124] = ~in[124];
  assign inbar[125] = ~in[125];
  assign inbar[126] = ~in[126];
  assign inbar[127] = ~in[127];
  assign inbar[128] = ~in[128];
  assign inbar[129] = ~in[129];
  assign inbar[130] = ~in[130];
  assign inbar[131] = ~in[131];
  assign inbar[132] = ~in[132];
  assign inbar[133] = ~in[133];
  assign inbar[134] = ~in[134];
  assign inbar[135] = ~in[135];
  assign inbar[136] = ~in[136];
  assign inbar[137] = ~in[137];
  assign inbar[138] = ~in[138];
  assign inbar[139] = ~in[139];
  assign inbar[140] = ~in[140];
  assign inbar[141] = ~in[141];
  assign inbar[142] = ~in[142];
  assign inbar[143] = ~in[143];
  assign inbar[144] = ~in[144];
  assign inbar[145] = ~in[145];
  assign inbar[146] = ~in[146];
  assign inbar[147] = ~in[147];
  assign inbar[148] = ~in[148];
  assign inbar[149] = ~in[149];
  assign inbar[150] = ~in[150];
  assign inbar[151] = ~in[151];
  assign inbar[152] = ~in[152];
  assign inbar[153] = ~in[153];
  assign inbar[154] = ~in[154];
  assign inbar[155] = ~in[155];
  assign inbar[156] = ~in[156];
  assign inbar[157] = ~in[157];
  assign inbar[158] = ~in[158];
  assign inbar[159] = ~in[159];
  assign inbar[160] = ~in[160];
  assign inbar[161] = ~in[161];
  assign inbar[162] = ~in[162];
  assign inbar[163] = ~in[163];
  assign inbar[164] = ~in[164];
  assign inbar[165] = ~in[165];
  assign inbar[166] = ~in[166];
  assign inbar[167] = ~in[167];
  assign inbar[168] = ~in[168];
  assign inbar[169] = ~in[169];
  assign inbar[170] = ~in[170];
  assign inbar[171] = ~in[171];
  assign inbar[172] = ~in[172];
  assign inbar[173] = ~in[173];
  assign inbar[174] = ~in[174];
  assign inbar[175] = ~in[175];
  assign inbar[176] = ~in[176];
  assign inbar[177] = ~in[177];
  assign inbar[178] = ~in[178];
  assign inbar[179] = ~in[179];
  assign inbar[180] = ~in[180];
  assign inbar[181] = ~in[181];
  assign inbar[182] = ~in[182];
  assign inbar[183] = ~in[183];
  assign inbar[184] = ~in[184];
  assign inbar[185] = ~in[185];
  assign inbar[186] = ~in[186];
  assign inbar[187] = ~in[187];
  assign inbar[188] = ~in[188];
  assign inbar[189] = ~in[189];
  assign inbar[190] = ~in[190];
  assign inbar[191] = ~in[191];
  assign inbar[192] = ~in[192];
  assign inbar[193] = ~in[193];
  assign inbar[194] = ~in[194];
  assign inbar[195] = ~in[195];
  assign inbar[196] = ~in[196];
  assign inbar[197] = ~in[197];
  assign inbar[198] = ~in[198];
  assign inbar[199] = ~in[199];
  assign inbar[200] = ~in[200];
  assign inbar[201] = ~in[201];
  assign inbar[202] = ~in[202];
  assign inbar[203] = ~in[203];
  assign inbar[204] = ~in[204];
  assign inbar[205] = ~in[205];
  assign inbar[206] = ~in[206];
  assign inbar[207] = ~in[207];
  assign inbar[208] = ~in[208];
  assign inbar[209] = ~in[209];
  assign inbar[210] = ~in[210];
  assign inbar[211] = ~in[211];
  assign inbar[212] = ~in[212];
  assign inbar[213] = ~in[213];
  assign inbar[214] = ~in[214];
  assign inbar[215] = ~in[215];
  assign inbar[216] = ~in[216];
  assign inbar[217] = ~in[217];
  assign inbar[218] = ~in[218];
  assign inbar[219] = ~in[219];
  assign inbar[220] = ~in[220];
  assign inbar[221] = ~in[221];
  assign inbar[222] = ~in[222];
  assign inbar[223] = ~in[223];
  assign inbar[224] = ~in[224];
  assign inbar[225] = ~in[225];
  assign inbar[226] = ~in[226];
  assign inbar[227] = ~in[227];
  assign inbar[228] = ~in[228];
  assign inbar[229] = ~in[229];
  assign inbar[230] = ~in[230];
  assign inbar[231] = ~in[231];
  assign inbar[232] = ~in[232];
  assign inbar[233] = ~in[233];
  assign inbar[234] = ~in[234];
  assign inbar[235] = ~in[235];
  assign inbar[236] = ~in[236];
  assign inbar[237] = ~in[237];
  assign inbar[238] = ~in[238];
  assign inbar[239] = ~in[239];
  assign inbar[240] = ~in[240];
  assign inbar[241] = ~in[241];
  assign inbar[242] = ~in[242];
  assign inbar[243] = ~in[243];
  assign inbar[244] = ~in[244];
  assign inbar[245] = ~in[245];
  assign inbar[246] = ~in[246];
  assign inbar[247] = ~in[247];
  assign inbar[248] = ~in[248];
  assign inbar[249] = ~in[249];
  assign inbar[250] = ~in[250];
  assign inbar[251] = ~in[251];
  assign inbar[252] = ~in[252];
  assign inbar[253] = ~in[253];
  assign inbar[254] = ~in[254];
  assign inbar[255] = ~in[255];
  //input_done

  output [7:0] out;
  reg [7:0] outbar;
  //output_done

  wire   in_81, in_80, in_79, in_78, in_77, in_76, in_75, in_74, in_73, in_72,
         in_71, in_70, in_69, in_68, in_67, in_66, in_65, in_64, in_63, in_62,
         in_61, in_60, in_59, in_58, in_57, in_56, in_55, in_54, in_53, in_52,
         in_51, in_50, in_49, in_48, in_47, in_46, in_45, in_44, in_43, in_42,
         in_41, in_40, in_39, in_38, in_37, in_36, in_35, in_34, in_33, in_32,
         in_31, in_30, in_29, in_28, in_27, in_26, in_25, in_24, in_23, in_22,
         in_21, in_20, in_19, in_18, in_17, in_16, in_15, in_14, in_13, in_12,
         in_11, in_10, in_9, in_8, in_7, in_6, in_5, in_4, in_3, in_2, in_1,
         in_0, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972;
  wire in_81bar, in_80bar, in_79bar, in_78bar, in_77bar, in_76bar, in_75bar, in_74bar, in_73bar, in_72bar, in_71bar, in_70bar, in_69bar, in_68bar, in_67bar, in_66bar, in_65bar, in_64bar, in_63bar, in_62bar, in_61bar, in_60bar, in_59bar, in_58bar, in_57bar, in_56bar, in_55bar, in_54bar, in_53bar, in_52bar, in_51bar, in_50bar, in_49bar, in_48bar, in_47bar, in_46bar, in_45bar, in_44bar, in_43bar, in_42bar, in_41bar, in_40bar, in_39bar, in_38bar, in_37bar, in_36bar, in_35bar, in_34bar, in_33bar, in_32bar, in_31bar, in_30bar, in_29bar, in_28bar, in_27bar, in_26bar, in_25bar, in_24bar, in_23bar, in_22bar, in_21bar, in_20bar, in_19bar, in_18bar, in_17bar, in_16bar, in_15bar, in_14bar, in_13bar, in_12bar, in_11bar, in_10bar, in_9bar, in_8bar, in_7bar, in_6bar, in_5bar, in_4bar, in_3bar, in_2bar, in_1bar, in_0bar, n487bar, n488bar, n489bar, n490bar, n491bar, n492bar, n493bar, n494bar, n495bar, n496bar, n497bar, n498bar, n499bar, n500bar, n501bar, n502bar, n503bar, n504bar, n505bar, n506bar, n507bar, n508bar, n509bar, n510bar, n511bar, n512bar, n513bar, n514bar, n515bar, n516bar, n517bar, n518bar, n519bar, n520bar, n521bar, n522bar, n523bar, n524bar, n525bar, n526bar, n527bar, n528bar, n529bar, n530bar, n531bar, n532bar, n533bar, n534bar, n535bar, n536bar, n537bar, n538bar, n539bar, n540bar, n541bar, n542bar, n543bar, n544bar, n545bar, n546bar, n547bar, n548bar, n549bar, n550bar, n551bar, n552bar, n553bar, n554bar, n555bar, n556bar, n557bar, n558bar, n559bar, n560bar, n561bar, n562bar, n563bar, n564bar, n565bar, n566bar, n567bar, n568bar, n569bar, n570bar, n571bar, n572bar, n573bar, n574bar, n575bar, n576bar, n577bar, n578bar, n579bar, n580bar, n581bar, n582bar, n583bar, n584bar, n585bar, n586bar, n587bar, n588bar, n589bar, n590bar, n591bar, n592bar, n593bar, n594bar, n595bar, n596bar, n597bar, n598bar, n599bar, n600bar, n601bar, n602bar, n603bar, n604bar, n605bar, n606bar, n607bar, n608bar, n609bar, n610bar, n611bar, n612bar, n613bar, n614bar, n615bar, n616bar, n617bar, n618bar, n619bar, n620bar, n621bar, n622bar, n623bar, n624bar, n625bar, n626bar, n627bar, n628bar, n629bar, n630bar, n631bar, n632bar, n633bar, n634bar, n635bar, n636bar, n637bar, n638bar, n639bar, n640bar, n641bar, n642bar, n643bar, n644bar, n645bar, n646bar, n647bar, n648bar, n649bar, n650bar, n651bar, n652bar, n653bar, n654bar, n655bar, n656bar, n657bar, n658bar, n659bar, n660bar, n661bar, n662bar, n663bar, n664bar, n665bar, n666bar, n667bar, n668bar, n669bar, n670bar, n671bar, n672bar, n673bar, n674bar, n675bar, n676bar, n677bar, n678bar, n679bar, n680bar, n681bar, n682bar, n683bar, n684bar, n685bar, n686bar, n687bar, n688bar, n689bar, n690bar, n691bar, n692bar, n693bar, n694bar, n695bar, n696bar, n697bar, n698bar, n699bar, n700bar, n701bar, n702bar, n703bar, n704bar, n705bar, n706bar, n707bar, n708bar, n709bar, n710bar, n711bar, n712bar, n713bar, n714bar, n715bar, n716bar, n717bar, n718bar, n719bar, n720bar, n721bar, n722bar, n723bar, n724bar, n725bar, n726bar, n727bar, n728bar, n729bar, n730bar, n731bar, n732bar, n733bar, n734bar, n735bar, n736bar, n737bar, n738bar, n739bar, n740bar, n741bar, n742bar, n743bar, n744bar, n745bar, n746bar, n747bar, n748bar, n749bar, n750bar, n751bar, n752bar, n753bar, n754bar, n755bar, n756bar, n757bar, n758bar, n759bar, n760bar, n761bar, n762bar, n763bar, n764bar, n765bar, n766bar, n767bar, n768bar, n769bar, n770bar, n771bar, n772bar, n773bar, n774bar, n775bar, n776bar, n777bar, n778bar, n779bar, n780bar, n781bar, n782bar, n783bar, n784bar, n785bar, n786bar, n787bar, n788bar, n789bar, n790bar, n791bar, n792bar, n793bar, n794bar, n795bar, n796bar, n797bar, n798bar, n799bar, n800bar, n801bar, n802bar, n803bar, n804bar, n805bar, n806bar, n807bar, n808bar, n809bar, n810bar, n811bar, n812bar, n813bar, n814bar, n815bar, n816bar, n817bar, n818bar, n819bar, n820bar, n821bar, n822bar, n823bar, n824bar, n825bar, n826bar, n827bar, n828bar, n829bar, n830bar, n831bar, n832bar, n833bar, n834bar, n835bar, n836bar, n837bar, n838bar, n839bar, n840bar, n841bar, n842bar, n843bar, n844bar, n845bar, n846bar, n847bar, n848bar, n849bar, n850bar, n851bar, n852bar, n853bar, n854bar, n855bar, n856bar, n857bar, n858bar, n859bar, n860bar, n861bar, n862bar, n863bar, n864bar, n865bar, n866bar, n867bar, n868bar, n869bar, n870bar, n871bar, n872bar, n873bar, n874bar, n875bar, n876bar, n877bar, n878bar, n879bar, n880bar, n881bar, n882bar, n883bar, n884bar, n885bar, n886bar, n887bar, n888bar, n889bar, n890bar, n891bar, n892bar, n893bar, n894bar, n895bar, n896bar, n897bar, n898bar, n899bar, n900bar, n901bar, n902bar, n903bar, n904bar, n905bar, n906bar, n907bar, n908bar, n909bar, n910bar, n911bar, n912bar, n913bar, n914bar, n915bar, n916bar, n917bar, n918bar, n919bar, n920bar, n921bar, n922bar, n923bar, n924bar, n925bar, n926bar, n927bar, n928bar, n929bar, n930bar, n931bar, n932bar, n933bar, n934bar, n935bar, n936bar, n937bar, n938bar, n939bar, n940bar, n941bar, n942bar, n943bar, n944bar, n945bar, n946bar, n947bar, n948bar, n949bar, n950bar, n951bar, n952bar, n953bar, n954bar, n955bar, n956bar, n957bar, n958bar, n959bar, n960bar, n961bar, n962bar, n963bar, n964bar, n965bar, n966bar, n967bar, n968bar, n969bar, n970bar, n971bar, n972bar;
  //wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];

  OR2_X1 U1 ( .A1(n972), .A2(n971), .ZN(out[7]) );
  AND2_X1 U1bar ( .A1(n972bar), .A2(n971bar), .ZN(outbar[7]);
  OR2_X1 U2 ( .A1(n970), .A2(n969), .ZN(n971) );
  AND2_X1 U2bar ( .A1(n970bar), .A2(n969bar), .ZN(n971bar);
  OR2_X1 U3 ( .A1(n968), .A2(n967), .ZN(n969) );
  AND2_X1 U3bar ( .A1(n968bar), .A2(n967bar), .ZN(n969bar);
  OR2_X1 U4 ( .A1(n966), .A2(n965), .ZN(n967) );
  AND2_X1 U4bar ( .A1(n966bar), .A2(n965bar), .ZN(n967bar);
  OR2_X1 U5 ( .A1(n964), .A2(n963), .ZN(n968) );
  AND2_X1 U5bar ( .A1(n964bar), .A2(n963bar), .ZN(n968bar);
  OR2_X1 U6 ( .A1(in[116]), .A2(n962), .ZN(n963) );
  AND2_X1 U6bar ( .A1(inbar[116]), .A2(n962bar), .ZN(n963bar);
  OR2_X1 U7 ( .A1(n961), .A2(n960), .ZN(n970) );
  AND2_X1 U7bar ( .A1(n961bar), .A2(n960bar), .ZN(n970bar);
  OR2_X1 U8 ( .A1(in[150]), .A2(in[127]), .ZN(n960) );
  AND2_X1 U8bar ( .A1(inbar[150]), .A2(inbar[127]), .ZN(n960bar);
  OR2_X1 U9 ( .A1(in[160]), .A2(n959), .ZN(n961) );
  AND2_X1 U9bar ( .A1(inbar[160]), .A2(n959bar), .ZN(n961bar);
  OR2_X1 U10 ( .A1(in[252]), .A2(in[168]), .ZN(n959) );
  AND2_X1 U10bar ( .A1(inbar[252]), .A2(inbar[168]), .ZN(n959bar);
  OR2_X1 U11 ( .A1(n958), .A2(n957), .ZN(n972) );
  AND2_X1 U11bar ( .A1(n958bar), .A2(n957bar), .ZN(n972bar);
  OR2_X1 U12 ( .A1(n956), .A2(n955), .ZN(n957) );
  AND2_X1 U12bar ( .A1(n956bar), .A2(n955bar), .ZN(n957bar);
  OR2_X1 U13 ( .A1(in_17), .A2(in[96]), .ZN(n955) );
  AND2_X1 U13bar ( .A1(in_17bar), .A2(inbar[96]), .ZN(n955bar);
  OR2_X1 U14 ( .A1(in_23), .A2(n954), .ZN(n956) );
  AND2_X1 U14bar ( .A1(in_23bar), .A2(n954bar), .ZN(n956bar);
  OR2_X1 U15 ( .A1(in_31), .A2(in_26), .ZN(n954) );
  AND2_X1 U15bar ( .A1(in_31bar), .A2(in_26bar), .ZN(n954bar);
  OR2_X1 U16 ( .A1(n953), .A2(n952), .ZN(n958) );
  AND2_X1 U16bar ( .A1(n953bar), .A2(n952bar), .ZN(n958bar);
  OR2_X1 U17 ( .A1(in_58), .A2(in_4), .ZN(n952) );
  AND2_X1 U17bar ( .A1(in_58bar), .A2(in_4bar), .ZN(n952bar);
  OR2_X1 U18 ( .A1(in_59), .A2(n951), .ZN(n953) );
  AND2_X1 U18bar ( .A1(in_59bar), .A2(n951bar), .ZN(n953bar);
  OR2_X1 U19 ( .A1(in_71), .A2(in_62), .ZN(n951) );
  AND2_X1 U19bar ( .A1(in_71bar), .A2(in_62bar), .ZN(n951bar);
  OR2_X1 U20 ( .A1(n950), .A2(n949), .ZN(out[6]) );
  AND2_X1 U20bar ( .A1(n950bar), .A2(n949bar), .ZN(outbar[6]);
  OR2_X1 U21 ( .A1(n948), .A2(n947), .ZN(n949) );
  AND2_X1 U21bar ( .A1(n948bar), .A2(n947bar), .ZN(n949bar);
  OR2_X1 U22 ( .A1(n946), .A2(n945), .ZN(n947) );
  AND2_X1 U22bar ( .A1(n946bar), .A2(n945bar), .ZN(n947bar);
  OR2_X1 U23 ( .A1(n944), .A2(n943), .ZN(n945) );
  AND2_X1 U23bar ( .A1(n944bar), .A2(n943bar), .ZN(n945bar);
  OR2_X1 U24 ( .A1(n942), .A2(n941), .ZN(n946) );
  AND2_X1 U24bar ( .A1(n942bar), .A2(n941bar), .ZN(n946bar);
  OR2_X1 U25 ( .A1(in[101]), .A2(n940), .ZN(n941) );
  AND2_X1 U25bar ( .A1(inbar[101]), .A2(n940bar), .ZN(n941bar);
  OR2_X1 U26 ( .A1(n939), .A2(n938), .ZN(n948) );
  AND2_X1 U26bar ( .A1(n939bar), .A2(n938bar), .ZN(n948bar);
  OR2_X1 U27 ( .A1(in[114]), .A2(in[104]), .ZN(n938) );
  AND2_X1 U27bar ( .A1(inbar[114]), .A2(inbar[104]), .ZN(n938bar);
  OR2_X1 U28 ( .A1(in[128]), .A2(n937), .ZN(n939) );
  AND2_X1 U28bar ( .A1(inbar[128]), .A2(n937bar), .ZN(n939bar);
  OR2_X1 U29 ( .A1(in[136]), .A2(in[134]), .ZN(n937) );
  AND2_X1 U29bar ( .A1(inbar[136]), .A2(inbar[134]), .ZN(n937bar);
  OR2_X1 U30 ( .A1(n936), .A2(n935), .ZN(n950) );
  AND2_X1 U30bar ( .A1(n936bar), .A2(n935bar), .ZN(n950bar);
  OR2_X1 U31 ( .A1(n934), .A2(n933), .ZN(n935) );
  AND2_X1 U31bar ( .A1(n934bar), .A2(n933bar), .ZN(n935bar);
  OR2_X1 U32 ( .A1(in[177]), .A2(in[164]), .ZN(n933) );
  AND2_X1 U32bar ( .A1(inbar[177]), .A2(inbar[164]), .ZN(n933bar);
  OR2_X1 U33 ( .A1(in[212]), .A2(n932), .ZN(n934) );
  AND2_X1 U33bar ( .A1(inbar[212]), .A2(n932bar), .ZN(n934bar);
  OR2_X1 U34 ( .A1(in[248]), .A2(in[221]), .ZN(n932) );
  AND2_X1 U34bar ( .A1(inbar[248]), .A2(inbar[221]), .ZN(n932bar);
  OR2_X1 U35 ( .A1(n931), .A2(n930), .ZN(n936) );
  AND2_X1 U35bar ( .A1(n931bar), .A2(n930bar), .ZN(n936bar);
  OR2_X1 U36 ( .A1(in_18), .A2(in[93]), .ZN(n930) );
  AND2_X1 U36bar ( .A1(in_18bar), .A2(inbar[93]), .ZN(n930bar);
  OR2_X1 U37 ( .A1(in_31), .A2(n929), .ZN(n931) );
  AND2_X1 U37bar ( .A1(in_31bar), .A2(n929bar), .ZN(n931bar);
  OR2_X1 U38 ( .A1(in_7), .A2(in_39), .ZN(n929) );
  AND2_X1 U38bar ( .A1(in_7bar), .A2(in_39bar), .ZN(n929bar);
  OR2_X1 U39 ( .A1(n928), .A2(n927), .ZN(out[5]) );
  AND2_X1 U39bar ( .A1(n928bar), .A2(n927bar), .ZN(outbar[5]);
  OR2_X1 U40 ( .A1(n926), .A2(n925), .ZN(n927) );
  AND2_X1 U40bar ( .A1(n926bar), .A2(n925bar), .ZN(n927bar);
  OR2_X1 U41 ( .A1(n924), .A2(n923), .ZN(n925) );
  AND2_X1 U41bar ( .A1(n924bar), .A2(n923bar), .ZN(n925bar);
  OR2_X1 U42 ( .A1(n922), .A2(n921), .ZN(n923) );
  AND2_X1 U42bar ( .A1(n922bar), .A2(n921bar), .ZN(n923bar);
  OR2_X1 U43 ( .A1(n940), .A2(n920), .ZN(n924) );
  AND2_X1 U43bar ( .A1(n940bar), .A2(n920bar), .ZN(n924bar);
  OR2_X1 U44 ( .A1(in[111]), .A2(n919), .ZN(n920) );
  AND2_X1 U44bar ( .A1(inbar[111]), .A2(n919bar), .ZN(n920bar);
  OR2_X1 U45 ( .A1(n918), .A2(n917), .ZN(n940) );
  AND2_X1 U45bar ( .A1(n918bar), .A2(n917bar), .ZN(n940bar);
  OR2_X1 U46 ( .A1(n916), .A2(n915), .ZN(n917) );
  AND2_X1 U46bar ( .A1(n916bar), .A2(n915bar), .ZN(n917bar);
  OR2_X1 U47 ( .A1(n914), .A2(n913), .ZN(n915) );
  AND2_X1 U47bar ( .A1(n914bar), .A2(n913bar), .ZN(n915bar);
  OR2_X1 U48 ( .A1(in[140]), .A2(in[131]), .ZN(n913) );
  AND2_X1 U48bar ( .A1(inbar[140]), .A2(inbar[131]), .ZN(n913bar);
  OR2_X1 U49 ( .A1(in[160]), .A2(in[144]), .ZN(n914) );
  AND2_X1 U49bar ( .A1(inbar[160]), .A2(inbar[144]), .ZN(n914bar);
  OR2_X1 U50 ( .A1(n912), .A2(n911), .ZN(n916) );
  AND2_X1 U50bar ( .A1(n912bar), .A2(n911bar), .ZN(n916bar);
  OR2_X1 U51 ( .A1(in[179]), .A2(in[174]), .ZN(n911) );
  AND2_X1 U51bar ( .A1(inbar[179]), .A2(inbar[174]), .ZN(n911bar);
  OR2_X1 U52 ( .A1(in[188]), .A2(in[184]), .ZN(n912) );
  AND2_X1 U52bar ( .A1(inbar[188]), .A2(inbar[184]), .ZN(n912bar);
  OR2_X1 U53 ( .A1(n910), .A2(n909), .ZN(n918) );
  AND2_X1 U53bar ( .A1(n910bar), .A2(n909bar), .ZN(n918bar);
  OR2_X1 U54 ( .A1(n908), .A2(n907), .ZN(n909) );
  AND2_X1 U54bar ( .A1(n908bar), .A2(n907bar), .ZN(n909bar);
  OR2_X1 U55 ( .A1(in[216]), .A2(in[200]), .ZN(n907) );
  AND2_X1 U55bar ( .A1(inbar[216]), .A2(inbar[200]), .ZN(n907bar);
  OR2_X1 U56 ( .A1(in[228]), .A2(in[224]), .ZN(n908) );
  AND2_X1 U56bar ( .A1(inbar[228]), .A2(inbar[224]), .ZN(n908bar);
  OR2_X1 U57 ( .A1(n906), .A2(n905), .ZN(n910) );
  AND2_X1 U57bar ( .A1(n906bar), .A2(n905bar), .ZN(n910bar);
  OR2_X1 U58 ( .A1(in[247]), .A2(in[235]), .ZN(n905) );
  AND2_X1 U58bar ( .A1(inbar[247]), .A2(inbar[235]), .ZN(n905bar);
  OR2_X1 U59 ( .A1(in_42), .A2(in[83]), .ZN(n906) );
  AND2_X1 U59bar ( .A1(in_42bar), .A2(inbar[83]), .ZN(n906bar);
  OR2_X1 U60 ( .A1(n904), .A2(n903), .ZN(n926) );
  AND2_X1 U60bar ( .A1(n904bar), .A2(n903bar), .ZN(n926bar);
  OR2_X1 U61 ( .A1(in[166]), .A2(in[123]), .ZN(n903) );
  AND2_X1 U61bar ( .A1(inbar[166]), .A2(inbar[123]), .ZN(n903bar);
  OR2_X1 U62 ( .A1(in[170]), .A2(n902), .ZN(n904) );
  AND2_X1 U62bar ( .A1(inbar[170]), .A2(n902bar), .ZN(n904bar);
  OR2_X1 U63 ( .A1(in[194]), .A2(in[183]), .ZN(n902) );
  AND2_X1 U63bar ( .A1(inbar[194]), .A2(inbar[183]), .ZN(n902bar);
  OR2_X1 U64 ( .A1(n901), .A2(n900), .ZN(n928) );
  AND2_X1 U64bar ( .A1(n901bar), .A2(n900bar), .ZN(n928bar);
  OR2_X1 U65 ( .A1(n899), .A2(n898), .ZN(n900) );
  AND2_X1 U65bar ( .A1(n899bar), .A2(n898bar), .ZN(n900bar);
  OR2_X1 U66 ( .A1(in[241]), .A2(in[238]), .ZN(n898) );
  AND2_X1 U66bar ( .A1(inbar[241]), .A2(inbar[238]), .ZN(n898bar);
  OR2_X1 U67 ( .A1(in[250]), .A2(n897), .ZN(n899) );
  AND2_X1 U67bar ( .A1(inbar[250]), .A2(n897bar), .ZN(n899bar);
  OR2_X1 U68 ( .A1(in_24), .A2(in[84]), .ZN(n897) );
  AND2_X1 U68bar ( .A1(in_24bar), .A2(inbar[84]), .ZN(n897bar);
  OR2_X1 U69 ( .A1(n896), .A2(n895), .ZN(n901) );
  AND2_X1 U69bar ( .A1(n896bar), .A2(n895bar), .ZN(n901bar);
  OR2_X1 U70 ( .A1(in_41), .A2(in_29), .ZN(n895) );
  AND2_X1 U70bar ( .A1(in_41bar), .A2(in_29bar), .ZN(n895bar);
  OR2_X1 U71 ( .A1(in_66), .A2(n894), .ZN(n896) );
  AND2_X1 U71bar ( .A1(in_66bar), .A2(n894bar), .ZN(n896bar);
  OR2_X1 U72 ( .A1(in_76), .A2(in_71), .ZN(n894) );
  AND2_X1 U72bar ( .A1(in_76bar), .A2(in_71bar), .ZN(n894bar);
  OR2_X1 U73 ( .A1(n893), .A2(n892), .ZN(out[4]) );
  AND2_X1 U73bar ( .A1(n893bar), .A2(n892bar), .ZN(outbar[4]);
  OR2_X1 U74 ( .A1(n891), .A2(n890), .ZN(n892) );
  AND2_X1 U74bar ( .A1(n891bar), .A2(n890bar), .ZN(n892bar);
  OR2_X1 U75 ( .A1(n889), .A2(n888), .ZN(n890) );
  AND2_X1 U75bar ( .A1(n889bar), .A2(n888bar), .ZN(n890bar);
  OR2_X1 U76 ( .A1(n922), .A2(n887), .ZN(n888) );
  AND2_X1 U76bar ( .A1(n922bar), .A2(n887bar), .ZN(n888bar);
  OR2_X1 U77 ( .A1(n886), .A2(n885), .ZN(n922) );
  AND2_X1 U77bar ( .A1(n886bar), .A2(n885bar), .ZN(n922bar);
  OR2_X1 U78 ( .A1(n884), .A2(n883), .ZN(n885) );
  AND2_X1 U78bar ( .A1(n884bar), .A2(n883bar), .ZN(n885bar);
  OR2_X1 U79 ( .A1(n882), .A2(n881), .ZN(n883) );
  AND2_X1 U79bar ( .A1(n882bar), .A2(n881bar), .ZN(n883bar);
  OR2_X1 U80 ( .A1(in[118]), .A2(in[109]), .ZN(n881) );
  AND2_X1 U80bar ( .A1(inbar[118]), .A2(inbar[109]), .ZN(n881bar);
  OR2_X1 U81 ( .A1(in[139]), .A2(in[120]), .ZN(n882) );
  AND2_X1 U81bar ( .A1(inbar[139]), .A2(inbar[120]), .ZN(n882bar);
  OR2_X1 U82 ( .A1(n880), .A2(n879), .ZN(n884) );
  AND2_X1 U82bar ( .A1(n880bar), .A2(n879bar), .ZN(n884bar);
  OR2_X1 U83 ( .A1(in[198]), .A2(in[154]), .ZN(n879) );
  AND2_X1 U83bar ( .A1(inbar[198]), .A2(inbar[154]), .ZN(n879bar);
  OR2_X1 U84 ( .A1(in[210]), .A2(in[205]), .ZN(n880) );
  AND2_X1 U84bar ( .A1(inbar[210]), .A2(inbar[205]), .ZN(n880bar);
  OR2_X1 U85 ( .A1(n878), .A2(n877), .ZN(n886) );
  AND2_X1 U85bar ( .A1(n878bar), .A2(n877bar), .ZN(n886bar);
  OR2_X1 U86 ( .A1(n876), .A2(n875), .ZN(n877) );
  AND2_X1 U86bar ( .A1(n876bar), .A2(n875bar), .ZN(n877bar);
  OR2_X1 U87 ( .A1(in[219]), .A2(in[217]), .ZN(n875) );
  AND2_X1 U87bar ( .A1(inbar[219]), .A2(inbar[217]), .ZN(n875bar);
  OR2_X1 U88 ( .A1(in[86]), .A2(in[252]), .ZN(n876) );
  AND2_X1 U88bar ( .A1(inbar[86]), .A2(inbar[252]), .ZN(n876bar);
  OR2_X1 U89 ( .A1(n874), .A2(n873), .ZN(n878) );
  AND2_X1 U89bar ( .A1(n874bar), .A2(n873bar), .ZN(n878bar);
  OR2_X1 U90 ( .A1(in_40), .A2(in[91]), .ZN(n873) );
  AND2_X1 U90bar ( .A1(in_40bar), .A2(inbar[91]), .ZN(n873bar);
  OR2_X1 U91 ( .A1(in_8), .A2(in_46), .ZN(n874) );
  AND2_X1 U91bar ( .A1(in_8bar), .A2(in_46bar), .ZN(n874bar);
  OR2_X1 U92 ( .A1(n872), .A2(n871), .ZN(n889) );
  AND2_X1 U92bar ( .A1(n872bar), .A2(n871bar), .ZN(n889bar);
  OR2_X1 U93 ( .A1(in[117]), .A2(n943), .ZN(n871) );
  AND2_X1 U93bar ( .A1(inbar[117]), .A2(n943bar), .ZN(n871bar);
  OR2_X1 U94 ( .A1(n870), .A2(n869), .ZN(n943) );
  AND2_X1 U94bar ( .A1(n870bar), .A2(n869bar), .ZN(n943bar);
  OR2_X1 U95 ( .A1(n868), .A2(n867), .ZN(n869) );
  AND2_X1 U95bar ( .A1(n868bar), .A2(n867bar), .ZN(n869bar);
  OR2_X1 U96 ( .A1(n866), .A2(n865), .ZN(n867) );
  AND2_X1 U96bar ( .A1(n866bar), .A2(n865bar), .ZN(n867bar);
  OR2_X1 U97 ( .A1(n864), .A2(n863), .ZN(n865) );
  AND2_X1 U97bar ( .A1(n864bar), .A2(n863bar), .ZN(n865bar);
  OR2_X1 U98 ( .A1(in[108]), .A2(n919), .ZN(n866) );
  AND2_X1 U98bar ( .A1(inbar[108]), .A2(n919bar), .ZN(n866bar);
  OR2_X1 U99 ( .A1(n862), .A2(n861), .ZN(n919) );
  AND2_X1 U99bar ( .A1(n862bar), .A2(n861bar), .ZN(n919bar);
  OR2_X1 U100 ( .A1(n860), .A2(n859), .ZN(n861) );
  AND2_X1 U100bar ( .A1(n860bar), .A2(n859bar), .ZN(n861bar);
  OR2_X1 U101 ( .A1(n858), .A2(n857), .ZN(n859) );
  AND2_X1 U101bar ( .A1(n858bar), .A2(n857bar), .ZN(n859bar);
  OR2_X1 U102 ( .A1(in[119]), .A2(in[105]), .ZN(n857) );
  AND2_X1 U102bar ( .A1(inbar[119]), .A2(inbar[105]), .ZN(n857bar);
  OR2_X1 U103 ( .A1(in[186]), .A2(in[175]), .ZN(n858) );
  AND2_X1 U103bar ( .A1(inbar[186]), .A2(inbar[175]), .ZN(n858bar);
  OR2_X1 U104 ( .A1(n856), .A2(n855), .ZN(n860) );
  AND2_X1 U104bar ( .A1(n856bar), .A2(n855bar), .ZN(n860bar);
  OR2_X1 U105 ( .A1(in[202]), .A2(in[193]), .ZN(n855) );
  AND2_X1 U105bar ( .A1(inbar[202]), .A2(inbar[193]), .ZN(n855bar);
  OR2_X1 U106 ( .A1(in[225]), .A2(in[208]), .ZN(n856) );
  AND2_X1 U106bar ( .A1(inbar[225]), .A2(inbar[208]), .ZN(n856bar);
  OR2_X1 U107 ( .A1(n854), .A2(n853), .ZN(n862) );
  AND2_X1 U107bar ( .A1(n854bar), .A2(n853bar), .ZN(n862bar);
  OR2_X1 U108 ( .A1(n852), .A2(n851), .ZN(n853) );
  AND2_X1 U108bar ( .A1(n852bar), .A2(n851bar), .ZN(n853bar);
  OR2_X1 U109 ( .A1(in_1), .A2(in[85]), .ZN(n851) );
  AND2_X1 U109bar ( .A1(in_1bar), .A2(inbar[85]), .ZN(n851bar);
  OR2_X1 U110 ( .A1(in_23), .A2(in_19), .ZN(n852) );
  AND2_X1 U110bar ( .A1(in_23bar), .A2(in_19bar), .ZN(n852bar);
  OR2_X1 U111 ( .A1(n850), .A2(n849), .ZN(n854) );
  AND2_X1 U111bar ( .A1(n850bar), .A2(n849bar), .ZN(n854bar);
  OR2_X1 U112 ( .A1(in_43), .A2(in_33), .ZN(n849) );
  AND2_X1 U112bar ( .A1(in_43bar), .A2(in_33bar), .ZN(n849bar);
  OR2_X1 U113 ( .A1(in_63), .A2(in_44), .ZN(n850) );
  AND2_X1 U113bar ( .A1(in_63bar), .A2(in_44bar), .ZN(n850bar);
  OR2_X1 U114 ( .A1(n848), .A2(n847), .ZN(n868) );
  AND2_X1 U114bar ( .A1(n848bar), .A2(n847bar), .ZN(n868bar);
  OR2_X1 U115 ( .A1(in[141]), .A2(in[112]), .ZN(n847) );
  AND2_X1 U115bar ( .A1(inbar[141]), .A2(inbar[112]), .ZN(n847bar);
  OR2_X1 U116 ( .A1(in[147]), .A2(n846), .ZN(n848) );
  AND2_X1 U116bar ( .A1(inbar[147]), .A2(n846bar), .ZN(n848bar);
  OR2_X1 U117 ( .A1(in[181]), .A2(in[167]), .ZN(n846) );
  AND2_X1 U117bar ( .A1(inbar[181]), .A2(inbar[167]), .ZN(n846bar);
  OR2_X1 U118 ( .A1(n845), .A2(n844), .ZN(n870) );
  AND2_X1 U118bar ( .A1(n845bar), .A2(n844bar), .ZN(n870bar);
  OR2_X1 U119 ( .A1(n843), .A2(n842), .ZN(n844) );
  AND2_X1 U119bar ( .A1(n843bar), .A2(n842bar), .ZN(n844bar);
  OR2_X1 U120 ( .A1(in[229]), .A2(in[201]), .ZN(n842) );
  AND2_X1 U120bar ( .A1(inbar[229]), .A2(inbar[201]), .ZN(n842bar);
  OR2_X1 U121 ( .A1(in[237]), .A2(n841), .ZN(n843) );
  AND2_X1 U121bar ( .A1(inbar[237]), .A2(n841bar), .ZN(n843bar);
  OR2_X1 U122 ( .A1(in[94]), .A2(in[253]), .ZN(n841) );
  AND2_X1 U122bar ( .A1(inbar[94]), .A2(inbar[253]), .ZN(n841bar);
  OR2_X1 U123 ( .A1(n840), .A2(n839), .ZN(n845) );
  AND2_X1 U123bar ( .A1(n840bar), .A2(n839bar), .ZN(n845bar);
  OR2_X1 U124 ( .A1(in_21), .A2(in[96]), .ZN(n839) );
  AND2_X1 U124bar ( .A1(in_21bar), .A2(inbar[96]), .ZN(n839bar);
  OR2_X1 U125 ( .A1(in_25), .A2(n838), .ZN(n840) );
  AND2_X1 U125bar ( .A1(in_25bar), .A2(n838bar), .ZN(n840bar);
  OR2_X1 U126 ( .A1(in_81), .A2(in_45), .ZN(n838) );
  AND2_X1 U126bar ( .A1(in_81bar), .A2(in_45bar), .ZN(n838bar);
  OR2_X1 U127 ( .A1(n837), .A2(n836), .ZN(n891) );
  AND2_X1 U127bar ( .A1(n837bar), .A2(n836bar), .ZN(n891bar);
  OR2_X1 U128 ( .A1(in[142]), .A2(in[124]), .ZN(n836) );
  AND2_X1 U128bar ( .A1(inbar[142]), .A2(inbar[124]), .ZN(n836bar);
  OR2_X1 U129 ( .A1(in[150]), .A2(n835), .ZN(n837) );
  AND2_X1 U129bar ( .A1(inbar[150]), .A2(n835bar), .ZN(n837bar);
  OR2_X1 U130 ( .A1(in[172]), .A2(in[155]), .ZN(n835) );
  AND2_X1 U130bar ( .A1(inbar[172]), .A2(inbar[155]), .ZN(n835bar);
  OR2_X1 U131 ( .A1(n834), .A2(n833), .ZN(n893) );
  AND2_X1 U131bar ( .A1(n834bar), .A2(n833bar), .ZN(n893bar);
  OR2_X1 U132 ( .A1(n832), .A2(n831), .ZN(n833) );
  AND2_X1 U132bar ( .A1(n832bar), .A2(n831bar), .ZN(n833bar);
  OR2_X1 U133 ( .A1(in[196]), .A2(in[173]), .ZN(n831) );
  AND2_X1 U133bar ( .A1(inbar[196]), .A2(inbar[173]), .ZN(n831bar);
  OR2_X1 U134 ( .A1(in[222]), .A2(n830), .ZN(n832) );
  AND2_X1 U134bar ( .A1(inbar[222]), .A2(n830bar), .ZN(n832bar);
  OR2_X1 U135 ( .A1(in[227]), .A2(in[226]), .ZN(n830) );
  AND2_X1 U135bar ( .A1(inbar[227]), .A2(inbar[226]), .ZN(n830bar);
  OR2_X1 U136 ( .A1(n829), .A2(n828), .ZN(n834) );
  AND2_X1 U136bar ( .A1(n829bar), .A2(n828bar), .ZN(n834bar);
  OR2_X1 U137 ( .A1(in[249]), .A2(in[231]), .ZN(n828) );
  AND2_X1 U137bar ( .A1(inbar[249]), .A2(inbar[231]), .ZN(n828bar);
  OR2_X1 U138 ( .A1(in_28), .A2(n827), .ZN(n829) );
  AND2_X1 U138bar ( .A1(in_28bar), .A2(n827bar), .ZN(n829bar);
  OR2_X1 U139 ( .A1(in_52), .A2(in_47), .ZN(n827) );
  AND2_X1 U139bar ( .A1(in_52bar), .A2(in_47bar), .ZN(n827bar);
  OR2_X1 U140 ( .A1(n826), .A2(n825), .ZN(out[3]) );
  AND2_X1 U140bar ( .A1(n826bar), .A2(n825bar), .ZN(outbar[3]);
  OR2_X1 U141 ( .A1(n824), .A2(n823), .ZN(n825) );
  AND2_X1 U141bar ( .A1(n824bar), .A2(n823bar), .ZN(n825bar);
  OR2_X1 U142 ( .A1(n822), .A2(n821), .ZN(n823) );
  AND2_X1 U142bar ( .A1(n822bar), .A2(n821bar), .ZN(n823bar);
  OR2_X1 U143 ( .A1(n820), .A2(n819), .ZN(n821) );
  AND2_X1 U143bar ( .A1(n820bar), .A2(n819bar), .ZN(n821bar);
  OR2_X1 U144 ( .A1(n964), .A2(n818), .ZN(n822) );
  AND2_X1 U144bar ( .A1(n964bar), .A2(n818bar), .ZN(n822bar);
  OR2_X1 U145 ( .A1(in[118]), .A2(n817), .ZN(n818) );
  AND2_X1 U145bar ( .A1(inbar[118]), .A2(n817bar), .ZN(n818bar);
  OR2_X1 U146 ( .A1(n816), .A2(n815), .ZN(n964) );
  AND2_X1 U146bar ( .A1(n816bar), .A2(n815bar), .ZN(n964bar);
  OR2_X1 U147 ( .A1(n814), .A2(n813), .ZN(n815) );
  AND2_X1 U147bar ( .A1(n814bar), .A2(n813bar), .ZN(n815bar);
  OR2_X1 U148 ( .A1(n812), .A2(n811), .ZN(n813) );
  AND2_X1 U148bar ( .A1(n812bar), .A2(n811bar), .ZN(n813bar);
  OR2_X1 U149 ( .A1(in[122]), .A2(in[111]), .ZN(n811) );
  AND2_X1 U149bar ( .A1(inbar[122]), .A2(inbar[111]), .ZN(n811bar);
  OR2_X1 U150 ( .A1(in[154]), .A2(in[151]), .ZN(n812) );
  AND2_X1 U150bar ( .A1(inbar[154]), .A2(inbar[151]), .ZN(n812bar);
  OR2_X1 U151 ( .A1(n810), .A2(n809), .ZN(n814) );
  AND2_X1 U151bar ( .A1(n810bar), .A2(n809bar), .ZN(n814bar);
  OR2_X1 U152 ( .A1(in[187]), .A2(in[177]), .ZN(n809) );
  AND2_X1 U152bar ( .A1(inbar[187]), .A2(inbar[177]), .ZN(n809bar);
  OR2_X1 U153 ( .A1(in[200]), .A2(in[192]), .ZN(n810) );
  AND2_X1 U153bar ( .A1(inbar[200]), .A2(inbar[192]), .ZN(n810bar);
  OR2_X1 U154 ( .A1(n808), .A2(n807), .ZN(n816) );
  AND2_X1 U154bar ( .A1(n808bar), .A2(n807bar), .ZN(n816bar);
  OR2_X1 U155 ( .A1(n806), .A2(n805), .ZN(n807) );
  AND2_X1 U155bar ( .A1(n806bar), .A2(n805bar), .ZN(n807bar);
  OR2_X1 U156 ( .A1(in[225]), .A2(in[207]), .ZN(n805) );
  AND2_X1 U156bar ( .A1(inbar[225]), .A2(inbar[207]), .ZN(n805bar);
  OR2_X1 U157 ( .A1(in[98]), .A2(in[226]), .ZN(n806) );
  AND2_X1 U157bar ( .A1(inbar[98]), .A2(inbar[226]), .ZN(n806bar);
  OR2_X1 U158 ( .A1(n804), .A2(n803), .ZN(n808) );
  AND2_X1 U158bar ( .A1(n804bar), .A2(n803bar), .ZN(n808bar);
  OR2_X1 U159 ( .A1(in_20), .A2(in_16), .ZN(n803) );
  AND2_X1 U159bar ( .A1(in_20bar), .A2(in_16bar), .ZN(n803bar);
  OR2_X1 U160 ( .A1(in_55), .A2(in_45), .ZN(n804) );
  AND2_X1 U160bar ( .A1(in_55bar), .A2(in_45bar), .ZN(n804bar);
  OR2_X1 U161 ( .A1(n802), .A2(n801), .ZN(n824) );
  AND2_X1 U161bar ( .A1(n802bar), .A2(n801bar), .ZN(n824bar);
  OR2_X1 U162 ( .A1(in[162]), .A2(in[149]), .ZN(n801) );
  AND2_X1 U162bar ( .A1(inbar[162]), .A2(inbar[149]), .ZN(n801bar);
  OR2_X1 U163 ( .A1(in[163]), .A2(n800), .ZN(n802) );
  AND2_X1 U163bar ( .A1(inbar[163]), .A2(n800bar), .ZN(n802bar);
  OR2_X1 U164 ( .A1(in[191]), .A2(in[189]), .ZN(n800) );
  AND2_X1 U164bar ( .A1(inbar[191]), .A2(inbar[189]), .ZN(n800bar);
  OR2_X1 U165 ( .A1(n799), .A2(n798), .ZN(n826) );
  AND2_X1 U165bar ( .A1(n799bar), .A2(n798bar), .ZN(n826bar);
  OR2_X1 U166 ( .A1(n797), .A2(n796), .ZN(n798) );
  AND2_X1 U166bar ( .A1(n797bar), .A2(n796bar), .ZN(n798bar);
  OR2_X1 U167 ( .A1(in[212]), .A2(in[193]), .ZN(n796) );
  AND2_X1 U167bar ( .A1(inbar[212]), .A2(inbar[193]), .ZN(n796bar);
  OR2_X1 U168 ( .A1(in[238]), .A2(n795), .ZN(n797) );
  AND2_X1 U168bar ( .A1(inbar[238]), .A2(n795bar), .ZN(n797bar);
  OR2_X1 U169 ( .A1(in[88]), .A2(in[247]), .ZN(n795) );
  AND2_X1 U169bar ( .A1(inbar[88]), .A2(inbar[247]), .ZN(n795bar);
  OR2_X1 U170 ( .A1(n794), .A2(n793), .ZN(n799) );
  AND2_X1 U170bar ( .A1(n794bar), .A2(n793bar), .ZN(n799bar);
  OR2_X1 U171 ( .A1(in[94]), .A2(in[92]), .ZN(n793) );
  AND2_X1 U171bar ( .A1(inbar[94]), .A2(inbar[92]), .ZN(n793bar);
  OR2_X1 U172 ( .A1(in_52), .A2(n792), .ZN(n794) );
  AND2_X1 U172bar ( .A1(in_52bar), .A2(n792bar), .ZN(n794bar);
  OR2_X1 U173 ( .A1(in_70), .A2(in_67), .ZN(n792) );
  AND2_X1 U173bar ( .A1(in_70bar), .A2(in_67bar), .ZN(n792bar);
  OR2_X1 U174 ( .A1(n791), .A2(n790), .ZN(out[2]) );
  AND2_X1 U174bar ( .A1(n791bar), .A2(n790bar), .ZN(outbar[2]);
  OR2_X1 U175 ( .A1(n789), .A2(n788), .ZN(n790) );
  AND2_X1 U175bar ( .A1(n789bar), .A2(n788bar), .ZN(n790bar);
  OR2_X1 U176 ( .A1(n787), .A2(n786), .ZN(n788) );
  AND2_X1 U176bar ( .A1(n787bar), .A2(n786bar), .ZN(n788bar);
  OR2_X1 U177 ( .A1(n819), .A2(n785), .ZN(n786) );
  AND2_X1 U177bar ( .A1(n819bar), .A2(n785bar), .ZN(n786bar);
  OR2_X1 U178 ( .A1(n784), .A2(n783), .ZN(n819) );
  AND2_X1 U178bar ( .A1(n784bar), .A2(n783bar), .ZN(n819bar);
  OR2_X1 U179 ( .A1(n782), .A2(n781), .ZN(n783) );
  AND2_X1 U179bar ( .A1(n782bar), .A2(n781bar), .ZN(n783bar);
  OR2_X1 U180 ( .A1(n780), .A2(n779), .ZN(n781) );
  AND2_X1 U180bar ( .A1(n780bar), .A2(n779bar), .ZN(n781bar);
  OR2_X1 U181 ( .A1(n962), .A2(n778), .ZN(n779) );
  AND2_X1 U181bar ( .A1(n962bar), .A2(n778bar), .ZN(n779bar);
  OR2_X1 U182 ( .A1(n777), .A2(n776), .ZN(n962) );
  AND2_X1 U182bar ( .A1(n777bar), .A2(n776bar), .ZN(n962bar);
  OR2_X1 U183 ( .A1(n775), .A2(n774), .ZN(n776) );
  AND2_X1 U183bar ( .A1(n775bar), .A2(n774bar), .ZN(n776bar);
  OR2_X1 U184 ( .A1(n773), .A2(n772), .ZN(n774) );
  AND2_X1 U184bar ( .A1(n773bar), .A2(n772bar), .ZN(n774bar);
  OR2_X1 U185 ( .A1(in[131]), .A2(in[120]), .ZN(n772) );
  AND2_X1 U185bar ( .A1(inbar[131]), .A2(inbar[120]), .ZN(n772bar);
  OR2_X1 U186 ( .A1(in[153]), .A2(in[147]), .ZN(n773) );
  AND2_X1 U186bar ( .A1(inbar[153]), .A2(inbar[147]), .ZN(n773bar);
  OR2_X1 U187 ( .A1(n771), .A2(n770), .ZN(n775) );
  AND2_X1 U187bar ( .A1(n771bar), .A2(n770bar), .ZN(n775bar);
  OR2_X1 U188 ( .A1(in[170]), .A2(in[156]), .ZN(n770) );
  AND2_X1 U188bar ( .A1(inbar[170]), .A2(inbar[156]), .ZN(n770bar);
  OR2_X1 U189 ( .A1(in[223]), .A2(in[190]), .ZN(n771) );
  AND2_X1 U189bar ( .A1(inbar[223]), .A2(inbar[190]), .ZN(n771bar);
  OR2_X1 U190 ( .A1(n769), .A2(n768), .ZN(n777) );
  AND2_X1 U190bar ( .A1(n769bar), .A2(n768bar), .ZN(n777bar);
  OR2_X1 U191 ( .A1(n767), .A2(n766), .ZN(n768) );
  AND2_X1 U191bar ( .A1(n767bar), .A2(n766bar), .ZN(n768bar);
  OR2_X1 U192 ( .A1(in[236]), .A2(in[230]), .ZN(n766) );
  AND2_X1 U192bar ( .A1(inbar[236]), .A2(inbar[230]), .ZN(n766bar);
  OR2_X1 U193 ( .A1(in[85]), .A2(in[240]), .ZN(n767) );
  AND2_X1 U193bar ( .A1(inbar[85]), .A2(inbar[240]), .ZN(n767bar);
  OR2_X1 U194 ( .A1(n765), .A2(n764), .ZN(n769) );
  AND2_X1 U194bar ( .A1(n765bar), .A2(n764bar), .ZN(n769bar);
  OR2_X1 U195 ( .A1(in_12), .A2(in[90]), .ZN(n764) );
  AND2_X1 U195bar ( .A1(in_12bar), .A2(inbar[90]), .ZN(n764bar);
  OR2_X1 U196 ( .A1(in_39), .A2(in_28), .ZN(n765) );
  AND2_X1 U196bar ( .A1(in_39bar), .A2(in_28bar), .ZN(n765bar);
  OR2_X1 U197 ( .A1(in[109]), .A2(n763), .ZN(n780) );
  AND2_X1 U197bar ( .A1(inbar[109]), .A2(n763bar), .ZN(n780bar);
  OR2_X1 U198 ( .A1(n762), .A2(n761), .ZN(n782) );
  AND2_X1 U198bar ( .A1(n762bar), .A2(n761bar), .ZN(n782bar);
  OR2_X1 U199 ( .A1(in[138]), .A2(in[129]), .ZN(n761) );
  AND2_X1 U199bar ( .A1(inbar[138]), .A2(inbar[129]), .ZN(n761bar);
  OR2_X1 U200 ( .A1(in[157]), .A2(n760), .ZN(n762) );
  AND2_X1 U200bar ( .A1(inbar[157]), .A2(n760bar), .ZN(n762bar);
  OR2_X1 U201 ( .A1(in[182]), .A2(in[167]), .ZN(n760) );
  AND2_X1 U201bar ( .A1(inbar[182]), .A2(inbar[167]), .ZN(n760bar);
  OR2_X1 U202 ( .A1(n759), .A2(n758), .ZN(n784) );
  AND2_X1 U202bar ( .A1(n759bar), .A2(n758bar), .ZN(n784bar);
  OR2_X1 U203 ( .A1(n757), .A2(n756), .ZN(n758) );
  AND2_X1 U203bar ( .A1(n757bar), .A2(n756bar), .ZN(n758bar);
  OR2_X1 U204 ( .A1(in[195]), .A2(in[184]), .ZN(n756) );
  AND2_X1 U204bar ( .A1(inbar[195]), .A2(inbar[184]), .ZN(n756bar);
  OR2_X1 U205 ( .A1(in[196]), .A2(n755), .ZN(n757) );
  AND2_X1 U205bar ( .A1(inbar[196]), .A2(n755bar), .ZN(n757bar);
  OR2_X1 U206 ( .A1(in[215]), .A2(in[209]), .ZN(n755) );
  AND2_X1 U206bar ( .A1(inbar[215]), .A2(inbar[209]), .ZN(n755bar);
  OR2_X1 U207 ( .A1(n754), .A2(n753), .ZN(n759) );
  AND2_X1 U207bar ( .A1(n754bar), .A2(n753bar), .ZN(n759bar);
  OR2_X1 U208 ( .A1(in[93]), .A2(in[233]), .ZN(n753) );
  AND2_X1 U208bar ( .A1(inbar[93]), .A2(inbar[233]), .ZN(n753bar);
  OR2_X1 U209 ( .A1(in_1), .A2(n752), .ZN(n754) );
  AND2_X1 U209bar ( .A1(in_1bar), .A2(n752bar), .ZN(n754bar);
  OR2_X1 U210 ( .A1(in_69), .A2(in_66), .ZN(n752) );
  AND2_X1 U210bar ( .A1(in_69bar), .A2(in_66bar), .ZN(n752bar);
  OR2_X1 U211 ( .A1(n966), .A2(n751), .ZN(n787) );
  AND2_X1 U211bar ( .A1(n966bar), .A2(n751bar), .ZN(n787bar);
  OR2_X1 U212 ( .A1(in[134]), .A2(n750), .ZN(n751) );
  AND2_X1 U212bar ( .A1(inbar[134]), .A2(n750bar), .ZN(n751bar);
  OR2_X1 U213 ( .A1(n749), .A2(n748), .ZN(n966) );
  AND2_X1 U213bar ( .A1(n749bar), .A2(n748bar), .ZN(n966bar);
  OR2_X1 U214 ( .A1(n747), .A2(n746), .ZN(n748) );
  AND2_X1 U214bar ( .A1(n747bar), .A2(n746bar), .ZN(n748bar);
  OR2_X1 U215 ( .A1(n745), .A2(n744), .ZN(n746) );
  AND2_X1 U215bar ( .A1(n745bar), .A2(n744bar), .ZN(n746bar);
  OR2_X1 U216 ( .A1(in[136]), .A2(in[121]), .ZN(n744) );
  AND2_X1 U216bar ( .A1(inbar[136]), .A2(inbar[121]), .ZN(n744bar);
  OR2_X1 U217 ( .A1(in[186]), .A2(in[174]), .ZN(n745) );
  AND2_X1 U217bar ( .A1(inbar[186]), .A2(inbar[174]), .ZN(n745bar);
  OR2_X1 U218 ( .A1(n743), .A2(n742), .ZN(n747) );
  AND2_X1 U218bar ( .A1(n743bar), .A2(n742bar), .ZN(n747bar);
  OR2_X1 U219 ( .A1(in[198]), .A2(in[197]), .ZN(n742) );
  AND2_X1 U219bar ( .A1(inbar[198]), .A2(inbar[197]), .ZN(n742bar);
  OR2_X1 U220 ( .A1(in[214]), .A2(in[199]), .ZN(n743) );
  AND2_X1 U220bar ( .A1(inbar[214]), .A2(inbar[199]), .ZN(n743bar);
  OR2_X1 U221 ( .A1(n741), .A2(n740), .ZN(n749) );
  AND2_X1 U221bar ( .A1(n741bar), .A2(n740bar), .ZN(n749bar);
  OR2_X1 U222 ( .A1(n739), .A2(n738), .ZN(n740) );
  AND2_X1 U222bar ( .A1(n739bar), .A2(n738bar), .ZN(n740bar);
  OR2_X1 U223 ( .A1(in[231]), .A2(in[220]), .ZN(n738) );
  AND2_X1 U223bar ( .A1(inbar[231]), .A2(inbar[220]), .ZN(n738bar);
  OR2_X1 U224 ( .A1(in_25), .A2(in[245]), .ZN(n739) );
  AND2_X1 U224bar ( .A1(in_25bar), .A2(inbar[245]), .ZN(n739bar);
  OR2_X1 U225 ( .A1(n737), .A2(n736), .ZN(n741) );
  AND2_X1 U225bar ( .A1(n737bar), .A2(n736bar), .ZN(n741bar);
  OR2_X1 U226 ( .A1(in_53), .A2(in_29), .ZN(n736) );
  AND2_X1 U226bar ( .A1(in_53bar), .A2(in_29bar), .ZN(n736bar);
  OR2_X1 U227 ( .A1(in_79), .A2(in_74), .ZN(n737) );
  AND2_X1 U227bar ( .A1(in_79bar), .A2(in_74bar), .ZN(n737bar);
  OR2_X1 U228 ( .A1(n735), .A2(n734), .ZN(n789) );
  AND2_X1 U228bar ( .A1(n735bar), .A2(n734bar), .ZN(n789bar);
  OR2_X1 U229 ( .A1(in[152]), .A2(in[140]), .ZN(n734) );
  AND2_X1 U229bar ( .A1(inbar[152]), .A2(inbar[140]), .ZN(n734bar);
  OR2_X1 U230 ( .A1(in[155]), .A2(n733), .ZN(n735) );
  AND2_X1 U230bar ( .A1(inbar[155]), .A2(n733bar), .ZN(n735bar);
  OR2_X1 U231 ( .A1(in[166]), .A2(in[165]), .ZN(n733) );
  AND2_X1 U231bar ( .A1(inbar[166]), .A2(inbar[165]), .ZN(n733bar);
  OR2_X1 U232 ( .A1(n732), .A2(n731), .ZN(n791) );
  AND2_X1 U232bar ( .A1(n732bar), .A2(n731bar), .ZN(n791bar);
  OR2_X1 U233 ( .A1(n730), .A2(n729), .ZN(n731) );
  AND2_X1 U233bar ( .A1(n730bar), .A2(n729bar), .ZN(n731bar);
  OR2_X1 U234 ( .A1(in[202]), .A2(in[185]), .ZN(n729) );
  AND2_X1 U234bar ( .A1(inbar[202]), .A2(inbar[185]), .ZN(n729bar);
  OR2_X1 U235 ( .A1(in[211]), .A2(n728), .ZN(n730) );
  AND2_X1 U235bar ( .A1(inbar[211]), .A2(n728bar), .ZN(n730bar);
  OR2_X1 U236 ( .A1(in[255]), .A2(in[253]), .ZN(n728) );
  AND2_X1 U236bar ( .A1(inbar[255]), .A2(inbar[253]), .ZN(n728bar);
  OR2_X1 U237 ( .A1(n727), .A2(n726), .ZN(n732) );
  AND2_X1 U237bar ( .A1(n727bar), .A2(n726bar), .ZN(n732bar);
  OR2_X1 U238 ( .A1(in_35), .A2(in_15), .ZN(n726) );
  AND2_X1 U238bar ( .A1(in_35bar), .A2(in_15bar), .ZN(n726bar);
  OR2_X1 U239 ( .A1(in_36), .A2(n725), .ZN(n727) );
  AND2_X1 U239bar ( .A1(in_36bar), .A2(n725bar), .ZN(n727bar);
  OR2_X1 U240 ( .A1(in_48), .A2(in_40), .ZN(n725) );
  AND2_X1 U240bar ( .A1(in_48bar), .A2(in_40bar), .ZN(n725bar);
  OR2_X1 U241 ( .A1(n724), .A2(n723), .ZN(out[1]) );
  AND2_X1 U241bar ( .A1(n724bar), .A2(n723bar), .ZN(outbar[1]);
  OR2_X1 U242 ( .A1(n722), .A2(n721), .ZN(n723) );
  AND2_X1 U242bar ( .A1(n722bar), .A2(n721bar), .ZN(n723bar);
  OR2_X1 U243 ( .A1(n720), .A2(n719), .ZN(n721) );
  AND2_X1 U243bar ( .A1(n720bar), .A2(n719bar), .ZN(n721bar);
  OR2_X1 U244 ( .A1(n921), .A2(n887), .ZN(n719) );
  AND2_X1 U244bar ( .A1(n921bar), .A2(n887bar), .ZN(n719bar);
  OR2_X1 U245 ( .A1(n718), .A2(n717), .ZN(n887) );
  AND2_X1 U245bar ( .A1(n718bar), .A2(n717bar), .ZN(n887bar);
  OR2_X1 U246 ( .A1(n716), .A2(n715), .ZN(n717) );
  AND2_X1 U246bar ( .A1(n716bar), .A2(n715bar), .ZN(n717bar);
  OR2_X1 U247 ( .A1(n714), .A2(n713), .ZN(n715) );
  AND2_X1 U247bar ( .A1(n714bar), .A2(n713bar), .ZN(n715bar);
  OR2_X1 U248 ( .A1(in[116]), .A2(in[110]), .ZN(n713) );
  AND2_X1 U248bar ( .A1(inbar[116]), .A2(inbar[110]), .ZN(n713bar);
  OR2_X1 U249 ( .A1(in[133]), .A2(in[130]), .ZN(n714) );
  AND2_X1 U249bar ( .A1(inbar[133]), .A2(inbar[130]), .ZN(n714bar);
  OR2_X1 U250 ( .A1(n712), .A2(n711), .ZN(n716) );
  AND2_X1 U250bar ( .A1(n712bar), .A2(n711bar), .ZN(n716bar);
  OR2_X1 U251 ( .A1(in[203]), .A2(in[135]), .ZN(n711) );
  AND2_X1 U251bar ( .A1(inbar[203]), .A2(inbar[135]), .ZN(n711bar);
  OR2_X1 U252 ( .A1(in[232]), .A2(in[223]), .ZN(n712) );
  AND2_X1 U252bar ( .A1(inbar[232]), .A2(inbar[223]), .ZN(n712bar);
  OR2_X1 U253 ( .A1(n710), .A2(n709), .ZN(n718) );
  AND2_X1 U253bar ( .A1(n710bar), .A2(n709bar), .ZN(n718bar);
  OR2_X1 U254 ( .A1(n708), .A2(n707), .ZN(n709) );
  AND2_X1 U254bar ( .A1(n708bar), .A2(n707bar), .ZN(n709bar);
  OR2_X1 U255 ( .A1(in[255]), .A2(in[233]), .ZN(n707) );
  AND2_X1 U255bar ( .A1(inbar[255]), .A2(inbar[233]), .ZN(n707bar);
  OR2_X1 U256 ( .A1(in_53), .A2(in_34), .ZN(n708) );
  AND2_X1 U256bar ( .A1(in_53bar), .A2(in_34bar), .ZN(n708bar);
  OR2_X1 U257 ( .A1(n706), .A2(n705), .ZN(n710) );
  AND2_X1 U257bar ( .A1(n706bar), .A2(n705bar), .ZN(n710bar);
  OR2_X1 U258 ( .A1(in_57), .A2(in_55), .ZN(n705) );
  AND2_X1 U258bar ( .A1(in_57bar), .A2(in_55bar), .ZN(n705bar);
  OR2_X1 U259 ( .A1(in_68), .A2(in_67), .ZN(n706) );
  AND2_X1 U259bar ( .A1(in_68bar), .A2(in_67bar), .ZN(n706bar);
  OR2_X1 U260 ( .A1(n704), .A2(n703), .ZN(n921) );
  AND2_X1 U260bar ( .A1(n704bar), .A2(n703bar), .ZN(n921bar);
  OR2_X1 U261 ( .A1(n702), .A2(n701), .ZN(n703) );
  AND2_X1 U261bar ( .A1(n702bar), .A2(n701bar), .ZN(n703bar);
  OR2_X1 U262 ( .A1(n700), .A2(n699), .ZN(n701) );
  AND2_X1 U262bar ( .A1(n700bar), .A2(n699bar), .ZN(n701bar);
  OR2_X1 U263 ( .A1(n944), .A2(n872), .ZN(n699) );
  AND2_X1 U263bar ( .A1(n944bar), .A2(n872bar), .ZN(n699bar);
  OR2_X1 U264 ( .A1(n698), .A2(n697), .ZN(n872) );
  AND2_X1 U264bar ( .A1(n698bar), .A2(n697bar), .ZN(n872bar);
  OR2_X1 U265 ( .A1(n696), .A2(n695), .ZN(n697) );
  AND2_X1 U265bar ( .A1(n696bar), .A2(n695bar), .ZN(n697bar);
  OR2_X1 U266 ( .A1(n694), .A2(n693), .ZN(n695) );
  AND2_X1 U266bar ( .A1(n694bar), .A2(n693bar), .ZN(n695bar);
  OR2_X1 U267 ( .A1(in[121]), .A2(in[102]), .ZN(n693) );
  AND2_X1 U267bar ( .A1(inbar[121]), .A2(inbar[102]), .ZN(n693bar);
  OR2_X1 U268 ( .A1(in[162]), .A2(in[161]), .ZN(n694) );
  AND2_X1 U268bar ( .A1(inbar[162]), .A2(inbar[161]), .ZN(n694bar);
  OR2_X1 U269 ( .A1(n692), .A2(n691), .ZN(n696) );
  AND2_X1 U269bar ( .A1(n692bar), .A2(n691bar), .ZN(n696bar);
  OR2_X1 U270 ( .A1(in[192]), .A2(in[178]), .ZN(n691) );
  AND2_X1 U270bar ( .A1(inbar[192]), .A2(inbar[178]), .ZN(n691bar);
  OR2_X1 U271 ( .A1(in[244]), .A2(in[209]), .ZN(n692) );
  AND2_X1 U271bar ( .A1(inbar[244]), .A2(inbar[209]), .ZN(n692bar);
  OR2_X1 U272 ( .A1(n690), .A2(n689), .ZN(n698) );
  AND2_X1 U272bar ( .A1(n690bar), .A2(n689bar), .ZN(n698bar);
  OR2_X1 U273 ( .A1(n688), .A2(n687), .ZN(n689) );
  AND2_X1 U273bar ( .A1(n688bar), .A2(n687bar), .ZN(n689bar);
  OR2_X1 U274 ( .A1(in[90]), .A2(in[254]), .ZN(n687) );
  AND2_X1 U274bar ( .A1(inbar[90]), .A2(inbar[254]), .ZN(n687bar);
  OR2_X1 U275 ( .A1(in_36), .A2(in_32), .ZN(n688) );
  AND2_X1 U275bar ( .A1(in_36bar), .A2(in_32bar), .ZN(n688bar);
  OR2_X1 U276 ( .A1(n686), .A2(n685), .ZN(n690) );
  AND2_X1 U276bar ( .A1(n686bar), .A2(n685bar), .ZN(n690bar);
  OR2_X1 U277 ( .A1(in_62), .A2(in_37), .ZN(n685) );
  AND2_X1 U277bar ( .A1(in_62bar), .A2(in_37bar), .ZN(n685bar);
  OR2_X1 U278 ( .A1(in_75), .A2(in_73), .ZN(n686) );
  AND2_X1 U278bar ( .A1(in_75bar), .A2(in_73bar), .ZN(n686bar);
  OR2_X1 U279 ( .A1(n684), .A2(n683), .ZN(n944) );
  AND2_X1 U279bar ( .A1(n684bar), .A2(n683bar), .ZN(n944bar);
  OR2_X1 U280 ( .A1(n682), .A2(n681), .ZN(n683) );
  AND2_X1 U280bar ( .A1(n682bar), .A2(n681bar), .ZN(n683bar);
  OR2_X1 U281 ( .A1(n680), .A2(n679), .ZN(n681) );
  AND2_X1 U281bar ( .A1(n680bar), .A2(n679bar), .ZN(n681bar);
  OR2_X1 U282 ( .A1(in[171]), .A2(in[153]), .ZN(n679) );
  AND2_X1 U282bar ( .A1(inbar[171]), .A2(inbar[153]), .ZN(n679bar);
  OR2_X1 U283 ( .A1(in[187]), .A2(in[176]), .ZN(n680) );
  AND2_X1 U283bar ( .A1(inbar[187]), .A2(inbar[176]), .ZN(n680bar);
  OR2_X1 U284 ( .A1(n678), .A2(n677), .ZN(n682) );
  AND2_X1 U284bar ( .A1(n678bar), .A2(n677bar), .ZN(n682bar);
  OR2_X1 U285 ( .A1(in[245]), .A2(in[211]), .ZN(n677) );
  AND2_X1 U285bar ( .A1(inbar[245]), .A2(inbar[211]), .ZN(n677bar);
  OR2_X1 U286 ( .A1(in[97]), .A2(in[88]), .ZN(n678) );
  AND2_X1 U286bar ( .A1(inbar[97]), .A2(inbar[88]), .ZN(n678bar);
  OR2_X1 U287 ( .A1(n676), .A2(n675), .ZN(n684) );
  AND2_X1 U287bar ( .A1(n676bar), .A2(n675bar), .ZN(n684bar);
  OR2_X1 U288 ( .A1(n674), .A2(n673), .ZN(n675) );
  AND2_X1 U288bar ( .A1(n674bar), .A2(n673bar), .ZN(n675bar);
  OR2_X1 U289 ( .A1(in_10), .A2(in_0), .ZN(n673) );
  AND2_X1 U289bar ( .A1(in_10bar), .A2(in_0bar), .ZN(n673bar);
  OR2_X1 U290 ( .A1(in_59), .A2(in_5), .ZN(n674) );
  AND2_X1 U290bar ( .A1(in_59bar), .A2(in_5bar), .ZN(n674bar);
  OR2_X1 U291 ( .A1(n672), .A2(n671), .ZN(n676) );
  AND2_X1 U291bar ( .A1(n672bar), .A2(n671bar), .ZN(n676bar);
  OR2_X1 U292 ( .A1(in_60), .A2(in_6), .ZN(n671) );
  AND2_X1 U292bar ( .A1(in_60bar), .A2(in_6bar), .ZN(n671bar);
  OR2_X1 U293 ( .A1(in_77), .A2(in_69), .ZN(n672) );
  AND2_X1 U293bar ( .A1(in_77bar), .A2(in_69bar), .ZN(n672bar);
  OR2_X1 U294 ( .A1(in[113]), .A2(n864), .ZN(n700) );
  AND2_X1 U294bar ( .A1(inbar[113]), .A2(n864bar), .ZN(n700bar);
  OR2_X1 U295 ( .A1(n670), .A2(n669), .ZN(n864) );
  AND2_X1 U295bar ( .A1(n670bar), .A2(n669bar), .ZN(n864bar);
  OR2_X1 U296 ( .A1(n668), .A2(n667), .ZN(n669) );
  AND2_X1 U296bar ( .A1(n668bar), .A2(n667bar), .ZN(n669bar);
  OR2_X1 U297 ( .A1(n666), .A2(n665), .ZN(n667) );
  AND2_X1 U297bar ( .A1(n666bar), .A2(n665bar), .ZN(n667bar);
  OR2_X1 U298 ( .A1(in[125]), .A2(in[107]), .ZN(n665) );
  AND2_X1 U298bar ( .A1(inbar[125]), .A2(inbar[107]), .ZN(n665bar);
  OR2_X1 U299 ( .A1(in[138]), .A2(in[126]), .ZN(n666) );
  AND2_X1 U299bar ( .A1(inbar[138]), .A2(inbar[126]), .ZN(n666bar);
  OR2_X1 U300 ( .A1(n664), .A2(n663), .ZN(n668) );
  AND2_X1 U300bar ( .A1(n664bar), .A2(n663bar), .ZN(n668bar);
  OR2_X1 U301 ( .A1(in[189]), .A2(in[143]), .ZN(n663) );
  AND2_X1 U301bar ( .A1(inbar[189]), .A2(inbar[143]), .ZN(n663bar);
  OR2_X1 U302 ( .A1(in[99]), .A2(in[214]), .ZN(n664) );
  AND2_X1 U302bar ( .A1(inbar[99]), .A2(inbar[214]), .ZN(n664bar);
  OR2_X1 U303 ( .A1(n662), .A2(n661), .ZN(n670) );
  AND2_X1 U303bar ( .A1(n662bar), .A2(n661bar), .ZN(n670bar);
  OR2_X1 U304 ( .A1(n660), .A2(n659), .ZN(n661) );
  AND2_X1 U304bar ( .A1(n660bar), .A2(n659bar), .ZN(n661bar);
  OR2_X1 U305 ( .A1(in_15), .A2(in_12), .ZN(n659) );
  AND2_X1 U305bar ( .A1(in_15bar), .A2(in_12bar), .ZN(n659bar);
  OR2_X1 U306 ( .A1(in_20), .A2(in_2), .ZN(n660) );
  AND2_X1 U306bar ( .A1(in_20bar), .A2(in_2bar), .ZN(n660bar);
  OR2_X1 U307 ( .A1(n658), .A2(n657), .ZN(n662) );
  AND2_X1 U307bar ( .A1(n658bar), .A2(n657bar), .ZN(n662bar);
  OR2_X1 U308 ( .A1(in_30), .A2(in_3), .ZN(n657) );
  AND2_X1 U308bar ( .A1(in_30bar), .A2(in_3bar), .ZN(n657bar);
  OR2_X1 U309 ( .A1(in_4), .A2(in_38), .ZN(n658) );
  AND2_X1 U309bar ( .A1(in_4bar), .A2(in_38bar), .ZN(n658bar);
  OR2_X1 U310 ( .A1(n656), .A2(n655), .ZN(n702) );
  AND2_X1 U310bar ( .A1(n656bar), .A2(n655bar), .ZN(n702bar);
  OR2_X1 U311 ( .A1(in[148]), .A2(in[137]), .ZN(n655) );
  AND2_X1 U311bar ( .A1(inbar[148]), .A2(inbar[137]), .ZN(n655bar);
  OR2_X1 U312 ( .A1(in[149]), .A2(n654), .ZN(n656) );
  AND2_X1 U312bar ( .A1(inbar[149]), .A2(n654bar), .ZN(n656bar);
  OR2_X1 U313 ( .A1(in[195]), .A2(in[190]), .ZN(n654) );
  AND2_X1 U313bar ( .A1(inbar[195]), .A2(inbar[190]), .ZN(n654bar);
  OR2_X1 U314 ( .A1(n653), .A2(n652), .ZN(n704) );
  AND2_X1 U314bar ( .A1(n653bar), .A2(n652bar), .ZN(n704bar);
  OR2_X1 U315 ( .A1(n651), .A2(n650), .ZN(n652) );
  AND2_X1 U315bar ( .A1(n651bar), .A2(n650bar), .ZN(n652bar);
  OR2_X1 U316 ( .A1(in[98]), .A2(in[197]), .ZN(n650) );
  AND2_X1 U316bar ( .A1(inbar[98]), .A2(inbar[197]), .ZN(n650bar);
  OR2_X1 U317 ( .A1(in_11), .A2(n649), .ZN(n651) );
  AND2_X1 U317bar ( .A1(in_11bar), .A2(n649bar), .ZN(n651bar);
  OR2_X1 U318 ( .A1(in_26), .A2(in_14), .ZN(n649) );
  AND2_X1 U318bar ( .A1(in_26bar), .A2(in_14bar), .ZN(n649bar);
  OR2_X1 U319 ( .A1(n648), .A2(n647), .ZN(n653) );
  AND2_X1 U319bar ( .A1(n648bar), .A2(n647bar), .ZN(n653bar);
  OR2_X1 U320 ( .A1(in_35), .A2(in_27), .ZN(n647) );
  AND2_X1 U320bar ( .A1(in_35bar), .A2(in_27bar), .ZN(n647bar);
  OR2_X1 U321 ( .A1(in_50), .A2(n646), .ZN(n648) );
  AND2_X1 U321bar ( .A1(in_50bar), .A2(n646bar), .ZN(n648bar);
  OR2_X1 U322 ( .A1(in_78), .A2(in_61), .ZN(n646) );
  AND2_X1 U322bar ( .A1(in_78bar), .A2(in_61bar), .ZN(n646bar);
  OR2_X1 U323 ( .A1(n942), .A2(n645), .ZN(n720) );
  AND2_X1 U323bar ( .A1(n942bar), .A2(n645bar), .ZN(n720bar);
  OR2_X1 U324 ( .A1(in[106]), .A2(n863), .ZN(n645) );
  AND2_X1 U324bar ( .A1(inbar[106]), .A2(n863bar), .ZN(n645bar);
  OR2_X1 U325 ( .A1(n644), .A2(n643), .ZN(n863) );
  AND2_X1 U325bar ( .A1(n644bar), .A2(n643bar), .ZN(n863bar);
  OR2_X1 U326 ( .A1(n642), .A2(n641), .ZN(n643) );
  AND2_X1 U326bar ( .A1(n642bar), .A2(n641bar), .ZN(n643bar);
  OR2_X1 U327 ( .A1(n640), .A2(n639), .ZN(n641) );
  AND2_X1 U327bar ( .A1(n640bar), .A2(n639bar), .ZN(n641bar);
  OR2_X1 U328 ( .A1(in[127]), .A2(in[122]), .ZN(n639) );
  AND2_X1 U328bar ( .A1(inbar[127]), .A2(inbar[122]), .ZN(n639bar);
  OR2_X1 U329 ( .A1(in[156]), .A2(in[132]), .ZN(n640) );
  AND2_X1 U329bar ( .A1(inbar[156]), .A2(inbar[132]), .ZN(n640bar);
  OR2_X1 U330 ( .A1(n638), .A2(n637), .ZN(n642) );
  AND2_X1 U330bar ( .A1(n638bar), .A2(n637bar), .ZN(n642bar);
  OR2_X1 U331 ( .A1(in[159]), .A2(in[157]), .ZN(n637) );
  AND2_X1 U331bar ( .A1(inbar[159]), .A2(inbar[157]), .ZN(n637bar);
  OR2_X1 U332 ( .A1(in[185]), .A2(in[169]), .ZN(n638) );
  AND2_X1 U332bar ( .A1(inbar[185]), .A2(inbar[169]), .ZN(n638bar);
  OR2_X1 U333 ( .A1(n636), .A2(n635), .ZN(n644) );
  AND2_X1 U333bar ( .A1(n636bar), .A2(n635bar), .ZN(n644bar);
  OR2_X1 U334 ( .A1(n634), .A2(n633), .ZN(n635) );
  AND2_X1 U334bar ( .A1(n634bar), .A2(n633bar), .ZN(n635bar);
  OR2_X1 U335 ( .A1(in[239]), .A2(in[218]), .ZN(n633) );
  AND2_X1 U335bar ( .A1(inbar[239]), .A2(inbar[218]), .ZN(n633bar);
  OR2_X1 U336 ( .A1(in_13), .A2(in[87]), .ZN(n634) );
  AND2_X1 U336bar ( .A1(in_13bar), .A2(inbar[87]), .ZN(n634bar);
  OR2_X1 U337 ( .A1(n632), .A2(n631), .ZN(n636) );
  AND2_X1 U337bar ( .A1(n632bar), .A2(n631bar), .ZN(n636bar);
  OR2_X1 U338 ( .A1(in_72), .A2(in_70), .ZN(n631) );
  AND2_X1 U338bar ( .A1(in_72bar), .A2(in_70bar), .ZN(n631bar);
  OR2_X1 U339 ( .A1(in_80), .A2(in_74), .ZN(n632) );
  AND2_X1 U339bar ( .A1(in_80bar), .A2(in_74bar), .ZN(n632bar);
  OR2_X1 U340 ( .A1(n630), .A2(n629), .ZN(n942) );
  AND2_X1 U340bar ( .A1(n630bar), .A2(n629bar), .ZN(n942bar);
  OR2_X1 U341 ( .A1(n628), .A2(n627), .ZN(n629) );
  AND2_X1 U341bar ( .A1(n628bar), .A2(n627bar), .ZN(n629bar);
  OR2_X1 U342 ( .A1(n626), .A2(n625), .ZN(n627) );
  AND2_X1 U342bar ( .A1(n626bar), .A2(n625bar), .ZN(n627bar);
  OR2_X1 U343 ( .A1(in[146]), .A2(in[100]), .ZN(n625) );
  AND2_X1 U343bar ( .A1(inbar[146]), .A2(inbar[100]), .ZN(n625bar);
  OR2_X1 U344 ( .A1(in[168]), .A2(in[152]), .ZN(n626) );
  AND2_X1 U344bar ( .A1(inbar[168]), .A2(inbar[152]), .ZN(n626bar);
  OR2_X1 U345 ( .A1(n624), .A2(n623), .ZN(n628) );
  AND2_X1 U345bar ( .A1(n624bar), .A2(n623bar), .ZN(n628bar);
  OR2_X1 U346 ( .A1(in[199]), .A2(in[182]), .ZN(n623) );
  AND2_X1 U346bar ( .A1(inbar[199]), .A2(inbar[182]), .ZN(n623bar);
  OR2_X1 U347 ( .A1(in[236]), .A2(in[204]), .ZN(n624) );
  AND2_X1 U347bar ( .A1(inbar[236]), .A2(inbar[204]), .ZN(n624bar);
  OR2_X1 U348 ( .A1(n622), .A2(n621), .ZN(n630) );
  AND2_X1 U348bar ( .A1(n622bar), .A2(n621bar), .ZN(n630bar);
  OR2_X1 U349 ( .A1(n620), .A2(n619), .ZN(n621) );
  AND2_X1 U349bar ( .A1(n620bar), .A2(n619bar), .ZN(n621bar);
  OR2_X1 U350 ( .A1(in[89]), .A2(in[246]), .ZN(n619) );
  AND2_X1 U350bar ( .A1(inbar[89]), .A2(inbar[246]), .ZN(n619bar);
  OR2_X1 U351 ( .A1(in[95]), .A2(in[92]), .ZN(n620) );
  AND2_X1 U351bar ( .A1(inbar[95]), .A2(inbar[92]), .ZN(n620bar);
  OR2_X1 U352 ( .A1(n618), .A2(n617), .ZN(n622) );
  AND2_X1 U352bar ( .A1(n618bar), .A2(n617bar), .ZN(n622bar);
  OR2_X1 U353 ( .A1(in_22), .A2(in_16), .ZN(n617) );
  AND2_X1 U353bar ( .A1(in_22bar), .A2(in_16bar), .ZN(n617bar);
  OR2_X1 U354 ( .A1(in_51), .A2(in_49), .ZN(n618) );
  AND2_X1 U354bar ( .A1(in_51bar), .A2(in_49bar), .ZN(n618bar);
  OR2_X1 U355 ( .A1(n616), .A2(n615), .ZN(n722) );
  AND2_X1 U355bar ( .A1(n616bar), .A2(n615bar), .ZN(n722bar);
  OR2_X1 U356 ( .A1(in[158]), .A2(in[115]), .ZN(n615) );
  AND2_X1 U356bar ( .A1(inbar[158]), .A2(inbar[115]), .ZN(n615bar);
  OR2_X1 U357 ( .A1(in[163]), .A2(n614), .ZN(n616) );
  AND2_X1 U357bar ( .A1(inbar[163]), .A2(n614bar), .ZN(n616bar);
  OR2_X1 U358 ( .A1(in[206]), .A2(in[165]), .ZN(n614) );
  AND2_X1 U358bar ( .A1(inbar[206]), .A2(inbar[165]), .ZN(n614bar);
  OR2_X1 U359 ( .A1(n613), .A2(n612), .ZN(n724) );
  AND2_X1 U359bar ( .A1(n613bar), .A2(n612bar), .ZN(n724bar);
  OR2_X1 U360 ( .A1(n611), .A2(n610), .ZN(n612) );
  AND2_X1 U360bar ( .A1(n611bar), .A2(n610bar), .ZN(n612bar);
  OR2_X1 U361 ( .A1(in[213]), .A2(in[207]), .ZN(n610) );
  AND2_X1 U361bar ( .A1(inbar[213]), .A2(inbar[207]), .ZN(n610bar);
  OR2_X1 U362 ( .A1(in[215]), .A2(n609), .ZN(n611) );
  AND2_X1 U362bar ( .A1(inbar[215]), .A2(n609bar), .ZN(n611bar);
  OR2_X1 U363 ( .A1(in[230]), .A2(in[220]), .ZN(n609) );
  AND2_X1 U363bar ( .A1(inbar[230]), .A2(inbar[220]), .ZN(n609bar);
  OR2_X1 U364 ( .A1(n608), .A2(n607), .ZN(n613) );
  AND2_X1 U364bar ( .A1(n608bar), .A2(n607bar), .ZN(n613bar);
  OR2_X1 U365 ( .A1(in[251]), .A2(in[234]), .ZN(n607) );
  AND2_X1 U365bar ( .A1(inbar[251]), .A2(inbar[234]), .ZN(n607bar);
  OR2_X1 U366 ( .A1(in_17), .A2(n606), .ZN(n608) );
  AND2_X1 U366bar ( .A1(in_17bar), .A2(n606bar), .ZN(n608bar);
  OR2_X1 U367 ( .A1(in_65), .A2(in_56), .ZN(n606) );
  AND2_X1 U367bar ( .A1(in_65bar), .A2(in_56bar), .ZN(n606bar);
  OR2_X1 U368 ( .A1(n605), .A2(n604), .ZN(out[0]) );
  AND2_X1 U368bar ( .A1(n605bar), .A2(n604bar), .ZN(outbar[0]);
  OR2_X1 U369 ( .A1(n603), .A2(n602), .ZN(n604) );
  AND2_X1 U369bar ( .A1(n603bar), .A2(n602bar), .ZN(n604bar);
  OR2_X1 U370 ( .A1(n601), .A2(n600), .ZN(n602) );
  AND2_X1 U370bar ( .A1(n601bar), .A2(n600bar), .ZN(n602bar);
  OR2_X1 U371 ( .A1(n820), .A2(n785), .ZN(n600) );
  AND2_X1 U371bar ( .A1(n820bar), .A2(n785bar), .ZN(n600bar);
  OR2_X1 U372 ( .A1(n599), .A2(n598), .ZN(n785) );
  AND2_X1 U372bar ( .A1(n599bar), .A2(n598bar), .ZN(n785bar);
  OR2_X1 U373 ( .A1(n597), .A2(n596), .ZN(n598) );
  AND2_X1 U373bar ( .A1(n597bar), .A2(n596bar), .ZN(n598bar);
  OR2_X1 U374 ( .A1(n595), .A2(n594), .ZN(n596) );
  AND2_X1 U374bar ( .A1(n595bar), .A2(n594bar), .ZN(n596bar);
  OR2_X1 U375 ( .A1(in[135]), .A2(in[104]), .ZN(n594) );
  AND2_X1 U375bar ( .A1(inbar[135]), .A2(inbar[104]), .ZN(n594bar);
  OR2_X1 U376 ( .A1(in[188]), .A2(in[178]), .ZN(n595) );
  AND2_X1 U376bar ( .A1(inbar[188]), .A2(inbar[178]), .ZN(n595bar);
  OR2_X1 U377 ( .A1(n593), .A2(n592), .ZN(n597) );
  AND2_X1 U377bar ( .A1(n593bar), .A2(n592bar), .ZN(n597bar);
  OR2_X1 U378 ( .A1(in[217]), .A2(in[194]), .ZN(n592) );
  AND2_X1 U378bar ( .A1(inbar[217]), .A2(inbar[194]), .ZN(n592bar);
  OR2_X1 U379 ( .A1(in[237]), .A2(in[218]), .ZN(n593) );
  AND2_X1 U379bar ( .A1(inbar[237]), .A2(inbar[218]), .ZN(n593bar);
  OR2_X1 U380 ( .A1(n591), .A2(n590), .ZN(n599) );
  AND2_X1 U380bar ( .A1(n591bar), .A2(n590bar), .ZN(n599bar);
  OR2_X1 U381 ( .A1(n589), .A2(n588), .ZN(n590) );
  AND2_X1 U381bar ( .A1(n589bar), .A2(n588bar), .ZN(n590bar);
  OR2_X1 U382 ( .A1(in_2), .A2(in_10), .ZN(n588) );
  AND2_X1 U382bar ( .A1(in_2bar), .A2(in_10bar), .ZN(n588bar);
  OR2_X1 U383 ( .A1(in_47), .A2(in_22), .ZN(n589) );
  AND2_X1 U383bar ( .A1(in_47bar), .A2(in_22bar), .ZN(n589bar);
  OR2_X1 U384 ( .A1(n587), .A2(n586), .ZN(n591) );
  AND2_X1 U384bar ( .A1(n587bar), .A2(n586bar), .ZN(n591bar);
  OR2_X1 U385 ( .A1(in_56), .A2(in_54), .ZN(n586) );
  AND2_X1 U385bar ( .A1(in_56bar), .A2(in_54bar), .ZN(n586bar);
  OR2_X1 U386 ( .A1(in_63), .A2(in_61), .ZN(n587) );
  AND2_X1 U386bar ( .A1(in_63bar), .A2(in_61bar), .ZN(n587bar);
  OR2_X1 U387 ( .A1(n585), .A2(n584), .ZN(n820) );
  AND2_X1 U387bar ( .A1(n585bar), .A2(n584bar), .ZN(n820bar);
  OR2_X1 U388 ( .A1(n583), .A2(n582), .ZN(n584) );
  AND2_X1 U388bar ( .A1(n583bar), .A2(n582bar), .ZN(n584bar);
  OR2_X1 U389 ( .A1(n581), .A2(n580), .ZN(n582) );
  AND2_X1 U389bar ( .A1(n581bar), .A2(n580bar), .ZN(n582bar);
  OR2_X1 U390 ( .A1(in[158]), .A2(in[142]), .ZN(n580) );
  AND2_X1 U390bar ( .A1(inbar[158]), .A2(inbar[142]), .ZN(n580bar);
  OR2_X1 U391 ( .A1(in[175]), .A2(in[164]), .ZN(n581) );
  AND2_X1 U391bar ( .A1(inbar[175]), .A2(inbar[164]), .ZN(n581bar);
  OR2_X1 U392 ( .A1(n579), .A2(n578), .ZN(n583) );
  AND2_X1 U392bar ( .A1(n579bar), .A2(n578bar), .ZN(n583bar);
  OR2_X1 U393 ( .A1(in[228]), .A2(in[204]), .ZN(n578) );
  AND2_X1 U393bar ( .A1(inbar[228]), .A2(inbar[204]), .ZN(n578bar);
  OR2_X1 U394 ( .A1(in[91]), .A2(in[87]), .ZN(n579) );
  AND2_X1 U394bar ( .A1(inbar[91]), .A2(inbar[87]), .ZN(n579bar);
  OR2_X1 U395 ( .A1(n577), .A2(n576), .ZN(n585) );
  AND2_X1 U395bar ( .A1(n577bar), .A2(n576bar), .ZN(n585bar);
  OR2_X1 U396 ( .A1(n575), .A2(n574), .ZN(n576) );
  AND2_X1 U396bar ( .A1(n575bar), .A2(n574bar), .ZN(n576bar);
  OR2_X1 U397 ( .A1(in_21), .A2(in_11), .ZN(n574) );
  AND2_X1 U397bar ( .A1(in_21bar), .A2(in_11bar), .ZN(n574bar);
  OR2_X1 U398 ( .A1(in_5), .A2(in_3), .ZN(n575) );
  AND2_X1 U398bar ( .A1(in_5bar), .A2(in_3bar), .ZN(n575bar);
  OR2_X1 U399 ( .A1(n573), .A2(n572), .ZN(n577) );
  AND2_X1 U399bar ( .A1(n573bar), .A2(n572bar), .ZN(n577bar);
  OR2_X1 U400 ( .A1(in_68), .A2(in_64), .ZN(n572) );
  AND2_X1 U400bar ( .A1(in_68bar), .A2(in_64bar), .ZN(n572bar);
  OR2_X1 U401 ( .A1(in_76), .A2(in_73), .ZN(n573) );
  AND2_X1 U401bar ( .A1(in_76bar), .A2(in_73bar), .ZN(n573bar);
  OR2_X1 U402 ( .A1(n778), .A2(n571), .ZN(n601) );
  AND2_X1 U402bar ( .A1(n778bar), .A2(n571bar), .ZN(n601bar);
  OR2_X1 U403 ( .A1(in[100]), .A2(n965), .ZN(n571) );
  AND2_X1 U403bar ( .A1(inbar[100]), .A2(n965bar), .ZN(n571bar);
  OR2_X1 U404 ( .A1(n570), .A2(n569), .ZN(n965) );
  AND2_X1 U404bar ( .A1(n570bar), .A2(n569bar), .ZN(n965bar);
  OR2_X1 U405 ( .A1(n568), .A2(n567), .ZN(n569) );
  AND2_X1 U405bar ( .A1(n568bar), .A2(n567bar), .ZN(n569bar);
  OR2_X1 U406 ( .A1(n566), .A2(n565), .ZN(n567) );
  AND2_X1 U406bar ( .A1(n566bar), .A2(n565bar), .ZN(n567bar);
  OR2_X1 U407 ( .A1(n817), .A2(n750), .ZN(n565) );
  AND2_X1 U407bar ( .A1(n817bar), .A2(n750bar), .ZN(n565bar);
  OR2_X1 U408 ( .A1(n564), .A2(n563), .ZN(n750) );
  AND2_X1 U408bar ( .A1(n564bar), .A2(n563bar), .ZN(n750bar);
  OR2_X1 U409 ( .A1(n562), .A2(n561), .ZN(n563) );
  AND2_X1 U409bar ( .A1(n562bar), .A2(n561bar), .ZN(n563bar);
  OR2_X1 U410 ( .A1(n560), .A2(n559), .ZN(n561) );
  AND2_X1 U410bar ( .A1(n560bar), .A2(n559bar), .ZN(n561bar);
  OR2_X1 U411 ( .A1(in[119]), .A2(in[103]), .ZN(n559) );
  AND2_X1 U411bar ( .A1(inbar[119]), .A2(inbar[103]), .ZN(n559bar);
  OR2_X1 U412 ( .A1(in[137]), .A2(in[133]), .ZN(n560) );
  AND2_X1 U412bar ( .A1(inbar[137]), .A2(inbar[133]), .ZN(n560bar);
  OR2_X1 U413 ( .A1(n558), .A2(n557), .ZN(n562) );
  AND2_X1 U413bar ( .A1(n558bar), .A2(n557bar), .ZN(n562bar);
  OR2_X1 U414 ( .A1(in[176]), .A2(in[173]), .ZN(n557) );
  AND2_X1 U414bar ( .A1(inbar[176]), .A2(inbar[173]), .ZN(n557bar);
  OR2_X1 U415 ( .A1(in[210]), .A2(in[181]), .ZN(n558) );
  AND2_X1 U415bar ( .A1(inbar[210]), .A2(inbar[181]), .ZN(n558bar);
  OR2_X1 U416 ( .A1(n556), .A2(n555), .ZN(n564) );
  AND2_X1 U416bar ( .A1(n556bar), .A2(n555bar), .ZN(n564bar);
  OR2_X1 U417 ( .A1(n554), .A2(n553), .ZN(n555) );
  AND2_X1 U417bar ( .A1(n554bar), .A2(n553bar), .ZN(n555bar);
  OR2_X1 U418 ( .A1(in_13), .A2(in[234]), .ZN(n553) );
  AND2_X1 U418bar ( .A1(in_13bar), .A2(inbar[234]), .ZN(n553bar);
  OR2_X1 U419 ( .A1(in_38), .A2(in_32), .ZN(n554) );
  AND2_X1 U419bar ( .A1(in_38bar), .A2(in_32bar), .ZN(n554bar);
  OR2_X1 U420 ( .A1(n552), .A2(n551), .ZN(n556) );
  AND2_X1 U420bar ( .A1(n552bar), .A2(n551bar), .ZN(n556bar);
  OR2_X1 U421 ( .A1(in_42), .A2(in_41), .ZN(n551) );
  AND2_X1 U421bar ( .A1(in_42bar), .A2(in_41bar), .ZN(n551bar);
  OR2_X1 U422 ( .A1(in_7), .A2(in_49), .ZN(n552) );
  AND2_X1 U422bar ( .A1(in_7bar), .A2(in_49bar), .ZN(n552bar);
  OR2_X1 U423 ( .A1(n550), .A2(n549), .ZN(n817) );
  AND2_X1 U423bar ( .A1(n550bar), .A2(n549bar), .ZN(n817bar);
  OR2_X1 U424 ( .A1(n548), .A2(n547), .ZN(n549) );
  AND2_X1 U424bar ( .A1(n548bar), .A2(n547bar), .ZN(n549bar);
  OR2_X1 U425 ( .A1(n546), .A2(n545), .ZN(n547) );
  AND2_X1 U425bar ( .A1(n546bar), .A2(n545bar), .ZN(n547bar);
  OR2_X1 U426 ( .A1(in[159]), .A2(in[105]), .ZN(n545) );
  AND2_X1 U426bar ( .A1(inbar[159]), .A2(inbar[105]), .ZN(n545bar);
  OR2_X1 U427 ( .A1(in[206]), .A2(in[183]), .ZN(n546) );
  AND2_X1 U427bar ( .A1(inbar[206]), .A2(inbar[183]), .ZN(n546bar);
  OR2_X1 U428 ( .A1(n544), .A2(n543), .ZN(n548) );
  AND2_X1 U428bar ( .A1(n544bar), .A2(n543bar), .ZN(n548bar);
  OR2_X1 U429 ( .A1(in[229]), .A2(in[219]), .ZN(n543) );
  AND2_X1 U429bar ( .A1(inbar[229]), .A2(inbar[219]), .ZN(n543bar);
  OR2_X1 U430 ( .A1(in[235]), .A2(in[232]), .ZN(n544) );
  AND2_X1 U430bar ( .A1(inbar[235]), .A2(inbar[232]), .ZN(n544bar);
  OR2_X1 U431 ( .A1(n542), .A2(n541), .ZN(n550) );
  AND2_X1 U431bar ( .A1(n542bar), .A2(n541bar), .ZN(n550bar);
  OR2_X1 U432 ( .A1(n540), .A2(n539), .ZN(n541) );
  AND2_X1 U432bar ( .A1(n540bar), .A2(n539bar), .ZN(n541bar);
  OR2_X1 U433 ( .A1(in[249]), .A2(in[242]), .ZN(n539) );
  AND2_X1 U433bar ( .A1(inbar[249]), .A2(inbar[242]), .ZN(n539bar);
  OR2_X1 U434 ( .A1(in[89]), .A2(in[254]), .ZN(n540) );
  AND2_X1 U434bar ( .A1(inbar[89]), .A2(inbar[254]), .ZN(n540bar);
  OR2_X1 U435 ( .A1(n538), .A2(n537), .ZN(n542) );
  AND2_X1 U435bar ( .A1(n538bar), .A2(n537bar), .ZN(n542bar);
  OR2_X1 U436 ( .A1(in_14), .A2(in[99]), .ZN(n537) );
  AND2_X1 U436bar ( .A1(in_14bar), .A2(inbar[99]), .ZN(n537bar);
  OR2_X1 U437 ( .A1(in_60), .A2(in_18), .ZN(n538) );
  AND2_X1 U437bar ( .A1(in_60bar), .A2(in_18bar), .ZN(n538bar);
  OR2_X1 U438 ( .A1(in[113]), .A2(n763), .ZN(n566) );
  AND2_X1 U438bar ( .A1(inbar[113]), .A2(n763bar), .ZN(n566bar);
  OR2_X1 U439 ( .A1(n536), .A2(n535), .ZN(n763) );
  AND2_X1 U439bar ( .A1(n536bar), .A2(n535bar), .ZN(n763bar);
  OR2_X1 U440 ( .A1(n534), .A2(n533), .ZN(n535) );
  AND2_X1 U440bar ( .A1(n534bar), .A2(n533bar), .ZN(n535bar);
  OR2_X1 U441 ( .A1(n532), .A2(n531), .ZN(n533) );
  AND2_X1 U441bar ( .A1(n532bar), .A2(n531bar), .ZN(n533bar);
  OR2_X1 U442 ( .A1(in[115]), .A2(in[110]), .ZN(n531) );
  AND2_X1 U442bar ( .A1(inbar[115]), .A2(inbar[110]), .ZN(n531bar);
  OR2_X1 U443 ( .A1(in[125]), .A2(in[117]), .ZN(n532) );
  AND2_X1 U443bar ( .A1(inbar[125]), .A2(inbar[117]), .ZN(n532bar);
  OR2_X1 U444 ( .A1(n530), .A2(n529), .ZN(n534) );
  AND2_X1 U444bar ( .A1(n530bar), .A2(n529bar), .ZN(n534bar);
  OR2_X1 U445 ( .A1(in[180]), .A2(in[128]), .ZN(n529) );
  AND2_X1 U445bar ( .A1(inbar[180]), .A2(inbar[128]), .ZN(n529bar);
  OR2_X1 U446 ( .A1(in[205]), .A2(in[201]), .ZN(n530) );
  AND2_X1 U446bar ( .A1(inbar[205]), .A2(inbar[201]), .ZN(n530bar);
  OR2_X1 U447 ( .A1(n528), .A2(n527), .ZN(n536) );
  AND2_X1 U447bar ( .A1(n528bar), .A2(n527bar), .ZN(n536bar);
  OR2_X1 U448 ( .A1(n526), .A2(n525), .ZN(n527) );
  AND2_X1 U448bar ( .A1(n526bar), .A2(n525bar), .ZN(n527bar);
  OR2_X1 U449 ( .A1(in[244]), .A2(in[239]), .ZN(n525) );
  AND2_X1 U449bar ( .A1(inbar[244]), .A2(inbar[239]), .ZN(n525bar);
  OR2_X1 U450 ( .A1(in[95]), .A2(in[83]), .ZN(n526) );
  AND2_X1 U450bar ( .A1(inbar[95]), .A2(inbar[83]), .ZN(n526bar);
  OR2_X1 U451 ( .A1(n524), .A2(n523), .ZN(n528) );
  AND2_X1 U451bar ( .A1(n524bar), .A2(n523bar), .ZN(n528bar);
  OR2_X1 U452 ( .A1(in_24), .A2(in[97]), .ZN(n523) );
  AND2_X1 U452bar ( .A1(in_24bar), .A2(inbar[97]), .ZN(n523bar);
  OR2_X1 U453 ( .A1(in_33), .A2(in_27), .ZN(n524) );
  AND2_X1 U453bar ( .A1(in_33bar), .A2(in_27bar), .ZN(n524bar);
  OR2_X1 U454 ( .A1(n522), .A2(n521), .ZN(n568) );
  AND2_X1 U454bar ( .A1(n522bar), .A2(n521bar), .ZN(n568bar);
  OR2_X1 U455 ( .A1(in[145]), .A2(in[126]), .ZN(n521) );
  AND2_X1 U455bar ( .A1(inbar[145]), .A2(inbar[126]), .ZN(n521bar);
  OR2_X1 U456 ( .A1(in[169]), .A2(n520), .ZN(n522) );
  AND2_X1 U456bar ( .A1(inbar[169]), .A2(n520bar), .ZN(n522bar);
  OR2_X1 U457 ( .A1(in[221]), .A2(in[172]), .ZN(n520) );
  AND2_X1 U457bar ( .A1(inbar[221]), .A2(inbar[172]), .ZN(n520bar);
  OR2_X1 U458 ( .A1(n519), .A2(n518), .ZN(n570) );
  AND2_X1 U458bar ( .A1(n519bar), .A2(n518bar), .ZN(n570bar);
  OR2_X1 U459 ( .A1(n517), .A2(n516), .ZN(n518) );
  AND2_X1 U459bar ( .A1(n517bar), .A2(n516bar), .ZN(n518bar);
  OR2_X1 U460 ( .A1(in[241]), .A2(in[224]), .ZN(n516) );
  AND2_X1 U460bar ( .A1(inbar[241]), .A2(inbar[224]), .ZN(n516bar);
  OR2_X1 U461 ( .A1(in[86]), .A2(n515), .ZN(n517) );
  AND2_X1 U461bar ( .A1(inbar[86]), .A2(n515bar), .ZN(n517bar);
  OR2_X1 U462 ( .A1(in_43), .A2(in_34), .ZN(n515) );
  AND2_X1 U462bar ( .A1(in_43bar), .A2(in_34bar), .ZN(n515bar);
  OR2_X1 U463 ( .A1(n514), .A2(n513), .ZN(n519) );
  AND2_X1 U463bar ( .A1(n514bar), .A2(n513bar), .ZN(n519bar);
  OR2_X1 U464 ( .A1(in_65), .A2(in_51), .ZN(n513) );
  AND2_X1 U464bar ( .A1(in_65bar), .A2(in_51bar), .ZN(n513bar);
  OR2_X1 U465 ( .A1(in_75), .A2(n512), .ZN(n514) );
  AND2_X1 U465bar ( .A1(in_75bar), .A2(n512bar), .ZN(n514bar);
  OR2_X1 U466 ( .A1(in_81), .A2(in_77), .ZN(n512) );
  AND2_X1 U466bar ( .A1(in_81bar), .A2(in_77bar), .ZN(n512bar);
  OR2_X1 U467 ( .A1(n511), .A2(n510), .ZN(n778) );
  AND2_X1 U467bar ( .A1(n511bar), .A2(n510bar), .ZN(n778bar);
  OR2_X1 U468 ( .A1(n509), .A2(n508), .ZN(n510) );
  AND2_X1 U468bar ( .A1(n509bar), .A2(n508bar), .ZN(n510bar);
  OR2_X1 U469 ( .A1(n507), .A2(n506), .ZN(n508) );
  AND2_X1 U469bar ( .A1(n507bar), .A2(n506bar), .ZN(n508bar);
  OR2_X1 U470 ( .A1(in[107]), .A2(in[101]), .ZN(n506) );
  AND2_X1 U470bar ( .A1(inbar[107]), .A2(inbar[101]), .ZN(n506bar);
  OR2_X1 U471 ( .A1(in[139]), .A2(in[132]), .ZN(n507) );
  AND2_X1 U471bar ( .A1(inbar[139]), .A2(inbar[132]), .ZN(n507bar);
  OR2_X1 U472 ( .A1(n505), .A2(n504), .ZN(n509) );
  AND2_X1 U472bar ( .A1(n505bar), .A2(n504bar), .ZN(n509bar);
  OR2_X1 U473 ( .A1(in[146]), .A2(in[141]), .ZN(n504) );
  AND2_X1 U473bar ( .A1(inbar[146]), .A2(inbar[141]), .ZN(n504bar);
  OR2_X1 U474 ( .A1(in[203]), .A2(in[179]), .ZN(n505) );
  AND2_X1 U474bar ( .A1(inbar[203]), .A2(inbar[179]), .ZN(n505bar);
  OR2_X1 U475 ( .A1(n503), .A2(n502), .ZN(n511) );
  AND2_X1 U475bar ( .A1(n503bar), .A2(n502bar), .ZN(n511bar);
  OR2_X1 U476 ( .A1(n501), .A2(n500), .ZN(n502) );
  AND2_X1 U476bar ( .A1(n501bar), .A2(n500bar), .ZN(n502bar);
  OR2_X1 U477 ( .A1(in[243]), .A2(in[222]), .ZN(n500) );
  AND2_X1 U477bar ( .A1(inbar[243]), .A2(inbar[222]), .ZN(n500bar);
  OR2_X1 U478 ( .A1(in[251]), .A2(in[250]), .ZN(n501) );
  AND2_X1 U478bar ( .A1(inbar[251]), .A2(inbar[250]), .ZN(n501bar);
  OR2_X1 U479 ( .A1(n499), .A2(n498), .ZN(n503) );
  AND2_X1 U479bar ( .A1(n499bar), .A2(n498bar), .ZN(n503bar);
  OR2_X1 U480 ( .A1(in_37), .A2(in_19), .ZN(n498) );
  AND2_X1 U480bar ( .A1(in_37bar), .A2(in_19bar), .ZN(n498bar);
  OR2_X1 U481 ( .A1(in_78), .A2(in_6), .ZN(n499) );
  AND2_X1 U481bar ( .A1(in_78bar), .A2(in_6bar), .ZN(n499bar);
  OR2_X1 U482 ( .A1(n497), .A2(n496), .ZN(n603) );
  AND2_X1 U482bar ( .A1(n497bar), .A2(n496bar), .ZN(n603bar);
  OR2_X1 U483 ( .A1(in[112]), .A2(in[102]), .ZN(n496) );
  AND2_X1 U483bar ( .A1(inbar[112]), .A2(inbar[102]), .ZN(n496bar);
  OR2_X1 U484 ( .A1(in[123]), .A2(n495), .ZN(n497) );
  AND2_X1 U484bar ( .A1(inbar[123]), .A2(n495bar), .ZN(n497bar);
  OR2_X1 U485 ( .A1(in[143]), .A2(in[130]), .ZN(n495) );
  AND2_X1 U485bar ( .A1(inbar[143]), .A2(inbar[130]), .ZN(n495bar);
  OR2_X1 U486 ( .A1(n494), .A2(n493), .ZN(n605) );
  AND2_X1 U486bar ( .A1(n494bar), .A2(n493bar), .ZN(n605bar);
  OR2_X1 U487 ( .A1(n492), .A2(n491), .ZN(n493) );
  AND2_X1 U487bar ( .A1(n492bar), .A2(n491bar), .ZN(n493bar);
  OR2_X1 U488 ( .A1(in[216]), .A2(in[213]), .ZN(n491) );
  AND2_X1 U488bar ( .A1(inbar[216]), .A2(inbar[213]), .ZN(n491bar);
  OR2_X1 U489 ( .A1(in[227]), .A2(n490), .ZN(n492) );
  AND2_X1 U489bar ( .A1(inbar[227]), .A2(n490bar), .ZN(n492bar);
  OR2_X1 U490 ( .A1(in_0), .A2(in[248]), .ZN(n490) );
  AND2_X1 U490bar ( .A1(in_0bar), .A2(inbar[248]), .ZN(n490bar);
  OR2_X1 U491 ( .A1(n489), .A2(n488), .ZN(n494) );
  AND2_X1 U491bar ( .A1(n489bar), .A2(n488bar), .ZN(n494bar);
  OR2_X1 U492 ( .A1(in_46), .A2(in_44), .ZN(n488) );
  AND2_X1 U492bar ( .A1(in_46bar), .A2(in_44bar), .ZN(n488bar);
  OR2_X1 U493 ( .A1(in_50), .A2(n487), .ZN(n489) );
  AND2_X1 U493bar ( .A1(in_50bar), .A2(n487bar), .ZN(n489bar);
  OR2_X1 U494 ( .A1(in_9), .A2(in_80), .ZN(n487) );
  AND2_X1 U494bar ( .A1(in_9bar), .A2(in_80bar), .ZN(n487bar);
endmodule




module sBox_1 ( in, out );
  input [7:0] in;
  //input_done

  output [7:0] out;
  //output_done

  wire   [255:0] decodeOut;
  //wire_done

  decode_1 dec ( .in(in), .out(decodeOut) );
  encode_1 enc ( .in(decodeOut), .out(out) );
endmodule


module CD2_5 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  //ooutput_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_6 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_7 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_8 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD4_3 ( a, b, y );
  input [3:0] a;
  input [3:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  //input_done

  output [15:0] y;
  reg [15:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]);
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]);
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]);
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]);
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]);
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]);
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]);
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]);
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]);
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]);
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]);
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]);
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]);
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]);
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]);
endmodule




module CD4_4 ( a, b, y );
  input [3:0] a;
  input [3:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  //input_done

  output [15:0] y;
  reg [15:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]);
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]);
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]);
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]);
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]);
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]);
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]);
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]);
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]);
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]);
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]);
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]);
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]);
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]);
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]);
endmodule




module CD16_2 ( a, b, y );
  input [15:0] a;
  input [15:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign abar[8] = ~a[8];
  assign abar[9] = ~a[9];
  assign abar[10] = ~a[10];
  assign abar[11] = ~a[11];
  assign abar[12] = ~a[12];
  assign abar[13] = ~a[13];
  assign abar[14] = ~a[14];
  assign abar[15] = ~a[15];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign bbar[8] = ~b[8];
  assign bbar[9] = ~b[9];
  assign bbar[10] = ~b[10];
  assign bbar[11] = ~b[11];
  assign bbar[12] = ~b[12];
  assign bbar[13] = ~b[13];
  assign bbar[14] = ~b[14];
  assign bbar[15] = ~b[15];
  //input_done

  output [255:0] y;
  reg [255:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[9]), .A2(a[0]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[9]), .A2(abar[0]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[3]), .A2(a[6]), .ZN(y[99]) );
  OR2_X1 U2bar ( .A1(bbar[3]), .A2(abar[6]), .ZN(ybar[99]);
  AND2_X1 U3 ( .A1(b[2]), .A2(a[6]), .ZN(y[98]) );
  OR2_X1 U3bar ( .A1(bbar[2]), .A2(abar[6]), .ZN(ybar[98]);
  AND2_X1 U4 ( .A1(b[1]), .A2(a[6]), .ZN(y[97]) );
  OR2_X1 U4bar ( .A1(bbar[1]), .A2(abar[6]), .ZN(ybar[97]);
  AND2_X1 U5 ( .A1(b[0]), .A2(a[6]), .ZN(y[96]) );
  OR2_X1 U5bar ( .A1(bbar[0]), .A2(abar[6]), .ZN(ybar[96]);
  AND2_X1 U6 ( .A1(b[15]), .A2(a[5]), .ZN(y[95]) );
  OR2_X1 U6bar ( .A1(bbar[15]), .A2(abar[5]), .ZN(ybar[95]);
  AND2_X1 U7 ( .A1(b[14]), .A2(a[5]), .ZN(y[94]) );
  OR2_X1 U7bar ( .A1(bbar[14]), .A2(abar[5]), .ZN(ybar[94]);
  AND2_X1 U8 ( .A1(b[13]), .A2(a[5]), .ZN(y[93]) );
  OR2_X1 U8bar ( .A1(bbar[13]), .A2(abar[5]), .ZN(ybar[93]);
  AND2_X1 U9 ( .A1(b[12]), .A2(a[5]), .ZN(y[92]) );
  OR2_X1 U9bar ( .A1(bbar[12]), .A2(abar[5]), .ZN(ybar[92]);
  AND2_X1 U10 ( .A1(b[11]), .A2(a[5]), .ZN(y[91]) );
  OR2_X1 U10bar ( .A1(bbar[11]), .A2(abar[5]), .ZN(ybar[91]);
  AND2_X1 U11 ( .A1(b[10]), .A2(a[5]), .ZN(y[90]) );
  OR2_X1 U11bar ( .A1(bbar[10]), .A2(abar[5]), .ZN(ybar[90]);
  AND2_X1 U12 ( .A1(b[8]), .A2(a[0]), .ZN(y[8]) );
  OR2_X1 U12bar ( .A1(bbar[8]), .A2(abar[0]), .ZN(ybar[8]);
  AND2_X1 U13 ( .A1(a[5]), .A2(b[9]), .ZN(y[89]) );
  OR2_X1 U13bar ( .A1(abar[5]), .A2(bbar[9]), .ZN(ybar[89]);
  AND2_X1 U14 ( .A1(b[8]), .A2(a[5]), .ZN(y[88]) );
  OR2_X1 U14bar ( .A1(bbar[8]), .A2(abar[5]), .ZN(ybar[88]);
  AND2_X1 U15 ( .A1(b[7]), .A2(a[5]), .ZN(y[87]) );
  OR2_X1 U15bar ( .A1(bbar[7]), .A2(abar[5]), .ZN(ybar[87]);
  AND2_X1 U16 ( .A1(b[6]), .A2(a[5]), .ZN(y[86]) );
  OR2_X1 U16bar ( .A1(bbar[6]), .A2(abar[5]), .ZN(ybar[86]);
  AND2_X1 U17 ( .A1(b[5]), .A2(a[5]), .ZN(y[85]) );
  OR2_X1 U17bar ( .A1(bbar[5]), .A2(abar[5]), .ZN(ybar[85]);
  AND2_X1 U18 ( .A1(b[4]), .A2(a[5]), .ZN(y[84]) );
  OR2_X1 U18bar ( .A1(bbar[4]), .A2(abar[5]), .ZN(ybar[84]);
  AND2_X1 U19 ( .A1(a[5]), .A2(b[3]), .ZN(y[83]) );
  OR2_X1 U19bar ( .A1(abar[5]), .A2(bbar[3]), .ZN(ybar[83]);
  AND2_X1 U20 ( .A1(a[5]), .A2(b[2]), .ZN(y[82]) );
  OR2_X1 U20bar ( .A1(abar[5]), .A2(bbar[2]), .ZN(ybar[82]);
  AND2_X1 U21 ( .A1(a[5]), .A2(b[1]), .ZN(y[81]) );
  OR2_X1 U21bar ( .A1(abar[5]), .A2(bbar[1]), .ZN(ybar[81]);
  AND2_X1 U22 ( .A1(a[5]), .A2(b[0]), .ZN(y[80]) );
  OR2_X1 U22bar ( .A1(abar[5]), .A2(bbar[0]), .ZN(ybar[80]);
  AND2_X1 U23 ( .A1(b[7]), .A2(a[0]), .ZN(y[7]) );
  OR2_X1 U23bar ( .A1(bbar[7]), .A2(abar[0]), .ZN(ybar[7]);
  AND2_X1 U24 ( .A1(a[4]), .A2(b[15]), .ZN(y[79]) );
  OR2_X1 U24bar ( .A1(abar[4]), .A2(bbar[15]), .ZN(ybar[79]);
  AND2_X1 U25 ( .A1(a[4]), .A2(b[14]), .ZN(y[78]) );
  OR2_X1 U25bar ( .A1(abar[4]), .A2(bbar[14]), .ZN(ybar[78]);
  AND2_X1 U26 ( .A1(a[4]), .A2(b[13]), .ZN(y[77]) );
  OR2_X1 U26bar ( .A1(abar[4]), .A2(bbar[13]), .ZN(ybar[77]);
  AND2_X1 U27 ( .A1(a[4]), .A2(b[12]), .ZN(y[76]) );
  OR2_X1 U27bar ( .A1(abar[4]), .A2(bbar[12]), .ZN(ybar[76]);
  AND2_X1 U28 ( .A1(a[4]), .A2(b[11]), .ZN(y[75]) );
  OR2_X1 U28bar ( .A1(abar[4]), .A2(bbar[11]), .ZN(ybar[75]);
  AND2_X1 U29 ( .A1(a[4]), .A2(b[10]), .ZN(y[74]) );
  OR2_X1 U29bar ( .A1(abar[4]), .A2(bbar[10]), .ZN(ybar[74]);
  AND2_X1 U30 ( .A1(a[4]), .A2(b[9]), .ZN(y[73]) );
  OR2_X1 U30bar ( .A1(abar[4]), .A2(bbar[9]), .ZN(ybar[73]);
  AND2_X1 U31 ( .A1(a[4]), .A2(b[8]), .ZN(y[72]) );
  OR2_X1 U31bar ( .A1(abar[4]), .A2(bbar[8]), .ZN(ybar[72]);
  AND2_X1 U32 ( .A1(a[4]), .A2(b[7]), .ZN(y[71]) );
  OR2_X1 U32bar ( .A1(abar[4]), .A2(bbar[7]), .ZN(ybar[71]);
  AND2_X1 U33 ( .A1(a[4]), .A2(b[6]), .ZN(y[70]) );
  OR2_X1 U33bar ( .A1(abar[4]), .A2(bbar[6]), .ZN(ybar[70]);
  AND2_X1 U34 ( .A1(b[6]), .A2(a[0]), .ZN(y[6]) );
  OR2_X1 U34bar ( .A1(bbar[6]), .A2(abar[0]), .ZN(ybar[6]);
  AND2_X1 U35 ( .A1(a[4]), .A2(b[5]), .ZN(y[69]) );
  OR2_X1 U35bar ( .A1(abar[4]), .A2(bbar[5]), .ZN(ybar[69]);
  AND2_X1 U36 ( .A1(a[4]), .A2(b[4]), .ZN(y[68]) );
  OR2_X1 U36bar ( .A1(abar[4]), .A2(bbar[4]), .ZN(ybar[68]);
  AND2_X1 U37 ( .A1(a[4]), .A2(b[3]), .ZN(y[67]) );
  OR2_X1 U37bar ( .A1(abar[4]), .A2(bbar[3]), .ZN(ybar[67]);
  AND2_X1 U38 ( .A1(a[4]), .A2(b[2]), .ZN(y[66]) );
  OR2_X1 U38bar ( .A1(abar[4]), .A2(bbar[2]), .ZN(ybar[66]);
  AND2_X1 U39 ( .A1(a[4]), .A2(b[1]), .ZN(y[65]) );
  OR2_X1 U39bar ( .A1(abar[4]), .A2(bbar[1]), .ZN(ybar[65]);
  AND2_X1 U40 ( .A1(a[4]), .A2(b[0]), .ZN(y[64]) );
  OR2_X1 U40bar ( .A1(abar[4]), .A2(bbar[0]), .ZN(ybar[64]);
  AND2_X1 U41 ( .A1(a[3]), .A2(b[15]), .ZN(y[63]) );
  OR2_X1 U41bar ( .A1(abar[3]), .A2(bbar[15]), .ZN(ybar[63]);
  AND2_X1 U42 ( .A1(a[3]), .A2(b[14]), .ZN(y[62]) );
  OR2_X1 U42bar ( .A1(abar[3]), .A2(bbar[14]), .ZN(ybar[62]);
  AND2_X1 U43 ( .A1(a[3]), .A2(b[13]), .ZN(y[61]) );
  OR2_X1 U43bar ( .A1(abar[3]), .A2(bbar[13]), .ZN(ybar[61]);
  AND2_X1 U44 ( .A1(a[3]), .A2(b[12]), .ZN(y[60]) );
  OR2_X1 U44bar ( .A1(abar[3]), .A2(bbar[12]), .ZN(ybar[60]);
  AND2_X1 U45 ( .A1(b[5]), .A2(a[0]), .ZN(y[5]) );
  OR2_X1 U45bar ( .A1(bbar[5]), .A2(abar[0]), .ZN(ybar[5]);
  AND2_X1 U46 ( .A1(a[3]), .A2(b[11]), .ZN(y[59]) );
  OR2_X1 U46bar ( .A1(abar[3]), .A2(bbar[11]), .ZN(ybar[59]);
  AND2_X1 U47 ( .A1(a[3]), .A2(b[10]), .ZN(y[58]) );
  OR2_X1 U47bar ( .A1(abar[3]), .A2(bbar[10]), .ZN(ybar[58]);
  AND2_X1 U48 ( .A1(a[3]), .A2(b[9]), .ZN(y[57]) );
  OR2_X1 U48bar ( .A1(abar[3]), .A2(bbar[9]), .ZN(ybar[57]);
  AND2_X1 U49 ( .A1(a[3]), .A2(b[8]), .ZN(y[56]) );
  OR2_X1 U49bar ( .A1(abar[3]), .A2(bbar[8]), .ZN(ybar[56]);
  AND2_X1 U50 ( .A1(a[3]), .A2(b[7]), .ZN(y[55]) );
  OR2_X1 U50bar ( .A1(abar[3]), .A2(bbar[7]), .ZN(ybar[55]);
  AND2_X1 U51 ( .A1(a[3]), .A2(b[6]), .ZN(y[54]) );
  OR2_X1 U51bar ( .A1(abar[3]), .A2(bbar[6]), .ZN(ybar[54]);
  AND2_X1 U52 ( .A1(a[3]), .A2(b[5]), .ZN(y[53]) );
  OR2_X1 U52bar ( .A1(abar[3]), .A2(bbar[5]), .ZN(ybar[53]);
  AND2_X1 U53 ( .A1(a[3]), .A2(b[4]), .ZN(y[52]) );
  OR2_X1 U53bar ( .A1(abar[3]), .A2(bbar[4]), .ZN(ybar[52]);
  AND2_X1 U54 ( .A1(a[3]), .A2(b[3]), .ZN(y[51]) );
  OR2_X1 U54bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[51]);
  AND2_X1 U55 ( .A1(a[3]), .A2(b[2]), .ZN(y[50]) );
  OR2_X1 U55bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[50]);
  AND2_X1 U56 ( .A1(b[4]), .A2(a[0]), .ZN(y[4]) );
  OR2_X1 U56bar ( .A1(bbar[4]), .A2(abar[0]), .ZN(ybar[4]);
  AND2_X1 U57 ( .A1(a[3]), .A2(b[1]), .ZN(y[49]) );
  OR2_X1 U57bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[49]);
  AND2_X1 U58 ( .A1(a[3]), .A2(b[0]), .ZN(y[48]) );
  OR2_X1 U58bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[48]);
  AND2_X1 U59 ( .A1(a[2]), .A2(b[15]), .ZN(y[47]) );
  OR2_X1 U59bar ( .A1(abar[2]), .A2(bbar[15]), .ZN(ybar[47]);
  AND2_X1 U60 ( .A1(a[2]), .A2(b[14]), .ZN(y[46]) );
  OR2_X1 U60bar ( .A1(abar[2]), .A2(bbar[14]), .ZN(ybar[46]);
  AND2_X1 U61 ( .A1(a[2]), .A2(b[13]), .ZN(y[45]) );
  OR2_X1 U61bar ( .A1(abar[2]), .A2(bbar[13]), .ZN(ybar[45]);
  AND2_X1 U62 ( .A1(a[2]), .A2(b[12]), .ZN(y[44]) );
  OR2_X1 U62bar ( .A1(abar[2]), .A2(bbar[12]), .ZN(ybar[44]);
  AND2_X1 U63 ( .A1(a[2]), .A2(b[11]), .ZN(y[43]) );
  OR2_X1 U63bar ( .A1(abar[2]), .A2(bbar[11]), .ZN(ybar[43]);
  AND2_X1 U64 ( .A1(a[2]), .A2(b[10]), .ZN(y[42]) );
  OR2_X1 U64bar ( .A1(abar[2]), .A2(bbar[10]), .ZN(ybar[42]);
  AND2_X1 U65 ( .A1(a[2]), .A2(b[9]), .ZN(y[41]) );
  OR2_X1 U65bar ( .A1(abar[2]), .A2(bbar[9]), .ZN(ybar[41]);
  AND2_X1 U66 ( .A1(a[2]), .A2(b[8]), .ZN(y[40]) );
  OR2_X1 U66bar ( .A1(abar[2]), .A2(bbar[8]), .ZN(ybar[40]);
  AND2_X1 U67 ( .A1(b[3]), .A2(a[0]), .ZN(y[3]) );
  OR2_X1 U67bar ( .A1(bbar[3]), .A2(abar[0]), .ZN(ybar[3]);
  AND2_X1 U68 ( .A1(a[2]), .A2(b[7]), .ZN(y[39]) );
  OR2_X1 U68bar ( .A1(abar[2]), .A2(bbar[7]), .ZN(ybar[39]);
  AND2_X1 U69 ( .A1(a[2]), .A2(b[6]), .ZN(y[38]) );
  OR2_X1 U69bar ( .A1(abar[2]), .A2(bbar[6]), .ZN(ybar[38]);
  AND2_X1 U70 ( .A1(a[2]), .A2(b[5]), .ZN(y[37]) );
  OR2_X1 U70bar ( .A1(abar[2]), .A2(bbar[5]), .ZN(ybar[37]);
  AND2_X1 U71 ( .A1(a[2]), .A2(b[4]), .ZN(y[36]) );
  OR2_X1 U71bar ( .A1(abar[2]), .A2(bbar[4]), .ZN(ybar[36]);
  AND2_X1 U72 ( .A1(a[2]), .A2(b[3]), .ZN(y[35]) );
  OR2_X1 U72bar ( .A1(abar[2]), .A2(bbar[3]), .ZN(ybar[35]);
  AND2_X1 U73 ( .A1(a[2]), .A2(b[2]), .ZN(y[34]) );
  OR2_X1 U73bar ( .A1(abar[2]), .A2(bbar[2]), .ZN(ybar[34]);
  AND2_X1 U74 ( .A1(a[2]), .A2(b[1]), .ZN(y[33]) );
  OR2_X1 U74bar ( .A1(abar[2]), .A2(bbar[1]), .ZN(ybar[33]);
  AND2_X1 U75 ( .A1(a[2]), .A2(b[0]), .ZN(y[32]) );
  OR2_X1 U75bar ( .A1(abar[2]), .A2(bbar[0]), .ZN(ybar[32]);
  AND2_X1 U76 ( .A1(a[1]), .A2(b[15]), .ZN(y[31]) );
  OR2_X1 U76bar ( .A1(abar[1]), .A2(bbar[15]), .ZN(ybar[31]);
  AND2_X1 U77 ( .A1(a[1]), .A2(b[14]), .ZN(y[30]) );
  OR2_X1 U77bar ( .A1(abar[1]), .A2(bbar[14]), .ZN(ybar[30]);
  AND2_X1 U78 ( .A1(b[2]), .A2(a[0]), .ZN(y[2]) );
  OR2_X1 U78bar ( .A1(bbar[2]), .A2(abar[0]), .ZN(ybar[2]);
  AND2_X1 U79 ( .A1(a[1]), .A2(b[13]), .ZN(y[29]) );
  OR2_X1 U79bar ( .A1(abar[1]), .A2(bbar[13]), .ZN(ybar[29]);
  AND2_X1 U80 ( .A1(a[1]), .A2(b[12]), .ZN(y[28]) );
  OR2_X1 U80bar ( .A1(abar[1]), .A2(bbar[12]), .ZN(ybar[28]);
  AND2_X1 U81 ( .A1(a[1]), .A2(b[11]), .ZN(y[27]) );
  OR2_X1 U81bar ( .A1(abar[1]), .A2(bbar[11]), .ZN(ybar[27]);
  AND2_X1 U82 ( .A1(a[1]), .A2(b[10]), .ZN(y[26]) );
  OR2_X1 U82bar ( .A1(abar[1]), .A2(bbar[10]), .ZN(ybar[26]);
  AND2_X1 U83 ( .A1(a[1]), .A2(b[9]), .ZN(y[25]) );
  OR2_X1 U83bar ( .A1(abar[1]), .A2(bbar[9]), .ZN(ybar[25]);
  AND2_X1 U84 ( .A1(a[15]), .A2(b[15]), .ZN(y[255]) );
  OR2_X1 U84bar ( .A1(abar[15]), .A2(bbar[15]), .ZN(ybar[255]);
  AND2_X1 U85 ( .A1(a[15]), .A2(b[14]), .ZN(y[254]) );
  OR2_X1 U85bar ( .A1(abar[15]), .A2(bbar[14]), .ZN(ybar[254]);
  AND2_X1 U86 ( .A1(a[15]), .A2(b[13]), .ZN(y[253]) );
  OR2_X1 U86bar ( .A1(abar[15]), .A2(bbar[13]), .ZN(ybar[253]);
  AND2_X1 U87 ( .A1(a[15]), .A2(b[12]), .ZN(y[252]) );
  OR2_X1 U87bar ( .A1(abar[15]), .A2(bbar[12]), .ZN(ybar[252]);
  AND2_X1 U88 ( .A1(a[15]), .A2(b[11]), .ZN(y[251]) );
  OR2_X1 U88bar ( .A1(abar[15]), .A2(bbar[11]), .ZN(ybar[251]);
  AND2_X1 U89 ( .A1(a[15]), .A2(b[10]), .ZN(y[250]) );
  OR2_X1 U89bar ( .A1(abar[15]), .A2(bbar[10]), .ZN(ybar[250]);
  AND2_X1 U90 ( .A1(a[1]), .A2(b[8]), .ZN(y[24]) );
  OR2_X1 U90bar ( .A1(abar[1]), .A2(bbar[8]), .ZN(ybar[24]);
  AND2_X1 U91 ( .A1(a[15]), .A2(b[9]), .ZN(y[249]) );
  OR2_X1 U91bar ( .A1(abar[15]), .A2(bbar[9]), .ZN(ybar[249]);
  AND2_X1 U92 ( .A1(a[15]), .A2(b[8]), .ZN(y[248]) );
  OR2_X1 U92bar ( .A1(abar[15]), .A2(bbar[8]), .ZN(ybar[248]);
  AND2_X1 U93 ( .A1(a[15]), .A2(b[7]), .ZN(y[247]) );
  OR2_X1 U93bar ( .A1(abar[15]), .A2(bbar[7]), .ZN(ybar[247]);
  AND2_X1 U94 ( .A1(a[15]), .A2(b[6]), .ZN(y[246]) );
  OR2_X1 U94bar ( .A1(abar[15]), .A2(bbar[6]), .ZN(ybar[246]);
  AND2_X1 U95 ( .A1(a[15]), .A2(b[5]), .ZN(y[245]) );
  OR2_X1 U95bar ( .A1(abar[15]), .A2(bbar[5]), .ZN(ybar[245]);
  AND2_X1 U96 ( .A1(a[15]), .A2(b[4]), .ZN(y[244]) );
  OR2_X1 U96bar ( .A1(abar[15]), .A2(bbar[4]), .ZN(ybar[244]);
  AND2_X1 U97 ( .A1(a[15]), .A2(b[3]), .ZN(y[243]) );
  OR2_X1 U97bar ( .A1(abar[15]), .A2(bbar[3]), .ZN(ybar[243]);
  AND2_X1 U98 ( .A1(a[15]), .A2(b[2]), .ZN(y[242]) );
  OR2_X1 U98bar ( .A1(abar[15]), .A2(bbar[2]), .ZN(ybar[242]);
  AND2_X1 U99 ( .A1(a[15]), .A2(b[1]), .ZN(y[241]) );
  OR2_X1 U99bar ( .A1(abar[15]), .A2(bbar[1]), .ZN(ybar[241]);
  AND2_X1 U100 ( .A1(a[15]), .A2(b[0]), .ZN(y[240]) );
  OR2_X1 U100bar ( .A1(abar[15]), .A2(bbar[0]), .ZN(ybar[240]);
  AND2_X1 U101 ( .A1(a[1]), .A2(b[7]), .ZN(y[23]) );
  OR2_X1 U101bar ( .A1(abar[1]), .A2(bbar[7]), .ZN(ybar[23]);
  AND2_X1 U102 ( .A1(a[14]), .A2(b[15]), .ZN(y[239]) );
  OR2_X1 U102bar ( .A1(abar[14]), .A2(bbar[15]), .ZN(ybar[239]);
  AND2_X1 U103 ( .A1(a[14]), .A2(b[14]), .ZN(y[238]) );
  OR2_X1 U103bar ( .A1(abar[14]), .A2(bbar[14]), .ZN(ybar[238]);
  AND2_X1 U104 ( .A1(a[14]), .A2(b[13]), .ZN(y[237]) );
  OR2_X1 U104bar ( .A1(abar[14]), .A2(bbar[13]), .ZN(ybar[237]);
  AND2_X1 U105 ( .A1(a[14]), .A2(b[12]), .ZN(y[236]) );
  OR2_X1 U105bar ( .A1(abar[14]), .A2(bbar[12]), .ZN(ybar[236]);
  AND2_X1 U106 ( .A1(a[14]), .A2(b[11]), .ZN(y[235]) );
  OR2_X1 U106bar ( .A1(abar[14]), .A2(bbar[11]), .ZN(ybar[235]);
  AND2_X1 U107 ( .A1(a[14]), .A2(b[10]), .ZN(y[234]) );
  OR2_X1 U107bar ( .A1(abar[14]), .A2(bbar[10]), .ZN(ybar[234]);
  AND2_X1 U108 ( .A1(a[14]), .A2(b[9]), .ZN(y[233]) );
  OR2_X1 U108bar ( .A1(abar[14]), .A2(bbar[9]), .ZN(ybar[233]);
  AND2_X1 U109 ( .A1(a[14]), .A2(b[8]), .ZN(y[232]) );
  OR2_X1 U109bar ( .A1(abar[14]), .A2(bbar[8]), .ZN(ybar[232]);
  AND2_X1 U110 ( .A1(a[14]), .A2(b[7]), .ZN(y[231]) );
  OR2_X1 U110bar ( .A1(abar[14]), .A2(bbar[7]), .ZN(ybar[231]);
  AND2_X1 U111 ( .A1(a[14]), .A2(b[6]), .ZN(y[230]) );
  OR2_X1 U111bar ( .A1(abar[14]), .A2(bbar[6]), .ZN(ybar[230]);
  AND2_X1 U112 ( .A1(a[1]), .A2(b[6]), .ZN(y[22]) );
  OR2_X1 U112bar ( .A1(abar[1]), .A2(bbar[6]), .ZN(ybar[22]);
  AND2_X1 U113 ( .A1(a[14]), .A2(b[5]), .ZN(y[229]) );
  OR2_X1 U113bar ( .A1(abar[14]), .A2(bbar[5]), .ZN(ybar[229]);
  AND2_X1 U114 ( .A1(a[14]), .A2(b[4]), .ZN(y[228]) );
  OR2_X1 U114bar ( .A1(abar[14]), .A2(bbar[4]), .ZN(ybar[228]);
  AND2_X1 U115 ( .A1(a[14]), .A2(b[3]), .ZN(y[227]) );
  OR2_X1 U115bar ( .A1(abar[14]), .A2(bbar[3]), .ZN(ybar[227]);
  AND2_X1 U116 ( .A1(a[14]), .A2(b[2]), .ZN(y[226]) );
  OR2_X1 U116bar ( .A1(abar[14]), .A2(bbar[2]), .ZN(ybar[226]);
  AND2_X1 U117 ( .A1(a[14]), .A2(b[1]), .ZN(y[225]) );
  OR2_X1 U117bar ( .A1(abar[14]), .A2(bbar[1]), .ZN(ybar[225]);
  AND2_X1 U118 ( .A1(a[14]), .A2(b[0]), .ZN(y[224]) );
  OR2_X1 U118bar ( .A1(abar[14]), .A2(bbar[0]), .ZN(ybar[224]);
  AND2_X1 U119 ( .A1(a[13]), .A2(b[15]), .ZN(y[223]) );
  OR2_X1 U119bar ( .A1(abar[13]), .A2(bbar[15]), .ZN(ybar[223]);
  AND2_X1 U120 ( .A1(a[13]), .A2(b[14]), .ZN(y[222]) );
  OR2_X1 U120bar ( .A1(abar[13]), .A2(bbar[14]), .ZN(ybar[222]);
  AND2_X1 U121 ( .A1(a[13]), .A2(b[13]), .ZN(y[221]) );
  OR2_X1 U121bar ( .A1(abar[13]), .A2(bbar[13]), .ZN(ybar[221]);
  AND2_X1 U122 ( .A1(a[13]), .A2(b[12]), .ZN(y[220]) );
  OR2_X1 U122bar ( .A1(abar[13]), .A2(bbar[12]), .ZN(ybar[220]);
  AND2_X1 U123 ( .A1(a[1]), .A2(b[5]), .ZN(y[21]) );
  OR2_X1 U123bar ( .A1(abar[1]), .A2(bbar[5]), .ZN(ybar[21]);
  AND2_X1 U124 ( .A1(a[13]), .A2(b[11]), .ZN(y[219]) );
  OR2_X1 U124bar ( .A1(abar[13]), .A2(bbar[11]), .ZN(ybar[219]);
  AND2_X1 U125 ( .A1(a[13]), .A2(b[10]), .ZN(y[218]) );
  OR2_X1 U125bar ( .A1(abar[13]), .A2(bbar[10]), .ZN(ybar[218]);
  AND2_X1 U126 ( .A1(a[13]), .A2(b[9]), .ZN(y[217]) );
  OR2_X1 U126bar ( .A1(abar[13]), .A2(bbar[9]), .ZN(ybar[217]);
  AND2_X1 U127 ( .A1(a[13]), .A2(b[8]), .ZN(y[216]) );
  OR2_X1 U127bar ( .A1(abar[13]), .A2(bbar[8]), .ZN(ybar[216]);
  AND2_X1 U128 ( .A1(a[13]), .A2(b[7]), .ZN(y[215]) );
  OR2_X1 U128bar ( .A1(abar[13]), .A2(bbar[7]), .ZN(ybar[215]);
  AND2_X1 U129 ( .A1(a[13]), .A2(b[6]), .ZN(y[214]) );
  OR2_X1 U129bar ( .A1(abar[13]), .A2(bbar[6]), .ZN(ybar[214]);
  AND2_X1 U130 ( .A1(a[13]), .A2(b[5]), .ZN(y[213]) );
  OR2_X1 U130bar ( .A1(abar[13]), .A2(bbar[5]), .ZN(ybar[213]);
  AND2_X1 U131 ( .A1(a[13]), .A2(b[4]), .ZN(y[212]) );
  OR2_X1 U131bar ( .A1(abar[13]), .A2(bbar[4]), .ZN(ybar[212]);
  AND2_X1 U132 ( .A1(a[13]), .A2(b[3]), .ZN(y[211]) );
  OR2_X1 U132bar ( .A1(abar[13]), .A2(bbar[3]), .ZN(ybar[211]);
  AND2_X1 U133 ( .A1(a[13]), .A2(b[2]), .ZN(y[210]) );
  OR2_X1 U133bar ( .A1(abar[13]), .A2(bbar[2]), .ZN(ybar[210]);
  AND2_X1 U134 ( .A1(a[1]), .A2(b[4]), .ZN(y[20]) );
  OR2_X1 U134bar ( .A1(abar[1]), .A2(bbar[4]), .ZN(ybar[20]);
  AND2_X1 U135 ( .A1(a[13]), .A2(b[1]), .ZN(y[209]) );
  OR2_X1 U135bar ( .A1(abar[13]), .A2(bbar[1]), .ZN(ybar[209]);
  AND2_X1 U136 ( .A1(a[13]), .A2(b[0]), .ZN(y[208]) );
  OR2_X1 U136bar ( .A1(abar[13]), .A2(bbar[0]), .ZN(ybar[208]);
  AND2_X1 U137 ( .A1(a[12]), .A2(b[15]), .ZN(y[207]) );
  OR2_X1 U137bar ( .A1(abar[12]), .A2(bbar[15]), .ZN(ybar[207]);
  AND2_X1 U138 ( .A1(a[12]), .A2(b[14]), .ZN(y[206]) );
  OR2_X1 U138bar ( .A1(abar[12]), .A2(bbar[14]), .ZN(ybar[206]);
  AND2_X1 U139 ( .A1(a[12]), .A2(b[13]), .ZN(y[205]) );
  OR2_X1 U139bar ( .A1(abar[12]), .A2(bbar[13]), .ZN(ybar[205]);
  AND2_X1 U140 ( .A1(a[12]), .A2(b[12]), .ZN(y[204]) );
  OR2_X1 U140bar ( .A1(abar[12]), .A2(bbar[12]), .ZN(ybar[204]);
  AND2_X1 U141 ( .A1(a[12]), .A2(b[11]), .ZN(y[203]) );
  OR2_X1 U141bar ( .A1(abar[12]), .A2(bbar[11]), .ZN(ybar[203]);
  AND2_X1 U142 ( .A1(a[12]), .A2(b[10]), .ZN(y[202]) );
  OR2_X1 U142bar ( .A1(abar[12]), .A2(bbar[10]), .ZN(ybar[202]);
  AND2_X1 U143 ( .A1(a[12]), .A2(b[9]), .ZN(y[201]) );
  OR2_X1 U143bar ( .A1(abar[12]), .A2(bbar[9]), .ZN(ybar[201]);
  AND2_X1 U144 ( .A1(a[12]), .A2(b[8]), .ZN(y[200]) );
  OR2_X1 U144bar ( .A1(abar[12]), .A2(bbar[8]), .ZN(ybar[200]);
  AND2_X1 U145 ( .A1(b[1]), .A2(a[0]), .ZN(y[1]) );
  OR2_X1 U145bar ( .A1(bbar[1]), .A2(abar[0]), .ZN(ybar[1]);
  AND2_X1 U146 ( .A1(a[1]), .A2(b[3]), .ZN(y[19]) );
  OR2_X1 U146bar ( .A1(abar[1]), .A2(bbar[3]), .ZN(ybar[19]);
  AND2_X1 U147 ( .A1(a[12]), .A2(b[7]), .ZN(y[199]) );
  OR2_X1 U147bar ( .A1(abar[12]), .A2(bbar[7]), .ZN(ybar[199]);
  AND2_X1 U148 ( .A1(a[12]), .A2(b[6]), .ZN(y[198]) );
  OR2_X1 U148bar ( .A1(abar[12]), .A2(bbar[6]), .ZN(ybar[198]);
  AND2_X1 U149 ( .A1(a[12]), .A2(b[5]), .ZN(y[197]) );
  OR2_X1 U149bar ( .A1(abar[12]), .A2(bbar[5]), .ZN(ybar[197]);
  AND2_X1 U150 ( .A1(a[12]), .A2(b[4]), .ZN(y[196]) );
  OR2_X1 U150bar ( .A1(abar[12]), .A2(bbar[4]), .ZN(ybar[196]);
  AND2_X1 U151 ( .A1(a[12]), .A2(b[3]), .ZN(y[195]) );
  OR2_X1 U151bar ( .A1(abar[12]), .A2(bbar[3]), .ZN(ybar[195]);
  AND2_X1 U152 ( .A1(a[12]), .A2(b[2]), .ZN(y[194]) );
  OR2_X1 U152bar ( .A1(abar[12]), .A2(bbar[2]), .ZN(ybar[194]);
  AND2_X1 U153 ( .A1(a[12]), .A2(b[1]), .ZN(y[193]) );
  OR2_X1 U153bar ( .A1(abar[12]), .A2(bbar[1]), .ZN(ybar[193]);
  AND2_X1 U154 ( .A1(a[12]), .A2(b[0]), .ZN(y[192]) );
  OR2_X1 U154bar ( .A1(abar[12]), .A2(bbar[0]), .ZN(ybar[192]);
  AND2_X1 U155 ( .A1(a[11]), .A2(b[15]), .ZN(y[191]) );
  OR2_X1 U155bar ( .A1(abar[11]), .A2(bbar[15]), .ZN(ybar[191]);
  AND2_X1 U156 ( .A1(a[11]), .A2(b[14]), .ZN(y[190]) );
  OR2_X1 U156bar ( .A1(abar[11]), .A2(bbar[14]), .ZN(ybar[190]);
  AND2_X1 U157 ( .A1(a[1]), .A2(b[2]), .ZN(y[18]) );
  OR2_X1 U157bar ( .A1(abar[1]), .A2(bbar[2]), .ZN(ybar[18]);
  AND2_X1 U158 ( .A1(a[11]), .A2(b[13]), .ZN(y[189]) );
  OR2_X1 U158bar ( .A1(abar[11]), .A2(bbar[13]), .ZN(ybar[189]);
  AND2_X1 U159 ( .A1(a[11]), .A2(b[12]), .ZN(y[188]) );
  OR2_X1 U159bar ( .A1(abar[11]), .A2(bbar[12]), .ZN(ybar[188]);
  AND2_X1 U160 ( .A1(a[11]), .A2(b[11]), .ZN(y[187]) );
  OR2_X1 U160bar ( .A1(abar[11]), .A2(bbar[11]), .ZN(ybar[187]);
  AND2_X1 U161 ( .A1(a[11]), .A2(b[10]), .ZN(y[186]) );
  OR2_X1 U161bar ( .A1(abar[11]), .A2(bbar[10]), .ZN(ybar[186]);
  AND2_X1 U162 ( .A1(a[11]), .A2(b[9]), .ZN(y[185]) );
  OR2_X1 U162bar ( .A1(abar[11]), .A2(bbar[9]), .ZN(ybar[185]);
  AND2_X1 U163 ( .A1(a[11]), .A2(b[8]), .ZN(y[184]) );
  OR2_X1 U163bar ( .A1(abar[11]), .A2(bbar[8]), .ZN(ybar[184]);
  AND2_X1 U164 ( .A1(a[11]), .A2(b[7]), .ZN(y[183]) );
  OR2_X1 U164bar ( .A1(abar[11]), .A2(bbar[7]), .ZN(ybar[183]);
  AND2_X1 U165 ( .A1(a[11]), .A2(b[6]), .ZN(y[182]) );
  OR2_X1 U165bar ( .A1(abar[11]), .A2(bbar[6]), .ZN(ybar[182]);
  AND2_X1 U166 ( .A1(a[11]), .A2(b[5]), .ZN(y[181]) );
  OR2_X1 U166bar ( .A1(abar[11]), .A2(bbar[5]), .ZN(ybar[181]);
  AND2_X1 U167 ( .A1(a[11]), .A2(b[4]), .ZN(y[180]) );
  OR2_X1 U167bar ( .A1(abar[11]), .A2(bbar[4]), .ZN(ybar[180]);
  AND2_X1 U168 ( .A1(a[1]), .A2(b[1]), .ZN(y[17]) );
  OR2_X1 U168bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[17]);
  AND2_X1 U169 ( .A1(a[11]), .A2(b[3]), .ZN(y[179]) );
  OR2_X1 U169bar ( .A1(abar[11]), .A2(bbar[3]), .ZN(ybar[179]);
  AND2_X1 U170 ( .A1(a[11]), .A2(b[2]), .ZN(y[178]) );
  OR2_X1 U170bar ( .A1(abar[11]), .A2(bbar[2]), .ZN(ybar[178]);
  AND2_X1 U171 ( .A1(a[11]), .A2(b[1]), .ZN(y[177]) );
  OR2_X1 U171bar ( .A1(abar[11]), .A2(bbar[1]), .ZN(ybar[177]);
  AND2_X1 U172 ( .A1(a[11]), .A2(b[0]), .ZN(y[176]) );
  OR2_X1 U172bar ( .A1(abar[11]), .A2(bbar[0]), .ZN(ybar[176]);
  AND2_X1 U173 ( .A1(a[10]), .A2(b[15]), .ZN(y[175]) );
  OR2_X1 U173bar ( .A1(abar[10]), .A2(bbar[15]), .ZN(ybar[175]);
  AND2_X1 U174 ( .A1(a[10]), .A2(b[14]), .ZN(y[174]) );
  OR2_X1 U174bar ( .A1(abar[10]), .A2(bbar[14]), .ZN(ybar[174]);
  AND2_X1 U175 ( .A1(a[10]), .A2(b[13]), .ZN(y[173]) );
  OR2_X1 U175bar ( .A1(abar[10]), .A2(bbar[13]), .ZN(ybar[173]);
  AND2_X1 U176 ( .A1(a[10]), .A2(b[12]), .ZN(y[172]) );
  OR2_X1 U176bar ( .A1(abar[10]), .A2(bbar[12]), .ZN(ybar[172]);
  AND2_X1 U177 ( .A1(a[10]), .A2(b[11]), .ZN(y[171]) );
  OR2_X1 U177bar ( .A1(abar[10]), .A2(bbar[11]), .ZN(ybar[171]);
  AND2_X1 U178 ( .A1(a[10]), .A2(b[10]), .ZN(y[170]) );
  OR2_X1 U178bar ( .A1(abar[10]), .A2(bbar[10]), .ZN(ybar[170]);
  AND2_X1 U179 ( .A1(a[1]), .A2(b[0]), .ZN(y[16]) );
  OR2_X1 U179bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[16]);
  AND2_X1 U180 ( .A1(a[10]), .A2(b[9]), .ZN(y[169]) );
  OR2_X1 U180bar ( .A1(abar[10]), .A2(bbar[9]), .ZN(ybar[169]);
  AND2_X1 U181 ( .A1(a[10]), .A2(b[8]), .ZN(y[168]) );
  OR2_X1 U181bar ( .A1(abar[10]), .A2(bbar[8]), .ZN(ybar[168]);
  AND2_X1 U182 ( .A1(a[10]), .A2(b[7]), .ZN(y[167]) );
  OR2_X1 U182bar ( .A1(abar[10]), .A2(bbar[7]), .ZN(ybar[167]);
  AND2_X1 U183 ( .A1(a[10]), .A2(b[6]), .ZN(y[166]) );
  OR2_X1 U183bar ( .A1(abar[10]), .A2(bbar[6]), .ZN(ybar[166]);
  AND2_X1 U184 ( .A1(a[10]), .A2(b[5]), .ZN(y[165]) );
  OR2_X1 U184bar ( .A1(abar[10]), .A2(bbar[5]), .ZN(ybar[165]);
  AND2_X1 U185 ( .A1(a[10]), .A2(b[4]), .ZN(y[164]) );
  OR2_X1 U185bar ( .A1(abar[10]), .A2(bbar[4]), .ZN(ybar[164]);
  AND2_X1 U186 ( .A1(a[10]), .A2(b[3]), .ZN(y[163]) );
  OR2_X1 U186bar ( .A1(abar[10]), .A2(bbar[3]), .ZN(ybar[163]);
  AND2_X1 U187 ( .A1(a[10]), .A2(b[2]), .ZN(y[162]) );
  OR2_X1 U187bar ( .A1(abar[10]), .A2(bbar[2]), .ZN(ybar[162]);
  AND2_X1 U188 ( .A1(a[10]), .A2(b[1]), .ZN(y[161]) );
  OR2_X1 U188bar ( .A1(abar[10]), .A2(bbar[1]), .ZN(ybar[161]);
  AND2_X1 U189 ( .A1(a[10]), .A2(b[0]), .ZN(y[160]) );
  OR2_X1 U189bar ( .A1(abar[10]), .A2(bbar[0]), .ZN(ybar[160]);
  AND2_X1 U190 ( .A1(b[15]), .A2(a[0]), .ZN(y[15]) );
  OR2_X1 U190bar ( .A1(bbar[15]), .A2(abar[0]), .ZN(ybar[15]);
  AND2_X1 U191 ( .A1(a[9]), .A2(b[15]), .ZN(y[159]) );
  OR2_X1 U191bar ( .A1(abar[9]), .A2(bbar[15]), .ZN(ybar[159]);
  AND2_X1 U192 ( .A1(a[9]), .A2(b[14]), .ZN(y[158]) );
  OR2_X1 U192bar ( .A1(abar[9]), .A2(bbar[14]), .ZN(ybar[158]);
  AND2_X1 U193 ( .A1(a[9]), .A2(b[13]), .ZN(y[157]) );
  OR2_X1 U193bar ( .A1(abar[9]), .A2(bbar[13]), .ZN(ybar[157]);
  AND2_X1 U194 ( .A1(a[9]), .A2(b[12]), .ZN(y[156]) );
  OR2_X1 U194bar ( .A1(abar[9]), .A2(bbar[12]), .ZN(ybar[156]);
  AND2_X1 U195 ( .A1(a[9]), .A2(b[11]), .ZN(y[155]) );
  OR2_X1 U195bar ( .A1(abar[9]), .A2(bbar[11]), .ZN(ybar[155]);
  AND2_X1 U196 ( .A1(a[9]), .A2(b[10]), .ZN(y[154]) );
  OR2_X1 U196bar ( .A1(abar[9]), .A2(bbar[10]), .ZN(ybar[154]);
  AND2_X1 U197 ( .A1(a[9]), .A2(b[9]), .ZN(y[153]) );
  OR2_X1 U197bar ( .A1(abar[9]), .A2(bbar[9]), .ZN(ybar[153]);
  AND2_X1 U198 ( .A1(a[9]), .A2(b[8]), .ZN(y[152]) );
  OR2_X1 U198bar ( .A1(abar[9]), .A2(bbar[8]), .ZN(ybar[152]);
  AND2_X1 U199 ( .A1(a[9]), .A2(b[7]), .ZN(y[151]) );
  OR2_X1 U199bar ( .A1(abar[9]), .A2(bbar[7]), .ZN(ybar[151]);
  AND2_X1 U200 ( .A1(a[9]), .A2(b[6]), .ZN(y[150]) );
  OR2_X1 U200bar ( .A1(abar[9]), .A2(bbar[6]), .ZN(ybar[150]);
  AND2_X1 U201 ( .A1(b[14]), .A2(a[0]), .ZN(y[14]) );
  OR2_X1 U201bar ( .A1(bbar[14]), .A2(abar[0]), .ZN(ybar[14]);
  AND2_X1 U202 ( .A1(a[9]), .A2(b[5]), .ZN(y[149]) );
  OR2_X1 U202bar ( .A1(abar[9]), .A2(bbar[5]), .ZN(ybar[149]);
  AND2_X1 U203 ( .A1(a[9]), .A2(b[4]), .ZN(y[148]) );
  OR2_X1 U203bar ( .A1(abar[9]), .A2(bbar[4]), .ZN(ybar[148]);
  AND2_X1 U204 ( .A1(a[9]), .A2(b[3]), .ZN(y[147]) );
  OR2_X1 U204bar ( .A1(abar[9]), .A2(bbar[3]), .ZN(ybar[147]);
  AND2_X1 U205 ( .A1(a[9]), .A2(b[2]), .ZN(y[146]) );
  OR2_X1 U205bar ( .A1(abar[9]), .A2(bbar[2]), .ZN(ybar[146]);
  AND2_X1 U206 ( .A1(a[9]), .A2(b[1]), .ZN(y[145]) );
  OR2_X1 U206bar ( .A1(abar[9]), .A2(bbar[1]), .ZN(ybar[145]);
  AND2_X1 U207 ( .A1(a[9]), .A2(b[0]), .ZN(y[144]) );
  OR2_X1 U207bar ( .A1(abar[9]), .A2(bbar[0]), .ZN(ybar[144]);
  AND2_X1 U208 ( .A1(a[8]), .A2(b[15]), .ZN(y[143]) );
  OR2_X1 U208bar ( .A1(abar[8]), .A2(bbar[15]), .ZN(ybar[143]);
  AND2_X1 U209 ( .A1(a[8]), .A2(b[14]), .ZN(y[142]) );
  OR2_X1 U209bar ( .A1(abar[8]), .A2(bbar[14]), .ZN(ybar[142]);
  AND2_X1 U210 ( .A1(a[8]), .A2(b[13]), .ZN(y[141]) );
  OR2_X1 U210bar ( .A1(abar[8]), .A2(bbar[13]), .ZN(ybar[141]);
  AND2_X1 U211 ( .A1(a[8]), .A2(b[12]), .ZN(y[140]) );
  OR2_X1 U211bar ( .A1(abar[8]), .A2(bbar[12]), .ZN(ybar[140]);
  AND2_X1 U212 ( .A1(b[13]), .A2(a[0]), .ZN(y[13]) );
  OR2_X1 U212bar ( .A1(bbar[13]), .A2(abar[0]), .ZN(ybar[13]);
  AND2_X1 U213 ( .A1(a[8]), .A2(b[11]), .ZN(y[139]) );
  OR2_X1 U213bar ( .A1(abar[8]), .A2(bbar[11]), .ZN(ybar[139]);
  AND2_X1 U214 ( .A1(a[8]), .A2(b[10]), .ZN(y[138]) );
  OR2_X1 U214bar ( .A1(abar[8]), .A2(bbar[10]), .ZN(ybar[138]);
  AND2_X1 U215 ( .A1(a[8]), .A2(b[9]), .ZN(y[137]) );
  OR2_X1 U215bar ( .A1(abar[8]), .A2(bbar[9]), .ZN(ybar[137]);
  AND2_X1 U216 ( .A1(a[8]), .A2(b[8]), .ZN(y[136]) );
  OR2_X1 U216bar ( .A1(abar[8]), .A2(bbar[8]), .ZN(ybar[136]);
  AND2_X1 U217 ( .A1(a[8]), .A2(b[7]), .ZN(y[135]) );
  OR2_X1 U217bar ( .A1(abar[8]), .A2(bbar[7]), .ZN(ybar[135]);
  AND2_X1 U218 ( .A1(a[8]), .A2(b[6]), .ZN(y[134]) );
  OR2_X1 U218bar ( .A1(abar[8]), .A2(bbar[6]), .ZN(ybar[134]);
  AND2_X1 U219 ( .A1(a[8]), .A2(b[5]), .ZN(y[133]) );
  OR2_X1 U219bar ( .A1(abar[8]), .A2(bbar[5]), .ZN(ybar[133]);
  AND2_X1 U220 ( .A1(a[8]), .A2(b[4]), .ZN(y[132]) );
  OR2_X1 U220bar ( .A1(abar[8]), .A2(bbar[4]), .ZN(ybar[132]);
  AND2_X1 U221 ( .A1(a[8]), .A2(b[3]), .ZN(y[131]) );
  OR2_X1 U221bar ( .A1(abar[8]), .A2(bbar[3]), .ZN(ybar[131]);
  AND2_X1 U222 ( .A1(a[8]), .A2(b[2]), .ZN(y[130]) );
  OR2_X1 U222bar ( .A1(abar[8]), .A2(bbar[2]), .ZN(ybar[130]);
  AND2_X1 U223 ( .A1(b[12]), .A2(a[0]), .ZN(y[12]) );
  OR2_X1 U223bar ( .A1(bbar[12]), .A2(abar[0]), .ZN(ybar[12]);
  AND2_X1 U224 ( .A1(a[8]), .A2(b[1]), .ZN(y[129]) );
  OR2_X1 U224bar ( .A1(abar[8]), .A2(bbar[1]), .ZN(ybar[129]);
  AND2_X1 U225 ( .A1(a[8]), .A2(b[0]), .ZN(y[128]) );
  OR2_X1 U225bar ( .A1(abar[8]), .A2(bbar[0]), .ZN(ybar[128]);
  AND2_X1 U226 ( .A1(a[7]), .A2(b[15]), .ZN(y[127]) );
  OR2_X1 U226bar ( .A1(abar[7]), .A2(bbar[15]), .ZN(ybar[127]);
  AND2_X1 U227 ( .A1(a[7]), .A2(b[14]), .ZN(y[126]) );
  OR2_X1 U227bar ( .A1(abar[7]), .A2(bbar[14]), .ZN(ybar[126]);
  AND2_X1 U228 ( .A1(a[7]), .A2(b[13]), .ZN(y[125]) );
  OR2_X1 U228bar ( .A1(abar[7]), .A2(bbar[13]), .ZN(ybar[125]);
  AND2_X1 U229 ( .A1(a[7]), .A2(b[12]), .ZN(y[124]) );
  OR2_X1 U229bar ( .A1(abar[7]), .A2(bbar[12]), .ZN(ybar[124]);
  AND2_X1 U230 ( .A1(a[7]), .A2(b[11]), .ZN(y[123]) );
  OR2_X1 U230bar ( .A1(abar[7]), .A2(bbar[11]), .ZN(ybar[123]);
  AND2_X1 U231 ( .A1(a[7]), .A2(b[10]), .ZN(y[122]) );
  OR2_X1 U231bar ( .A1(abar[7]), .A2(bbar[10]), .ZN(ybar[122]);
  AND2_X1 U232 ( .A1(a[7]), .A2(b[9]), .ZN(y[121]) );
  OR2_X1 U232bar ( .A1(abar[7]), .A2(bbar[9]), .ZN(ybar[121]);
  AND2_X1 U233 ( .A1(a[7]), .A2(b[8]), .ZN(y[120]) );
  OR2_X1 U233bar ( .A1(abar[7]), .A2(bbar[8]), .ZN(ybar[120]);
  AND2_X1 U234 ( .A1(b[11]), .A2(a[0]), .ZN(y[11]) );
  OR2_X1 U234bar ( .A1(bbar[11]), .A2(abar[0]), .ZN(ybar[11]);
  AND2_X1 U235 ( .A1(a[7]), .A2(b[7]), .ZN(y[119]) );
  OR2_X1 U235bar ( .A1(abar[7]), .A2(bbar[7]), .ZN(ybar[119]);
  AND2_X1 U236 ( .A1(a[7]), .A2(b[6]), .ZN(y[118]) );
  OR2_X1 U236bar ( .A1(abar[7]), .A2(bbar[6]), .ZN(ybar[118]);
  AND2_X1 U237 ( .A1(a[7]), .A2(b[5]), .ZN(y[117]) );
  OR2_X1 U237bar ( .A1(abar[7]), .A2(bbar[5]), .ZN(ybar[117]);
  AND2_X1 U238 ( .A1(a[7]), .A2(b[4]), .ZN(y[116]) );
  OR2_X1 U238bar ( .A1(abar[7]), .A2(bbar[4]), .ZN(ybar[116]);
  AND2_X1 U239 ( .A1(a[7]), .A2(b[3]), .ZN(y[115]) );
  OR2_X1 U239bar ( .A1(abar[7]), .A2(bbar[3]), .ZN(ybar[115]);
  AND2_X1 U240 ( .A1(a[7]), .A2(b[2]), .ZN(y[114]) );
  OR2_X1 U240bar ( .A1(abar[7]), .A2(bbar[2]), .ZN(ybar[114]);
  AND2_X1 U241 ( .A1(a[7]), .A2(b[1]), .ZN(y[113]) );
  OR2_X1 U241bar ( .A1(abar[7]), .A2(bbar[1]), .ZN(ybar[113]);
  AND2_X1 U242 ( .A1(a[7]), .A2(b[0]), .ZN(y[112]) );
  OR2_X1 U242bar ( .A1(abar[7]), .A2(bbar[0]), .ZN(ybar[112]);
  AND2_X1 U243 ( .A1(b[15]), .A2(a[6]), .ZN(y[111]) );
  OR2_X1 U243bar ( .A1(bbar[15]), .A2(abar[6]), .ZN(ybar[111]);
  AND2_X1 U244 ( .A1(b[14]), .A2(a[6]), .ZN(y[110]) );
  OR2_X1 U244bar ( .A1(bbar[14]), .A2(abar[6]), .ZN(ybar[110]);
  AND2_X1 U245 ( .A1(b[10]), .A2(a[0]), .ZN(y[10]) );
  OR2_X1 U245bar ( .A1(bbar[10]), .A2(abar[0]), .ZN(ybar[10]);
  AND2_X1 U246 ( .A1(b[13]), .A2(a[6]), .ZN(y[109]) );
  OR2_X1 U246bar ( .A1(bbar[13]), .A2(abar[6]), .ZN(ybar[109]);
  AND2_X1 U247 ( .A1(b[12]), .A2(a[6]), .ZN(y[108]) );
  OR2_X1 U247bar ( .A1(bbar[12]), .A2(abar[6]), .ZN(ybar[108]);
  AND2_X1 U248 ( .A1(b[11]), .A2(a[6]), .ZN(y[107]) );
  OR2_X1 U248bar ( .A1(bbar[11]), .A2(abar[6]), .ZN(ybar[107]);
  AND2_X1 U249 ( .A1(b[10]), .A2(a[6]), .ZN(y[106]) );
  OR2_X1 U249bar ( .A1(bbar[10]), .A2(abar[6]), .ZN(ybar[106]);
  AND2_X1 U250 ( .A1(a[6]), .A2(b[9]), .ZN(y[105]) );
  OR2_X1 U250bar ( .A1(abar[6]), .A2(bbar[9]), .ZN(ybar[105]);
  AND2_X1 U251 ( .A1(b[8]), .A2(a[6]), .ZN(y[104]) );
  OR2_X1 U251bar ( .A1(bbar[8]), .A2(abar[6]), .ZN(ybar[104]);
  AND2_X1 U252 ( .A1(b[7]), .A2(a[6]), .ZN(y[103]) );
  OR2_X1 U252bar ( .A1(bbar[7]), .A2(abar[6]), .ZN(ybar[103]);
  AND2_X1 U253 ( .A1(b[6]), .A2(a[6]), .ZN(y[102]) );
  OR2_X1 U253bar ( .A1(bbar[6]), .A2(abar[6]), .ZN(ybar[102]);
  AND2_X1 U254 ( .A1(b[5]), .A2(a[6]), .ZN(y[101]) );
  OR2_X1 U254bar ( .A1(bbar[5]), .A2(abar[6]), .ZN(ybar[101]);
  AND2_X1 U255 ( .A1(b[4]), .A2(a[6]), .ZN(y[100]) );
  OR2_X1 U255bar ( .A1(bbar[4]), .A2(abar[6]), .ZN(ybar[100]);
  AND2_X1 U256 ( .A1(b[0]), .A2(a[0]), .ZN(y[0]) );
  OR2_X1 U256bar ( .A1(bbar[0]), .A2(abar[0]), .ZN(ybar[0]);
endmodule




module decode_2 ( in, out );
  input [7:0] in;
  //input_done

  output [255:0] out;
  //output_done

  wire   [15:0] level1;
  wire   [31:0] level2;
  //wire_done

  CD2_8 cd_l1_1 ( .a(in[1]), .b(in[0]), .y(level1[3:0]) );
  CD2_7 cd_l1_2 ( .a(in[3]), .b(in[2]), .y(level1[7:4]) );
  CD2_6 cd_l1_3 ( .a(in[5]), .b(in[4]), .y(level1[11:8]) );
  CD2_5 cd_l1_4 ( .a(in[7]), .b(in[6]), .y(level1[15:12]) );
  CD4_4 cd_l2_1 ( .a(level1[7:4]), .b(level1[3:0]), .y(level2[15:0]) );
  CD4_3 cd_l2_2 ( .a(level1[15:12]), .b(level1[11:8]), .y(level2[31:16]) );
  CD16_2 cd_l3 ( .a(level2[31:16]), .b(level2[15:0]), .y(out) );
endmodule


module encode_2 ( in, out );
  input [255:0] in;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
  assign inbar[8] = ~in[8];
  assign inbar[9] = ~in[9];
  assign inbar[10] = ~in[10];
  assign inbar[11] = ~in[11];
  assign inbar[12] = ~in[12];
  assign inbar[13] = ~in[13];
  assign inbar[14] = ~in[14];
  assign inbar[15] = ~in[15];
  assign inbar[16] = ~in[16];
  assign inbar[17] = ~in[17];
  assign inbar[18] = ~in[18];
  assign inbar[19] = ~in[19];
  assign inbar[20] = ~in[20];
  assign inbar[21] = ~in[21];
  assign inbar[22] = ~in[22];
  assign inbar[23] = ~in[23];
  assign inbar[24] = ~in[24];
  assign inbar[25] = ~in[25];
  assign inbar[26] = ~in[26];
  assign inbar[27] = ~in[27];
  assign inbar[28] = ~in[28];
  assign inbar[29] = ~in[29];
  assign inbar[30] = ~in[30];
  assign inbar[31] = ~in[31];
  assign inbar[32] = ~in[32];
  assign inbar[33] = ~in[33];
  assign inbar[34] = ~in[34];
  assign inbar[35] = ~in[35];
  assign inbar[36] = ~in[36];
  assign inbar[37] = ~in[37];
  assign inbar[38] = ~in[38];
  assign inbar[39] = ~in[39];
  assign inbar[40] = ~in[40];
  assign inbar[41] = ~in[41];
  assign inbar[42] = ~in[42];
  assign inbar[43] = ~in[43];
  assign inbar[44] = ~in[44];
  assign inbar[45] = ~in[45];
  assign inbar[46] = ~in[46];
  assign inbar[47] = ~in[47];
  assign inbar[48] = ~in[48];
  assign inbar[49] = ~in[49];
  assign inbar[50] = ~in[50];
  assign inbar[51] = ~in[51];
  assign inbar[52] = ~in[52];
  assign inbar[53] = ~in[53];
  assign inbar[54] = ~in[54];
  assign inbar[55] = ~in[55];
  assign inbar[56] = ~in[56];
  assign inbar[57] = ~in[57];
  assign inbar[58] = ~in[58];
  assign inbar[59] = ~in[59];
  assign inbar[60] = ~in[60];
  assign inbar[61] = ~in[61];
  assign inbar[62] = ~in[62];
  assign inbar[63] = ~in[63];
  assign inbar[64] = ~in[64];
  assign inbar[65] = ~in[65];
  assign inbar[66] = ~in[66];
  assign inbar[67] = ~in[67];
  assign inbar[68] = ~in[68];
  assign inbar[69] = ~in[69];
  assign inbar[70] = ~in[70];
  assign inbar[71] = ~in[71];
  assign inbar[72] = ~in[72];
  assign inbar[73] = ~in[73];
  assign inbar[74] = ~in[74];
  assign inbar[75] = ~in[75];
  assign inbar[76] = ~in[76];
  assign inbar[77] = ~in[77];
  assign inbar[78] = ~in[78];
  assign inbar[79] = ~in[79];
  assign inbar[80] = ~in[80];
  assign inbar[81] = ~in[81];
  assign inbar[82] = ~in[82];
  assign inbar[83] = ~in[83];
  assign inbar[84] = ~in[84];
  assign inbar[85] = ~in[85];
  assign inbar[86] = ~in[86];
  assign inbar[87] = ~in[87];
  assign inbar[88] = ~in[88];
  assign inbar[89] = ~in[89];
  assign inbar[90] = ~in[90];
  assign inbar[91] = ~in[91];
  assign inbar[92] = ~in[92];
  assign inbar[93] = ~in[93];
  assign inbar[94] = ~in[94];
  assign inbar[95] = ~in[95];
  assign inbar[96] = ~in[96];
  assign inbar[97] = ~in[97];
  assign inbar[98] = ~in[98];
  assign inbar[99] = ~in[99];
  assign inbar[100] = ~in[100];
  assign inbar[101] = ~in[101];
  assign inbar[102] = ~in[102];
  assign inbar[103] = ~in[103];
  assign inbar[104] = ~in[104];
  assign inbar[105] = ~in[105];
  assign inbar[106] = ~in[106];
  assign inbar[107] = ~in[107];
  assign inbar[108] = ~in[108];
  assign inbar[109] = ~in[109];
  assign inbar[110] = ~in[110];
  assign inbar[111] = ~in[111];
  assign inbar[112] = ~in[112];
  assign inbar[113] = ~in[113];
  assign inbar[114] = ~in[114];
  assign inbar[115] = ~in[115];
  assign inbar[116] = ~in[116];
  assign inbar[117] = ~in[117];
  assign inbar[118] = ~in[118];
  assign inbar[119] = ~in[119];
  assign inbar[120] = ~in[120];
  assign inbar[121] = ~in[121];
  assign inbar[122] = ~in[122];
  assign inbar[123] = ~in[123];
  assign inbar[124] = ~in[124];
  assign inbar[125] = ~in[125];
  assign inbar[126] = ~in[126];
  assign inbar[127] = ~in[127];
  assign inbar[128] = ~in[128];
  assign inbar[129] = ~in[129];
  assign inbar[130] = ~in[130];
  assign inbar[131] = ~in[131];
  assign inbar[132] = ~in[132];
  assign inbar[133] = ~in[133];
  assign inbar[134] = ~in[134];
  assign inbar[135] = ~in[135];
  assign inbar[136] = ~in[136];
  assign inbar[137] = ~in[137];
  assign inbar[138] = ~in[138];
  assign inbar[139] = ~in[139];
  assign inbar[140] = ~in[140];
  assign inbar[141] = ~in[141];
  assign inbar[142] = ~in[142];
  assign inbar[143] = ~in[143];
  assign inbar[144] = ~in[144];
  assign inbar[145] = ~in[145];
  assign inbar[146] = ~in[146];
  assign inbar[147] = ~in[147];
  assign inbar[148] = ~in[148];
  assign inbar[149] = ~in[149];
  assign inbar[150] = ~in[150];
  assign inbar[151] = ~in[151];
  assign inbar[152] = ~in[152];
  assign inbar[153] = ~in[153];
  assign inbar[154] = ~in[154];
  assign inbar[155] = ~in[155];
  assign inbar[156] = ~in[156];
  assign inbar[157] = ~in[157];
  assign inbar[158] = ~in[158];
  assign inbar[159] = ~in[159];
  assign inbar[160] = ~in[160];
  assign inbar[161] = ~in[161];
  assign inbar[162] = ~in[162];
  assign inbar[163] = ~in[163];
  assign inbar[164] = ~in[164];
  assign inbar[165] = ~in[165];
  assign inbar[166] = ~in[166];
  assign inbar[167] = ~in[167];
  assign inbar[168] = ~in[168];
  assign inbar[169] = ~in[169];
  assign inbar[170] = ~in[170];
  assign inbar[171] = ~in[171];
  assign inbar[172] = ~in[172];
  assign inbar[173] = ~in[173];
  assign inbar[174] = ~in[174];
  assign inbar[175] = ~in[175];
  assign inbar[176] = ~in[176];
  assign inbar[177] = ~in[177];
  assign inbar[178] = ~in[178];
  assign inbar[179] = ~in[179];
  assign inbar[180] = ~in[180];
  assign inbar[181] = ~in[181];
  assign inbar[182] = ~in[182];
  assign inbar[183] = ~in[183];
  assign inbar[184] = ~in[184];
  assign inbar[185] = ~in[185];
  assign inbar[186] = ~in[186];
  assign inbar[187] = ~in[187];
  assign inbar[188] = ~in[188];
  assign inbar[189] = ~in[189];
  assign inbar[190] = ~in[190];
  assign inbar[191] = ~in[191];
  assign inbar[192] = ~in[192];
  assign inbar[193] = ~in[193];
  assign inbar[194] = ~in[194];
  assign inbar[195] = ~in[195];
  assign inbar[196] = ~in[196];
  assign inbar[197] = ~in[197];
  assign inbar[198] = ~in[198];
  assign inbar[199] = ~in[199];
  assign inbar[200] = ~in[200];
  assign inbar[201] = ~in[201];
  assign inbar[202] = ~in[202];
  assign inbar[203] = ~in[203];
  assign inbar[204] = ~in[204];
  assign inbar[205] = ~in[205];
  assign inbar[206] = ~in[206];
  assign inbar[207] = ~in[207];
  assign inbar[208] = ~in[208];
  assign inbar[209] = ~in[209];
  assign inbar[210] = ~in[210];
  assign inbar[211] = ~in[211];
  assign inbar[212] = ~in[212];
  assign inbar[213] = ~in[213];
  assign inbar[214] = ~in[214];
  assign inbar[215] = ~in[215];
  assign inbar[216] = ~in[216];
  assign inbar[217] = ~in[217];
  assign inbar[218] = ~in[218];
  assign inbar[219] = ~in[219];
  assign inbar[220] = ~in[220];
  assign inbar[221] = ~in[221];
  assign inbar[222] = ~in[222];
  assign inbar[223] = ~in[223];
  assign inbar[224] = ~in[224];
  assign inbar[225] = ~in[225];
  assign inbar[226] = ~in[226];
  assign inbar[227] = ~in[227];
  assign inbar[228] = ~in[228];
  assign inbar[229] = ~in[229];
  assign inbar[230] = ~in[230];
  assign inbar[231] = ~in[231];
  assign inbar[232] = ~in[232];
  assign inbar[233] = ~in[233];
  assign inbar[234] = ~in[234];
  assign inbar[235] = ~in[235];
  assign inbar[236] = ~in[236];
  assign inbar[237] = ~in[237];
  assign inbar[238] = ~in[238];
  assign inbar[239] = ~in[239];
  assign inbar[240] = ~in[240];
  assign inbar[241] = ~in[241];
  assign inbar[242] = ~in[242];
  assign inbar[243] = ~in[243];
  assign inbar[244] = ~in[244];
  assign inbar[245] = ~in[245];
  assign inbar[246] = ~in[246];
  assign inbar[247] = ~in[247];
  assign inbar[248] = ~in[248];
  assign inbar[249] = ~in[249];
  assign inbar[250] = ~in[250];
  assign inbar[251] = ~in[251];
  assign inbar[252] = ~in[252];
  assign inbar[253] = ~in[253];
  assign inbar[254] = ~in[254];
  assign inbar[255] = ~in[255];
  //input_done

  output [7:0] out;
  reg [7:0] outbar;
  //output_done

  wire   in_81, in_80, in_79, in_78, in_77, in_76, in_75, in_74, in_73, in_72,
         in_71, in_70, in_69, in_68, in_67, in_66, in_65, in_64, in_63, in_62,
         in_61, in_60, in_59, in_58, in_57, in_56, in_55, in_54, in_53, in_52,
         in_51, in_50, in_49, in_48, in_47, in_46, in_45, in_44, in_43, in_42,
         in_41, in_40, in_39, in_38, in_37, in_36, in_35, in_34, in_33, in_32,
         in_31, in_30, in_29, in_28, in_27, in_26, in_25, in_24, in_23, in_22,
         in_21, in_20, in_19, in_18, in_17, in_16, in_15, in_14, in_13, in_12,
         in_11, in_10, in_9, in_8, in_7, in_6, in_5, in_4, in_3, in_2, in_1,
         in_0, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972;
  wire in_81bar, in_80bar, in_79bar, in_78bar, in_77bar, in_76bar, in_75bar, in_74bar, in_73bar, in_72bar, in_71bar, in_70bar, in_69bar, in_68bar, in_67bar, in_66bar, in_65bar, in_64bar, in_63bar, in_62bar, in_61bar, in_60bar, in_59bar, in_58bar, in_57bar, in_56bar, in_55bar, in_54bar, in_53bar, in_52bar, in_51bar, in_50bar, in_49bar, in_48bar, in_47bar, in_46bar, in_45bar, in_44bar, in_43bar, in_42bar, in_41bar, in_40bar, in_39bar, in_38bar, in_37bar, in_36bar, in_35bar, in_34bar, in_33bar, in_32bar, in_31bar, in_30bar, in_29bar, in_28bar, in_27bar, in_26bar, in_25bar, in_24bar, in_23bar, in_22bar, in_21bar, in_20bar, in_19bar, in_18bar, in_17bar, in_16bar, in_15bar, in_14bar, in_13bar, in_12bar, in_11bar, in_10bar, in_9bar, in_8bar, in_7bar, in_6bar, in_5bar, in_4bar, in_3bar, in_2bar, in_1bar, in_0bar, n487bar, n488bar, n489bar, n490bar, n491bar, n492bar, n493bar, n494bar, n495bar, n496bar, n497bar, n498bar, n499bar, n500bar, n501bar, n502bar, n503bar, n504bar, n505bar, n506bar, n507bar, n508bar, n509bar, n510bar, n511bar, n512bar, n513bar, n514bar, n515bar, n516bar, n517bar, n518bar, n519bar, n520bar, n521bar, n522bar, n523bar, n524bar, n525bar, n526bar, n527bar, n528bar, n529bar, n530bar, n531bar, n532bar, n533bar, n534bar, n535bar, n536bar, n537bar, n538bar, n539bar, n540bar, n541bar, n542bar, n543bar, n544bar, n545bar, n546bar, n547bar, n548bar, n549bar, n550bar, n551bar, n552bar, n553bar, n554bar, n555bar, n556bar, n557bar, n558bar, n559bar, n560bar, n561bar, n562bar, n563bar, n564bar, n565bar, n566bar, n567bar, n568bar, n569bar, n570bar, n571bar, n572bar, n573bar, n574bar, n575bar, n576bar, n577bar, n578bar, n579bar, n580bar, n581bar, n582bar, n583bar, n584bar, n585bar, n586bar, n587bar, n588bar, n589bar, n590bar, n591bar, n592bar, n593bar, n594bar, n595bar, n596bar, n597bar, n598bar, n599bar, n600bar, n601bar, n602bar, n603bar, n604bar, n605bar, n606bar, n607bar, n608bar, n609bar, n610bar, n611bar, n612bar, n613bar, n614bar, n615bar, n616bar, n617bar, n618bar, n619bar, n620bar, n621bar, n622bar, n623bar, n624bar, n625bar, n626bar, n627bar, n628bar, n629bar, n630bar, n631bar, n632bar, n633bar, n634bar, n635bar, n636bar, n637bar, n638bar, n639bar, n640bar, n641bar, n642bar, n643bar, n644bar, n645bar, n646bar, n647bar, n648bar, n649bar, n650bar, n651bar, n652bar, n653bar, n654bar, n655bar, n656bar, n657bar, n658bar, n659bar, n660bar, n661bar, n662bar, n663bar, n664bar, n665bar, n666bar, n667bar, n668bar, n669bar, n670bar, n671bar, n672bar, n673bar, n674bar, n675bar, n676bar, n677bar, n678bar, n679bar, n680bar, n681bar, n682bar, n683bar, n684bar, n685bar, n686bar, n687bar, n688bar, n689bar, n690bar, n691bar, n692bar, n693bar, n694bar, n695bar, n696bar, n697bar, n698bar, n699bar, n700bar, n701bar, n702bar, n703bar, n704bar, n705bar, n706bar, n707bar, n708bar, n709bar, n710bar, n711bar, n712bar, n713bar, n714bar, n715bar, n716bar, n717bar, n718bar, n719bar, n720bar, n721bar, n722bar, n723bar, n724bar, n725bar, n726bar, n727bar, n728bar, n729bar, n730bar, n731bar, n732bar, n733bar, n734bar, n735bar, n736bar, n737bar, n738bar, n739bar, n740bar, n741bar, n742bar, n743bar, n744bar, n745bar, n746bar, n747bar, n748bar, n749bar, n750bar, n751bar, n752bar, n753bar, n754bar, n755bar, n756bar, n757bar, n758bar, n759bar, n760bar, n761bar, n762bar, n763bar, n764bar, n765bar, n766bar, n767bar, n768bar, n769bar, n770bar, n771bar, n772bar, n773bar, n774bar, n775bar, n776bar, n777bar, n778bar, n779bar, n780bar, n781bar, n782bar, n783bar, n784bar, n785bar, n786bar, n787bar, n788bar, n789bar, n790bar, n791bar, n792bar, n793bar, n794bar, n795bar, n796bar, n797bar, n798bar, n799bar, n800bar, n801bar, n802bar, n803bar, n804bar, n805bar, n806bar, n807bar, n808bar, n809bar, n810bar, n811bar, n812bar, n813bar, n814bar, n815bar, n816bar, n817bar, n818bar, n819bar, n820bar, n821bar, n822bar, n823bar, n824bar, n825bar, n826bar, n827bar, n828bar, n829bar, n830bar, n831bar, n832bar, n833bar, n834bar, n835bar, n836bar, n837bar, n838bar, n839bar, n840bar, n841bar, n842bar, n843bar, n844bar, n845bar, n846bar, n847bar, n848bar, n849bar, n850bar, n851bar, n852bar, n853bar, n854bar, n855bar, n856bar, n857bar, n858bar, n859bar, n860bar, n861bar, n862bar, n863bar, n864bar, n865bar, n866bar, n867bar, n868bar, n869bar, n870bar, n871bar, n872bar, n873bar, n874bar, n875bar, n876bar, n877bar, n878bar, n879bar, n880bar, n881bar, n882bar, n883bar, n884bar, n885bar, n886bar, n887bar, n888bar, n889bar, n890bar, n891bar, n892bar, n893bar, n894bar, n895bar, n896bar, n897bar, n898bar, n899bar, n900bar, n901bar, n902bar, n903bar, n904bar, n905bar, n906bar, n907bar, n908bar, n909bar, n910bar, n911bar, n912bar, n913bar, n914bar, n915bar, n916bar, n917bar, n918bar, n919bar, n920bar, n921bar, n922bar, n923bar, n924bar, n925bar, n926bar, n927bar, n928bar, n929bar, n930bar, n931bar, n932bar, n933bar, n934bar, n935bar, n936bar, n937bar, n938bar, n939bar, n940bar, n941bar, n942bar, n943bar, n944bar, n945bar, n946bar, n947bar, n948bar, n949bar, n950bar, n951bar, n952bar, n953bar, n954bar, n955bar, n956bar, n957bar, n958bar, n959bar, n960bar, n961bar, n962bar, n963bar, n964bar, n965bar, n966bar, n967bar, n968bar, n969bar, n970bar, n971bar, n972bar;
  //wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];

  OR2_X1 U1 ( .A1(n972), .A2(n971), .ZN(out[7]) );
  AND2_X1 U1bar ( .A1(n972bar), .A2(n971bar), .ZN(outbar[7]);
  OR2_X1 U2 ( .A1(n970), .A2(n969), .ZN(n971) );
  AND2_X1 U2bar ( .A1(n970bar), .A2(n969bar), .ZN(n971bar);
  OR2_X1 U3 ( .A1(n968), .A2(n967), .ZN(n969) );
  AND2_X1 U3bar ( .A1(n968bar), .A2(n967bar), .ZN(n969bar);
  OR2_X1 U4 ( .A1(n966), .A2(n965), .ZN(n967) );
  AND2_X1 U4bar ( .A1(n966bar), .A2(n965bar), .ZN(n967bar);
  OR2_X1 U5 ( .A1(n964), .A2(n963), .ZN(n968) );
  AND2_X1 U5bar ( .A1(n964bar), .A2(n963bar), .ZN(n968bar);
  OR2_X1 U6 ( .A1(in[116]), .A2(n962), .ZN(n963) );
  AND2_X1 U6bar ( .A1(inbar[116]), .A2(n962bar), .ZN(n963bar);
  OR2_X1 U7 ( .A1(n961), .A2(n960), .ZN(n970) );
  AND2_X1 U7bar ( .A1(n961bar), .A2(n960bar), .ZN(n970bar);
  OR2_X1 U8 ( .A1(in[150]), .A2(in[127]), .ZN(n960) );
  AND2_X1 U8bar ( .A1(inbar[150]), .A2(inbar[127]), .ZN(n960bar);
  OR2_X1 U9 ( .A1(in[160]), .A2(n959), .ZN(n961) );
  AND2_X1 U9bar ( .A1(inbar[160]), .A2(n959bar), .ZN(n961bar);
  OR2_X1 U10 ( .A1(in[252]), .A2(in[168]), .ZN(n959) );
  AND2_X1 U10bar ( .A1(inbar[252]), .A2(inbar[168]), .ZN(n959bar);
  OR2_X1 U11 ( .A1(n958), .A2(n957), .ZN(n972) );
  AND2_X1 U11bar ( .A1(n958bar), .A2(n957bar), .ZN(n972bar);
  OR2_X1 U12 ( .A1(n956), .A2(n955), .ZN(n957) );
  AND2_X1 U12bar ( .A1(n956bar), .A2(n955bar), .ZN(n957bar);
  OR2_X1 U13 ( .A1(in_17), .A2(in[96]), .ZN(n955) );
  AND2_X1 U13bar ( .A1(in_17bar), .A2(inbar[96]), .ZN(n955bar);
  OR2_X1 U14 ( .A1(in_23), .A2(n954), .ZN(n956) );
  AND2_X1 U14bar ( .A1(in_23bar), .A2(n954bar), .ZN(n956bar);
  OR2_X1 U15 ( .A1(in_31), .A2(in_26), .ZN(n954) );
  AND2_X1 U15bar ( .A1(in_31bar), .A2(in_26bar), .ZN(n954bar);
  OR2_X1 U16 ( .A1(n953), .A2(n952), .ZN(n958) );
  AND2_X1 U16bar ( .A1(n953bar), .A2(n952bar), .ZN(n958bar);
  OR2_X1 U17 ( .A1(in_58), .A2(in_4), .ZN(n952) );
  AND2_X1 U17bar ( .A1(in_58bar), .A2(in_4bar), .ZN(n952bar);
  OR2_X1 U18 ( .A1(in_59), .A2(n951), .ZN(n953) );
  AND2_X1 U18bar ( .A1(in_59bar), .A2(n951bar), .ZN(n953bar);
  OR2_X1 U19 ( .A1(in_71), .A2(in_62), .ZN(n951) );
  AND2_X1 U19bar ( .A1(in_71bar), .A2(in_62bar), .ZN(n951bar);
  OR2_X1 U20 ( .A1(n950), .A2(n949), .ZN(out[6]) );
  AND2_X1 U20bar ( .A1(n950bar), .A2(n949bar), .ZN(outbar[6]);
  OR2_X1 U21 ( .A1(n948), .A2(n947), .ZN(n949) );
  AND2_X1 U21bar ( .A1(n948bar), .A2(n947bar), .ZN(n949bar);
  OR2_X1 U22 ( .A1(n946), .A2(n945), .ZN(n947) );
  AND2_X1 U22bar ( .A1(n946bar), .A2(n945bar), .ZN(n947bar);
  OR2_X1 U23 ( .A1(n944), .A2(n943), .ZN(n945) );
  AND2_X1 U23bar ( .A1(n944bar), .A2(n943bar), .ZN(n945bar);
  OR2_X1 U24 ( .A1(n942), .A2(n941), .ZN(n946) );
  AND2_X1 U24bar ( .A1(n942bar), .A2(n941bar), .ZN(n946bar);
  OR2_X1 U25 ( .A1(in[101]), .A2(n940), .ZN(n941) );
  AND2_X1 U25bar ( .A1(inbar[101]), .A2(n940bar), .ZN(n941bar);
  OR2_X1 U26 ( .A1(n939), .A2(n938), .ZN(n948) );
  AND2_X1 U26bar ( .A1(n939bar), .A2(n938bar), .ZN(n948bar);
  OR2_X1 U27 ( .A1(in[114]), .A2(in[104]), .ZN(n938) );
  AND2_X1 U27bar ( .A1(inbar[114]), .A2(inbar[104]), .ZN(n938bar);
  OR2_X1 U28 ( .A1(in[128]), .A2(n937), .ZN(n939) );
  AND2_X1 U28bar ( .A1(inbar[128]), .A2(n937bar), .ZN(n939bar);
  OR2_X1 U29 ( .A1(in[136]), .A2(in[134]), .ZN(n937) );
  AND2_X1 U29bar ( .A1(inbar[136]), .A2(inbar[134]), .ZN(n937bar);
  OR2_X1 U30 ( .A1(n936), .A2(n935), .ZN(n950) );
  AND2_X1 U30bar ( .A1(n936bar), .A2(n935bar), .ZN(n950bar);
  OR2_X1 U31 ( .A1(n934), .A2(n933), .ZN(n935) );
  AND2_X1 U31bar ( .A1(n934bar), .A2(n933bar), .ZN(n935bar);
  OR2_X1 U32 ( .A1(in[177]), .A2(in[164]), .ZN(n933) );
  AND2_X1 U32bar ( .A1(inbar[177]), .A2(inbar[164]), .ZN(n933bar);
  OR2_X1 U33 ( .A1(in[212]), .A2(n932), .ZN(n934) );
  AND2_X1 U33bar ( .A1(inbar[212]), .A2(n932bar), .ZN(n934bar);
  OR2_X1 U34 ( .A1(in[248]), .A2(in[221]), .ZN(n932) );
  AND2_X1 U34bar ( .A1(inbar[248]), .A2(inbar[221]), .ZN(n932bar);
  OR2_X1 U35 ( .A1(n931), .A2(n930), .ZN(n936) );
  AND2_X1 U35bar ( .A1(n931bar), .A2(n930bar), .ZN(n936bar);
  OR2_X1 U36 ( .A1(in_18), .A2(in[93]), .ZN(n930) );
  AND2_X1 U36bar ( .A1(in_18bar), .A2(inbar[93]), .ZN(n930bar);
  OR2_X1 U37 ( .A1(in_31), .A2(n929), .ZN(n931) );
  AND2_X1 U37bar ( .A1(in_31bar), .A2(n929bar), .ZN(n931bar);
  OR2_X1 U38 ( .A1(in_7), .A2(in_39), .ZN(n929) );
  AND2_X1 U38bar ( .A1(in_7bar), .A2(in_39bar), .ZN(n929bar);
  OR2_X1 U39 ( .A1(n928), .A2(n927), .ZN(out[5]) );
  AND2_X1 U39bar ( .A1(n928bar), .A2(n927bar), .ZN(outbar[5]);
  OR2_X1 U40 ( .A1(n926), .A2(n925), .ZN(n927) );
  AND2_X1 U40bar ( .A1(n926bar), .A2(n925bar), .ZN(n927bar);
  OR2_X1 U41 ( .A1(n924), .A2(n923), .ZN(n925) );
  AND2_X1 U41bar ( .A1(n924bar), .A2(n923bar), .ZN(n925bar);
  OR2_X1 U42 ( .A1(n922), .A2(n921), .ZN(n923) );
  AND2_X1 U42bar ( .A1(n922bar), .A2(n921bar), .ZN(n923bar);
  OR2_X1 U43 ( .A1(n940), .A2(n920), .ZN(n924) );
  AND2_X1 U43bar ( .A1(n940bar), .A2(n920bar), .ZN(n924bar);
  OR2_X1 U44 ( .A1(in[111]), .A2(n919), .ZN(n920) );
  AND2_X1 U44bar ( .A1(inbar[111]), .A2(n919bar), .ZN(n920bar);
  OR2_X1 U45 ( .A1(n918), .A2(n917), .ZN(n940) );
  AND2_X1 U45bar ( .A1(n918bar), .A2(n917bar), .ZN(n940bar);
  OR2_X1 U46 ( .A1(n916), .A2(n915), .ZN(n917) );
  AND2_X1 U46bar ( .A1(n916bar), .A2(n915bar), .ZN(n917bar);
  OR2_X1 U47 ( .A1(n914), .A2(n913), .ZN(n915) );
  AND2_X1 U47bar ( .A1(n914bar), .A2(n913bar), .ZN(n915bar);
  OR2_X1 U48 ( .A1(in[140]), .A2(in[131]), .ZN(n913) );
  AND2_X1 U48bar ( .A1(inbar[140]), .A2(inbar[131]), .ZN(n913bar);
  OR2_X1 U49 ( .A1(in[160]), .A2(in[144]), .ZN(n914) );
  AND2_X1 U49bar ( .A1(inbar[160]), .A2(inbar[144]), .ZN(n914bar);
  OR2_X1 U50 ( .A1(n912), .A2(n911), .ZN(n916) );
  AND2_X1 U50bar ( .A1(n912bar), .A2(n911bar), .ZN(n916bar);
  OR2_X1 U51 ( .A1(in[179]), .A2(in[174]), .ZN(n911) );
  AND2_X1 U51bar ( .A1(inbar[179]), .A2(inbar[174]), .ZN(n911bar);
  OR2_X1 U52 ( .A1(in[188]), .A2(in[184]), .ZN(n912) );
  AND2_X1 U52bar ( .A1(inbar[188]), .A2(inbar[184]), .ZN(n912bar);
  OR2_X1 U53 ( .A1(n910), .A2(n909), .ZN(n918) );
  AND2_X1 U53bar ( .A1(n910bar), .A2(n909bar), .ZN(n918bar);
  OR2_X1 U54 ( .A1(n908), .A2(n907), .ZN(n909) );
  AND2_X1 U54bar ( .A1(n908bar), .A2(n907bar), .ZN(n909bar);
  OR2_X1 U55 ( .A1(in[216]), .A2(in[200]), .ZN(n907) );
  AND2_X1 U55bar ( .A1(inbar[216]), .A2(inbar[200]), .ZN(n907bar);
  OR2_X1 U56 ( .A1(in[228]), .A2(in[224]), .ZN(n908) );
  AND2_X1 U56bar ( .A1(inbar[228]), .A2(inbar[224]), .ZN(n908bar);
  OR2_X1 U57 ( .A1(n906), .A2(n905), .ZN(n910) );
  AND2_X1 U57bar ( .A1(n906bar), .A2(n905bar), .ZN(n910bar);
  OR2_X1 U58 ( .A1(in[247]), .A2(in[235]), .ZN(n905) );
  AND2_X1 U58bar ( .A1(inbar[247]), .A2(inbar[235]), .ZN(n905bar);
  OR2_X1 U59 ( .A1(in_42), .A2(in[83]), .ZN(n906) );
  AND2_X1 U59bar ( .A1(in_42bar), .A2(inbar[83]), .ZN(n906bar);
  OR2_X1 U60 ( .A1(n904), .A2(n903), .ZN(n926) );
  AND2_X1 U60bar ( .A1(n904bar), .A2(n903bar), .ZN(n926bar);
  OR2_X1 U61 ( .A1(in[166]), .A2(in[123]), .ZN(n903) );
  AND2_X1 U61bar ( .A1(inbar[166]), .A2(inbar[123]), .ZN(n903bar);
  OR2_X1 U62 ( .A1(in[170]), .A2(n902), .ZN(n904) );
  AND2_X1 U62bar ( .A1(inbar[170]), .A2(n902bar), .ZN(n904bar);
  OR2_X1 U63 ( .A1(in[194]), .A2(in[183]), .ZN(n902) );
  AND2_X1 U63bar ( .A1(inbar[194]), .A2(inbar[183]), .ZN(n902bar);
  OR2_X1 U64 ( .A1(n901), .A2(n900), .ZN(n928) );
  AND2_X1 U64bar ( .A1(n901bar), .A2(n900bar), .ZN(n928bar);
  OR2_X1 U65 ( .A1(n899), .A2(n898), .ZN(n900) );
  AND2_X1 U65bar ( .A1(n899bar), .A2(n898bar), .ZN(n900bar);
  OR2_X1 U66 ( .A1(in[241]), .A2(in[238]), .ZN(n898) );
  AND2_X1 U66bar ( .A1(inbar[241]), .A2(inbar[238]), .ZN(n898bar);
  OR2_X1 U67 ( .A1(in[250]), .A2(n897), .ZN(n899) );
  AND2_X1 U67bar ( .A1(inbar[250]), .A2(n897bar), .ZN(n899bar);
  OR2_X1 U68 ( .A1(in_24), .A2(in[84]), .ZN(n897) );
  AND2_X1 U68bar ( .A1(in_24bar), .A2(inbar[84]), .ZN(n897bar);
  OR2_X1 U69 ( .A1(n896), .A2(n895), .ZN(n901) );
  AND2_X1 U69bar ( .A1(n896bar), .A2(n895bar), .ZN(n901bar);
  OR2_X1 U70 ( .A1(in_41), .A2(in_29), .ZN(n895) );
  AND2_X1 U70bar ( .A1(in_41bar), .A2(in_29bar), .ZN(n895bar);
  OR2_X1 U71 ( .A1(in_66), .A2(n894), .ZN(n896) );
  AND2_X1 U71bar ( .A1(in_66bar), .A2(n894bar), .ZN(n896bar);
  OR2_X1 U72 ( .A1(in_76), .A2(in_71), .ZN(n894) );
  AND2_X1 U72bar ( .A1(in_76bar), .A2(in_71bar), .ZN(n894bar);
  OR2_X1 U73 ( .A1(n893), .A2(n892), .ZN(out[4]) );
  AND2_X1 U73bar ( .A1(n893bar), .A2(n892bar), .ZN(outbar[4]);
  OR2_X1 U74 ( .A1(n891), .A2(n890), .ZN(n892) );
  AND2_X1 U74bar ( .A1(n891bar), .A2(n890bar), .ZN(n892bar);
  OR2_X1 U75 ( .A1(n889), .A2(n888), .ZN(n890) );
  AND2_X1 U75bar ( .A1(n889bar), .A2(n888bar), .ZN(n890bar);
  OR2_X1 U76 ( .A1(n922), .A2(n887), .ZN(n888) );
  AND2_X1 U76bar ( .A1(n922bar), .A2(n887bar), .ZN(n888bar);
  OR2_X1 U77 ( .A1(n886), .A2(n885), .ZN(n922) );
  AND2_X1 U77bar ( .A1(n886bar), .A2(n885bar), .ZN(n922bar);
  OR2_X1 U78 ( .A1(n884), .A2(n883), .ZN(n885) );
  AND2_X1 U78bar ( .A1(n884bar), .A2(n883bar), .ZN(n885bar);
  OR2_X1 U79 ( .A1(n882), .A2(n881), .ZN(n883) );
  AND2_X1 U79bar ( .A1(n882bar), .A2(n881bar), .ZN(n883bar);
  OR2_X1 U80 ( .A1(in[118]), .A2(in[109]), .ZN(n881) );
  AND2_X1 U80bar ( .A1(inbar[118]), .A2(inbar[109]), .ZN(n881bar);
  OR2_X1 U81 ( .A1(in[139]), .A2(in[120]), .ZN(n882) );
  AND2_X1 U81bar ( .A1(inbar[139]), .A2(inbar[120]), .ZN(n882bar);
  OR2_X1 U82 ( .A1(n880), .A2(n879), .ZN(n884) );
  AND2_X1 U82bar ( .A1(n880bar), .A2(n879bar), .ZN(n884bar);
  OR2_X1 U83 ( .A1(in[198]), .A2(in[154]), .ZN(n879) );
  AND2_X1 U83bar ( .A1(inbar[198]), .A2(inbar[154]), .ZN(n879bar);
  OR2_X1 U84 ( .A1(in[210]), .A2(in[205]), .ZN(n880) );
  AND2_X1 U84bar ( .A1(inbar[210]), .A2(inbar[205]), .ZN(n880bar);
  OR2_X1 U85 ( .A1(n878), .A2(n877), .ZN(n886) );
  AND2_X1 U85bar ( .A1(n878bar), .A2(n877bar), .ZN(n886bar);
  OR2_X1 U86 ( .A1(n876), .A2(n875), .ZN(n877) );
  AND2_X1 U86bar ( .A1(n876bar), .A2(n875bar), .ZN(n877bar);
  OR2_X1 U87 ( .A1(in[219]), .A2(in[217]), .ZN(n875) );
  AND2_X1 U87bar ( .A1(inbar[219]), .A2(inbar[217]), .ZN(n875bar);
  OR2_X1 U88 ( .A1(in[86]), .A2(in[252]), .ZN(n876) );
  AND2_X1 U88bar ( .A1(inbar[86]), .A2(inbar[252]), .ZN(n876bar);
  OR2_X1 U89 ( .A1(n874), .A2(n873), .ZN(n878) );
  AND2_X1 U89bar ( .A1(n874bar), .A2(n873bar), .ZN(n878bar);
  OR2_X1 U90 ( .A1(in_40), .A2(in[91]), .ZN(n873) );
  AND2_X1 U90bar ( .A1(in_40bar), .A2(inbar[91]), .ZN(n873bar);
  OR2_X1 U91 ( .A1(in_8), .A2(in_46), .ZN(n874) );
  AND2_X1 U91bar ( .A1(in_8bar), .A2(in_46bar), .ZN(n874bar);
  OR2_X1 U92 ( .A1(n872), .A2(n871), .ZN(n889) );
  AND2_X1 U92bar ( .A1(n872bar), .A2(n871bar), .ZN(n889bar);
  OR2_X1 U93 ( .A1(in[117]), .A2(n943), .ZN(n871) );
  AND2_X1 U93bar ( .A1(inbar[117]), .A2(n943bar), .ZN(n871bar);
  OR2_X1 U94 ( .A1(n870), .A2(n869), .ZN(n943) );
  AND2_X1 U94bar ( .A1(n870bar), .A2(n869bar), .ZN(n943bar);
  OR2_X1 U95 ( .A1(n868), .A2(n867), .ZN(n869) );
  AND2_X1 U95bar ( .A1(n868bar), .A2(n867bar), .ZN(n869bar);
  OR2_X1 U96 ( .A1(n866), .A2(n865), .ZN(n867) );
  AND2_X1 U96bar ( .A1(n866bar), .A2(n865bar), .ZN(n867bar);
  OR2_X1 U97 ( .A1(n864), .A2(n863), .ZN(n865) );
  AND2_X1 U97bar ( .A1(n864bar), .A2(n863bar), .ZN(n865bar);
  OR2_X1 U98 ( .A1(in[108]), .A2(n919), .ZN(n866) );
  AND2_X1 U98bar ( .A1(inbar[108]), .A2(n919bar), .ZN(n866bar);
  OR2_X1 U99 ( .A1(n862), .A2(n861), .ZN(n919) );
  AND2_X1 U99bar ( .A1(n862bar), .A2(n861bar), .ZN(n919bar);
  OR2_X1 U100 ( .A1(n860), .A2(n859), .ZN(n861) );
  AND2_X1 U100bar ( .A1(n860bar), .A2(n859bar), .ZN(n861bar);
  OR2_X1 U101 ( .A1(n858), .A2(n857), .ZN(n859) );
  AND2_X1 U101bar ( .A1(n858bar), .A2(n857bar), .ZN(n859bar);
  OR2_X1 U102 ( .A1(in[119]), .A2(in[105]), .ZN(n857) );
  AND2_X1 U102bar ( .A1(inbar[119]), .A2(inbar[105]), .ZN(n857bar);
  OR2_X1 U103 ( .A1(in[186]), .A2(in[175]), .ZN(n858) );
  AND2_X1 U103bar ( .A1(inbar[186]), .A2(inbar[175]), .ZN(n858bar);
  OR2_X1 U104 ( .A1(n856), .A2(n855), .ZN(n860) );
  AND2_X1 U104bar ( .A1(n856bar), .A2(n855bar), .ZN(n860bar);
  OR2_X1 U105 ( .A1(in[202]), .A2(in[193]), .ZN(n855) );
  AND2_X1 U105bar ( .A1(inbar[202]), .A2(inbar[193]), .ZN(n855bar);
  OR2_X1 U106 ( .A1(in[225]), .A2(in[208]), .ZN(n856) );
  AND2_X1 U106bar ( .A1(inbar[225]), .A2(inbar[208]), .ZN(n856bar);
  OR2_X1 U107 ( .A1(n854), .A2(n853), .ZN(n862) );
  AND2_X1 U107bar ( .A1(n854bar), .A2(n853bar), .ZN(n862bar);
  OR2_X1 U108 ( .A1(n852), .A2(n851), .ZN(n853) );
  AND2_X1 U108bar ( .A1(n852bar), .A2(n851bar), .ZN(n853bar);
  OR2_X1 U109 ( .A1(in_1), .A2(in[85]), .ZN(n851) );
  AND2_X1 U109bar ( .A1(in_1bar), .A2(inbar[85]), .ZN(n851bar);
  OR2_X1 U110 ( .A1(in_23), .A2(in_19), .ZN(n852) );
  AND2_X1 U110bar ( .A1(in_23bar), .A2(in_19bar), .ZN(n852bar);
  OR2_X1 U111 ( .A1(n850), .A2(n849), .ZN(n854) );
  AND2_X1 U111bar ( .A1(n850bar), .A2(n849bar), .ZN(n854bar);
  OR2_X1 U112 ( .A1(in_43), .A2(in_33), .ZN(n849) );
  AND2_X1 U112bar ( .A1(in_43bar), .A2(in_33bar), .ZN(n849bar);
  OR2_X1 U113 ( .A1(in_63), .A2(in_44), .ZN(n850) );
  AND2_X1 U113bar ( .A1(in_63bar), .A2(in_44bar), .ZN(n850bar);
  OR2_X1 U114 ( .A1(n848), .A2(n847), .ZN(n868) );
  AND2_X1 U114bar ( .A1(n848bar), .A2(n847bar), .ZN(n868bar);
  OR2_X1 U115 ( .A1(in[141]), .A2(in[112]), .ZN(n847) );
  AND2_X1 U115bar ( .A1(inbar[141]), .A2(inbar[112]), .ZN(n847bar);
  OR2_X1 U116 ( .A1(in[147]), .A2(n846), .ZN(n848) );
  AND2_X1 U116bar ( .A1(inbar[147]), .A2(n846bar), .ZN(n848bar);
  OR2_X1 U117 ( .A1(in[181]), .A2(in[167]), .ZN(n846) );
  AND2_X1 U117bar ( .A1(inbar[181]), .A2(inbar[167]), .ZN(n846bar);
  OR2_X1 U118 ( .A1(n845), .A2(n844), .ZN(n870) );
  AND2_X1 U118bar ( .A1(n845bar), .A2(n844bar), .ZN(n870bar);
  OR2_X1 U119 ( .A1(n843), .A2(n842), .ZN(n844) );
  AND2_X1 U119bar ( .A1(n843bar), .A2(n842bar), .ZN(n844bar);
  OR2_X1 U120 ( .A1(in[229]), .A2(in[201]), .ZN(n842) );
  AND2_X1 U120bar ( .A1(inbar[229]), .A2(inbar[201]), .ZN(n842bar);
  OR2_X1 U121 ( .A1(in[237]), .A2(n841), .ZN(n843) );
  AND2_X1 U121bar ( .A1(inbar[237]), .A2(n841bar), .ZN(n843bar);
  OR2_X1 U122 ( .A1(in[94]), .A2(in[253]), .ZN(n841) );
  AND2_X1 U122bar ( .A1(inbar[94]), .A2(inbar[253]), .ZN(n841bar);
  OR2_X1 U123 ( .A1(n840), .A2(n839), .ZN(n845) );
  AND2_X1 U123bar ( .A1(n840bar), .A2(n839bar), .ZN(n845bar);
  OR2_X1 U124 ( .A1(in_21), .A2(in[96]), .ZN(n839) );
  AND2_X1 U124bar ( .A1(in_21bar), .A2(inbar[96]), .ZN(n839bar);
  OR2_X1 U125 ( .A1(in_25), .A2(n838), .ZN(n840) );
  AND2_X1 U125bar ( .A1(in_25bar), .A2(n838bar), .ZN(n840bar);
  OR2_X1 U126 ( .A1(in_81), .A2(in_45), .ZN(n838) );
  AND2_X1 U126bar ( .A1(in_81bar), .A2(in_45bar), .ZN(n838bar);
  OR2_X1 U127 ( .A1(n837), .A2(n836), .ZN(n891) );
  AND2_X1 U127bar ( .A1(n837bar), .A2(n836bar), .ZN(n891bar);
  OR2_X1 U128 ( .A1(in[142]), .A2(in[124]), .ZN(n836) );
  AND2_X1 U128bar ( .A1(inbar[142]), .A2(inbar[124]), .ZN(n836bar);
  OR2_X1 U129 ( .A1(in[150]), .A2(n835), .ZN(n837) );
  AND2_X1 U129bar ( .A1(inbar[150]), .A2(n835bar), .ZN(n837bar);
  OR2_X1 U130 ( .A1(in[172]), .A2(in[155]), .ZN(n835) );
  AND2_X1 U130bar ( .A1(inbar[172]), .A2(inbar[155]), .ZN(n835bar);
  OR2_X1 U131 ( .A1(n834), .A2(n833), .ZN(n893) );
  AND2_X1 U131bar ( .A1(n834bar), .A2(n833bar), .ZN(n893bar);
  OR2_X1 U132 ( .A1(n832), .A2(n831), .ZN(n833) );
  AND2_X1 U132bar ( .A1(n832bar), .A2(n831bar), .ZN(n833bar);
  OR2_X1 U133 ( .A1(in[196]), .A2(in[173]), .ZN(n831) );
  AND2_X1 U133bar ( .A1(inbar[196]), .A2(inbar[173]), .ZN(n831bar);
  OR2_X1 U134 ( .A1(in[222]), .A2(n830), .ZN(n832) );
  AND2_X1 U134bar ( .A1(inbar[222]), .A2(n830bar), .ZN(n832bar);
  OR2_X1 U135 ( .A1(in[227]), .A2(in[226]), .ZN(n830) );
  AND2_X1 U135bar ( .A1(inbar[227]), .A2(inbar[226]), .ZN(n830bar);
  OR2_X1 U136 ( .A1(n829), .A2(n828), .ZN(n834) );
  AND2_X1 U136bar ( .A1(n829bar), .A2(n828bar), .ZN(n834bar);
  OR2_X1 U137 ( .A1(in[249]), .A2(in[231]), .ZN(n828) );
  AND2_X1 U137bar ( .A1(inbar[249]), .A2(inbar[231]), .ZN(n828bar);
  OR2_X1 U138 ( .A1(in_28), .A2(n827), .ZN(n829) );
  AND2_X1 U138bar ( .A1(in_28bar), .A2(n827bar), .ZN(n829bar);
  OR2_X1 U139 ( .A1(in_52), .A2(in_47), .ZN(n827) );
  AND2_X1 U139bar ( .A1(in_52bar), .A2(in_47bar), .ZN(n827bar);
  OR2_X1 U140 ( .A1(n826), .A2(n825), .ZN(out[3]) );
  AND2_X1 U140bar ( .A1(n826bar), .A2(n825bar), .ZN(outbar[3]);
  OR2_X1 U141 ( .A1(n824), .A2(n823), .ZN(n825) );
  AND2_X1 U141bar ( .A1(n824bar), .A2(n823bar), .ZN(n825bar);
  OR2_X1 U142 ( .A1(n822), .A2(n821), .ZN(n823) );
  AND2_X1 U142bar ( .A1(n822bar), .A2(n821bar), .ZN(n823bar);
  OR2_X1 U143 ( .A1(n820), .A2(n819), .ZN(n821) );
  AND2_X1 U143bar ( .A1(n820bar), .A2(n819bar), .ZN(n821bar);
  OR2_X1 U144 ( .A1(n964), .A2(n818), .ZN(n822) );
  AND2_X1 U144bar ( .A1(n964bar), .A2(n818bar), .ZN(n822bar);
  OR2_X1 U145 ( .A1(in[118]), .A2(n817), .ZN(n818) );
  AND2_X1 U145bar ( .A1(inbar[118]), .A2(n817bar), .ZN(n818bar);
  OR2_X1 U146 ( .A1(n816), .A2(n815), .ZN(n964) );
  AND2_X1 U146bar ( .A1(n816bar), .A2(n815bar), .ZN(n964bar);
  OR2_X1 U147 ( .A1(n814), .A2(n813), .ZN(n815) );
  AND2_X1 U147bar ( .A1(n814bar), .A2(n813bar), .ZN(n815bar);
  OR2_X1 U148 ( .A1(n812), .A2(n811), .ZN(n813) );
  AND2_X1 U148bar ( .A1(n812bar), .A2(n811bar), .ZN(n813bar);
  OR2_X1 U149 ( .A1(in[122]), .A2(in[111]), .ZN(n811) );
  AND2_X1 U149bar ( .A1(inbar[122]), .A2(inbar[111]), .ZN(n811bar);
  OR2_X1 U150 ( .A1(in[154]), .A2(in[151]), .ZN(n812) );
  AND2_X1 U150bar ( .A1(inbar[154]), .A2(inbar[151]), .ZN(n812bar);
  OR2_X1 U151 ( .A1(n810), .A2(n809), .ZN(n814) );
  AND2_X1 U151bar ( .A1(n810bar), .A2(n809bar), .ZN(n814bar);
  OR2_X1 U152 ( .A1(in[187]), .A2(in[177]), .ZN(n809) );
  AND2_X1 U152bar ( .A1(inbar[187]), .A2(inbar[177]), .ZN(n809bar);
  OR2_X1 U153 ( .A1(in[200]), .A2(in[192]), .ZN(n810) );
  AND2_X1 U153bar ( .A1(inbar[200]), .A2(inbar[192]), .ZN(n810bar);
  OR2_X1 U154 ( .A1(n808), .A2(n807), .ZN(n816) );
  AND2_X1 U154bar ( .A1(n808bar), .A2(n807bar), .ZN(n816bar);
  OR2_X1 U155 ( .A1(n806), .A2(n805), .ZN(n807) );
  AND2_X1 U155bar ( .A1(n806bar), .A2(n805bar), .ZN(n807bar);
  OR2_X1 U156 ( .A1(in[225]), .A2(in[207]), .ZN(n805) );
  AND2_X1 U156bar ( .A1(inbar[225]), .A2(inbar[207]), .ZN(n805bar);
  OR2_X1 U157 ( .A1(in[98]), .A2(in[226]), .ZN(n806) );
  AND2_X1 U157bar ( .A1(inbar[98]), .A2(inbar[226]), .ZN(n806bar);
  OR2_X1 U158 ( .A1(n804), .A2(n803), .ZN(n808) );
  AND2_X1 U158bar ( .A1(n804bar), .A2(n803bar), .ZN(n808bar);
  OR2_X1 U159 ( .A1(in_20), .A2(in_16), .ZN(n803) );
  AND2_X1 U159bar ( .A1(in_20bar), .A2(in_16bar), .ZN(n803bar);
  OR2_X1 U160 ( .A1(in_55), .A2(in_45), .ZN(n804) );
  AND2_X1 U160bar ( .A1(in_55bar), .A2(in_45bar), .ZN(n804bar);
  OR2_X1 U161 ( .A1(n802), .A2(n801), .ZN(n824) );
  AND2_X1 U161bar ( .A1(n802bar), .A2(n801bar), .ZN(n824bar);
  OR2_X1 U162 ( .A1(in[162]), .A2(in[149]), .ZN(n801) );
  AND2_X1 U162bar ( .A1(inbar[162]), .A2(inbar[149]), .ZN(n801bar);
  OR2_X1 U163 ( .A1(in[163]), .A2(n800), .ZN(n802) );
  AND2_X1 U163bar ( .A1(inbar[163]), .A2(n800bar), .ZN(n802bar);
  OR2_X1 U164 ( .A1(in[191]), .A2(in[189]), .ZN(n800) );
  AND2_X1 U164bar ( .A1(inbar[191]), .A2(inbar[189]), .ZN(n800bar);
  OR2_X1 U165 ( .A1(n799), .A2(n798), .ZN(n826) );
  AND2_X1 U165bar ( .A1(n799bar), .A2(n798bar), .ZN(n826bar);
  OR2_X1 U166 ( .A1(n797), .A2(n796), .ZN(n798) );
  AND2_X1 U166bar ( .A1(n797bar), .A2(n796bar), .ZN(n798bar);
  OR2_X1 U167 ( .A1(in[212]), .A2(in[193]), .ZN(n796) );
  AND2_X1 U167bar ( .A1(inbar[212]), .A2(inbar[193]), .ZN(n796bar);
  OR2_X1 U168 ( .A1(in[238]), .A2(n795), .ZN(n797) );
  AND2_X1 U168bar ( .A1(inbar[238]), .A2(n795bar), .ZN(n797bar);
  OR2_X1 U169 ( .A1(in[88]), .A2(in[247]), .ZN(n795) );
  AND2_X1 U169bar ( .A1(inbar[88]), .A2(inbar[247]), .ZN(n795bar);
  OR2_X1 U170 ( .A1(n794), .A2(n793), .ZN(n799) );
  AND2_X1 U170bar ( .A1(n794bar), .A2(n793bar), .ZN(n799bar);
  OR2_X1 U171 ( .A1(in[94]), .A2(in[92]), .ZN(n793) );
  AND2_X1 U171bar ( .A1(inbar[94]), .A2(inbar[92]), .ZN(n793bar);
  OR2_X1 U172 ( .A1(in_52), .A2(n792), .ZN(n794) );
  AND2_X1 U172bar ( .A1(in_52bar), .A2(n792bar), .ZN(n794bar);
  OR2_X1 U173 ( .A1(in_70), .A2(in_67), .ZN(n792) );
  AND2_X1 U173bar ( .A1(in_70bar), .A2(in_67bar), .ZN(n792bar);
  OR2_X1 U174 ( .A1(n791), .A2(n790), .ZN(out[2]) );
  AND2_X1 U174bar ( .A1(n791bar), .A2(n790bar), .ZN(outbar[2]);
  OR2_X1 U175 ( .A1(n789), .A2(n788), .ZN(n790) );
  AND2_X1 U175bar ( .A1(n789bar), .A2(n788bar), .ZN(n790bar);
  OR2_X1 U176 ( .A1(n787), .A2(n786), .ZN(n788) );
  AND2_X1 U176bar ( .A1(n787bar), .A2(n786bar), .ZN(n788bar);
  OR2_X1 U177 ( .A1(n819), .A2(n785), .ZN(n786) );
  AND2_X1 U177bar ( .A1(n819bar), .A2(n785bar), .ZN(n786bar);
  OR2_X1 U178 ( .A1(n784), .A2(n783), .ZN(n819) );
  AND2_X1 U178bar ( .A1(n784bar), .A2(n783bar), .ZN(n819bar);
  OR2_X1 U179 ( .A1(n782), .A2(n781), .ZN(n783) );
  AND2_X1 U179bar ( .A1(n782bar), .A2(n781bar), .ZN(n783bar);
  OR2_X1 U180 ( .A1(n780), .A2(n779), .ZN(n781) );
  AND2_X1 U180bar ( .A1(n780bar), .A2(n779bar), .ZN(n781bar);
  OR2_X1 U181 ( .A1(n962), .A2(n778), .ZN(n779) );
  AND2_X1 U181bar ( .A1(n962bar), .A2(n778bar), .ZN(n779bar);
  OR2_X1 U182 ( .A1(n777), .A2(n776), .ZN(n962) );
  AND2_X1 U182bar ( .A1(n777bar), .A2(n776bar), .ZN(n962bar);
  OR2_X1 U183 ( .A1(n775), .A2(n774), .ZN(n776) );
  AND2_X1 U183bar ( .A1(n775bar), .A2(n774bar), .ZN(n776bar);
  OR2_X1 U184 ( .A1(n773), .A2(n772), .ZN(n774) );
  AND2_X1 U184bar ( .A1(n773bar), .A2(n772bar), .ZN(n774bar);
  OR2_X1 U185 ( .A1(in[131]), .A2(in[120]), .ZN(n772) );
  AND2_X1 U185bar ( .A1(inbar[131]), .A2(inbar[120]), .ZN(n772bar);
  OR2_X1 U186 ( .A1(in[153]), .A2(in[147]), .ZN(n773) );
  AND2_X1 U186bar ( .A1(inbar[153]), .A2(inbar[147]), .ZN(n773bar);
  OR2_X1 U187 ( .A1(n771), .A2(n770), .ZN(n775) );
  AND2_X1 U187bar ( .A1(n771bar), .A2(n770bar), .ZN(n775bar);
  OR2_X1 U188 ( .A1(in[170]), .A2(in[156]), .ZN(n770) );
  AND2_X1 U188bar ( .A1(inbar[170]), .A2(inbar[156]), .ZN(n770bar);
  OR2_X1 U189 ( .A1(in[223]), .A2(in[190]), .ZN(n771) );
  AND2_X1 U189bar ( .A1(inbar[223]), .A2(inbar[190]), .ZN(n771bar);
  OR2_X1 U190 ( .A1(n769), .A2(n768), .ZN(n777) );
  AND2_X1 U190bar ( .A1(n769bar), .A2(n768bar), .ZN(n777bar);
  OR2_X1 U191 ( .A1(n767), .A2(n766), .ZN(n768) );
  AND2_X1 U191bar ( .A1(n767bar), .A2(n766bar), .ZN(n768bar);
  OR2_X1 U192 ( .A1(in[236]), .A2(in[230]), .ZN(n766) );
  AND2_X1 U192bar ( .A1(inbar[236]), .A2(inbar[230]), .ZN(n766bar);
  OR2_X1 U193 ( .A1(in[85]), .A2(in[240]), .ZN(n767) );
  AND2_X1 U193bar ( .A1(inbar[85]), .A2(inbar[240]), .ZN(n767bar);
  OR2_X1 U194 ( .A1(n765), .A2(n764), .ZN(n769) );
  AND2_X1 U194bar ( .A1(n765bar), .A2(n764bar), .ZN(n769bar);
  OR2_X1 U195 ( .A1(in_12), .A2(in[90]), .ZN(n764) );
  AND2_X1 U195bar ( .A1(in_12bar), .A2(inbar[90]), .ZN(n764bar);
  OR2_X1 U196 ( .A1(in_39), .A2(in_28), .ZN(n765) );
  AND2_X1 U196bar ( .A1(in_39bar), .A2(in_28bar), .ZN(n765bar);
  OR2_X1 U197 ( .A1(in[109]), .A2(n763), .ZN(n780) );
  AND2_X1 U197bar ( .A1(inbar[109]), .A2(n763bar), .ZN(n780bar);
  OR2_X1 U198 ( .A1(n762), .A2(n761), .ZN(n782) );
  AND2_X1 U198bar ( .A1(n762bar), .A2(n761bar), .ZN(n782bar);
  OR2_X1 U199 ( .A1(in[138]), .A2(in[129]), .ZN(n761) );
  AND2_X1 U199bar ( .A1(inbar[138]), .A2(inbar[129]), .ZN(n761bar);
  OR2_X1 U200 ( .A1(in[157]), .A2(n760), .ZN(n762) );
  AND2_X1 U200bar ( .A1(inbar[157]), .A2(n760bar), .ZN(n762bar);
  OR2_X1 U201 ( .A1(in[182]), .A2(in[167]), .ZN(n760) );
  AND2_X1 U201bar ( .A1(inbar[182]), .A2(inbar[167]), .ZN(n760bar);
  OR2_X1 U202 ( .A1(n759), .A2(n758), .ZN(n784) );
  AND2_X1 U202bar ( .A1(n759bar), .A2(n758bar), .ZN(n784bar);
  OR2_X1 U203 ( .A1(n757), .A2(n756), .ZN(n758) );
  AND2_X1 U203bar ( .A1(n757bar), .A2(n756bar), .ZN(n758bar);
  OR2_X1 U204 ( .A1(in[195]), .A2(in[184]), .ZN(n756) );
  AND2_X1 U204bar ( .A1(inbar[195]), .A2(inbar[184]), .ZN(n756bar);
  OR2_X1 U205 ( .A1(in[196]), .A2(n755), .ZN(n757) );
  AND2_X1 U205bar ( .A1(inbar[196]), .A2(n755bar), .ZN(n757bar);
  OR2_X1 U206 ( .A1(in[215]), .A2(in[209]), .ZN(n755) );
  AND2_X1 U206bar ( .A1(inbar[215]), .A2(inbar[209]), .ZN(n755bar);
  OR2_X1 U207 ( .A1(n754), .A2(n753), .ZN(n759) );
  AND2_X1 U207bar ( .A1(n754bar), .A2(n753bar), .ZN(n759bar);
  OR2_X1 U208 ( .A1(in[93]), .A2(in[233]), .ZN(n753) );
  AND2_X1 U208bar ( .A1(inbar[93]), .A2(inbar[233]), .ZN(n753bar);
  OR2_X1 U209 ( .A1(in_1), .A2(n752), .ZN(n754) );
  AND2_X1 U209bar ( .A1(in_1bar), .A2(n752bar), .ZN(n754bar);
  OR2_X1 U210 ( .A1(in_69), .A2(in_66), .ZN(n752) );
  AND2_X1 U210bar ( .A1(in_69bar), .A2(in_66bar), .ZN(n752bar);
  OR2_X1 U211 ( .A1(n966), .A2(n751), .ZN(n787) );
  AND2_X1 U211bar ( .A1(n966bar), .A2(n751bar), .ZN(n787bar);
  OR2_X1 U212 ( .A1(in[134]), .A2(n750), .ZN(n751) );
  AND2_X1 U212bar ( .A1(inbar[134]), .A2(n750bar), .ZN(n751bar);
  OR2_X1 U213 ( .A1(n749), .A2(n748), .ZN(n966) );
  AND2_X1 U213bar ( .A1(n749bar), .A2(n748bar), .ZN(n966bar);
  OR2_X1 U214 ( .A1(n747), .A2(n746), .ZN(n748) );
  AND2_X1 U214bar ( .A1(n747bar), .A2(n746bar), .ZN(n748bar);
  OR2_X1 U215 ( .A1(n745), .A2(n744), .ZN(n746) );
  AND2_X1 U215bar ( .A1(n745bar), .A2(n744bar), .ZN(n746bar);
  OR2_X1 U216 ( .A1(in[136]), .A2(in[121]), .ZN(n744) );
  AND2_X1 U216bar ( .A1(inbar[136]), .A2(inbar[121]), .ZN(n744bar);
  OR2_X1 U217 ( .A1(in[186]), .A2(in[174]), .ZN(n745) );
  AND2_X1 U217bar ( .A1(inbar[186]), .A2(inbar[174]), .ZN(n745bar);
  OR2_X1 U218 ( .A1(n743), .A2(n742), .ZN(n747) );
  AND2_X1 U218bar ( .A1(n743bar), .A2(n742bar), .ZN(n747bar);
  OR2_X1 U219 ( .A1(in[198]), .A2(in[197]), .ZN(n742) );
  AND2_X1 U219bar ( .A1(inbar[198]), .A2(inbar[197]), .ZN(n742bar);
  OR2_X1 U220 ( .A1(in[214]), .A2(in[199]), .ZN(n743) );
  AND2_X1 U220bar ( .A1(inbar[214]), .A2(inbar[199]), .ZN(n743bar);
  OR2_X1 U221 ( .A1(n741), .A2(n740), .ZN(n749) );
  AND2_X1 U221bar ( .A1(n741bar), .A2(n740bar), .ZN(n749bar);
  OR2_X1 U222 ( .A1(n739), .A2(n738), .ZN(n740) );
  AND2_X1 U222bar ( .A1(n739bar), .A2(n738bar), .ZN(n740bar);
  OR2_X1 U223 ( .A1(in[231]), .A2(in[220]), .ZN(n738) );
  AND2_X1 U223bar ( .A1(inbar[231]), .A2(inbar[220]), .ZN(n738bar);
  OR2_X1 U224 ( .A1(in_25), .A2(in[245]), .ZN(n739) );
  AND2_X1 U224bar ( .A1(in_25bar), .A2(inbar[245]), .ZN(n739bar);
  OR2_X1 U225 ( .A1(n737), .A2(n736), .ZN(n741) );
  AND2_X1 U225bar ( .A1(n737bar), .A2(n736bar), .ZN(n741bar);
  OR2_X1 U226 ( .A1(in_53), .A2(in_29), .ZN(n736) );
  AND2_X1 U226bar ( .A1(in_53bar), .A2(in_29bar), .ZN(n736bar);
  OR2_X1 U227 ( .A1(in_79), .A2(in_74), .ZN(n737) );
  AND2_X1 U227bar ( .A1(in_79bar), .A2(in_74bar), .ZN(n737bar);
  OR2_X1 U228 ( .A1(n735), .A2(n734), .ZN(n789) );
  AND2_X1 U228bar ( .A1(n735bar), .A2(n734bar), .ZN(n789bar);
  OR2_X1 U229 ( .A1(in[152]), .A2(in[140]), .ZN(n734) );
  AND2_X1 U229bar ( .A1(inbar[152]), .A2(inbar[140]), .ZN(n734bar);
  OR2_X1 U230 ( .A1(in[155]), .A2(n733), .ZN(n735) );
  AND2_X1 U230bar ( .A1(inbar[155]), .A2(n733bar), .ZN(n735bar);
  OR2_X1 U231 ( .A1(in[166]), .A2(in[165]), .ZN(n733) );
  AND2_X1 U231bar ( .A1(inbar[166]), .A2(inbar[165]), .ZN(n733bar);
  OR2_X1 U232 ( .A1(n732), .A2(n731), .ZN(n791) );
  AND2_X1 U232bar ( .A1(n732bar), .A2(n731bar), .ZN(n791bar);
  OR2_X1 U233 ( .A1(n730), .A2(n729), .ZN(n731) );
  AND2_X1 U233bar ( .A1(n730bar), .A2(n729bar), .ZN(n731bar);
  OR2_X1 U234 ( .A1(in[202]), .A2(in[185]), .ZN(n729) );
  AND2_X1 U234bar ( .A1(inbar[202]), .A2(inbar[185]), .ZN(n729bar);
  OR2_X1 U235 ( .A1(in[211]), .A2(n728), .ZN(n730) );
  AND2_X1 U235bar ( .A1(inbar[211]), .A2(n728bar), .ZN(n730bar);
  OR2_X1 U236 ( .A1(in[255]), .A2(in[253]), .ZN(n728) );
  AND2_X1 U236bar ( .A1(inbar[255]), .A2(inbar[253]), .ZN(n728bar);
  OR2_X1 U237 ( .A1(n727), .A2(n726), .ZN(n732) );
  AND2_X1 U237bar ( .A1(n727bar), .A2(n726bar), .ZN(n732bar);
  OR2_X1 U238 ( .A1(in_35), .A2(in_15), .ZN(n726) );
  AND2_X1 U238bar ( .A1(in_35bar), .A2(in_15bar), .ZN(n726bar);
  OR2_X1 U239 ( .A1(in_36), .A2(n725), .ZN(n727) );
  AND2_X1 U239bar ( .A1(in_36bar), .A2(n725bar), .ZN(n727bar);
  OR2_X1 U240 ( .A1(in_48), .A2(in_40), .ZN(n725) );
  AND2_X1 U240bar ( .A1(in_48bar), .A2(in_40bar), .ZN(n725bar);
  OR2_X1 U241 ( .A1(n724), .A2(n723), .ZN(out[1]) );
  AND2_X1 U241bar ( .A1(n724bar), .A2(n723bar), .ZN(outbar[1]);
  OR2_X1 U242 ( .A1(n722), .A2(n721), .ZN(n723) );
  AND2_X1 U242bar ( .A1(n722bar), .A2(n721bar), .ZN(n723bar);
  OR2_X1 U243 ( .A1(n720), .A2(n719), .ZN(n721) );
  AND2_X1 U243bar ( .A1(n720bar), .A2(n719bar), .ZN(n721bar);
  OR2_X1 U244 ( .A1(n921), .A2(n887), .ZN(n719) );
  AND2_X1 U244bar ( .A1(n921bar), .A2(n887bar), .ZN(n719bar);
  OR2_X1 U245 ( .A1(n718), .A2(n717), .ZN(n887) );
  AND2_X1 U245bar ( .A1(n718bar), .A2(n717bar), .ZN(n887bar);
  OR2_X1 U246 ( .A1(n716), .A2(n715), .ZN(n717) );
  AND2_X1 U246bar ( .A1(n716bar), .A2(n715bar), .ZN(n717bar);
  OR2_X1 U247 ( .A1(n714), .A2(n713), .ZN(n715) );
  AND2_X1 U247bar ( .A1(n714bar), .A2(n713bar), .ZN(n715bar);
  OR2_X1 U248 ( .A1(in[116]), .A2(in[110]), .ZN(n713) );
  AND2_X1 U248bar ( .A1(inbar[116]), .A2(inbar[110]), .ZN(n713bar);
  OR2_X1 U249 ( .A1(in[133]), .A2(in[130]), .ZN(n714) );
  AND2_X1 U249bar ( .A1(inbar[133]), .A2(inbar[130]), .ZN(n714bar);
  OR2_X1 U250 ( .A1(n712), .A2(n711), .ZN(n716) );
  AND2_X1 U250bar ( .A1(n712bar), .A2(n711bar), .ZN(n716bar);
  OR2_X1 U251 ( .A1(in[203]), .A2(in[135]), .ZN(n711) );
  AND2_X1 U251bar ( .A1(inbar[203]), .A2(inbar[135]), .ZN(n711bar);
  OR2_X1 U252 ( .A1(in[232]), .A2(in[223]), .ZN(n712) );
  AND2_X1 U252bar ( .A1(inbar[232]), .A2(inbar[223]), .ZN(n712bar);
  OR2_X1 U253 ( .A1(n710), .A2(n709), .ZN(n718) );
  AND2_X1 U253bar ( .A1(n710bar), .A2(n709bar), .ZN(n718bar);
  OR2_X1 U254 ( .A1(n708), .A2(n707), .ZN(n709) );
  AND2_X1 U254bar ( .A1(n708bar), .A2(n707bar), .ZN(n709bar);
  OR2_X1 U255 ( .A1(in[255]), .A2(in[233]), .ZN(n707) );
  AND2_X1 U255bar ( .A1(inbar[255]), .A2(inbar[233]), .ZN(n707bar);
  OR2_X1 U256 ( .A1(in_53), .A2(in_34), .ZN(n708) );
  AND2_X1 U256bar ( .A1(in_53bar), .A2(in_34bar), .ZN(n708bar);
  OR2_X1 U257 ( .A1(n706), .A2(n705), .ZN(n710) );
  AND2_X1 U257bar ( .A1(n706bar), .A2(n705bar), .ZN(n710bar);
  OR2_X1 U258 ( .A1(in_57), .A2(in_55), .ZN(n705) );
  AND2_X1 U258bar ( .A1(in_57bar), .A2(in_55bar), .ZN(n705bar);
  OR2_X1 U259 ( .A1(in_68), .A2(in_67), .ZN(n706) );
  AND2_X1 U259bar ( .A1(in_68bar), .A2(in_67bar), .ZN(n706bar);
  OR2_X1 U260 ( .A1(n704), .A2(n703), .ZN(n921) );
  AND2_X1 U260bar ( .A1(n704bar), .A2(n703bar), .ZN(n921bar);
  OR2_X1 U261 ( .A1(n702), .A2(n701), .ZN(n703) );
  AND2_X1 U261bar ( .A1(n702bar), .A2(n701bar), .ZN(n703bar);
  OR2_X1 U262 ( .A1(n700), .A2(n699), .ZN(n701) );
  AND2_X1 U262bar ( .A1(n700bar), .A2(n699bar), .ZN(n701bar);
  OR2_X1 U263 ( .A1(n944), .A2(n872), .ZN(n699) );
  AND2_X1 U263bar ( .A1(n944bar), .A2(n872bar), .ZN(n699bar);
  OR2_X1 U264 ( .A1(n698), .A2(n697), .ZN(n872) );
  AND2_X1 U264bar ( .A1(n698bar), .A2(n697bar), .ZN(n872bar);
  OR2_X1 U265 ( .A1(n696), .A2(n695), .ZN(n697) );
  AND2_X1 U265bar ( .A1(n696bar), .A2(n695bar), .ZN(n697bar);
  OR2_X1 U266 ( .A1(n694), .A2(n693), .ZN(n695) );
  AND2_X1 U266bar ( .A1(n694bar), .A2(n693bar), .ZN(n695bar);
  OR2_X1 U267 ( .A1(in[121]), .A2(in[102]), .ZN(n693) );
  AND2_X1 U267bar ( .A1(inbar[121]), .A2(inbar[102]), .ZN(n693bar);
  OR2_X1 U268 ( .A1(in[162]), .A2(in[161]), .ZN(n694) );
  AND2_X1 U268bar ( .A1(inbar[162]), .A2(inbar[161]), .ZN(n694bar);
  OR2_X1 U269 ( .A1(n692), .A2(n691), .ZN(n696) );
  AND2_X1 U269bar ( .A1(n692bar), .A2(n691bar), .ZN(n696bar);
  OR2_X1 U270 ( .A1(in[192]), .A2(in[178]), .ZN(n691) );
  AND2_X1 U270bar ( .A1(inbar[192]), .A2(inbar[178]), .ZN(n691bar);
  OR2_X1 U271 ( .A1(in[244]), .A2(in[209]), .ZN(n692) );
  AND2_X1 U271bar ( .A1(inbar[244]), .A2(inbar[209]), .ZN(n692bar);
  OR2_X1 U272 ( .A1(n690), .A2(n689), .ZN(n698) );
  AND2_X1 U272bar ( .A1(n690bar), .A2(n689bar), .ZN(n698bar);
  OR2_X1 U273 ( .A1(n688), .A2(n687), .ZN(n689) );
  AND2_X1 U273bar ( .A1(n688bar), .A2(n687bar), .ZN(n689bar);
  OR2_X1 U274 ( .A1(in[90]), .A2(in[254]), .ZN(n687) );
  AND2_X1 U274bar ( .A1(inbar[90]), .A2(inbar[254]), .ZN(n687bar);
  OR2_X1 U275 ( .A1(in_36), .A2(in_32), .ZN(n688) );
  AND2_X1 U275bar ( .A1(in_36bar), .A2(in_32bar), .ZN(n688bar);
  OR2_X1 U276 ( .A1(n686), .A2(n685), .ZN(n690) );
  AND2_X1 U276bar ( .A1(n686bar), .A2(n685bar), .ZN(n690bar);
  OR2_X1 U277 ( .A1(in_62), .A2(in_37), .ZN(n685) );
  AND2_X1 U277bar ( .A1(in_62bar), .A2(in_37bar), .ZN(n685bar);
  OR2_X1 U278 ( .A1(in_75), .A2(in_73), .ZN(n686) );
  AND2_X1 U278bar ( .A1(in_75bar), .A2(in_73bar), .ZN(n686bar);
  OR2_X1 U279 ( .A1(n684), .A2(n683), .ZN(n944) );
  AND2_X1 U279bar ( .A1(n684bar), .A2(n683bar), .ZN(n944bar);
  OR2_X1 U280 ( .A1(n682), .A2(n681), .ZN(n683) );
  AND2_X1 U280bar ( .A1(n682bar), .A2(n681bar), .ZN(n683bar);
  OR2_X1 U281 ( .A1(n680), .A2(n679), .ZN(n681) );
  AND2_X1 U281bar ( .A1(n680bar), .A2(n679bar), .ZN(n681bar);
  OR2_X1 U282 ( .A1(in[171]), .A2(in[153]), .ZN(n679) );
  AND2_X1 U282bar ( .A1(inbar[171]), .A2(inbar[153]), .ZN(n679bar);
  OR2_X1 U283 ( .A1(in[187]), .A2(in[176]), .ZN(n680) );
  AND2_X1 U283bar ( .A1(inbar[187]), .A2(inbar[176]), .ZN(n680bar);
  OR2_X1 U284 ( .A1(n678), .A2(n677), .ZN(n682) );
  AND2_X1 U284bar ( .A1(n678bar), .A2(n677bar), .ZN(n682bar);
  OR2_X1 U285 ( .A1(in[245]), .A2(in[211]), .ZN(n677) );
  AND2_X1 U285bar ( .A1(inbar[245]), .A2(inbar[211]), .ZN(n677bar);
  OR2_X1 U286 ( .A1(in[97]), .A2(in[88]), .ZN(n678) );
  AND2_X1 U286bar ( .A1(inbar[97]), .A2(inbar[88]), .ZN(n678bar);
  OR2_X1 U287 ( .A1(n676), .A2(n675), .ZN(n684) );
  AND2_X1 U287bar ( .A1(n676bar), .A2(n675bar), .ZN(n684bar);
  OR2_X1 U288 ( .A1(n674), .A2(n673), .ZN(n675) );
  AND2_X1 U288bar ( .A1(n674bar), .A2(n673bar), .ZN(n675bar);
  OR2_X1 U289 ( .A1(in_10), .A2(in_0), .ZN(n673) );
  AND2_X1 U289bar ( .A1(in_10bar), .A2(in_0bar), .ZN(n673bar);
  OR2_X1 U290 ( .A1(in_59), .A2(in_5), .ZN(n674) );
  AND2_X1 U290bar ( .A1(in_59bar), .A2(in_5bar), .ZN(n674bar);
  OR2_X1 U291 ( .A1(n672), .A2(n671), .ZN(n676) );
  AND2_X1 U291bar ( .A1(n672bar), .A2(n671bar), .ZN(n676bar);
  OR2_X1 U292 ( .A1(in_60), .A2(in_6), .ZN(n671) );
  AND2_X1 U292bar ( .A1(in_60bar), .A2(in_6bar), .ZN(n671bar);
  OR2_X1 U293 ( .A1(in_77), .A2(in_69), .ZN(n672) );
  AND2_X1 U293bar ( .A1(in_77bar), .A2(in_69bar), .ZN(n672bar);
  OR2_X1 U294 ( .A1(in[113]), .A2(n864), .ZN(n700) );
  AND2_X1 U294bar ( .A1(inbar[113]), .A2(n864bar), .ZN(n700bar);
  OR2_X1 U295 ( .A1(n670), .A2(n669), .ZN(n864) );
  AND2_X1 U295bar ( .A1(n670bar), .A2(n669bar), .ZN(n864bar);
  OR2_X1 U296 ( .A1(n668), .A2(n667), .ZN(n669) );
  AND2_X1 U296bar ( .A1(n668bar), .A2(n667bar), .ZN(n669bar);
  OR2_X1 U297 ( .A1(n666), .A2(n665), .ZN(n667) );
  AND2_X1 U297bar ( .A1(n666bar), .A2(n665bar), .ZN(n667bar);
  OR2_X1 U298 ( .A1(in[125]), .A2(in[107]), .ZN(n665) );
  AND2_X1 U298bar ( .A1(inbar[125]), .A2(inbar[107]), .ZN(n665bar);
  OR2_X1 U299 ( .A1(in[138]), .A2(in[126]), .ZN(n666) );
  AND2_X1 U299bar ( .A1(inbar[138]), .A2(inbar[126]), .ZN(n666bar);
  OR2_X1 U300 ( .A1(n664), .A2(n663), .ZN(n668) );
  AND2_X1 U300bar ( .A1(n664bar), .A2(n663bar), .ZN(n668bar);
  OR2_X1 U301 ( .A1(in[189]), .A2(in[143]), .ZN(n663) );
  AND2_X1 U301bar ( .A1(inbar[189]), .A2(inbar[143]), .ZN(n663bar);
  OR2_X1 U302 ( .A1(in[99]), .A2(in[214]), .ZN(n664) );
  AND2_X1 U302bar ( .A1(inbar[99]), .A2(inbar[214]), .ZN(n664bar);
  OR2_X1 U303 ( .A1(n662), .A2(n661), .ZN(n670) );
  AND2_X1 U303bar ( .A1(n662bar), .A2(n661bar), .ZN(n670bar);
  OR2_X1 U304 ( .A1(n660), .A2(n659), .ZN(n661) );
  AND2_X1 U304bar ( .A1(n660bar), .A2(n659bar), .ZN(n661bar);
  OR2_X1 U305 ( .A1(in_15), .A2(in_12), .ZN(n659) );
  AND2_X1 U305bar ( .A1(in_15bar), .A2(in_12bar), .ZN(n659bar);
  OR2_X1 U306 ( .A1(in_20), .A2(in_2), .ZN(n660) );
  AND2_X1 U306bar ( .A1(in_20bar), .A2(in_2bar), .ZN(n660bar);
  OR2_X1 U307 ( .A1(n658), .A2(n657), .ZN(n662) );
  AND2_X1 U307bar ( .A1(n658bar), .A2(n657bar), .ZN(n662bar);
  OR2_X1 U308 ( .A1(in_30), .A2(in_3), .ZN(n657) );
  AND2_X1 U308bar ( .A1(in_30bar), .A2(in_3bar), .ZN(n657bar);
  OR2_X1 U309 ( .A1(in_4), .A2(in_38), .ZN(n658) );
  AND2_X1 U309bar ( .A1(in_4bar), .A2(in_38bar), .ZN(n658bar);
  OR2_X1 U310 ( .A1(n656), .A2(n655), .ZN(n702) );
  AND2_X1 U310bar ( .A1(n656bar), .A2(n655bar), .ZN(n702bar);
  OR2_X1 U311 ( .A1(in[148]), .A2(in[137]), .ZN(n655) );
  AND2_X1 U311bar ( .A1(inbar[148]), .A2(inbar[137]), .ZN(n655bar);
  OR2_X1 U312 ( .A1(in[149]), .A2(n654), .ZN(n656) );
  AND2_X1 U312bar ( .A1(inbar[149]), .A2(n654bar), .ZN(n656bar);
  OR2_X1 U313 ( .A1(in[195]), .A2(in[190]), .ZN(n654) );
  AND2_X1 U313bar ( .A1(inbar[195]), .A2(inbar[190]), .ZN(n654bar);
  OR2_X1 U314 ( .A1(n653), .A2(n652), .ZN(n704) );
  AND2_X1 U314bar ( .A1(n653bar), .A2(n652bar), .ZN(n704bar);
  OR2_X1 U315 ( .A1(n651), .A2(n650), .ZN(n652) );
  AND2_X1 U315bar ( .A1(n651bar), .A2(n650bar), .ZN(n652bar);
  OR2_X1 U316 ( .A1(in[98]), .A2(in[197]), .ZN(n650) );
  AND2_X1 U316bar ( .A1(inbar[98]), .A2(inbar[197]), .ZN(n650bar);
  OR2_X1 U317 ( .A1(in_11), .A2(n649), .ZN(n651) );
  AND2_X1 U317bar ( .A1(in_11bar), .A2(n649bar), .ZN(n651bar);
  OR2_X1 U318 ( .A1(in_26), .A2(in_14), .ZN(n649) );
  AND2_X1 U318bar ( .A1(in_26bar), .A2(in_14bar), .ZN(n649bar);
  OR2_X1 U319 ( .A1(n648), .A2(n647), .ZN(n653) );
  AND2_X1 U319bar ( .A1(n648bar), .A2(n647bar), .ZN(n653bar);
  OR2_X1 U320 ( .A1(in_35), .A2(in_27), .ZN(n647) );
  AND2_X1 U320bar ( .A1(in_35bar), .A2(in_27bar), .ZN(n647bar);
  OR2_X1 U321 ( .A1(in_50), .A2(n646), .ZN(n648) );
  AND2_X1 U321bar ( .A1(in_50bar), .A2(n646bar), .ZN(n648bar);
  OR2_X1 U322 ( .A1(in_78), .A2(in_61), .ZN(n646) );
  AND2_X1 U322bar ( .A1(in_78bar), .A2(in_61bar), .ZN(n646bar);
  OR2_X1 U323 ( .A1(n942), .A2(n645), .ZN(n720) );
  AND2_X1 U323bar ( .A1(n942bar), .A2(n645bar), .ZN(n720bar);
  OR2_X1 U324 ( .A1(in[106]), .A2(n863), .ZN(n645) );
  AND2_X1 U324bar ( .A1(inbar[106]), .A2(n863bar), .ZN(n645bar);
  OR2_X1 U325 ( .A1(n644), .A2(n643), .ZN(n863) );
  AND2_X1 U325bar ( .A1(n644bar), .A2(n643bar), .ZN(n863bar);
  OR2_X1 U326 ( .A1(n642), .A2(n641), .ZN(n643) );
  AND2_X1 U326bar ( .A1(n642bar), .A2(n641bar), .ZN(n643bar);
  OR2_X1 U327 ( .A1(n640), .A2(n639), .ZN(n641) );
  AND2_X1 U327bar ( .A1(n640bar), .A2(n639bar), .ZN(n641bar);
  OR2_X1 U328 ( .A1(in[127]), .A2(in[122]), .ZN(n639) );
  AND2_X1 U328bar ( .A1(inbar[127]), .A2(inbar[122]), .ZN(n639bar);
  OR2_X1 U329 ( .A1(in[156]), .A2(in[132]), .ZN(n640) );
  AND2_X1 U329bar ( .A1(inbar[156]), .A2(inbar[132]), .ZN(n640bar);
  OR2_X1 U330 ( .A1(n638), .A2(n637), .ZN(n642) );
  AND2_X1 U330bar ( .A1(n638bar), .A2(n637bar), .ZN(n642bar);
  OR2_X1 U331 ( .A1(in[159]), .A2(in[157]), .ZN(n637) );
  AND2_X1 U331bar ( .A1(inbar[159]), .A2(inbar[157]), .ZN(n637bar);
  OR2_X1 U332 ( .A1(in[185]), .A2(in[169]), .ZN(n638) );
  AND2_X1 U332bar ( .A1(inbar[185]), .A2(inbar[169]), .ZN(n638bar);
  OR2_X1 U333 ( .A1(n636), .A2(n635), .ZN(n644) );
  AND2_X1 U333bar ( .A1(n636bar), .A2(n635bar), .ZN(n644bar);
  OR2_X1 U334 ( .A1(n634), .A2(n633), .ZN(n635) );
  AND2_X1 U334bar ( .A1(n634bar), .A2(n633bar), .ZN(n635bar);
  OR2_X1 U335 ( .A1(in[239]), .A2(in[218]), .ZN(n633) );
  AND2_X1 U335bar ( .A1(inbar[239]), .A2(inbar[218]), .ZN(n633bar);
  OR2_X1 U336 ( .A1(in_13), .A2(in[87]), .ZN(n634) );
  AND2_X1 U336bar ( .A1(in_13bar), .A2(inbar[87]), .ZN(n634bar);
  OR2_X1 U337 ( .A1(n632), .A2(n631), .ZN(n636) );
  AND2_X1 U337bar ( .A1(n632bar), .A2(n631bar), .ZN(n636bar);
  OR2_X1 U338 ( .A1(in_72), .A2(in_70), .ZN(n631) );
  AND2_X1 U338bar ( .A1(in_72bar), .A2(in_70bar), .ZN(n631bar);
  OR2_X1 U339 ( .A1(in_80), .A2(in_74), .ZN(n632) );
  AND2_X1 U339bar ( .A1(in_80bar), .A2(in_74bar), .ZN(n632bar);
  OR2_X1 U340 ( .A1(n630), .A2(n629), .ZN(n942) );
  AND2_X1 U340bar ( .A1(n630bar), .A2(n629bar), .ZN(n942bar);
  OR2_X1 U341 ( .A1(n628), .A2(n627), .ZN(n629) );
  AND2_X1 U341bar ( .A1(n628bar), .A2(n627bar), .ZN(n629bar);
  OR2_X1 U342 ( .A1(n626), .A2(n625), .ZN(n627) );
  AND2_X1 U342bar ( .A1(n626bar), .A2(n625bar), .ZN(n627bar);
  OR2_X1 U343 ( .A1(in[146]), .A2(in[100]), .ZN(n625) );
  AND2_X1 U343bar ( .A1(inbar[146]), .A2(inbar[100]), .ZN(n625bar);
  OR2_X1 U344 ( .A1(in[168]), .A2(in[152]), .ZN(n626) );
  AND2_X1 U344bar ( .A1(inbar[168]), .A2(inbar[152]), .ZN(n626bar);
  OR2_X1 U345 ( .A1(n624), .A2(n623), .ZN(n628) );
  AND2_X1 U345bar ( .A1(n624bar), .A2(n623bar), .ZN(n628bar);
  OR2_X1 U346 ( .A1(in[199]), .A2(in[182]), .ZN(n623) );
  AND2_X1 U346bar ( .A1(inbar[199]), .A2(inbar[182]), .ZN(n623bar);
  OR2_X1 U347 ( .A1(in[236]), .A2(in[204]), .ZN(n624) );
  AND2_X1 U347bar ( .A1(inbar[236]), .A2(inbar[204]), .ZN(n624bar);
  OR2_X1 U348 ( .A1(n622), .A2(n621), .ZN(n630) );
  AND2_X1 U348bar ( .A1(n622bar), .A2(n621bar), .ZN(n630bar);
  OR2_X1 U349 ( .A1(n620), .A2(n619), .ZN(n621) );
  AND2_X1 U349bar ( .A1(n620bar), .A2(n619bar), .ZN(n621bar);
  OR2_X1 U350 ( .A1(in[89]), .A2(in[246]), .ZN(n619) );
  AND2_X1 U350bar ( .A1(inbar[89]), .A2(inbar[246]), .ZN(n619bar);
  OR2_X1 U351 ( .A1(in[95]), .A2(in[92]), .ZN(n620) );
  AND2_X1 U351bar ( .A1(inbar[95]), .A2(inbar[92]), .ZN(n620bar);
  OR2_X1 U352 ( .A1(n618), .A2(n617), .ZN(n622) );
  AND2_X1 U352bar ( .A1(n618bar), .A2(n617bar), .ZN(n622bar);
  OR2_X1 U353 ( .A1(in_22), .A2(in_16), .ZN(n617) );
  AND2_X1 U353bar ( .A1(in_22bar), .A2(in_16bar), .ZN(n617bar);
  OR2_X1 U354 ( .A1(in_51), .A2(in_49), .ZN(n618) );
  AND2_X1 U354bar ( .A1(in_51bar), .A2(in_49bar), .ZN(n618bar);
  OR2_X1 U355 ( .A1(n616), .A2(n615), .ZN(n722) );
  AND2_X1 U355bar ( .A1(n616bar), .A2(n615bar), .ZN(n722bar);
  OR2_X1 U356 ( .A1(in[158]), .A2(in[115]), .ZN(n615) );
  AND2_X1 U356bar ( .A1(inbar[158]), .A2(inbar[115]), .ZN(n615bar);
  OR2_X1 U357 ( .A1(in[163]), .A2(n614), .ZN(n616) );
  AND2_X1 U357bar ( .A1(inbar[163]), .A2(n614bar), .ZN(n616bar);
  OR2_X1 U358 ( .A1(in[206]), .A2(in[165]), .ZN(n614) );
  AND2_X1 U358bar ( .A1(inbar[206]), .A2(inbar[165]), .ZN(n614bar);
  OR2_X1 U359 ( .A1(n613), .A2(n612), .ZN(n724) );
  AND2_X1 U359bar ( .A1(n613bar), .A2(n612bar), .ZN(n724bar);
  OR2_X1 U360 ( .A1(n611), .A2(n610), .ZN(n612) );
  AND2_X1 U360bar ( .A1(n611bar), .A2(n610bar), .ZN(n612bar);
  OR2_X1 U361 ( .A1(in[213]), .A2(in[207]), .ZN(n610) );
  AND2_X1 U361bar ( .A1(inbar[213]), .A2(inbar[207]), .ZN(n610bar);
  OR2_X1 U362 ( .A1(in[215]), .A2(n609), .ZN(n611) );
  AND2_X1 U362bar ( .A1(inbar[215]), .A2(n609bar), .ZN(n611bar);
  OR2_X1 U363 ( .A1(in[230]), .A2(in[220]), .ZN(n609) );
  AND2_X1 U363bar ( .A1(inbar[230]), .A2(inbar[220]), .ZN(n609bar);
  OR2_X1 U364 ( .A1(n608), .A2(n607), .ZN(n613) );
  AND2_X1 U364bar ( .A1(n608bar), .A2(n607bar), .ZN(n613bar);
  OR2_X1 U365 ( .A1(in[251]), .A2(in[234]), .ZN(n607) );
  AND2_X1 U365bar ( .A1(inbar[251]), .A2(inbar[234]), .ZN(n607bar);
  OR2_X1 U366 ( .A1(in_17), .A2(n606), .ZN(n608) );
  AND2_X1 U366bar ( .A1(in_17bar), .A2(n606bar), .ZN(n608bar);
  OR2_X1 U367 ( .A1(in_65), .A2(in_56), .ZN(n606) );
  AND2_X1 U367bar ( .A1(in_65bar), .A2(in_56bar), .ZN(n606bar);
  OR2_X1 U368 ( .A1(n605), .A2(n604), .ZN(out[0]) );
  AND2_X1 U368bar ( .A1(n605bar), .A2(n604bar), .ZN(outbar[0]);
  OR2_X1 U369 ( .A1(n603), .A2(n602), .ZN(n604) );
  AND2_X1 U369bar ( .A1(n603bar), .A2(n602bar), .ZN(n604bar);
  OR2_X1 U370 ( .A1(n601), .A2(n600), .ZN(n602) );
  AND2_X1 U370bar ( .A1(n601bar), .A2(n600bar), .ZN(n602bar);
  OR2_X1 U371 ( .A1(n820), .A2(n785), .ZN(n600) );
  AND2_X1 U371bar ( .A1(n820bar), .A2(n785bar), .ZN(n600bar);
  OR2_X1 U372 ( .A1(n599), .A2(n598), .ZN(n785) );
  AND2_X1 U372bar ( .A1(n599bar), .A2(n598bar), .ZN(n785bar);
  OR2_X1 U373 ( .A1(n597), .A2(n596), .ZN(n598) );
  AND2_X1 U373bar ( .A1(n597bar), .A2(n596bar), .ZN(n598bar);
  OR2_X1 U374 ( .A1(n595), .A2(n594), .ZN(n596) );
  AND2_X1 U374bar ( .A1(n595bar), .A2(n594bar), .ZN(n596bar);
  OR2_X1 U375 ( .A1(in[135]), .A2(in[104]), .ZN(n594) );
  AND2_X1 U375bar ( .A1(inbar[135]), .A2(inbar[104]), .ZN(n594bar);
  OR2_X1 U376 ( .A1(in[188]), .A2(in[178]), .ZN(n595) );
  AND2_X1 U376bar ( .A1(inbar[188]), .A2(inbar[178]), .ZN(n595bar);
  OR2_X1 U377 ( .A1(n593), .A2(n592), .ZN(n597) );
  AND2_X1 U377bar ( .A1(n593bar), .A2(n592bar), .ZN(n597bar);
  OR2_X1 U378 ( .A1(in[217]), .A2(in[194]), .ZN(n592) );
  AND2_X1 U378bar ( .A1(inbar[217]), .A2(inbar[194]), .ZN(n592bar);
  OR2_X1 U379 ( .A1(in[237]), .A2(in[218]), .ZN(n593) );
  AND2_X1 U379bar ( .A1(inbar[237]), .A2(inbar[218]), .ZN(n593bar);
  OR2_X1 U380 ( .A1(n591), .A2(n590), .ZN(n599) );
  AND2_X1 U380bar ( .A1(n591bar), .A2(n590bar), .ZN(n599bar);
  OR2_X1 U381 ( .A1(n589), .A2(n588), .ZN(n590) );
  AND2_X1 U381bar ( .A1(n589bar), .A2(n588bar), .ZN(n590bar);
  OR2_X1 U382 ( .A1(in_2), .A2(in_10), .ZN(n588) );
  AND2_X1 U382bar ( .A1(in_2bar), .A2(in_10bar), .ZN(n588bar);
  OR2_X1 U383 ( .A1(in_47), .A2(in_22), .ZN(n589) );
  AND2_X1 U383bar ( .A1(in_47bar), .A2(in_22bar), .ZN(n589bar);
  OR2_X1 U384 ( .A1(n587), .A2(n586), .ZN(n591) );
  AND2_X1 U384bar ( .A1(n587bar), .A2(n586bar), .ZN(n591bar);
  OR2_X1 U385 ( .A1(in_56), .A2(in_54), .ZN(n586) );
  AND2_X1 U385bar ( .A1(in_56bar), .A2(in_54bar), .ZN(n586bar);
  OR2_X1 U386 ( .A1(in_63), .A2(in_61), .ZN(n587) );
  AND2_X1 U386bar ( .A1(in_63bar), .A2(in_61bar), .ZN(n587bar);
  OR2_X1 U387 ( .A1(n585), .A2(n584), .ZN(n820) );
  AND2_X1 U387bar ( .A1(n585bar), .A2(n584bar), .ZN(n820bar);
  OR2_X1 U388 ( .A1(n583), .A2(n582), .ZN(n584) );
  AND2_X1 U388bar ( .A1(n583bar), .A2(n582bar), .ZN(n584bar);
  OR2_X1 U389 ( .A1(n581), .A2(n580), .ZN(n582) );
  AND2_X1 U389bar ( .A1(n581bar), .A2(n580bar), .ZN(n582bar);
  OR2_X1 U390 ( .A1(in[158]), .A2(in[142]), .ZN(n580) );
  AND2_X1 U390bar ( .A1(inbar[158]), .A2(inbar[142]), .ZN(n580bar);
  OR2_X1 U391 ( .A1(in[175]), .A2(in[164]), .ZN(n581) );
  AND2_X1 U391bar ( .A1(inbar[175]), .A2(inbar[164]), .ZN(n581bar);
  OR2_X1 U392 ( .A1(n579), .A2(n578), .ZN(n583) );
  AND2_X1 U392bar ( .A1(n579bar), .A2(n578bar), .ZN(n583bar);
  OR2_X1 U393 ( .A1(in[228]), .A2(in[204]), .ZN(n578) );
  AND2_X1 U393bar ( .A1(inbar[228]), .A2(inbar[204]), .ZN(n578bar);
  OR2_X1 U394 ( .A1(in[91]), .A2(in[87]), .ZN(n579) );
  AND2_X1 U394bar ( .A1(inbar[91]), .A2(inbar[87]), .ZN(n579bar);
  OR2_X1 U395 ( .A1(n577), .A2(n576), .ZN(n585) );
  AND2_X1 U395bar ( .A1(n577bar), .A2(n576bar), .ZN(n585bar);
  OR2_X1 U396 ( .A1(n575), .A2(n574), .ZN(n576) );
  AND2_X1 U396bar ( .A1(n575bar), .A2(n574bar), .ZN(n576bar);
  OR2_X1 U397 ( .A1(in_21), .A2(in_11), .ZN(n574) );
  AND2_X1 U397bar ( .A1(in_21bar), .A2(in_11bar), .ZN(n574bar);
  OR2_X1 U398 ( .A1(in_5), .A2(in_3), .ZN(n575) );
  AND2_X1 U398bar ( .A1(in_5bar), .A2(in_3bar), .ZN(n575bar);
  OR2_X1 U399 ( .A1(n573), .A2(n572), .ZN(n577) );
  AND2_X1 U399bar ( .A1(n573bar), .A2(n572bar), .ZN(n577bar);
  OR2_X1 U400 ( .A1(in_68), .A2(in_64), .ZN(n572) );
  AND2_X1 U400bar ( .A1(in_68bar), .A2(in_64bar), .ZN(n572bar);
  OR2_X1 U401 ( .A1(in_76), .A2(in_73), .ZN(n573) );
  AND2_X1 U401bar ( .A1(in_76bar), .A2(in_73bar), .ZN(n573bar);
  OR2_X1 U402 ( .A1(n778), .A2(n571), .ZN(n601) );
  AND2_X1 U402bar ( .A1(n778bar), .A2(n571bar), .ZN(n601bar);
  OR2_X1 U403 ( .A1(in[100]), .A2(n965), .ZN(n571) );
  AND2_X1 U403bar ( .A1(inbar[100]), .A2(n965bar), .ZN(n571bar);
  OR2_X1 U404 ( .A1(n570), .A2(n569), .ZN(n965) );
  AND2_X1 U404bar ( .A1(n570bar), .A2(n569bar), .ZN(n965bar);
  OR2_X1 U405 ( .A1(n568), .A2(n567), .ZN(n569) );
  AND2_X1 U405bar ( .A1(n568bar), .A2(n567bar), .ZN(n569bar);
  OR2_X1 U406 ( .A1(n566), .A2(n565), .ZN(n567) );
  AND2_X1 U406bar ( .A1(n566bar), .A2(n565bar), .ZN(n567bar);
  OR2_X1 U407 ( .A1(n817), .A2(n750), .ZN(n565) );
  AND2_X1 U407bar ( .A1(n817bar), .A2(n750bar), .ZN(n565bar);
  OR2_X1 U408 ( .A1(n564), .A2(n563), .ZN(n750) );
  AND2_X1 U408bar ( .A1(n564bar), .A2(n563bar), .ZN(n750bar);
  OR2_X1 U409 ( .A1(n562), .A2(n561), .ZN(n563) );
  AND2_X1 U409bar ( .A1(n562bar), .A2(n561bar), .ZN(n563bar);
  OR2_X1 U410 ( .A1(n560), .A2(n559), .ZN(n561) );
  AND2_X1 U410bar ( .A1(n560bar), .A2(n559bar), .ZN(n561bar);
  OR2_X1 U411 ( .A1(in[119]), .A2(in[103]), .ZN(n559) );
  AND2_X1 U411bar ( .A1(inbar[119]), .A2(inbar[103]), .ZN(n559bar);
  OR2_X1 U412 ( .A1(in[137]), .A2(in[133]), .ZN(n560) );
  AND2_X1 U412bar ( .A1(inbar[137]), .A2(inbar[133]), .ZN(n560bar);
  OR2_X1 U413 ( .A1(n558), .A2(n557), .ZN(n562) );
  AND2_X1 U413bar ( .A1(n558bar), .A2(n557bar), .ZN(n562bar);
  OR2_X1 U414 ( .A1(in[176]), .A2(in[173]), .ZN(n557) );
  AND2_X1 U414bar ( .A1(inbar[176]), .A2(inbar[173]), .ZN(n557bar);
  OR2_X1 U415 ( .A1(in[210]), .A2(in[181]), .ZN(n558) );
  AND2_X1 U415bar ( .A1(inbar[210]), .A2(inbar[181]), .ZN(n558bar);
  OR2_X1 U416 ( .A1(n556), .A2(n555), .ZN(n564) );
  AND2_X1 U416bar ( .A1(n556bar), .A2(n555bar), .ZN(n564bar);
  OR2_X1 U417 ( .A1(n554), .A2(n553), .ZN(n555) );
  AND2_X1 U417bar ( .A1(n554bar), .A2(n553bar), .ZN(n555bar);
  OR2_X1 U418 ( .A1(in_13), .A2(in[234]), .ZN(n553) );
  AND2_X1 U418bar ( .A1(in_13bar), .A2(inbar[234]), .ZN(n553bar);
  OR2_X1 U419 ( .A1(in_38), .A2(in_32), .ZN(n554) );
  AND2_X1 U419bar ( .A1(in_38bar), .A2(in_32bar), .ZN(n554bar);
  OR2_X1 U420 ( .A1(n552), .A2(n551), .ZN(n556) );
  AND2_X1 U420bar ( .A1(n552bar), .A2(n551bar), .ZN(n556bar);
  OR2_X1 U421 ( .A1(in_42), .A2(in_41), .ZN(n551) );
  AND2_X1 U421bar ( .A1(in_42bar), .A2(in_41bar), .ZN(n551bar);
  OR2_X1 U422 ( .A1(in_7), .A2(in_49), .ZN(n552) );
  AND2_X1 U422bar ( .A1(in_7bar), .A2(in_49bar), .ZN(n552bar);
  OR2_X1 U423 ( .A1(n550), .A2(n549), .ZN(n817) );
  AND2_X1 U423bar ( .A1(n550bar), .A2(n549bar), .ZN(n817bar);
  OR2_X1 U424 ( .A1(n548), .A2(n547), .ZN(n549) );
  AND2_X1 U424bar ( .A1(n548bar), .A2(n547bar), .ZN(n549bar);
  OR2_X1 U425 ( .A1(n546), .A2(n545), .ZN(n547) );
  AND2_X1 U425bar ( .A1(n546bar), .A2(n545bar), .ZN(n547bar);
  OR2_X1 U426 ( .A1(in[159]), .A2(in[105]), .ZN(n545) );
  AND2_X1 U426bar ( .A1(inbar[159]), .A2(inbar[105]), .ZN(n545bar);
  OR2_X1 U427 ( .A1(in[206]), .A2(in[183]), .ZN(n546) );
  AND2_X1 U427bar ( .A1(inbar[206]), .A2(inbar[183]), .ZN(n546bar);
  OR2_X1 U428 ( .A1(n544), .A2(n543), .ZN(n548) );
  AND2_X1 U428bar ( .A1(n544bar), .A2(n543bar), .ZN(n548bar);
  OR2_X1 U429 ( .A1(in[229]), .A2(in[219]), .ZN(n543) );
  AND2_X1 U429bar ( .A1(inbar[229]), .A2(inbar[219]), .ZN(n543bar);
  OR2_X1 U430 ( .A1(in[235]), .A2(in[232]), .ZN(n544) );
  AND2_X1 U430bar ( .A1(inbar[235]), .A2(inbar[232]), .ZN(n544bar);
  OR2_X1 U431 ( .A1(n542), .A2(n541), .ZN(n550) );
  AND2_X1 U431bar ( .A1(n542bar), .A2(n541bar), .ZN(n550bar);
  OR2_X1 U432 ( .A1(n540), .A2(n539), .ZN(n541) );
  AND2_X1 U432bar ( .A1(n540bar), .A2(n539bar), .ZN(n541bar);
  OR2_X1 U433 ( .A1(in[249]), .A2(in[242]), .ZN(n539) );
  AND2_X1 U433bar ( .A1(inbar[249]), .A2(inbar[242]), .ZN(n539bar);
  OR2_X1 U434 ( .A1(in[89]), .A2(in[254]), .ZN(n540) );
  AND2_X1 U434bar ( .A1(inbar[89]), .A2(inbar[254]), .ZN(n540bar);
  OR2_X1 U435 ( .A1(n538), .A2(n537), .ZN(n542) );
  AND2_X1 U435bar ( .A1(n538bar), .A2(n537bar), .ZN(n542bar);
  OR2_X1 U436 ( .A1(in_14), .A2(in[99]), .ZN(n537) );
  AND2_X1 U436bar ( .A1(in_14bar), .A2(inbar[99]), .ZN(n537bar);
  OR2_X1 U437 ( .A1(in_60), .A2(in_18), .ZN(n538) );
  AND2_X1 U437bar ( .A1(in_60bar), .A2(in_18bar), .ZN(n538bar);
  OR2_X1 U438 ( .A1(in[113]), .A2(n763), .ZN(n566) );
  AND2_X1 U438bar ( .A1(inbar[113]), .A2(n763bar), .ZN(n566bar);
  OR2_X1 U439 ( .A1(n536), .A2(n535), .ZN(n763) );
  AND2_X1 U439bar ( .A1(n536bar), .A2(n535bar), .ZN(n763bar);
  OR2_X1 U440 ( .A1(n534), .A2(n533), .ZN(n535) );
  AND2_X1 U440bar ( .A1(n534bar), .A2(n533bar), .ZN(n535bar);
  OR2_X1 U441 ( .A1(n532), .A2(n531), .ZN(n533) );
  AND2_X1 U441bar ( .A1(n532bar), .A2(n531bar), .ZN(n533bar);
  OR2_X1 U442 ( .A1(in[115]), .A2(in[110]), .ZN(n531) );
  AND2_X1 U442bar ( .A1(inbar[115]), .A2(inbar[110]), .ZN(n531bar);
  OR2_X1 U443 ( .A1(in[125]), .A2(in[117]), .ZN(n532) );
  AND2_X1 U443bar ( .A1(inbar[125]), .A2(inbar[117]), .ZN(n532bar);
  OR2_X1 U444 ( .A1(n530), .A2(n529), .ZN(n534) );
  AND2_X1 U444bar ( .A1(n530bar), .A2(n529bar), .ZN(n534bar);
  OR2_X1 U445 ( .A1(in[180]), .A2(in[128]), .ZN(n529) );
  AND2_X1 U445bar ( .A1(inbar[180]), .A2(inbar[128]), .ZN(n529bar);
  OR2_X1 U446 ( .A1(in[205]), .A2(in[201]), .ZN(n530) );
  AND2_X1 U446bar ( .A1(inbar[205]), .A2(inbar[201]), .ZN(n530bar);
  OR2_X1 U447 ( .A1(n528), .A2(n527), .ZN(n536) );
  AND2_X1 U447bar ( .A1(n528bar), .A2(n527bar), .ZN(n536bar);
  OR2_X1 U448 ( .A1(n526), .A2(n525), .ZN(n527) );
  AND2_X1 U448bar ( .A1(n526bar), .A2(n525bar), .ZN(n527bar);
  OR2_X1 U449 ( .A1(in[244]), .A2(in[239]), .ZN(n525) );
  AND2_X1 U449bar ( .A1(inbar[244]), .A2(inbar[239]), .ZN(n525bar);
  OR2_X1 U450 ( .A1(in[95]), .A2(in[83]), .ZN(n526) );
  AND2_X1 U450bar ( .A1(inbar[95]), .A2(inbar[83]), .ZN(n526bar);
  OR2_X1 U451 ( .A1(n524), .A2(n523), .ZN(n528) );
  AND2_X1 U451bar ( .A1(n524bar), .A2(n523bar), .ZN(n528bar);
  OR2_X1 U452 ( .A1(in_24), .A2(in[97]), .ZN(n523) );
  AND2_X1 U452bar ( .A1(in_24bar), .A2(inbar[97]), .ZN(n523bar);
  OR2_X1 U453 ( .A1(in_33), .A2(in_27), .ZN(n524) );
  AND2_X1 U453bar ( .A1(in_33bar), .A2(in_27bar), .ZN(n524bar);
  OR2_X1 U454 ( .A1(n522), .A2(n521), .ZN(n568) );
  AND2_X1 U454bar ( .A1(n522bar), .A2(n521bar), .ZN(n568bar);
  OR2_X1 U455 ( .A1(in[145]), .A2(in[126]), .ZN(n521) );
  AND2_X1 U455bar ( .A1(inbar[145]), .A2(inbar[126]), .ZN(n521bar);
  OR2_X1 U456 ( .A1(in[169]), .A2(n520), .ZN(n522) );
  AND2_X1 U456bar ( .A1(inbar[169]), .A2(n520bar), .ZN(n522bar);
  OR2_X1 U457 ( .A1(in[221]), .A2(in[172]), .ZN(n520) );
  AND2_X1 U457bar ( .A1(inbar[221]), .A2(inbar[172]), .ZN(n520bar);
  OR2_X1 U458 ( .A1(n519), .A2(n518), .ZN(n570) );
  AND2_X1 U458bar ( .A1(n519bar), .A2(n518bar), .ZN(n570bar);
  OR2_X1 U459 ( .A1(n517), .A2(n516), .ZN(n518) );
  AND2_X1 U459bar ( .A1(n517bar), .A2(n516bar), .ZN(n518bar);
  OR2_X1 U460 ( .A1(in[241]), .A2(in[224]), .ZN(n516) );
  AND2_X1 U460bar ( .A1(inbar[241]), .A2(inbar[224]), .ZN(n516bar);
  OR2_X1 U461 ( .A1(in[86]), .A2(n515), .ZN(n517) );
  AND2_X1 U461bar ( .A1(inbar[86]), .A2(n515bar), .ZN(n517bar);
  OR2_X1 U462 ( .A1(in_43), .A2(in_34), .ZN(n515) );
  AND2_X1 U462bar ( .A1(in_43bar), .A2(in_34bar), .ZN(n515bar);
  OR2_X1 U463 ( .A1(n514), .A2(n513), .ZN(n519) );
  AND2_X1 U463bar ( .A1(n514bar), .A2(n513bar), .ZN(n519bar);
  OR2_X1 U464 ( .A1(in_65), .A2(in_51), .ZN(n513) );
  AND2_X1 U464bar ( .A1(in_65bar), .A2(in_51bar), .ZN(n513bar);
  OR2_X1 U465 ( .A1(in_75), .A2(n512), .ZN(n514) );
  AND2_X1 U465bar ( .A1(in_75bar), .A2(n512bar), .ZN(n514bar);
  OR2_X1 U466 ( .A1(in_81), .A2(in_77), .ZN(n512) );
  AND2_X1 U466bar ( .A1(in_81bar), .A2(in_77bar), .ZN(n512bar);
  OR2_X1 U467 ( .A1(n511), .A2(n510), .ZN(n778) );
  AND2_X1 U467bar ( .A1(n511bar), .A2(n510bar), .ZN(n778bar);
  OR2_X1 U468 ( .A1(n509), .A2(n508), .ZN(n510) );
  AND2_X1 U468bar ( .A1(n509bar), .A2(n508bar), .ZN(n510bar);
  OR2_X1 U469 ( .A1(n507), .A2(n506), .ZN(n508) );
  AND2_X1 U469bar ( .A1(n507bar), .A2(n506bar), .ZN(n508bar);
  OR2_X1 U470 ( .A1(in[107]), .A2(in[101]), .ZN(n506) );
  AND2_X1 U470bar ( .A1(inbar[107]), .A2(inbar[101]), .ZN(n506bar);
  OR2_X1 U471 ( .A1(in[139]), .A2(in[132]), .ZN(n507) );
  AND2_X1 U471bar ( .A1(inbar[139]), .A2(inbar[132]), .ZN(n507bar);
  OR2_X1 U472 ( .A1(n505), .A2(n504), .ZN(n509) );
  AND2_X1 U472bar ( .A1(n505bar), .A2(n504bar), .ZN(n509bar);
  OR2_X1 U473 ( .A1(in[146]), .A2(in[141]), .ZN(n504) );
  AND2_X1 U473bar ( .A1(inbar[146]), .A2(inbar[141]), .ZN(n504bar);
  OR2_X1 U474 ( .A1(in[203]), .A2(in[179]), .ZN(n505) );
  AND2_X1 U474bar ( .A1(inbar[203]), .A2(inbar[179]), .ZN(n505bar);
  OR2_X1 U475 ( .A1(n503), .A2(n502), .ZN(n511) );
  AND2_X1 U475bar ( .A1(n503bar), .A2(n502bar), .ZN(n511bar);
  OR2_X1 U476 ( .A1(n501), .A2(n500), .ZN(n502) );
  AND2_X1 U476bar ( .A1(n501bar), .A2(n500bar), .ZN(n502bar);
  OR2_X1 U477 ( .A1(in[243]), .A2(in[222]), .ZN(n500) );
  AND2_X1 U477bar ( .A1(inbar[243]), .A2(inbar[222]), .ZN(n500bar);
  OR2_X1 U478 ( .A1(in[251]), .A2(in[250]), .ZN(n501) );
  AND2_X1 U478bar ( .A1(inbar[251]), .A2(inbar[250]), .ZN(n501bar);
  OR2_X1 U479 ( .A1(n499), .A2(n498), .ZN(n503) );
  AND2_X1 U479bar ( .A1(n499bar), .A2(n498bar), .ZN(n503bar);
  OR2_X1 U480 ( .A1(in_37), .A2(in_19), .ZN(n498) );
  AND2_X1 U480bar ( .A1(in_37bar), .A2(in_19bar), .ZN(n498bar);
  OR2_X1 U481 ( .A1(in_78), .A2(in_6), .ZN(n499) );
  AND2_X1 U481bar ( .A1(in_78bar), .A2(in_6bar), .ZN(n499bar);
  OR2_X1 U482 ( .A1(n497), .A2(n496), .ZN(n603) );
  AND2_X1 U482bar ( .A1(n497bar), .A2(n496bar), .ZN(n603bar);
  OR2_X1 U483 ( .A1(in[112]), .A2(in[102]), .ZN(n496) );
  AND2_X1 U483bar ( .A1(inbar[112]), .A2(inbar[102]), .ZN(n496bar);
  OR2_X1 U484 ( .A1(in[123]), .A2(n495), .ZN(n497) );
  AND2_X1 U484bar ( .A1(inbar[123]), .A2(n495bar), .ZN(n497bar);
  OR2_X1 U485 ( .A1(in[143]), .A2(in[130]), .ZN(n495) );
  AND2_X1 U485bar ( .A1(inbar[143]), .A2(inbar[130]), .ZN(n495bar);
  OR2_X1 U486 ( .A1(n494), .A2(n493), .ZN(n605) );
  AND2_X1 U486bar ( .A1(n494bar), .A2(n493bar), .ZN(n605bar);
  OR2_X1 U487 ( .A1(n492), .A2(n491), .ZN(n493) );
  AND2_X1 U487bar ( .A1(n492bar), .A2(n491bar), .ZN(n493bar);
  OR2_X1 U488 ( .A1(in[216]), .A2(in[213]), .ZN(n491) );
  AND2_X1 U488bar ( .A1(inbar[216]), .A2(inbar[213]), .ZN(n491bar);
  OR2_X1 U489 ( .A1(in[227]), .A2(n490), .ZN(n492) );
  AND2_X1 U489bar ( .A1(inbar[227]), .A2(n490bar), .ZN(n492bar);
  OR2_X1 U490 ( .A1(in_0), .A2(in[248]), .ZN(n490) );
  AND2_X1 U490bar ( .A1(in_0bar), .A2(inbar[248]), .ZN(n490bar);
  OR2_X1 U491 ( .A1(n489), .A2(n488), .ZN(n494) );
  AND2_X1 U491bar ( .A1(n489bar), .A2(n488bar), .ZN(n494bar);
  OR2_X1 U492 ( .A1(in_46), .A2(in_44), .ZN(n488) );
  AND2_X1 U492bar ( .A1(in_46bar), .A2(in_44bar), .ZN(n488bar);
  OR2_X1 U493 ( .A1(in_50), .A2(n487), .ZN(n489) );
  AND2_X1 U493bar ( .A1(in_50bar), .A2(n487bar), .ZN(n489bar);
  OR2_X1 U494 ( .A1(in_9), .A2(in_80), .ZN(n487) );
  AND2_X1 U494bar ( .A1(in_9bar), .A2(in_80bar), .ZN(n487bar);
endmodule




module sBox_2 ( in, out );
  input [7:0] in;
  //input_done

  output [7:0] out;
  //output_done

  wire   [255:0] decodeOut;
  //wire_done

  decode_2 dec ( .in(in), .out(decodeOut) );
  encode_2 enc ( .in(decodeOut), .out(out) );
endmodule


module CD2_9 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_10 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_11 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_12 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD4_5 ( a, b, y );
  input [3:0] a;
  input [3:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  //input_done

  output [15:0] y;
  reg [15:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]);
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]);
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]);
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]);
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]);
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]);
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]);
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]);
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]);
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]);
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]);
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]);
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]);
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]);
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]);
endmodule




module CD4_6 ( a, b, y );
  input [3:0] a;
  input [3:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  //input_done

  output [15:0] y;
  reg [15:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]);
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]);
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]);
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]);
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]);
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]);
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]);
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]);
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]);
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]);
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]);
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]);
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]);
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]);
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]);
endmodule




module CD16_3 ( a, b, y );
  input [15:0] a;
  input [15:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign abar[8] = ~a[8];
  assign abar[9] = ~a[9];
  assign abar[10] = ~a[10];
  assign abar[11] = ~a[11];
  assign abar[12] = ~a[12];
  assign abar[13] = ~a[13];
  assign abar[14] = ~a[14];
  assign abar[15] = ~a[15];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign bbar[8] = ~b[8];
  assign bbar[9] = ~b[9];
  assign bbar[10] = ~b[10];
  assign bbar[11] = ~b[11];
  assign bbar[12] = ~b[12];
  assign bbar[13] = ~b[13];
  assign bbar[14] = ~b[14];
  assign bbar[15] = ~b[15];
  //input_done

  output [255:0] y;
  reg [255:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[9]), .A2(a[0]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[9]), .A2(abar[0]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[3]), .A2(a[6]), .ZN(y[99]) );
  OR2_X1 U2bar ( .A1(bbar[3]), .A2(abar[6]), .ZN(ybar[99]);
  AND2_X1 U3 ( .A1(b[2]), .A2(a[6]), .ZN(y[98]) );
  OR2_X1 U3bar ( .A1(bbar[2]), .A2(abar[6]), .ZN(ybar[98]);
  AND2_X1 U4 ( .A1(b[1]), .A2(a[6]), .ZN(y[97]) );
  OR2_X1 U4bar ( .A1(bbar[1]), .A2(abar[6]), .ZN(ybar[97]);
  AND2_X1 U5 ( .A1(b[0]), .A2(a[6]), .ZN(y[96]) );
  OR2_X1 U5bar ( .A1(bbar[0]), .A2(abar[6]), .ZN(ybar[96]);
  AND2_X1 U6 ( .A1(b[15]), .A2(a[5]), .ZN(y[95]) );
  OR2_X1 U6bar ( .A1(bbar[15]), .A2(abar[5]), .ZN(ybar[95]);
  AND2_X1 U7 ( .A1(b[14]), .A2(a[5]), .ZN(y[94]) );
  OR2_X1 U7bar ( .A1(bbar[14]), .A2(abar[5]), .ZN(ybar[94]);
  AND2_X1 U8 ( .A1(b[13]), .A2(a[5]), .ZN(y[93]) );
  OR2_X1 U8bar ( .A1(bbar[13]), .A2(abar[5]), .ZN(ybar[93]);
  AND2_X1 U9 ( .A1(b[12]), .A2(a[5]), .ZN(y[92]) );
  OR2_X1 U9bar ( .A1(bbar[12]), .A2(abar[5]), .ZN(ybar[92]);
  AND2_X1 U10 ( .A1(b[11]), .A2(a[5]), .ZN(y[91]) );
  OR2_X1 U10bar ( .A1(bbar[11]), .A2(abar[5]), .ZN(ybar[91]);
  AND2_X1 U11 ( .A1(b[10]), .A2(a[5]), .ZN(y[90]) );
  OR2_X1 U11bar ( .A1(bbar[10]), .A2(abar[5]), .ZN(ybar[90]);
  AND2_X1 U12 ( .A1(b[8]), .A2(a[0]), .ZN(y[8]) );
  OR2_X1 U12bar ( .A1(bbar[8]), .A2(abar[0]), .ZN(ybar[8]);
  AND2_X1 U13 ( .A1(a[5]), .A2(b[9]), .ZN(y[89]) );
  OR2_X1 U13bar ( .A1(abar[5]), .A2(bbar[9]), .ZN(ybar[89]);
  AND2_X1 U14 ( .A1(b[8]), .A2(a[5]), .ZN(y[88]) );
  OR2_X1 U14bar ( .A1(bbar[8]), .A2(abar[5]), .ZN(ybar[88]);
  AND2_X1 U15 ( .A1(b[7]), .A2(a[5]), .ZN(y[87]) );
  OR2_X1 U15bar ( .A1(bbar[7]), .A2(abar[5]), .ZN(ybar[87]);
  AND2_X1 U16 ( .A1(b[6]), .A2(a[5]), .ZN(y[86]) );
  OR2_X1 U16bar ( .A1(bbar[6]), .A2(abar[5]), .ZN(ybar[86]);
  AND2_X1 U17 ( .A1(b[5]), .A2(a[5]), .ZN(y[85]) );
  OR2_X1 U17bar ( .A1(bbar[5]), .A2(abar[5]), .ZN(ybar[85]);
  AND2_X1 U18 ( .A1(b[4]), .A2(a[5]), .ZN(y[84]) );
  OR2_X1 U18bar ( .A1(bbar[4]), .A2(abar[5]), .ZN(ybar[84]);
  AND2_X1 U19 ( .A1(a[5]), .A2(b[3]), .ZN(y[83]) );
  OR2_X1 U19bar ( .A1(abar[5]), .A2(bbar[3]), .ZN(ybar[83]);
  AND2_X1 U20 ( .A1(a[5]), .A2(b[2]), .ZN(y[82]) );
  OR2_X1 U20bar ( .A1(abar[5]), .A2(bbar[2]), .ZN(ybar[82]);
  AND2_X1 U21 ( .A1(a[5]), .A2(b[1]), .ZN(y[81]) );
  OR2_X1 U21bar ( .A1(abar[5]), .A2(bbar[1]), .ZN(ybar[81]);
  AND2_X1 U22 ( .A1(a[5]), .A2(b[0]), .ZN(y[80]) );
  OR2_X1 U22bar ( .A1(abar[5]), .A2(bbar[0]), .ZN(ybar[80]);
  AND2_X1 U23 ( .A1(b[7]), .A2(a[0]), .ZN(y[7]) );
  OR2_X1 U23bar ( .A1(bbar[7]), .A2(abar[0]), .ZN(ybar[7]);
  AND2_X1 U24 ( .A1(a[4]), .A2(b[15]), .ZN(y[79]) );
  OR2_X1 U24bar ( .A1(abar[4]), .A2(bbar[15]), .ZN(ybar[79]);
  AND2_X1 U25 ( .A1(a[4]), .A2(b[14]), .ZN(y[78]) );
  OR2_X1 U25bar ( .A1(abar[4]), .A2(bbar[14]), .ZN(ybar[78]);
  AND2_X1 U26 ( .A1(a[4]), .A2(b[13]), .ZN(y[77]) );
  OR2_X1 U26bar ( .A1(abar[4]), .A2(bbar[13]), .ZN(ybar[77]);
  AND2_X1 U27 ( .A1(a[4]), .A2(b[12]), .ZN(y[76]) );
  OR2_X1 U27bar ( .A1(abar[4]), .A2(bbar[12]), .ZN(ybar[76]);
  AND2_X1 U28 ( .A1(a[4]), .A2(b[11]), .ZN(y[75]) );
  OR2_X1 U28bar ( .A1(abar[4]), .A2(bbar[11]), .ZN(ybar[75]);
  AND2_X1 U29 ( .A1(a[4]), .A2(b[10]), .ZN(y[74]) );
  OR2_X1 U29bar ( .A1(abar[4]), .A2(bbar[10]), .ZN(ybar[74]);
  AND2_X1 U30 ( .A1(a[4]), .A2(b[9]), .ZN(y[73]) );
  OR2_X1 U30bar ( .A1(abar[4]), .A2(bbar[9]), .ZN(ybar[73]);
  AND2_X1 U31 ( .A1(a[4]), .A2(b[8]), .ZN(y[72]) );
  OR2_X1 U31bar ( .A1(abar[4]), .A2(bbar[8]), .ZN(ybar[72]);
  AND2_X1 U32 ( .A1(a[4]), .A2(b[7]), .ZN(y[71]) );
  OR2_X1 U32bar ( .A1(abar[4]), .A2(bbar[7]), .ZN(ybar[71]);
  AND2_X1 U33 ( .A1(a[4]), .A2(b[6]), .ZN(y[70]) );
  OR2_X1 U33bar ( .A1(abar[4]), .A2(bbar[6]), .ZN(ybar[70]);
  AND2_X1 U34 ( .A1(b[6]), .A2(a[0]), .ZN(y[6]) );
  OR2_X1 U34bar ( .A1(bbar[6]), .A2(abar[0]), .ZN(ybar[6]);
  AND2_X1 U35 ( .A1(a[4]), .A2(b[5]), .ZN(y[69]) );
  OR2_X1 U35bar ( .A1(abar[4]), .A2(bbar[5]), .ZN(ybar[69]);
  AND2_X1 U36 ( .A1(a[4]), .A2(b[4]), .ZN(y[68]) );
  OR2_X1 U36bar ( .A1(abar[4]), .A2(bbar[4]), .ZN(ybar[68]);
  AND2_X1 U37 ( .A1(a[4]), .A2(b[3]), .ZN(y[67]) );
  OR2_X1 U37bar ( .A1(abar[4]), .A2(bbar[3]), .ZN(ybar[67]);
  AND2_X1 U38 ( .A1(a[4]), .A2(b[2]), .ZN(y[66]) );
  OR2_X1 U38bar ( .A1(abar[4]), .A2(bbar[2]), .ZN(ybar[66]);
  AND2_X1 U39 ( .A1(a[4]), .A2(b[1]), .ZN(y[65]) );
  OR2_X1 U39bar ( .A1(abar[4]), .A2(bbar[1]), .ZN(ybar[65]);
  AND2_X1 U40 ( .A1(a[4]), .A2(b[0]), .ZN(y[64]) );
  OR2_X1 U40bar ( .A1(abar[4]), .A2(bbar[0]), .ZN(ybar[64]);
  AND2_X1 U41 ( .A1(a[3]), .A2(b[15]), .ZN(y[63]) );
  OR2_X1 U41bar ( .A1(abar[3]), .A2(bbar[15]), .ZN(ybar[63]);
  AND2_X1 U42 ( .A1(a[3]), .A2(b[14]), .ZN(y[62]) );
  OR2_X1 U42bar ( .A1(abar[3]), .A2(bbar[14]), .ZN(ybar[62]);
  AND2_X1 U43 ( .A1(a[3]), .A2(b[13]), .ZN(y[61]) );
  OR2_X1 U43bar ( .A1(abar[3]), .A2(bbar[13]), .ZN(ybar[61]);
  AND2_X1 U44 ( .A1(a[3]), .A2(b[12]), .ZN(y[60]) );
  OR2_X1 U44bar ( .A1(abar[3]), .A2(bbar[12]), .ZN(ybar[60]);
  AND2_X1 U45 ( .A1(b[5]), .A2(a[0]), .ZN(y[5]) );
  OR2_X1 U45bar ( .A1(bbar[5]), .A2(abar[0]), .ZN(ybar[5]);
  AND2_X1 U46 ( .A1(a[3]), .A2(b[11]), .ZN(y[59]) );
  OR2_X1 U46bar ( .A1(abar[3]), .A2(bbar[11]), .ZN(ybar[59]);
  AND2_X1 U47 ( .A1(a[3]), .A2(b[10]), .ZN(y[58]) );
  OR2_X1 U47bar ( .A1(abar[3]), .A2(bbar[10]), .ZN(ybar[58]);
  AND2_X1 U48 ( .A1(a[3]), .A2(b[9]), .ZN(y[57]) );
  OR2_X1 U48bar ( .A1(abar[3]), .A2(bbar[9]), .ZN(ybar[57]);
  AND2_X1 U49 ( .A1(a[3]), .A2(b[8]), .ZN(y[56]) );
  OR2_X1 U49bar ( .A1(abar[3]), .A2(bbar[8]), .ZN(ybar[56]);
  AND2_X1 U50 ( .A1(a[3]), .A2(b[7]), .ZN(y[55]) );
  OR2_X1 U50bar ( .A1(abar[3]), .A2(bbar[7]), .ZN(ybar[55]);
  AND2_X1 U51 ( .A1(a[3]), .A2(b[6]), .ZN(y[54]) );
  OR2_X1 U51bar ( .A1(abar[3]), .A2(bbar[6]), .ZN(ybar[54]);
  AND2_X1 U52 ( .A1(a[3]), .A2(b[5]), .ZN(y[53]) );
  OR2_X1 U52bar ( .A1(abar[3]), .A2(bbar[5]), .ZN(ybar[53]);
  AND2_X1 U53 ( .A1(a[3]), .A2(b[4]), .ZN(y[52]) );
  OR2_X1 U53bar ( .A1(abar[3]), .A2(bbar[4]), .ZN(ybar[52]);
  AND2_X1 U54 ( .A1(a[3]), .A2(b[3]), .ZN(y[51]) );
  OR2_X1 U54bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[51]);
  AND2_X1 U55 ( .A1(a[3]), .A2(b[2]), .ZN(y[50]) );
  OR2_X1 U55bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[50]);
  AND2_X1 U56 ( .A1(b[4]), .A2(a[0]), .ZN(y[4]) );
  OR2_X1 U56bar ( .A1(bbar[4]), .A2(abar[0]), .ZN(ybar[4]);
  AND2_X1 U57 ( .A1(a[3]), .A2(b[1]), .ZN(y[49]) );
  OR2_X1 U57bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[49]);
  AND2_X1 U58 ( .A1(a[3]), .A2(b[0]), .ZN(y[48]) );
  OR2_X1 U58bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[48]);
  AND2_X1 U59 ( .A1(a[2]), .A2(b[15]), .ZN(y[47]) );
  OR2_X1 U59bar ( .A1(abar[2]), .A2(bbar[15]), .ZN(ybar[47]);
  AND2_X1 U60 ( .A1(a[2]), .A2(b[14]), .ZN(y[46]) );
  OR2_X1 U60bar ( .A1(abar[2]), .A2(bbar[14]), .ZN(ybar[46]);
  AND2_X1 U61 ( .A1(a[2]), .A2(b[13]), .ZN(y[45]) );
  OR2_X1 U61bar ( .A1(abar[2]), .A2(bbar[13]), .ZN(ybar[45]);
  AND2_X1 U62 ( .A1(a[2]), .A2(b[12]), .ZN(y[44]) );
  OR2_X1 U62bar ( .A1(abar[2]), .A2(bbar[12]), .ZN(ybar[44]);
  AND2_X1 U63 ( .A1(a[2]), .A2(b[11]), .ZN(y[43]) );
  OR2_X1 U63bar ( .A1(abar[2]), .A2(bbar[11]), .ZN(ybar[43]);
  AND2_X1 U64 ( .A1(a[2]), .A2(b[10]), .ZN(y[42]) );
  OR2_X1 U64bar ( .A1(abar[2]), .A2(bbar[10]), .ZN(ybar[42]);
  AND2_X1 U65 ( .A1(a[2]), .A2(b[9]), .ZN(y[41]) );
  OR2_X1 U65bar ( .A1(abar[2]), .A2(bbar[9]), .ZN(ybar[41]);
  AND2_X1 U66 ( .A1(a[2]), .A2(b[8]), .ZN(y[40]) );
  OR2_X1 U66bar ( .A1(abar[2]), .A2(bbar[8]), .ZN(ybar[40]);
  AND2_X1 U67 ( .A1(b[3]), .A2(a[0]), .ZN(y[3]) );
  OR2_X1 U67bar ( .A1(bbar[3]), .A2(abar[0]), .ZN(ybar[3]);
  AND2_X1 U68 ( .A1(a[2]), .A2(b[7]), .ZN(y[39]) );
  OR2_X1 U68bar ( .A1(abar[2]), .A2(bbar[7]), .ZN(ybar[39]);
  AND2_X1 U69 ( .A1(a[2]), .A2(b[6]), .ZN(y[38]) );
  OR2_X1 U69bar ( .A1(abar[2]), .A2(bbar[6]), .ZN(ybar[38]);
  AND2_X1 U70 ( .A1(a[2]), .A2(b[5]), .ZN(y[37]) );
  OR2_X1 U70bar ( .A1(abar[2]), .A2(bbar[5]), .ZN(ybar[37]);
  AND2_X1 U71 ( .A1(a[2]), .A2(b[4]), .ZN(y[36]) );
  OR2_X1 U71bar ( .A1(abar[2]), .A2(bbar[4]), .ZN(ybar[36]);
  AND2_X1 U72 ( .A1(a[2]), .A2(b[3]), .ZN(y[35]) );
  OR2_X1 U72bar ( .A1(abar[2]), .A2(bbar[3]), .ZN(ybar[35]);
  AND2_X1 U73 ( .A1(a[2]), .A2(b[2]), .ZN(y[34]) );
  OR2_X1 U73bar ( .A1(abar[2]), .A2(bbar[2]), .ZN(ybar[34]);
  AND2_X1 U74 ( .A1(a[2]), .A2(b[1]), .ZN(y[33]) );
  OR2_X1 U74bar ( .A1(abar[2]), .A2(bbar[1]), .ZN(ybar[33]);
  AND2_X1 U75 ( .A1(a[2]), .A2(b[0]), .ZN(y[32]) );
  OR2_X1 U75bar ( .A1(abar[2]), .A2(bbar[0]), .ZN(ybar[32]);
  AND2_X1 U76 ( .A1(a[1]), .A2(b[15]), .ZN(y[31]) );
  OR2_X1 U76bar ( .A1(abar[1]), .A2(bbar[15]), .ZN(ybar[31]);
  AND2_X1 U77 ( .A1(a[1]), .A2(b[14]), .ZN(y[30]) );
  OR2_X1 U77bar ( .A1(abar[1]), .A2(bbar[14]), .ZN(ybar[30]);
  AND2_X1 U78 ( .A1(b[2]), .A2(a[0]), .ZN(y[2]) );
  OR2_X1 U78bar ( .A1(bbar[2]), .A2(abar[0]), .ZN(ybar[2]);
  AND2_X1 U79 ( .A1(a[1]), .A2(b[13]), .ZN(y[29]) );
  OR2_X1 U79bar ( .A1(abar[1]), .A2(bbar[13]), .ZN(ybar[29]);
  AND2_X1 U80 ( .A1(a[1]), .A2(b[12]), .ZN(y[28]) );
  OR2_X1 U80bar ( .A1(abar[1]), .A2(bbar[12]), .ZN(ybar[28]);
  AND2_X1 U81 ( .A1(a[1]), .A2(b[11]), .ZN(y[27]) );
  OR2_X1 U81bar ( .A1(abar[1]), .A2(bbar[11]), .ZN(ybar[27]);
  AND2_X1 U82 ( .A1(a[1]), .A2(b[10]), .ZN(y[26]) );
  OR2_X1 U82bar ( .A1(abar[1]), .A2(bbar[10]), .ZN(ybar[26]);
  AND2_X1 U83 ( .A1(a[1]), .A2(b[9]), .ZN(y[25]) );
  OR2_X1 U83bar ( .A1(abar[1]), .A2(bbar[9]), .ZN(ybar[25]);
  AND2_X1 U84 ( .A1(a[15]), .A2(b[15]), .ZN(y[255]) );
  OR2_X1 U84bar ( .A1(abar[15]), .A2(bbar[15]), .ZN(ybar[255]);
  AND2_X1 U85 ( .A1(a[15]), .A2(b[14]), .ZN(y[254]) );
  OR2_X1 U85bar ( .A1(abar[15]), .A2(bbar[14]), .ZN(ybar[254]);
  AND2_X1 U86 ( .A1(a[15]), .A2(b[13]), .ZN(y[253]) );
  OR2_X1 U86bar ( .A1(abar[15]), .A2(bbar[13]), .ZN(ybar[253]);
  AND2_X1 U87 ( .A1(a[15]), .A2(b[12]), .ZN(y[252]) );
  OR2_X1 U87bar ( .A1(abar[15]), .A2(bbar[12]), .ZN(ybar[252]);
  AND2_X1 U88 ( .A1(a[15]), .A2(b[11]), .ZN(y[251]) );
  OR2_X1 U88bar ( .A1(abar[15]), .A2(bbar[11]), .ZN(ybar[251]);
  AND2_X1 U89 ( .A1(a[15]), .A2(b[10]), .ZN(y[250]) );
  OR2_X1 U89bar ( .A1(abar[15]), .A2(bbar[10]), .ZN(ybar[250]);
  AND2_X1 U90 ( .A1(a[1]), .A2(b[8]), .ZN(y[24]) );
  OR2_X1 U90bar ( .A1(abar[1]), .A2(bbar[8]), .ZN(ybar[24]);
  AND2_X1 U91 ( .A1(a[15]), .A2(b[9]), .ZN(y[249]) );
  OR2_X1 U91bar ( .A1(abar[15]), .A2(bbar[9]), .ZN(ybar[249]);
  AND2_X1 U92 ( .A1(a[15]), .A2(b[8]), .ZN(y[248]) );
  OR2_X1 U92bar ( .A1(abar[15]), .A2(bbar[8]), .ZN(ybar[248]);
  AND2_X1 U93 ( .A1(a[15]), .A2(b[7]), .ZN(y[247]) );
  OR2_X1 U93bar ( .A1(abar[15]), .A2(bbar[7]), .ZN(ybar[247]);
  AND2_X1 U94 ( .A1(a[15]), .A2(b[6]), .ZN(y[246]) );
  OR2_X1 U94bar ( .A1(abar[15]), .A2(bbar[6]), .ZN(ybar[246]);
  AND2_X1 U95 ( .A1(a[15]), .A2(b[5]), .ZN(y[245]) );
  OR2_X1 U95bar ( .A1(abar[15]), .A2(bbar[5]), .ZN(ybar[245]);
  AND2_X1 U96 ( .A1(a[15]), .A2(b[4]), .ZN(y[244]) );
  OR2_X1 U96bar ( .A1(abar[15]), .A2(bbar[4]), .ZN(ybar[244]);
  AND2_X1 U97 ( .A1(a[15]), .A2(b[3]), .ZN(y[243]) );
  OR2_X1 U97bar ( .A1(abar[15]), .A2(bbar[3]), .ZN(ybar[243]);
  AND2_X1 U98 ( .A1(a[15]), .A2(b[2]), .ZN(y[242]) );
  OR2_X1 U98bar ( .A1(abar[15]), .A2(bbar[2]), .ZN(ybar[242]);
  AND2_X1 U99 ( .A1(a[15]), .A2(b[1]), .ZN(y[241]) );
  OR2_X1 U99bar ( .A1(abar[15]), .A2(bbar[1]), .ZN(ybar[241]);
  AND2_X1 U100 ( .A1(a[15]), .A2(b[0]), .ZN(y[240]) );
  OR2_X1 U100bar ( .A1(abar[15]), .A2(bbar[0]), .ZN(ybar[240]);
  AND2_X1 U101 ( .A1(a[1]), .A2(b[7]), .ZN(y[23]) );
  OR2_X1 U101bar ( .A1(abar[1]), .A2(bbar[7]), .ZN(ybar[23]);
  AND2_X1 U102 ( .A1(a[14]), .A2(b[15]), .ZN(y[239]) );
  OR2_X1 U102bar ( .A1(abar[14]), .A2(bbar[15]), .ZN(ybar[239]);
  AND2_X1 U103 ( .A1(a[14]), .A2(b[14]), .ZN(y[238]) );
  OR2_X1 U103bar ( .A1(abar[14]), .A2(bbar[14]), .ZN(ybar[238]);
  AND2_X1 U104 ( .A1(a[14]), .A2(b[13]), .ZN(y[237]) );
  OR2_X1 U104bar ( .A1(abar[14]), .A2(bbar[13]), .ZN(ybar[237]);
  AND2_X1 U105 ( .A1(a[14]), .A2(b[12]), .ZN(y[236]) );
  OR2_X1 U105bar ( .A1(abar[14]), .A2(bbar[12]), .ZN(ybar[236]);
  AND2_X1 U106 ( .A1(a[14]), .A2(b[11]), .ZN(y[235]) );
  OR2_X1 U106bar ( .A1(abar[14]), .A2(bbar[11]), .ZN(ybar[235]);
  AND2_X1 U107 ( .A1(a[14]), .A2(b[10]), .ZN(y[234]) );
  OR2_X1 U107bar ( .A1(abar[14]), .A2(bbar[10]), .ZN(ybar[234]);
  AND2_X1 U108 ( .A1(a[14]), .A2(b[9]), .ZN(y[233]) );
  OR2_X1 U108bar ( .A1(abar[14]), .A2(bbar[9]), .ZN(ybar[233]);
  AND2_X1 U109 ( .A1(a[14]), .A2(b[8]), .ZN(y[232]) );
  OR2_X1 U109bar ( .A1(abar[14]), .A2(bbar[8]), .ZN(ybar[232]);
  AND2_X1 U110 ( .A1(a[14]), .A2(b[7]), .ZN(y[231]) );
  OR2_X1 U110bar ( .A1(abar[14]), .A2(bbar[7]), .ZN(ybar[231]);
  AND2_X1 U111 ( .A1(a[14]), .A2(b[6]), .ZN(y[230]) );
  OR2_X1 U111bar ( .A1(abar[14]), .A2(bbar[6]), .ZN(ybar[230]);
  AND2_X1 U112 ( .A1(a[1]), .A2(b[6]), .ZN(y[22]) );
  OR2_X1 U112bar ( .A1(abar[1]), .A2(bbar[6]), .ZN(ybar[22]);
  AND2_X1 U113 ( .A1(a[14]), .A2(b[5]), .ZN(y[229]) );
  OR2_X1 U113bar ( .A1(abar[14]), .A2(bbar[5]), .ZN(ybar[229]);
  AND2_X1 U114 ( .A1(a[14]), .A2(b[4]), .ZN(y[228]) );
  OR2_X1 U114bar ( .A1(abar[14]), .A2(bbar[4]), .ZN(ybar[228]);
  AND2_X1 U115 ( .A1(a[14]), .A2(b[3]), .ZN(y[227]) );
  OR2_X1 U115bar ( .A1(abar[14]), .A2(bbar[3]), .ZN(ybar[227]);
  AND2_X1 U116 ( .A1(a[14]), .A2(b[2]), .ZN(y[226]) );
  OR2_X1 U116bar ( .A1(abar[14]), .A2(bbar[2]), .ZN(ybar[226]);
  AND2_X1 U117 ( .A1(a[14]), .A2(b[1]), .ZN(y[225]) );
  OR2_X1 U117bar ( .A1(abar[14]), .A2(bbar[1]), .ZN(ybar[225]);
  AND2_X1 U118 ( .A1(a[14]), .A2(b[0]), .ZN(y[224]) );
  OR2_X1 U118bar ( .A1(abar[14]), .A2(bbar[0]), .ZN(ybar[224]);
  AND2_X1 U119 ( .A1(a[13]), .A2(b[15]), .ZN(y[223]) );
  OR2_X1 U119bar ( .A1(abar[13]), .A2(bbar[15]), .ZN(ybar[223]);
  AND2_X1 U120 ( .A1(a[13]), .A2(b[14]), .ZN(y[222]) );
  OR2_X1 U120bar ( .A1(abar[13]), .A2(bbar[14]), .ZN(ybar[222]);
  AND2_X1 U121 ( .A1(a[13]), .A2(b[13]), .ZN(y[221]) );
  OR2_X1 U121bar ( .A1(abar[13]), .A2(bbar[13]), .ZN(ybar[221]);
  AND2_X1 U122 ( .A1(a[13]), .A2(b[12]), .ZN(y[220]) );
  OR2_X1 U122bar ( .A1(abar[13]), .A2(bbar[12]), .ZN(ybar[220]);
  AND2_X1 U123 ( .A1(a[1]), .A2(b[5]), .ZN(y[21]) );
  OR2_X1 U123bar ( .A1(abar[1]), .A2(bbar[5]), .ZN(ybar[21]);
  AND2_X1 U124 ( .A1(a[13]), .A2(b[11]), .ZN(y[219]) );
  OR2_X1 U124bar ( .A1(abar[13]), .A2(bbar[11]), .ZN(ybar[219]);
  AND2_X1 U125 ( .A1(a[13]), .A2(b[10]), .ZN(y[218]) );
  OR2_X1 U125bar ( .A1(abar[13]), .A2(bbar[10]), .ZN(ybar[218]);
  AND2_X1 U126 ( .A1(a[13]), .A2(b[9]), .ZN(y[217]) );
  OR2_X1 U126bar ( .A1(abar[13]), .A2(bbar[9]), .ZN(ybar[217]);
  AND2_X1 U127 ( .A1(a[13]), .A2(b[8]), .ZN(y[216]) );
  OR2_X1 U127bar ( .A1(abar[13]), .A2(bbar[8]), .ZN(ybar[216]);
  AND2_X1 U128 ( .A1(a[13]), .A2(b[7]), .ZN(y[215]) );
  OR2_X1 U128bar ( .A1(abar[13]), .A2(bbar[7]), .ZN(ybar[215]);
  AND2_X1 U129 ( .A1(a[13]), .A2(b[6]), .ZN(y[214]) );
  OR2_X1 U129bar ( .A1(abar[13]), .A2(bbar[6]), .ZN(ybar[214]);
  AND2_X1 U130 ( .A1(a[13]), .A2(b[5]), .ZN(y[213]) );
  OR2_X1 U130bar ( .A1(abar[13]), .A2(bbar[5]), .ZN(ybar[213]);
  AND2_X1 U131 ( .A1(a[13]), .A2(b[4]), .ZN(y[212]) );
  OR2_X1 U131bar ( .A1(abar[13]), .A2(bbar[4]), .ZN(ybar[212]);
  AND2_X1 U132 ( .A1(a[13]), .A2(b[3]), .ZN(y[211]) );
  OR2_X1 U132bar ( .A1(abar[13]), .A2(bbar[3]), .ZN(ybar[211]);
  AND2_X1 U133 ( .A1(a[13]), .A2(b[2]), .ZN(y[210]) );
  OR2_X1 U133bar ( .A1(abar[13]), .A2(bbar[2]), .ZN(ybar[210]);
  AND2_X1 U134 ( .A1(a[1]), .A2(b[4]), .ZN(y[20]) );
  OR2_X1 U134bar ( .A1(abar[1]), .A2(bbar[4]), .ZN(ybar[20]);
  AND2_X1 U135 ( .A1(a[13]), .A2(b[1]), .ZN(y[209]) );
  OR2_X1 U135bar ( .A1(abar[13]), .A2(bbar[1]), .ZN(ybar[209]);
  AND2_X1 U136 ( .A1(a[13]), .A2(b[0]), .ZN(y[208]) );
  OR2_X1 U136bar ( .A1(abar[13]), .A2(bbar[0]), .ZN(ybar[208]);
  AND2_X1 U137 ( .A1(a[12]), .A2(b[15]), .ZN(y[207]) );
  OR2_X1 U137bar ( .A1(abar[12]), .A2(bbar[15]), .ZN(ybar[207]);
  AND2_X1 U138 ( .A1(a[12]), .A2(b[14]), .ZN(y[206]) );
  OR2_X1 U138bar ( .A1(abar[12]), .A2(bbar[14]), .ZN(ybar[206]);
  AND2_X1 U139 ( .A1(a[12]), .A2(b[13]), .ZN(y[205]) );
  OR2_X1 U139bar ( .A1(abar[12]), .A2(bbar[13]), .ZN(ybar[205]);
  AND2_X1 U140 ( .A1(a[12]), .A2(b[12]), .ZN(y[204]) );
  OR2_X1 U140bar ( .A1(abar[12]), .A2(bbar[12]), .ZN(ybar[204]);
  AND2_X1 U141 ( .A1(a[12]), .A2(b[11]), .ZN(y[203]) );
  OR2_X1 U141bar ( .A1(abar[12]), .A2(bbar[11]), .ZN(ybar[203]);
  AND2_X1 U142 ( .A1(a[12]), .A2(b[10]), .ZN(y[202]) );
  OR2_X1 U142bar ( .A1(abar[12]), .A2(bbar[10]), .ZN(ybar[202]);
  AND2_X1 U143 ( .A1(a[12]), .A2(b[9]), .ZN(y[201]) );
  OR2_X1 U143bar ( .A1(abar[12]), .A2(bbar[9]), .ZN(ybar[201]);
  AND2_X1 U144 ( .A1(a[12]), .A2(b[8]), .ZN(y[200]) );
  OR2_X1 U144bar ( .A1(abar[12]), .A2(bbar[8]), .ZN(ybar[200]);
  AND2_X1 U145 ( .A1(b[1]), .A2(a[0]), .ZN(y[1]) );
  OR2_X1 U145bar ( .A1(bbar[1]), .A2(abar[0]), .ZN(ybar[1]);
  AND2_X1 U146 ( .A1(a[1]), .A2(b[3]), .ZN(y[19]) );
  OR2_X1 U146bar ( .A1(abar[1]), .A2(bbar[3]), .ZN(ybar[19]);
  AND2_X1 U147 ( .A1(a[12]), .A2(b[7]), .ZN(y[199]) );
  OR2_X1 U147bar ( .A1(abar[12]), .A2(bbar[7]), .ZN(ybar[199]);
  AND2_X1 U148 ( .A1(a[12]), .A2(b[6]), .ZN(y[198]) );
  OR2_X1 U148bar ( .A1(abar[12]), .A2(bbar[6]), .ZN(ybar[198]);
  AND2_X1 U149 ( .A1(a[12]), .A2(b[5]), .ZN(y[197]) );
  OR2_X1 U149bar ( .A1(abar[12]), .A2(bbar[5]), .ZN(ybar[197]);
  AND2_X1 U150 ( .A1(a[12]), .A2(b[4]), .ZN(y[196]) );
  OR2_X1 U150bar ( .A1(abar[12]), .A2(bbar[4]), .ZN(ybar[196]);
  AND2_X1 U151 ( .A1(a[12]), .A2(b[3]), .ZN(y[195]) );
  OR2_X1 U151bar ( .A1(abar[12]), .A2(bbar[3]), .ZN(ybar[195]);
  AND2_X1 U152 ( .A1(a[12]), .A2(b[2]), .ZN(y[194]) );
  OR2_X1 U152bar ( .A1(abar[12]), .A2(bbar[2]), .ZN(ybar[194]);
  AND2_X1 U153 ( .A1(a[12]), .A2(b[1]), .ZN(y[193]) );
  OR2_X1 U153bar ( .A1(abar[12]), .A2(bbar[1]), .ZN(ybar[193]);
  AND2_X1 U154 ( .A1(a[12]), .A2(b[0]), .ZN(y[192]) );
  OR2_X1 U154bar ( .A1(abar[12]), .A2(bbar[0]), .ZN(ybar[192]);
  AND2_X1 U155 ( .A1(a[11]), .A2(b[15]), .ZN(y[191]) );
  OR2_X1 U155bar ( .A1(abar[11]), .A2(bbar[15]), .ZN(ybar[191]);
  AND2_X1 U156 ( .A1(a[11]), .A2(b[14]), .ZN(y[190]) );
  OR2_X1 U156bar ( .A1(abar[11]), .A2(bbar[14]), .ZN(ybar[190]);
  AND2_X1 U157 ( .A1(a[1]), .A2(b[2]), .ZN(y[18]) );
  OR2_X1 U157bar ( .A1(abar[1]), .A2(bbar[2]), .ZN(ybar[18]);
  AND2_X1 U158 ( .A1(a[11]), .A2(b[13]), .ZN(y[189]) );
  OR2_X1 U158bar ( .A1(abar[11]), .A2(bbar[13]), .ZN(ybar[189]);
  AND2_X1 U159 ( .A1(a[11]), .A2(b[12]), .ZN(y[188]) );
  OR2_X1 U159bar ( .A1(abar[11]), .A2(bbar[12]), .ZN(ybar[188]);
  AND2_X1 U160 ( .A1(a[11]), .A2(b[11]), .ZN(y[187]) );
  OR2_X1 U160bar ( .A1(abar[11]), .A2(bbar[11]), .ZN(ybar[187]);
  AND2_X1 U161 ( .A1(a[11]), .A2(b[10]), .ZN(y[186]) );
  OR2_X1 U161bar ( .A1(abar[11]), .A2(bbar[10]), .ZN(ybar[186]);
  AND2_X1 U162 ( .A1(a[11]), .A2(b[9]), .ZN(y[185]) );
  OR2_X1 U162bar ( .A1(abar[11]), .A2(bbar[9]), .ZN(ybar[185]);
  AND2_X1 U163 ( .A1(a[11]), .A2(b[8]), .ZN(y[184]) );
  OR2_X1 U163bar ( .A1(abar[11]), .A2(bbar[8]), .ZN(ybar[184]);
  AND2_X1 U164 ( .A1(a[11]), .A2(b[7]), .ZN(y[183]) );
  OR2_X1 U164bar ( .A1(abar[11]), .A2(bbar[7]), .ZN(ybar[183]);
  AND2_X1 U165 ( .A1(a[11]), .A2(b[6]), .ZN(y[182]) );
  OR2_X1 U165bar ( .A1(abar[11]), .A2(bbar[6]), .ZN(ybar[182]);
  AND2_X1 U166 ( .A1(a[11]), .A2(b[5]), .ZN(y[181]) );
  OR2_X1 U166bar ( .A1(abar[11]), .A2(bbar[5]), .ZN(ybar[181]);
  AND2_X1 U167 ( .A1(a[11]), .A2(b[4]), .ZN(y[180]) );
  OR2_X1 U167bar ( .A1(abar[11]), .A2(bbar[4]), .ZN(ybar[180]);
  AND2_X1 U168 ( .A1(a[1]), .A2(b[1]), .ZN(y[17]) );
  OR2_X1 U168bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[17]);
  AND2_X1 U169 ( .A1(a[11]), .A2(b[3]), .ZN(y[179]) );
  OR2_X1 U169bar ( .A1(abar[11]), .A2(bbar[3]), .ZN(ybar[179]);
  AND2_X1 U170 ( .A1(a[11]), .A2(b[2]), .ZN(y[178]) );
  OR2_X1 U170bar ( .A1(abar[11]), .A2(bbar[2]), .ZN(ybar[178]);
  AND2_X1 U171 ( .A1(a[11]), .A2(b[1]), .ZN(y[177]) );
  OR2_X1 U171bar ( .A1(abar[11]), .A2(bbar[1]), .ZN(ybar[177]);
  AND2_X1 U172 ( .A1(a[11]), .A2(b[0]), .ZN(y[176]) );
  OR2_X1 U172bar ( .A1(abar[11]), .A2(bbar[0]), .ZN(ybar[176]);
  AND2_X1 U173 ( .A1(a[10]), .A2(b[15]), .ZN(y[175]) );
  OR2_X1 U173bar ( .A1(abar[10]), .A2(bbar[15]), .ZN(ybar[175]);
  AND2_X1 U174 ( .A1(a[10]), .A2(b[14]), .ZN(y[174]) );
  OR2_X1 U174bar ( .A1(abar[10]), .A2(bbar[14]), .ZN(ybar[174]);
  AND2_X1 U175 ( .A1(a[10]), .A2(b[13]), .ZN(y[173]) );
  OR2_X1 U175bar ( .A1(abar[10]), .A2(bbar[13]), .ZN(ybar[173]);
  AND2_X1 U176 ( .A1(a[10]), .A2(b[12]), .ZN(y[172]) );
  OR2_X1 U176bar ( .A1(abar[10]), .A2(bbar[12]), .ZN(ybar[172]);
  AND2_X1 U177 ( .A1(a[10]), .A2(b[11]), .ZN(y[171]) );
  OR2_X1 U177bar ( .A1(abar[10]), .A2(bbar[11]), .ZN(ybar[171]);
  AND2_X1 U178 ( .A1(a[10]), .A2(b[10]), .ZN(y[170]) );
  OR2_X1 U178bar ( .A1(abar[10]), .A2(bbar[10]), .ZN(ybar[170]);
  AND2_X1 U179 ( .A1(a[1]), .A2(b[0]), .ZN(y[16]) );
  OR2_X1 U179bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[16]);
  AND2_X1 U180 ( .A1(a[10]), .A2(b[9]), .ZN(y[169]) );
  OR2_X1 U180bar ( .A1(abar[10]), .A2(bbar[9]), .ZN(ybar[169]);
  AND2_X1 U181 ( .A1(a[10]), .A2(b[8]), .ZN(y[168]) );
  OR2_X1 U181bar ( .A1(abar[10]), .A2(bbar[8]), .ZN(ybar[168]);
  AND2_X1 U182 ( .A1(a[10]), .A2(b[7]), .ZN(y[167]) );
  OR2_X1 U182bar ( .A1(abar[10]), .A2(bbar[7]), .ZN(ybar[167]);
  AND2_X1 U183 ( .A1(a[10]), .A2(b[6]), .ZN(y[166]) );
  OR2_X1 U183bar ( .A1(abar[10]), .A2(bbar[6]), .ZN(ybar[166]);
  AND2_X1 U184 ( .A1(a[10]), .A2(b[5]), .ZN(y[165]) );
  OR2_X1 U184bar ( .A1(abar[10]), .A2(bbar[5]), .ZN(ybar[165]);
  AND2_X1 U185 ( .A1(a[10]), .A2(b[4]), .ZN(y[164]) );
  OR2_X1 U185bar ( .A1(abar[10]), .A2(bbar[4]), .ZN(ybar[164]);
  AND2_X1 U186 ( .A1(a[10]), .A2(b[3]), .ZN(y[163]) );
  OR2_X1 U186bar ( .A1(abar[10]), .A2(bbar[3]), .ZN(ybar[163]);
  AND2_X1 U187 ( .A1(a[10]), .A2(b[2]), .ZN(y[162]) );
  OR2_X1 U187bar ( .A1(abar[10]), .A2(bbar[2]), .ZN(ybar[162]);
  AND2_X1 U188 ( .A1(a[10]), .A2(b[1]), .ZN(y[161]) );
  OR2_X1 U188bar ( .A1(abar[10]), .A2(bbar[1]), .ZN(ybar[161]);
  AND2_X1 U189 ( .A1(a[10]), .A2(b[0]), .ZN(y[160]) );
  OR2_X1 U189bar ( .A1(abar[10]), .A2(bbar[0]), .ZN(ybar[160]);
  AND2_X1 U190 ( .A1(b[15]), .A2(a[0]), .ZN(y[15]) );
  OR2_X1 U190bar ( .A1(bbar[15]), .A2(abar[0]), .ZN(ybar[15]);
  AND2_X1 U191 ( .A1(a[9]), .A2(b[15]), .ZN(y[159]) );
  OR2_X1 U191bar ( .A1(abar[9]), .A2(bbar[15]), .ZN(ybar[159]);
  AND2_X1 U192 ( .A1(a[9]), .A2(b[14]), .ZN(y[158]) );
  OR2_X1 U192bar ( .A1(abar[9]), .A2(bbar[14]), .ZN(ybar[158]);
  AND2_X1 U193 ( .A1(a[9]), .A2(b[13]), .ZN(y[157]) );
  OR2_X1 U193bar ( .A1(abar[9]), .A2(bbar[13]), .ZN(ybar[157]);
  AND2_X1 U194 ( .A1(a[9]), .A2(b[12]), .ZN(y[156]) );
  OR2_X1 U194bar ( .A1(abar[9]), .A2(bbar[12]), .ZN(ybar[156]);
  AND2_X1 U195 ( .A1(a[9]), .A2(b[11]), .ZN(y[155]) );
  OR2_X1 U195bar ( .A1(abar[9]), .A2(bbar[11]), .ZN(ybar[155]);
  AND2_X1 U196 ( .A1(a[9]), .A2(b[10]), .ZN(y[154]) );
  OR2_X1 U196bar ( .A1(abar[9]), .A2(bbar[10]), .ZN(ybar[154]);
  AND2_X1 U197 ( .A1(a[9]), .A2(b[9]), .ZN(y[153]) );
  OR2_X1 U197bar ( .A1(abar[9]), .A2(bbar[9]), .ZN(ybar[153]);
  AND2_X1 U198 ( .A1(a[9]), .A2(b[8]), .ZN(y[152]) );
  OR2_X1 U198bar ( .A1(abar[9]), .A2(bbar[8]), .ZN(ybar[152]);
  AND2_X1 U199 ( .A1(a[9]), .A2(b[7]), .ZN(y[151]) );
  OR2_X1 U199bar ( .A1(abar[9]), .A2(bbar[7]), .ZN(ybar[151]);
  AND2_X1 U200 ( .A1(a[9]), .A2(b[6]), .ZN(y[150]) );
  OR2_X1 U200bar ( .A1(abar[9]), .A2(bbar[6]), .ZN(ybar[150]);
  AND2_X1 U201 ( .A1(b[14]), .A2(a[0]), .ZN(y[14]) );
  OR2_X1 U201bar ( .A1(bbar[14]), .A2(abar[0]), .ZN(ybar[14]);
  AND2_X1 U202 ( .A1(a[9]), .A2(b[5]), .ZN(y[149]) );
  OR2_X1 U202bar ( .A1(abar[9]), .A2(bbar[5]), .ZN(ybar[149]);
  AND2_X1 U203 ( .A1(a[9]), .A2(b[4]), .ZN(y[148]) );
  OR2_X1 U203bar ( .A1(abar[9]), .A2(bbar[4]), .ZN(ybar[148]);
  AND2_X1 U204 ( .A1(a[9]), .A2(b[3]), .ZN(y[147]) );
  OR2_X1 U204bar ( .A1(abar[9]), .A2(bbar[3]), .ZN(ybar[147]);
  AND2_X1 U205 ( .A1(a[9]), .A2(b[2]), .ZN(y[146]) );
  OR2_X1 U205bar ( .A1(abar[9]), .A2(bbar[2]), .ZN(ybar[146]);
  AND2_X1 U206 ( .A1(a[9]), .A2(b[1]), .ZN(y[145]) );
  OR2_X1 U206bar ( .A1(abar[9]), .A2(bbar[1]), .ZN(ybar[145]);
  AND2_X1 U207 ( .A1(a[9]), .A2(b[0]), .ZN(y[144]) );
  OR2_X1 U207bar ( .A1(abar[9]), .A2(bbar[0]), .ZN(ybar[144]);
  AND2_X1 U208 ( .A1(a[8]), .A2(b[15]), .ZN(y[143]) );
  OR2_X1 U208bar ( .A1(abar[8]), .A2(bbar[15]), .ZN(ybar[143]);
  AND2_X1 U209 ( .A1(a[8]), .A2(b[14]), .ZN(y[142]) );
  OR2_X1 U209bar ( .A1(abar[8]), .A2(bbar[14]), .ZN(ybar[142]);
  AND2_X1 U210 ( .A1(a[8]), .A2(b[13]), .ZN(y[141]) );
  OR2_X1 U210bar ( .A1(abar[8]), .A2(bbar[13]), .ZN(ybar[141]);
  AND2_X1 U211 ( .A1(a[8]), .A2(b[12]), .ZN(y[140]) );
  OR2_X1 U211bar ( .A1(abar[8]), .A2(bbar[12]), .ZN(ybar[140]);
  AND2_X1 U212 ( .A1(b[13]), .A2(a[0]), .ZN(y[13]) );
  OR2_X1 U212bar ( .A1(bbar[13]), .A2(abar[0]), .ZN(ybar[13]);
  AND2_X1 U213 ( .A1(a[8]), .A2(b[11]), .ZN(y[139]) );
  OR2_X1 U213bar ( .A1(abar[8]), .A2(bbar[11]), .ZN(ybar[139]);
  AND2_X1 U214 ( .A1(a[8]), .A2(b[10]), .ZN(y[138]) );
  OR2_X1 U214bar ( .A1(abar[8]), .A2(bbar[10]), .ZN(ybar[138]);
  AND2_X1 U215 ( .A1(a[8]), .A2(b[9]), .ZN(y[137]) );
  OR2_X1 U215bar ( .A1(abar[8]), .A2(bbar[9]), .ZN(ybar[137]);
  AND2_X1 U216 ( .A1(a[8]), .A2(b[8]), .ZN(y[136]) );
  OR2_X1 U216bar ( .A1(abar[8]), .A2(bbar[8]), .ZN(ybar[136]);
  AND2_X1 U217 ( .A1(a[8]), .A2(b[7]), .ZN(y[135]) );
  OR2_X1 U217bar ( .A1(abar[8]), .A2(bbar[7]), .ZN(ybar[135]);
  AND2_X1 U218 ( .A1(a[8]), .A2(b[6]), .ZN(y[134]) );
  OR2_X1 U218bar ( .A1(abar[8]), .A2(bbar[6]), .ZN(ybar[134]);
  AND2_X1 U219 ( .A1(a[8]), .A2(b[5]), .ZN(y[133]) );
  OR2_X1 U219bar ( .A1(abar[8]), .A2(bbar[5]), .ZN(ybar[133]);
  AND2_X1 U220 ( .A1(a[8]), .A2(b[4]), .ZN(y[132]) );
  OR2_X1 U220bar ( .A1(abar[8]), .A2(bbar[4]), .ZN(ybar[132]);
  AND2_X1 U221 ( .A1(a[8]), .A2(b[3]), .ZN(y[131]) );
  OR2_X1 U221bar ( .A1(abar[8]), .A2(bbar[3]), .ZN(ybar[131]);
  AND2_X1 U222 ( .A1(a[8]), .A2(b[2]), .ZN(y[130]) );
  OR2_X1 U222bar ( .A1(abar[8]), .A2(bbar[2]), .ZN(ybar[130]);
  AND2_X1 U223 ( .A1(b[12]), .A2(a[0]), .ZN(y[12]) );
  OR2_X1 U223bar ( .A1(bbar[12]), .A2(abar[0]), .ZN(ybar[12]);
  AND2_X1 U224 ( .A1(a[8]), .A2(b[1]), .ZN(y[129]) );
  OR2_X1 U224bar ( .A1(abar[8]), .A2(bbar[1]), .ZN(ybar[129]);
  AND2_X1 U225 ( .A1(a[8]), .A2(b[0]), .ZN(y[128]) );
  OR2_X1 U225bar ( .A1(abar[8]), .A2(bbar[0]), .ZN(ybar[128]);
  AND2_X1 U226 ( .A1(a[7]), .A2(b[15]), .ZN(y[127]) );
  OR2_X1 U226bar ( .A1(abar[7]), .A2(bbar[15]), .ZN(ybar[127]);
  AND2_X1 U227 ( .A1(a[7]), .A2(b[14]), .ZN(y[126]) );
  OR2_X1 U227bar ( .A1(abar[7]), .A2(bbar[14]), .ZN(ybar[126]);
  AND2_X1 U228 ( .A1(a[7]), .A2(b[13]), .ZN(y[125]) );
  OR2_X1 U228bar ( .A1(abar[7]), .A2(bbar[13]), .ZN(ybar[125]);
  AND2_X1 U229 ( .A1(a[7]), .A2(b[12]), .ZN(y[124]) );
  OR2_X1 U229bar ( .A1(abar[7]), .A2(bbar[12]), .ZN(ybar[124]);
  AND2_X1 U230 ( .A1(a[7]), .A2(b[11]), .ZN(y[123]) );
  OR2_X1 U230bar ( .A1(abar[7]), .A2(bbar[11]), .ZN(ybar[123]);
  AND2_X1 U231 ( .A1(a[7]), .A2(b[10]), .ZN(y[122]) );
  OR2_X1 U231bar ( .A1(abar[7]), .A2(bbar[10]), .ZN(ybar[122]);
  AND2_X1 U232 ( .A1(a[7]), .A2(b[9]), .ZN(y[121]) );
  OR2_X1 U232bar ( .A1(abar[7]), .A2(bbar[9]), .ZN(ybar[121]);
  AND2_X1 U233 ( .A1(a[7]), .A2(b[8]), .ZN(y[120]) );
  OR2_X1 U233bar ( .A1(abar[7]), .A2(bbar[8]), .ZN(ybar[120]);
  AND2_X1 U234 ( .A1(b[11]), .A2(a[0]), .ZN(y[11]) );
  OR2_X1 U234bar ( .A1(bbar[11]), .A2(abar[0]), .ZN(ybar[11]);
  AND2_X1 U235 ( .A1(a[7]), .A2(b[7]), .ZN(y[119]) );
  OR2_X1 U235bar ( .A1(abar[7]), .A2(bbar[7]), .ZN(ybar[119]);
  AND2_X1 U236 ( .A1(a[7]), .A2(b[6]), .ZN(y[118]) );
  OR2_X1 U236bar ( .A1(abar[7]), .A2(bbar[6]), .ZN(ybar[118]);
  AND2_X1 U237 ( .A1(a[7]), .A2(b[5]), .ZN(y[117]) );
  OR2_X1 U237bar ( .A1(abar[7]), .A2(bbar[5]), .ZN(ybar[117]);
  AND2_X1 U238 ( .A1(a[7]), .A2(b[4]), .ZN(y[116]) );
  OR2_X1 U238bar ( .A1(abar[7]), .A2(bbar[4]), .ZN(ybar[116]);
  AND2_X1 U239 ( .A1(a[7]), .A2(b[3]), .ZN(y[115]) );
  OR2_X1 U239bar ( .A1(abar[7]), .A2(bbar[3]), .ZN(ybar[115]);
  AND2_X1 U240 ( .A1(a[7]), .A2(b[2]), .ZN(y[114]) );
  OR2_X1 U240bar ( .A1(abar[7]), .A2(bbar[2]), .ZN(ybar[114]);
  AND2_X1 U241 ( .A1(a[7]), .A2(b[1]), .ZN(y[113]) );
  OR2_X1 U241bar ( .A1(abar[7]), .A2(bbar[1]), .ZN(ybar[113]);
  AND2_X1 U242 ( .A1(a[7]), .A2(b[0]), .ZN(y[112]) );
  OR2_X1 U242bar ( .A1(abar[7]), .A2(bbar[0]), .ZN(ybar[112]);
  AND2_X1 U243 ( .A1(b[15]), .A2(a[6]), .ZN(y[111]) );
  OR2_X1 U243bar ( .A1(bbar[15]), .A2(abar[6]), .ZN(ybar[111]);
  AND2_X1 U244 ( .A1(b[14]), .A2(a[6]), .ZN(y[110]) );
  OR2_X1 U244bar ( .A1(bbar[14]), .A2(abar[6]), .ZN(ybar[110]);
  AND2_X1 U245 ( .A1(b[10]), .A2(a[0]), .ZN(y[10]) );
  OR2_X1 U245bar ( .A1(bbar[10]), .A2(abar[0]), .ZN(ybar[10]);
  AND2_X1 U246 ( .A1(b[13]), .A2(a[6]), .ZN(y[109]) );
  OR2_X1 U246bar ( .A1(bbar[13]), .A2(abar[6]), .ZN(ybar[109]);
  AND2_X1 U247 ( .A1(b[12]), .A2(a[6]), .ZN(y[108]) );
  OR2_X1 U247bar ( .A1(bbar[12]), .A2(abar[6]), .ZN(ybar[108]);
  AND2_X1 U248 ( .A1(b[11]), .A2(a[6]), .ZN(y[107]) );
  OR2_X1 U248bar ( .A1(bbar[11]), .A2(abar[6]), .ZN(ybar[107]);
  AND2_X1 U249 ( .A1(b[10]), .A2(a[6]), .ZN(y[106]) );
  OR2_X1 U249bar ( .A1(bbar[10]), .A2(abar[6]), .ZN(ybar[106]);
  AND2_X1 U250 ( .A1(a[6]), .A2(b[9]), .ZN(y[105]) );
  OR2_X1 U250bar ( .A1(abar[6]), .A2(bbar[9]), .ZN(ybar[105]);
  AND2_X1 U251 ( .A1(b[8]), .A2(a[6]), .ZN(y[104]) );
  OR2_X1 U251bar ( .A1(bbar[8]), .A2(abar[6]), .ZN(ybar[104]);
  AND2_X1 U252 ( .A1(b[7]), .A2(a[6]), .ZN(y[103]) );
  OR2_X1 U252bar ( .A1(bbar[7]), .A2(abar[6]), .ZN(ybar[103]);
  AND2_X1 U253 ( .A1(b[6]), .A2(a[6]), .ZN(y[102]) );
  OR2_X1 U253bar ( .A1(bbar[6]), .A2(abar[6]), .ZN(ybar[102]);
  AND2_X1 U254 ( .A1(b[5]), .A2(a[6]), .ZN(y[101]) );
  OR2_X1 U254bar ( .A1(bbar[5]), .A2(abar[6]), .ZN(ybar[101]);
  AND2_X1 U255 ( .A1(b[4]), .A2(a[6]), .ZN(y[100]) );
  OR2_X1 U255bar ( .A1(bbar[4]), .A2(abar[6]), .ZN(ybar[100]);
  AND2_X1 U256 ( .A1(b[0]), .A2(a[0]), .ZN(y[0]) );
  OR2_X1 U256bar ( .A1(bbar[0]), .A2(abar[0]), .ZN(ybar[0]);
endmodule




module decode_3 ( in, out );
  input [7:0] in;
  //input_done

  output [255:0] out;
  //output_done

  wire   [15:0] level1;
  wire   [31:0] level2;
  //wire_done

  CD2_12 cd_l1_1 ( .a(in[1]), .b(in[0]), .y(level1[3:0]) );
  CD2_11 cd_l1_2 ( .a(in[3]), .b(in[2]), .y(level1[7:4]) );
  CD2_10 cd_l1_3 ( .a(in[5]), .b(in[4]), .y(level1[11:8]) );
  CD2_9 cd_l1_4 ( .a(in[7]), .b(in[6]), .y(level1[15:12]) );
  CD4_6 cd_l2_1 ( .a(level1[7:4]), .b(level1[3:0]), .y(level2[15:0]) );
  CD4_5 cd_l2_2 ( .a(level1[15:12]), .b(level1[11:8]), .y(level2[31:16]) );
  CD16_3 cd_l3 ( .a(level2[31:16]), .b(level2[15:0]), .y(out) );
endmodule


module encode_3 ( in, out );
  input [255:0] in;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
  assign inbar[8] = ~in[8];
  assign inbar[9] = ~in[9];
  assign inbar[10] = ~in[10];
  assign inbar[11] = ~in[11];
  assign inbar[12] = ~in[12];
  assign inbar[13] = ~in[13];
  assign inbar[14] = ~in[14];
  assign inbar[15] = ~in[15];
  assign inbar[16] = ~in[16];
  assign inbar[17] = ~in[17];
  assign inbar[18] = ~in[18];
  assign inbar[19] = ~in[19];
  assign inbar[20] = ~in[20];
  assign inbar[21] = ~in[21];
  assign inbar[22] = ~in[22];
  assign inbar[23] = ~in[23];
  assign inbar[24] = ~in[24];
  assign inbar[25] = ~in[25];
  assign inbar[26] = ~in[26];
  assign inbar[27] = ~in[27];
  assign inbar[28] = ~in[28];
  assign inbar[29] = ~in[29];
  assign inbar[30] = ~in[30];
  assign inbar[31] = ~in[31];
  assign inbar[32] = ~in[32];
  assign inbar[33] = ~in[33];
  assign inbar[34] = ~in[34];
  assign inbar[35] = ~in[35];
  assign inbar[36] = ~in[36];
  assign inbar[37] = ~in[37];
  assign inbar[38] = ~in[38];
  assign inbar[39] = ~in[39];
  assign inbar[40] = ~in[40];
  assign inbar[41] = ~in[41];
  assign inbar[42] = ~in[42];
  assign inbar[43] = ~in[43];
  assign inbar[44] = ~in[44];
  assign inbar[45] = ~in[45];
  assign inbar[46] = ~in[46];
  assign inbar[47] = ~in[47];
  assign inbar[48] = ~in[48];
  assign inbar[49] = ~in[49];
  assign inbar[50] = ~in[50];
  assign inbar[51] = ~in[51];
  assign inbar[52] = ~in[52];
  assign inbar[53] = ~in[53];
  assign inbar[54] = ~in[54];
  assign inbar[55] = ~in[55];
  assign inbar[56] = ~in[56];
  assign inbar[57] = ~in[57];
  assign inbar[58] = ~in[58];
  assign inbar[59] = ~in[59];
  assign inbar[60] = ~in[60];
  assign inbar[61] = ~in[61];
  assign inbar[62] = ~in[62];
  assign inbar[63] = ~in[63];
  assign inbar[64] = ~in[64];
  assign inbar[65] = ~in[65];
  assign inbar[66] = ~in[66];
  assign inbar[67] = ~in[67];
  assign inbar[68] = ~in[68];
  assign inbar[69] = ~in[69];
  assign inbar[70] = ~in[70];
  assign inbar[71] = ~in[71];
  assign inbar[72] = ~in[72];
  assign inbar[73] = ~in[73];
  assign inbar[74] = ~in[74];
  assign inbar[75] = ~in[75];
  assign inbar[76] = ~in[76];
  assign inbar[77] = ~in[77];
  assign inbar[78] = ~in[78];
  assign inbar[79] = ~in[79];
  assign inbar[80] = ~in[80];
  assign inbar[81] = ~in[81];
  assign inbar[82] = ~in[82];
  assign inbar[83] = ~in[83];
  assign inbar[84] = ~in[84];
  assign inbar[85] = ~in[85];
  assign inbar[86] = ~in[86];
  assign inbar[87] = ~in[87];
  assign inbar[88] = ~in[88];
  assign inbar[89] = ~in[89];
  assign inbar[90] = ~in[90];
  assign inbar[91] = ~in[91];
  assign inbar[92] = ~in[92];
  assign inbar[93] = ~in[93];
  assign inbar[94] = ~in[94];
  assign inbar[95] = ~in[95];
  assign inbar[96] = ~in[96];
  assign inbar[97] = ~in[97];
  assign inbar[98] = ~in[98];
  assign inbar[99] = ~in[99];
  assign inbar[100] = ~in[100];
  assign inbar[101] = ~in[101];
  assign inbar[102] = ~in[102];
  assign inbar[103] = ~in[103];
  assign inbar[104] = ~in[104];
  assign inbar[105] = ~in[105];
  assign inbar[106] = ~in[106];
  assign inbar[107] = ~in[107];
  assign inbar[108] = ~in[108];
  assign inbar[109] = ~in[109];
  assign inbar[110] = ~in[110];
  assign inbar[111] = ~in[111];
  assign inbar[112] = ~in[112];
  assign inbar[113] = ~in[113];
  assign inbar[114] = ~in[114];
  assign inbar[115] = ~in[115];
  assign inbar[116] = ~in[116];
  assign inbar[117] = ~in[117];
  assign inbar[118] = ~in[118];
  assign inbar[119] = ~in[119];
  assign inbar[120] = ~in[120];
  assign inbar[121] = ~in[121];
  assign inbar[122] = ~in[122];
  assign inbar[123] = ~in[123];
  assign inbar[124] = ~in[124];
  assign inbar[125] = ~in[125];
  assign inbar[126] = ~in[126];
  assign inbar[127] = ~in[127];
  assign inbar[128] = ~in[128];
  assign inbar[129] = ~in[129];
  assign inbar[130] = ~in[130];
  assign inbar[131] = ~in[131];
  assign inbar[132] = ~in[132];
  assign inbar[133] = ~in[133];
  assign inbar[134] = ~in[134];
  assign inbar[135] = ~in[135];
  assign inbar[136] = ~in[136];
  assign inbar[137] = ~in[137];
  assign inbar[138] = ~in[138];
  assign inbar[139] = ~in[139];
  assign inbar[140] = ~in[140];
  assign inbar[141] = ~in[141];
  assign inbar[142] = ~in[142];
  assign inbar[143] = ~in[143];
  assign inbar[144] = ~in[144];
  assign inbar[145] = ~in[145];
  assign inbar[146] = ~in[146];
  assign inbar[147] = ~in[147];
  assign inbar[148] = ~in[148];
  assign inbar[149] = ~in[149];
  assign inbar[150] = ~in[150];
  assign inbar[151] = ~in[151];
  assign inbar[152] = ~in[152];
  assign inbar[153] = ~in[153];
  assign inbar[154] = ~in[154];
  assign inbar[155] = ~in[155];
  assign inbar[156] = ~in[156];
  assign inbar[157] = ~in[157];
  assign inbar[158] = ~in[158];
  assign inbar[159] = ~in[159];
  assign inbar[160] = ~in[160];
  assign inbar[161] = ~in[161];
  assign inbar[162] = ~in[162];
  assign inbar[163] = ~in[163];
  assign inbar[164] = ~in[164];
  assign inbar[165] = ~in[165];
  assign inbar[166] = ~in[166];
  assign inbar[167] = ~in[167];
  assign inbar[168] = ~in[168];
  assign inbar[169] = ~in[169];
  assign inbar[170] = ~in[170];
  assign inbar[171] = ~in[171];
  assign inbar[172] = ~in[172];
  assign inbar[173] = ~in[173];
  assign inbar[174] = ~in[174];
  assign inbar[175] = ~in[175];
  assign inbar[176] = ~in[176];
  assign inbar[177] = ~in[177];
  assign inbar[178] = ~in[178];
  assign inbar[179] = ~in[179];
  assign inbar[180] = ~in[180];
  assign inbar[181] = ~in[181];
  assign inbar[182] = ~in[182];
  assign inbar[183] = ~in[183];
  assign inbar[184] = ~in[184];
  assign inbar[185] = ~in[185];
  assign inbar[186] = ~in[186];
  assign inbar[187] = ~in[187];
  assign inbar[188] = ~in[188];
  assign inbar[189] = ~in[189];
  assign inbar[190] = ~in[190];
  assign inbar[191] = ~in[191];
  assign inbar[192] = ~in[192];
  assign inbar[193] = ~in[193];
  assign inbar[194] = ~in[194];
  assign inbar[195] = ~in[195];
  assign inbar[196] = ~in[196];
  assign inbar[197] = ~in[197];
  assign inbar[198] = ~in[198];
  assign inbar[199] = ~in[199];
  assign inbar[200] = ~in[200];
  assign inbar[201] = ~in[201];
  assign inbar[202] = ~in[202];
  assign inbar[203] = ~in[203];
  assign inbar[204] = ~in[204];
  assign inbar[205] = ~in[205];
  assign inbar[206] = ~in[206];
  assign inbar[207] = ~in[207];
  assign inbar[208] = ~in[208];
  assign inbar[209] = ~in[209];
  assign inbar[210] = ~in[210];
  assign inbar[211] = ~in[211];
  assign inbar[212] = ~in[212];
  assign inbar[213] = ~in[213];
  assign inbar[214] = ~in[214];
  assign inbar[215] = ~in[215];
  assign inbar[216] = ~in[216];
  assign inbar[217] = ~in[217];
  assign inbar[218] = ~in[218];
  assign inbar[219] = ~in[219];
  assign inbar[220] = ~in[220];
  assign inbar[221] = ~in[221];
  assign inbar[222] = ~in[222];
  assign inbar[223] = ~in[223];
  assign inbar[224] = ~in[224];
  assign inbar[225] = ~in[225];
  assign inbar[226] = ~in[226];
  assign inbar[227] = ~in[227];
  assign inbar[228] = ~in[228];
  assign inbar[229] = ~in[229];
  assign inbar[230] = ~in[230];
  assign inbar[231] = ~in[231];
  assign inbar[232] = ~in[232];
  assign inbar[233] = ~in[233];
  assign inbar[234] = ~in[234];
  assign inbar[235] = ~in[235];
  assign inbar[236] = ~in[236];
  assign inbar[237] = ~in[237];
  assign inbar[238] = ~in[238];
  assign inbar[239] = ~in[239];
  assign inbar[240] = ~in[240];
  assign inbar[241] = ~in[241];
  assign inbar[242] = ~in[242];
  assign inbar[243] = ~in[243];
  assign inbar[244] = ~in[244];
  assign inbar[245] = ~in[245];
  assign inbar[246] = ~in[246];
  assign inbar[247] = ~in[247];
  assign inbar[248] = ~in[248];
  assign inbar[249] = ~in[249];
  assign inbar[250] = ~in[250];
  assign inbar[251] = ~in[251];
  assign inbar[252] = ~in[252];
  assign inbar[253] = ~in[253];
  assign inbar[254] = ~in[254];
  assign inbar[255] = ~in[255];
  //input_done

  output [7:0] out;
  reg [7:0] outbar;
  //output_done

  wire   in_81, in_80, in_79, in_78, in_77, in_76, in_75, in_74, in_73, in_72,
         in_71, in_70, in_69, in_68, in_67, in_66, in_65, in_64, in_63, in_62,
         in_61, in_60, in_59, in_58, in_57, in_56, in_55, in_54, in_53, in_52,
         in_51, in_50, in_49, in_48, in_47, in_46, in_45, in_44, in_43, in_42,
         in_41, in_40, in_39, in_38, in_37, in_36, in_35, in_34, in_33, in_32,
         in_31, in_30, in_29, in_28, in_27, in_26, in_25, in_24, in_23, in_22,
         in_21, in_20, in_19, in_18, in_17, in_16, in_15, in_14, in_13, in_12,
         in_11, in_10, in_9, in_8, in_7, in_6, in_5, in_4, in_3, in_2, in_1,
         in_0, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972;
  wire in_81bar, in_80bar, in_79bar, in_78bar, in_77bar, in_76bar, in_75bar, in_74bar, in_73bar, in_72bar, in_71bar, in_70bar, in_69bar, in_68bar, in_67bar, in_66bar, in_65bar, in_64bar, in_63bar, in_62bar, in_61bar, in_60bar, in_59bar, in_58bar, in_57bar, in_56bar, in_55bar, in_54bar, in_53bar, in_52bar, in_51bar, in_50bar, in_49bar, in_48bar, in_47bar, in_46bar, in_45bar, in_44bar, in_43bar, in_42bar, in_41bar, in_40bar, in_39bar, in_38bar, in_37bar, in_36bar, in_35bar, in_34bar, in_33bar, in_32bar, in_31bar, in_30bar, in_29bar, in_28bar, in_27bar, in_26bar, in_25bar, in_24bar, in_23bar, in_22bar, in_21bar, in_20bar, in_19bar, in_18bar, in_17bar, in_16bar, in_15bar, in_14bar, in_13bar, in_12bar, in_11bar, in_10bar, in_9bar, in_8bar, in_7bar, in_6bar, in_5bar, in_4bar, in_3bar, in_2bar, in_1bar, in_0bar, n487bar, n488bar, n489bar, n490bar, n491bar, n492bar, n493bar, n494bar, n495bar, n496bar, n497bar, n498bar, n499bar, n500bar, n501bar, n502bar, n503bar, n504bar, n505bar, n506bar, n507bar, n508bar, n509bar, n510bar, n511bar, n512bar, n513bar, n514bar, n515bar, n516bar, n517bar, n518bar, n519bar, n520bar, n521bar, n522bar, n523bar, n524bar, n525bar, n526bar, n527bar, n528bar, n529bar, n530bar, n531bar, n532bar, n533bar, n534bar, n535bar, n536bar, n537bar, n538bar, n539bar, n540bar, n541bar, n542bar, n543bar, n544bar, n545bar, n546bar, n547bar, n548bar, n549bar, n550bar, n551bar, n552bar, n553bar, n554bar, n555bar, n556bar, n557bar, n558bar, n559bar, n560bar, n561bar, n562bar, n563bar, n564bar, n565bar, n566bar, n567bar, n568bar, n569bar, n570bar, n571bar, n572bar, n573bar, n574bar, n575bar, n576bar, n577bar, n578bar, n579bar, n580bar, n581bar, n582bar, n583bar, n584bar, n585bar, n586bar, n587bar, n588bar, n589bar, n590bar, n591bar, n592bar, n593bar, n594bar, n595bar, n596bar, n597bar, n598bar, n599bar, n600bar, n601bar, n602bar, n603bar, n604bar, n605bar, n606bar, n607bar, n608bar, n609bar, n610bar, n611bar, n612bar, n613bar, n614bar, n615bar, n616bar, n617bar, n618bar, n619bar, n620bar, n621bar, n622bar, n623bar, n624bar, n625bar, n626bar, n627bar, n628bar, n629bar, n630bar, n631bar, n632bar, n633bar, n634bar, n635bar, n636bar, n637bar, n638bar, n639bar, n640bar, n641bar, n642bar, n643bar, n644bar, n645bar, n646bar, n647bar, n648bar, n649bar, n650bar, n651bar, n652bar, n653bar, n654bar, n655bar, n656bar, n657bar, n658bar, n659bar, n660bar, n661bar, n662bar, n663bar, n664bar, n665bar, n666bar, n667bar, n668bar, n669bar, n670bar, n671bar, n672bar, n673bar, n674bar, n675bar, n676bar, n677bar, n678bar, n679bar, n680bar, n681bar, n682bar, n683bar, n684bar, n685bar, n686bar, n687bar, n688bar, n689bar, n690bar, n691bar, n692bar, n693bar, n694bar, n695bar, n696bar, n697bar, n698bar, n699bar, n700bar, n701bar, n702bar, n703bar, n704bar, n705bar, n706bar, n707bar, n708bar, n709bar, n710bar, n711bar, n712bar, n713bar, n714bar, n715bar, n716bar, n717bar, n718bar, n719bar, n720bar, n721bar, n722bar, n723bar, n724bar, n725bar, n726bar, n727bar, n728bar, n729bar, n730bar, n731bar, n732bar, n733bar, n734bar, n735bar, n736bar, n737bar, n738bar, n739bar, n740bar, n741bar, n742bar, n743bar, n744bar, n745bar, n746bar, n747bar, n748bar, n749bar, n750bar, n751bar, n752bar, n753bar, n754bar, n755bar, n756bar, n757bar, n758bar, n759bar, n760bar, n761bar, n762bar, n763bar, n764bar, n765bar, n766bar, n767bar, n768bar, n769bar, n770bar, n771bar, n772bar, n773bar, n774bar, n775bar, n776bar, n777bar, n778bar, n779bar, n780bar, n781bar, n782bar, n783bar, n784bar, n785bar, n786bar, n787bar, n788bar, n789bar, n790bar, n791bar, n792bar, n793bar, n794bar, n795bar, n796bar, n797bar, n798bar, n799bar, n800bar, n801bar, n802bar, n803bar, n804bar, n805bar, n806bar, n807bar, n808bar, n809bar, n810bar, n811bar, n812bar, n813bar, n814bar, n815bar, n816bar, n817bar, n818bar, n819bar, n820bar, n821bar, n822bar, n823bar, n824bar, n825bar, n826bar, n827bar, n828bar, n829bar, n830bar, n831bar, n832bar, n833bar, n834bar, n835bar, n836bar, n837bar, n838bar, n839bar, n840bar, n841bar, n842bar, n843bar, n844bar, n845bar, n846bar, n847bar, n848bar, n849bar, n850bar, n851bar, n852bar, n853bar, n854bar, n855bar, n856bar, n857bar, n858bar, n859bar, n860bar, n861bar, n862bar, n863bar, n864bar, n865bar, n866bar, n867bar, n868bar, n869bar, n870bar, n871bar, n872bar, n873bar, n874bar, n875bar, n876bar, n877bar, n878bar, n879bar, n880bar, n881bar, n882bar, n883bar, n884bar, n885bar, n886bar, n887bar, n888bar, n889bar, n890bar, n891bar, n892bar, n893bar, n894bar, n895bar, n896bar, n897bar, n898bar, n899bar, n900bar, n901bar, n902bar, n903bar, n904bar, n905bar, n906bar, n907bar, n908bar, n909bar, n910bar, n911bar, n912bar, n913bar, n914bar, n915bar, n916bar, n917bar, n918bar, n919bar, n920bar, n921bar, n922bar, n923bar, n924bar, n925bar, n926bar, n927bar, n928bar, n929bar, n930bar, n931bar, n932bar, n933bar, n934bar, n935bar, n936bar, n937bar, n938bar, n939bar, n940bar, n941bar, n942bar, n943bar, n944bar, n945bar, n946bar, n947bar, n948bar, n949bar, n950bar, n951bar, n952bar, n953bar, n954bar, n955bar, n956bar, n957bar, n958bar, n959bar, n960bar, n961bar, n962bar, n963bar, n964bar, n965bar, n966bar, n967bar, n968bar, n969bar, n970bar, n971bar, n972bar;
  //wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];

  OR2_X1 U1 ( .A1(n972), .A2(n971), .ZN(out[7]) );
  AND2_X1 U1bar ( .A1(n972bar), .A2(n971bar), .ZN(outbar[7]);
  OR2_X1 U2 ( .A1(n970), .A2(n969), .ZN(n971) );
  AND2_X1 U2bar ( .A1(n970bar), .A2(n969bar), .ZN(n971bar);
  OR2_X1 U3 ( .A1(n968), .A2(n967), .ZN(n969) );
  AND2_X1 U3bar ( .A1(n968bar), .A2(n967bar), .ZN(n969bar);
  OR2_X1 U4 ( .A1(n966), .A2(n965), .ZN(n967) );
  AND2_X1 U4bar ( .A1(n966bar), .A2(n965bar), .ZN(n967bar);
  OR2_X1 U5 ( .A1(n964), .A2(n963), .ZN(n968) );
  AND2_X1 U5bar ( .A1(n964bar), .A2(n963bar), .ZN(n968bar);
  OR2_X1 U6 ( .A1(in[116]), .A2(n962), .ZN(n963) );
  AND2_X1 U6bar ( .A1(inbar[116]), .A2(n962bar), .ZN(n963bar);
  OR2_X1 U7 ( .A1(n961), .A2(n960), .ZN(n970) );
  AND2_X1 U7bar ( .A1(n961bar), .A2(n960bar), .ZN(n970bar);
  OR2_X1 U8 ( .A1(in[150]), .A2(in[127]), .ZN(n960) );
  AND2_X1 U8bar ( .A1(inbar[150]), .A2(inbar[127]), .ZN(n960bar);
  OR2_X1 U9 ( .A1(in[160]), .A2(n959), .ZN(n961) );
  AND2_X1 U9bar ( .A1(inbar[160]), .A2(n959bar), .ZN(n961bar);
  OR2_X1 U10 ( .A1(in[252]), .A2(in[168]), .ZN(n959) );
  AND2_X1 U10bar ( .A1(inbar[252]), .A2(inbar[168]), .ZN(n959bar);
  OR2_X1 U11 ( .A1(n958), .A2(n957), .ZN(n972) );
  AND2_X1 U11bar ( .A1(n958bar), .A2(n957bar), .ZN(n972bar);
  OR2_X1 U12 ( .A1(n956), .A2(n955), .ZN(n957) );
  AND2_X1 U12bar ( .A1(n956bar), .A2(n955bar), .ZN(n957bar);
  OR2_X1 U13 ( .A1(in_17), .A2(in[96]), .ZN(n955) );
  AND2_X1 U13bar ( .A1(in_17bar), .A2(inbar[96]), .ZN(n955bar);
  OR2_X1 U14 ( .A1(in_23), .A2(n954), .ZN(n956) );
  AND2_X1 U14bar ( .A1(in_23bar), .A2(n954bar), .ZN(n956bar);
  OR2_X1 U15 ( .A1(in_31), .A2(in_26), .ZN(n954) );
  AND2_X1 U15bar ( .A1(in_31bar), .A2(in_26bar), .ZN(n954bar);
  OR2_X1 U16 ( .A1(n953), .A2(n952), .ZN(n958) );
  AND2_X1 U16bar ( .A1(n953bar), .A2(n952bar), .ZN(n958bar);
  OR2_X1 U17 ( .A1(in_58), .A2(in_4), .ZN(n952) );
  AND2_X1 U17bar ( .A1(in_58bar), .A2(in_4bar), .ZN(n952bar);
  OR2_X1 U18 ( .A1(in_59), .A2(n951), .ZN(n953) );
  AND2_X1 U18bar ( .A1(in_59bar), .A2(n951bar), .ZN(n953bar);
  OR2_X1 U19 ( .A1(in_71), .A2(in_62), .ZN(n951) );
  AND2_X1 U19bar ( .A1(in_71bar), .A2(in_62bar), .ZN(n951bar);
  OR2_X1 U20 ( .A1(n950), .A2(n949), .ZN(out[6]) );
  AND2_X1 U20bar ( .A1(n950bar), .A2(n949bar), .ZN(outbar[6]);
  OR2_X1 U21 ( .A1(n948), .A2(n947), .ZN(n949) );
  AND2_X1 U21bar ( .A1(n948bar), .A2(n947bar), .ZN(n949bar);
  OR2_X1 U22 ( .A1(n946), .A2(n945), .ZN(n947) );
  AND2_X1 U22bar ( .A1(n946bar), .A2(n945bar), .ZN(n947bar);
  OR2_X1 U23 ( .A1(n944), .A2(n943), .ZN(n945) );
  AND2_X1 U23bar ( .A1(n944bar), .A2(n943bar), .ZN(n945bar);
  OR2_X1 U24 ( .A1(n942), .A2(n941), .ZN(n946) );
  AND2_X1 U24bar ( .A1(n942bar), .A2(n941bar), .ZN(n946bar);
  OR2_X1 U25 ( .A1(in[101]), .A2(n940), .ZN(n941) );
  AND2_X1 U25bar ( .A1(inbar[101]), .A2(n940bar), .ZN(n941bar);
  OR2_X1 U26 ( .A1(n939), .A2(n938), .ZN(n948) );
  AND2_X1 U26bar ( .A1(n939bar), .A2(n938bar), .ZN(n948bar);
  OR2_X1 U27 ( .A1(in[114]), .A2(in[104]), .ZN(n938) );
  AND2_X1 U27bar ( .A1(inbar[114]), .A2(inbar[104]), .ZN(n938bar);
  OR2_X1 U28 ( .A1(in[128]), .A2(n937), .ZN(n939) );
  AND2_X1 U28bar ( .A1(inbar[128]), .A2(n937bar), .ZN(n939bar);
  OR2_X1 U29 ( .A1(in[136]), .A2(in[134]), .ZN(n937) );
  AND2_X1 U29bar ( .A1(inbar[136]), .A2(inbar[134]), .ZN(n937bar);
  OR2_X1 U30 ( .A1(n936), .A2(n935), .ZN(n950) );
  AND2_X1 U30bar ( .A1(n936bar), .A2(n935bar), .ZN(n950bar);
  OR2_X1 U31 ( .A1(n934), .A2(n933), .ZN(n935) );
  AND2_X1 U31bar ( .A1(n934bar), .A2(n933bar), .ZN(n935bar);
  OR2_X1 U32 ( .A1(in[177]), .A2(in[164]), .ZN(n933) );
  AND2_X1 U32bar ( .A1(inbar[177]), .A2(inbar[164]), .ZN(n933bar);
  OR2_X1 U33 ( .A1(in[212]), .A2(n932), .ZN(n934) );
  AND2_X1 U33bar ( .A1(inbar[212]), .A2(n932bar), .ZN(n934bar);
  OR2_X1 U34 ( .A1(in[248]), .A2(in[221]), .ZN(n932) );
  AND2_X1 U34bar ( .A1(inbar[248]), .A2(inbar[221]), .ZN(n932bar);
  OR2_X1 U35 ( .A1(n931), .A2(n930), .ZN(n936) );
  AND2_X1 U35bar ( .A1(n931bar), .A2(n930bar), .ZN(n936bar);
  OR2_X1 U36 ( .A1(in_18), .A2(in[93]), .ZN(n930) );
  AND2_X1 U36bar ( .A1(in_18bar), .A2(inbar[93]), .ZN(n930bar);
  OR2_X1 U37 ( .A1(in_31), .A2(n929), .ZN(n931) );
  AND2_X1 U37bar ( .A1(in_31bar), .A2(n929bar), .ZN(n931bar);
  OR2_X1 U38 ( .A1(in_7), .A2(in_39), .ZN(n929) );
  AND2_X1 U38bar ( .A1(in_7bar), .A2(in_39bar), .ZN(n929bar);
  OR2_X1 U39 ( .A1(n928), .A2(n927), .ZN(out[5]) );
  AND2_X1 U39bar ( .A1(n928bar), .A2(n927bar), .ZN(outbar[5]);
  OR2_X1 U40 ( .A1(n926), .A2(n925), .ZN(n927) );
  AND2_X1 U40bar ( .A1(n926bar), .A2(n925bar), .ZN(n927bar);
  OR2_X1 U41 ( .A1(n924), .A2(n923), .ZN(n925) );
  AND2_X1 U41bar ( .A1(n924bar), .A2(n923bar), .ZN(n925bar);
  OR2_X1 U42 ( .A1(n922), .A2(n921), .ZN(n923) );
  AND2_X1 U42bar ( .A1(n922bar), .A2(n921bar), .ZN(n923bar);
  OR2_X1 U43 ( .A1(n940), .A2(n920), .ZN(n924) );
  AND2_X1 U43bar ( .A1(n940bar), .A2(n920bar), .ZN(n924bar);
  OR2_X1 U44 ( .A1(in[111]), .A2(n919), .ZN(n920) );
  AND2_X1 U44bar ( .A1(inbar[111]), .A2(n919bar), .ZN(n920bar);
  OR2_X1 U45 ( .A1(n918), .A2(n917), .ZN(n940) );
  AND2_X1 U45bar ( .A1(n918bar), .A2(n917bar), .ZN(n940bar);
  OR2_X1 U46 ( .A1(n916), .A2(n915), .ZN(n917) );
  AND2_X1 U46bar ( .A1(n916bar), .A2(n915bar), .ZN(n917bar);
  OR2_X1 U47 ( .A1(n914), .A2(n913), .ZN(n915) );
  AND2_X1 U47bar ( .A1(n914bar), .A2(n913bar), .ZN(n915bar);
  OR2_X1 U48 ( .A1(in[140]), .A2(in[131]), .ZN(n913) );
  AND2_X1 U48bar ( .A1(inbar[140]), .A2(inbar[131]), .ZN(n913bar);
  OR2_X1 U49 ( .A1(in[160]), .A2(in[144]), .ZN(n914) );
  AND2_X1 U49bar ( .A1(inbar[160]), .A2(inbar[144]), .ZN(n914bar);
  OR2_X1 U50 ( .A1(n912), .A2(n911), .ZN(n916) );
  AND2_X1 U50bar ( .A1(n912bar), .A2(n911bar), .ZN(n916bar);
  OR2_X1 U51 ( .A1(in[179]), .A2(in[174]), .ZN(n911) );
  AND2_X1 U51bar ( .A1(inbar[179]), .A2(inbar[174]), .ZN(n911bar);
  OR2_X1 U52 ( .A1(in[188]), .A2(in[184]), .ZN(n912) );
  AND2_X1 U52bar ( .A1(inbar[188]), .A2(inbar[184]), .ZN(n912bar);
  OR2_X1 U53 ( .A1(n910), .A2(n909), .ZN(n918) );
  AND2_X1 U53bar ( .A1(n910bar), .A2(n909bar), .ZN(n918bar);
  OR2_X1 U54 ( .A1(n908), .A2(n907), .ZN(n909) );
  AND2_X1 U54bar ( .A1(n908bar), .A2(n907bar), .ZN(n909bar);
  OR2_X1 U55 ( .A1(in[216]), .A2(in[200]), .ZN(n907) );
  AND2_X1 U55bar ( .A1(inbar[216]), .A2(inbar[200]), .ZN(n907bar);
  OR2_X1 U56 ( .A1(in[228]), .A2(in[224]), .ZN(n908) );
  AND2_X1 U56bar ( .A1(inbar[228]), .A2(inbar[224]), .ZN(n908bar);
  OR2_X1 U57 ( .A1(n906), .A2(n905), .ZN(n910) );
  AND2_X1 U57bar ( .A1(n906bar), .A2(n905bar), .ZN(n910bar);
  OR2_X1 U58 ( .A1(in[247]), .A2(in[235]), .ZN(n905) );
  AND2_X1 U58bar ( .A1(inbar[247]), .A2(inbar[235]), .ZN(n905bar);
  OR2_X1 U59 ( .A1(in_42), .A2(in[83]), .ZN(n906) );
  AND2_X1 U59bar ( .A1(in_42bar), .A2(inbar[83]), .ZN(n906bar);
  OR2_X1 U60 ( .A1(n904), .A2(n903), .ZN(n926) );
  AND2_X1 U60bar ( .A1(n904bar), .A2(n903bar), .ZN(n926bar);
  OR2_X1 U61 ( .A1(in[166]), .A2(in[123]), .ZN(n903) );
  AND2_X1 U61bar ( .A1(inbar[166]), .A2(inbar[123]), .ZN(n903bar);
  OR2_X1 U62 ( .A1(in[170]), .A2(n902), .ZN(n904) );
  AND2_X1 U62bar ( .A1(inbar[170]), .A2(n902bar), .ZN(n904bar);
  OR2_X1 U63 ( .A1(in[194]), .A2(in[183]), .ZN(n902) );
  AND2_X1 U63bar ( .A1(inbar[194]), .A2(inbar[183]), .ZN(n902bar);
  OR2_X1 U64 ( .A1(n901), .A2(n900), .ZN(n928) );
  AND2_X1 U64bar ( .A1(n901bar), .A2(n900bar), .ZN(n928bar);
  OR2_X1 U65 ( .A1(n899), .A2(n898), .ZN(n900) );
  AND2_X1 U65bar ( .A1(n899bar), .A2(n898bar), .ZN(n900bar);
  OR2_X1 U66 ( .A1(in[241]), .A2(in[238]), .ZN(n898) );
  AND2_X1 U66bar ( .A1(inbar[241]), .A2(inbar[238]), .ZN(n898bar);
  OR2_X1 U67 ( .A1(in[250]), .A2(n897), .ZN(n899) );
  AND2_X1 U67bar ( .A1(inbar[250]), .A2(n897bar), .ZN(n899bar);
  OR2_X1 U68 ( .A1(in_24), .A2(in[84]), .ZN(n897) );
  AND2_X1 U68bar ( .A1(in_24bar), .A2(inbar[84]), .ZN(n897bar);
  OR2_X1 U69 ( .A1(n896), .A2(n895), .ZN(n901) );
  AND2_X1 U69bar ( .A1(n896bar), .A2(n895bar), .ZN(n901bar);
  OR2_X1 U70 ( .A1(in_41), .A2(in_29), .ZN(n895) );
  AND2_X1 U70bar ( .A1(in_41bar), .A2(in_29bar), .ZN(n895bar);
  OR2_X1 U71 ( .A1(in_66), .A2(n894), .ZN(n896) );
  AND2_X1 U71bar ( .A1(in_66bar), .A2(n894bar), .ZN(n896bar);
  OR2_X1 U72 ( .A1(in_76), .A2(in_71), .ZN(n894) );
  AND2_X1 U72bar ( .A1(in_76bar), .A2(in_71bar), .ZN(n894bar);
  OR2_X1 U73 ( .A1(n893), .A2(n892), .ZN(out[4]) );
  AND2_X1 U73bar ( .A1(n893bar), .A2(n892bar), .ZN(outbar[4]);
  OR2_X1 U74 ( .A1(n891), .A2(n890), .ZN(n892) );
  AND2_X1 U74bar ( .A1(n891bar), .A2(n890bar), .ZN(n892bar);
  OR2_X1 U75 ( .A1(n889), .A2(n888), .ZN(n890) );
  AND2_X1 U75bar ( .A1(n889bar), .A2(n888bar), .ZN(n890bar);
  OR2_X1 U76 ( .A1(n922), .A2(n887), .ZN(n888) );
  AND2_X1 U76bar ( .A1(n922bar), .A2(n887bar), .ZN(n888bar);
  OR2_X1 U77 ( .A1(n886), .A2(n885), .ZN(n922) );
  AND2_X1 U77bar ( .A1(n886bar), .A2(n885bar), .ZN(n922bar);
  OR2_X1 U78 ( .A1(n884), .A2(n883), .ZN(n885) );
  AND2_X1 U78bar ( .A1(n884bar), .A2(n883bar), .ZN(n885bar);
  OR2_X1 U79 ( .A1(n882), .A2(n881), .ZN(n883) );
  AND2_X1 U79bar ( .A1(n882bar), .A2(n881bar), .ZN(n883bar);
  OR2_X1 U80 ( .A1(in[118]), .A2(in[109]), .ZN(n881) );
  AND2_X1 U80bar ( .A1(inbar[118]), .A2(inbar[109]), .ZN(n881bar);
  OR2_X1 U81 ( .A1(in[139]), .A2(in[120]), .ZN(n882) );
  AND2_X1 U81bar ( .A1(inbar[139]), .A2(inbar[120]), .ZN(n882bar);
  OR2_X1 U82 ( .A1(n880), .A2(n879), .ZN(n884) );
  AND2_X1 U82bar ( .A1(n880bar), .A2(n879bar), .ZN(n884bar);
  OR2_X1 U83 ( .A1(in[198]), .A2(in[154]), .ZN(n879) );
  AND2_X1 U83bar ( .A1(inbar[198]), .A2(inbar[154]), .ZN(n879bar);
  OR2_X1 U84 ( .A1(in[210]), .A2(in[205]), .ZN(n880) );
  AND2_X1 U84bar ( .A1(inbar[210]), .A2(inbar[205]), .ZN(n880bar);
  OR2_X1 U85 ( .A1(n878), .A2(n877), .ZN(n886) );
  AND2_X1 U85bar ( .A1(n878bar), .A2(n877bar), .ZN(n886bar);
  OR2_X1 U86 ( .A1(n876), .A2(n875), .ZN(n877) );
  AND2_X1 U86bar ( .A1(n876bar), .A2(n875bar), .ZN(n877bar);
  OR2_X1 U87 ( .A1(in[219]), .A2(in[217]), .ZN(n875) );
  AND2_X1 U87bar ( .A1(inbar[219]), .A2(inbar[217]), .ZN(n875bar);
  OR2_X1 U88 ( .A1(in[86]), .A2(in[252]), .ZN(n876) );
  AND2_X1 U88bar ( .A1(inbar[86]), .A2(inbar[252]), .ZN(n876bar);
  OR2_X1 U89 ( .A1(n874), .A2(n873), .ZN(n878) );
  AND2_X1 U89bar ( .A1(n874bar), .A2(n873bar), .ZN(n878bar);
  OR2_X1 U90 ( .A1(in_40), .A2(in[91]), .ZN(n873) );
  AND2_X1 U90bar ( .A1(in_40bar), .A2(inbar[91]), .ZN(n873bar);
  OR2_X1 U91 ( .A1(in_8), .A2(in_46), .ZN(n874) );
  AND2_X1 U91bar ( .A1(in_8bar), .A2(in_46bar), .ZN(n874bar);
  OR2_X1 U92 ( .A1(n872), .A2(n871), .ZN(n889) );
  AND2_X1 U92bar ( .A1(n872bar), .A2(n871bar), .ZN(n889bar);
  OR2_X1 U93 ( .A1(in[117]), .A2(n943), .ZN(n871) );
  AND2_X1 U93bar ( .A1(inbar[117]), .A2(n943bar), .ZN(n871bar);
  OR2_X1 U94 ( .A1(n870), .A2(n869), .ZN(n943) );
  AND2_X1 U94bar ( .A1(n870bar), .A2(n869bar), .ZN(n943bar);
  OR2_X1 U95 ( .A1(n868), .A2(n867), .ZN(n869) );
  AND2_X1 U95bar ( .A1(n868bar), .A2(n867bar), .ZN(n869bar);
  OR2_X1 U96 ( .A1(n866), .A2(n865), .ZN(n867) );
  AND2_X1 U96bar ( .A1(n866bar), .A2(n865bar), .ZN(n867bar);
  OR2_X1 U97 ( .A1(n864), .A2(n863), .ZN(n865) );
  AND2_X1 U97bar ( .A1(n864bar), .A2(n863bar), .ZN(n865bar);
  OR2_X1 U98 ( .A1(in[108]), .A2(n919), .ZN(n866) );
  AND2_X1 U98bar ( .A1(inbar[108]), .A2(n919bar), .ZN(n866bar);
  OR2_X1 U99 ( .A1(n862), .A2(n861), .ZN(n919) );
  AND2_X1 U99bar ( .A1(n862bar), .A2(n861bar), .ZN(n919bar);
  OR2_X1 U100 ( .A1(n860), .A2(n859), .ZN(n861) );
  AND2_X1 U100bar ( .A1(n860bar), .A2(n859bar), .ZN(n861bar);
  OR2_X1 U101 ( .A1(n858), .A2(n857), .ZN(n859) );
  AND2_X1 U101bar ( .A1(n858bar), .A2(n857bar), .ZN(n859bar);
  OR2_X1 U102 ( .A1(in[119]), .A2(in[105]), .ZN(n857) );
  AND2_X1 U102bar ( .A1(inbar[119]), .A2(inbar[105]), .ZN(n857bar);
  OR2_X1 U103 ( .A1(in[186]), .A2(in[175]), .ZN(n858) );
  AND2_X1 U103bar ( .A1(inbar[186]), .A2(inbar[175]), .ZN(n858bar);
  OR2_X1 U104 ( .A1(n856), .A2(n855), .ZN(n860) );
  AND2_X1 U104bar ( .A1(n856bar), .A2(n855bar), .ZN(n860bar);
  OR2_X1 U105 ( .A1(in[202]), .A2(in[193]), .ZN(n855) );
  AND2_X1 U105bar ( .A1(inbar[202]), .A2(inbar[193]), .ZN(n855bar);
  OR2_X1 U106 ( .A1(in[225]), .A2(in[208]), .ZN(n856) );
  AND2_X1 U106bar ( .A1(inbar[225]), .A2(inbar[208]), .ZN(n856bar);
  OR2_X1 U107 ( .A1(n854), .A2(n853), .ZN(n862) );
  AND2_X1 U107bar ( .A1(n854bar), .A2(n853bar), .ZN(n862bar);
  OR2_X1 U108 ( .A1(n852), .A2(n851), .ZN(n853) );
  AND2_X1 U108bar ( .A1(n852bar), .A2(n851bar), .ZN(n853bar);
  OR2_X1 U109 ( .A1(in_1), .A2(in[85]), .ZN(n851) );
  AND2_X1 U109bar ( .A1(in_1bar), .A2(inbar[85]), .ZN(n851bar);
  OR2_X1 U110 ( .A1(in_23), .A2(in_19), .ZN(n852) );
  AND2_X1 U110bar ( .A1(in_23bar), .A2(in_19bar), .ZN(n852bar);
  OR2_X1 U111 ( .A1(n850), .A2(n849), .ZN(n854) );
  AND2_X1 U111bar ( .A1(n850bar), .A2(n849bar), .ZN(n854bar);
  OR2_X1 U112 ( .A1(in_43), .A2(in_33), .ZN(n849) );
  AND2_X1 U112bar ( .A1(in_43bar), .A2(in_33bar), .ZN(n849bar);
  OR2_X1 U113 ( .A1(in_63), .A2(in_44), .ZN(n850) );
  AND2_X1 U113bar ( .A1(in_63bar), .A2(in_44bar), .ZN(n850bar);
  OR2_X1 U114 ( .A1(n848), .A2(n847), .ZN(n868) );
  AND2_X1 U114bar ( .A1(n848bar), .A2(n847bar), .ZN(n868bar);
  OR2_X1 U115 ( .A1(in[141]), .A2(in[112]), .ZN(n847) );
  AND2_X1 U115bar ( .A1(inbar[141]), .A2(inbar[112]), .ZN(n847bar);
  OR2_X1 U116 ( .A1(in[147]), .A2(n846), .ZN(n848) );
  AND2_X1 U116bar ( .A1(inbar[147]), .A2(n846bar), .ZN(n848bar);
  OR2_X1 U117 ( .A1(in[181]), .A2(in[167]), .ZN(n846) );
  AND2_X1 U117bar ( .A1(inbar[181]), .A2(inbar[167]), .ZN(n846bar);
  OR2_X1 U118 ( .A1(n845), .A2(n844), .ZN(n870) );
  AND2_X1 U118bar ( .A1(n845bar), .A2(n844bar), .ZN(n870bar);
  OR2_X1 U119 ( .A1(n843), .A2(n842), .ZN(n844) );
  AND2_X1 U119bar ( .A1(n843bar), .A2(n842bar), .ZN(n844bar);
  OR2_X1 U120 ( .A1(in[229]), .A2(in[201]), .ZN(n842) );
  AND2_X1 U120bar ( .A1(inbar[229]), .A2(inbar[201]), .ZN(n842bar);
  OR2_X1 U121 ( .A1(in[237]), .A2(n841), .ZN(n843) );
  AND2_X1 U121bar ( .A1(inbar[237]), .A2(n841bar), .ZN(n843bar);
  OR2_X1 U122 ( .A1(in[94]), .A2(in[253]), .ZN(n841) );
  AND2_X1 U122bar ( .A1(inbar[94]), .A2(inbar[253]), .ZN(n841bar);
  OR2_X1 U123 ( .A1(n840), .A2(n839), .ZN(n845) );
  AND2_X1 U123bar ( .A1(n840bar), .A2(n839bar), .ZN(n845bar);
  OR2_X1 U124 ( .A1(in_21), .A2(in[96]), .ZN(n839) );
  AND2_X1 U124bar ( .A1(in_21bar), .A2(inbar[96]), .ZN(n839bar);
  OR2_X1 U125 ( .A1(in_25), .A2(n838), .ZN(n840) );
  AND2_X1 U125bar ( .A1(in_25bar), .A2(n838bar), .ZN(n840bar);
  OR2_X1 U126 ( .A1(in_81), .A2(in_45), .ZN(n838) );
  AND2_X1 U126bar ( .A1(in_81bar), .A2(in_45bar), .ZN(n838bar);
  OR2_X1 U127 ( .A1(n837), .A2(n836), .ZN(n891) );
  AND2_X1 U127bar ( .A1(n837bar), .A2(n836bar), .ZN(n891bar);
  OR2_X1 U128 ( .A1(in[142]), .A2(in[124]), .ZN(n836) );
  AND2_X1 U128bar ( .A1(inbar[142]), .A2(inbar[124]), .ZN(n836bar);
  OR2_X1 U129 ( .A1(in[150]), .A2(n835), .ZN(n837) );
  AND2_X1 U129bar ( .A1(inbar[150]), .A2(n835bar), .ZN(n837bar);
  OR2_X1 U130 ( .A1(in[172]), .A2(in[155]), .ZN(n835) );
  AND2_X1 U130bar ( .A1(inbar[172]), .A2(inbar[155]), .ZN(n835bar);
  OR2_X1 U131 ( .A1(n834), .A2(n833), .ZN(n893) );
  AND2_X1 U131bar ( .A1(n834bar), .A2(n833bar), .ZN(n893bar);
  OR2_X1 U132 ( .A1(n832), .A2(n831), .ZN(n833) );
  AND2_X1 U132bar ( .A1(n832bar), .A2(n831bar), .ZN(n833bar);
  OR2_X1 U133 ( .A1(in[196]), .A2(in[173]), .ZN(n831) );
  AND2_X1 U133bar ( .A1(inbar[196]), .A2(inbar[173]), .ZN(n831bar);
  OR2_X1 U134 ( .A1(in[222]), .A2(n830), .ZN(n832) );
  AND2_X1 U134bar ( .A1(inbar[222]), .A2(n830bar), .ZN(n832bar);
  OR2_X1 U135 ( .A1(in[227]), .A2(in[226]), .ZN(n830) );
  AND2_X1 U135bar ( .A1(inbar[227]), .A2(inbar[226]), .ZN(n830bar);
  OR2_X1 U136 ( .A1(n829), .A2(n828), .ZN(n834) );
  AND2_X1 U136bar ( .A1(n829bar), .A2(n828bar), .ZN(n834bar);
  OR2_X1 U137 ( .A1(in[249]), .A2(in[231]), .ZN(n828) );
  AND2_X1 U137bar ( .A1(inbar[249]), .A2(inbar[231]), .ZN(n828bar);
  OR2_X1 U138 ( .A1(in_28), .A2(n827), .ZN(n829) );
  AND2_X1 U138bar ( .A1(in_28bar), .A2(n827bar), .ZN(n829bar);
  OR2_X1 U139 ( .A1(in_52), .A2(in_47), .ZN(n827) );
  AND2_X1 U139bar ( .A1(in_52bar), .A2(in_47bar), .ZN(n827bar);
  OR2_X1 U140 ( .A1(n826), .A2(n825), .ZN(out[3]) );
  AND2_X1 U140bar ( .A1(n826bar), .A2(n825bar), .ZN(outbar[3]);
  OR2_X1 U141 ( .A1(n824), .A2(n823), .ZN(n825) );
  AND2_X1 U141bar ( .A1(n824bar), .A2(n823bar), .ZN(n825bar);
  OR2_X1 U142 ( .A1(n822), .A2(n821), .ZN(n823) );
  AND2_X1 U142bar ( .A1(n822bar), .A2(n821bar), .ZN(n823bar);
  OR2_X1 U143 ( .A1(n820), .A2(n819), .ZN(n821) );
  AND2_X1 U143bar ( .A1(n820bar), .A2(n819bar), .ZN(n821bar);
  OR2_X1 U144 ( .A1(n964), .A2(n818), .ZN(n822) );
  AND2_X1 U144bar ( .A1(n964bar), .A2(n818bar), .ZN(n822bar);
  OR2_X1 U145 ( .A1(in[118]), .A2(n817), .ZN(n818) );
  AND2_X1 U145bar ( .A1(inbar[118]), .A2(n817bar), .ZN(n818bar);
  OR2_X1 U146 ( .A1(n816), .A2(n815), .ZN(n964) );
  AND2_X1 U146bar ( .A1(n816bar), .A2(n815bar), .ZN(n964bar);
  OR2_X1 U147 ( .A1(n814), .A2(n813), .ZN(n815) );
  AND2_X1 U147bar ( .A1(n814bar), .A2(n813bar), .ZN(n815bar);
  OR2_X1 U148 ( .A1(n812), .A2(n811), .ZN(n813) );
  AND2_X1 U148bar ( .A1(n812bar), .A2(n811bar), .ZN(n813bar);
  OR2_X1 U149 ( .A1(in[122]), .A2(in[111]), .ZN(n811) );
  AND2_X1 U149bar ( .A1(inbar[122]), .A2(inbar[111]), .ZN(n811bar);
  OR2_X1 U150 ( .A1(in[154]), .A2(in[151]), .ZN(n812) );
  AND2_X1 U150bar ( .A1(inbar[154]), .A2(inbar[151]), .ZN(n812bar);
  OR2_X1 U151 ( .A1(n810), .A2(n809), .ZN(n814) );
  AND2_X1 U151bar ( .A1(n810bar), .A2(n809bar), .ZN(n814bar);
  OR2_X1 U152 ( .A1(in[187]), .A2(in[177]), .ZN(n809) );
  AND2_X1 U152bar ( .A1(inbar[187]), .A2(inbar[177]), .ZN(n809bar);
  OR2_X1 U153 ( .A1(in[200]), .A2(in[192]), .ZN(n810) );
  AND2_X1 U153bar ( .A1(inbar[200]), .A2(inbar[192]), .ZN(n810bar);
  OR2_X1 U154 ( .A1(n808), .A2(n807), .ZN(n816) );
  AND2_X1 U154bar ( .A1(n808bar), .A2(n807bar), .ZN(n816bar);
  OR2_X1 U155 ( .A1(n806), .A2(n805), .ZN(n807) );
  AND2_X1 U155bar ( .A1(n806bar), .A2(n805bar), .ZN(n807bar);
  OR2_X1 U156 ( .A1(in[225]), .A2(in[207]), .ZN(n805) );
  AND2_X1 U156bar ( .A1(inbar[225]), .A2(inbar[207]), .ZN(n805bar);
  OR2_X1 U157 ( .A1(in[98]), .A2(in[226]), .ZN(n806) );
  AND2_X1 U157bar ( .A1(inbar[98]), .A2(inbar[226]), .ZN(n806bar);
  OR2_X1 U158 ( .A1(n804), .A2(n803), .ZN(n808) );
  AND2_X1 U158bar ( .A1(n804bar), .A2(n803bar), .ZN(n808bar);
  OR2_X1 U159 ( .A1(in_20), .A2(in_16), .ZN(n803) );
  AND2_X1 U159bar ( .A1(in_20bar), .A2(in_16bar), .ZN(n803bar);
  OR2_X1 U160 ( .A1(in_55), .A2(in_45), .ZN(n804) );
  AND2_X1 U160bar ( .A1(in_55bar), .A2(in_45bar), .ZN(n804bar);
  OR2_X1 U161 ( .A1(n802), .A2(n801), .ZN(n824) );
  AND2_X1 U161bar ( .A1(n802bar), .A2(n801bar), .ZN(n824bar);
  OR2_X1 U162 ( .A1(in[162]), .A2(in[149]), .ZN(n801) );
  AND2_X1 U162bar ( .A1(inbar[162]), .A2(inbar[149]), .ZN(n801bar);
  OR2_X1 U163 ( .A1(in[163]), .A2(n800), .ZN(n802) );
  AND2_X1 U163bar ( .A1(inbar[163]), .A2(n800bar), .ZN(n802bar);
  OR2_X1 U164 ( .A1(in[191]), .A2(in[189]), .ZN(n800) );
  AND2_X1 U164bar ( .A1(inbar[191]), .A2(inbar[189]), .ZN(n800bar);
  OR2_X1 U165 ( .A1(n799), .A2(n798), .ZN(n826) );
  AND2_X1 U165bar ( .A1(n799bar), .A2(n798bar), .ZN(n826bar);
  OR2_X1 U166 ( .A1(n797), .A2(n796), .ZN(n798) );
  AND2_X1 U166bar ( .A1(n797bar), .A2(n796bar), .ZN(n798bar);
  OR2_X1 U167 ( .A1(in[212]), .A2(in[193]), .ZN(n796) );
  AND2_X1 U167bar ( .A1(inbar[212]), .A2(inbar[193]), .ZN(n796bar);
  OR2_X1 U168 ( .A1(in[238]), .A2(n795), .ZN(n797) );
  AND2_X1 U168bar ( .A1(inbar[238]), .A2(n795bar), .ZN(n797bar);
  OR2_X1 U169 ( .A1(in[88]), .A2(in[247]), .ZN(n795) );
  AND2_X1 U169bar ( .A1(inbar[88]), .A2(inbar[247]), .ZN(n795bar);
  OR2_X1 U170 ( .A1(n794), .A2(n793), .ZN(n799) );
  AND2_X1 U170bar ( .A1(n794bar), .A2(n793bar), .ZN(n799bar);
  OR2_X1 U171 ( .A1(in[94]), .A2(in[92]), .ZN(n793) );
  AND2_X1 U171bar ( .A1(inbar[94]), .A2(inbar[92]), .ZN(n793bar);
  OR2_X1 U172 ( .A1(in_52), .A2(n792), .ZN(n794) );
  AND2_X1 U172bar ( .A1(in_52bar), .A2(n792bar), .ZN(n794bar);
  OR2_X1 U173 ( .A1(in_70), .A2(in_67), .ZN(n792) );
  AND2_X1 U173bar ( .A1(in_70bar), .A2(in_67bar), .ZN(n792bar);
  OR2_X1 U174 ( .A1(n791), .A2(n790), .ZN(out[2]) );
  AND2_X1 U174bar ( .A1(n791bar), .A2(n790bar), .ZN(outbar[2]);
  OR2_X1 U175 ( .A1(n789), .A2(n788), .ZN(n790) );
  AND2_X1 U175bar ( .A1(n789bar), .A2(n788bar), .ZN(n790bar);
  OR2_X1 U176 ( .A1(n787), .A2(n786), .ZN(n788) );
  AND2_X1 U176bar ( .A1(n787bar), .A2(n786bar), .ZN(n788bar);
  OR2_X1 U177 ( .A1(n819), .A2(n785), .ZN(n786) );
  AND2_X1 U177bar ( .A1(n819bar), .A2(n785bar), .ZN(n786bar);
  OR2_X1 U178 ( .A1(n784), .A2(n783), .ZN(n819) );
  AND2_X1 U178bar ( .A1(n784bar), .A2(n783bar), .ZN(n819bar);
  OR2_X1 U179 ( .A1(n782), .A2(n781), .ZN(n783) );
  AND2_X1 U179bar ( .A1(n782bar), .A2(n781bar), .ZN(n783bar);
  OR2_X1 U180 ( .A1(n780), .A2(n779), .ZN(n781) );
  AND2_X1 U180bar ( .A1(n780bar), .A2(n779bar), .ZN(n781bar);
  OR2_X1 U181 ( .A1(n962), .A2(n778), .ZN(n779) );
  AND2_X1 U181bar ( .A1(n962bar), .A2(n778bar), .ZN(n779bar);
  OR2_X1 U182 ( .A1(n777), .A2(n776), .ZN(n962) );
  AND2_X1 U182bar ( .A1(n777bar), .A2(n776bar), .ZN(n962bar);
  OR2_X1 U183 ( .A1(n775), .A2(n774), .ZN(n776) );
  AND2_X1 U183bar ( .A1(n775bar), .A2(n774bar), .ZN(n776bar);
  OR2_X1 U184 ( .A1(n773), .A2(n772), .ZN(n774) );
  AND2_X1 U184bar ( .A1(n773bar), .A2(n772bar), .ZN(n774bar);
  OR2_X1 U185 ( .A1(in[131]), .A2(in[120]), .ZN(n772) );
  AND2_X1 U185bar ( .A1(inbar[131]), .A2(inbar[120]), .ZN(n772bar);
  OR2_X1 U186 ( .A1(in[153]), .A2(in[147]), .ZN(n773) );
  AND2_X1 U186bar ( .A1(inbar[153]), .A2(inbar[147]), .ZN(n773bar);
  OR2_X1 U187 ( .A1(n771), .A2(n770), .ZN(n775) );
  AND2_X1 U187bar ( .A1(n771bar), .A2(n770bar), .ZN(n775bar);
  OR2_X1 U188 ( .A1(in[170]), .A2(in[156]), .ZN(n770) );
  AND2_X1 U188bar ( .A1(inbar[170]), .A2(inbar[156]), .ZN(n770bar);
  OR2_X1 U189 ( .A1(in[223]), .A2(in[190]), .ZN(n771) );
  AND2_X1 U189bar ( .A1(inbar[223]), .A2(inbar[190]), .ZN(n771bar);
  OR2_X1 U190 ( .A1(n769), .A2(n768), .ZN(n777) );
  AND2_X1 U190bar ( .A1(n769bar), .A2(n768bar), .ZN(n777bar);
  OR2_X1 U191 ( .A1(n767), .A2(n766), .ZN(n768) );
  AND2_X1 U191bar ( .A1(n767bar), .A2(n766bar), .ZN(n768bar);
  OR2_X1 U192 ( .A1(in[236]), .A2(in[230]), .ZN(n766) );
  AND2_X1 U192bar ( .A1(inbar[236]), .A2(inbar[230]), .ZN(n766bar);
  OR2_X1 U193 ( .A1(in[85]), .A2(in[240]), .ZN(n767) );
  AND2_X1 U193bar ( .A1(inbar[85]), .A2(inbar[240]), .ZN(n767bar);
  OR2_X1 U194 ( .A1(n765), .A2(n764), .ZN(n769) );
  AND2_X1 U194bar ( .A1(n765bar), .A2(n764bar), .ZN(n769bar);
  OR2_X1 U195 ( .A1(in_12), .A2(in[90]), .ZN(n764) );
  AND2_X1 U195bar ( .A1(in_12bar), .A2(inbar[90]), .ZN(n764bar);
  OR2_X1 U196 ( .A1(in_39), .A2(in_28), .ZN(n765) );
  AND2_X1 U196bar ( .A1(in_39bar), .A2(in_28bar), .ZN(n765bar);
  OR2_X1 U197 ( .A1(in[109]), .A2(n763), .ZN(n780) );
  AND2_X1 U197bar ( .A1(inbar[109]), .A2(n763bar), .ZN(n780bar);
  OR2_X1 U198 ( .A1(n762), .A2(n761), .ZN(n782) );
  AND2_X1 U198bar ( .A1(n762bar), .A2(n761bar), .ZN(n782bar);
  OR2_X1 U199 ( .A1(in[138]), .A2(in[129]), .ZN(n761) );
  AND2_X1 U199bar ( .A1(inbar[138]), .A2(inbar[129]), .ZN(n761bar);
  OR2_X1 U200 ( .A1(in[157]), .A2(n760), .ZN(n762) );
  AND2_X1 U200bar ( .A1(inbar[157]), .A2(n760bar), .ZN(n762bar);
  OR2_X1 U201 ( .A1(in[182]), .A2(in[167]), .ZN(n760) );
  AND2_X1 U201bar ( .A1(inbar[182]), .A2(inbar[167]), .ZN(n760bar);
  OR2_X1 U202 ( .A1(n759), .A2(n758), .ZN(n784) );
  AND2_X1 U202bar ( .A1(n759bar), .A2(n758bar), .ZN(n784bar);
  OR2_X1 U203 ( .A1(n757), .A2(n756), .ZN(n758) );
  AND2_X1 U203bar ( .A1(n757bar), .A2(n756bar), .ZN(n758bar);
  OR2_X1 U204 ( .A1(in[195]), .A2(in[184]), .ZN(n756) );
  AND2_X1 U204bar ( .A1(inbar[195]), .A2(inbar[184]), .ZN(n756bar);
  OR2_X1 U205 ( .A1(in[196]), .A2(n755), .ZN(n757) );
  AND2_X1 U205bar ( .A1(inbar[196]), .A2(n755bar), .ZN(n757bar);
  OR2_X1 U206 ( .A1(in[215]), .A2(in[209]), .ZN(n755) );
  AND2_X1 U206bar ( .A1(inbar[215]), .A2(inbar[209]), .ZN(n755bar);
  OR2_X1 U207 ( .A1(n754), .A2(n753), .ZN(n759) );
  AND2_X1 U207bar ( .A1(n754bar), .A2(n753bar), .ZN(n759bar);
  OR2_X1 U208 ( .A1(in[93]), .A2(in[233]), .ZN(n753) );
  AND2_X1 U208bar ( .A1(inbar[93]), .A2(inbar[233]), .ZN(n753bar);
  OR2_X1 U209 ( .A1(in_1), .A2(n752), .ZN(n754) );
  AND2_X1 U209bar ( .A1(in_1bar), .A2(n752bar), .ZN(n754bar);
  OR2_X1 U210 ( .A1(in_69), .A2(in_66), .ZN(n752) );
  AND2_X1 U210bar ( .A1(in_69bar), .A2(in_66bar), .ZN(n752bar);
  OR2_X1 U211 ( .A1(n966), .A2(n751), .ZN(n787) );
  AND2_X1 U211bar ( .A1(n966bar), .A2(n751bar), .ZN(n787bar);
  OR2_X1 U212 ( .A1(in[134]), .A2(n750), .ZN(n751) );
  AND2_X1 U212bar ( .A1(inbar[134]), .A2(n750bar), .ZN(n751bar);
  OR2_X1 U213 ( .A1(n749), .A2(n748), .ZN(n966) );
  AND2_X1 U213bar ( .A1(n749bar), .A2(n748bar), .ZN(n966bar);
  OR2_X1 U214 ( .A1(n747), .A2(n746), .ZN(n748) );
  AND2_X1 U214bar ( .A1(n747bar), .A2(n746bar), .ZN(n748bar);
  OR2_X1 U215 ( .A1(n745), .A2(n744), .ZN(n746) );
  AND2_X1 U215bar ( .A1(n745bar), .A2(n744bar), .ZN(n746bar);
  OR2_X1 U216 ( .A1(in[136]), .A2(in[121]), .ZN(n744) );
  AND2_X1 U216bar ( .A1(inbar[136]), .A2(inbar[121]), .ZN(n744bar);
  OR2_X1 U217 ( .A1(in[186]), .A2(in[174]), .ZN(n745) );
  AND2_X1 U217bar ( .A1(inbar[186]), .A2(inbar[174]), .ZN(n745bar);
  OR2_X1 U218 ( .A1(n743), .A2(n742), .ZN(n747) );
  AND2_X1 U218bar ( .A1(n743bar), .A2(n742bar), .ZN(n747bar);
  OR2_X1 U219 ( .A1(in[198]), .A2(in[197]), .ZN(n742) );
  AND2_X1 U219bar ( .A1(inbar[198]), .A2(inbar[197]), .ZN(n742bar);
  OR2_X1 U220 ( .A1(in[214]), .A2(in[199]), .ZN(n743) );
  AND2_X1 U220bar ( .A1(inbar[214]), .A2(inbar[199]), .ZN(n743bar);
  OR2_X1 U221 ( .A1(n741), .A2(n740), .ZN(n749) );
  AND2_X1 U221bar ( .A1(n741bar), .A2(n740bar), .ZN(n749bar);
  OR2_X1 U222 ( .A1(n739), .A2(n738), .ZN(n740) );
  AND2_X1 U222bar ( .A1(n739bar), .A2(n738bar), .ZN(n740bar);
  OR2_X1 U223 ( .A1(in[231]), .A2(in[220]), .ZN(n738) );
  AND2_X1 U223bar ( .A1(inbar[231]), .A2(inbar[220]), .ZN(n738bar);
  OR2_X1 U224 ( .A1(in_25), .A2(in[245]), .ZN(n739) );
  AND2_X1 U224bar ( .A1(in_25bar), .A2(inbar[245]), .ZN(n739bar);
  OR2_X1 U225 ( .A1(n737), .A2(n736), .ZN(n741) );
  AND2_X1 U225bar ( .A1(n737bar), .A2(n736bar), .ZN(n741bar);
  OR2_X1 U226 ( .A1(in_53), .A2(in_29), .ZN(n736) );
  AND2_X1 U226bar ( .A1(in_53bar), .A2(in_29bar), .ZN(n736bar);
  OR2_X1 U227 ( .A1(in_79), .A2(in_74), .ZN(n737) );
  AND2_X1 U227bar ( .A1(in_79bar), .A2(in_74bar), .ZN(n737bar);
  OR2_X1 U228 ( .A1(n735), .A2(n734), .ZN(n789) );
  AND2_X1 U228bar ( .A1(n735bar), .A2(n734bar), .ZN(n789bar);
  OR2_X1 U229 ( .A1(in[152]), .A2(in[140]), .ZN(n734) );
  AND2_X1 U229bar ( .A1(inbar[152]), .A2(inbar[140]), .ZN(n734bar);
  OR2_X1 U230 ( .A1(in[155]), .A2(n733), .ZN(n735) );
  AND2_X1 U230bar ( .A1(inbar[155]), .A2(n733bar), .ZN(n735bar);
  OR2_X1 U231 ( .A1(in[166]), .A2(in[165]), .ZN(n733) );
  AND2_X1 U231bar ( .A1(inbar[166]), .A2(inbar[165]), .ZN(n733bar);
  OR2_X1 U232 ( .A1(n732), .A2(n731), .ZN(n791) );
  AND2_X1 U232bar ( .A1(n732bar), .A2(n731bar), .ZN(n791bar);
  OR2_X1 U233 ( .A1(n730), .A2(n729), .ZN(n731) );
  AND2_X1 U233bar ( .A1(n730bar), .A2(n729bar), .ZN(n731bar);
  OR2_X1 U234 ( .A1(in[202]), .A2(in[185]), .ZN(n729) );
  AND2_X1 U234bar ( .A1(inbar[202]), .A2(inbar[185]), .ZN(n729bar);
  OR2_X1 U235 ( .A1(in[211]), .A2(n728), .ZN(n730) );
  AND2_X1 U235bar ( .A1(inbar[211]), .A2(n728bar), .ZN(n730bar);
  OR2_X1 U236 ( .A1(in[255]), .A2(in[253]), .ZN(n728) );
  AND2_X1 U236bar ( .A1(inbar[255]), .A2(inbar[253]), .ZN(n728bar);
  OR2_X1 U237 ( .A1(n727), .A2(n726), .ZN(n732) );
  AND2_X1 U237bar ( .A1(n727bar), .A2(n726bar), .ZN(n732bar);
  OR2_X1 U238 ( .A1(in_35), .A2(in_15), .ZN(n726) );
  AND2_X1 U238bar ( .A1(in_35bar), .A2(in_15bar), .ZN(n726bar);
  OR2_X1 U239 ( .A1(in_36), .A2(n725), .ZN(n727) );
  AND2_X1 U239bar ( .A1(in_36bar), .A2(n725bar), .ZN(n727bar);
  OR2_X1 U240 ( .A1(in_48), .A2(in_40), .ZN(n725) );
  AND2_X1 U240bar ( .A1(in_48bar), .A2(in_40bar), .ZN(n725bar);
  OR2_X1 U241 ( .A1(n724), .A2(n723), .ZN(out[1]) );
  AND2_X1 U241bar ( .A1(n724bar), .A2(n723bar), .ZN(outbar[1]);
  OR2_X1 U242 ( .A1(n722), .A2(n721), .ZN(n723) );
  AND2_X1 U242bar ( .A1(n722bar), .A2(n721bar), .ZN(n723bar);
  OR2_X1 U243 ( .A1(n720), .A2(n719), .ZN(n721) );
  AND2_X1 U243bar ( .A1(n720bar), .A2(n719bar), .ZN(n721bar);
  OR2_X1 U244 ( .A1(n921), .A2(n887), .ZN(n719) );
  AND2_X1 U244bar ( .A1(n921bar), .A2(n887bar), .ZN(n719bar);
  OR2_X1 U245 ( .A1(n718), .A2(n717), .ZN(n887) );
  AND2_X1 U245bar ( .A1(n718bar), .A2(n717bar), .ZN(n887bar);
  OR2_X1 U246 ( .A1(n716), .A2(n715), .ZN(n717) );
  AND2_X1 U246bar ( .A1(n716bar), .A2(n715bar), .ZN(n717bar);
  OR2_X1 U247 ( .A1(n714), .A2(n713), .ZN(n715) );
  AND2_X1 U247bar ( .A1(n714bar), .A2(n713bar), .ZN(n715bar);
  OR2_X1 U248 ( .A1(in[116]), .A2(in[110]), .ZN(n713) );
  AND2_X1 U248bar ( .A1(inbar[116]), .A2(inbar[110]), .ZN(n713bar);
  OR2_X1 U249 ( .A1(in[133]), .A2(in[130]), .ZN(n714) );
  AND2_X1 U249bar ( .A1(inbar[133]), .A2(inbar[130]), .ZN(n714bar);
  OR2_X1 U250 ( .A1(n712), .A2(n711), .ZN(n716) );
  AND2_X1 U250bar ( .A1(n712bar), .A2(n711bar), .ZN(n716bar);
  OR2_X1 U251 ( .A1(in[203]), .A2(in[135]), .ZN(n711) );
  AND2_X1 U251bar ( .A1(inbar[203]), .A2(inbar[135]), .ZN(n711bar);
  OR2_X1 U252 ( .A1(in[232]), .A2(in[223]), .ZN(n712) );
  AND2_X1 U252bar ( .A1(inbar[232]), .A2(inbar[223]), .ZN(n712bar);
  OR2_X1 U253 ( .A1(n710), .A2(n709), .ZN(n718) );
  AND2_X1 U253bar ( .A1(n710bar), .A2(n709bar), .ZN(n718bar);
  OR2_X1 U254 ( .A1(n708), .A2(n707), .ZN(n709) );
  AND2_X1 U254bar ( .A1(n708bar), .A2(n707bar), .ZN(n709bar);
  OR2_X1 U255 ( .A1(in[255]), .A2(in[233]), .ZN(n707) );
  AND2_X1 U255bar ( .A1(inbar[255]), .A2(inbar[233]), .ZN(n707bar);
  OR2_X1 U256 ( .A1(in_53), .A2(in_34), .ZN(n708) );
  AND2_X1 U256bar ( .A1(in_53bar), .A2(in_34bar), .ZN(n708bar);
  OR2_X1 U257 ( .A1(n706), .A2(n705), .ZN(n710) );
  AND2_X1 U257bar ( .A1(n706bar), .A2(n705bar), .ZN(n710bar);
  OR2_X1 U258 ( .A1(in_57), .A2(in_55), .ZN(n705) );
  AND2_X1 U258bar ( .A1(in_57bar), .A2(in_55bar), .ZN(n705bar);
  OR2_X1 U259 ( .A1(in_68), .A2(in_67), .ZN(n706) );
  AND2_X1 U259bar ( .A1(in_68bar), .A2(in_67bar), .ZN(n706bar);
  OR2_X1 U260 ( .A1(n704), .A2(n703), .ZN(n921) );
  AND2_X1 U260bar ( .A1(n704bar), .A2(n703bar), .ZN(n921bar);
  OR2_X1 U261 ( .A1(n702), .A2(n701), .ZN(n703) );
  AND2_X1 U261bar ( .A1(n702bar), .A2(n701bar), .ZN(n703bar);
  OR2_X1 U262 ( .A1(n700), .A2(n699), .ZN(n701) );
  AND2_X1 U262bar ( .A1(n700bar), .A2(n699bar), .ZN(n701bar);
  OR2_X1 U263 ( .A1(n944), .A2(n872), .ZN(n699) );
  AND2_X1 U263bar ( .A1(n944bar), .A2(n872bar), .ZN(n699bar);
  OR2_X1 U264 ( .A1(n698), .A2(n697), .ZN(n872) );
  AND2_X1 U264bar ( .A1(n698bar), .A2(n697bar), .ZN(n872bar);
  OR2_X1 U265 ( .A1(n696), .A2(n695), .ZN(n697) );
  AND2_X1 U265bar ( .A1(n696bar), .A2(n695bar), .ZN(n697bar);
  OR2_X1 U266 ( .A1(n694), .A2(n693), .ZN(n695) );
  AND2_X1 U266bar ( .A1(n694bar), .A2(n693bar), .ZN(n695bar);
  OR2_X1 U267 ( .A1(in[121]), .A2(in[102]), .ZN(n693) );
  AND2_X1 U267bar ( .A1(inbar[121]), .A2(inbar[102]), .ZN(n693bar);
  OR2_X1 U268 ( .A1(in[162]), .A2(in[161]), .ZN(n694) );
  AND2_X1 U268bar ( .A1(inbar[162]), .A2(inbar[161]), .ZN(n694bar);
  OR2_X1 U269 ( .A1(n692), .A2(n691), .ZN(n696) );
  AND2_X1 U269bar ( .A1(n692bar), .A2(n691bar), .ZN(n696bar);
  OR2_X1 U270 ( .A1(in[192]), .A2(in[178]), .ZN(n691) );
  AND2_X1 U270bar ( .A1(inbar[192]), .A2(inbar[178]), .ZN(n691bar);
  OR2_X1 U271 ( .A1(in[244]), .A2(in[209]), .ZN(n692) );
  AND2_X1 U271bar ( .A1(inbar[244]), .A2(inbar[209]), .ZN(n692bar);
  OR2_X1 U272 ( .A1(n690), .A2(n689), .ZN(n698) );
  AND2_X1 U272bar ( .A1(n690bar), .A2(n689bar), .ZN(n698bar);
  OR2_X1 U273 ( .A1(n688), .A2(n687), .ZN(n689) );
  AND2_X1 U273bar ( .A1(n688bar), .A2(n687bar), .ZN(n689bar);
  OR2_X1 U274 ( .A1(in[90]), .A2(in[254]), .ZN(n687) );
  AND2_X1 U274bar ( .A1(inbar[90]), .A2(inbar[254]), .ZN(n687bar);
  OR2_X1 U275 ( .A1(in_36), .A2(in_32), .ZN(n688) );
  AND2_X1 U275bar ( .A1(in_36bar), .A2(in_32bar), .ZN(n688bar);
  OR2_X1 U276 ( .A1(n686), .A2(n685), .ZN(n690) );
  AND2_X1 U276bar ( .A1(n686bar), .A2(n685bar), .ZN(n690bar);
  OR2_X1 U277 ( .A1(in_62), .A2(in_37), .ZN(n685) );
  AND2_X1 U277bar ( .A1(in_62bar), .A2(in_37bar), .ZN(n685bar);
  OR2_X1 U278 ( .A1(in_75), .A2(in_73), .ZN(n686) );
  AND2_X1 U278bar ( .A1(in_75bar), .A2(in_73bar), .ZN(n686bar);
  OR2_X1 U279 ( .A1(n684), .A2(n683), .ZN(n944) );
  AND2_X1 U279bar ( .A1(n684bar), .A2(n683bar), .ZN(n944bar);
  OR2_X1 U280 ( .A1(n682), .A2(n681), .ZN(n683) );
  AND2_X1 U280bar ( .A1(n682bar), .A2(n681bar), .ZN(n683bar);
  OR2_X1 U281 ( .A1(n680), .A2(n679), .ZN(n681) );
  AND2_X1 U281bar ( .A1(n680bar), .A2(n679bar), .ZN(n681bar);
  OR2_X1 U282 ( .A1(in[171]), .A2(in[153]), .ZN(n679) );
  AND2_X1 U282bar ( .A1(inbar[171]), .A2(inbar[153]), .ZN(n679bar);
  OR2_X1 U283 ( .A1(in[187]), .A2(in[176]), .ZN(n680) );
  AND2_X1 U283bar ( .A1(inbar[187]), .A2(inbar[176]), .ZN(n680bar);
  OR2_X1 U284 ( .A1(n678), .A2(n677), .ZN(n682) );
  AND2_X1 U284bar ( .A1(n678bar), .A2(n677bar), .ZN(n682bar);
  OR2_X1 U285 ( .A1(in[245]), .A2(in[211]), .ZN(n677) );
  AND2_X1 U285bar ( .A1(inbar[245]), .A2(inbar[211]), .ZN(n677bar);
  OR2_X1 U286 ( .A1(in[97]), .A2(in[88]), .ZN(n678) );
  AND2_X1 U286bar ( .A1(inbar[97]), .A2(inbar[88]), .ZN(n678bar);
  OR2_X1 U287 ( .A1(n676), .A2(n675), .ZN(n684) );
  AND2_X1 U287bar ( .A1(n676bar), .A2(n675bar), .ZN(n684bar);
  OR2_X1 U288 ( .A1(n674), .A2(n673), .ZN(n675) );
  AND2_X1 U288bar ( .A1(n674bar), .A2(n673bar), .ZN(n675bar);
  OR2_X1 U289 ( .A1(in_10), .A2(in_0), .ZN(n673) );
  AND2_X1 U289bar ( .A1(in_10bar), .A2(in_0bar), .ZN(n673bar);
  OR2_X1 U290 ( .A1(in_59), .A2(in_5), .ZN(n674) );
  AND2_X1 U290bar ( .A1(in_59bar), .A2(in_5bar), .ZN(n674bar);
  OR2_X1 U291 ( .A1(n672), .A2(n671), .ZN(n676) );
  AND2_X1 U291bar ( .A1(n672bar), .A2(n671bar), .ZN(n676bar);
  OR2_X1 U292 ( .A1(in_60), .A2(in_6), .ZN(n671) );
  AND2_X1 U292bar ( .A1(in_60bar), .A2(in_6bar), .ZN(n671bar);
  OR2_X1 U293 ( .A1(in_77), .A2(in_69), .ZN(n672) );
  AND2_X1 U293bar ( .A1(in_77bar), .A2(in_69bar), .ZN(n672bar);
  OR2_X1 U294 ( .A1(in[113]), .A2(n864), .ZN(n700) );
  AND2_X1 U294bar ( .A1(inbar[113]), .A2(n864bar), .ZN(n700bar);
  OR2_X1 U295 ( .A1(n670), .A2(n669), .ZN(n864) );
  AND2_X1 U295bar ( .A1(n670bar), .A2(n669bar), .ZN(n864bar);
  OR2_X1 U296 ( .A1(n668), .A2(n667), .ZN(n669) );
  AND2_X1 U296bar ( .A1(n668bar), .A2(n667bar), .ZN(n669bar);
  OR2_X1 U297 ( .A1(n666), .A2(n665), .ZN(n667) );
  AND2_X1 U297bar ( .A1(n666bar), .A2(n665bar), .ZN(n667bar);
  OR2_X1 U298 ( .A1(in[125]), .A2(in[107]), .ZN(n665) );
  AND2_X1 U298bar ( .A1(inbar[125]), .A2(inbar[107]), .ZN(n665bar);
  OR2_X1 U299 ( .A1(in[138]), .A2(in[126]), .ZN(n666) );
  AND2_X1 U299bar ( .A1(inbar[138]), .A2(inbar[126]), .ZN(n666bar);
  OR2_X1 U300 ( .A1(n664), .A2(n663), .ZN(n668) );
  AND2_X1 U300bar ( .A1(n664bar), .A2(n663bar), .ZN(n668bar);
  OR2_X1 U301 ( .A1(in[189]), .A2(in[143]), .ZN(n663) );
  AND2_X1 U301bar ( .A1(inbar[189]), .A2(inbar[143]), .ZN(n663bar);
  OR2_X1 U302 ( .A1(in[99]), .A2(in[214]), .ZN(n664) );
  AND2_X1 U302bar ( .A1(inbar[99]), .A2(inbar[214]), .ZN(n664bar);
  OR2_X1 U303 ( .A1(n662), .A2(n661), .ZN(n670) );
  AND2_X1 U303bar ( .A1(n662bar), .A2(n661bar), .ZN(n670bar);
  OR2_X1 U304 ( .A1(n660), .A2(n659), .ZN(n661) );
  AND2_X1 U304bar ( .A1(n660bar), .A2(n659bar), .ZN(n661bar);
  OR2_X1 U305 ( .A1(in_15), .A2(in_12), .ZN(n659) );
  AND2_X1 U305bar ( .A1(in_15bar), .A2(in_12bar), .ZN(n659bar);
  OR2_X1 U306 ( .A1(in_20), .A2(in_2), .ZN(n660) );
  AND2_X1 U306bar ( .A1(in_20bar), .A2(in_2bar), .ZN(n660bar);
  OR2_X1 U307 ( .A1(n658), .A2(n657), .ZN(n662) );
  AND2_X1 U307bar ( .A1(n658bar), .A2(n657bar), .ZN(n662bar);
  OR2_X1 U308 ( .A1(in_30), .A2(in_3), .ZN(n657) );
  AND2_X1 U308bar ( .A1(in_30bar), .A2(in_3bar), .ZN(n657bar);
  OR2_X1 U309 ( .A1(in_4), .A2(in_38), .ZN(n658) );
  AND2_X1 U309bar ( .A1(in_4bar), .A2(in_38bar), .ZN(n658bar);
  OR2_X1 U310 ( .A1(n656), .A2(n655), .ZN(n702) );
  AND2_X1 U310bar ( .A1(n656bar), .A2(n655bar), .ZN(n702bar);
  OR2_X1 U311 ( .A1(in[148]), .A2(in[137]), .ZN(n655) );
  AND2_X1 U311bar ( .A1(inbar[148]), .A2(inbar[137]), .ZN(n655bar);
  OR2_X1 U312 ( .A1(in[149]), .A2(n654), .ZN(n656) );
  AND2_X1 U312bar ( .A1(inbar[149]), .A2(n654bar), .ZN(n656bar);
  OR2_X1 U313 ( .A1(in[195]), .A2(in[190]), .ZN(n654) );
  AND2_X1 U313bar ( .A1(inbar[195]), .A2(inbar[190]), .ZN(n654bar);
  OR2_X1 U314 ( .A1(n653), .A2(n652), .ZN(n704) );
  AND2_X1 U314bar ( .A1(n653bar), .A2(n652bar), .ZN(n704bar);
  OR2_X1 U315 ( .A1(n651), .A2(n650), .ZN(n652) );
  AND2_X1 U315bar ( .A1(n651bar), .A2(n650bar), .ZN(n652bar);
  OR2_X1 U316 ( .A1(in[98]), .A2(in[197]), .ZN(n650) );
  AND2_X1 U316bar ( .A1(inbar[98]), .A2(inbar[197]), .ZN(n650bar);
  OR2_X1 U317 ( .A1(in_11), .A2(n649), .ZN(n651) );
  AND2_X1 U317bar ( .A1(in_11bar), .A2(n649bar), .ZN(n651bar);
  OR2_X1 U318 ( .A1(in_26), .A2(in_14), .ZN(n649) );
  AND2_X1 U318bar ( .A1(in_26bar), .A2(in_14bar), .ZN(n649bar);
  OR2_X1 U319 ( .A1(n648), .A2(n647), .ZN(n653) );
  AND2_X1 U319bar ( .A1(n648bar), .A2(n647bar), .ZN(n653bar);
  OR2_X1 U320 ( .A1(in_35), .A2(in_27), .ZN(n647) );
  AND2_X1 U320bar ( .A1(in_35bar), .A2(in_27bar), .ZN(n647bar);
  OR2_X1 U321 ( .A1(in_50), .A2(n646), .ZN(n648) );
  AND2_X1 U321bar ( .A1(in_50bar), .A2(n646bar), .ZN(n648bar);
  OR2_X1 U322 ( .A1(in_78), .A2(in_61), .ZN(n646) );
  AND2_X1 U322bar ( .A1(in_78bar), .A2(in_61bar), .ZN(n646bar);
  OR2_X1 U323 ( .A1(n942), .A2(n645), .ZN(n720) );
  AND2_X1 U323bar ( .A1(n942bar), .A2(n645bar), .ZN(n720bar);
  OR2_X1 U324 ( .A1(in[106]), .A2(n863), .ZN(n645) );
  AND2_X1 U324bar ( .A1(inbar[106]), .A2(n863bar), .ZN(n645bar);
  OR2_X1 U325 ( .A1(n644), .A2(n643), .ZN(n863) );
  AND2_X1 U325bar ( .A1(n644bar), .A2(n643bar), .ZN(n863bar);
  OR2_X1 U326 ( .A1(n642), .A2(n641), .ZN(n643) );
  AND2_X1 U326bar ( .A1(n642bar), .A2(n641bar), .ZN(n643bar);
  OR2_X1 U327 ( .A1(n640), .A2(n639), .ZN(n641) );
  AND2_X1 U327bar ( .A1(n640bar), .A2(n639bar), .ZN(n641bar);
  OR2_X1 U328 ( .A1(in[127]), .A2(in[122]), .ZN(n639) );
  AND2_X1 U328bar ( .A1(inbar[127]), .A2(inbar[122]), .ZN(n639bar);
  OR2_X1 U329 ( .A1(in[156]), .A2(in[132]), .ZN(n640) );
  AND2_X1 U329bar ( .A1(inbar[156]), .A2(inbar[132]), .ZN(n640bar);
  OR2_X1 U330 ( .A1(n638), .A2(n637), .ZN(n642) );
  AND2_X1 U330bar ( .A1(n638bar), .A2(n637bar), .ZN(n642bar);
  OR2_X1 U331 ( .A1(in[159]), .A2(in[157]), .ZN(n637) );
  AND2_X1 U331bar ( .A1(inbar[159]), .A2(inbar[157]), .ZN(n637bar);
  OR2_X1 U332 ( .A1(in[185]), .A2(in[169]), .ZN(n638) );
  AND2_X1 U332bar ( .A1(inbar[185]), .A2(inbar[169]), .ZN(n638bar);
  OR2_X1 U333 ( .A1(n636), .A2(n635), .ZN(n644) );
  AND2_X1 U333bar ( .A1(n636bar), .A2(n635bar), .ZN(n644bar);
  OR2_X1 U334 ( .A1(n634), .A2(n633), .ZN(n635) );
  AND2_X1 U334bar ( .A1(n634bar), .A2(n633bar), .ZN(n635bar);
  OR2_X1 U335 ( .A1(in[239]), .A2(in[218]), .ZN(n633) );
  AND2_X1 U335bar ( .A1(inbar[239]), .A2(inbar[218]), .ZN(n633bar);
  OR2_X1 U336 ( .A1(in_13), .A2(in[87]), .ZN(n634) );
  AND2_X1 U336bar ( .A1(in_13bar), .A2(inbar[87]), .ZN(n634bar);
  OR2_X1 U337 ( .A1(n632), .A2(n631), .ZN(n636) );
  AND2_X1 U337bar ( .A1(n632bar), .A2(n631bar), .ZN(n636bar);
  OR2_X1 U338 ( .A1(in_72), .A2(in_70), .ZN(n631) );
  AND2_X1 U338bar ( .A1(in_72bar), .A2(in_70bar), .ZN(n631bar);
  OR2_X1 U339 ( .A1(in_80), .A2(in_74), .ZN(n632) );
  AND2_X1 U339bar ( .A1(in_80bar), .A2(in_74bar), .ZN(n632bar);
  OR2_X1 U340 ( .A1(n630), .A2(n629), .ZN(n942) );
  AND2_X1 U340bar ( .A1(n630bar), .A2(n629bar), .ZN(n942bar);
  OR2_X1 U341 ( .A1(n628), .A2(n627), .ZN(n629) );
  AND2_X1 U341bar ( .A1(n628bar), .A2(n627bar), .ZN(n629bar);
  OR2_X1 U342 ( .A1(n626), .A2(n625), .ZN(n627) );
  AND2_X1 U342bar ( .A1(n626bar), .A2(n625bar), .ZN(n627bar);
  OR2_X1 U343 ( .A1(in[146]), .A2(in[100]), .ZN(n625) );
  AND2_X1 U343bar ( .A1(inbar[146]), .A2(inbar[100]), .ZN(n625bar);
  OR2_X1 U344 ( .A1(in[168]), .A2(in[152]), .ZN(n626) );
  AND2_X1 U344bar ( .A1(inbar[168]), .A2(inbar[152]), .ZN(n626bar);
  OR2_X1 U345 ( .A1(n624), .A2(n623), .ZN(n628) );
  AND2_X1 U345bar ( .A1(n624bar), .A2(n623bar), .ZN(n628bar);
  OR2_X1 U346 ( .A1(in[199]), .A2(in[182]), .ZN(n623) );
  AND2_X1 U346bar ( .A1(inbar[199]), .A2(inbar[182]), .ZN(n623bar);
  OR2_X1 U347 ( .A1(in[236]), .A2(in[204]), .ZN(n624) );
  AND2_X1 U347bar ( .A1(inbar[236]), .A2(inbar[204]), .ZN(n624bar);
  OR2_X1 U348 ( .A1(n622), .A2(n621), .ZN(n630) );
  AND2_X1 U348bar ( .A1(n622bar), .A2(n621bar), .ZN(n630bar);
  OR2_X1 U349 ( .A1(n620), .A2(n619), .ZN(n621) );
  AND2_X1 U349bar ( .A1(n620bar), .A2(n619bar), .ZN(n621bar);
  OR2_X1 U350 ( .A1(in[89]), .A2(in[246]), .ZN(n619) );
  AND2_X1 U350bar ( .A1(inbar[89]), .A2(inbar[246]), .ZN(n619bar);
  OR2_X1 U351 ( .A1(in[95]), .A2(in[92]), .ZN(n620) );
  AND2_X1 U351bar ( .A1(inbar[95]), .A2(inbar[92]), .ZN(n620bar);
  OR2_X1 U352 ( .A1(n618), .A2(n617), .ZN(n622) );
  AND2_X1 U352bar ( .A1(n618bar), .A2(n617bar), .ZN(n622bar);
  OR2_X1 U353 ( .A1(in_22), .A2(in_16), .ZN(n617) );
  AND2_X1 U353bar ( .A1(in_22bar), .A2(in_16bar), .ZN(n617bar);
  OR2_X1 U354 ( .A1(in_51), .A2(in_49), .ZN(n618) );
  AND2_X1 U354bar ( .A1(in_51bar), .A2(in_49bar), .ZN(n618bar);
  OR2_X1 U355 ( .A1(n616), .A2(n615), .ZN(n722) );
  AND2_X1 U355bar ( .A1(n616bar), .A2(n615bar), .ZN(n722bar);
  OR2_X1 U356 ( .A1(in[158]), .A2(in[115]), .ZN(n615) );
  AND2_X1 U356bar ( .A1(inbar[158]), .A2(inbar[115]), .ZN(n615bar);
  OR2_X1 U357 ( .A1(in[163]), .A2(n614), .ZN(n616) );
  AND2_X1 U357bar ( .A1(inbar[163]), .A2(n614bar), .ZN(n616bar);
  OR2_X1 U358 ( .A1(in[206]), .A2(in[165]), .ZN(n614) );
  AND2_X1 U358bar ( .A1(inbar[206]), .A2(inbar[165]), .ZN(n614bar);
  OR2_X1 U359 ( .A1(n613), .A2(n612), .ZN(n724) );
  AND2_X1 U359bar ( .A1(n613bar), .A2(n612bar), .ZN(n724bar);
  OR2_X1 U360 ( .A1(n611), .A2(n610), .ZN(n612) );
  AND2_X1 U360bar ( .A1(n611bar), .A2(n610bar), .ZN(n612bar);
  OR2_X1 U361 ( .A1(in[213]), .A2(in[207]), .ZN(n610) );
  AND2_X1 U361bar ( .A1(inbar[213]), .A2(inbar[207]), .ZN(n610bar);
  OR2_X1 U362 ( .A1(in[215]), .A2(n609), .ZN(n611) );
  AND2_X1 U362bar ( .A1(inbar[215]), .A2(n609bar), .ZN(n611bar);
  OR2_X1 U363 ( .A1(in[230]), .A2(in[220]), .ZN(n609) );
  AND2_X1 U363bar ( .A1(inbar[230]), .A2(inbar[220]), .ZN(n609bar);
  OR2_X1 U364 ( .A1(n608), .A2(n607), .ZN(n613) );
  AND2_X1 U364bar ( .A1(n608bar), .A2(n607bar), .ZN(n613bar);
  OR2_X1 U365 ( .A1(in[251]), .A2(in[234]), .ZN(n607) );
  AND2_X1 U365bar ( .A1(inbar[251]), .A2(inbar[234]), .ZN(n607bar);
  OR2_X1 U366 ( .A1(in_17), .A2(n606), .ZN(n608) );
  AND2_X1 U366bar ( .A1(in_17bar), .A2(n606bar), .ZN(n608bar);
  OR2_X1 U367 ( .A1(in_65), .A2(in_56), .ZN(n606) );
  AND2_X1 U367bar ( .A1(in_65bar), .A2(in_56bar), .ZN(n606bar);
  OR2_X1 U368 ( .A1(n605), .A2(n604), .ZN(out[0]) );
  AND2_X1 U368bar ( .A1(n605bar), .A2(n604bar), .ZN(outbar[0]);
  OR2_X1 U369 ( .A1(n603), .A2(n602), .ZN(n604) );
  AND2_X1 U369bar ( .A1(n603bar), .A2(n602bar), .ZN(n604bar);
  OR2_X1 U370 ( .A1(n601), .A2(n600), .ZN(n602) );
  AND2_X1 U370bar ( .A1(n601bar), .A2(n600bar), .ZN(n602bar);
  OR2_X1 U371 ( .A1(n820), .A2(n785), .ZN(n600) );
  AND2_X1 U371bar ( .A1(n820bar), .A2(n785bar), .ZN(n600bar);
  OR2_X1 U372 ( .A1(n599), .A2(n598), .ZN(n785) );
  AND2_X1 U372bar ( .A1(n599bar), .A2(n598bar), .ZN(n785bar);
  OR2_X1 U373 ( .A1(n597), .A2(n596), .ZN(n598) );
  AND2_X1 U373bar ( .A1(n597bar), .A2(n596bar), .ZN(n598bar);
  OR2_X1 U374 ( .A1(n595), .A2(n594), .ZN(n596) );
  AND2_X1 U374bar ( .A1(n595bar), .A2(n594bar), .ZN(n596bar);
  OR2_X1 U375 ( .A1(in[135]), .A2(in[104]), .ZN(n594) );
  AND2_X1 U375bar ( .A1(inbar[135]), .A2(inbar[104]), .ZN(n594bar);
  OR2_X1 U376 ( .A1(in[188]), .A2(in[178]), .ZN(n595) );
  AND2_X1 U376bar ( .A1(inbar[188]), .A2(inbar[178]), .ZN(n595bar);
  OR2_X1 U377 ( .A1(n593), .A2(n592), .ZN(n597) );
  AND2_X1 U377bar ( .A1(n593bar), .A2(n592bar), .ZN(n597bar);
  OR2_X1 U378 ( .A1(in[217]), .A2(in[194]), .ZN(n592) );
  AND2_X1 U378bar ( .A1(inbar[217]), .A2(inbar[194]), .ZN(n592bar);
  OR2_X1 U379 ( .A1(in[237]), .A2(in[218]), .ZN(n593) );
  AND2_X1 U379bar ( .A1(inbar[237]), .A2(inbar[218]), .ZN(n593bar);
  OR2_X1 U380 ( .A1(n591), .A2(n590), .ZN(n599) );
  AND2_X1 U380bar ( .A1(n591bar), .A2(n590bar), .ZN(n599bar);
  OR2_X1 U381 ( .A1(n589), .A2(n588), .ZN(n590) );
  AND2_X1 U381bar ( .A1(n589bar), .A2(n588bar), .ZN(n590bar);
  OR2_X1 U382 ( .A1(in_2), .A2(in_10), .ZN(n588) );
  AND2_X1 U382bar ( .A1(in_2bar), .A2(in_10bar), .ZN(n588bar);
  OR2_X1 U383 ( .A1(in_47), .A2(in_22), .ZN(n589) );
  AND2_X1 U383bar ( .A1(in_47bar), .A2(in_22bar), .ZN(n589bar);
  OR2_X1 U384 ( .A1(n587), .A2(n586), .ZN(n591) );
  AND2_X1 U384bar ( .A1(n587bar), .A2(n586bar), .ZN(n591bar);
  OR2_X1 U385 ( .A1(in_56), .A2(in_54), .ZN(n586) );
  AND2_X1 U385bar ( .A1(in_56bar), .A2(in_54bar), .ZN(n586bar);
  OR2_X1 U386 ( .A1(in_63), .A2(in_61), .ZN(n587) );
  AND2_X1 U386bar ( .A1(in_63bar), .A2(in_61bar), .ZN(n587bar);
  OR2_X1 U387 ( .A1(n585), .A2(n584), .ZN(n820) );
  AND2_X1 U387bar ( .A1(n585bar), .A2(n584bar), .ZN(n820bar);
  OR2_X1 U388 ( .A1(n583), .A2(n582), .ZN(n584) );
  AND2_X1 U388bar ( .A1(n583bar), .A2(n582bar), .ZN(n584bar);
  OR2_X1 U389 ( .A1(n581), .A2(n580), .ZN(n582) );
  AND2_X1 U389bar ( .A1(n581bar), .A2(n580bar), .ZN(n582bar);
  OR2_X1 U390 ( .A1(in[158]), .A2(in[142]), .ZN(n580) );
  AND2_X1 U390bar ( .A1(inbar[158]), .A2(inbar[142]), .ZN(n580bar);
  OR2_X1 U391 ( .A1(in[175]), .A2(in[164]), .ZN(n581) );
  AND2_X1 U391bar ( .A1(inbar[175]), .A2(inbar[164]), .ZN(n581bar);
  OR2_X1 U392 ( .A1(n579), .A2(n578), .ZN(n583) );
  AND2_X1 U392bar ( .A1(n579bar), .A2(n578bar), .ZN(n583bar);
  OR2_X1 U393 ( .A1(in[228]), .A2(in[204]), .ZN(n578) );
  AND2_X1 U393bar ( .A1(inbar[228]), .A2(inbar[204]), .ZN(n578bar);
  OR2_X1 U394 ( .A1(in[91]), .A2(in[87]), .ZN(n579) );
  AND2_X1 U394bar ( .A1(inbar[91]), .A2(inbar[87]), .ZN(n579bar);
  OR2_X1 U395 ( .A1(n577), .A2(n576), .ZN(n585) );
  AND2_X1 U395bar ( .A1(n577bar), .A2(n576bar), .ZN(n585bar);
  OR2_X1 U396 ( .A1(n575), .A2(n574), .ZN(n576) );
  AND2_X1 U396bar ( .A1(n575bar), .A2(n574bar), .ZN(n576bar);
  OR2_X1 U397 ( .A1(in_21), .A2(in_11), .ZN(n574) );
  AND2_X1 U397bar ( .A1(in_21bar), .A2(in_11bar), .ZN(n574bar);
  OR2_X1 U398 ( .A1(in_5), .A2(in_3), .ZN(n575) );
  AND2_X1 U398bar ( .A1(in_5bar), .A2(in_3bar), .ZN(n575bar);
  OR2_X1 U399 ( .A1(n573), .A2(n572), .ZN(n577) );
  AND2_X1 U399bar ( .A1(n573bar), .A2(n572bar), .ZN(n577bar);
  OR2_X1 U400 ( .A1(in_68), .A2(in_64), .ZN(n572) );
  AND2_X1 U400bar ( .A1(in_68bar), .A2(in_64bar), .ZN(n572bar);
  OR2_X1 U401 ( .A1(in_76), .A2(in_73), .ZN(n573) );
  AND2_X1 U401bar ( .A1(in_76bar), .A2(in_73bar), .ZN(n573bar);
  OR2_X1 U402 ( .A1(n778), .A2(n571), .ZN(n601) );
  AND2_X1 U402bar ( .A1(n778bar), .A2(n571bar), .ZN(n601bar);
  OR2_X1 U403 ( .A1(in[100]), .A2(n965), .ZN(n571) );
  AND2_X1 U403bar ( .A1(inbar[100]), .A2(n965bar), .ZN(n571bar);
  OR2_X1 U404 ( .A1(n570), .A2(n569), .ZN(n965) );
  AND2_X1 U404bar ( .A1(n570bar), .A2(n569bar), .ZN(n965bar);
  OR2_X1 U405 ( .A1(n568), .A2(n567), .ZN(n569) );
  AND2_X1 U405bar ( .A1(n568bar), .A2(n567bar), .ZN(n569bar);
  OR2_X1 U406 ( .A1(n566), .A2(n565), .ZN(n567) );
  AND2_X1 U406bar ( .A1(n566bar), .A2(n565bar), .ZN(n567bar);
  OR2_X1 U407 ( .A1(n817), .A2(n750), .ZN(n565) );
  AND2_X1 U407bar ( .A1(n817bar), .A2(n750bar), .ZN(n565bar);
  OR2_X1 U408 ( .A1(n564), .A2(n563), .ZN(n750) );
  AND2_X1 U408bar ( .A1(n564bar), .A2(n563bar), .ZN(n750bar);
  OR2_X1 U409 ( .A1(n562), .A2(n561), .ZN(n563) );
  AND2_X1 U409bar ( .A1(n562bar), .A2(n561bar), .ZN(n563bar);
  OR2_X1 U410 ( .A1(n560), .A2(n559), .ZN(n561) );
  AND2_X1 U410bar ( .A1(n560bar), .A2(n559bar), .ZN(n561bar);
  OR2_X1 U411 ( .A1(in[119]), .A2(in[103]), .ZN(n559) );
  AND2_X1 U411bar ( .A1(inbar[119]), .A2(inbar[103]), .ZN(n559bar);
  OR2_X1 U412 ( .A1(in[137]), .A2(in[133]), .ZN(n560) );
  AND2_X1 U412bar ( .A1(inbar[137]), .A2(inbar[133]), .ZN(n560bar);
  OR2_X1 U413 ( .A1(n558), .A2(n557), .ZN(n562) );
  AND2_X1 U413bar ( .A1(n558bar), .A2(n557bar), .ZN(n562bar);
  OR2_X1 U414 ( .A1(in[176]), .A2(in[173]), .ZN(n557) );
  AND2_X1 U414bar ( .A1(inbar[176]), .A2(inbar[173]), .ZN(n557bar);
  OR2_X1 U415 ( .A1(in[210]), .A2(in[181]), .ZN(n558) );
  AND2_X1 U415bar ( .A1(inbar[210]), .A2(inbar[181]), .ZN(n558bar);
  OR2_X1 U416 ( .A1(n556), .A2(n555), .ZN(n564) );
  AND2_X1 U416bar ( .A1(n556bar), .A2(n555bar), .ZN(n564bar);
  OR2_X1 U417 ( .A1(n554), .A2(n553), .ZN(n555) );
  AND2_X1 U417bar ( .A1(n554bar), .A2(n553bar), .ZN(n555bar);
  OR2_X1 U418 ( .A1(in_13), .A2(in[234]), .ZN(n553) );
  AND2_X1 U418bar ( .A1(in_13bar), .A2(inbar[234]), .ZN(n553bar);
  OR2_X1 U419 ( .A1(in_38), .A2(in_32), .ZN(n554) );
  AND2_X1 U419bar ( .A1(in_38bar), .A2(in_32bar), .ZN(n554bar);
  OR2_X1 U420 ( .A1(n552), .A2(n551), .ZN(n556) );
  AND2_X1 U420bar ( .A1(n552bar), .A2(n551bar), .ZN(n556bar);
  OR2_X1 U421 ( .A1(in_42), .A2(in_41), .ZN(n551) );
  AND2_X1 U421bar ( .A1(in_42bar), .A2(in_41bar), .ZN(n551bar);
  OR2_X1 U422 ( .A1(in_7), .A2(in_49), .ZN(n552) );
  AND2_X1 U422bar ( .A1(in_7bar), .A2(in_49bar), .ZN(n552bar);
  OR2_X1 U423 ( .A1(n550), .A2(n549), .ZN(n817) );
  AND2_X1 U423bar ( .A1(n550bar), .A2(n549bar), .ZN(n817bar);
  OR2_X1 U424 ( .A1(n548), .A2(n547), .ZN(n549) );
  AND2_X1 U424bar ( .A1(n548bar), .A2(n547bar), .ZN(n549bar);
  OR2_X1 U425 ( .A1(n546), .A2(n545), .ZN(n547) );
  AND2_X1 U425bar ( .A1(n546bar), .A2(n545bar), .ZN(n547bar);
  OR2_X1 U426 ( .A1(in[159]), .A2(in[105]), .ZN(n545) );
  AND2_X1 U426bar ( .A1(inbar[159]), .A2(inbar[105]), .ZN(n545bar);
  OR2_X1 U427 ( .A1(in[206]), .A2(in[183]), .ZN(n546) );
  AND2_X1 U427bar ( .A1(inbar[206]), .A2(inbar[183]), .ZN(n546bar);
  OR2_X1 U428 ( .A1(n544), .A2(n543), .ZN(n548) );
  AND2_X1 U428bar ( .A1(n544bar), .A2(n543bar), .ZN(n548bar);
  OR2_X1 U429 ( .A1(in[229]), .A2(in[219]), .ZN(n543) );
  AND2_X1 U429bar ( .A1(inbar[229]), .A2(inbar[219]), .ZN(n543bar);
  OR2_X1 U430 ( .A1(in[235]), .A2(in[232]), .ZN(n544) );
  AND2_X1 U430bar ( .A1(inbar[235]), .A2(inbar[232]), .ZN(n544bar);
  OR2_X1 U431 ( .A1(n542), .A2(n541), .ZN(n550) );
  AND2_X1 U431bar ( .A1(n542bar), .A2(n541bar), .ZN(n550bar);
  OR2_X1 U432 ( .A1(n540), .A2(n539), .ZN(n541) );
  AND2_X1 U432bar ( .A1(n540bar), .A2(n539bar), .ZN(n541bar);
  OR2_X1 U433 ( .A1(in[249]), .A2(in[242]), .ZN(n539) );
  AND2_X1 U433bar ( .A1(inbar[249]), .A2(inbar[242]), .ZN(n539bar);
  OR2_X1 U434 ( .A1(in[89]), .A2(in[254]), .ZN(n540) );
  AND2_X1 U434bar ( .A1(inbar[89]), .A2(inbar[254]), .ZN(n540bar);
  OR2_X1 U435 ( .A1(n538), .A2(n537), .ZN(n542) );
  AND2_X1 U435bar ( .A1(n538bar), .A2(n537bar), .ZN(n542bar);
  OR2_X1 U436 ( .A1(in_14), .A2(in[99]), .ZN(n537) );
  AND2_X1 U436bar ( .A1(in_14bar), .A2(inbar[99]), .ZN(n537bar);
  OR2_X1 U437 ( .A1(in_60), .A2(in_18), .ZN(n538) );
  AND2_X1 U437bar ( .A1(in_60bar), .A2(in_18bar), .ZN(n538bar);
  OR2_X1 U438 ( .A1(in[113]), .A2(n763), .ZN(n566) );
  AND2_X1 U438bar ( .A1(inbar[113]), .A2(n763bar), .ZN(n566bar);
  OR2_X1 U439 ( .A1(n536), .A2(n535), .ZN(n763) );
  AND2_X1 U439bar ( .A1(n536bar), .A2(n535bar), .ZN(n763bar);
  OR2_X1 U440 ( .A1(n534), .A2(n533), .ZN(n535) );
  AND2_X1 U440bar ( .A1(n534bar), .A2(n533bar), .ZN(n535bar);
  OR2_X1 U441 ( .A1(n532), .A2(n531), .ZN(n533) );
  AND2_X1 U441bar ( .A1(n532bar), .A2(n531bar), .ZN(n533bar);
  OR2_X1 U442 ( .A1(in[115]), .A2(in[110]), .ZN(n531) );
  AND2_X1 U442bar ( .A1(inbar[115]), .A2(inbar[110]), .ZN(n531bar);
  OR2_X1 U443 ( .A1(in[125]), .A2(in[117]), .ZN(n532) );
  AND2_X1 U443bar ( .A1(inbar[125]), .A2(inbar[117]), .ZN(n532bar);
  OR2_X1 U444 ( .A1(n530), .A2(n529), .ZN(n534) );
  AND2_X1 U444bar ( .A1(n530bar), .A2(n529bar), .ZN(n534bar);
  OR2_X1 U445 ( .A1(in[180]), .A2(in[128]), .ZN(n529) );
  AND2_X1 U445bar ( .A1(inbar[180]), .A2(inbar[128]), .ZN(n529bar);
  OR2_X1 U446 ( .A1(in[205]), .A2(in[201]), .ZN(n530) );
  AND2_X1 U446bar ( .A1(inbar[205]), .A2(inbar[201]), .ZN(n530bar);
  OR2_X1 U447 ( .A1(n528), .A2(n527), .ZN(n536) );
  AND2_X1 U447bar ( .A1(n528bar), .A2(n527bar), .ZN(n536bar);
  OR2_X1 U448 ( .A1(n526), .A2(n525), .ZN(n527) );
  AND2_X1 U448bar ( .A1(n526bar), .A2(n525bar), .ZN(n527bar);
  OR2_X1 U449 ( .A1(in[244]), .A2(in[239]), .ZN(n525) );
  AND2_X1 U449bar ( .A1(inbar[244]), .A2(inbar[239]), .ZN(n525bar);
  OR2_X1 U450 ( .A1(in[95]), .A2(in[83]), .ZN(n526) );
  AND2_X1 U450bar ( .A1(inbar[95]), .A2(inbar[83]), .ZN(n526bar);
  OR2_X1 U451 ( .A1(n524), .A2(n523), .ZN(n528) );
  AND2_X1 U451bar ( .A1(n524bar), .A2(n523bar), .ZN(n528bar);
  OR2_X1 U452 ( .A1(in_24), .A2(in[97]), .ZN(n523) );
  AND2_X1 U452bar ( .A1(in_24bar), .A2(inbar[97]), .ZN(n523bar);
  OR2_X1 U453 ( .A1(in_33), .A2(in_27), .ZN(n524) );
  AND2_X1 U453bar ( .A1(in_33bar), .A2(in_27bar), .ZN(n524bar);
  OR2_X1 U454 ( .A1(n522), .A2(n521), .ZN(n568) );
  AND2_X1 U454bar ( .A1(n522bar), .A2(n521bar), .ZN(n568bar);
  OR2_X1 U455 ( .A1(in[145]), .A2(in[126]), .ZN(n521) );
  AND2_X1 U455bar ( .A1(inbar[145]), .A2(inbar[126]), .ZN(n521bar);
  OR2_X1 U456 ( .A1(in[169]), .A2(n520), .ZN(n522) );
  AND2_X1 U456bar ( .A1(inbar[169]), .A2(n520bar), .ZN(n522bar);
  OR2_X1 U457 ( .A1(in[221]), .A2(in[172]), .ZN(n520) );
  AND2_X1 U457bar ( .A1(inbar[221]), .A2(inbar[172]), .ZN(n520bar);
  OR2_X1 U458 ( .A1(n519), .A2(n518), .ZN(n570) );
  AND2_X1 U458bar ( .A1(n519bar), .A2(n518bar), .ZN(n570bar);
  OR2_X1 U459 ( .A1(n517), .A2(n516), .ZN(n518) );
  AND2_X1 U459bar ( .A1(n517bar), .A2(n516bar), .ZN(n518bar);
  OR2_X1 U460 ( .A1(in[241]), .A2(in[224]), .ZN(n516) );
  AND2_X1 U460bar ( .A1(inbar[241]), .A2(inbar[224]), .ZN(n516bar);
  OR2_X1 U461 ( .A1(in[86]), .A2(n515), .ZN(n517) );
  AND2_X1 U461bar ( .A1(inbar[86]), .A2(n515bar), .ZN(n517bar);
  OR2_X1 U462 ( .A1(in_43), .A2(in_34), .ZN(n515) );
  AND2_X1 U462bar ( .A1(in_43bar), .A2(in_34bar), .ZN(n515bar);
  OR2_X1 U463 ( .A1(n514), .A2(n513), .ZN(n519) );
  AND2_X1 U463bar ( .A1(n514bar), .A2(n513bar), .ZN(n519bar);
  OR2_X1 U464 ( .A1(in_65), .A2(in_51), .ZN(n513) );
  AND2_X1 U464bar ( .A1(in_65bar), .A2(in_51bar), .ZN(n513bar);
  OR2_X1 U465 ( .A1(in_75), .A2(n512), .ZN(n514) );
  AND2_X1 U465bar ( .A1(in_75bar), .A2(n512bar), .ZN(n514bar);
  OR2_X1 U466 ( .A1(in_81), .A2(in_77), .ZN(n512) );
  AND2_X1 U466bar ( .A1(in_81bar), .A2(in_77bar), .ZN(n512bar);
  OR2_X1 U467 ( .A1(n511), .A2(n510), .ZN(n778) );
  AND2_X1 U467bar ( .A1(n511bar), .A2(n510bar), .ZN(n778bar);
  OR2_X1 U468 ( .A1(n509), .A2(n508), .ZN(n510) );
  AND2_X1 U468bar ( .A1(n509bar), .A2(n508bar), .ZN(n510bar);
  OR2_X1 U469 ( .A1(n507), .A2(n506), .ZN(n508) );
  AND2_X1 U469bar ( .A1(n507bar), .A2(n506bar), .ZN(n508bar);
  OR2_X1 U470 ( .A1(in[107]), .A2(in[101]), .ZN(n506) );
  AND2_X1 U470bar ( .A1(inbar[107]), .A2(inbar[101]), .ZN(n506bar);
  OR2_X1 U471 ( .A1(in[139]), .A2(in[132]), .ZN(n507) );
  AND2_X1 U471bar ( .A1(inbar[139]), .A2(inbar[132]), .ZN(n507bar);
  OR2_X1 U472 ( .A1(n505), .A2(n504), .ZN(n509) );
  AND2_X1 U472bar ( .A1(n505bar), .A2(n504bar), .ZN(n509bar);
  OR2_X1 U473 ( .A1(in[146]), .A2(in[141]), .ZN(n504) );
  AND2_X1 U473bar ( .A1(inbar[146]), .A2(inbar[141]), .ZN(n504bar);
  OR2_X1 U474 ( .A1(in[203]), .A2(in[179]), .ZN(n505) );
  AND2_X1 U474bar ( .A1(inbar[203]), .A2(inbar[179]), .ZN(n505bar);
  OR2_X1 U475 ( .A1(n503), .A2(n502), .ZN(n511) );
  AND2_X1 U475bar ( .A1(n503bar), .A2(n502bar), .ZN(n511bar);
  OR2_X1 U476 ( .A1(n501), .A2(n500), .ZN(n502) );
  AND2_X1 U476bar ( .A1(n501bar), .A2(n500bar), .ZN(n502bar);
  OR2_X1 U477 ( .A1(in[243]), .A2(in[222]), .ZN(n500) );
  AND2_X1 U477bar ( .A1(inbar[243]), .A2(inbar[222]), .ZN(n500bar);
  OR2_X1 U478 ( .A1(in[251]), .A2(in[250]), .ZN(n501) );
  AND2_X1 U478bar ( .A1(inbar[251]), .A2(inbar[250]), .ZN(n501bar);
  OR2_X1 U479 ( .A1(n499), .A2(n498), .ZN(n503) );
  AND2_X1 U479bar ( .A1(n499bar), .A2(n498bar), .ZN(n503bar);
  OR2_X1 U480 ( .A1(in_37), .A2(in_19), .ZN(n498) );
  AND2_X1 U480bar ( .A1(in_37bar), .A2(in_19bar), .ZN(n498bar);
  OR2_X1 U481 ( .A1(in_78), .A2(in_6), .ZN(n499) );
  AND2_X1 U481bar ( .A1(in_78bar), .A2(in_6bar), .ZN(n499bar);
  OR2_X1 U482 ( .A1(n497), .A2(n496), .ZN(n603) );
  AND2_X1 U482bar ( .A1(n497bar), .A2(n496bar), .ZN(n603bar);
  OR2_X1 U483 ( .A1(in[112]), .A2(in[102]), .ZN(n496) );
  AND2_X1 U483bar ( .A1(inbar[112]), .A2(inbar[102]), .ZN(n496bar);
  OR2_X1 U484 ( .A1(in[123]), .A2(n495), .ZN(n497) );
  AND2_X1 U484bar ( .A1(inbar[123]), .A2(n495bar), .ZN(n497bar);
  OR2_X1 U485 ( .A1(in[143]), .A2(in[130]), .ZN(n495) );
  AND2_X1 U485bar ( .A1(inbar[143]), .A2(inbar[130]), .ZN(n495bar);
  OR2_X1 U486 ( .A1(n494), .A2(n493), .ZN(n605) );
  AND2_X1 U486bar ( .A1(n494bar), .A2(n493bar), .ZN(n605bar);
  OR2_X1 U487 ( .A1(n492), .A2(n491), .ZN(n493) );
  AND2_X1 U487bar ( .A1(n492bar), .A2(n491bar), .ZN(n493bar);
  OR2_X1 U488 ( .A1(in[216]), .A2(in[213]), .ZN(n491) );
  AND2_X1 U488bar ( .A1(inbar[216]), .A2(inbar[213]), .ZN(n491bar);
  OR2_X1 U489 ( .A1(in[227]), .A2(n490), .ZN(n492) );
  AND2_X1 U489bar ( .A1(inbar[227]), .A2(n490bar), .ZN(n492bar);
  OR2_X1 U490 ( .A1(in_0), .A2(in[248]), .ZN(n490) );
  AND2_X1 U490bar ( .A1(in_0bar), .A2(inbar[248]), .ZN(n490bar);
  OR2_X1 U491 ( .A1(n489), .A2(n488), .ZN(n494) );
  AND2_X1 U491bar ( .A1(n489bar), .A2(n488bar), .ZN(n494bar);
  OR2_X1 U492 ( .A1(in_46), .A2(in_44), .ZN(n488) );
  AND2_X1 U492bar ( .A1(in_46bar), .A2(in_44bar), .ZN(n488bar);
  OR2_X1 U493 ( .A1(in_50), .A2(n487), .ZN(n489) );
  AND2_X1 U493bar ( .A1(in_50bar), .A2(n487bar), .ZN(n489bar);
  OR2_X1 U494 ( .A1(in_9), .A2(in_80), .ZN(n487) );
  AND2_X1 U494bar ( .A1(in_9bar), .A2(in_80bar), .ZN(n487bar);
endmodule




module sBox_3 ( in, out );
  input [7:0] in;
  //input_done

  output [7:0] out;
  //output_done

  wire   [255:0] decodeOut;
  //wire_done

  decode_3 dec ( .in(in), .out(decodeOut) );
  encode_3 enc ( .in(decodeOut), .out(out) );
endmodule


module CD2_13 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_14 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_15 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_16 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD4_7 ( a, b, y );
  input [3:0] a;
  input [3:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  //input_done

  output [15:0] y;
  reg [15:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]);
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]);
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]);
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]);
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]);
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]);
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]);
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]);
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]);
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]);
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]);
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]);
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]);
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]);
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]);
endmodule




module CD4_8 ( a, b, y );
  input [3:0] a;
  input [3:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  //input_done

  output [15:0] y;
  reg [15:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]);
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]);
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]);
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]);
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]);
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]);
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]);
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]);
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]);
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]);
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]);
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]);
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]);
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]);
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]);
endmodule




module CD16_4 ( a, b, y );
  input [15:0] a;
  input [15:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign abar[8] = ~a[8];
  assign abar[9] = ~a[9];
  assign abar[10] = ~a[10];
  assign abar[11] = ~a[11];
  assign abar[12] = ~a[12];
  assign abar[13] = ~a[13];
  assign abar[14] = ~a[14];
  assign abar[15] = ~a[15];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign bbar[8] = ~b[8];
  assign bbar[9] = ~b[9];
  assign bbar[10] = ~b[10];
  assign bbar[11] = ~b[11];
  assign bbar[12] = ~b[12];
  assign bbar[13] = ~b[13];
  assign bbar[14] = ~b[14];
  assign bbar[15] = ~b[15];
  //input_done

  output [255:0] y;
  reg [255:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[9]), .A2(a[0]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[9]), .A2(abar[0]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[3]), .A2(a[6]), .ZN(y[99]) );
  OR2_X1 U2bar ( .A1(bbar[3]), .A2(abar[6]), .ZN(ybar[99]);
  AND2_X1 U3 ( .A1(b[2]), .A2(a[6]), .ZN(y[98]) );
  OR2_X1 U3bar ( .A1(bbar[2]), .A2(abar[6]), .ZN(ybar[98]);
  AND2_X1 U4 ( .A1(b[1]), .A2(a[6]), .ZN(y[97]) );
  OR2_X1 U4bar ( .A1(bbar[1]), .A2(abar[6]), .ZN(ybar[97]);
  AND2_X1 U5 ( .A1(b[0]), .A2(a[6]), .ZN(y[96]) );
  OR2_X1 U5bar ( .A1(bbar[0]), .A2(abar[6]), .ZN(ybar[96]);
  AND2_X1 U6 ( .A1(b[15]), .A2(a[5]), .ZN(y[95]) );
  OR2_X1 U6bar ( .A1(bbar[15]), .A2(abar[5]), .ZN(ybar[95]);
  AND2_X1 U7 ( .A1(b[14]), .A2(a[5]), .ZN(y[94]) );
  OR2_X1 U7bar ( .A1(bbar[14]), .A2(abar[5]), .ZN(ybar[94]);
  AND2_X1 U8 ( .A1(b[13]), .A2(a[5]), .ZN(y[93]) );
  OR2_X1 U8bar ( .A1(bbar[13]), .A2(abar[5]), .ZN(ybar[93]);
  AND2_X1 U9 ( .A1(b[12]), .A2(a[5]), .ZN(y[92]) );
  OR2_X1 U9bar ( .A1(bbar[12]), .A2(abar[5]), .ZN(ybar[92]);
  AND2_X1 U10 ( .A1(b[11]), .A2(a[5]), .ZN(y[91]) );
  OR2_X1 U10bar ( .A1(bbar[11]), .A2(abar[5]), .ZN(ybar[91]);
  AND2_X1 U11 ( .A1(b[10]), .A2(a[5]), .ZN(y[90]) );
  OR2_X1 U11bar ( .A1(bbar[10]), .A2(abar[5]), .ZN(ybar[90]);
  AND2_X1 U12 ( .A1(b[8]), .A2(a[0]), .ZN(y[8]) );
  OR2_X1 U12bar ( .A1(bbar[8]), .A2(abar[0]), .ZN(ybar[8]);
  AND2_X1 U13 ( .A1(a[5]), .A2(b[9]), .ZN(y[89]) );
  OR2_X1 U13bar ( .A1(abar[5]), .A2(bbar[9]), .ZN(ybar[89]);
  AND2_X1 U14 ( .A1(b[8]), .A2(a[5]), .ZN(y[88]) );
  OR2_X1 U14bar ( .A1(bbar[8]), .A2(abar[5]), .ZN(ybar[88]);
  AND2_X1 U15 ( .A1(b[7]), .A2(a[5]), .ZN(y[87]) );
  OR2_X1 U15bar ( .A1(bbar[7]), .A2(abar[5]), .ZN(ybar[87]);
  AND2_X1 U16 ( .A1(b[6]), .A2(a[5]), .ZN(y[86]) );
  OR2_X1 U16bar ( .A1(bbar[6]), .A2(abar[5]), .ZN(ybar[86]);
  AND2_X1 U17 ( .A1(b[5]), .A2(a[5]), .ZN(y[85]) );
  OR2_X1 U17bar ( .A1(bbar[5]), .A2(abar[5]), .ZN(ybar[85]);
  AND2_X1 U18 ( .A1(b[4]), .A2(a[5]), .ZN(y[84]) );
  OR2_X1 U18bar ( .A1(bbar[4]), .A2(abar[5]), .ZN(ybar[84]);
  AND2_X1 U19 ( .A1(a[5]), .A2(b[3]), .ZN(y[83]) );
  OR2_X1 U19bar ( .A1(abar[5]), .A2(bbar[3]), .ZN(ybar[83]);
  AND2_X1 U20 ( .A1(a[5]), .A2(b[2]), .ZN(y[82]) );
  OR2_X1 U20bar ( .A1(abar[5]), .A2(bbar[2]), .ZN(ybar[82]);
  AND2_X1 U21 ( .A1(a[5]), .A2(b[1]), .ZN(y[81]) );
  OR2_X1 U21bar ( .A1(abar[5]), .A2(bbar[1]), .ZN(ybar[81]);
  AND2_X1 U22 ( .A1(a[5]), .A2(b[0]), .ZN(y[80]) );
  OR2_X1 U22bar ( .A1(abar[5]), .A2(bbar[0]), .ZN(ybar[80]);
  AND2_X1 U23 ( .A1(b[7]), .A2(a[0]), .ZN(y[7]) );
  OR2_X1 U23bar ( .A1(bbar[7]), .A2(abar[0]), .ZN(ybar[7]);
  AND2_X1 U24 ( .A1(a[4]), .A2(b[15]), .ZN(y[79]) );
  OR2_X1 U24bar ( .A1(abar[4]), .A2(bbar[15]), .ZN(ybar[79]);
  AND2_X1 U25 ( .A1(a[4]), .A2(b[14]), .ZN(y[78]) );
  OR2_X1 U25bar ( .A1(abar[4]), .A2(bbar[14]), .ZN(ybar[78]);
  AND2_X1 U26 ( .A1(a[4]), .A2(b[13]), .ZN(y[77]) );
  OR2_X1 U26bar ( .A1(abar[4]), .A2(bbar[13]), .ZN(ybar[77]);
  AND2_X1 U27 ( .A1(a[4]), .A2(b[12]), .ZN(y[76]) );
  OR2_X1 U27bar ( .A1(abar[4]), .A2(bbar[12]), .ZN(ybar[76]);
  AND2_X1 U28 ( .A1(a[4]), .A2(b[11]), .ZN(y[75]) );
  OR2_X1 U28bar ( .A1(abar[4]), .A2(bbar[11]), .ZN(ybar[75]);
  AND2_X1 U29 ( .A1(a[4]), .A2(b[10]), .ZN(y[74]) );
  OR2_X1 U29bar ( .A1(abar[4]), .A2(bbar[10]), .ZN(ybar[74]);
  AND2_X1 U30 ( .A1(a[4]), .A2(b[9]), .ZN(y[73]) );
  OR2_X1 U30bar ( .A1(abar[4]), .A2(bbar[9]), .ZN(ybar[73]);
  AND2_X1 U31 ( .A1(a[4]), .A2(b[8]), .ZN(y[72]) );
  OR2_X1 U31bar ( .A1(abar[4]), .A2(bbar[8]), .ZN(ybar[72]);
  AND2_X1 U32 ( .A1(a[4]), .A2(b[7]), .ZN(y[71]) );
  OR2_X1 U32bar ( .A1(abar[4]), .A2(bbar[7]), .ZN(ybar[71]);
  AND2_X1 U33 ( .A1(a[4]), .A2(b[6]), .ZN(y[70]) );
  OR2_X1 U33bar ( .A1(abar[4]), .A2(bbar[6]), .ZN(ybar[70]);
  AND2_X1 U34 ( .A1(b[6]), .A2(a[0]), .ZN(y[6]) );
  OR2_X1 U34bar ( .A1(bbar[6]), .A2(abar[0]), .ZN(ybar[6]);
  AND2_X1 U35 ( .A1(a[4]), .A2(b[5]), .ZN(y[69]) );
  OR2_X1 U35bar ( .A1(abar[4]), .A2(bbar[5]), .ZN(ybar[69]);
  AND2_X1 U36 ( .A1(a[4]), .A2(b[4]), .ZN(y[68]) );
  OR2_X1 U36bar ( .A1(abar[4]), .A2(bbar[4]), .ZN(ybar[68]);
  AND2_X1 U37 ( .A1(a[4]), .A2(b[3]), .ZN(y[67]) );
  OR2_X1 U37bar ( .A1(abar[4]), .A2(bbar[3]), .ZN(ybar[67]);
  AND2_X1 U38 ( .A1(a[4]), .A2(b[2]), .ZN(y[66]) );
  OR2_X1 U38bar ( .A1(abar[4]), .A2(bbar[2]), .ZN(ybar[66]);
  AND2_X1 U39 ( .A1(a[4]), .A2(b[1]), .ZN(y[65]) );
  OR2_X1 U39bar ( .A1(abar[4]), .A2(bbar[1]), .ZN(ybar[65]);
  AND2_X1 U40 ( .A1(a[4]), .A2(b[0]), .ZN(y[64]) );
  OR2_X1 U40bar ( .A1(abar[4]), .A2(bbar[0]), .ZN(ybar[64]);
  AND2_X1 U41 ( .A1(a[3]), .A2(b[15]), .ZN(y[63]) );
  OR2_X1 U41bar ( .A1(abar[3]), .A2(bbar[15]), .ZN(ybar[63]);
  AND2_X1 U42 ( .A1(a[3]), .A2(b[14]), .ZN(y[62]) );
  OR2_X1 U42bar ( .A1(abar[3]), .A2(bbar[14]), .ZN(ybar[62]);
  AND2_X1 U43 ( .A1(a[3]), .A2(b[13]), .ZN(y[61]) );
  OR2_X1 U43bar ( .A1(abar[3]), .A2(bbar[13]), .ZN(ybar[61]);
  AND2_X1 U44 ( .A1(a[3]), .A2(b[12]), .ZN(y[60]) );
  OR2_X1 U44bar ( .A1(abar[3]), .A2(bbar[12]), .ZN(ybar[60]);
  AND2_X1 U45 ( .A1(b[5]), .A2(a[0]), .ZN(y[5]) );
  OR2_X1 U45bar ( .A1(bbar[5]), .A2(abar[0]), .ZN(ybar[5]);
  AND2_X1 U46 ( .A1(a[3]), .A2(b[11]), .ZN(y[59]) );
  OR2_X1 U46bar ( .A1(abar[3]), .A2(bbar[11]), .ZN(ybar[59]);
  AND2_X1 U47 ( .A1(a[3]), .A2(b[10]), .ZN(y[58]) );
  OR2_X1 U47bar ( .A1(abar[3]), .A2(bbar[10]), .ZN(ybar[58]);
  AND2_X1 U48 ( .A1(a[3]), .A2(b[9]), .ZN(y[57]) );
  OR2_X1 U48bar ( .A1(abar[3]), .A2(bbar[9]), .ZN(ybar[57]);
  AND2_X1 U49 ( .A1(a[3]), .A2(b[8]), .ZN(y[56]) );
  OR2_X1 U49bar ( .A1(abar[3]), .A2(bbar[8]), .ZN(ybar[56]);
  AND2_X1 U50 ( .A1(a[3]), .A2(b[7]), .ZN(y[55]) );
  OR2_X1 U50bar ( .A1(abar[3]), .A2(bbar[7]), .ZN(ybar[55]);
  AND2_X1 U51 ( .A1(a[3]), .A2(b[6]), .ZN(y[54]) );
  OR2_X1 U51bar ( .A1(abar[3]), .A2(bbar[6]), .ZN(ybar[54]);
  AND2_X1 U52 ( .A1(a[3]), .A2(b[5]), .ZN(y[53]) );
  OR2_X1 U52bar ( .A1(abar[3]), .A2(bbar[5]), .ZN(ybar[53]);
  AND2_X1 U53 ( .A1(a[3]), .A2(b[4]), .ZN(y[52]) );
  OR2_X1 U53bar ( .A1(abar[3]), .A2(bbar[4]), .ZN(ybar[52]);
  AND2_X1 U54 ( .A1(a[3]), .A2(b[3]), .ZN(y[51]) );
  OR2_X1 U54bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[51]);
  AND2_X1 U55 ( .A1(a[3]), .A2(b[2]), .ZN(y[50]) );
  OR2_X1 U55bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[50]);
  AND2_X1 U56 ( .A1(b[4]), .A2(a[0]), .ZN(y[4]) );
  OR2_X1 U56bar ( .A1(bbar[4]), .A2(abar[0]), .ZN(ybar[4]);
  AND2_X1 U57 ( .A1(a[3]), .A2(b[1]), .ZN(y[49]) );
  OR2_X1 U57bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[49]);
  AND2_X1 U58 ( .A1(a[3]), .A2(b[0]), .ZN(y[48]) );
  OR2_X1 U58bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[48]);
  AND2_X1 U59 ( .A1(a[2]), .A2(b[15]), .ZN(y[47]) );
  OR2_X1 U59bar ( .A1(abar[2]), .A2(bbar[15]), .ZN(ybar[47]);
  AND2_X1 U60 ( .A1(a[2]), .A2(b[14]), .ZN(y[46]) );
  OR2_X1 U60bar ( .A1(abar[2]), .A2(bbar[14]), .ZN(ybar[46]);
  AND2_X1 U61 ( .A1(a[2]), .A2(b[13]), .ZN(y[45]) );
  OR2_X1 U61bar ( .A1(abar[2]), .A2(bbar[13]), .ZN(ybar[45]);
  AND2_X1 U62 ( .A1(a[2]), .A2(b[12]), .ZN(y[44]) );
  OR2_X1 U62bar ( .A1(abar[2]), .A2(bbar[12]), .ZN(ybar[44]);
  AND2_X1 U63 ( .A1(a[2]), .A2(b[11]), .ZN(y[43]) );
  OR2_X1 U63bar ( .A1(abar[2]), .A2(bbar[11]), .ZN(ybar[43]);
  AND2_X1 U64 ( .A1(a[2]), .A2(b[10]), .ZN(y[42]) );
  OR2_X1 U64bar ( .A1(abar[2]), .A2(bbar[10]), .ZN(ybar[42]);
  AND2_X1 U65 ( .A1(a[2]), .A2(b[9]), .ZN(y[41]) );
  OR2_X1 U65bar ( .A1(abar[2]), .A2(bbar[9]), .ZN(ybar[41]);
  AND2_X1 U66 ( .A1(a[2]), .A2(b[8]), .ZN(y[40]) );
  OR2_X1 U66bar ( .A1(abar[2]), .A2(bbar[8]), .ZN(ybar[40]);
  AND2_X1 U67 ( .A1(b[3]), .A2(a[0]), .ZN(y[3]) );
  OR2_X1 U67bar ( .A1(bbar[3]), .A2(abar[0]), .ZN(ybar[3]);
  AND2_X1 U68 ( .A1(a[2]), .A2(b[7]), .ZN(y[39]) );
  OR2_X1 U68bar ( .A1(abar[2]), .A2(bbar[7]), .ZN(ybar[39]);
  AND2_X1 U69 ( .A1(a[2]), .A2(b[6]), .ZN(y[38]) );
  OR2_X1 U69bar ( .A1(abar[2]), .A2(bbar[6]), .ZN(ybar[38]);
  AND2_X1 U70 ( .A1(a[2]), .A2(b[5]), .ZN(y[37]) );
  OR2_X1 U70bar ( .A1(abar[2]), .A2(bbar[5]), .ZN(ybar[37]);
  AND2_X1 U71 ( .A1(a[2]), .A2(b[4]), .ZN(y[36]) );
  OR2_X1 U71bar ( .A1(abar[2]), .A2(bbar[4]), .ZN(ybar[36]);
  AND2_X1 U72 ( .A1(a[2]), .A2(b[3]), .ZN(y[35]) );
  OR2_X1 U72bar ( .A1(abar[2]), .A2(bbar[3]), .ZN(ybar[35]);
  AND2_X1 U73 ( .A1(a[2]), .A2(b[2]), .ZN(y[34]) );
  OR2_X1 U73bar ( .A1(abar[2]), .A2(bbar[2]), .ZN(ybar[34]);
  AND2_X1 U74 ( .A1(a[2]), .A2(b[1]), .ZN(y[33]) );
  OR2_X1 U74bar ( .A1(abar[2]), .A2(bbar[1]), .ZN(ybar[33]);
  AND2_X1 U75 ( .A1(a[2]), .A2(b[0]), .ZN(y[32]) );
  OR2_X1 U75bar ( .A1(abar[2]), .A2(bbar[0]), .ZN(ybar[32]);
  AND2_X1 U76 ( .A1(a[1]), .A2(b[15]), .ZN(y[31]) );
  OR2_X1 U76bar ( .A1(abar[1]), .A2(bbar[15]), .ZN(ybar[31]);
  AND2_X1 U77 ( .A1(a[1]), .A2(b[14]), .ZN(y[30]) );
  OR2_X1 U77bar ( .A1(abar[1]), .A2(bbar[14]), .ZN(ybar[30]);
  AND2_X1 U78 ( .A1(b[2]), .A2(a[0]), .ZN(y[2]) );
  OR2_X1 U78bar ( .A1(bbar[2]), .A2(abar[0]), .ZN(ybar[2]);
  AND2_X1 U79 ( .A1(a[1]), .A2(b[13]), .ZN(y[29]) );
  OR2_X1 U79bar ( .A1(abar[1]), .A2(bbar[13]), .ZN(ybar[29]);
  AND2_X1 U80 ( .A1(a[1]), .A2(b[12]), .ZN(y[28]) );
  OR2_X1 U80bar ( .A1(abar[1]), .A2(bbar[12]), .ZN(ybar[28]);
  AND2_X1 U81 ( .A1(a[1]), .A2(b[11]), .ZN(y[27]) );
  OR2_X1 U81bar ( .A1(abar[1]), .A2(bbar[11]), .ZN(ybar[27]);
  AND2_X1 U82 ( .A1(a[1]), .A2(b[10]), .ZN(y[26]) );
  OR2_X1 U82bar ( .A1(abar[1]), .A2(bbar[10]), .ZN(ybar[26]);
  AND2_X1 U83 ( .A1(a[1]), .A2(b[9]), .ZN(y[25]) );
  OR2_X1 U83bar ( .A1(abar[1]), .A2(bbar[9]), .ZN(ybar[25]);
  AND2_X1 U84 ( .A1(a[15]), .A2(b[15]), .ZN(y[255]) );
  OR2_X1 U84bar ( .A1(abar[15]), .A2(bbar[15]), .ZN(ybar[255]);
  AND2_X1 U85 ( .A1(a[15]), .A2(b[14]), .ZN(y[254]) );
  OR2_X1 U85bar ( .A1(abar[15]), .A2(bbar[14]), .ZN(ybar[254]);
  AND2_X1 U86 ( .A1(a[15]), .A2(b[13]), .ZN(y[253]) );
  OR2_X1 U86bar ( .A1(abar[15]), .A2(bbar[13]), .ZN(ybar[253]);
  AND2_X1 U87 ( .A1(a[15]), .A2(b[12]), .ZN(y[252]) );
  OR2_X1 U87bar ( .A1(abar[15]), .A2(bbar[12]), .ZN(ybar[252]);
  AND2_X1 U88 ( .A1(a[15]), .A2(b[11]), .ZN(y[251]) );
  OR2_X1 U88bar ( .A1(abar[15]), .A2(bbar[11]), .ZN(ybar[251]);
  AND2_X1 U89 ( .A1(a[15]), .A2(b[10]), .ZN(y[250]) );
  OR2_X1 U89bar ( .A1(abar[15]), .A2(bbar[10]), .ZN(ybar[250]);
  AND2_X1 U90 ( .A1(a[1]), .A2(b[8]), .ZN(y[24]) );
  OR2_X1 U90bar ( .A1(abar[1]), .A2(bbar[8]), .ZN(ybar[24]);
  AND2_X1 U91 ( .A1(a[15]), .A2(b[9]), .ZN(y[249]) );
  OR2_X1 U91bar ( .A1(abar[15]), .A2(bbar[9]), .ZN(ybar[249]);
  AND2_X1 U92 ( .A1(a[15]), .A2(b[8]), .ZN(y[248]) );
  OR2_X1 U92bar ( .A1(abar[15]), .A2(bbar[8]), .ZN(ybar[248]);
  AND2_X1 U93 ( .A1(a[15]), .A2(b[7]), .ZN(y[247]) );
  OR2_X1 U93bar ( .A1(abar[15]), .A2(bbar[7]), .ZN(ybar[247]);
  AND2_X1 U94 ( .A1(a[15]), .A2(b[6]), .ZN(y[246]) );
  OR2_X1 U94bar ( .A1(abar[15]), .A2(bbar[6]), .ZN(ybar[246]);
  AND2_X1 U95 ( .A1(a[15]), .A2(b[5]), .ZN(y[245]) );
  OR2_X1 U95bar ( .A1(abar[15]), .A2(bbar[5]), .ZN(ybar[245]);
  AND2_X1 U96 ( .A1(a[15]), .A2(b[4]), .ZN(y[244]) );
  OR2_X1 U96bar ( .A1(abar[15]), .A2(bbar[4]), .ZN(ybar[244]);
  AND2_X1 U97 ( .A1(a[15]), .A2(b[3]), .ZN(y[243]) );
  OR2_X1 U97bar ( .A1(abar[15]), .A2(bbar[3]), .ZN(ybar[243]);
  AND2_X1 U98 ( .A1(a[15]), .A2(b[2]), .ZN(y[242]) );
  OR2_X1 U98bar ( .A1(abar[15]), .A2(bbar[2]), .ZN(ybar[242]);
  AND2_X1 U99 ( .A1(a[15]), .A2(b[1]), .ZN(y[241]) );
  OR2_X1 U99bar ( .A1(abar[15]), .A2(bbar[1]), .ZN(ybar[241]);
  AND2_X1 U100 ( .A1(a[15]), .A2(b[0]), .ZN(y[240]) );
  OR2_X1 U100bar ( .A1(abar[15]), .A2(bbar[0]), .ZN(ybar[240]);
  AND2_X1 U101 ( .A1(a[1]), .A2(b[7]), .ZN(y[23]) );
  OR2_X1 U101bar ( .A1(abar[1]), .A2(bbar[7]), .ZN(ybar[23]);
  AND2_X1 U102 ( .A1(a[14]), .A2(b[15]), .ZN(y[239]) );
  OR2_X1 U102bar ( .A1(abar[14]), .A2(bbar[15]), .ZN(ybar[239]);
  AND2_X1 U103 ( .A1(a[14]), .A2(b[14]), .ZN(y[238]) );
  OR2_X1 U103bar ( .A1(abar[14]), .A2(bbar[14]), .ZN(ybar[238]);
  AND2_X1 U104 ( .A1(a[14]), .A2(b[13]), .ZN(y[237]) );
  OR2_X1 U104bar ( .A1(abar[14]), .A2(bbar[13]), .ZN(ybar[237]);
  AND2_X1 U105 ( .A1(a[14]), .A2(b[12]), .ZN(y[236]) );
  OR2_X1 U105bar ( .A1(abar[14]), .A2(bbar[12]), .ZN(ybar[236]);
  AND2_X1 U106 ( .A1(a[14]), .A2(b[11]), .ZN(y[235]) );
  OR2_X1 U106bar ( .A1(abar[14]), .A2(bbar[11]), .ZN(ybar[235]);
  AND2_X1 U107 ( .A1(a[14]), .A2(b[10]), .ZN(y[234]) );
  OR2_X1 U107bar ( .A1(abar[14]), .A2(bbar[10]), .ZN(ybar[234]);
  AND2_X1 U108 ( .A1(a[14]), .A2(b[9]), .ZN(y[233]) );
  OR2_X1 U108bar ( .A1(abar[14]), .A2(bbar[9]), .ZN(ybar[233]);
  AND2_X1 U109 ( .A1(a[14]), .A2(b[8]), .ZN(y[232]) );
  OR2_X1 U109bar ( .A1(abar[14]), .A2(bbar[8]), .ZN(ybar[232]);
  AND2_X1 U110 ( .A1(a[14]), .A2(b[7]), .ZN(y[231]) );
  OR2_X1 U110bar ( .A1(abar[14]), .A2(bbar[7]), .ZN(ybar[231]);
  AND2_X1 U111 ( .A1(a[14]), .A2(b[6]), .ZN(y[230]) );
  OR2_X1 U111bar ( .A1(abar[14]), .A2(bbar[6]), .ZN(ybar[230]);
  AND2_X1 U112 ( .A1(a[1]), .A2(b[6]), .ZN(y[22]) );
  OR2_X1 U112bar ( .A1(abar[1]), .A2(bbar[6]), .ZN(ybar[22]);
  AND2_X1 U113 ( .A1(a[14]), .A2(b[5]), .ZN(y[229]) );
  OR2_X1 U113bar ( .A1(abar[14]), .A2(bbar[5]), .ZN(ybar[229]);
  AND2_X1 U114 ( .A1(a[14]), .A2(b[4]), .ZN(y[228]) );
  OR2_X1 U114bar ( .A1(abar[14]), .A2(bbar[4]), .ZN(ybar[228]);
  AND2_X1 U115 ( .A1(a[14]), .A2(b[3]), .ZN(y[227]) );
  OR2_X1 U115bar ( .A1(abar[14]), .A2(bbar[3]), .ZN(ybar[227]);
  AND2_X1 U116 ( .A1(a[14]), .A2(b[2]), .ZN(y[226]) );
  OR2_X1 U116bar ( .A1(abar[14]), .A2(bbar[2]), .ZN(ybar[226]);
  AND2_X1 U117 ( .A1(a[14]), .A2(b[1]), .ZN(y[225]) );
  OR2_X1 U117bar ( .A1(abar[14]), .A2(bbar[1]), .ZN(ybar[225]);
  AND2_X1 U118 ( .A1(a[14]), .A2(b[0]), .ZN(y[224]) );
  OR2_X1 U118bar ( .A1(abar[14]), .A2(bbar[0]), .ZN(ybar[224]);
  AND2_X1 U119 ( .A1(a[13]), .A2(b[15]), .ZN(y[223]) );
  OR2_X1 U119bar ( .A1(abar[13]), .A2(bbar[15]), .ZN(ybar[223]);
  AND2_X1 U120 ( .A1(a[13]), .A2(b[14]), .ZN(y[222]) );
  OR2_X1 U120bar ( .A1(abar[13]), .A2(bbar[14]), .ZN(ybar[222]);
  AND2_X1 U121 ( .A1(a[13]), .A2(b[13]), .ZN(y[221]) );
  OR2_X1 U121bar ( .A1(abar[13]), .A2(bbar[13]), .ZN(ybar[221]);
  AND2_X1 U122 ( .A1(a[13]), .A2(b[12]), .ZN(y[220]) );
  OR2_X1 U122bar ( .A1(abar[13]), .A2(bbar[12]), .ZN(ybar[220]);
  AND2_X1 U123 ( .A1(a[1]), .A2(b[5]), .ZN(y[21]) );
  OR2_X1 U123bar ( .A1(abar[1]), .A2(bbar[5]), .ZN(ybar[21]);
  AND2_X1 U124 ( .A1(a[13]), .A2(b[11]), .ZN(y[219]) );
  OR2_X1 U124bar ( .A1(abar[13]), .A2(bbar[11]), .ZN(ybar[219]);
  AND2_X1 U125 ( .A1(a[13]), .A2(b[10]), .ZN(y[218]) );
  OR2_X1 U125bar ( .A1(abar[13]), .A2(bbar[10]), .ZN(ybar[218]);
  AND2_X1 U126 ( .A1(a[13]), .A2(b[9]), .ZN(y[217]) );
  OR2_X1 U126bar ( .A1(abar[13]), .A2(bbar[9]), .ZN(ybar[217]);
  AND2_X1 U127 ( .A1(a[13]), .A2(b[8]), .ZN(y[216]) );
  OR2_X1 U127bar ( .A1(abar[13]), .A2(bbar[8]), .ZN(ybar[216]);
  AND2_X1 U128 ( .A1(a[13]), .A2(b[7]), .ZN(y[215]) );
  OR2_X1 U128bar ( .A1(abar[13]), .A2(bbar[7]), .ZN(ybar[215]);
  AND2_X1 U129 ( .A1(a[13]), .A2(b[6]), .ZN(y[214]) );
  OR2_X1 U129bar ( .A1(abar[13]), .A2(bbar[6]), .ZN(ybar[214]);
  AND2_X1 U130 ( .A1(a[13]), .A2(b[5]), .ZN(y[213]) );
  OR2_X1 U130bar ( .A1(abar[13]), .A2(bbar[5]), .ZN(ybar[213]);
  AND2_X1 U131 ( .A1(a[13]), .A2(b[4]), .ZN(y[212]) );
  OR2_X1 U131bar ( .A1(abar[13]), .A2(bbar[4]), .ZN(ybar[212]);
  AND2_X1 U132 ( .A1(a[13]), .A2(b[3]), .ZN(y[211]) );
  OR2_X1 U132bar ( .A1(abar[13]), .A2(bbar[3]), .ZN(ybar[211]);
  AND2_X1 U133 ( .A1(a[13]), .A2(b[2]), .ZN(y[210]) );
  OR2_X1 U133bar ( .A1(abar[13]), .A2(bbar[2]), .ZN(ybar[210]);
  AND2_X1 U134 ( .A1(a[1]), .A2(b[4]), .ZN(y[20]) );
  OR2_X1 U134bar ( .A1(abar[1]), .A2(bbar[4]), .ZN(ybar[20]);
  AND2_X1 U135 ( .A1(a[13]), .A2(b[1]), .ZN(y[209]) );
  OR2_X1 U135bar ( .A1(abar[13]), .A2(bbar[1]), .ZN(ybar[209]);
  AND2_X1 U136 ( .A1(a[13]), .A2(b[0]), .ZN(y[208]) );
  OR2_X1 U136bar ( .A1(abar[13]), .A2(bbar[0]), .ZN(ybar[208]);
  AND2_X1 U137 ( .A1(a[12]), .A2(b[15]), .ZN(y[207]) );
  OR2_X1 U137bar ( .A1(abar[12]), .A2(bbar[15]), .ZN(ybar[207]);
  AND2_X1 U138 ( .A1(a[12]), .A2(b[14]), .ZN(y[206]) );
  OR2_X1 U138bar ( .A1(abar[12]), .A2(bbar[14]), .ZN(ybar[206]);
  AND2_X1 U139 ( .A1(a[12]), .A2(b[13]), .ZN(y[205]) );
  OR2_X1 U139bar ( .A1(abar[12]), .A2(bbar[13]), .ZN(ybar[205]);
  AND2_X1 U140 ( .A1(a[12]), .A2(b[12]), .ZN(y[204]) );
  OR2_X1 U140bar ( .A1(abar[12]), .A2(bbar[12]), .ZN(ybar[204]);
  AND2_X1 U141 ( .A1(a[12]), .A2(b[11]), .ZN(y[203]) );
  OR2_X1 U141bar ( .A1(abar[12]), .A2(bbar[11]), .ZN(ybar[203]);
  AND2_X1 U142 ( .A1(a[12]), .A2(b[10]), .ZN(y[202]) );
  OR2_X1 U142bar ( .A1(abar[12]), .A2(bbar[10]), .ZN(ybar[202]);
  AND2_X1 U143 ( .A1(a[12]), .A2(b[9]), .ZN(y[201]) );
  OR2_X1 U143bar ( .A1(abar[12]), .A2(bbar[9]), .ZN(ybar[201]);
  AND2_X1 U144 ( .A1(a[12]), .A2(b[8]), .ZN(y[200]) );
  OR2_X1 U144bar ( .A1(abar[12]), .A2(bbar[8]), .ZN(ybar[200]);
  AND2_X1 U145 ( .A1(b[1]), .A2(a[0]), .ZN(y[1]) );
  OR2_X1 U145bar ( .A1(bbar[1]), .A2(abar[0]), .ZN(ybar[1]);
  AND2_X1 U146 ( .A1(a[1]), .A2(b[3]), .ZN(y[19]) );
  OR2_X1 U146bar ( .A1(abar[1]), .A2(bbar[3]), .ZN(ybar[19]);
  AND2_X1 U147 ( .A1(a[12]), .A2(b[7]), .ZN(y[199]) );
  OR2_X1 U147bar ( .A1(abar[12]), .A2(bbar[7]), .ZN(ybar[199]);
  AND2_X1 U148 ( .A1(a[12]), .A2(b[6]), .ZN(y[198]) );
  OR2_X1 U148bar ( .A1(abar[12]), .A2(bbar[6]), .ZN(ybar[198]);
  AND2_X1 U149 ( .A1(a[12]), .A2(b[5]), .ZN(y[197]) );
  OR2_X1 U149bar ( .A1(abar[12]), .A2(bbar[5]), .ZN(ybar[197]);
  AND2_X1 U150 ( .A1(a[12]), .A2(b[4]), .ZN(y[196]) );
  OR2_X1 U150bar ( .A1(abar[12]), .A2(bbar[4]), .ZN(ybar[196]);
  AND2_X1 U151 ( .A1(a[12]), .A2(b[3]), .ZN(y[195]) );
  OR2_X1 U151bar ( .A1(abar[12]), .A2(bbar[3]), .ZN(ybar[195]);
  AND2_X1 U152 ( .A1(a[12]), .A2(b[2]), .ZN(y[194]) );
  OR2_X1 U152bar ( .A1(abar[12]), .A2(bbar[2]), .ZN(ybar[194]);
  AND2_X1 U153 ( .A1(a[12]), .A2(b[1]), .ZN(y[193]) );
  OR2_X1 U153bar ( .A1(abar[12]), .A2(bbar[1]), .ZN(ybar[193]);
  AND2_X1 U154 ( .A1(a[12]), .A2(b[0]), .ZN(y[192]) );
  OR2_X1 U154bar ( .A1(abar[12]), .A2(bbar[0]), .ZN(ybar[192]);
  AND2_X1 U155 ( .A1(a[11]), .A2(b[15]), .ZN(y[191]) );
  OR2_X1 U155bar ( .A1(abar[11]), .A2(bbar[15]), .ZN(ybar[191]);
  AND2_X1 U156 ( .A1(a[11]), .A2(b[14]), .ZN(y[190]) );
  OR2_X1 U156bar ( .A1(abar[11]), .A2(bbar[14]), .ZN(ybar[190]);
  AND2_X1 U157 ( .A1(a[1]), .A2(b[2]), .ZN(y[18]) );
  OR2_X1 U157bar ( .A1(abar[1]), .A2(bbar[2]), .ZN(ybar[18]);
  AND2_X1 U158 ( .A1(a[11]), .A2(b[13]), .ZN(y[189]) );
  OR2_X1 U158bar ( .A1(abar[11]), .A2(bbar[13]), .ZN(ybar[189]);
  AND2_X1 U159 ( .A1(a[11]), .A2(b[12]), .ZN(y[188]) );
  OR2_X1 U159bar ( .A1(abar[11]), .A2(bbar[12]), .ZN(ybar[188]);
  AND2_X1 U160 ( .A1(a[11]), .A2(b[11]), .ZN(y[187]) );
  OR2_X1 U160bar ( .A1(abar[11]), .A2(bbar[11]), .ZN(ybar[187]);
  AND2_X1 U161 ( .A1(a[11]), .A2(b[10]), .ZN(y[186]) );
  OR2_X1 U161bar ( .A1(abar[11]), .A2(bbar[10]), .ZN(ybar[186]);
  AND2_X1 U162 ( .A1(a[11]), .A2(b[9]), .ZN(y[185]) );
  OR2_X1 U162bar ( .A1(abar[11]), .A2(bbar[9]), .ZN(ybar[185]);
  AND2_X1 U163 ( .A1(a[11]), .A2(b[8]), .ZN(y[184]) );
  OR2_X1 U163bar ( .A1(abar[11]), .A2(bbar[8]), .ZN(ybar[184]);
  AND2_X1 U164 ( .A1(a[11]), .A2(b[7]), .ZN(y[183]) );
  OR2_X1 U164bar ( .A1(abar[11]), .A2(bbar[7]), .ZN(ybar[183]);
  AND2_X1 U165 ( .A1(a[11]), .A2(b[6]), .ZN(y[182]) );
  OR2_X1 U165bar ( .A1(abar[11]), .A2(bbar[6]), .ZN(ybar[182]);
  AND2_X1 U166 ( .A1(a[11]), .A2(b[5]), .ZN(y[181]) );
  OR2_X1 U166bar ( .A1(abar[11]), .A2(bbar[5]), .ZN(ybar[181]);
  AND2_X1 U167 ( .A1(a[11]), .A2(b[4]), .ZN(y[180]) );
  OR2_X1 U167bar ( .A1(abar[11]), .A2(bbar[4]), .ZN(ybar[180]);
  AND2_X1 U168 ( .A1(a[1]), .A2(b[1]), .ZN(y[17]) );
  OR2_X1 U168bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[17]);
  AND2_X1 U169 ( .A1(a[11]), .A2(b[3]), .ZN(y[179]) );
  OR2_X1 U169bar ( .A1(abar[11]), .A2(bbar[3]), .ZN(ybar[179]);
  AND2_X1 U170 ( .A1(a[11]), .A2(b[2]), .ZN(y[178]) );
  OR2_X1 U170bar ( .A1(abar[11]), .A2(bbar[2]), .ZN(ybar[178]);
  AND2_X1 U171 ( .A1(a[11]), .A2(b[1]), .ZN(y[177]) );
  OR2_X1 U171bar ( .A1(abar[11]), .A2(bbar[1]), .ZN(ybar[177]);
  AND2_X1 U172 ( .A1(a[11]), .A2(b[0]), .ZN(y[176]) );
  OR2_X1 U172bar ( .A1(abar[11]), .A2(bbar[0]), .ZN(ybar[176]);
  AND2_X1 U173 ( .A1(a[10]), .A2(b[15]), .ZN(y[175]) );
  OR2_X1 U173bar ( .A1(abar[10]), .A2(bbar[15]), .ZN(ybar[175]);
  AND2_X1 U174 ( .A1(a[10]), .A2(b[14]), .ZN(y[174]) );
  OR2_X1 U174bar ( .A1(abar[10]), .A2(bbar[14]), .ZN(ybar[174]);
  AND2_X1 U175 ( .A1(a[10]), .A2(b[13]), .ZN(y[173]) );
  OR2_X1 U175bar ( .A1(abar[10]), .A2(bbar[13]), .ZN(ybar[173]);
  AND2_X1 U176 ( .A1(a[10]), .A2(b[12]), .ZN(y[172]) );
  OR2_X1 U176bar ( .A1(abar[10]), .A2(bbar[12]), .ZN(ybar[172]);
  AND2_X1 U177 ( .A1(a[10]), .A2(b[11]), .ZN(y[171]) );
  OR2_X1 U177bar ( .A1(abar[10]), .A2(bbar[11]), .ZN(ybar[171]);
  AND2_X1 U178 ( .A1(a[10]), .A2(b[10]), .ZN(y[170]) );
  OR2_X1 U178bar ( .A1(abar[10]), .A2(bbar[10]), .ZN(ybar[170]);
  AND2_X1 U179 ( .A1(a[1]), .A2(b[0]), .ZN(y[16]) );
  OR2_X1 U179bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[16]);
  AND2_X1 U180 ( .A1(a[10]), .A2(b[9]), .ZN(y[169]) );
  OR2_X1 U180bar ( .A1(abar[10]), .A2(bbar[9]), .ZN(ybar[169]);
  AND2_X1 U181 ( .A1(a[10]), .A2(b[8]), .ZN(y[168]) );
  OR2_X1 U181bar ( .A1(abar[10]), .A2(bbar[8]), .ZN(ybar[168]);
  AND2_X1 U182 ( .A1(a[10]), .A2(b[7]), .ZN(y[167]) );
  OR2_X1 U182bar ( .A1(abar[10]), .A2(bbar[7]), .ZN(ybar[167]);
  AND2_X1 U183 ( .A1(a[10]), .A2(b[6]), .ZN(y[166]) );
  OR2_X1 U183bar ( .A1(abar[10]), .A2(bbar[6]), .ZN(ybar[166]);
  AND2_X1 U184 ( .A1(a[10]), .A2(b[5]), .ZN(y[165]) );
  OR2_X1 U184bar ( .A1(abar[10]), .A2(bbar[5]), .ZN(ybar[165]);
  AND2_X1 U185 ( .A1(a[10]), .A2(b[4]), .ZN(y[164]) );
  OR2_X1 U185bar ( .A1(abar[10]), .A2(bbar[4]), .ZN(ybar[164]);
  AND2_X1 U186 ( .A1(a[10]), .A2(b[3]), .ZN(y[163]) );
  OR2_X1 U186bar ( .A1(abar[10]), .A2(bbar[3]), .ZN(ybar[163]);
  AND2_X1 U187 ( .A1(a[10]), .A2(b[2]), .ZN(y[162]) );
  OR2_X1 U187bar ( .A1(abar[10]), .A2(bbar[2]), .ZN(ybar[162]);
  AND2_X1 U188 ( .A1(a[10]), .A2(b[1]), .ZN(y[161]) );
  OR2_X1 U188bar ( .A1(abar[10]), .A2(bbar[1]), .ZN(ybar[161]);
  AND2_X1 U189 ( .A1(a[10]), .A2(b[0]), .ZN(y[160]) );
  OR2_X1 U189bar ( .A1(abar[10]), .A2(bbar[0]), .ZN(ybar[160]);
  AND2_X1 U190 ( .A1(b[15]), .A2(a[0]), .ZN(y[15]) );
  OR2_X1 U190bar ( .A1(bbar[15]), .A2(abar[0]), .ZN(ybar[15]);
  AND2_X1 U191 ( .A1(a[9]), .A2(b[15]), .ZN(y[159]) );
  OR2_X1 U191bar ( .A1(abar[9]), .A2(bbar[15]), .ZN(ybar[159]);
  AND2_X1 U192 ( .A1(a[9]), .A2(b[14]), .ZN(y[158]) );
  OR2_X1 U192bar ( .A1(abar[9]), .A2(bbar[14]), .ZN(ybar[158]);
  AND2_X1 U193 ( .A1(a[9]), .A2(b[13]), .ZN(y[157]) );
  OR2_X1 U193bar ( .A1(abar[9]), .A2(bbar[13]), .ZN(ybar[157]);
  AND2_X1 U194 ( .A1(a[9]), .A2(b[12]), .ZN(y[156]) );
  OR2_X1 U194bar ( .A1(abar[9]), .A2(bbar[12]), .ZN(ybar[156]);
  AND2_X1 U195 ( .A1(a[9]), .A2(b[11]), .ZN(y[155]) );
  OR2_X1 U195bar ( .A1(abar[9]), .A2(bbar[11]), .ZN(ybar[155]);
  AND2_X1 U196 ( .A1(a[9]), .A2(b[10]), .ZN(y[154]) );
  OR2_X1 U196bar ( .A1(abar[9]), .A2(bbar[10]), .ZN(ybar[154]);
  AND2_X1 U197 ( .A1(a[9]), .A2(b[9]), .ZN(y[153]) );
  OR2_X1 U197bar ( .A1(abar[9]), .A2(bbar[9]), .ZN(ybar[153]);
  AND2_X1 U198 ( .A1(a[9]), .A2(b[8]), .ZN(y[152]) );
  OR2_X1 U198bar ( .A1(abar[9]), .A2(bbar[8]), .ZN(ybar[152]);
  AND2_X1 U199 ( .A1(a[9]), .A2(b[7]), .ZN(y[151]) );
  OR2_X1 U199bar ( .A1(abar[9]), .A2(bbar[7]), .ZN(ybar[151]);
  AND2_X1 U200 ( .A1(a[9]), .A2(b[6]), .ZN(y[150]) );
  OR2_X1 U200bar ( .A1(abar[9]), .A2(bbar[6]), .ZN(ybar[150]);
  AND2_X1 U201 ( .A1(b[14]), .A2(a[0]), .ZN(y[14]) );
  OR2_X1 U201bar ( .A1(bbar[14]), .A2(abar[0]), .ZN(ybar[14]);
  AND2_X1 U202 ( .A1(a[9]), .A2(b[5]), .ZN(y[149]) );
  OR2_X1 U202bar ( .A1(abar[9]), .A2(bbar[5]), .ZN(ybar[149]);
  AND2_X1 U203 ( .A1(a[9]), .A2(b[4]), .ZN(y[148]) );
  OR2_X1 U203bar ( .A1(abar[9]), .A2(bbar[4]), .ZN(ybar[148]);
  AND2_X1 U204 ( .A1(a[9]), .A2(b[3]), .ZN(y[147]) );
  OR2_X1 U204bar ( .A1(abar[9]), .A2(bbar[3]), .ZN(ybar[147]);
  AND2_X1 U205 ( .A1(a[9]), .A2(b[2]), .ZN(y[146]) );
  OR2_X1 U205bar ( .A1(abar[9]), .A2(bbar[2]), .ZN(ybar[146]);
  AND2_X1 U206 ( .A1(a[9]), .A2(b[1]), .ZN(y[145]) );
  OR2_X1 U206bar ( .A1(abar[9]), .A2(bbar[1]), .ZN(ybar[145]);
  AND2_X1 U207 ( .A1(a[9]), .A2(b[0]), .ZN(y[144]) );
  OR2_X1 U207bar ( .A1(abar[9]), .A2(bbar[0]), .ZN(ybar[144]);
  AND2_X1 U208 ( .A1(a[8]), .A2(b[15]), .ZN(y[143]) );
  OR2_X1 U208bar ( .A1(abar[8]), .A2(bbar[15]), .ZN(ybar[143]);
  AND2_X1 U209 ( .A1(a[8]), .A2(b[14]), .ZN(y[142]) );
  OR2_X1 U209bar ( .A1(abar[8]), .A2(bbar[14]), .ZN(ybar[142]);
  AND2_X1 U210 ( .A1(a[8]), .A2(b[13]), .ZN(y[141]) );
  OR2_X1 U210bar ( .A1(abar[8]), .A2(bbar[13]), .ZN(ybar[141]);
  AND2_X1 U211 ( .A1(a[8]), .A2(b[12]), .ZN(y[140]) );
  OR2_X1 U211bar ( .A1(abar[8]), .A2(bbar[12]), .ZN(ybar[140]);
  AND2_X1 U212 ( .A1(b[13]), .A2(a[0]), .ZN(y[13]) );
  OR2_X1 U212bar ( .A1(bbar[13]), .A2(abar[0]), .ZN(ybar[13]);
  AND2_X1 U213 ( .A1(a[8]), .A2(b[11]), .ZN(y[139]) );
  OR2_X1 U213bar ( .A1(abar[8]), .A2(bbar[11]), .ZN(ybar[139]);
  AND2_X1 U214 ( .A1(a[8]), .A2(b[10]), .ZN(y[138]) );
  OR2_X1 U214bar ( .A1(abar[8]), .A2(bbar[10]), .ZN(ybar[138]);
  AND2_X1 U215 ( .A1(a[8]), .A2(b[9]), .ZN(y[137]) );
  OR2_X1 U215bar ( .A1(abar[8]), .A2(bbar[9]), .ZN(ybar[137]);
  AND2_X1 U216 ( .A1(a[8]), .A2(b[8]), .ZN(y[136]) );
  OR2_X1 U216bar ( .A1(abar[8]), .A2(bbar[8]), .ZN(ybar[136]);
  AND2_X1 U217 ( .A1(a[8]), .A2(b[7]), .ZN(y[135]) );
  OR2_X1 U217bar ( .A1(abar[8]), .A2(bbar[7]), .ZN(ybar[135]);
  AND2_X1 U218 ( .A1(a[8]), .A2(b[6]), .ZN(y[134]) );
  OR2_X1 U218bar ( .A1(abar[8]), .A2(bbar[6]), .ZN(ybar[134]);
  AND2_X1 U219 ( .A1(a[8]), .A2(b[5]), .ZN(y[133]) );
  OR2_X1 U219bar ( .A1(abar[8]), .A2(bbar[5]), .ZN(ybar[133]);
  AND2_X1 U220 ( .A1(a[8]), .A2(b[4]), .ZN(y[132]) );
  OR2_X1 U220bar ( .A1(abar[8]), .A2(bbar[4]), .ZN(ybar[132]);
  AND2_X1 U221 ( .A1(a[8]), .A2(b[3]), .ZN(y[131]) );
  OR2_X1 U221bar ( .A1(abar[8]), .A2(bbar[3]), .ZN(ybar[131]);
  AND2_X1 U222 ( .A1(a[8]), .A2(b[2]), .ZN(y[130]) );
  OR2_X1 U222bar ( .A1(abar[8]), .A2(bbar[2]), .ZN(ybar[130]);
  AND2_X1 U223 ( .A1(b[12]), .A2(a[0]), .ZN(y[12]) );
  OR2_X1 U223bar ( .A1(bbar[12]), .A2(abar[0]), .ZN(ybar[12]);
  AND2_X1 U224 ( .A1(a[8]), .A2(b[1]), .ZN(y[129]) );
  OR2_X1 U224bar ( .A1(abar[8]), .A2(bbar[1]), .ZN(ybar[129]);
  AND2_X1 U225 ( .A1(a[8]), .A2(b[0]), .ZN(y[128]) );
  OR2_X1 U225bar ( .A1(abar[8]), .A2(bbar[0]), .ZN(ybar[128]);
  AND2_X1 U226 ( .A1(a[7]), .A2(b[15]), .ZN(y[127]) );
  OR2_X1 U226bar ( .A1(abar[7]), .A2(bbar[15]), .ZN(ybar[127]);
  AND2_X1 U227 ( .A1(a[7]), .A2(b[14]), .ZN(y[126]) );
  OR2_X1 U227bar ( .A1(abar[7]), .A2(bbar[14]), .ZN(ybar[126]);
  AND2_X1 U228 ( .A1(a[7]), .A2(b[13]), .ZN(y[125]) );
  OR2_X1 U228bar ( .A1(abar[7]), .A2(bbar[13]), .ZN(ybar[125]);
  AND2_X1 U229 ( .A1(a[7]), .A2(b[12]), .ZN(y[124]) );
  OR2_X1 U229bar ( .A1(abar[7]), .A2(bbar[12]), .ZN(ybar[124]);
  AND2_X1 U230 ( .A1(a[7]), .A2(b[11]), .ZN(y[123]) );
  OR2_X1 U230bar ( .A1(abar[7]), .A2(bbar[11]), .ZN(ybar[123]);
  AND2_X1 U231 ( .A1(a[7]), .A2(b[10]), .ZN(y[122]) );
  OR2_X1 U231bar ( .A1(abar[7]), .A2(bbar[10]), .ZN(ybar[122]);
  AND2_X1 U232 ( .A1(a[7]), .A2(b[9]), .ZN(y[121]) );
  OR2_X1 U232bar ( .A1(abar[7]), .A2(bbar[9]), .ZN(ybar[121]);
  AND2_X1 U233 ( .A1(a[7]), .A2(b[8]), .ZN(y[120]) );
  OR2_X1 U233bar ( .A1(abar[7]), .A2(bbar[8]), .ZN(ybar[120]);
  AND2_X1 U234 ( .A1(b[11]), .A2(a[0]), .ZN(y[11]) );
  OR2_X1 U234bar ( .A1(bbar[11]), .A2(abar[0]), .ZN(ybar[11]);
  AND2_X1 U235 ( .A1(a[7]), .A2(b[7]), .ZN(y[119]) );
  OR2_X1 U235bar ( .A1(abar[7]), .A2(bbar[7]), .ZN(ybar[119]);
  AND2_X1 U236 ( .A1(a[7]), .A2(b[6]), .ZN(y[118]) );
  OR2_X1 U236bar ( .A1(abar[7]), .A2(bbar[6]), .ZN(ybar[118]);
  AND2_X1 U237 ( .A1(a[7]), .A2(b[5]), .ZN(y[117]) );
  OR2_X1 U237bar ( .A1(abar[7]), .A2(bbar[5]), .ZN(ybar[117]);
  AND2_X1 U238 ( .A1(a[7]), .A2(b[4]), .ZN(y[116]) );
  OR2_X1 U238bar ( .A1(abar[7]), .A2(bbar[4]), .ZN(ybar[116]);
  AND2_X1 U239 ( .A1(a[7]), .A2(b[3]), .ZN(y[115]) );
  OR2_X1 U239bar ( .A1(abar[7]), .A2(bbar[3]), .ZN(ybar[115]);
  AND2_X1 U240 ( .A1(a[7]), .A2(b[2]), .ZN(y[114]) );
  OR2_X1 U240bar ( .A1(abar[7]), .A2(bbar[2]), .ZN(ybar[114]);
  AND2_X1 U241 ( .A1(a[7]), .A2(b[1]), .ZN(y[113]) );
  OR2_X1 U241bar ( .A1(abar[7]), .A2(bbar[1]), .ZN(ybar[113]);
  AND2_X1 U242 ( .A1(a[7]), .A2(b[0]), .ZN(y[112]) );
  OR2_X1 U242bar ( .A1(abar[7]), .A2(bbar[0]), .ZN(ybar[112]);
  AND2_X1 U243 ( .A1(b[15]), .A2(a[6]), .ZN(y[111]) );
  OR2_X1 U243bar ( .A1(bbar[15]), .A2(abar[6]), .ZN(ybar[111]);
  AND2_X1 U244 ( .A1(b[14]), .A2(a[6]), .ZN(y[110]) );
  OR2_X1 U244bar ( .A1(bbar[14]), .A2(abar[6]), .ZN(ybar[110]);
  AND2_X1 U245 ( .A1(b[10]), .A2(a[0]), .ZN(y[10]) );
  OR2_X1 U245bar ( .A1(bbar[10]), .A2(abar[0]), .ZN(ybar[10]);
  AND2_X1 U246 ( .A1(b[13]), .A2(a[6]), .ZN(y[109]) );
  OR2_X1 U246bar ( .A1(bbar[13]), .A2(abar[6]), .ZN(ybar[109]);
  AND2_X1 U247 ( .A1(b[12]), .A2(a[6]), .ZN(y[108]) );
  OR2_X1 U247bar ( .A1(bbar[12]), .A2(abar[6]), .ZN(ybar[108]);
  AND2_X1 U248 ( .A1(b[11]), .A2(a[6]), .ZN(y[107]) );
  OR2_X1 U248bar ( .A1(bbar[11]), .A2(abar[6]), .ZN(ybar[107]);
  AND2_X1 U249 ( .A1(b[10]), .A2(a[6]), .ZN(y[106]) );
  OR2_X1 U249bar ( .A1(bbar[10]), .A2(abar[6]), .ZN(ybar[106]);
  AND2_X1 U250 ( .A1(a[6]), .A2(b[9]), .ZN(y[105]) );
  OR2_X1 U250bar ( .A1(abar[6]), .A2(bbar[9]), .ZN(ybar[105]);
  AND2_X1 U251 ( .A1(b[8]), .A2(a[6]), .ZN(y[104]) );
  OR2_X1 U251bar ( .A1(bbar[8]), .A2(abar[6]), .ZN(ybar[104]);
  AND2_X1 U252 ( .A1(b[7]), .A2(a[6]), .ZN(y[103]) );
  OR2_X1 U252bar ( .A1(bbar[7]), .A2(abar[6]), .ZN(ybar[103]);
  AND2_X1 U253 ( .A1(b[6]), .A2(a[6]), .ZN(y[102]) );
  OR2_X1 U253bar ( .A1(bbar[6]), .A2(abar[6]), .ZN(ybar[102]);
  AND2_X1 U254 ( .A1(b[5]), .A2(a[6]), .ZN(y[101]) );
  OR2_X1 U254bar ( .A1(bbar[5]), .A2(abar[6]), .ZN(ybar[101]);
  AND2_X1 U255 ( .A1(b[4]), .A2(a[6]), .ZN(y[100]) );
  OR2_X1 U255bar ( .A1(bbar[4]), .A2(abar[6]), .ZN(ybar[100]);
  AND2_X1 U256 ( .A1(b[0]), .A2(a[0]), .ZN(y[0]) );
  OR2_X1 U256bar ( .A1(bbar[0]), .A2(abar[0]), .ZN(ybar[0]);
endmodule




module decode_4 ( in, out );
  input [7:0] in;
  //input_done

  output [255:0] out;
  //output_done

  wire   [15:0] level1;
  wire   [31:0] level2;
  //wire_done

  CD2_16 cd_l1_1 ( .a(in[1]), .b(in[0]), .y(level1[3:0]) );
  CD2_15 cd_l1_2 ( .a(in[3]), .b(in[2]), .y(level1[7:4]) );
  CD2_14 cd_l1_3 ( .a(in[5]), .b(in[4]), .y(level1[11:8]) );
  CD2_13 cd_l1_4 ( .a(in[7]), .b(in[6]), .y(level1[15:12]) );
  CD4_8 cd_l2_1 ( .a(level1[7:4]), .b(level1[3:0]), .y(level2[15:0]) );
  CD4_7 cd_l2_2 ( .a(level1[15:12]), .b(level1[11:8]), .y(level2[31:16]) );
  CD16_4 cd_l3 ( .a(level2[31:16]), .b(level2[15:0]), .y(out) );
endmodule


module encode_4 ( in, out );
  input [255:0] in;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
  assign inbar[8] = ~in[8];
  assign inbar[9] = ~in[9];
  assign inbar[10] = ~in[10];
  assign inbar[11] = ~in[11];
  assign inbar[12] = ~in[12];
  assign inbar[13] = ~in[13];
  assign inbar[14] = ~in[14];
  assign inbar[15] = ~in[15];
  assign inbar[16] = ~in[16];
  assign inbar[17] = ~in[17];
  assign inbar[18] = ~in[18];
  assign inbar[19] = ~in[19];
  assign inbar[20] = ~in[20];
  assign inbar[21] = ~in[21];
  assign inbar[22] = ~in[22];
  assign inbar[23] = ~in[23];
  assign inbar[24] = ~in[24];
  assign inbar[25] = ~in[25];
  assign inbar[26] = ~in[26];
  assign inbar[27] = ~in[27];
  assign inbar[28] = ~in[28];
  assign inbar[29] = ~in[29];
  assign inbar[30] = ~in[30];
  assign inbar[31] = ~in[31];
  assign inbar[32] = ~in[32];
  assign inbar[33] = ~in[33];
  assign inbar[34] = ~in[34];
  assign inbar[35] = ~in[35];
  assign inbar[36] = ~in[36];
  assign inbar[37] = ~in[37];
  assign inbar[38] = ~in[38];
  assign inbar[39] = ~in[39];
  assign inbar[40] = ~in[40];
  assign inbar[41] = ~in[41];
  assign inbar[42] = ~in[42];
  assign inbar[43] = ~in[43];
  assign inbar[44] = ~in[44];
  assign inbar[45] = ~in[45];
  assign inbar[46] = ~in[46];
  assign inbar[47] = ~in[47];
  assign inbar[48] = ~in[48];
  assign inbar[49] = ~in[49];
  assign inbar[50] = ~in[50];
  assign inbar[51] = ~in[51];
  assign inbar[52] = ~in[52];
  assign inbar[53] = ~in[53];
  assign inbar[54] = ~in[54];
  assign inbar[55] = ~in[55];
  assign inbar[56] = ~in[56];
  assign inbar[57] = ~in[57];
  assign inbar[58] = ~in[58];
  assign inbar[59] = ~in[59];
  assign inbar[60] = ~in[60];
  assign inbar[61] = ~in[61];
  assign inbar[62] = ~in[62];
  assign inbar[63] = ~in[63];
  assign inbar[64] = ~in[64];
  assign inbar[65] = ~in[65];
  assign inbar[66] = ~in[66];
  assign inbar[67] = ~in[67];
  assign inbar[68] = ~in[68];
  assign inbar[69] = ~in[69];
  assign inbar[70] = ~in[70];
  assign inbar[71] = ~in[71];
  assign inbar[72] = ~in[72];
  assign inbar[73] = ~in[73];
  assign inbar[74] = ~in[74];
  assign inbar[75] = ~in[75];
  assign inbar[76] = ~in[76];
  assign inbar[77] = ~in[77];
  assign inbar[78] = ~in[78];
  assign inbar[79] = ~in[79];
  assign inbar[80] = ~in[80];
  assign inbar[81] = ~in[81];
  assign inbar[82] = ~in[82];
  assign inbar[83] = ~in[83];
  assign inbar[84] = ~in[84];
  assign inbar[85] = ~in[85];
  assign inbar[86] = ~in[86];
  assign inbar[87] = ~in[87];
  assign inbar[88] = ~in[88];
  assign inbar[89] = ~in[89];
  assign inbar[90] = ~in[90];
  assign inbar[91] = ~in[91];
  assign inbar[92] = ~in[92];
  assign inbar[93] = ~in[93];
  assign inbar[94] = ~in[94];
  assign inbar[95] = ~in[95];
  assign inbar[96] = ~in[96];
  assign inbar[97] = ~in[97];
  assign inbar[98] = ~in[98];
  assign inbar[99] = ~in[99];
  assign inbar[100] = ~in[100];
  assign inbar[101] = ~in[101];
  assign inbar[102] = ~in[102];
  assign inbar[103] = ~in[103];
  assign inbar[104] = ~in[104];
  assign inbar[105] = ~in[105];
  assign inbar[106] = ~in[106];
  assign inbar[107] = ~in[107];
  assign inbar[108] = ~in[108];
  assign inbar[109] = ~in[109];
  assign inbar[110] = ~in[110];
  assign inbar[111] = ~in[111];
  assign inbar[112] = ~in[112];
  assign inbar[113] = ~in[113];
  assign inbar[114] = ~in[114];
  assign inbar[115] = ~in[115];
  assign inbar[116] = ~in[116];
  assign inbar[117] = ~in[117];
  assign inbar[118] = ~in[118];
  assign inbar[119] = ~in[119];
  assign inbar[120] = ~in[120];
  assign inbar[121] = ~in[121];
  assign inbar[122] = ~in[122];
  assign inbar[123] = ~in[123];
  assign inbar[124] = ~in[124];
  assign inbar[125] = ~in[125];
  assign inbar[126] = ~in[126];
  assign inbar[127] = ~in[127];
  assign inbar[128] = ~in[128];
  assign inbar[129] = ~in[129];
  assign inbar[130] = ~in[130];
  assign inbar[131] = ~in[131];
  assign inbar[132] = ~in[132];
  assign inbar[133] = ~in[133];
  assign inbar[134] = ~in[134];
  assign inbar[135] = ~in[135];
  assign inbar[136] = ~in[136];
  assign inbar[137] = ~in[137];
  assign inbar[138] = ~in[138];
  assign inbar[139] = ~in[139];
  assign inbar[140] = ~in[140];
  assign inbar[141] = ~in[141];
  assign inbar[142] = ~in[142];
  assign inbar[143] = ~in[143];
  assign inbar[144] = ~in[144];
  assign inbar[145] = ~in[145];
  assign inbar[146] = ~in[146];
  assign inbar[147] = ~in[147];
  assign inbar[148] = ~in[148];
  assign inbar[149] = ~in[149];
  assign inbar[150] = ~in[150];
  assign inbar[151] = ~in[151];
  assign inbar[152] = ~in[152];
  assign inbar[153] = ~in[153];
  assign inbar[154] = ~in[154];
  assign inbar[155] = ~in[155];
  assign inbar[156] = ~in[156];
  assign inbar[157] = ~in[157];
  assign inbar[158] = ~in[158];
  assign inbar[159] = ~in[159];
  assign inbar[160] = ~in[160];
  assign inbar[161] = ~in[161];
  assign inbar[162] = ~in[162];
  assign inbar[163] = ~in[163];
  assign inbar[164] = ~in[164];
  assign inbar[165] = ~in[165];
  assign inbar[166] = ~in[166];
  assign inbar[167] = ~in[167];
  assign inbar[168] = ~in[168];
  assign inbar[169] = ~in[169];
  assign inbar[170] = ~in[170];
  assign inbar[171] = ~in[171];
  assign inbar[172] = ~in[172];
  assign inbar[173] = ~in[173];
  assign inbar[174] = ~in[174];
  assign inbar[175] = ~in[175];
  assign inbar[176] = ~in[176];
  assign inbar[177] = ~in[177];
  assign inbar[178] = ~in[178];
  assign inbar[179] = ~in[179];
  assign inbar[180] = ~in[180];
  assign inbar[181] = ~in[181];
  assign inbar[182] = ~in[182];
  assign inbar[183] = ~in[183];
  assign inbar[184] = ~in[184];
  assign inbar[185] = ~in[185];
  assign inbar[186] = ~in[186];
  assign inbar[187] = ~in[187];
  assign inbar[188] = ~in[188];
  assign inbar[189] = ~in[189];
  assign inbar[190] = ~in[190];
  assign inbar[191] = ~in[191];
  assign inbar[192] = ~in[192];
  assign inbar[193] = ~in[193];
  assign inbar[194] = ~in[194];
  assign inbar[195] = ~in[195];
  assign inbar[196] = ~in[196];
  assign inbar[197] = ~in[197];
  assign inbar[198] = ~in[198];
  assign inbar[199] = ~in[199];
  assign inbar[200] = ~in[200];
  assign inbar[201] = ~in[201];
  assign inbar[202] = ~in[202];
  assign inbar[203] = ~in[203];
  assign inbar[204] = ~in[204];
  assign inbar[205] = ~in[205];
  assign inbar[206] = ~in[206];
  assign inbar[207] = ~in[207];
  assign inbar[208] = ~in[208];
  assign inbar[209] = ~in[209];
  assign inbar[210] = ~in[210];
  assign inbar[211] = ~in[211];
  assign inbar[212] = ~in[212];
  assign inbar[213] = ~in[213];
  assign inbar[214] = ~in[214];
  assign inbar[215] = ~in[215];
  assign inbar[216] = ~in[216];
  assign inbar[217] = ~in[217];
  assign inbar[218] = ~in[218];
  assign inbar[219] = ~in[219];
  assign inbar[220] = ~in[220];
  assign inbar[221] = ~in[221];
  assign inbar[222] = ~in[222];
  assign inbar[223] = ~in[223];
  assign inbar[224] = ~in[224];
  assign inbar[225] = ~in[225];
  assign inbar[226] = ~in[226];
  assign inbar[227] = ~in[227];
  assign inbar[228] = ~in[228];
  assign inbar[229] = ~in[229];
  assign inbar[230] = ~in[230];
  assign inbar[231] = ~in[231];
  assign inbar[232] = ~in[232];
  assign inbar[233] = ~in[233];
  assign inbar[234] = ~in[234];
  assign inbar[235] = ~in[235];
  assign inbar[236] = ~in[236];
  assign inbar[237] = ~in[237];
  assign inbar[238] = ~in[238];
  assign inbar[239] = ~in[239];
  assign inbar[240] = ~in[240];
  assign inbar[241] = ~in[241];
  assign inbar[242] = ~in[242];
  assign inbar[243] = ~in[243];
  assign inbar[244] = ~in[244];
  assign inbar[245] = ~in[245];
  assign inbar[246] = ~in[246];
  assign inbar[247] = ~in[247];
  assign inbar[248] = ~in[248];
  assign inbar[249] = ~in[249];
  assign inbar[250] = ~in[250];
  assign inbar[251] = ~in[251];
  assign inbar[252] = ~in[252];
  assign inbar[253] = ~in[253];
  assign inbar[254] = ~in[254];
  assign inbar[255] = ~in[255];
  //input_done

  output [7:0] out;
  reg [7:0] outbar;
  //output_done

  wire   in_81, in_80, in_79, in_78, in_77, in_76, in_75, in_74, in_73, in_72,
         in_71, in_70, in_69, in_68, in_67, in_66, in_65, in_64, in_63, in_62,
         in_61, in_60, in_59, in_58, in_57, in_56, in_55, in_54, in_53, in_52,
         in_51, in_50, in_49, in_48, in_47, in_46, in_45, in_44, in_43, in_42,
         in_41, in_40, in_39, in_38, in_37, in_36, in_35, in_34, in_33, in_32,
         in_31, in_30, in_29, in_28, in_27, in_26, in_25, in_24, in_23, in_22,
         in_21, in_20, in_19, in_18, in_17, in_16, in_15, in_14, in_13, in_12,
         in_11, in_10, in_9, in_8, in_7, in_6, in_5, in_4, in_3, in_2, in_1,
         in_0, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972;
  wire in_81bar, in_80bar, in_79bar, in_78bar, in_77bar, in_76bar, in_75bar, in_74bar, in_73bar, in_72bar, in_71bar, in_70bar, in_69bar, in_68bar, in_67bar, in_66bar, in_65bar, in_64bar, in_63bar, in_62bar, in_61bar, in_60bar, in_59bar, in_58bar, in_57bar, in_56bar, in_55bar, in_54bar, in_53bar, in_52bar, in_51bar, in_50bar, in_49bar, in_48bar, in_47bar, in_46bar, in_45bar, in_44bar, in_43bar, in_42bar, in_41bar, in_40bar, in_39bar, in_38bar, in_37bar, in_36bar, in_35bar, in_34bar, in_33bar, in_32bar, in_31bar, in_30bar, in_29bar, in_28bar, in_27bar, in_26bar, in_25bar, in_24bar, in_23bar, in_22bar, in_21bar, in_20bar, in_19bar, in_18bar, in_17bar, in_16bar, in_15bar, in_14bar, in_13bar, in_12bar, in_11bar, in_10bar, in_9bar, in_8bar, in_7bar, in_6bar, in_5bar, in_4bar, in_3bar, in_2bar, in_1bar, in_0bar, n487bar, n488bar, n489bar, n490bar, n491bar, n492bar, n493bar, n494bar, n495bar, n496bar, n497bar, n498bar, n499bar, n500bar, n501bar, n502bar, n503bar, n504bar, n505bar, n506bar, n507bar, n508bar, n509bar, n510bar, n511bar, n512bar, n513bar, n514bar, n515bar, n516bar, n517bar, n518bar, n519bar, n520bar, n521bar, n522bar, n523bar, n524bar, n525bar, n526bar, n527bar, n528bar, n529bar, n530bar, n531bar, n532bar, n533bar, n534bar, n535bar, n536bar, n537bar, n538bar, n539bar, n540bar, n541bar, n542bar, n543bar, n544bar, n545bar, n546bar, n547bar, n548bar, n549bar, n550bar, n551bar, n552bar, n553bar, n554bar, n555bar, n556bar, n557bar, n558bar, n559bar, n560bar, n561bar, n562bar, n563bar, n564bar, n565bar, n566bar, n567bar, n568bar, n569bar, n570bar, n571bar, n572bar, n573bar, n574bar, n575bar, n576bar, n577bar, n578bar, n579bar, n580bar, n581bar, n582bar, n583bar, n584bar, n585bar, n586bar, n587bar, n588bar, n589bar, n590bar, n591bar, n592bar, n593bar, n594bar, n595bar, n596bar, n597bar, n598bar, n599bar, n600bar, n601bar, n602bar, n603bar, n604bar, n605bar, n606bar, n607bar, n608bar, n609bar, n610bar, n611bar, n612bar, n613bar, n614bar, n615bar, n616bar, n617bar, n618bar, n619bar, n620bar, n621bar, n622bar, n623bar, n624bar, n625bar, n626bar, n627bar, n628bar, n629bar, n630bar, n631bar, n632bar, n633bar, n634bar, n635bar, n636bar, n637bar, n638bar, n639bar, n640bar, n641bar, n642bar, n643bar, n644bar, n645bar, n646bar, n647bar, n648bar, n649bar, n650bar, n651bar, n652bar, n653bar, n654bar, n655bar, n656bar, n657bar, n658bar, n659bar, n660bar, n661bar, n662bar, n663bar, n664bar, n665bar, n666bar, n667bar, n668bar, n669bar, n670bar, n671bar, n672bar, n673bar, n674bar, n675bar, n676bar, n677bar, n678bar, n679bar, n680bar, n681bar, n682bar, n683bar, n684bar, n685bar, n686bar, n687bar, n688bar, n689bar, n690bar, n691bar, n692bar, n693bar, n694bar, n695bar, n696bar, n697bar, n698bar, n699bar, n700bar, n701bar, n702bar, n703bar, n704bar, n705bar, n706bar, n707bar, n708bar, n709bar, n710bar, n711bar, n712bar, n713bar, n714bar, n715bar, n716bar, n717bar, n718bar, n719bar, n720bar, n721bar, n722bar, n723bar, n724bar, n725bar, n726bar, n727bar, n728bar, n729bar, n730bar, n731bar, n732bar, n733bar, n734bar, n735bar, n736bar, n737bar, n738bar, n739bar, n740bar, n741bar, n742bar, n743bar, n744bar, n745bar, n746bar, n747bar, n748bar, n749bar, n750bar, n751bar, n752bar, n753bar, n754bar, n755bar, n756bar, n757bar, n758bar, n759bar, n760bar, n761bar, n762bar, n763bar, n764bar, n765bar, n766bar, n767bar, n768bar, n769bar, n770bar, n771bar, n772bar, n773bar, n774bar, n775bar, n776bar, n777bar, n778bar, n779bar, n780bar, n781bar, n782bar, n783bar, n784bar, n785bar, n786bar, n787bar, n788bar, n789bar, n790bar, n791bar, n792bar, n793bar, n794bar, n795bar, n796bar, n797bar, n798bar, n799bar, n800bar, n801bar, n802bar, n803bar, n804bar, n805bar, n806bar, n807bar, n808bar, n809bar, n810bar, n811bar, n812bar, n813bar, n814bar, n815bar, n816bar, n817bar, n818bar, n819bar, n820bar, n821bar, n822bar, n823bar, n824bar, n825bar, n826bar, n827bar, n828bar, n829bar, n830bar, n831bar, n832bar, n833bar, n834bar, n835bar, n836bar, n837bar, n838bar, n839bar, n840bar, n841bar, n842bar, n843bar, n844bar, n845bar, n846bar, n847bar, n848bar, n849bar, n850bar, n851bar, n852bar, n853bar, n854bar, n855bar, n856bar, n857bar, n858bar, n859bar, n860bar, n861bar, n862bar, n863bar, n864bar, n865bar, n866bar, n867bar, n868bar, n869bar, n870bar, n871bar, n872bar, n873bar, n874bar, n875bar, n876bar, n877bar, n878bar, n879bar, n880bar, n881bar, n882bar, n883bar, n884bar, n885bar, n886bar, n887bar, n888bar, n889bar, n890bar, n891bar, n892bar, n893bar, n894bar, n895bar, n896bar, n897bar, n898bar, n899bar, n900bar, n901bar, n902bar, n903bar, n904bar, n905bar, n906bar, n907bar, n908bar, n909bar, n910bar, n911bar, n912bar, n913bar, n914bar, n915bar, n916bar, n917bar, n918bar, n919bar, n920bar, n921bar, n922bar, n923bar, n924bar, n925bar, n926bar, n927bar, n928bar, n929bar, n930bar, n931bar, n932bar, n933bar, n934bar, n935bar, n936bar, n937bar, n938bar, n939bar, n940bar, n941bar, n942bar, n943bar, n944bar, n945bar, n946bar, n947bar, n948bar, n949bar, n950bar, n951bar, n952bar, n953bar, n954bar, n955bar, n956bar, n957bar, n958bar, n959bar, n960bar, n961bar, n962bar, n963bar, n964bar, n965bar, n966bar, n967bar, n968bar, n969bar, n970bar, n971bar, n972bar;
  //wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];

  OR2_X1 U1 ( .A1(n972), .A2(n971), .ZN(out[7]) );
  AND2_X1 U1bar ( .A1(n972bar), .A2(n971bar), .ZN(outbar[7]);
  OR2_X1 U2 ( .A1(n970), .A2(n969), .ZN(n971) );
  AND2_X1 U2bar ( .A1(n970bar), .A2(n969bar), .ZN(n971bar);
  OR2_X1 U3 ( .A1(n968), .A2(n967), .ZN(n969) );
  AND2_X1 U3bar ( .A1(n968bar), .A2(n967bar), .ZN(n969bar);
  OR2_X1 U4 ( .A1(n966), .A2(n965), .ZN(n967) );
  AND2_X1 U4bar ( .A1(n966bar), .A2(n965bar), .ZN(n967bar);
  OR2_X1 U5 ( .A1(n964), .A2(n963), .ZN(n968) );
  AND2_X1 U5bar ( .A1(n964bar), .A2(n963bar), .ZN(n968bar);
  OR2_X1 U6 ( .A1(in[116]), .A2(n962), .ZN(n963) );
  AND2_X1 U6bar ( .A1(inbar[116]), .A2(n962bar), .ZN(n963bar);
  OR2_X1 U7 ( .A1(n961), .A2(n960), .ZN(n970) );
  AND2_X1 U7bar ( .A1(n961bar), .A2(n960bar), .ZN(n970bar);
  OR2_X1 U8 ( .A1(in[150]), .A2(in[127]), .ZN(n960) );
  AND2_X1 U8bar ( .A1(inbar[150]), .A2(inbar[127]), .ZN(n960bar);
  OR2_X1 U9 ( .A1(in[160]), .A2(n959), .ZN(n961) );
  AND2_X1 U9bar ( .A1(inbar[160]), .A2(n959bar), .ZN(n961bar);
  OR2_X1 U10 ( .A1(in[252]), .A2(in[168]), .ZN(n959) );
  AND2_X1 U10bar ( .A1(inbar[252]), .A2(inbar[168]), .ZN(n959bar);
  OR2_X1 U11 ( .A1(n958), .A2(n957), .ZN(n972) );
  AND2_X1 U11bar ( .A1(n958bar), .A2(n957bar), .ZN(n972bar);
  OR2_X1 U12 ( .A1(n956), .A2(n955), .ZN(n957) );
  AND2_X1 U12bar ( .A1(n956bar), .A2(n955bar), .ZN(n957bar);
  OR2_X1 U13 ( .A1(in_17), .A2(in[96]), .ZN(n955) );
  AND2_X1 U13bar ( .A1(in_17bar), .A2(inbar[96]), .ZN(n955bar);
  OR2_X1 U14 ( .A1(in_23), .A2(n954), .ZN(n956) );
  AND2_X1 U14bar ( .A1(in_23bar), .A2(n954bar), .ZN(n956bar);
  OR2_X1 U15 ( .A1(in_31), .A2(in_26), .ZN(n954) );
  AND2_X1 U15bar ( .A1(in_31bar), .A2(in_26bar), .ZN(n954bar);
  OR2_X1 U16 ( .A1(n953), .A2(n952), .ZN(n958) );
  AND2_X1 U16bar ( .A1(n953bar), .A2(n952bar), .ZN(n958bar);
  OR2_X1 U17 ( .A1(in_58), .A2(in_4), .ZN(n952) );
  AND2_X1 U17bar ( .A1(in_58bar), .A2(in_4bar), .ZN(n952bar);
  OR2_X1 U18 ( .A1(in_59), .A2(n951), .ZN(n953) );
  AND2_X1 U18bar ( .A1(in_59bar), .A2(n951bar), .ZN(n953bar);
  OR2_X1 U19 ( .A1(in_71), .A2(in_62), .ZN(n951) );
  AND2_X1 U19bar ( .A1(in_71bar), .A2(in_62bar), .ZN(n951bar);
  OR2_X1 U20 ( .A1(n950), .A2(n949), .ZN(out[6]) );
  AND2_X1 U20bar ( .A1(n950bar), .A2(n949bar), .ZN(outbar[6]);
  OR2_X1 U21 ( .A1(n948), .A2(n947), .ZN(n949) );
  AND2_X1 U21bar ( .A1(n948bar), .A2(n947bar), .ZN(n949bar);
  OR2_X1 U22 ( .A1(n946), .A2(n945), .ZN(n947) );
  AND2_X1 U22bar ( .A1(n946bar), .A2(n945bar), .ZN(n947bar);
  OR2_X1 U23 ( .A1(n944), .A2(n943), .ZN(n945) );
  AND2_X1 U23bar ( .A1(n944bar), .A2(n943bar), .ZN(n945bar);
  OR2_X1 U24 ( .A1(n942), .A2(n941), .ZN(n946) );
  AND2_X1 U24bar ( .A1(n942bar), .A2(n941bar), .ZN(n946bar);
  OR2_X1 U25 ( .A1(in[101]), .A2(n940), .ZN(n941) );
  AND2_X1 U25bar ( .A1(inbar[101]), .A2(n940bar), .ZN(n941bar);
  OR2_X1 U26 ( .A1(n939), .A2(n938), .ZN(n948) );
  AND2_X1 U26bar ( .A1(n939bar), .A2(n938bar), .ZN(n948bar);
  OR2_X1 U27 ( .A1(in[114]), .A2(in[104]), .ZN(n938) );
  AND2_X1 U27bar ( .A1(inbar[114]), .A2(inbar[104]), .ZN(n938bar);
  OR2_X1 U28 ( .A1(in[128]), .A2(n937), .ZN(n939) );
  AND2_X1 U28bar ( .A1(inbar[128]), .A2(n937bar), .ZN(n939bar);
  OR2_X1 U29 ( .A1(in[136]), .A2(in[134]), .ZN(n937) );
  AND2_X1 U29bar ( .A1(inbar[136]), .A2(inbar[134]), .ZN(n937bar);
  OR2_X1 U30 ( .A1(n936), .A2(n935), .ZN(n950) );
  AND2_X1 U30bar ( .A1(n936bar), .A2(n935bar), .ZN(n950bar);
  OR2_X1 U31 ( .A1(n934), .A2(n933), .ZN(n935) );
  AND2_X1 U31bar ( .A1(n934bar), .A2(n933bar), .ZN(n935bar);
  OR2_X1 U32 ( .A1(in[177]), .A2(in[164]), .ZN(n933) );
  AND2_X1 U32bar ( .A1(inbar[177]), .A2(inbar[164]), .ZN(n933bar);
  OR2_X1 U33 ( .A1(in[212]), .A2(n932), .ZN(n934) );
  AND2_X1 U33bar ( .A1(inbar[212]), .A2(n932bar), .ZN(n934bar);
  OR2_X1 U34 ( .A1(in[248]), .A2(in[221]), .ZN(n932) );
  AND2_X1 U34bar ( .A1(inbar[248]), .A2(inbar[221]), .ZN(n932bar);
  OR2_X1 U35 ( .A1(n931), .A2(n930), .ZN(n936) );
  AND2_X1 U35bar ( .A1(n931bar), .A2(n930bar), .ZN(n936bar);
  OR2_X1 U36 ( .A1(in_18), .A2(in[93]), .ZN(n930) );
  AND2_X1 U36bar ( .A1(in_18bar), .A2(inbar[93]), .ZN(n930bar);
  OR2_X1 U37 ( .A1(in_31), .A2(n929), .ZN(n931) );
  AND2_X1 U37bar ( .A1(in_31bar), .A2(n929bar), .ZN(n931bar);
  OR2_X1 U38 ( .A1(in_7), .A2(in_39), .ZN(n929) );
  AND2_X1 U38bar ( .A1(in_7bar), .A2(in_39bar), .ZN(n929bar);
  OR2_X1 U39 ( .A1(n928), .A2(n927), .ZN(out[5]) );
  AND2_X1 U39bar ( .A1(n928bar), .A2(n927bar), .ZN(outbar[5]);
  OR2_X1 U40 ( .A1(n926), .A2(n925), .ZN(n927) );
  AND2_X1 U40bar ( .A1(n926bar), .A2(n925bar), .ZN(n927bar);
  OR2_X1 U41 ( .A1(n924), .A2(n923), .ZN(n925) );
  AND2_X1 U41bar ( .A1(n924bar), .A2(n923bar), .ZN(n925bar);
  OR2_X1 U42 ( .A1(n922), .A2(n921), .ZN(n923) );
  AND2_X1 U42bar ( .A1(n922bar), .A2(n921bar), .ZN(n923bar);
  OR2_X1 U43 ( .A1(n940), .A2(n920), .ZN(n924) );
  AND2_X1 U43bar ( .A1(n940bar), .A2(n920bar), .ZN(n924bar);
  OR2_X1 U44 ( .A1(in[111]), .A2(n919), .ZN(n920) );
  AND2_X1 U44bar ( .A1(inbar[111]), .A2(n919bar), .ZN(n920bar);
  OR2_X1 U45 ( .A1(n918), .A2(n917), .ZN(n940) );
  AND2_X1 U45bar ( .A1(n918bar), .A2(n917bar), .ZN(n940bar);
  OR2_X1 U46 ( .A1(n916), .A2(n915), .ZN(n917) );
  AND2_X1 U46bar ( .A1(n916bar), .A2(n915bar), .ZN(n917bar);
  OR2_X1 U47 ( .A1(n914), .A2(n913), .ZN(n915) );
  AND2_X1 U47bar ( .A1(n914bar), .A2(n913bar), .ZN(n915bar);
  OR2_X1 U48 ( .A1(in[140]), .A2(in[131]), .ZN(n913) );
  AND2_X1 U48bar ( .A1(inbar[140]), .A2(inbar[131]), .ZN(n913bar);
  OR2_X1 U49 ( .A1(in[160]), .A2(in[144]), .ZN(n914) );
  AND2_X1 U49bar ( .A1(inbar[160]), .A2(inbar[144]), .ZN(n914bar);
  OR2_X1 U50 ( .A1(n912), .A2(n911), .ZN(n916) );
  AND2_X1 U50bar ( .A1(n912bar), .A2(n911bar), .ZN(n916bar);
  OR2_X1 U51 ( .A1(in[179]), .A2(in[174]), .ZN(n911) );
  AND2_X1 U51bar ( .A1(inbar[179]), .A2(inbar[174]), .ZN(n911bar);
  OR2_X1 U52 ( .A1(in[188]), .A2(in[184]), .ZN(n912) );
  AND2_X1 U52bar ( .A1(inbar[188]), .A2(inbar[184]), .ZN(n912bar);
  OR2_X1 U53 ( .A1(n910), .A2(n909), .ZN(n918) );
  AND2_X1 U53bar ( .A1(n910bar), .A2(n909bar), .ZN(n918bar);
  OR2_X1 U54 ( .A1(n908), .A2(n907), .ZN(n909) );
  AND2_X1 U54bar ( .A1(n908bar), .A2(n907bar), .ZN(n909bar);
  OR2_X1 U55 ( .A1(in[216]), .A2(in[200]), .ZN(n907) );
  AND2_X1 U55bar ( .A1(inbar[216]), .A2(inbar[200]), .ZN(n907bar);
  OR2_X1 U56 ( .A1(in[228]), .A2(in[224]), .ZN(n908) );
  AND2_X1 U56bar ( .A1(inbar[228]), .A2(inbar[224]), .ZN(n908bar);
  OR2_X1 U57 ( .A1(n906), .A2(n905), .ZN(n910) );
  AND2_X1 U57bar ( .A1(n906bar), .A2(n905bar), .ZN(n910bar);
  OR2_X1 U58 ( .A1(in[247]), .A2(in[235]), .ZN(n905) );
  AND2_X1 U58bar ( .A1(inbar[247]), .A2(inbar[235]), .ZN(n905bar);
  OR2_X1 U59 ( .A1(in_42), .A2(in[83]), .ZN(n906) );
  AND2_X1 U59bar ( .A1(in_42bar), .A2(inbar[83]), .ZN(n906bar);
  OR2_X1 U60 ( .A1(n904), .A2(n903), .ZN(n926) );
  AND2_X1 U60bar ( .A1(n904bar), .A2(n903bar), .ZN(n926bar);
  OR2_X1 U61 ( .A1(in[166]), .A2(in[123]), .ZN(n903) );
  AND2_X1 U61bar ( .A1(inbar[166]), .A2(inbar[123]), .ZN(n903bar);
  OR2_X1 U62 ( .A1(in[170]), .A2(n902), .ZN(n904) );
  AND2_X1 U62bar ( .A1(inbar[170]), .A2(n902bar), .ZN(n904bar);
  OR2_X1 U63 ( .A1(in[194]), .A2(in[183]), .ZN(n902) );
  AND2_X1 U63bar ( .A1(inbar[194]), .A2(inbar[183]), .ZN(n902bar);
  OR2_X1 U64 ( .A1(n901), .A2(n900), .ZN(n928) );
  AND2_X1 U64bar ( .A1(n901bar), .A2(n900bar), .ZN(n928bar);
  OR2_X1 U65 ( .A1(n899), .A2(n898), .ZN(n900) );
  AND2_X1 U65bar ( .A1(n899bar), .A2(n898bar), .ZN(n900bar);
  OR2_X1 U66 ( .A1(in[241]), .A2(in[238]), .ZN(n898) );
  AND2_X1 U66bar ( .A1(inbar[241]), .A2(inbar[238]), .ZN(n898bar);
  OR2_X1 U67 ( .A1(in[250]), .A2(n897), .ZN(n899) );
  AND2_X1 U67bar ( .A1(inbar[250]), .A2(n897bar), .ZN(n899bar);
  OR2_X1 U68 ( .A1(in_24), .A2(in[84]), .ZN(n897) );
  AND2_X1 U68bar ( .A1(in_24bar), .A2(inbar[84]), .ZN(n897bar);
  OR2_X1 U69 ( .A1(n896), .A2(n895), .ZN(n901) );
  AND2_X1 U69bar ( .A1(n896bar), .A2(n895bar), .ZN(n901bar);
  OR2_X1 U70 ( .A1(in_41), .A2(in_29), .ZN(n895) );
  AND2_X1 U70bar ( .A1(in_41bar), .A2(in_29bar), .ZN(n895bar);
  OR2_X1 U71 ( .A1(in_66), .A2(n894), .ZN(n896) );
  AND2_X1 U71bar ( .A1(in_66bar), .A2(n894bar), .ZN(n896bar);
  OR2_X1 U72 ( .A1(in_76), .A2(in_71), .ZN(n894) );
  AND2_X1 U72bar ( .A1(in_76bar), .A2(in_71bar), .ZN(n894bar);
  OR2_X1 U73 ( .A1(n893), .A2(n892), .ZN(out[4]) );
  AND2_X1 U73bar ( .A1(n893bar), .A2(n892bar), .ZN(outbar[4]);
  OR2_X1 U74 ( .A1(n891), .A2(n890), .ZN(n892) );
  AND2_X1 U74bar ( .A1(n891bar), .A2(n890bar), .ZN(n892bar);
  OR2_X1 U75 ( .A1(n889), .A2(n888), .ZN(n890) );
  AND2_X1 U75bar ( .A1(n889bar), .A2(n888bar), .ZN(n890bar);
  OR2_X1 U76 ( .A1(n922), .A2(n887), .ZN(n888) );
  AND2_X1 U76bar ( .A1(n922bar), .A2(n887bar), .ZN(n888bar);
  OR2_X1 U77 ( .A1(n886), .A2(n885), .ZN(n922) );
  AND2_X1 U77bar ( .A1(n886bar), .A2(n885bar), .ZN(n922bar);
  OR2_X1 U78 ( .A1(n884), .A2(n883), .ZN(n885) );
  AND2_X1 U78bar ( .A1(n884bar), .A2(n883bar), .ZN(n885bar);
  OR2_X1 U79 ( .A1(n882), .A2(n881), .ZN(n883) );
  AND2_X1 U79bar ( .A1(n882bar), .A2(n881bar), .ZN(n883bar);
  OR2_X1 U80 ( .A1(in[118]), .A2(in[109]), .ZN(n881) );
  AND2_X1 U80bar ( .A1(inbar[118]), .A2(inbar[109]), .ZN(n881bar);
  OR2_X1 U81 ( .A1(in[139]), .A2(in[120]), .ZN(n882) );
  AND2_X1 U81bar ( .A1(inbar[139]), .A2(inbar[120]), .ZN(n882bar);
  OR2_X1 U82 ( .A1(n880), .A2(n879), .ZN(n884) );
  AND2_X1 U82bar ( .A1(n880bar), .A2(n879bar), .ZN(n884bar);
  OR2_X1 U83 ( .A1(in[198]), .A2(in[154]), .ZN(n879) );
  AND2_X1 U83bar ( .A1(inbar[198]), .A2(inbar[154]), .ZN(n879bar);
  OR2_X1 U84 ( .A1(in[210]), .A2(in[205]), .ZN(n880) );
  AND2_X1 U84bar ( .A1(inbar[210]), .A2(inbar[205]), .ZN(n880bar);
  OR2_X1 U85 ( .A1(n878), .A2(n877), .ZN(n886) );
  AND2_X1 U85bar ( .A1(n878bar), .A2(n877bar), .ZN(n886bar);
  OR2_X1 U86 ( .A1(n876), .A2(n875), .ZN(n877) );
  AND2_X1 U86bar ( .A1(n876bar), .A2(n875bar), .ZN(n877bar);
  OR2_X1 U87 ( .A1(in[219]), .A2(in[217]), .ZN(n875) );
  AND2_X1 U87bar ( .A1(inbar[219]), .A2(inbar[217]), .ZN(n875bar);
  OR2_X1 U88 ( .A1(in[86]), .A2(in[252]), .ZN(n876) );
  AND2_X1 U88bar ( .A1(inbar[86]), .A2(inbar[252]), .ZN(n876bar);
  OR2_X1 U89 ( .A1(n874), .A2(n873), .ZN(n878) );
  AND2_X1 U89bar ( .A1(n874bar), .A2(n873bar), .ZN(n878bar);
  OR2_X1 U90 ( .A1(in_40), .A2(in[91]), .ZN(n873) );
  AND2_X1 U90bar ( .A1(in_40bar), .A2(inbar[91]), .ZN(n873bar);
  OR2_X1 U91 ( .A1(in_8), .A2(in_46), .ZN(n874) );
  AND2_X1 U91bar ( .A1(in_8bar), .A2(in_46bar), .ZN(n874bar);
  OR2_X1 U92 ( .A1(n872), .A2(n871), .ZN(n889) );
  AND2_X1 U92bar ( .A1(n872bar), .A2(n871bar), .ZN(n889bar);
  OR2_X1 U93 ( .A1(in[117]), .A2(n943), .ZN(n871) );
  AND2_X1 U93bar ( .A1(inbar[117]), .A2(n943bar), .ZN(n871bar);
  OR2_X1 U94 ( .A1(n870), .A2(n869), .ZN(n943) );
  AND2_X1 U94bar ( .A1(n870bar), .A2(n869bar), .ZN(n943bar);
  OR2_X1 U95 ( .A1(n868), .A2(n867), .ZN(n869) );
  AND2_X1 U95bar ( .A1(n868bar), .A2(n867bar), .ZN(n869bar);
  OR2_X1 U96 ( .A1(n866), .A2(n865), .ZN(n867) );
  AND2_X1 U96bar ( .A1(n866bar), .A2(n865bar), .ZN(n867bar);
  OR2_X1 U97 ( .A1(n864), .A2(n863), .ZN(n865) );
  AND2_X1 U97bar ( .A1(n864bar), .A2(n863bar), .ZN(n865bar);
  OR2_X1 U98 ( .A1(in[108]), .A2(n919), .ZN(n866) );
  AND2_X1 U98bar ( .A1(inbar[108]), .A2(n919bar), .ZN(n866bar);
  OR2_X1 U99 ( .A1(n862), .A2(n861), .ZN(n919) );
  AND2_X1 U99bar ( .A1(n862bar), .A2(n861bar), .ZN(n919bar);
  OR2_X1 U100 ( .A1(n860), .A2(n859), .ZN(n861) );
  AND2_X1 U100bar ( .A1(n860bar), .A2(n859bar), .ZN(n861bar);
  OR2_X1 U101 ( .A1(n858), .A2(n857), .ZN(n859) );
  AND2_X1 U101bar ( .A1(n858bar), .A2(n857bar), .ZN(n859bar);
  OR2_X1 U102 ( .A1(in[119]), .A2(in[105]), .ZN(n857) );
  AND2_X1 U102bar ( .A1(inbar[119]), .A2(inbar[105]), .ZN(n857bar);
  OR2_X1 U103 ( .A1(in[186]), .A2(in[175]), .ZN(n858) );
  AND2_X1 U103bar ( .A1(inbar[186]), .A2(inbar[175]), .ZN(n858bar);
  OR2_X1 U104 ( .A1(n856), .A2(n855), .ZN(n860) );
  AND2_X1 U104bar ( .A1(n856bar), .A2(n855bar), .ZN(n860bar);
  OR2_X1 U105 ( .A1(in[202]), .A2(in[193]), .ZN(n855) );
  AND2_X1 U105bar ( .A1(inbar[202]), .A2(inbar[193]), .ZN(n855bar);
  OR2_X1 U106 ( .A1(in[225]), .A2(in[208]), .ZN(n856) );
  AND2_X1 U106bar ( .A1(inbar[225]), .A2(inbar[208]), .ZN(n856bar);
  OR2_X1 U107 ( .A1(n854), .A2(n853), .ZN(n862) );
  AND2_X1 U107bar ( .A1(n854bar), .A2(n853bar), .ZN(n862bar);
  OR2_X1 U108 ( .A1(n852), .A2(n851), .ZN(n853) );
  AND2_X1 U108bar ( .A1(n852bar), .A2(n851bar), .ZN(n853bar);
  OR2_X1 U109 ( .A1(in_1), .A2(in[85]), .ZN(n851) );
  AND2_X1 U109bar ( .A1(in_1bar), .A2(inbar[85]), .ZN(n851bar);
  OR2_X1 U110 ( .A1(in_23), .A2(in_19), .ZN(n852) );
  AND2_X1 U110bar ( .A1(in_23bar), .A2(in_19bar), .ZN(n852bar);
  OR2_X1 U111 ( .A1(n850), .A2(n849), .ZN(n854) );
  AND2_X1 U111bar ( .A1(n850bar), .A2(n849bar), .ZN(n854bar);
  OR2_X1 U112 ( .A1(in_43), .A2(in_33), .ZN(n849) );
  AND2_X1 U112bar ( .A1(in_43bar), .A2(in_33bar), .ZN(n849bar);
  OR2_X1 U113 ( .A1(in_63), .A2(in_44), .ZN(n850) );
  AND2_X1 U113bar ( .A1(in_63bar), .A2(in_44bar), .ZN(n850bar);
  OR2_X1 U114 ( .A1(n848), .A2(n847), .ZN(n868) );
  AND2_X1 U114bar ( .A1(n848bar), .A2(n847bar), .ZN(n868bar);
  OR2_X1 U115 ( .A1(in[141]), .A2(in[112]), .ZN(n847) );
  AND2_X1 U115bar ( .A1(inbar[141]), .A2(inbar[112]), .ZN(n847bar);
  OR2_X1 U116 ( .A1(in[147]), .A2(n846), .ZN(n848) );
  AND2_X1 U116bar ( .A1(inbar[147]), .A2(n846bar), .ZN(n848bar);
  OR2_X1 U117 ( .A1(in[181]), .A2(in[167]), .ZN(n846) );
  AND2_X1 U117bar ( .A1(inbar[181]), .A2(inbar[167]), .ZN(n846bar);
  OR2_X1 U118 ( .A1(n845), .A2(n844), .ZN(n870) );
  AND2_X1 U118bar ( .A1(n845bar), .A2(n844bar), .ZN(n870bar);
  OR2_X1 U119 ( .A1(n843), .A2(n842), .ZN(n844) );
  AND2_X1 U119bar ( .A1(n843bar), .A2(n842bar), .ZN(n844bar);
  OR2_X1 U120 ( .A1(in[229]), .A2(in[201]), .ZN(n842) );
  AND2_X1 U120bar ( .A1(inbar[229]), .A2(inbar[201]), .ZN(n842bar);
  OR2_X1 U121 ( .A1(in[237]), .A2(n841), .ZN(n843) );
  AND2_X1 U121bar ( .A1(inbar[237]), .A2(n841bar), .ZN(n843bar);
  OR2_X1 U122 ( .A1(in[94]), .A2(in[253]), .ZN(n841) );
  AND2_X1 U122bar ( .A1(inbar[94]), .A2(inbar[253]), .ZN(n841bar);
  OR2_X1 U123 ( .A1(n840), .A2(n839), .ZN(n845) );
  AND2_X1 U123bar ( .A1(n840bar), .A2(n839bar), .ZN(n845bar);
  OR2_X1 U124 ( .A1(in_21), .A2(in[96]), .ZN(n839) );
  AND2_X1 U124bar ( .A1(in_21bar), .A2(inbar[96]), .ZN(n839bar);
  OR2_X1 U125 ( .A1(in_25), .A2(n838), .ZN(n840) );
  AND2_X1 U125bar ( .A1(in_25bar), .A2(n838bar), .ZN(n840bar);
  OR2_X1 U126 ( .A1(in_81), .A2(in_45), .ZN(n838) );
  AND2_X1 U126bar ( .A1(in_81bar), .A2(in_45bar), .ZN(n838bar);
  OR2_X1 U127 ( .A1(n837), .A2(n836), .ZN(n891) );
  AND2_X1 U127bar ( .A1(n837bar), .A2(n836bar), .ZN(n891bar);
  OR2_X1 U128 ( .A1(in[142]), .A2(in[124]), .ZN(n836) );
  AND2_X1 U128bar ( .A1(inbar[142]), .A2(inbar[124]), .ZN(n836bar);
  OR2_X1 U129 ( .A1(in[150]), .A2(n835), .ZN(n837) );
  AND2_X1 U129bar ( .A1(inbar[150]), .A2(n835bar), .ZN(n837bar);
  OR2_X1 U130 ( .A1(in[172]), .A2(in[155]), .ZN(n835) );
  AND2_X1 U130bar ( .A1(inbar[172]), .A2(inbar[155]), .ZN(n835bar);
  OR2_X1 U131 ( .A1(n834), .A2(n833), .ZN(n893) );
  AND2_X1 U131bar ( .A1(n834bar), .A2(n833bar), .ZN(n893bar);
  OR2_X1 U132 ( .A1(n832), .A2(n831), .ZN(n833) );
  AND2_X1 U132bar ( .A1(n832bar), .A2(n831bar), .ZN(n833bar);
  OR2_X1 U133 ( .A1(in[196]), .A2(in[173]), .ZN(n831) );
  AND2_X1 U133bar ( .A1(inbar[196]), .A2(inbar[173]), .ZN(n831bar);
  OR2_X1 U134 ( .A1(in[222]), .A2(n830), .ZN(n832) );
  AND2_X1 U134bar ( .A1(inbar[222]), .A2(n830bar), .ZN(n832bar);
  OR2_X1 U135 ( .A1(in[227]), .A2(in[226]), .ZN(n830) );
  AND2_X1 U135bar ( .A1(inbar[227]), .A2(inbar[226]), .ZN(n830bar);
  OR2_X1 U136 ( .A1(n829), .A2(n828), .ZN(n834) );
  AND2_X1 U136bar ( .A1(n829bar), .A2(n828bar), .ZN(n834bar);
  OR2_X1 U137 ( .A1(in[249]), .A2(in[231]), .ZN(n828) );
  AND2_X1 U137bar ( .A1(inbar[249]), .A2(inbar[231]), .ZN(n828bar);
  OR2_X1 U138 ( .A1(in_28), .A2(n827), .ZN(n829) );
  AND2_X1 U138bar ( .A1(in_28bar), .A2(n827bar), .ZN(n829bar);
  OR2_X1 U139 ( .A1(in_52), .A2(in_47), .ZN(n827) );
  AND2_X1 U139bar ( .A1(in_52bar), .A2(in_47bar), .ZN(n827bar);
  OR2_X1 U140 ( .A1(n826), .A2(n825), .ZN(out[3]) );
  AND2_X1 U140bar ( .A1(n826bar), .A2(n825bar), .ZN(outbar[3]);
  OR2_X1 U141 ( .A1(n824), .A2(n823), .ZN(n825) );
  AND2_X1 U141bar ( .A1(n824bar), .A2(n823bar), .ZN(n825bar);
  OR2_X1 U142 ( .A1(n822), .A2(n821), .ZN(n823) );
  AND2_X1 U142bar ( .A1(n822bar), .A2(n821bar), .ZN(n823bar);
  OR2_X1 U143 ( .A1(n820), .A2(n819), .ZN(n821) );
  AND2_X1 U143bar ( .A1(n820bar), .A2(n819bar), .ZN(n821bar);
  OR2_X1 U144 ( .A1(n964), .A2(n818), .ZN(n822) );
  AND2_X1 U144bar ( .A1(n964bar), .A2(n818bar), .ZN(n822bar);
  OR2_X1 U145 ( .A1(in[118]), .A2(n817), .ZN(n818) );
  AND2_X1 U145bar ( .A1(inbar[118]), .A2(n817bar), .ZN(n818bar);
  OR2_X1 U146 ( .A1(n816), .A2(n815), .ZN(n964) );
  AND2_X1 U146bar ( .A1(n816bar), .A2(n815bar), .ZN(n964bar);
  OR2_X1 U147 ( .A1(n814), .A2(n813), .ZN(n815) );
  AND2_X1 U147bar ( .A1(n814bar), .A2(n813bar), .ZN(n815bar);
  OR2_X1 U148 ( .A1(n812), .A2(n811), .ZN(n813) );
  AND2_X1 U148bar ( .A1(n812bar), .A2(n811bar), .ZN(n813bar);
  OR2_X1 U149 ( .A1(in[122]), .A2(in[111]), .ZN(n811) );
  AND2_X1 U149bar ( .A1(inbar[122]), .A2(inbar[111]), .ZN(n811bar);
  OR2_X1 U150 ( .A1(in[154]), .A2(in[151]), .ZN(n812) );
  AND2_X1 U150bar ( .A1(inbar[154]), .A2(inbar[151]), .ZN(n812bar);
  OR2_X1 U151 ( .A1(n810), .A2(n809), .ZN(n814) );
  AND2_X1 U151bar ( .A1(n810bar), .A2(n809bar), .ZN(n814bar);
  OR2_X1 U152 ( .A1(in[187]), .A2(in[177]), .ZN(n809) );
  AND2_X1 U152bar ( .A1(inbar[187]), .A2(inbar[177]), .ZN(n809bar);
  OR2_X1 U153 ( .A1(in[200]), .A2(in[192]), .ZN(n810) );
  AND2_X1 U153bar ( .A1(inbar[200]), .A2(inbar[192]), .ZN(n810bar);
  OR2_X1 U154 ( .A1(n808), .A2(n807), .ZN(n816) );
  AND2_X1 U154bar ( .A1(n808bar), .A2(n807bar), .ZN(n816bar);
  OR2_X1 U155 ( .A1(n806), .A2(n805), .ZN(n807) );
  AND2_X1 U155bar ( .A1(n806bar), .A2(n805bar), .ZN(n807bar);
  OR2_X1 U156 ( .A1(in[225]), .A2(in[207]), .ZN(n805) );
  AND2_X1 U156bar ( .A1(inbar[225]), .A2(inbar[207]), .ZN(n805bar);
  OR2_X1 U157 ( .A1(in[98]), .A2(in[226]), .ZN(n806) );
  AND2_X1 U157bar ( .A1(inbar[98]), .A2(inbar[226]), .ZN(n806bar);
  OR2_X1 U158 ( .A1(n804), .A2(n803), .ZN(n808) );
  AND2_X1 U158bar ( .A1(n804bar), .A2(n803bar), .ZN(n808bar);
  OR2_X1 U159 ( .A1(in_20), .A2(in_16), .ZN(n803) );
  AND2_X1 U159bar ( .A1(in_20bar), .A2(in_16bar), .ZN(n803bar);
  OR2_X1 U160 ( .A1(in_55), .A2(in_45), .ZN(n804) );
  AND2_X1 U160bar ( .A1(in_55bar), .A2(in_45bar), .ZN(n804bar);
  OR2_X1 U161 ( .A1(n802), .A2(n801), .ZN(n824) );
  AND2_X1 U161bar ( .A1(n802bar), .A2(n801bar), .ZN(n824bar);
  OR2_X1 U162 ( .A1(in[162]), .A2(in[149]), .ZN(n801) );
  AND2_X1 U162bar ( .A1(inbar[162]), .A2(inbar[149]), .ZN(n801bar);
  OR2_X1 U163 ( .A1(in[163]), .A2(n800), .ZN(n802) );
  AND2_X1 U163bar ( .A1(inbar[163]), .A2(n800bar), .ZN(n802bar);
  OR2_X1 U164 ( .A1(in[191]), .A2(in[189]), .ZN(n800) );
  AND2_X1 U164bar ( .A1(inbar[191]), .A2(inbar[189]), .ZN(n800bar);
  OR2_X1 U165 ( .A1(n799), .A2(n798), .ZN(n826) );
  AND2_X1 U165bar ( .A1(n799bar), .A2(n798bar), .ZN(n826bar);
  OR2_X1 U166 ( .A1(n797), .A2(n796), .ZN(n798) );
  AND2_X1 U166bar ( .A1(n797bar), .A2(n796bar), .ZN(n798bar);
  OR2_X1 U167 ( .A1(in[212]), .A2(in[193]), .ZN(n796) );
  AND2_X1 U167bar ( .A1(inbar[212]), .A2(inbar[193]), .ZN(n796bar);
  OR2_X1 U168 ( .A1(in[238]), .A2(n795), .ZN(n797) );
  AND2_X1 U168bar ( .A1(inbar[238]), .A2(n795bar), .ZN(n797bar);
  OR2_X1 U169 ( .A1(in[88]), .A2(in[247]), .ZN(n795) );
  AND2_X1 U169bar ( .A1(inbar[88]), .A2(inbar[247]), .ZN(n795bar);
  OR2_X1 U170 ( .A1(n794), .A2(n793), .ZN(n799) );
  AND2_X1 U170bar ( .A1(n794bar), .A2(n793bar), .ZN(n799bar);
  OR2_X1 U171 ( .A1(in[94]), .A2(in[92]), .ZN(n793) );
  AND2_X1 U171bar ( .A1(inbar[94]), .A2(inbar[92]), .ZN(n793bar);
  OR2_X1 U172 ( .A1(in_52), .A2(n792), .ZN(n794) );
  AND2_X1 U172bar ( .A1(in_52bar), .A2(n792bar), .ZN(n794bar);
  OR2_X1 U173 ( .A1(in_70), .A2(in_67), .ZN(n792) );
  AND2_X1 U173bar ( .A1(in_70bar), .A2(in_67bar), .ZN(n792bar);
  OR2_X1 U174 ( .A1(n791), .A2(n790), .ZN(out[2]) );
  AND2_X1 U174bar ( .A1(n791bar), .A2(n790bar), .ZN(outbar[2]);
  OR2_X1 U175 ( .A1(n789), .A2(n788), .ZN(n790) );
  AND2_X1 U175bar ( .A1(n789bar), .A2(n788bar), .ZN(n790bar);
  OR2_X1 U176 ( .A1(n787), .A2(n786), .ZN(n788) );
  AND2_X1 U176bar ( .A1(n787bar), .A2(n786bar), .ZN(n788bar);
  OR2_X1 U177 ( .A1(n819), .A2(n785), .ZN(n786) );
  AND2_X1 U177bar ( .A1(n819bar), .A2(n785bar), .ZN(n786bar);
  OR2_X1 U178 ( .A1(n784), .A2(n783), .ZN(n819) );
  AND2_X1 U178bar ( .A1(n784bar), .A2(n783bar), .ZN(n819bar);
  OR2_X1 U179 ( .A1(n782), .A2(n781), .ZN(n783) );
  AND2_X1 U179bar ( .A1(n782bar), .A2(n781bar), .ZN(n783bar);
  OR2_X1 U180 ( .A1(n780), .A2(n779), .ZN(n781) );
  AND2_X1 U180bar ( .A1(n780bar), .A2(n779bar), .ZN(n781bar);
  OR2_X1 U181 ( .A1(n962), .A2(n778), .ZN(n779) );
  AND2_X1 U181bar ( .A1(n962bar), .A2(n778bar), .ZN(n779bar);
  OR2_X1 U182 ( .A1(n777), .A2(n776), .ZN(n962) );
  AND2_X1 U182bar ( .A1(n777bar), .A2(n776bar), .ZN(n962bar);
  OR2_X1 U183 ( .A1(n775), .A2(n774), .ZN(n776) );
  AND2_X1 U183bar ( .A1(n775bar), .A2(n774bar), .ZN(n776bar);
  OR2_X1 U184 ( .A1(n773), .A2(n772), .ZN(n774) );
  AND2_X1 U184bar ( .A1(n773bar), .A2(n772bar), .ZN(n774bar);
  OR2_X1 U185 ( .A1(in[131]), .A2(in[120]), .ZN(n772) );
  AND2_X1 U185bar ( .A1(inbar[131]), .A2(inbar[120]), .ZN(n772bar);
  OR2_X1 U186 ( .A1(in[153]), .A2(in[147]), .ZN(n773) );
  AND2_X1 U186bar ( .A1(inbar[153]), .A2(inbar[147]), .ZN(n773bar);
  OR2_X1 U187 ( .A1(n771), .A2(n770), .ZN(n775) );
  AND2_X1 U187bar ( .A1(n771bar), .A2(n770bar), .ZN(n775bar);
  OR2_X1 U188 ( .A1(in[170]), .A2(in[156]), .ZN(n770) );
  AND2_X1 U188bar ( .A1(inbar[170]), .A2(inbar[156]), .ZN(n770bar);
  OR2_X1 U189 ( .A1(in[223]), .A2(in[190]), .ZN(n771) );
  AND2_X1 U189bar ( .A1(inbar[223]), .A2(inbar[190]), .ZN(n771bar);
  OR2_X1 U190 ( .A1(n769), .A2(n768), .ZN(n777) );
  AND2_X1 U190bar ( .A1(n769bar), .A2(n768bar), .ZN(n777bar);
  OR2_X1 U191 ( .A1(n767), .A2(n766), .ZN(n768) );
  AND2_X1 U191bar ( .A1(n767bar), .A2(n766bar), .ZN(n768bar);
  OR2_X1 U192 ( .A1(in[236]), .A2(in[230]), .ZN(n766) );
  AND2_X1 U192bar ( .A1(inbar[236]), .A2(inbar[230]), .ZN(n766bar);
  OR2_X1 U193 ( .A1(in[85]), .A2(in[240]), .ZN(n767) );
  AND2_X1 U193bar ( .A1(inbar[85]), .A2(inbar[240]), .ZN(n767bar);
  OR2_X1 U194 ( .A1(n765), .A2(n764), .ZN(n769) );
  AND2_X1 U194bar ( .A1(n765bar), .A2(n764bar), .ZN(n769bar);
  OR2_X1 U195 ( .A1(in_12), .A2(in[90]), .ZN(n764) );
  AND2_X1 U195bar ( .A1(in_12bar), .A2(inbar[90]), .ZN(n764bar);
  OR2_X1 U196 ( .A1(in_39), .A2(in_28), .ZN(n765) );
  AND2_X1 U196bar ( .A1(in_39bar), .A2(in_28bar), .ZN(n765bar);
  OR2_X1 U197 ( .A1(in[109]), .A2(n763), .ZN(n780) );
  AND2_X1 U197bar ( .A1(inbar[109]), .A2(n763bar), .ZN(n780bar);
  OR2_X1 U198 ( .A1(n762), .A2(n761), .ZN(n782) );
  AND2_X1 U198bar ( .A1(n762bar), .A2(n761bar), .ZN(n782bar);
  OR2_X1 U199 ( .A1(in[138]), .A2(in[129]), .ZN(n761) );
  AND2_X1 U199bar ( .A1(inbar[138]), .A2(inbar[129]), .ZN(n761bar);
  OR2_X1 U200 ( .A1(in[157]), .A2(n760), .ZN(n762) );
  AND2_X1 U200bar ( .A1(inbar[157]), .A2(n760bar), .ZN(n762bar);
  OR2_X1 U201 ( .A1(in[182]), .A2(in[167]), .ZN(n760) );
  AND2_X1 U201bar ( .A1(inbar[182]), .A2(inbar[167]), .ZN(n760bar);
  OR2_X1 U202 ( .A1(n759), .A2(n758), .ZN(n784) );
  AND2_X1 U202bar ( .A1(n759bar), .A2(n758bar), .ZN(n784bar);
  OR2_X1 U203 ( .A1(n757), .A2(n756), .ZN(n758) );
  AND2_X1 U203bar ( .A1(n757bar), .A2(n756bar), .ZN(n758bar);
  OR2_X1 U204 ( .A1(in[195]), .A2(in[184]), .ZN(n756) );
  AND2_X1 U204bar ( .A1(inbar[195]), .A2(inbar[184]), .ZN(n756bar);
  OR2_X1 U205 ( .A1(in[196]), .A2(n755), .ZN(n757) );
  AND2_X1 U205bar ( .A1(inbar[196]), .A2(n755bar), .ZN(n757bar);
  OR2_X1 U206 ( .A1(in[215]), .A2(in[209]), .ZN(n755) );
  AND2_X1 U206bar ( .A1(inbar[215]), .A2(inbar[209]), .ZN(n755bar);
  OR2_X1 U207 ( .A1(n754), .A2(n753), .ZN(n759) );
  AND2_X1 U207bar ( .A1(n754bar), .A2(n753bar), .ZN(n759bar);
  OR2_X1 U208 ( .A1(in[93]), .A2(in[233]), .ZN(n753) );
  AND2_X1 U208bar ( .A1(inbar[93]), .A2(inbar[233]), .ZN(n753bar);
  OR2_X1 U209 ( .A1(in_1), .A2(n752), .ZN(n754) );
  AND2_X1 U209bar ( .A1(in_1bar), .A2(n752bar), .ZN(n754bar);
  OR2_X1 U210 ( .A1(in_69), .A2(in_66), .ZN(n752) );
  AND2_X1 U210bar ( .A1(in_69bar), .A2(in_66bar), .ZN(n752bar);
  OR2_X1 U211 ( .A1(n966), .A2(n751), .ZN(n787) );
  AND2_X1 U211bar ( .A1(n966bar), .A2(n751bar), .ZN(n787bar);
  OR2_X1 U212 ( .A1(in[134]), .A2(n750), .ZN(n751) );
  AND2_X1 U212bar ( .A1(inbar[134]), .A2(n750bar), .ZN(n751bar);
  OR2_X1 U213 ( .A1(n749), .A2(n748), .ZN(n966) );
  AND2_X1 U213bar ( .A1(n749bar), .A2(n748bar), .ZN(n966bar);
  OR2_X1 U214 ( .A1(n747), .A2(n746), .ZN(n748) );
  AND2_X1 U214bar ( .A1(n747bar), .A2(n746bar), .ZN(n748bar);
  OR2_X1 U215 ( .A1(n745), .A2(n744), .ZN(n746) );
  AND2_X1 U215bar ( .A1(n745bar), .A2(n744bar), .ZN(n746bar);
  OR2_X1 U216 ( .A1(in[136]), .A2(in[121]), .ZN(n744) );
  AND2_X1 U216bar ( .A1(inbar[136]), .A2(inbar[121]), .ZN(n744bar);
  OR2_X1 U217 ( .A1(in[186]), .A2(in[174]), .ZN(n745) );
  AND2_X1 U217bar ( .A1(inbar[186]), .A2(inbar[174]), .ZN(n745bar);
  OR2_X1 U218 ( .A1(n743), .A2(n742), .ZN(n747) );
  AND2_X1 U218bar ( .A1(n743bar), .A2(n742bar), .ZN(n747bar);
  OR2_X1 U219 ( .A1(in[198]), .A2(in[197]), .ZN(n742) );
  AND2_X1 U219bar ( .A1(inbar[198]), .A2(inbar[197]), .ZN(n742bar);
  OR2_X1 U220 ( .A1(in[214]), .A2(in[199]), .ZN(n743) );
  AND2_X1 U220bar ( .A1(inbar[214]), .A2(inbar[199]), .ZN(n743bar);
  OR2_X1 U221 ( .A1(n741), .A2(n740), .ZN(n749) );
  AND2_X1 U221bar ( .A1(n741bar), .A2(n740bar), .ZN(n749bar);
  OR2_X1 U222 ( .A1(n739), .A2(n738), .ZN(n740) );
  AND2_X1 U222bar ( .A1(n739bar), .A2(n738bar), .ZN(n740bar);
  OR2_X1 U223 ( .A1(in[231]), .A2(in[220]), .ZN(n738) );
  AND2_X1 U223bar ( .A1(inbar[231]), .A2(inbar[220]), .ZN(n738bar);
  OR2_X1 U224 ( .A1(in_25), .A2(in[245]), .ZN(n739) );
  AND2_X1 U224bar ( .A1(in_25bar), .A2(inbar[245]), .ZN(n739bar);
  OR2_X1 U225 ( .A1(n737), .A2(n736), .ZN(n741) );
  AND2_X1 U225bar ( .A1(n737bar), .A2(n736bar), .ZN(n741bar);
  OR2_X1 U226 ( .A1(in_53), .A2(in_29), .ZN(n736) );
  AND2_X1 U226bar ( .A1(in_53bar), .A2(in_29bar), .ZN(n736bar);
  OR2_X1 U227 ( .A1(in_79), .A2(in_74), .ZN(n737) );
  AND2_X1 U227bar ( .A1(in_79bar), .A2(in_74bar), .ZN(n737bar);
  OR2_X1 U228 ( .A1(n735), .A2(n734), .ZN(n789) );
  AND2_X1 U228bar ( .A1(n735bar), .A2(n734bar), .ZN(n789bar);
  OR2_X1 U229 ( .A1(in[152]), .A2(in[140]), .ZN(n734) );
  AND2_X1 U229bar ( .A1(inbar[152]), .A2(inbar[140]), .ZN(n734bar);
  OR2_X1 U230 ( .A1(in[155]), .A2(n733), .ZN(n735) );
  AND2_X1 U230bar ( .A1(inbar[155]), .A2(n733bar), .ZN(n735bar);
  OR2_X1 U231 ( .A1(in[166]), .A2(in[165]), .ZN(n733) );
  AND2_X1 U231bar ( .A1(inbar[166]), .A2(inbar[165]), .ZN(n733bar);
  OR2_X1 U232 ( .A1(n732), .A2(n731), .ZN(n791) );
  AND2_X1 U232bar ( .A1(n732bar), .A2(n731bar), .ZN(n791bar);
  OR2_X1 U233 ( .A1(n730), .A2(n729), .ZN(n731) );
  AND2_X1 U233bar ( .A1(n730bar), .A2(n729bar), .ZN(n731bar);
  OR2_X1 U234 ( .A1(in[202]), .A2(in[185]), .ZN(n729) );
  AND2_X1 U234bar ( .A1(inbar[202]), .A2(inbar[185]), .ZN(n729bar);
  OR2_X1 U235 ( .A1(in[211]), .A2(n728), .ZN(n730) );
  AND2_X1 U235bar ( .A1(inbar[211]), .A2(n728bar), .ZN(n730bar);
  OR2_X1 U236 ( .A1(in[255]), .A2(in[253]), .ZN(n728) );
  AND2_X1 U236bar ( .A1(inbar[255]), .A2(inbar[253]), .ZN(n728bar);
  OR2_X1 U237 ( .A1(n727), .A2(n726), .ZN(n732) );
  AND2_X1 U237bar ( .A1(n727bar), .A2(n726bar), .ZN(n732bar);
  OR2_X1 U238 ( .A1(in_35), .A2(in_15), .ZN(n726) );
  AND2_X1 U238bar ( .A1(in_35bar), .A2(in_15bar), .ZN(n726bar);
  OR2_X1 U239 ( .A1(in_36), .A2(n725), .ZN(n727) );
  AND2_X1 U239bar ( .A1(in_36bar), .A2(n725bar), .ZN(n727bar);
  OR2_X1 U240 ( .A1(in_48), .A2(in_40), .ZN(n725) );
  AND2_X1 U240bar ( .A1(in_48bar), .A2(in_40bar), .ZN(n725bar);
  OR2_X1 U241 ( .A1(n724), .A2(n723), .ZN(out[1]) );
  AND2_X1 U241bar ( .A1(n724bar), .A2(n723bar), .ZN(outbar[1]);
  OR2_X1 U242 ( .A1(n722), .A2(n721), .ZN(n723) );
  AND2_X1 U242bar ( .A1(n722bar), .A2(n721bar), .ZN(n723bar);
  OR2_X1 U243 ( .A1(n720), .A2(n719), .ZN(n721) );
  AND2_X1 U243bar ( .A1(n720bar), .A2(n719bar), .ZN(n721bar);
  OR2_X1 U244 ( .A1(n921), .A2(n887), .ZN(n719) );
  AND2_X1 U244bar ( .A1(n921bar), .A2(n887bar), .ZN(n719bar);
  OR2_X1 U245 ( .A1(n718), .A2(n717), .ZN(n887) );
  AND2_X1 U245bar ( .A1(n718bar), .A2(n717bar), .ZN(n887bar);
  OR2_X1 U246 ( .A1(n716), .A2(n715), .ZN(n717) );
  AND2_X1 U246bar ( .A1(n716bar), .A2(n715bar), .ZN(n717bar);
  OR2_X1 U247 ( .A1(n714), .A2(n713), .ZN(n715) );
  AND2_X1 U247bar ( .A1(n714bar), .A2(n713bar), .ZN(n715bar);
  OR2_X1 U248 ( .A1(in[116]), .A2(in[110]), .ZN(n713) );
  AND2_X1 U248bar ( .A1(inbar[116]), .A2(inbar[110]), .ZN(n713bar);
  OR2_X1 U249 ( .A1(in[133]), .A2(in[130]), .ZN(n714) );
  AND2_X1 U249bar ( .A1(inbar[133]), .A2(inbar[130]), .ZN(n714bar);
  OR2_X1 U250 ( .A1(n712), .A2(n711), .ZN(n716) );
  AND2_X1 U250bar ( .A1(n712bar), .A2(n711bar), .ZN(n716bar);
  OR2_X1 U251 ( .A1(in[203]), .A2(in[135]), .ZN(n711) );
  AND2_X1 U251bar ( .A1(inbar[203]), .A2(inbar[135]), .ZN(n711bar);
  OR2_X1 U252 ( .A1(in[232]), .A2(in[223]), .ZN(n712) );
  AND2_X1 U252bar ( .A1(inbar[232]), .A2(inbar[223]), .ZN(n712bar);
  OR2_X1 U253 ( .A1(n710), .A2(n709), .ZN(n718) );
  AND2_X1 U253bar ( .A1(n710bar), .A2(n709bar), .ZN(n718bar);
  OR2_X1 U254 ( .A1(n708), .A2(n707), .ZN(n709) );
  AND2_X1 U254bar ( .A1(n708bar), .A2(n707bar), .ZN(n709bar);
  OR2_X1 U255 ( .A1(in[255]), .A2(in[233]), .ZN(n707) );
  AND2_X1 U255bar ( .A1(inbar[255]), .A2(inbar[233]), .ZN(n707bar);
  OR2_X1 U256 ( .A1(in_53), .A2(in_34), .ZN(n708) );
  AND2_X1 U256bar ( .A1(in_53bar), .A2(in_34bar), .ZN(n708bar);
  OR2_X1 U257 ( .A1(n706), .A2(n705), .ZN(n710) );
  AND2_X1 U257bar ( .A1(n706bar), .A2(n705bar), .ZN(n710bar);
  OR2_X1 U258 ( .A1(in_57), .A2(in_55), .ZN(n705) );
  AND2_X1 U258bar ( .A1(in_57bar), .A2(in_55bar), .ZN(n705bar);
  OR2_X1 U259 ( .A1(in_68), .A2(in_67), .ZN(n706) );
  AND2_X1 U259bar ( .A1(in_68bar), .A2(in_67bar), .ZN(n706bar);
  OR2_X1 U260 ( .A1(n704), .A2(n703), .ZN(n921) );
  AND2_X1 U260bar ( .A1(n704bar), .A2(n703bar), .ZN(n921bar);
  OR2_X1 U261 ( .A1(n702), .A2(n701), .ZN(n703) );
  AND2_X1 U261bar ( .A1(n702bar), .A2(n701bar), .ZN(n703bar);
  OR2_X1 U262 ( .A1(n700), .A2(n699), .ZN(n701) );
  AND2_X1 U262bar ( .A1(n700bar), .A2(n699bar), .ZN(n701bar);
  OR2_X1 U263 ( .A1(n944), .A2(n872), .ZN(n699) );
  AND2_X1 U263bar ( .A1(n944bar), .A2(n872bar), .ZN(n699bar);
  OR2_X1 U264 ( .A1(n698), .A2(n697), .ZN(n872) );
  AND2_X1 U264bar ( .A1(n698bar), .A2(n697bar), .ZN(n872bar);
  OR2_X1 U265 ( .A1(n696), .A2(n695), .ZN(n697) );
  AND2_X1 U265bar ( .A1(n696bar), .A2(n695bar), .ZN(n697bar);
  OR2_X1 U266 ( .A1(n694), .A2(n693), .ZN(n695) );
  AND2_X1 U266bar ( .A1(n694bar), .A2(n693bar), .ZN(n695bar);
  OR2_X1 U267 ( .A1(in[121]), .A2(in[102]), .ZN(n693) );
  AND2_X1 U267bar ( .A1(inbar[121]), .A2(inbar[102]), .ZN(n693bar);
  OR2_X1 U268 ( .A1(in[162]), .A2(in[161]), .ZN(n694) );
  AND2_X1 U268bar ( .A1(inbar[162]), .A2(inbar[161]), .ZN(n694bar);
  OR2_X1 U269 ( .A1(n692), .A2(n691), .ZN(n696) );
  AND2_X1 U269bar ( .A1(n692bar), .A2(n691bar), .ZN(n696bar);
  OR2_X1 U270 ( .A1(in[192]), .A2(in[178]), .ZN(n691) );
  AND2_X1 U270bar ( .A1(inbar[192]), .A2(inbar[178]), .ZN(n691bar);
  OR2_X1 U271 ( .A1(in[244]), .A2(in[209]), .ZN(n692) );
  AND2_X1 U271bar ( .A1(inbar[244]), .A2(inbar[209]), .ZN(n692bar);
  OR2_X1 U272 ( .A1(n690), .A2(n689), .ZN(n698) );
  AND2_X1 U272bar ( .A1(n690bar), .A2(n689bar), .ZN(n698bar);
  OR2_X1 U273 ( .A1(n688), .A2(n687), .ZN(n689) );
  AND2_X1 U273bar ( .A1(n688bar), .A2(n687bar), .ZN(n689bar);
  OR2_X1 U274 ( .A1(in[90]), .A2(in[254]), .ZN(n687) );
  AND2_X1 U274bar ( .A1(inbar[90]), .A2(inbar[254]), .ZN(n687bar);
  OR2_X1 U275 ( .A1(in_36), .A2(in_32), .ZN(n688) );
  AND2_X1 U275bar ( .A1(in_36bar), .A2(in_32bar), .ZN(n688bar);
  OR2_X1 U276 ( .A1(n686), .A2(n685), .ZN(n690) );
  AND2_X1 U276bar ( .A1(n686bar), .A2(n685bar), .ZN(n690bar);
  OR2_X1 U277 ( .A1(in_62), .A2(in_37), .ZN(n685) );
  AND2_X1 U277bar ( .A1(in_62bar), .A2(in_37bar), .ZN(n685bar);
  OR2_X1 U278 ( .A1(in_75), .A2(in_73), .ZN(n686) );
  AND2_X1 U278bar ( .A1(in_75bar), .A2(in_73bar), .ZN(n686bar);
  OR2_X1 U279 ( .A1(n684), .A2(n683), .ZN(n944) );
  AND2_X1 U279bar ( .A1(n684bar), .A2(n683bar), .ZN(n944bar);
  OR2_X1 U280 ( .A1(n682), .A2(n681), .ZN(n683) );
  AND2_X1 U280bar ( .A1(n682bar), .A2(n681bar), .ZN(n683bar);
  OR2_X1 U281 ( .A1(n680), .A2(n679), .ZN(n681) );
  AND2_X1 U281bar ( .A1(n680bar), .A2(n679bar), .ZN(n681bar);
  OR2_X1 U282 ( .A1(in[171]), .A2(in[153]), .ZN(n679) );
  AND2_X1 U282bar ( .A1(inbar[171]), .A2(inbar[153]), .ZN(n679bar);
  OR2_X1 U283 ( .A1(in[187]), .A2(in[176]), .ZN(n680) );
  AND2_X1 U283bar ( .A1(inbar[187]), .A2(inbar[176]), .ZN(n680bar);
  OR2_X1 U284 ( .A1(n678), .A2(n677), .ZN(n682) );
  AND2_X1 U284bar ( .A1(n678bar), .A2(n677bar), .ZN(n682bar);
  OR2_X1 U285 ( .A1(in[245]), .A2(in[211]), .ZN(n677) );
  AND2_X1 U285bar ( .A1(inbar[245]), .A2(inbar[211]), .ZN(n677bar);
  OR2_X1 U286 ( .A1(in[97]), .A2(in[88]), .ZN(n678) );
  AND2_X1 U286bar ( .A1(inbar[97]), .A2(inbar[88]), .ZN(n678bar);
  OR2_X1 U287 ( .A1(n676), .A2(n675), .ZN(n684) );
  AND2_X1 U287bar ( .A1(n676bar), .A2(n675bar), .ZN(n684bar);
  OR2_X1 U288 ( .A1(n674), .A2(n673), .ZN(n675) );
  AND2_X1 U288bar ( .A1(n674bar), .A2(n673bar), .ZN(n675bar);
  OR2_X1 U289 ( .A1(in_10), .A2(in_0), .ZN(n673) );
  AND2_X1 U289bar ( .A1(in_10bar), .A2(in_0bar), .ZN(n673bar);
  OR2_X1 U290 ( .A1(in_59), .A2(in_5), .ZN(n674) );
  AND2_X1 U290bar ( .A1(in_59bar), .A2(in_5bar), .ZN(n674bar);
  OR2_X1 U291 ( .A1(n672), .A2(n671), .ZN(n676) );
  AND2_X1 U291bar ( .A1(n672bar), .A2(n671bar), .ZN(n676bar);
  OR2_X1 U292 ( .A1(in_60), .A2(in_6), .ZN(n671) );
  AND2_X1 U292bar ( .A1(in_60bar), .A2(in_6bar), .ZN(n671bar);
  OR2_X1 U293 ( .A1(in_77), .A2(in_69), .ZN(n672) );
  AND2_X1 U293bar ( .A1(in_77bar), .A2(in_69bar), .ZN(n672bar);
  OR2_X1 U294 ( .A1(in[113]), .A2(n864), .ZN(n700) );
  AND2_X1 U294bar ( .A1(inbar[113]), .A2(n864bar), .ZN(n700bar);
  OR2_X1 U295 ( .A1(n670), .A2(n669), .ZN(n864) );
  AND2_X1 U295bar ( .A1(n670bar), .A2(n669bar), .ZN(n864bar);
  OR2_X1 U296 ( .A1(n668), .A2(n667), .ZN(n669) );
  AND2_X1 U296bar ( .A1(n668bar), .A2(n667bar), .ZN(n669bar);
  OR2_X1 U297 ( .A1(n666), .A2(n665), .ZN(n667) );
  AND2_X1 U297bar ( .A1(n666bar), .A2(n665bar), .ZN(n667bar);
  OR2_X1 U298 ( .A1(in[125]), .A2(in[107]), .ZN(n665) );
  AND2_X1 U298bar ( .A1(inbar[125]), .A2(inbar[107]), .ZN(n665bar);
  OR2_X1 U299 ( .A1(in[138]), .A2(in[126]), .ZN(n666) );
  AND2_X1 U299bar ( .A1(inbar[138]), .A2(inbar[126]), .ZN(n666bar);
  OR2_X1 U300 ( .A1(n664), .A2(n663), .ZN(n668) );
  AND2_X1 U300bar ( .A1(n664bar), .A2(n663bar), .ZN(n668bar);
  OR2_X1 U301 ( .A1(in[189]), .A2(in[143]), .ZN(n663) );
  AND2_X1 U301bar ( .A1(inbar[189]), .A2(inbar[143]), .ZN(n663bar);
  OR2_X1 U302 ( .A1(in[99]), .A2(in[214]), .ZN(n664) );
  AND2_X1 U302bar ( .A1(inbar[99]), .A2(inbar[214]), .ZN(n664bar);
  OR2_X1 U303 ( .A1(n662), .A2(n661), .ZN(n670) );
  AND2_X1 U303bar ( .A1(n662bar), .A2(n661bar), .ZN(n670bar);
  OR2_X1 U304 ( .A1(n660), .A2(n659), .ZN(n661) );
  AND2_X1 U304bar ( .A1(n660bar), .A2(n659bar), .ZN(n661bar);
  OR2_X1 U305 ( .A1(in_15), .A2(in_12), .ZN(n659) );
  AND2_X1 U305bar ( .A1(in_15bar), .A2(in_12bar), .ZN(n659bar);
  OR2_X1 U306 ( .A1(in_20), .A2(in_2), .ZN(n660) );
  AND2_X1 U306bar ( .A1(in_20bar), .A2(in_2bar), .ZN(n660bar);
  OR2_X1 U307 ( .A1(n658), .A2(n657), .ZN(n662) );
  AND2_X1 U307bar ( .A1(n658bar), .A2(n657bar), .ZN(n662bar);
  OR2_X1 U308 ( .A1(in_30), .A2(in_3), .ZN(n657) );
  AND2_X1 U308bar ( .A1(in_30bar), .A2(in_3bar), .ZN(n657bar);
  OR2_X1 U309 ( .A1(in_4), .A2(in_38), .ZN(n658) );
  AND2_X1 U309bar ( .A1(in_4bar), .A2(in_38bar), .ZN(n658bar);
  OR2_X1 U310 ( .A1(n656), .A2(n655), .ZN(n702) );
  AND2_X1 U310bar ( .A1(n656bar), .A2(n655bar), .ZN(n702bar);
  OR2_X1 U311 ( .A1(in[148]), .A2(in[137]), .ZN(n655) );
  AND2_X1 U311bar ( .A1(inbar[148]), .A2(inbar[137]), .ZN(n655bar);
  OR2_X1 U312 ( .A1(in[149]), .A2(n654), .ZN(n656) );
  AND2_X1 U312bar ( .A1(inbar[149]), .A2(n654bar), .ZN(n656bar);
  OR2_X1 U313 ( .A1(in[195]), .A2(in[190]), .ZN(n654) );
  AND2_X1 U313bar ( .A1(inbar[195]), .A2(inbar[190]), .ZN(n654bar);
  OR2_X1 U314 ( .A1(n653), .A2(n652), .ZN(n704) );
  AND2_X1 U314bar ( .A1(n653bar), .A2(n652bar), .ZN(n704bar);
  OR2_X1 U315 ( .A1(n651), .A2(n650), .ZN(n652) );
  AND2_X1 U315bar ( .A1(n651bar), .A2(n650bar), .ZN(n652bar);
  OR2_X1 U316 ( .A1(in[98]), .A2(in[197]), .ZN(n650) );
  AND2_X1 U316bar ( .A1(inbar[98]), .A2(inbar[197]), .ZN(n650bar);
  OR2_X1 U317 ( .A1(in_11), .A2(n649), .ZN(n651) );
  AND2_X1 U317bar ( .A1(in_11bar), .A2(n649bar), .ZN(n651bar);
  OR2_X1 U318 ( .A1(in_26), .A2(in_14), .ZN(n649) );
  AND2_X1 U318bar ( .A1(in_26bar), .A2(in_14bar), .ZN(n649bar);
  OR2_X1 U319 ( .A1(n648), .A2(n647), .ZN(n653) );
  AND2_X1 U319bar ( .A1(n648bar), .A2(n647bar), .ZN(n653bar);
  OR2_X1 U320 ( .A1(in_35), .A2(in_27), .ZN(n647) );
  AND2_X1 U320bar ( .A1(in_35bar), .A2(in_27bar), .ZN(n647bar);
  OR2_X1 U321 ( .A1(in_50), .A2(n646), .ZN(n648) );
  AND2_X1 U321bar ( .A1(in_50bar), .A2(n646bar), .ZN(n648bar);
  OR2_X1 U322 ( .A1(in_78), .A2(in_61), .ZN(n646) );
  AND2_X1 U322bar ( .A1(in_78bar), .A2(in_61bar), .ZN(n646bar);
  OR2_X1 U323 ( .A1(n942), .A2(n645), .ZN(n720) );
  AND2_X1 U323bar ( .A1(n942bar), .A2(n645bar), .ZN(n720bar);
  OR2_X1 U324 ( .A1(in[106]), .A2(n863), .ZN(n645) );
  AND2_X1 U324bar ( .A1(inbar[106]), .A2(n863bar), .ZN(n645bar);
  OR2_X1 U325 ( .A1(n644), .A2(n643), .ZN(n863) );
  AND2_X1 U325bar ( .A1(n644bar), .A2(n643bar), .ZN(n863bar);
  OR2_X1 U326 ( .A1(n642), .A2(n641), .ZN(n643) );
  AND2_X1 U326bar ( .A1(n642bar), .A2(n641bar), .ZN(n643bar);
  OR2_X1 U327 ( .A1(n640), .A2(n639), .ZN(n641) );
  AND2_X1 U327bar ( .A1(n640bar), .A2(n639bar), .ZN(n641bar);
  OR2_X1 U328 ( .A1(in[127]), .A2(in[122]), .ZN(n639) );
  AND2_X1 U328bar ( .A1(inbar[127]), .A2(inbar[122]), .ZN(n639bar);
  OR2_X1 U329 ( .A1(in[156]), .A2(in[132]), .ZN(n640) );
  AND2_X1 U329bar ( .A1(inbar[156]), .A2(inbar[132]), .ZN(n640bar);
  OR2_X1 U330 ( .A1(n638), .A2(n637), .ZN(n642) );
  AND2_X1 U330bar ( .A1(n638bar), .A2(n637bar), .ZN(n642bar);
  OR2_X1 U331 ( .A1(in[159]), .A2(in[157]), .ZN(n637) );
  AND2_X1 U331bar ( .A1(inbar[159]), .A2(inbar[157]), .ZN(n637bar);
  OR2_X1 U332 ( .A1(in[185]), .A2(in[169]), .ZN(n638) );
  AND2_X1 U332bar ( .A1(inbar[185]), .A2(inbar[169]), .ZN(n638bar);
  OR2_X1 U333 ( .A1(n636), .A2(n635), .ZN(n644) );
  AND2_X1 U333bar ( .A1(n636bar), .A2(n635bar), .ZN(n644bar);
  OR2_X1 U334 ( .A1(n634), .A2(n633), .ZN(n635) );
  AND2_X1 U334bar ( .A1(n634bar), .A2(n633bar), .ZN(n635bar);
  OR2_X1 U335 ( .A1(in[239]), .A2(in[218]), .ZN(n633) );
  AND2_X1 U335bar ( .A1(inbar[239]), .A2(inbar[218]), .ZN(n633bar);
  OR2_X1 U336 ( .A1(in_13), .A2(in[87]), .ZN(n634) );
  AND2_X1 U336bar ( .A1(in_13bar), .A2(inbar[87]), .ZN(n634bar);
  OR2_X1 U337 ( .A1(n632), .A2(n631), .ZN(n636) );
  AND2_X1 U337bar ( .A1(n632bar), .A2(n631bar), .ZN(n636bar);
  OR2_X1 U338 ( .A1(in_72), .A2(in_70), .ZN(n631) );
  AND2_X1 U338bar ( .A1(in_72bar), .A2(in_70bar), .ZN(n631bar);
  OR2_X1 U339 ( .A1(in_80), .A2(in_74), .ZN(n632) );
  AND2_X1 U339bar ( .A1(in_80bar), .A2(in_74bar), .ZN(n632bar);
  OR2_X1 U340 ( .A1(n630), .A2(n629), .ZN(n942) );
  AND2_X1 U340bar ( .A1(n630bar), .A2(n629bar), .ZN(n942bar);
  OR2_X1 U341 ( .A1(n628), .A2(n627), .ZN(n629) );
  AND2_X1 U341bar ( .A1(n628bar), .A2(n627bar), .ZN(n629bar);
  OR2_X1 U342 ( .A1(n626), .A2(n625), .ZN(n627) );
  AND2_X1 U342bar ( .A1(n626bar), .A2(n625bar), .ZN(n627bar);
  OR2_X1 U343 ( .A1(in[146]), .A2(in[100]), .ZN(n625) );
  AND2_X1 U343bar ( .A1(inbar[146]), .A2(inbar[100]), .ZN(n625bar);
  OR2_X1 U344 ( .A1(in[168]), .A2(in[152]), .ZN(n626) );
  AND2_X1 U344bar ( .A1(inbar[168]), .A2(inbar[152]), .ZN(n626bar);
  OR2_X1 U345 ( .A1(n624), .A2(n623), .ZN(n628) );
  AND2_X1 U345bar ( .A1(n624bar), .A2(n623bar), .ZN(n628bar);
  OR2_X1 U346 ( .A1(in[199]), .A2(in[182]), .ZN(n623) );
  AND2_X1 U346bar ( .A1(inbar[199]), .A2(inbar[182]), .ZN(n623bar);
  OR2_X1 U347 ( .A1(in[236]), .A2(in[204]), .ZN(n624) );
  AND2_X1 U347bar ( .A1(inbar[236]), .A2(inbar[204]), .ZN(n624bar);
  OR2_X1 U348 ( .A1(n622), .A2(n621), .ZN(n630) );
  AND2_X1 U348bar ( .A1(n622bar), .A2(n621bar), .ZN(n630bar);
  OR2_X1 U349 ( .A1(n620), .A2(n619), .ZN(n621) );
  AND2_X1 U349bar ( .A1(n620bar), .A2(n619bar), .ZN(n621bar);
  OR2_X1 U350 ( .A1(in[89]), .A2(in[246]), .ZN(n619) );
  AND2_X1 U350bar ( .A1(inbar[89]), .A2(inbar[246]), .ZN(n619bar);
  OR2_X1 U351 ( .A1(in[95]), .A2(in[92]), .ZN(n620) );
  AND2_X1 U351bar ( .A1(inbar[95]), .A2(inbar[92]), .ZN(n620bar);
  OR2_X1 U352 ( .A1(n618), .A2(n617), .ZN(n622) );
  AND2_X1 U352bar ( .A1(n618bar), .A2(n617bar), .ZN(n622bar);
  OR2_X1 U353 ( .A1(in_22), .A2(in_16), .ZN(n617) );
  AND2_X1 U353bar ( .A1(in_22bar), .A2(in_16bar), .ZN(n617bar);
  OR2_X1 U354 ( .A1(in_51), .A2(in_49), .ZN(n618) );
  AND2_X1 U354bar ( .A1(in_51bar), .A2(in_49bar), .ZN(n618bar);
  OR2_X1 U355 ( .A1(n616), .A2(n615), .ZN(n722) );
  AND2_X1 U355bar ( .A1(n616bar), .A2(n615bar), .ZN(n722bar);
  OR2_X1 U356 ( .A1(in[158]), .A2(in[115]), .ZN(n615) );
  AND2_X1 U356bar ( .A1(inbar[158]), .A2(inbar[115]), .ZN(n615bar);
  OR2_X1 U357 ( .A1(in[163]), .A2(n614), .ZN(n616) );
  AND2_X1 U357bar ( .A1(inbar[163]), .A2(n614bar), .ZN(n616bar);
  OR2_X1 U358 ( .A1(in[206]), .A2(in[165]), .ZN(n614) );
  AND2_X1 U358bar ( .A1(inbar[206]), .A2(inbar[165]), .ZN(n614bar);
  OR2_X1 U359 ( .A1(n613), .A2(n612), .ZN(n724) );
  AND2_X1 U359bar ( .A1(n613bar), .A2(n612bar), .ZN(n724bar);
  OR2_X1 U360 ( .A1(n611), .A2(n610), .ZN(n612) );
  AND2_X1 U360bar ( .A1(n611bar), .A2(n610bar), .ZN(n612bar);
  OR2_X1 U361 ( .A1(in[213]), .A2(in[207]), .ZN(n610) );
  AND2_X1 U361bar ( .A1(inbar[213]), .A2(inbar[207]), .ZN(n610bar);
  OR2_X1 U362 ( .A1(in[215]), .A2(n609), .ZN(n611) );
  AND2_X1 U362bar ( .A1(inbar[215]), .A2(n609bar), .ZN(n611bar);
  OR2_X1 U363 ( .A1(in[230]), .A2(in[220]), .ZN(n609) );
  AND2_X1 U363bar ( .A1(inbar[230]), .A2(inbar[220]), .ZN(n609bar);
  OR2_X1 U364 ( .A1(n608), .A2(n607), .ZN(n613) );
  AND2_X1 U364bar ( .A1(n608bar), .A2(n607bar), .ZN(n613bar);
  OR2_X1 U365 ( .A1(in[251]), .A2(in[234]), .ZN(n607) );
  AND2_X1 U365bar ( .A1(inbar[251]), .A2(inbar[234]), .ZN(n607bar);
  OR2_X1 U366 ( .A1(in_17), .A2(n606), .ZN(n608) );
  AND2_X1 U366bar ( .A1(in_17bar), .A2(n606bar), .ZN(n608bar);
  OR2_X1 U367 ( .A1(in_65), .A2(in_56), .ZN(n606) );
  AND2_X1 U367bar ( .A1(in_65bar), .A2(in_56bar), .ZN(n606bar);
  OR2_X1 U368 ( .A1(n605), .A2(n604), .ZN(out[0]) );
  AND2_X1 U368bar ( .A1(n605bar), .A2(n604bar), .ZN(outbar[0]);
  OR2_X1 U369 ( .A1(n603), .A2(n602), .ZN(n604) );
  AND2_X1 U369bar ( .A1(n603bar), .A2(n602bar), .ZN(n604bar);
  OR2_X1 U370 ( .A1(n601), .A2(n600), .ZN(n602) );
  AND2_X1 U370bar ( .A1(n601bar), .A2(n600bar), .ZN(n602bar);
  OR2_X1 U371 ( .A1(n820), .A2(n785), .ZN(n600) );
  AND2_X1 U371bar ( .A1(n820bar), .A2(n785bar), .ZN(n600bar);
  OR2_X1 U372 ( .A1(n599), .A2(n598), .ZN(n785) );
  AND2_X1 U372bar ( .A1(n599bar), .A2(n598bar), .ZN(n785bar);
  OR2_X1 U373 ( .A1(n597), .A2(n596), .ZN(n598) );
  AND2_X1 U373bar ( .A1(n597bar), .A2(n596bar), .ZN(n598bar);
  OR2_X1 U374 ( .A1(n595), .A2(n594), .ZN(n596) );
  AND2_X1 U374bar ( .A1(n595bar), .A2(n594bar), .ZN(n596bar);
  OR2_X1 U375 ( .A1(in[135]), .A2(in[104]), .ZN(n594) );
  AND2_X1 U375bar ( .A1(inbar[135]), .A2(inbar[104]), .ZN(n594bar);
  OR2_X1 U376 ( .A1(in[188]), .A2(in[178]), .ZN(n595) );
  AND2_X1 U376bar ( .A1(inbar[188]), .A2(inbar[178]), .ZN(n595bar);
  OR2_X1 U377 ( .A1(n593), .A2(n592), .ZN(n597) );
  AND2_X1 U377bar ( .A1(n593bar), .A2(n592bar), .ZN(n597bar);
  OR2_X1 U378 ( .A1(in[217]), .A2(in[194]), .ZN(n592) );
  AND2_X1 U378bar ( .A1(inbar[217]), .A2(inbar[194]), .ZN(n592bar);
  OR2_X1 U379 ( .A1(in[237]), .A2(in[218]), .ZN(n593) );
  AND2_X1 U379bar ( .A1(inbar[237]), .A2(inbar[218]), .ZN(n593bar);
  OR2_X1 U380 ( .A1(n591), .A2(n590), .ZN(n599) );
  AND2_X1 U380bar ( .A1(n591bar), .A2(n590bar), .ZN(n599bar);
  OR2_X1 U381 ( .A1(n589), .A2(n588), .ZN(n590) );
  AND2_X1 U381bar ( .A1(n589bar), .A2(n588bar), .ZN(n590bar);
  OR2_X1 U382 ( .A1(in_2), .A2(in_10), .ZN(n588) );
  AND2_X1 U382bar ( .A1(in_2bar), .A2(in_10bar), .ZN(n588bar);
  OR2_X1 U383 ( .A1(in_47), .A2(in_22), .ZN(n589) );
  AND2_X1 U383bar ( .A1(in_47bar), .A2(in_22bar), .ZN(n589bar);
  OR2_X1 U384 ( .A1(n587), .A2(n586), .ZN(n591) );
  AND2_X1 U384bar ( .A1(n587bar), .A2(n586bar), .ZN(n591bar);
  OR2_X1 U385 ( .A1(in_56), .A2(in_54), .ZN(n586) );
  AND2_X1 U385bar ( .A1(in_56bar), .A2(in_54bar), .ZN(n586bar);
  OR2_X1 U386 ( .A1(in_63), .A2(in_61), .ZN(n587) );
  AND2_X1 U386bar ( .A1(in_63bar), .A2(in_61bar), .ZN(n587bar);
  OR2_X1 U387 ( .A1(n585), .A2(n584), .ZN(n820) );
  AND2_X1 U387bar ( .A1(n585bar), .A2(n584bar), .ZN(n820bar);
  OR2_X1 U388 ( .A1(n583), .A2(n582), .ZN(n584) );
  AND2_X1 U388bar ( .A1(n583bar), .A2(n582bar), .ZN(n584bar);
  OR2_X1 U389 ( .A1(n581), .A2(n580), .ZN(n582) );
  AND2_X1 U389bar ( .A1(n581bar), .A2(n580bar), .ZN(n582bar);
  OR2_X1 U390 ( .A1(in[158]), .A2(in[142]), .ZN(n580) );
  AND2_X1 U390bar ( .A1(inbar[158]), .A2(inbar[142]), .ZN(n580bar);
  OR2_X1 U391 ( .A1(in[175]), .A2(in[164]), .ZN(n581) );
  AND2_X1 U391bar ( .A1(inbar[175]), .A2(inbar[164]), .ZN(n581bar);
  OR2_X1 U392 ( .A1(n579), .A2(n578), .ZN(n583) );
  AND2_X1 U392bar ( .A1(n579bar), .A2(n578bar), .ZN(n583bar);
  OR2_X1 U393 ( .A1(in[228]), .A2(in[204]), .ZN(n578) );
  AND2_X1 U393bar ( .A1(inbar[228]), .A2(inbar[204]), .ZN(n578bar);
  OR2_X1 U394 ( .A1(in[91]), .A2(in[87]), .ZN(n579) );
  AND2_X1 U394bar ( .A1(inbar[91]), .A2(inbar[87]), .ZN(n579bar);
  OR2_X1 U395 ( .A1(n577), .A2(n576), .ZN(n585) );
  AND2_X1 U395bar ( .A1(n577bar), .A2(n576bar), .ZN(n585bar);
  OR2_X1 U396 ( .A1(n575), .A2(n574), .ZN(n576) );
  AND2_X1 U396bar ( .A1(n575bar), .A2(n574bar), .ZN(n576bar);
  OR2_X1 U397 ( .A1(in_21), .A2(in_11), .ZN(n574) );
  AND2_X1 U397bar ( .A1(in_21bar), .A2(in_11bar), .ZN(n574bar);
  OR2_X1 U398 ( .A1(in_5), .A2(in_3), .ZN(n575) );
  AND2_X1 U398bar ( .A1(in_5bar), .A2(in_3bar), .ZN(n575bar);
  OR2_X1 U399 ( .A1(n573), .A2(n572), .ZN(n577) );
  AND2_X1 U399bar ( .A1(n573bar), .A2(n572bar), .ZN(n577bar);
  OR2_X1 U400 ( .A1(in_68), .A2(in_64), .ZN(n572) );
  AND2_X1 U400bar ( .A1(in_68bar), .A2(in_64bar), .ZN(n572bar);
  OR2_X1 U401 ( .A1(in_76), .A2(in_73), .ZN(n573) );
  AND2_X1 U401bar ( .A1(in_76bar), .A2(in_73bar), .ZN(n573bar);
  OR2_X1 U402 ( .A1(n778), .A2(n571), .ZN(n601) );
  AND2_X1 U402bar ( .A1(n778bar), .A2(n571bar), .ZN(n601bar);
  OR2_X1 U403 ( .A1(in[100]), .A2(n965), .ZN(n571) );
  AND2_X1 U403bar ( .A1(inbar[100]), .A2(n965bar), .ZN(n571bar);
  OR2_X1 U404 ( .A1(n570), .A2(n569), .ZN(n965) );
  AND2_X1 U404bar ( .A1(n570bar), .A2(n569bar), .ZN(n965bar);
  OR2_X1 U405 ( .A1(n568), .A2(n567), .ZN(n569) );
  AND2_X1 U405bar ( .A1(n568bar), .A2(n567bar), .ZN(n569bar);
  OR2_X1 U406 ( .A1(n566), .A2(n565), .ZN(n567) );
  AND2_X1 U406bar ( .A1(n566bar), .A2(n565bar), .ZN(n567bar);
  OR2_X1 U407 ( .A1(n817), .A2(n750), .ZN(n565) );
  AND2_X1 U407bar ( .A1(n817bar), .A2(n750bar), .ZN(n565bar);
  OR2_X1 U408 ( .A1(n564), .A2(n563), .ZN(n750) );
  AND2_X1 U408bar ( .A1(n564bar), .A2(n563bar), .ZN(n750bar);
  OR2_X1 U409 ( .A1(n562), .A2(n561), .ZN(n563) );
  AND2_X1 U409bar ( .A1(n562bar), .A2(n561bar), .ZN(n563bar);
  OR2_X1 U410 ( .A1(n560), .A2(n559), .ZN(n561) );
  AND2_X1 U410bar ( .A1(n560bar), .A2(n559bar), .ZN(n561bar);
  OR2_X1 U411 ( .A1(in[119]), .A2(in[103]), .ZN(n559) );
  AND2_X1 U411bar ( .A1(inbar[119]), .A2(inbar[103]), .ZN(n559bar);
  OR2_X1 U412 ( .A1(in[137]), .A2(in[133]), .ZN(n560) );
  AND2_X1 U412bar ( .A1(inbar[137]), .A2(inbar[133]), .ZN(n560bar);
  OR2_X1 U413 ( .A1(n558), .A2(n557), .ZN(n562) );
  AND2_X1 U413bar ( .A1(n558bar), .A2(n557bar), .ZN(n562bar);
  OR2_X1 U414 ( .A1(in[176]), .A2(in[173]), .ZN(n557) );
  AND2_X1 U414bar ( .A1(inbar[176]), .A2(inbar[173]), .ZN(n557bar);
  OR2_X1 U415 ( .A1(in[210]), .A2(in[181]), .ZN(n558) );
  AND2_X1 U415bar ( .A1(inbar[210]), .A2(inbar[181]), .ZN(n558bar);
  OR2_X1 U416 ( .A1(n556), .A2(n555), .ZN(n564) );
  AND2_X1 U416bar ( .A1(n556bar), .A2(n555bar), .ZN(n564bar);
  OR2_X1 U417 ( .A1(n554), .A2(n553), .ZN(n555) );
  AND2_X1 U417bar ( .A1(n554bar), .A2(n553bar), .ZN(n555bar);
  OR2_X1 U418 ( .A1(in_13), .A2(in[234]), .ZN(n553) );
  AND2_X1 U418bar ( .A1(in_13bar), .A2(inbar[234]), .ZN(n553bar);
  OR2_X1 U419 ( .A1(in_38), .A2(in_32), .ZN(n554) );
  AND2_X1 U419bar ( .A1(in_38bar), .A2(in_32bar), .ZN(n554bar);
  OR2_X1 U420 ( .A1(n552), .A2(n551), .ZN(n556) );
  AND2_X1 U420bar ( .A1(n552bar), .A2(n551bar), .ZN(n556bar);
  OR2_X1 U421 ( .A1(in_42), .A2(in_41), .ZN(n551) );
  AND2_X1 U421bar ( .A1(in_42bar), .A2(in_41bar), .ZN(n551bar);
  OR2_X1 U422 ( .A1(in_7), .A2(in_49), .ZN(n552) );
  AND2_X1 U422bar ( .A1(in_7bar), .A2(in_49bar), .ZN(n552bar);
  OR2_X1 U423 ( .A1(n550), .A2(n549), .ZN(n817) );
  AND2_X1 U423bar ( .A1(n550bar), .A2(n549bar), .ZN(n817bar);
  OR2_X1 U424 ( .A1(n548), .A2(n547), .ZN(n549) );
  AND2_X1 U424bar ( .A1(n548bar), .A2(n547bar), .ZN(n549bar);
  OR2_X1 U425 ( .A1(n546), .A2(n545), .ZN(n547) );
  AND2_X1 U425bar ( .A1(n546bar), .A2(n545bar), .ZN(n547bar);
  OR2_X1 U426 ( .A1(in[159]), .A2(in[105]), .ZN(n545) );
  AND2_X1 U426bar ( .A1(inbar[159]), .A2(inbar[105]), .ZN(n545bar);
  OR2_X1 U427 ( .A1(in[206]), .A2(in[183]), .ZN(n546) );
  AND2_X1 U427bar ( .A1(inbar[206]), .A2(inbar[183]), .ZN(n546bar);
  OR2_X1 U428 ( .A1(n544), .A2(n543), .ZN(n548) );
  AND2_X1 U428bar ( .A1(n544bar), .A2(n543bar), .ZN(n548bar);
  OR2_X1 U429 ( .A1(in[229]), .A2(in[219]), .ZN(n543) );
  AND2_X1 U429bar ( .A1(inbar[229]), .A2(inbar[219]), .ZN(n543bar);
  OR2_X1 U430 ( .A1(in[235]), .A2(in[232]), .ZN(n544) );
  AND2_X1 U430bar ( .A1(inbar[235]), .A2(inbar[232]), .ZN(n544bar);
  OR2_X1 U431 ( .A1(n542), .A2(n541), .ZN(n550) );
  AND2_X1 U431bar ( .A1(n542bar), .A2(n541bar), .ZN(n550bar);
  OR2_X1 U432 ( .A1(n540), .A2(n539), .ZN(n541) );
  AND2_X1 U432bar ( .A1(n540bar), .A2(n539bar), .ZN(n541bar);
  OR2_X1 U433 ( .A1(in[249]), .A2(in[242]), .ZN(n539) );
  AND2_X1 U433bar ( .A1(inbar[249]), .A2(inbar[242]), .ZN(n539bar);
  OR2_X1 U434 ( .A1(in[89]), .A2(in[254]), .ZN(n540) );
  AND2_X1 U434bar ( .A1(inbar[89]), .A2(inbar[254]), .ZN(n540bar);
  OR2_X1 U435 ( .A1(n538), .A2(n537), .ZN(n542) );
  AND2_X1 U435bar ( .A1(n538bar), .A2(n537bar), .ZN(n542bar);
  OR2_X1 U436 ( .A1(in_14), .A2(in[99]), .ZN(n537) );
  AND2_X1 U436bar ( .A1(in_14bar), .A2(inbar[99]), .ZN(n537bar);
  OR2_X1 U437 ( .A1(in_60), .A2(in_18), .ZN(n538) );
  AND2_X1 U437bar ( .A1(in_60bar), .A2(in_18bar), .ZN(n538bar);
  OR2_X1 U438 ( .A1(in[113]), .A2(n763), .ZN(n566) );
  AND2_X1 U438bar ( .A1(inbar[113]), .A2(n763bar), .ZN(n566bar);
  OR2_X1 U439 ( .A1(n536), .A2(n535), .ZN(n763) );
  AND2_X1 U439bar ( .A1(n536bar), .A2(n535bar), .ZN(n763bar);
  OR2_X1 U440 ( .A1(n534), .A2(n533), .ZN(n535) );
  AND2_X1 U440bar ( .A1(n534bar), .A2(n533bar), .ZN(n535bar);
  OR2_X1 U441 ( .A1(n532), .A2(n531), .ZN(n533) );
  AND2_X1 U441bar ( .A1(n532bar), .A2(n531bar), .ZN(n533bar);
  OR2_X1 U442 ( .A1(in[115]), .A2(in[110]), .ZN(n531) );
  AND2_X1 U442bar ( .A1(inbar[115]), .A2(inbar[110]), .ZN(n531bar);
  OR2_X1 U443 ( .A1(in[125]), .A2(in[117]), .ZN(n532) );
  AND2_X1 U443bar ( .A1(inbar[125]), .A2(inbar[117]), .ZN(n532bar);
  OR2_X1 U444 ( .A1(n530), .A2(n529), .ZN(n534) );
  AND2_X1 U444bar ( .A1(n530bar), .A2(n529bar), .ZN(n534bar);
  OR2_X1 U445 ( .A1(in[180]), .A2(in[128]), .ZN(n529) );
  AND2_X1 U445bar ( .A1(inbar[180]), .A2(inbar[128]), .ZN(n529bar);
  OR2_X1 U446 ( .A1(in[205]), .A2(in[201]), .ZN(n530) );
  AND2_X1 U446bar ( .A1(inbar[205]), .A2(inbar[201]), .ZN(n530bar);
  OR2_X1 U447 ( .A1(n528), .A2(n527), .ZN(n536) );
  AND2_X1 U447bar ( .A1(n528bar), .A2(n527bar), .ZN(n536bar);
  OR2_X1 U448 ( .A1(n526), .A2(n525), .ZN(n527) );
  AND2_X1 U448bar ( .A1(n526bar), .A2(n525bar), .ZN(n527bar);
  OR2_X1 U449 ( .A1(in[244]), .A2(in[239]), .ZN(n525) );
  AND2_X1 U449bar ( .A1(inbar[244]), .A2(inbar[239]), .ZN(n525bar);
  OR2_X1 U450 ( .A1(in[95]), .A2(in[83]), .ZN(n526) );
  AND2_X1 U450bar ( .A1(inbar[95]), .A2(inbar[83]), .ZN(n526bar);
  OR2_X1 U451 ( .A1(n524), .A2(n523), .ZN(n528) );
  AND2_X1 U451bar ( .A1(n524bar), .A2(n523bar), .ZN(n528bar);
  OR2_X1 U452 ( .A1(in_24), .A2(in[97]), .ZN(n523) );
  AND2_X1 U452bar ( .A1(in_24bar), .A2(inbar[97]), .ZN(n523bar);
  OR2_X1 U453 ( .A1(in_33), .A2(in_27), .ZN(n524) );
  AND2_X1 U453bar ( .A1(in_33bar), .A2(in_27bar), .ZN(n524bar);
  OR2_X1 U454 ( .A1(n522), .A2(n521), .ZN(n568) );
  AND2_X1 U454bar ( .A1(n522bar), .A2(n521bar), .ZN(n568bar);
  OR2_X1 U455 ( .A1(in[145]), .A2(in[126]), .ZN(n521) );
  AND2_X1 U455bar ( .A1(inbar[145]), .A2(inbar[126]), .ZN(n521bar);
  OR2_X1 U456 ( .A1(in[169]), .A2(n520), .ZN(n522) );
  AND2_X1 U456bar ( .A1(inbar[169]), .A2(n520bar), .ZN(n522bar);
  OR2_X1 U457 ( .A1(in[221]), .A2(in[172]), .ZN(n520) );
  AND2_X1 U457bar ( .A1(inbar[221]), .A2(inbar[172]), .ZN(n520bar);
  OR2_X1 U458 ( .A1(n519), .A2(n518), .ZN(n570) );
  AND2_X1 U458bar ( .A1(n519bar), .A2(n518bar), .ZN(n570bar);
  OR2_X1 U459 ( .A1(n517), .A2(n516), .ZN(n518) );
  AND2_X1 U459bar ( .A1(n517bar), .A2(n516bar), .ZN(n518bar);
  OR2_X1 U460 ( .A1(in[241]), .A2(in[224]), .ZN(n516) );
  AND2_X1 U460bar ( .A1(inbar[241]), .A2(inbar[224]), .ZN(n516bar);
  OR2_X1 U461 ( .A1(in[86]), .A2(n515), .ZN(n517) );
  AND2_X1 U461bar ( .A1(inbar[86]), .A2(n515bar), .ZN(n517bar);
  OR2_X1 U462 ( .A1(in_43), .A2(in_34), .ZN(n515) );
  AND2_X1 U462bar ( .A1(in_43bar), .A2(in_34bar), .ZN(n515bar);
  OR2_X1 U463 ( .A1(n514), .A2(n513), .ZN(n519) );
  AND2_X1 U463bar ( .A1(n514bar), .A2(n513bar), .ZN(n519bar);
  OR2_X1 U464 ( .A1(in_65), .A2(in_51), .ZN(n513) );
  AND2_X1 U464bar ( .A1(in_65bar), .A2(in_51bar), .ZN(n513bar);
  OR2_X1 U465 ( .A1(in_75), .A2(n512), .ZN(n514) );
  AND2_X1 U465bar ( .A1(in_75bar), .A2(n512bar), .ZN(n514bar);
  OR2_X1 U466 ( .A1(in_81), .A2(in_77), .ZN(n512) );
  AND2_X1 U466bar ( .A1(in_81bar), .A2(in_77bar), .ZN(n512bar);
  OR2_X1 U467 ( .A1(n511), .A2(n510), .ZN(n778) );
  AND2_X1 U467bar ( .A1(n511bar), .A2(n510bar), .ZN(n778bar);
  OR2_X1 U468 ( .A1(n509), .A2(n508), .ZN(n510) );
  AND2_X1 U468bar ( .A1(n509bar), .A2(n508bar), .ZN(n510bar);
  OR2_X1 U469 ( .A1(n507), .A2(n506), .ZN(n508) );
  AND2_X1 U469bar ( .A1(n507bar), .A2(n506bar), .ZN(n508bar);
  OR2_X1 U470 ( .A1(in[107]), .A2(in[101]), .ZN(n506) );
  AND2_X1 U470bar ( .A1(inbar[107]), .A2(inbar[101]), .ZN(n506bar);
  OR2_X1 U471 ( .A1(in[139]), .A2(in[132]), .ZN(n507) );
  AND2_X1 U471bar ( .A1(inbar[139]), .A2(inbar[132]), .ZN(n507bar);
  OR2_X1 U472 ( .A1(n505), .A2(n504), .ZN(n509) );
  AND2_X1 U472bar ( .A1(n505bar), .A2(n504bar), .ZN(n509bar);
  OR2_X1 U473 ( .A1(in[146]), .A2(in[141]), .ZN(n504) );
  AND2_X1 U473bar ( .A1(inbar[146]), .A2(inbar[141]), .ZN(n504bar);
  OR2_X1 U474 ( .A1(in[203]), .A2(in[179]), .ZN(n505) );
  AND2_X1 U474bar ( .A1(inbar[203]), .A2(inbar[179]), .ZN(n505bar);
  OR2_X1 U475 ( .A1(n503), .A2(n502), .ZN(n511) );
  AND2_X1 U475bar ( .A1(n503bar), .A2(n502bar), .ZN(n511bar);
  OR2_X1 U476 ( .A1(n501), .A2(n500), .ZN(n502) );
  AND2_X1 U476bar ( .A1(n501bar), .A2(n500bar), .ZN(n502bar);
  OR2_X1 U477 ( .A1(in[243]), .A2(in[222]), .ZN(n500) );
  AND2_X1 U477bar ( .A1(inbar[243]), .A2(inbar[222]), .ZN(n500bar);
  OR2_X1 U478 ( .A1(in[251]), .A2(in[250]), .ZN(n501) );
  AND2_X1 U478bar ( .A1(inbar[251]), .A2(inbar[250]), .ZN(n501bar);
  OR2_X1 U479 ( .A1(n499), .A2(n498), .ZN(n503) );
  AND2_X1 U479bar ( .A1(n499bar), .A2(n498bar), .ZN(n503bar);
  OR2_X1 U480 ( .A1(in_37), .A2(in_19), .ZN(n498) );
  AND2_X1 U480bar ( .A1(in_37bar), .A2(in_19bar), .ZN(n498bar);
  OR2_X1 U481 ( .A1(in_78), .A2(in_6), .ZN(n499) );
  AND2_X1 U481bar ( .A1(in_78bar), .A2(in_6bar), .ZN(n499bar);
  OR2_X1 U482 ( .A1(n497), .A2(n496), .ZN(n603) );
  AND2_X1 U482bar ( .A1(n497bar), .A2(n496bar), .ZN(n603bar);
  OR2_X1 U483 ( .A1(in[112]), .A2(in[102]), .ZN(n496) );
  AND2_X1 U483bar ( .A1(inbar[112]), .A2(inbar[102]), .ZN(n496bar);
  OR2_X1 U484 ( .A1(in[123]), .A2(n495), .ZN(n497) );
  AND2_X1 U484bar ( .A1(inbar[123]), .A2(n495bar), .ZN(n497bar);
  OR2_X1 U485 ( .A1(in[143]), .A2(in[130]), .ZN(n495) );
  AND2_X1 U485bar ( .A1(inbar[143]), .A2(inbar[130]), .ZN(n495bar);
  OR2_X1 U486 ( .A1(n494), .A2(n493), .ZN(n605) );
  AND2_X1 U486bar ( .A1(n494bar), .A2(n493bar), .ZN(n605bar);
  OR2_X1 U487 ( .A1(n492), .A2(n491), .ZN(n493) );
  AND2_X1 U487bar ( .A1(n492bar), .A2(n491bar), .ZN(n493bar);
  OR2_X1 U488 ( .A1(in[216]), .A2(in[213]), .ZN(n491) );
  AND2_X1 U488bar ( .A1(inbar[216]), .A2(inbar[213]), .ZN(n491bar);
  OR2_X1 U489 ( .A1(in[227]), .A2(n490), .ZN(n492) );
  AND2_X1 U489bar ( .A1(inbar[227]), .A2(n490bar), .ZN(n492bar);
  OR2_X1 U490 ( .A1(in_0), .A2(in[248]), .ZN(n490) );
  AND2_X1 U490bar ( .A1(in_0bar), .A2(inbar[248]), .ZN(n490bar);
  OR2_X1 U491 ( .A1(n489), .A2(n488), .ZN(n494) );
  AND2_X1 U491bar ( .A1(n489bar), .A2(n488bar), .ZN(n494bar);
  OR2_X1 U492 ( .A1(in_46), .A2(in_44), .ZN(n488) );
  AND2_X1 U492bar ( .A1(in_46bar), .A2(in_44bar), .ZN(n488bar);
  OR2_X1 U493 ( .A1(in_50), .A2(n487), .ZN(n489) );
  AND2_X1 U493bar ( .A1(in_50bar), .A2(n487bar), .ZN(n489bar);
  OR2_X1 U494 ( .A1(in_9), .A2(in_80), .ZN(n487) );
  AND2_X1 U494bar ( .A1(in_9bar), .A2(in_80bar), .ZN(n487bar);
endmodule




module sBox_4 ( in, out );
  input [7:0] in;
  //input_done

  output [7:0] out;
  //output_done

  wire   [255:0] decodeOut;
  //wire_done

  decode_4 dec ( .in(in), .out(decodeOut) );
  encode_4 enc ( .in(decodeOut), .out(out) );
endmodule


module byteXor_1 ( a, b, y );
  input [7:0] a;
  input [7:0] b;
  //input_done

  output [7:0] y;
  //output_done
  
  wire   n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64;
  //wire_done

  INV_X1 U1 ( .A(n47), .ZN(n64) );
  INV_X1 U2 ( .A(a[7]), .ZN(n63) );
  INV_X1 U3 ( .A(n45), .ZN(n62) );
  INV_X1 U4 ( .A(a[6]), .ZN(n61) );
  INV_X1 U5 ( .A(n43), .ZN(n60) );
  INV_X1 U6 ( .A(a[5]), .ZN(n59) );
  INV_X1 U7 ( .A(n41), .ZN(n58) );
  INV_X1 U8 ( .A(a[4]), .ZN(n57) );
  INV_X1 U9 ( .A(n39), .ZN(n56) );
  INV_X1 U10 ( .A(a[3]), .ZN(n55) );
  INV_X1 U11 ( .A(n37), .ZN(n54) );
  INV_X1 U12 ( .A(a[2]), .ZN(n53) );
  INV_X1 U13 ( .A(n35), .ZN(n52) );
  INV_X1 U14 ( .A(a[1]), .ZN(n51) );
  INV_X1 U15 ( .A(n33), .ZN(n50) );
  INV_X1 U16 ( .A(a[0]), .ZN(n49) );
  OR2_X1 U17 ( .A1(n48), .A2(n64), .ZN(y[7]) );
  OR2_X1 U18 ( .A1(n63), .A2(b[7]), .ZN(n47) );
  AND2_X1 U19 ( .A1(b[7]), .A2(n63), .ZN(n48) );
  OR2_X1 U20 ( .A1(n46), .A2(n62), .ZN(y[6]) );
  OR2_X1 U21 ( .A1(n61), .A2(b[6]), .ZN(n45) );
  AND2_X1 U22 ( .A1(b[6]), .A2(n61), .ZN(n46) );
  OR2_X1 U23 ( .A1(n44), .A2(n60), .ZN(y[5]) );
  OR2_X1 U24 ( .A1(n59), .A2(b[5]), .ZN(n43) );
  AND2_X1 U25 ( .A1(b[5]), .A2(n59), .ZN(n44) );
  OR2_X1 U26 ( .A1(n42), .A2(n58), .ZN(y[4]) );
  OR2_X1 U27 ( .A1(n57), .A2(b[4]), .ZN(n41) );
  AND2_X1 U28 ( .A1(b[4]), .A2(n57), .ZN(n42) );
  OR2_X1 U29 ( .A1(n40), .A2(n56), .ZN(y[3]) );
  OR2_X1 U30 ( .A1(n55), .A2(b[3]), .ZN(n39) );
  AND2_X1 U31 ( .A1(b[3]), .A2(n55), .ZN(n40) );
  OR2_X1 U32 ( .A1(n38), .A2(n54), .ZN(y[2]) );
  OR2_X1 U33 ( .A1(n53), .A2(b[2]), .ZN(n37) );
  AND2_X1 U34 ( .A1(b[2]), .A2(n53), .ZN(n38) );
  OR2_X1 U35 ( .A1(n36), .A2(n52), .ZN(y[1]) );
  OR2_X1 U36 ( .A1(n51), .A2(b[1]), .ZN(n35) );
  AND2_X1 U37 ( .A1(b[1]), .A2(n51), .ZN(n36) );
  OR2_X1 U38 ( .A1(n34), .A2(n50), .ZN(y[0]) );
  OR2_X1 U39 ( .A1(n49), .A2(b[0]), .ZN(n33) );
  AND2_X1 U40 ( .A1(b[0]), .A2(n49), .ZN(n34) );
endmodule


module gFunction ( in, rc, out );
  input [31:0] in;
  input [7:0] rc;
  //input_done

  output [31:0] out;
  //output_done

  wire   [7:0] temp;
  //wire_done

  sBox_4 s0 ( .in(in[23:16]), .out(temp) );
  sBox_3 s1 ( .in(in[15:8]), .out(out[23:16]) );
  sBox_2 s2 ( .in(in[7:0]), .out(out[15:8]) );
  sBox_1 s3 ( .in(in[31:24]), .out(out[7:0]) );
  byteXor_1 bx0 ( .a(temp), .b(rc), .y(out[31:24]) );
endmodule


module wordXor_0 ( a, b, y );
  input [31:0] a;
  input [31:0] b;
  //input_done

  output [31:0] y;
  //output_done

  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128;
  //wire_done

  INV_X1 U1 ( .A(n80), .ZN(n1) );
  INV_X1 U2 ( .A(a[31]), .ZN(n2) );
  INV_X1 U3 ( .A(n82), .ZN(n3) );
  INV_X1 U4 ( .A(a[30]), .ZN(n4) );
  INV_X1 U5 ( .A(n86), .ZN(n5) );
  INV_X1 U6 ( .A(a[29]), .ZN(n6) );
  INV_X1 U7 ( .A(n88), .ZN(n7) );
  INV_X1 U8 ( .A(a[28]), .ZN(n8) );
  INV_X1 U9 ( .A(n90), .ZN(n9) );
  INV_X1 U10 ( .A(a[27]), .ZN(n10) );
  INV_X1 U11 ( .A(n92), .ZN(n11) );
  INV_X1 U12 ( .A(a[26]), .ZN(n12) );
  INV_X1 U13 ( .A(n94), .ZN(n13) );
  INV_X1 U14 ( .A(a[25]), .ZN(n14) );
  INV_X1 U15 ( .A(n96), .ZN(n15) );
  INV_X1 U16 ( .A(a[24]), .ZN(n16) );
  INV_X1 U17 ( .A(n98), .ZN(n17) );
  INV_X1 U18 ( .A(a[23]), .ZN(n18) );
  INV_X1 U19 ( .A(n100), .ZN(n19) );
  INV_X1 U20 ( .A(a[22]), .ZN(n20) );
  INV_X1 U21 ( .A(n102), .ZN(n21) );
  INV_X1 U22 ( .A(a[21]), .ZN(n22) );
  INV_X1 U23 ( .A(n104), .ZN(n23) );
  INV_X1 U24 ( .A(a[20]), .ZN(n24) );
  INV_X1 U25 ( .A(n108), .ZN(n25) );
  INV_X1 U26 ( .A(a[19]), .ZN(n26) );
  INV_X1 U27 ( .A(n110), .ZN(n27) );
  INV_X1 U28 ( .A(a[18]), .ZN(n28) );
  INV_X1 U29 ( .A(n112), .ZN(n29) );
  INV_X1 U30 ( .A(a[17]), .ZN(n30) );
  INV_X1 U31 ( .A(n114), .ZN(n31) );
  INV_X1 U32 ( .A(a[16]), .ZN(n32) );
  INV_X1 U33 ( .A(n116), .ZN(n33) );
  INV_X1 U34 ( .A(a[15]), .ZN(n34) );
  INV_X1 U35 ( .A(n118), .ZN(n35) );
  INV_X1 U36 ( .A(a[14]), .ZN(n36) );
  INV_X1 U37 ( .A(n120), .ZN(n37) );
  INV_X1 U38 ( .A(a[13]), .ZN(n38) );
  INV_X1 U39 ( .A(n122), .ZN(n39) );
  INV_X1 U40 ( .A(a[12]), .ZN(n40) );
  INV_X1 U41 ( .A(n124), .ZN(n41) );
  INV_X1 U42 ( .A(a[11]), .ZN(n42) );
  INV_X1 U43 ( .A(n126), .ZN(n43) );
  INV_X1 U44 ( .A(a[10]), .ZN(n44) );
  INV_X1 U45 ( .A(n66), .ZN(n45) );
  INV_X1 U46 ( .A(a[9]), .ZN(n46) );
  INV_X1 U47 ( .A(n68), .ZN(n47) );
  INV_X1 U48 ( .A(a[8]), .ZN(n48) );
  INV_X1 U49 ( .A(n70), .ZN(n49) );
  INV_X1 U50 ( .A(a[7]), .ZN(n50) );
  INV_X1 U51 ( .A(n72), .ZN(n51) );
  INV_X1 U52 ( .A(a[6]), .ZN(n52) );
  INV_X1 U53 ( .A(n74), .ZN(n53) );
  INV_X1 U54 ( .A(a[5]), .ZN(n54) );
  INV_X1 U55 ( .A(n76), .ZN(n55) );
  INV_X1 U56 ( .A(a[4]), .ZN(n56) );
  INV_X1 U57 ( .A(n78), .ZN(n57) );
  INV_X1 U58 ( .A(a[3]), .ZN(n58) );
  INV_X1 U59 ( .A(n84), .ZN(n59) );
  INV_X1 U60 ( .A(a[2]), .ZN(n60) );
  INV_X1 U61 ( .A(n106), .ZN(n61) );
  INV_X1 U62 ( .A(a[1]), .ZN(n62) );
  INV_X1 U63 ( .A(n128), .ZN(n63) );
  INV_X1 U64 ( .A(a[0]), .ZN(n64) );
  OR2_X1 U65 ( .A1(n65), .A2(n45), .ZN(y[9]) );
  OR2_X1 U66 ( .A1(n46), .A2(b[9]), .ZN(n66) );
  AND2_X1 U67 ( .A1(b[9]), .A2(n46), .ZN(n65) );
  OR2_X1 U68 ( .A1(n67), .A2(n47), .ZN(y[8]) );
  OR2_X1 U69 ( .A1(n48), .A2(b[8]), .ZN(n68) );
  AND2_X1 U70 ( .A1(b[8]), .A2(n48), .ZN(n67) );
  OR2_X1 U71 ( .A1(n69), .A2(n49), .ZN(y[7]) );
  OR2_X1 U72 ( .A1(n50), .A2(b[7]), .ZN(n70) );
  AND2_X1 U73 ( .A1(b[7]), .A2(n50), .ZN(n69) );
  OR2_X1 U74 ( .A1(n71), .A2(n51), .ZN(y[6]) );
  OR2_X1 U75 ( .A1(n52), .A2(b[6]), .ZN(n72) );
  AND2_X1 U76 ( .A1(b[6]), .A2(n52), .ZN(n71) );
  OR2_X1 U77 ( .A1(n73), .A2(n53), .ZN(y[5]) );
  OR2_X1 U78 ( .A1(n54), .A2(b[5]), .ZN(n74) );
  AND2_X1 U79 ( .A1(b[5]), .A2(n54), .ZN(n73) );
  OR2_X1 U80 ( .A1(n75), .A2(n55), .ZN(y[4]) );
  OR2_X1 U81 ( .A1(n56), .A2(b[4]), .ZN(n76) );
  AND2_X1 U82 ( .A1(b[4]), .A2(n56), .ZN(n75) );
  OR2_X1 U83 ( .A1(n77), .A2(n57), .ZN(y[3]) );
  OR2_X1 U84 ( .A1(n58), .A2(b[3]), .ZN(n78) );
  AND2_X1 U85 ( .A1(b[3]), .A2(n58), .ZN(n77) );
  OR2_X1 U86 ( .A1(n79), .A2(n1), .ZN(y[31]) );
  OR2_X1 U87 ( .A1(n2), .A2(b[31]), .ZN(n80) );
  AND2_X1 U88 ( .A1(b[31]), .A2(n2), .ZN(n79) );
  OR2_X1 U89 ( .A1(n81), .A2(n3), .ZN(y[30]) );
  OR2_X1 U90 ( .A1(n4), .A2(b[30]), .ZN(n82) );
  AND2_X1 U91 ( .A1(b[30]), .A2(n4), .ZN(n81) );
  OR2_X1 U92 ( .A1(n83), .A2(n59), .ZN(y[2]) );
  OR2_X1 U93 ( .A1(n60), .A2(b[2]), .ZN(n84) );
  AND2_X1 U94 ( .A1(b[2]), .A2(n60), .ZN(n83) );
  OR2_X1 U95 ( .A1(n85), .A2(n5), .ZN(y[29]) );
  OR2_X1 U96 ( .A1(n6), .A2(b[29]), .ZN(n86) );
  AND2_X1 U97 ( .A1(b[29]), .A2(n6), .ZN(n85) );
  OR2_X1 U98 ( .A1(n87), .A2(n7), .ZN(y[28]) );
  OR2_X1 U99 ( .A1(n8), .A2(b[28]), .ZN(n88) );
  AND2_X1 U100 ( .A1(b[28]), .A2(n8), .ZN(n87) );
  OR2_X1 U101 ( .A1(n89), .A2(n9), .ZN(y[27]) );
  OR2_X1 U102 ( .A1(n10), .A2(b[27]), .ZN(n90) );
  AND2_X1 U103 ( .A1(b[27]), .A2(n10), .ZN(n89) );
  OR2_X1 U104 ( .A1(n91), .A2(n11), .ZN(y[26]) );
  OR2_X1 U105 ( .A1(n12), .A2(b[26]), .ZN(n92) );
  AND2_X1 U106 ( .A1(b[26]), .A2(n12), .ZN(n91) );
  OR2_X1 U107 ( .A1(n93), .A2(n13), .ZN(y[25]) );
  OR2_X1 U108 ( .A1(n14), .A2(b[25]), .ZN(n94) );
  AND2_X1 U109 ( .A1(b[25]), .A2(n14), .ZN(n93) );
  OR2_X1 U110 ( .A1(n95), .A2(n15), .ZN(y[24]) );
  OR2_X1 U111 ( .A1(n16), .A2(b[24]), .ZN(n96) );
  AND2_X1 U112 ( .A1(b[24]), .A2(n16), .ZN(n95) );
  OR2_X1 U113 ( .A1(n97), .A2(n17), .ZN(y[23]) );
  OR2_X1 U114 ( .A1(n18), .A2(b[23]), .ZN(n98) );
  AND2_X1 U115 ( .A1(b[23]), .A2(n18), .ZN(n97) );
  OR2_X1 U116 ( .A1(n99), .A2(n19), .ZN(y[22]) );
  OR2_X1 U117 ( .A1(n20), .A2(b[22]), .ZN(n100) );
  AND2_X1 U118 ( .A1(b[22]), .A2(n20), .ZN(n99) );
  OR2_X1 U119 ( .A1(n101), .A2(n21), .ZN(y[21]) );
  OR2_X1 U120 ( .A1(n22), .A2(b[21]), .ZN(n102) );
  AND2_X1 U121 ( .A1(b[21]), .A2(n22), .ZN(n101) );
  OR2_X1 U122 ( .A1(n103), .A2(n23), .ZN(y[20]) );
  OR2_X1 U123 ( .A1(n24), .A2(b[20]), .ZN(n104) );
  AND2_X1 U124 ( .A1(b[20]), .A2(n24), .ZN(n103) );
  OR2_X1 U125 ( .A1(n105), .A2(n61), .ZN(y[1]) );
  OR2_X1 U126 ( .A1(n62), .A2(b[1]), .ZN(n106) );
  AND2_X1 U127 ( .A1(b[1]), .A2(n62), .ZN(n105) );
  OR2_X1 U128 ( .A1(n107), .A2(n25), .ZN(y[19]) );
  OR2_X1 U129 ( .A1(n26), .A2(b[19]), .ZN(n108) );
  AND2_X1 U130 ( .A1(b[19]), .A2(n26), .ZN(n107) );
  OR2_X1 U131 ( .A1(n109), .A2(n27), .ZN(y[18]) );
  OR2_X1 U132 ( .A1(n28), .A2(b[18]), .ZN(n110) );
  AND2_X1 U133 ( .A1(b[18]), .A2(n28), .ZN(n109) );
  OR2_X1 U134 ( .A1(n111), .A2(n29), .ZN(y[17]) );
  OR2_X1 U135 ( .A1(n30), .A2(b[17]), .ZN(n112) );
  AND2_X1 U136 ( .A1(b[17]), .A2(n30), .ZN(n111) );
  OR2_X1 U137 ( .A1(n113), .A2(n31), .ZN(y[16]) );
  OR2_X1 U138 ( .A1(n32), .A2(b[16]), .ZN(n114) );
  AND2_X1 U139 ( .A1(b[16]), .A2(n32), .ZN(n113) );
  OR2_X1 U140 ( .A1(n115), .A2(n33), .ZN(y[15]) );
  OR2_X1 U141 ( .A1(n34), .A2(b[15]), .ZN(n116) );
  AND2_X1 U142 ( .A1(b[15]), .A2(n34), .ZN(n115) );
  OR2_X1 U143 ( .A1(n117), .A2(n35), .ZN(y[14]) );
  OR2_X1 U144 ( .A1(n36), .A2(b[14]), .ZN(n118) );
  AND2_X1 U145 ( .A1(b[14]), .A2(n36), .ZN(n117) );
  OR2_X1 U146 ( .A1(n119), .A2(n37), .ZN(y[13]) );
  OR2_X1 U147 ( .A1(n38), .A2(b[13]), .ZN(n120) );
  AND2_X1 U148 ( .A1(b[13]), .A2(n38), .ZN(n119) );
  OR2_X1 U149 ( .A1(n121), .A2(n39), .ZN(y[12]) );
  OR2_X1 U150 ( .A1(n40), .A2(b[12]), .ZN(n122) );
  AND2_X1 U151 ( .A1(b[12]), .A2(n40), .ZN(n121) );
  OR2_X1 U152 ( .A1(n123), .A2(n41), .ZN(y[11]) );
  OR2_X1 U153 ( .A1(n42), .A2(b[11]), .ZN(n124) );
  AND2_X1 U154 ( .A1(b[11]), .A2(n42), .ZN(n123) );
  OR2_X1 U155 ( .A1(n125), .A2(n43), .ZN(y[10]) );
  OR2_X1 U156 ( .A1(n44), .A2(b[10]), .ZN(n126) );
  AND2_X1 U157 ( .A1(b[10]), .A2(n44), .ZN(n125) );
  OR2_X1 U158 ( .A1(n127), .A2(n63), .ZN(y[0]) );
  OR2_X1 U159 ( .A1(n64), .A2(b[0]), .ZN(n128) );
  AND2_X1 U160 ( .A1(b[0]), .A2(n64), .ZN(n127) );
endmodule


module mux128_1 ( a, b, sel, y );
  input [127:0] a;
  input [127:0] b;
  input sel;
  //input_done

  output [127:0] y;
  //output_done
  
  wire   n1, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516;
  //wire_done

  OR2_X1 U2 ( .A1(n516), .A2(n515), .ZN(y[9]) );
  AND2_X1 U3 ( .A1(sel), .A2(b[9]), .ZN(n515) );
  AND2_X1 U4 ( .A1(a[9]), .A2(n258), .ZN(n516) );
  OR2_X1 U5 ( .A1(n514), .A2(n513), .ZN(y[99]) );
  AND2_X1 U6 ( .A1(b[99]), .A2(sel), .ZN(n513) );
  AND2_X1 U7 ( .A1(a[99]), .A2(n258), .ZN(n514) );
  OR2_X1 U8 ( .A1(n512), .A2(n511), .ZN(y[98]) );
  AND2_X1 U9 ( .A1(b[98]), .A2(sel), .ZN(n511) );
  AND2_X1 U10 ( .A1(a[98]), .A2(n258), .ZN(n512) );
  OR2_X1 U11 ( .A1(n510), .A2(n509), .ZN(y[97]) );
  AND2_X1 U12 ( .A1(b[97]), .A2(sel), .ZN(n509) );
  AND2_X1 U13 ( .A1(a[97]), .A2(n258), .ZN(n510) );
  OR2_X1 U14 ( .A1(n508), .A2(n507), .ZN(y[96]) );
  AND2_X1 U15 ( .A1(b[96]), .A2(sel), .ZN(n507) );
  AND2_X1 U16 ( .A1(a[96]), .A2(n258), .ZN(n508) );
  OR2_X1 U17 ( .A1(n506), .A2(n505), .ZN(y[95]) );
  AND2_X1 U18 ( .A1(b[95]), .A2(sel), .ZN(n505) );
  AND2_X1 U19 ( .A1(a[95]), .A2(n258), .ZN(n506) );
  OR2_X1 U20 ( .A1(n504), .A2(n503), .ZN(y[94]) );
  AND2_X1 U21 ( .A1(b[94]), .A2(sel), .ZN(n503) );
  AND2_X1 U22 ( .A1(a[94]), .A2(n258), .ZN(n504) );
  OR2_X1 U23 ( .A1(n502), .A2(n501), .ZN(y[93]) );
  AND2_X1 U24 ( .A1(b[93]), .A2(sel), .ZN(n501) );
  AND2_X1 U25 ( .A1(a[93]), .A2(n258), .ZN(n502) );
  OR2_X1 U26 ( .A1(n500), .A2(n499), .ZN(y[92]) );
  AND2_X1 U27 ( .A1(b[92]), .A2(sel), .ZN(n499) );
  AND2_X1 U28 ( .A1(a[92]), .A2(n258), .ZN(n500) );
  OR2_X1 U29 ( .A1(n498), .A2(n497), .ZN(y[91]) );
  AND2_X1 U30 ( .A1(b[91]), .A2(sel), .ZN(n497) );
  AND2_X1 U31 ( .A1(a[91]), .A2(n258), .ZN(n498) );
  OR2_X1 U32 ( .A1(n496), .A2(n495), .ZN(y[90]) );
  AND2_X1 U33 ( .A1(b[90]), .A2(sel), .ZN(n495) );
  AND2_X1 U34 ( .A1(a[90]), .A2(n258), .ZN(n496) );
  OR2_X1 U35 ( .A1(n494), .A2(n493), .ZN(y[8]) );
  AND2_X1 U36 ( .A1(b[8]), .A2(sel), .ZN(n493) );
  AND2_X1 U37 ( .A1(a[8]), .A2(n260), .ZN(n494) );
  OR2_X1 U38 ( .A1(n492), .A2(n491), .ZN(y[89]) );
  AND2_X1 U39 ( .A1(b[89]), .A2(sel), .ZN(n491) );
  AND2_X1 U40 ( .A1(a[89]), .A2(n258), .ZN(n492) );
  OR2_X1 U41 ( .A1(n490), .A2(n489), .ZN(y[88]) );
  AND2_X1 U42 ( .A1(b[88]), .A2(sel), .ZN(n489) );
  AND2_X1 U43 ( .A1(a[88]), .A2(n1), .ZN(n490) );
  OR2_X1 U44 ( .A1(n488), .A2(n487), .ZN(y[87]) );
  AND2_X1 U45 ( .A1(b[87]), .A2(sel), .ZN(n487) );
  AND2_X1 U46 ( .A1(a[87]), .A2(n259), .ZN(n488) );
  OR2_X1 U47 ( .A1(n486), .A2(n485), .ZN(y[86]) );
  AND2_X1 U48 ( .A1(b[86]), .A2(sel), .ZN(n485) );
  AND2_X1 U49 ( .A1(a[86]), .A2(n260), .ZN(n486) );
  OR2_X1 U50 ( .A1(n484), .A2(n483), .ZN(y[85]) );
  AND2_X1 U51 ( .A1(b[85]), .A2(sel), .ZN(n483) );
  AND2_X1 U52 ( .A1(a[85]), .A2(n260), .ZN(n484) );
  OR2_X1 U53 ( .A1(n482), .A2(n481), .ZN(y[84]) );
  AND2_X1 U54 ( .A1(b[84]), .A2(sel), .ZN(n481) );
  AND2_X1 U55 ( .A1(a[84]), .A2(n258), .ZN(n482) );
  OR2_X1 U56 ( .A1(n480), .A2(n479), .ZN(y[83]) );
  AND2_X1 U57 ( .A1(b[83]), .A2(sel), .ZN(n479) );
  AND2_X1 U58 ( .A1(a[83]), .A2(n1), .ZN(n480) );
  OR2_X1 U59 ( .A1(n478), .A2(n477), .ZN(y[82]) );
  AND2_X1 U60 ( .A1(b[82]), .A2(sel), .ZN(n477) );
  AND2_X1 U61 ( .A1(a[82]), .A2(n259), .ZN(n478) );
  OR2_X1 U62 ( .A1(n476), .A2(n475), .ZN(y[81]) );
  AND2_X1 U63 ( .A1(b[81]), .A2(sel), .ZN(n475) );
  AND2_X1 U64 ( .A1(a[81]), .A2(n260), .ZN(n476) );
  OR2_X1 U65 ( .A1(n474), .A2(n473), .ZN(y[80]) );
  AND2_X1 U66 ( .A1(b[80]), .A2(sel), .ZN(n473) );
  AND2_X1 U67 ( .A1(a[80]), .A2(n1), .ZN(n474) );
  OR2_X1 U68 ( .A1(n472), .A2(n471), .ZN(y[7]) );
  AND2_X1 U69 ( .A1(b[7]), .A2(sel), .ZN(n471) );
  AND2_X1 U70 ( .A1(a[7]), .A2(n258), .ZN(n472) );
  OR2_X1 U71 ( .A1(n470), .A2(n469), .ZN(y[79]) );
  AND2_X1 U72 ( .A1(b[79]), .A2(sel), .ZN(n469) );
  AND2_X1 U73 ( .A1(a[79]), .A2(n258), .ZN(n470) );
  OR2_X1 U74 ( .A1(n468), .A2(n467), .ZN(y[78]) );
  AND2_X1 U75 ( .A1(b[78]), .A2(sel), .ZN(n467) );
  AND2_X1 U76 ( .A1(a[78]), .A2(n259), .ZN(n468) );
  OR2_X1 U77 ( .A1(n466), .A2(n465), .ZN(y[77]) );
  AND2_X1 U78 ( .A1(b[77]), .A2(sel), .ZN(n465) );
  AND2_X1 U79 ( .A1(a[77]), .A2(n1), .ZN(n466) );
  OR2_X1 U80 ( .A1(n464), .A2(n463), .ZN(y[76]) );
  AND2_X1 U81 ( .A1(b[76]), .A2(sel), .ZN(n463) );
  AND2_X1 U82 ( .A1(a[76]), .A2(n260), .ZN(n464) );
  OR2_X1 U83 ( .A1(n462), .A2(n461), .ZN(y[75]) );
  AND2_X1 U84 ( .A1(b[75]), .A2(sel), .ZN(n461) );
  AND2_X1 U85 ( .A1(a[75]), .A2(n260), .ZN(n462) );
  OR2_X1 U86 ( .A1(n460), .A2(n459), .ZN(y[74]) );
  AND2_X1 U87 ( .A1(b[74]), .A2(sel), .ZN(n459) );
  AND2_X1 U88 ( .A1(a[74]), .A2(n1), .ZN(n460) );
  OR2_X1 U89 ( .A1(n458), .A2(n457), .ZN(y[73]) );
  AND2_X1 U90 ( .A1(b[73]), .A2(sel), .ZN(n457) );
  AND2_X1 U91 ( .A1(a[73]), .A2(n258), .ZN(n458) );
  OR2_X1 U92 ( .A1(n456), .A2(n455), .ZN(y[72]) );
  AND2_X1 U93 ( .A1(b[72]), .A2(sel), .ZN(n455) );
  AND2_X1 U94 ( .A1(a[72]), .A2(n259), .ZN(n456) );
  OR2_X1 U95 ( .A1(n454), .A2(n453), .ZN(y[71]) );
  AND2_X1 U96 ( .A1(b[71]), .A2(sel), .ZN(n453) );
  AND2_X1 U97 ( .A1(a[71]), .A2(n1), .ZN(n454) );
  OR2_X1 U98 ( .A1(n452), .A2(n451), .ZN(y[70]) );
  AND2_X1 U99 ( .A1(b[70]), .A2(sel), .ZN(n451) );
  AND2_X1 U100 ( .A1(a[70]), .A2(n1), .ZN(n452) );
  OR2_X1 U101 ( .A1(n450), .A2(n449), .ZN(y[6]) );
  AND2_X1 U102 ( .A1(b[6]), .A2(sel), .ZN(n449) );
  AND2_X1 U103 ( .A1(a[6]), .A2(n260), .ZN(n450) );
  OR2_X1 U104 ( .A1(n448), .A2(n447), .ZN(y[69]) );
  AND2_X1 U105 ( .A1(b[69]), .A2(sel), .ZN(n447) );
  AND2_X1 U106 ( .A1(a[69]), .A2(n260), .ZN(n448) );
  OR2_X1 U107 ( .A1(n446), .A2(n445), .ZN(y[68]) );
  AND2_X1 U108 ( .A1(b[68]), .A2(sel), .ZN(n445) );
  AND2_X1 U109 ( .A1(a[68]), .A2(n1), .ZN(n446) );
  OR2_X1 U110 ( .A1(n444), .A2(n443), .ZN(y[67]) );
  AND2_X1 U111 ( .A1(b[67]), .A2(sel), .ZN(n443) );
  AND2_X1 U112 ( .A1(a[67]), .A2(n260), .ZN(n444) );
  OR2_X1 U113 ( .A1(n442), .A2(n441), .ZN(y[66]) );
  AND2_X1 U114 ( .A1(b[66]), .A2(sel), .ZN(n441) );
  AND2_X1 U115 ( .A1(a[66]), .A2(n258), .ZN(n442) );
  OR2_X1 U116 ( .A1(n440), .A2(n439), .ZN(y[65]) );
  AND2_X1 U117 ( .A1(b[65]), .A2(sel), .ZN(n439) );
  AND2_X1 U118 ( .A1(a[65]), .A2(n1), .ZN(n440) );
  OR2_X1 U119 ( .A1(n438), .A2(n437), .ZN(y[64]) );
  AND2_X1 U120 ( .A1(b[64]), .A2(sel), .ZN(n437) );
  AND2_X1 U121 ( .A1(a[64]), .A2(n260), .ZN(n438) );
  OR2_X1 U122 ( .A1(n436), .A2(n435), .ZN(y[63]) );
  AND2_X1 U123 ( .A1(b[63]), .A2(sel), .ZN(n435) );
  AND2_X1 U124 ( .A1(a[63]), .A2(n259), .ZN(n436) );
  OR2_X1 U125 ( .A1(n434), .A2(n433), .ZN(y[62]) );
  AND2_X1 U126 ( .A1(b[62]), .A2(sel), .ZN(n433) );
  AND2_X1 U127 ( .A1(a[62]), .A2(n258), .ZN(n434) );
  OR2_X1 U128 ( .A1(n432), .A2(n431), .ZN(y[61]) );
  AND2_X1 U129 ( .A1(b[61]), .A2(sel), .ZN(n431) );
  AND2_X1 U130 ( .A1(a[61]), .A2(n260), .ZN(n432) );
  OR2_X1 U131 ( .A1(n430), .A2(n429), .ZN(y[60]) );
  AND2_X1 U132 ( .A1(b[60]), .A2(sel), .ZN(n429) );
  AND2_X1 U133 ( .A1(a[60]), .A2(n259), .ZN(n430) );
  OR2_X1 U134 ( .A1(n428), .A2(n427), .ZN(y[5]) );
  AND2_X1 U135 ( .A1(b[5]), .A2(sel), .ZN(n427) );
  AND2_X1 U136 ( .A1(a[5]), .A2(n1), .ZN(n428) );
  OR2_X1 U137 ( .A1(n426), .A2(n425), .ZN(y[59]) );
  AND2_X1 U138 ( .A1(b[59]), .A2(sel), .ZN(n425) );
  AND2_X1 U139 ( .A1(a[59]), .A2(n259), .ZN(n426) );
  OR2_X1 U140 ( .A1(n424), .A2(n423), .ZN(y[58]) );
  AND2_X1 U141 ( .A1(b[58]), .A2(sel), .ZN(n423) );
  AND2_X1 U142 ( .A1(a[58]), .A2(n258), .ZN(n424) );
  OR2_X1 U143 ( .A1(n422), .A2(n421), .ZN(y[57]) );
  AND2_X1 U144 ( .A1(b[57]), .A2(sel), .ZN(n421) );
  AND2_X1 U145 ( .A1(a[57]), .A2(n1), .ZN(n422) );
  OR2_X1 U146 ( .A1(n420), .A2(n419), .ZN(y[56]) );
  AND2_X1 U147 ( .A1(b[56]), .A2(sel), .ZN(n419) );
  AND2_X1 U148 ( .A1(a[56]), .A2(n259), .ZN(n420) );
  OR2_X1 U149 ( .A1(n418), .A2(n417), .ZN(y[55]) );
  AND2_X1 U150 ( .A1(b[55]), .A2(sel), .ZN(n417) );
  AND2_X1 U151 ( .A1(a[55]), .A2(n1), .ZN(n418) );
  OR2_X1 U152 ( .A1(n416), .A2(n415), .ZN(y[54]) );
  AND2_X1 U153 ( .A1(b[54]), .A2(sel), .ZN(n415) );
  AND2_X1 U154 ( .A1(a[54]), .A2(n259), .ZN(n416) );
  OR2_X1 U155 ( .A1(n414), .A2(n413), .ZN(y[53]) );
  AND2_X1 U156 ( .A1(b[53]), .A2(sel), .ZN(n413) );
  AND2_X1 U157 ( .A1(a[53]), .A2(n259), .ZN(n414) );
  OR2_X1 U158 ( .A1(n412), .A2(n411), .ZN(y[52]) );
  AND2_X1 U159 ( .A1(b[52]), .A2(sel), .ZN(n411) );
  AND2_X1 U160 ( .A1(a[52]), .A2(n260), .ZN(n412) );
  OR2_X1 U161 ( .A1(n410), .A2(n409), .ZN(y[51]) );
  AND2_X1 U162 ( .A1(b[51]), .A2(sel), .ZN(n409) );
  AND2_X1 U163 ( .A1(a[51]), .A2(n259), .ZN(n410) );
  OR2_X1 U164 ( .A1(n408), .A2(n407), .ZN(y[50]) );
  AND2_X1 U165 ( .A1(b[50]), .A2(sel), .ZN(n407) );
  AND2_X1 U166 ( .A1(a[50]), .A2(n1), .ZN(n408) );
  OR2_X1 U167 ( .A1(n406), .A2(n405), .ZN(y[4]) );
  AND2_X1 U168 ( .A1(b[4]), .A2(sel), .ZN(n405) );
  AND2_X1 U169 ( .A1(a[4]), .A2(n260), .ZN(n406) );
  OR2_X1 U170 ( .A1(n404), .A2(n403), .ZN(y[49]) );
  AND2_X1 U171 ( .A1(b[49]), .A2(sel), .ZN(n403) );
  AND2_X1 U172 ( .A1(a[49]), .A2(n1), .ZN(n404) );
  OR2_X1 U173 ( .A1(n402), .A2(n401), .ZN(y[48]) );
  AND2_X1 U174 ( .A1(b[48]), .A2(sel), .ZN(n401) );
  AND2_X1 U175 ( .A1(a[48]), .A2(n258), .ZN(n402) );
  OR2_X1 U176 ( .A1(n400), .A2(n399), .ZN(y[47]) );
  AND2_X1 U177 ( .A1(b[47]), .A2(sel), .ZN(n399) );
  AND2_X1 U178 ( .A1(a[47]), .A2(n260), .ZN(n400) );
  OR2_X1 U179 ( .A1(n398), .A2(n397), .ZN(y[46]) );
  AND2_X1 U180 ( .A1(b[46]), .A2(sel), .ZN(n397) );
  AND2_X1 U181 ( .A1(a[46]), .A2(n260), .ZN(n398) );
  OR2_X1 U182 ( .A1(n396), .A2(n395), .ZN(y[45]) );
  AND2_X1 U183 ( .A1(b[45]), .A2(sel), .ZN(n395) );
  AND2_X1 U184 ( .A1(a[45]), .A2(n258), .ZN(n396) );
  OR2_X1 U185 ( .A1(n394), .A2(n393), .ZN(y[44]) );
  AND2_X1 U186 ( .A1(b[44]), .A2(sel), .ZN(n393) );
  AND2_X1 U187 ( .A1(a[44]), .A2(n259), .ZN(n394) );
  OR2_X1 U188 ( .A1(n392), .A2(n391), .ZN(y[43]) );
  AND2_X1 U189 ( .A1(b[43]), .A2(sel), .ZN(n391) );
  AND2_X1 U190 ( .A1(a[43]), .A2(n258), .ZN(n392) );
  OR2_X1 U191 ( .A1(n390), .A2(n389), .ZN(y[42]) );
  AND2_X1 U192 ( .A1(b[42]), .A2(sel), .ZN(n389) );
  AND2_X1 U193 ( .A1(a[42]), .A2(n1), .ZN(n390) );
  OR2_X1 U194 ( .A1(n388), .A2(n387), .ZN(y[41]) );
  AND2_X1 U195 ( .A1(b[41]), .A2(sel), .ZN(n387) );
  AND2_X1 U196 ( .A1(a[41]), .A2(n260), .ZN(n388) );
  OR2_X1 U197 ( .A1(n386), .A2(n385), .ZN(y[40]) );
  AND2_X1 U198 ( .A1(b[40]), .A2(sel), .ZN(n385) );
  AND2_X1 U199 ( .A1(a[40]), .A2(n260), .ZN(n386) );
  OR2_X1 U200 ( .A1(n384), .A2(n383), .ZN(y[3]) );
  AND2_X1 U201 ( .A1(b[3]), .A2(sel), .ZN(n383) );
  AND2_X1 U202 ( .A1(a[3]), .A2(n258), .ZN(n384) );
  OR2_X1 U203 ( .A1(n382), .A2(n381), .ZN(y[39]) );
  AND2_X1 U204 ( .A1(b[39]), .A2(sel), .ZN(n381) );
  AND2_X1 U205 ( .A1(a[39]), .A2(n259), .ZN(n382) );
  OR2_X1 U206 ( .A1(n380), .A2(n379), .ZN(y[38]) );
  AND2_X1 U207 ( .A1(b[38]), .A2(sel), .ZN(n379) );
  AND2_X1 U208 ( .A1(a[38]), .A2(n259), .ZN(n380) );
  OR2_X1 U209 ( .A1(n378), .A2(n377), .ZN(y[37]) );
  AND2_X1 U210 ( .A1(b[37]), .A2(sel), .ZN(n377) );
  AND2_X1 U211 ( .A1(a[37]), .A2(n1), .ZN(n378) );
  OR2_X1 U212 ( .A1(n376), .A2(n375), .ZN(y[36]) );
  AND2_X1 U213 ( .A1(b[36]), .A2(sel), .ZN(n375) );
  AND2_X1 U214 ( .A1(a[36]), .A2(n260), .ZN(n376) );
  OR2_X1 U215 ( .A1(n374), .A2(n373), .ZN(y[35]) );
  AND2_X1 U216 ( .A1(b[35]), .A2(sel), .ZN(n373) );
  AND2_X1 U217 ( .A1(a[35]), .A2(n260), .ZN(n374) );
  OR2_X1 U218 ( .A1(n372), .A2(n371), .ZN(y[34]) );
  AND2_X1 U219 ( .A1(b[34]), .A2(sel), .ZN(n371) );
  AND2_X1 U220 ( .A1(a[34]), .A2(n260), .ZN(n372) );
  OR2_X1 U221 ( .A1(n370), .A2(n369), .ZN(y[33]) );
  AND2_X1 U222 ( .A1(b[33]), .A2(sel), .ZN(n369) );
  AND2_X1 U223 ( .A1(a[33]), .A2(n260), .ZN(n370) );
  OR2_X1 U224 ( .A1(n368), .A2(n367), .ZN(y[32]) );
  AND2_X1 U225 ( .A1(b[32]), .A2(sel), .ZN(n367) );
  AND2_X1 U226 ( .A1(a[32]), .A2(n258), .ZN(n368) );
  OR2_X1 U227 ( .A1(n366), .A2(n365), .ZN(y[31]) );
  AND2_X1 U228 ( .A1(b[31]), .A2(sel), .ZN(n365) );
  AND2_X1 U229 ( .A1(a[31]), .A2(n259), .ZN(n366) );
  OR2_X1 U230 ( .A1(n364), .A2(n363), .ZN(y[30]) );
  AND2_X1 U231 ( .A1(b[30]), .A2(sel), .ZN(n363) );
  AND2_X1 U232 ( .A1(a[30]), .A2(n1), .ZN(n364) );
  OR2_X1 U233 ( .A1(n362), .A2(n361), .ZN(y[2]) );
  AND2_X1 U234 ( .A1(b[2]), .A2(sel), .ZN(n361) );
  AND2_X1 U235 ( .A1(a[2]), .A2(n258), .ZN(n362) );
  OR2_X1 U236 ( .A1(n360), .A2(n359), .ZN(y[29]) );
  AND2_X1 U237 ( .A1(b[29]), .A2(sel), .ZN(n359) );
  AND2_X1 U238 ( .A1(a[29]), .A2(n259), .ZN(n360) );
  OR2_X1 U239 ( .A1(n358), .A2(n357), .ZN(y[28]) );
  AND2_X1 U240 ( .A1(b[28]), .A2(sel), .ZN(n357) );
  AND2_X1 U241 ( .A1(a[28]), .A2(n1), .ZN(n358) );
  OR2_X1 U242 ( .A1(n356), .A2(n355), .ZN(y[27]) );
  AND2_X1 U243 ( .A1(b[27]), .A2(sel), .ZN(n355) );
  AND2_X1 U244 ( .A1(a[27]), .A2(n260), .ZN(n356) );
  OR2_X1 U245 ( .A1(n354), .A2(n353), .ZN(y[26]) );
  AND2_X1 U246 ( .A1(b[26]), .A2(sel), .ZN(n353) );
  AND2_X1 U247 ( .A1(a[26]), .A2(n259), .ZN(n354) );
  OR2_X1 U248 ( .A1(n352), .A2(n351), .ZN(y[25]) );
  AND2_X1 U249 ( .A1(b[25]), .A2(sel), .ZN(n351) );
  AND2_X1 U250 ( .A1(a[25]), .A2(n259), .ZN(n352) );
  OR2_X1 U251 ( .A1(n350), .A2(n349), .ZN(y[24]) );
  AND2_X1 U252 ( .A1(b[24]), .A2(sel), .ZN(n349) );
  AND2_X1 U253 ( .A1(a[24]), .A2(n260), .ZN(n350) );
  OR2_X1 U254 ( .A1(n348), .A2(n347), .ZN(y[23]) );
  AND2_X1 U255 ( .A1(b[23]), .A2(sel), .ZN(n347) );
  AND2_X1 U256 ( .A1(a[23]), .A2(n1), .ZN(n348) );
  OR2_X1 U257 ( .A1(n346), .A2(n345), .ZN(y[22]) );
  AND2_X1 U258 ( .A1(b[22]), .A2(sel), .ZN(n345) );
  AND2_X1 U259 ( .A1(a[22]), .A2(n258), .ZN(n346) );
  OR2_X1 U260 ( .A1(n344), .A2(n343), .ZN(y[21]) );
  AND2_X1 U261 ( .A1(b[21]), .A2(sel), .ZN(n343) );
  AND2_X1 U262 ( .A1(a[21]), .A2(n259), .ZN(n344) );
  OR2_X1 U263 ( .A1(n342), .A2(n341), .ZN(y[20]) );
  AND2_X1 U264 ( .A1(b[20]), .A2(sel), .ZN(n341) );
  AND2_X1 U265 ( .A1(a[20]), .A2(n1), .ZN(n342) );
  OR2_X1 U266 ( .A1(n340), .A2(n339), .ZN(y[1]) );
  AND2_X1 U267 ( .A1(b[1]), .A2(sel), .ZN(n339) );
  AND2_X1 U268 ( .A1(a[1]), .A2(n1), .ZN(n340) );
  OR2_X1 U269 ( .A1(n338), .A2(n337), .ZN(y[19]) );
  AND2_X1 U270 ( .A1(b[19]), .A2(sel), .ZN(n337) );
  AND2_X1 U271 ( .A1(a[19]), .A2(n260), .ZN(n338) );
  OR2_X1 U272 ( .A1(n336), .A2(n335), .ZN(y[18]) );
  AND2_X1 U273 ( .A1(b[18]), .A2(sel), .ZN(n335) );
  AND2_X1 U274 ( .A1(a[18]), .A2(n258), .ZN(n336) );
  OR2_X1 U275 ( .A1(n334), .A2(n333), .ZN(y[17]) );
  AND2_X1 U276 ( .A1(b[17]), .A2(sel), .ZN(n333) );
  AND2_X1 U277 ( .A1(a[17]), .A2(n258), .ZN(n334) );
  OR2_X1 U278 ( .A1(n332), .A2(n331), .ZN(y[16]) );
  AND2_X1 U279 ( .A1(b[16]), .A2(sel), .ZN(n331) );
  AND2_X1 U280 ( .A1(a[16]), .A2(n259), .ZN(n332) );
  OR2_X1 U281 ( .A1(n330), .A2(n329), .ZN(y[15]) );
  AND2_X1 U282 ( .A1(b[15]), .A2(sel), .ZN(n329) );
  AND2_X1 U283 ( .A1(a[15]), .A2(n259), .ZN(n330) );
  OR2_X1 U284 ( .A1(n328), .A2(n327), .ZN(y[14]) );
  AND2_X1 U285 ( .A1(b[14]), .A2(sel), .ZN(n327) );
  AND2_X1 U286 ( .A1(a[14]), .A2(n1), .ZN(n328) );
  OR2_X1 U287 ( .A1(n326), .A2(n325), .ZN(y[13]) );
  AND2_X1 U288 ( .A1(b[13]), .A2(sel), .ZN(n325) );
  AND2_X1 U289 ( .A1(a[13]), .A2(n259), .ZN(n326) );
  OR2_X1 U290 ( .A1(n324), .A2(n323), .ZN(y[12]) );
  AND2_X1 U291 ( .A1(b[12]), .A2(sel), .ZN(n323) );
  AND2_X1 U292 ( .A1(a[12]), .A2(n260), .ZN(n324) );
  OR2_X1 U293 ( .A1(n322), .A2(n321), .ZN(y[127]) );
  AND2_X1 U294 ( .A1(b[127]), .A2(sel), .ZN(n321) );
  AND2_X1 U295 ( .A1(a[127]), .A2(n1), .ZN(n322) );
  OR2_X1 U296 ( .A1(n320), .A2(n319), .ZN(y[126]) );
  AND2_X1 U297 ( .A1(b[126]), .A2(sel), .ZN(n319) );
  AND2_X1 U298 ( .A1(a[126]), .A2(n259), .ZN(n320) );
  OR2_X1 U299 ( .A1(n318), .A2(n317), .ZN(y[125]) );
  AND2_X1 U300 ( .A1(b[125]), .A2(sel), .ZN(n317) );
  AND2_X1 U301 ( .A1(a[125]), .A2(n1), .ZN(n318) );
  OR2_X1 U302 ( .A1(n316), .A2(n315), .ZN(y[124]) );
  AND2_X1 U303 ( .A1(b[124]), .A2(sel), .ZN(n315) );
  AND2_X1 U304 ( .A1(a[124]), .A2(n1), .ZN(n316) );
  OR2_X1 U305 ( .A1(n314), .A2(n313), .ZN(y[123]) );
  AND2_X1 U306 ( .A1(b[123]), .A2(sel), .ZN(n313) );
  AND2_X1 U307 ( .A1(a[123]), .A2(n259), .ZN(n314) );
  OR2_X1 U308 ( .A1(n312), .A2(n311), .ZN(y[122]) );
  AND2_X1 U309 ( .A1(b[122]), .A2(sel), .ZN(n311) );
  AND2_X1 U310 ( .A1(a[122]), .A2(n1), .ZN(n312) );
  OR2_X1 U311 ( .A1(n310), .A2(n309), .ZN(y[121]) );
  AND2_X1 U312 ( .A1(b[121]), .A2(sel), .ZN(n309) );
  AND2_X1 U313 ( .A1(a[121]), .A2(n259), .ZN(n310) );
  OR2_X1 U314 ( .A1(n308), .A2(n307), .ZN(y[120]) );
  AND2_X1 U315 ( .A1(b[120]), .A2(sel), .ZN(n307) );
  AND2_X1 U316 ( .A1(a[120]), .A2(n259), .ZN(n308) );
  OR2_X1 U317 ( .A1(n306), .A2(n305), .ZN(y[11]) );
  AND2_X1 U318 ( .A1(b[11]), .A2(sel), .ZN(n305) );
  AND2_X1 U319 ( .A1(a[11]), .A2(n260), .ZN(n306) );
  OR2_X1 U320 ( .A1(n304), .A2(n303), .ZN(y[119]) );
  AND2_X1 U321 ( .A1(b[119]), .A2(sel), .ZN(n303) );
  AND2_X1 U322 ( .A1(a[119]), .A2(n260), .ZN(n304) );
  OR2_X1 U323 ( .A1(n302), .A2(n301), .ZN(y[118]) );
  AND2_X1 U324 ( .A1(b[118]), .A2(sel), .ZN(n301) );
  AND2_X1 U325 ( .A1(a[118]), .A2(n1), .ZN(n302) );
  OR2_X1 U326 ( .A1(n300), .A2(n299), .ZN(y[117]) );
  AND2_X1 U327 ( .A1(b[117]), .A2(sel), .ZN(n299) );
  AND2_X1 U328 ( .A1(a[117]), .A2(n259), .ZN(n300) );
  OR2_X1 U329 ( .A1(n298), .A2(n297), .ZN(y[116]) );
  AND2_X1 U330 ( .A1(b[116]), .A2(sel), .ZN(n297) );
  AND2_X1 U331 ( .A1(a[116]), .A2(n1), .ZN(n298) );
  OR2_X1 U332 ( .A1(n296), .A2(n295), .ZN(y[115]) );
  AND2_X1 U333 ( .A1(b[115]), .A2(sel), .ZN(n295) );
  AND2_X1 U334 ( .A1(a[115]), .A2(n260), .ZN(n296) );
  OR2_X1 U335 ( .A1(n294), .A2(n293), .ZN(y[114]) );
  AND2_X1 U336 ( .A1(b[114]), .A2(sel), .ZN(n293) );
  AND2_X1 U337 ( .A1(a[114]), .A2(n258), .ZN(n294) );
  OR2_X1 U338 ( .A1(n292), .A2(n291), .ZN(y[113]) );
  AND2_X1 U339 ( .A1(b[113]), .A2(sel), .ZN(n291) );
  AND2_X1 U340 ( .A1(a[113]), .A2(n258), .ZN(n292) );
  OR2_X1 U341 ( .A1(n290), .A2(n289), .ZN(y[112]) );
  AND2_X1 U342 ( .A1(b[112]), .A2(sel), .ZN(n289) );
  AND2_X1 U343 ( .A1(a[112]), .A2(n260), .ZN(n290) );
  OR2_X1 U344 ( .A1(n288), .A2(n287), .ZN(y[111]) );
  AND2_X1 U345 ( .A1(b[111]), .A2(sel), .ZN(n287) );
  AND2_X1 U346 ( .A1(a[111]), .A2(n259), .ZN(n288) );
  OR2_X1 U347 ( .A1(n286), .A2(n285), .ZN(y[110]) );
  AND2_X1 U348 ( .A1(b[110]), .A2(sel), .ZN(n285) );
  AND2_X1 U349 ( .A1(a[110]), .A2(n259), .ZN(n286) );
  OR2_X1 U350 ( .A1(n284), .A2(n283), .ZN(y[10]) );
  AND2_X1 U351 ( .A1(b[10]), .A2(sel), .ZN(n283) );
  AND2_X1 U352 ( .A1(a[10]), .A2(n1), .ZN(n284) );
  OR2_X1 U353 ( .A1(n282), .A2(n281), .ZN(y[109]) );
  AND2_X1 U354 ( .A1(b[109]), .A2(sel), .ZN(n281) );
  AND2_X1 U355 ( .A1(a[109]), .A2(n259), .ZN(n282) );
  OR2_X1 U356 ( .A1(n280), .A2(n279), .ZN(y[108]) );
  AND2_X1 U357 ( .A1(b[108]), .A2(sel), .ZN(n279) );
  AND2_X1 U358 ( .A1(a[108]), .A2(n1), .ZN(n280) );
  OR2_X1 U359 ( .A1(n278), .A2(n277), .ZN(y[107]) );
  AND2_X1 U360 ( .A1(b[107]), .A2(sel), .ZN(n277) );
  AND2_X1 U361 ( .A1(a[107]), .A2(n260), .ZN(n278) );
  OR2_X1 U362 ( .A1(n276), .A2(n275), .ZN(y[106]) );
  AND2_X1 U363 ( .A1(b[106]), .A2(sel), .ZN(n275) );
  AND2_X1 U364 ( .A1(a[106]), .A2(n1), .ZN(n276) );
  OR2_X1 U365 ( .A1(n274), .A2(n273), .ZN(y[105]) );
  AND2_X1 U366 ( .A1(b[105]), .A2(sel), .ZN(n273) );
  AND2_X1 U367 ( .A1(a[105]), .A2(n260), .ZN(n274) );
  OR2_X1 U368 ( .A1(n272), .A2(n271), .ZN(y[104]) );
  AND2_X1 U369 ( .A1(b[104]), .A2(sel), .ZN(n271) );
  AND2_X1 U370 ( .A1(a[104]), .A2(n258), .ZN(n272) );
  OR2_X1 U371 ( .A1(n270), .A2(n269), .ZN(y[103]) );
  AND2_X1 U372 ( .A1(b[103]), .A2(sel), .ZN(n269) );
  AND2_X1 U373 ( .A1(a[103]), .A2(n258), .ZN(n270) );
  OR2_X1 U374 ( .A1(n268), .A2(n267), .ZN(y[102]) );
  AND2_X1 U375 ( .A1(b[102]), .A2(sel), .ZN(n267) );
  AND2_X1 U376 ( .A1(a[102]), .A2(n259), .ZN(n268) );
  OR2_X1 U377 ( .A1(n266), .A2(n265), .ZN(y[101]) );
  AND2_X1 U378 ( .A1(b[101]), .A2(sel), .ZN(n265) );
  AND2_X1 U379 ( .A1(a[101]), .A2(n260), .ZN(n266) );
  OR2_X1 U380 ( .A1(n264), .A2(n263), .ZN(y[100]) );
  AND2_X1 U381 ( .A1(b[100]), .A2(sel), .ZN(n263) );
  AND2_X1 U382 ( .A1(a[100]), .A2(n259), .ZN(n264) );
  OR2_X1 U383 ( .A1(n262), .A2(n261), .ZN(y[0]) );
  AND2_X1 U384 ( .A1(b[0]), .A2(sel), .ZN(n261) );
  AND2_X1 U385 ( .A1(a[0]), .A2(n1), .ZN(n262) );
  INV_X1 U1 ( .A(sel), .ZN(n1) );
  INV_X1 U386 ( .A(sel), .ZN(n258) );
  INV_X1 U387 ( .A(sel), .ZN(n259) );
  INV_X1 U388 ( .A(sel), .ZN(n260) );
endmodule


module wordXor_1 ( a, b, y );
  input [31:0] a;
  input [31:0] b;
  //input_done

  output [31:0] y;
  //output_done

  wire   n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256;
  //wire_done

  INV_X1 U1 ( .A(n177), .ZN(n256) );
  INV_X1 U2 ( .A(a[31]), .ZN(n255) );
  INV_X1 U3 ( .A(n175), .ZN(n254) );
  INV_X1 U4 ( .A(a[30]), .ZN(n253) );
  INV_X1 U5 ( .A(n171), .ZN(n252) );
  INV_X1 U6 ( .A(a[29]), .ZN(n251) );
  INV_X1 U7 ( .A(n169), .ZN(n250) );
  INV_X1 U8 ( .A(a[28]), .ZN(n249) );
  INV_X1 U9 ( .A(n167), .ZN(n248) );
  INV_X1 U10 ( .A(a[27]), .ZN(n247) );
  INV_X1 U11 ( .A(n165), .ZN(n246) );
  INV_X1 U12 ( .A(a[26]), .ZN(n245) );
  INV_X1 U13 ( .A(n163), .ZN(n244) );
  INV_X1 U14 ( .A(a[25]), .ZN(n243) );
  INV_X1 U15 ( .A(n161), .ZN(n242) );
  INV_X1 U16 ( .A(a[24]), .ZN(n241) );
  INV_X1 U17 ( .A(n159), .ZN(n240) );
  INV_X1 U18 ( .A(a[23]), .ZN(n239) );
  INV_X1 U19 ( .A(n157), .ZN(n238) );
  INV_X1 U20 ( .A(a[22]), .ZN(n237) );
  INV_X1 U21 ( .A(n155), .ZN(n236) );
  INV_X1 U22 ( .A(a[21]), .ZN(n235) );
  INV_X1 U23 ( .A(n153), .ZN(n234) );
  INV_X1 U24 ( .A(a[20]), .ZN(n233) );
  INV_X1 U25 ( .A(n149), .ZN(n232) );
  INV_X1 U26 ( .A(a[19]), .ZN(n231) );
  INV_X1 U27 ( .A(n147), .ZN(n230) );
  INV_X1 U28 ( .A(a[18]), .ZN(n229) );
  INV_X1 U29 ( .A(n145), .ZN(n228) );
  INV_X1 U30 ( .A(a[17]), .ZN(n227) );
  INV_X1 U31 ( .A(n143), .ZN(n226) );
  INV_X1 U32 ( .A(a[16]), .ZN(n225) );
  INV_X1 U33 ( .A(n141), .ZN(n224) );
  INV_X1 U34 ( .A(a[15]), .ZN(n223) );
  INV_X1 U35 ( .A(n139), .ZN(n222) );
  INV_X1 U36 ( .A(a[14]), .ZN(n221) );
  INV_X1 U37 ( .A(n137), .ZN(n220) );
  INV_X1 U38 ( .A(a[13]), .ZN(n219) );
  INV_X1 U39 ( .A(n135), .ZN(n218) );
  INV_X1 U40 ( .A(a[12]), .ZN(n217) );
  INV_X1 U41 ( .A(n133), .ZN(n216) );
  INV_X1 U42 ( .A(a[11]), .ZN(n215) );
  INV_X1 U43 ( .A(n131), .ZN(n214) );
  INV_X1 U44 ( .A(a[10]), .ZN(n213) );
  INV_X1 U45 ( .A(n191), .ZN(n212) );
  INV_X1 U46 ( .A(a[9]), .ZN(n211) );
  INV_X1 U47 ( .A(n189), .ZN(n210) );
  INV_X1 U48 ( .A(a[8]), .ZN(n209) );
  INV_X1 U49 ( .A(n187), .ZN(n208) );
  INV_X1 U50 ( .A(a[7]), .ZN(n207) );
  INV_X1 U51 ( .A(n185), .ZN(n206) );
  INV_X1 U52 ( .A(a[6]), .ZN(n205) );
  INV_X1 U53 ( .A(n183), .ZN(n204) );
  INV_X1 U54 ( .A(a[5]), .ZN(n203) );
  INV_X1 U55 ( .A(n181), .ZN(n202) );
  INV_X1 U56 ( .A(a[4]), .ZN(n201) );
  INV_X1 U57 ( .A(n179), .ZN(n200) );
  INV_X1 U58 ( .A(a[3]), .ZN(n199) );
  INV_X1 U59 ( .A(n173), .ZN(n198) );
  INV_X1 U60 ( .A(a[2]), .ZN(n197) );
  INV_X1 U61 ( .A(n151), .ZN(n196) );
  INV_X1 U62 ( .A(a[1]), .ZN(n195) );
  INV_X1 U63 ( .A(n129), .ZN(n194) );
  INV_X1 U64 ( .A(a[0]), .ZN(n193) );
  OR2_X1 U65 ( .A1(n192), .A2(n212), .ZN(y[9]) );
  OR2_X1 U66 ( .A1(n211), .A2(b[9]), .ZN(n191) );
  AND2_X1 U67 ( .A1(b[9]), .A2(n211), .ZN(n192) );
  OR2_X1 U68 ( .A1(n190), .A2(n210), .ZN(y[8]) );
  OR2_X1 U69 ( .A1(n209), .A2(b[8]), .ZN(n189) );
  AND2_X1 U70 ( .A1(b[8]), .A2(n209), .ZN(n190) );
  OR2_X1 U71 ( .A1(n188), .A2(n208), .ZN(y[7]) );
  OR2_X1 U72 ( .A1(n207), .A2(b[7]), .ZN(n187) );
  AND2_X1 U73 ( .A1(b[7]), .A2(n207), .ZN(n188) );
  OR2_X1 U74 ( .A1(n186), .A2(n206), .ZN(y[6]) );
  OR2_X1 U75 ( .A1(n205), .A2(b[6]), .ZN(n185) );
  AND2_X1 U76 ( .A1(b[6]), .A2(n205), .ZN(n186) );
  OR2_X1 U77 ( .A1(n184), .A2(n204), .ZN(y[5]) );
  OR2_X1 U78 ( .A1(n203), .A2(b[5]), .ZN(n183) );
  AND2_X1 U79 ( .A1(b[5]), .A2(n203), .ZN(n184) );
  OR2_X1 U80 ( .A1(n182), .A2(n202), .ZN(y[4]) );
  OR2_X1 U81 ( .A1(n201), .A2(b[4]), .ZN(n181) );
  AND2_X1 U82 ( .A1(b[4]), .A2(n201), .ZN(n182) );
  OR2_X1 U83 ( .A1(n180), .A2(n200), .ZN(y[3]) );
  OR2_X1 U84 ( .A1(n199), .A2(b[3]), .ZN(n179) );
  AND2_X1 U85 ( .A1(b[3]), .A2(n199), .ZN(n180) );
  OR2_X1 U86 ( .A1(n178), .A2(n256), .ZN(y[31]) );
  OR2_X1 U87 ( .A1(n255), .A2(b[31]), .ZN(n177) );
  AND2_X1 U88 ( .A1(b[31]), .A2(n255), .ZN(n178) );
  OR2_X1 U89 ( .A1(n176), .A2(n254), .ZN(y[30]) );
  OR2_X1 U90 ( .A1(n253), .A2(b[30]), .ZN(n175) );
  AND2_X1 U91 ( .A1(b[30]), .A2(n253), .ZN(n176) );
  OR2_X1 U92 ( .A1(n174), .A2(n198), .ZN(y[2]) );
  OR2_X1 U93 ( .A1(n197), .A2(b[2]), .ZN(n173) );
  AND2_X1 U94 ( .A1(b[2]), .A2(n197), .ZN(n174) );
  OR2_X1 U95 ( .A1(n172), .A2(n252), .ZN(y[29]) );
  OR2_X1 U96 ( .A1(n251), .A2(b[29]), .ZN(n171) );
  AND2_X1 U97 ( .A1(b[29]), .A2(n251), .ZN(n172) );
  OR2_X1 U98 ( .A1(n170), .A2(n250), .ZN(y[28]) );
  OR2_X1 U99 ( .A1(n249), .A2(b[28]), .ZN(n169) );
  AND2_X1 U100 ( .A1(b[28]), .A2(n249), .ZN(n170) );
  OR2_X1 U101 ( .A1(n168), .A2(n248), .ZN(y[27]) );
  OR2_X1 U102 ( .A1(n247), .A2(b[27]), .ZN(n167) );
  AND2_X1 U103 ( .A1(b[27]), .A2(n247), .ZN(n168) );
  OR2_X1 U104 ( .A1(n166), .A2(n246), .ZN(y[26]) );
  OR2_X1 U105 ( .A1(n245), .A2(b[26]), .ZN(n165) );
  AND2_X1 U106 ( .A1(b[26]), .A2(n245), .ZN(n166) );
  OR2_X1 U107 ( .A1(n164), .A2(n244), .ZN(y[25]) );
  OR2_X1 U108 ( .A1(n243), .A2(b[25]), .ZN(n163) );
  AND2_X1 U109 ( .A1(b[25]), .A2(n243), .ZN(n164) );
  OR2_X1 U110 ( .A1(n162), .A2(n242), .ZN(y[24]) );
  OR2_X1 U111 ( .A1(n241), .A2(b[24]), .ZN(n161) );
  AND2_X1 U112 ( .A1(b[24]), .A2(n241), .ZN(n162) );
  OR2_X1 U113 ( .A1(n160), .A2(n240), .ZN(y[23]) );
  OR2_X1 U114 ( .A1(n239), .A2(b[23]), .ZN(n159) );
  AND2_X1 U115 ( .A1(b[23]), .A2(n239), .ZN(n160) );
  OR2_X1 U116 ( .A1(n158), .A2(n238), .ZN(y[22]) );
  OR2_X1 U117 ( .A1(n237), .A2(b[22]), .ZN(n157) );
  AND2_X1 U118 ( .A1(b[22]), .A2(n237), .ZN(n158) );
  OR2_X1 U119 ( .A1(n156), .A2(n236), .ZN(y[21]) );
  OR2_X1 U120 ( .A1(n235), .A2(b[21]), .ZN(n155) );
  AND2_X1 U121 ( .A1(b[21]), .A2(n235), .ZN(n156) );
  OR2_X1 U122 ( .A1(n154), .A2(n234), .ZN(y[20]) );
  OR2_X1 U123 ( .A1(n233), .A2(b[20]), .ZN(n153) );
  AND2_X1 U124 ( .A1(b[20]), .A2(n233), .ZN(n154) );
  OR2_X1 U125 ( .A1(n152), .A2(n196), .ZN(y[1]) );
  OR2_X1 U126 ( .A1(n195), .A2(b[1]), .ZN(n151) );
  AND2_X1 U127 ( .A1(b[1]), .A2(n195), .ZN(n152) );
  OR2_X1 U128 ( .A1(n150), .A2(n232), .ZN(y[19]) );
  OR2_X1 U129 ( .A1(n231), .A2(b[19]), .ZN(n149) );
  AND2_X1 U130 ( .A1(b[19]), .A2(n231), .ZN(n150) );
  OR2_X1 U131 ( .A1(n148), .A2(n230), .ZN(y[18]) );
  OR2_X1 U132 ( .A1(n229), .A2(b[18]), .ZN(n147) );
  AND2_X1 U133 ( .A1(b[18]), .A2(n229), .ZN(n148) );
  OR2_X1 U134 ( .A1(n146), .A2(n228), .ZN(y[17]) );
  OR2_X1 U135 ( .A1(n227), .A2(b[17]), .ZN(n145) );
  AND2_X1 U136 ( .A1(b[17]), .A2(n227), .ZN(n146) );
  OR2_X1 U137 ( .A1(n144), .A2(n226), .ZN(y[16]) );
  OR2_X1 U138 ( .A1(n225), .A2(b[16]), .ZN(n143) );
  AND2_X1 U139 ( .A1(b[16]), .A2(n225), .ZN(n144) );
  OR2_X1 U140 ( .A1(n142), .A2(n224), .ZN(y[15]) );
  OR2_X1 U141 ( .A1(n223), .A2(b[15]), .ZN(n141) );
  AND2_X1 U142 ( .A1(b[15]), .A2(n223), .ZN(n142) );
  OR2_X1 U143 ( .A1(n140), .A2(n222), .ZN(y[14]) );
  OR2_X1 U144 ( .A1(n221), .A2(b[14]), .ZN(n139) );
  AND2_X1 U145 ( .A1(b[14]), .A2(n221), .ZN(n140) );
  OR2_X1 U146 ( .A1(n138), .A2(n220), .ZN(y[13]) );
  OR2_X1 U147 ( .A1(n219), .A2(b[13]), .ZN(n137) );
  AND2_X1 U148 ( .A1(b[13]), .A2(n219), .ZN(n138) );
  OR2_X1 U149 ( .A1(n136), .A2(n218), .ZN(y[12]) );
  OR2_X1 U150 ( .A1(n217), .A2(b[12]), .ZN(n135) );
  AND2_X1 U151 ( .A1(b[12]), .A2(n217), .ZN(n136) );
  OR2_X1 U152 ( .A1(n134), .A2(n216), .ZN(y[11]) );
  OR2_X1 U153 ( .A1(n215), .A2(b[11]), .ZN(n133) );
  AND2_X1 U154 ( .A1(b[11]), .A2(n215), .ZN(n134) );
  OR2_X1 U155 ( .A1(n132), .A2(n214), .ZN(y[10]) );
  OR2_X1 U156 ( .A1(n213), .A2(b[10]), .ZN(n131) );
  AND2_X1 U157 ( .A1(b[10]), .A2(n213), .ZN(n132) );
  OR2_X1 U158 ( .A1(n130), .A2(n194), .ZN(y[0]) );
  OR2_X1 U159 ( .A1(n193), .A2(b[0]), .ZN(n129) );
  AND2_X1 U160 ( .A1(b[0]), .A2(n193), .ZN(n130) );
endmodule


module wordXor_2 ( a, b, y );
  input [31:0] a;
  input [31:0] b;
  //input_done

  output [31:0] y;
  //output_done

  wire   n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256;
  //wire_done

  INV_X1 U1 ( .A(n177), .ZN(n256) );
  INV_X1 U2 ( .A(a[31]), .ZN(n255) );
  INV_X1 U3 ( .A(n175), .ZN(n254) );
  INV_X1 U4 ( .A(a[30]), .ZN(n253) );
  INV_X1 U5 ( .A(n171), .ZN(n252) );
  INV_X1 U6 ( .A(a[29]), .ZN(n251) );
  INV_X1 U7 ( .A(n169), .ZN(n250) );
  INV_X1 U8 ( .A(a[28]), .ZN(n249) );
  INV_X1 U9 ( .A(n167), .ZN(n248) );
  INV_X1 U10 ( .A(a[27]), .ZN(n247) );
  INV_X1 U11 ( .A(n165), .ZN(n246) );
  INV_X1 U12 ( .A(a[26]), .ZN(n245) );
  INV_X1 U13 ( .A(n163), .ZN(n244) );
  INV_X1 U14 ( .A(a[25]), .ZN(n243) );
  INV_X1 U15 ( .A(n161), .ZN(n242) );
  INV_X1 U16 ( .A(a[24]), .ZN(n241) );
  INV_X1 U17 ( .A(n159), .ZN(n240) );
  INV_X1 U18 ( .A(a[23]), .ZN(n239) );
  INV_X1 U19 ( .A(n157), .ZN(n238) );
  INV_X1 U20 ( .A(a[22]), .ZN(n237) );
  INV_X1 U21 ( .A(n155), .ZN(n236) );
  INV_X1 U22 ( .A(a[21]), .ZN(n235) );
  INV_X1 U23 ( .A(n153), .ZN(n234) );
  INV_X1 U24 ( .A(a[20]), .ZN(n233) );
  INV_X1 U25 ( .A(n149), .ZN(n232) );
  INV_X1 U26 ( .A(a[19]), .ZN(n231) );
  INV_X1 U27 ( .A(n147), .ZN(n230) );
  INV_X1 U28 ( .A(a[18]), .ZN(n229) );
  INV_X1 U29 ( .A(n145), .ZN(n228) );
  INV_X1 U30 ( .A(a[17]), .ZN(n227) );
  INV_X1 U31 ( .A(n143), .ZN(n226) );
  INV_X1 U32 ( .A(a[16]), .ZN(n225) );
  INV_X1 U33 ( .A(n141), .ZN(n224) );
  INV_X1 U34 ( .A(a[15]), .ZN(n223) );
  INV_X1 U35 ( .A(n139), .ZN(n222) );
  INV_X1 U36 ( .A(a[14]), .ZN(n221) );
  INV_X1 U37 ( .A(n137), .ZN(n220) );
  INV_X1 U38 ( .A(a[13]), .ZN(n219) );
  INV_X1 U39 ( .A(n135), .ZN(n218) );
  INV_X1 U40 ( .A(a[12]), .ZN(n217) );
  INV_X1 U41 ( .A(n133), .ZN(n216) );
  INV_X1 U42 ( .A(a[11]), .ZN(n215) );
  INV_X1 U43 ( .A(n131), .ZN(n214) );
  INV_X1 U44 ( .A(a[10]), .ZN(n213) );
  INV_X1 U45 ( .A(n191), .ZN(n212) );
  INV_X1 U46 ( .A(a[9]), .ZN(n211) );
  INV_X1 U47 ( .A(n189), .ZN(n210) );
  INV_X1 U48 ( .A(a[8]), .ZN(n209) );
  INV_X1 U49 ( .A(n187), .ZN(n208) );
  INV_X1 U50 ( .A(a[7]), .ZN(n207) );
  INV_X1 U51 ( .A(n185), .ZN(n206) );
  INV_X1 U52 ( .A(a[6]), .ZN(n205) );
  INV_X1 U53 ( .A(n183), .ZN(n204) );
  INV_X1 U54 ( .A(a[5]), .ZN(n203) );
  INV_X1 U55 ( .A(n181), .ZN(n202) );
  INV_X1 U56 ( .A(a[4]), .ZN(n201) );
  INV_X1 U57 ( .A(n179), .ZN(n200) );
  INV_X1 U58 ( .A(a[3]), .ZN(n199) );
  INV_X1 U59 ( .A(n173), .ZN(n198) );
  INV_X1 U60 ( .A(a[2]), .ZN(n197) );
  INV_X1 U61 ( .A(n151), .ZN(n196) );
  INV_X1 U62 ( .A(a[1]), .ZN(n195) );
  INV_X1 U63 ( .A(n129), .ZN(n194) );
  INV_X1 U64 ( .A(a[0]), .ZN(n193) );
  OR2_X1 U65 ( .A1(n192), .A2(n212), .ZN(y[9]) );
  OR2_X1 U66 ( .A1(n211), .A2(b[9]), .ZN(n191) );
  AND2_X1 U67 ( .A1(b[9]), .A2(n211), .ZN(n192) );
  OR2_X1 U68 ( .A1(n190), .A2(n210), .ZN(y[8]) );
  OR2_X1 U69 ( .A1(n209), .A2(b[8]), .ZN(n189) );
  AND2_X1 U70 ( .A1(b[8]), .A2(n209), .ZN(n190) );
  OR2_X1 U71 ( .A1(n188), .A2(n208), .ZN(y[7]) );
  OR2_X1 U72 ( .A1(n207), .A2(b[7]), .ZN(n187) );
  AND2_X1 U73 ( .A1(b[7]), .A2(n207), .ZN(n188) );
  OR2_X1 U74 ( .A1(n186), .A2(n206), .ZN(y[6]) );
  OR2_X1 U75 ( .A1(n205), .A2(b[6]), .ZN(n185) );
  AND2_X1 U76 ( .A1(b[6]), .A2(n205), .ZN(n186) );
  OR2_X1 U77 ( .A1(n184), .A2(n204), .ZN(y[5]) );
  OR2_X1 U78 ( .A1(n203), .A2(b[5]), .ZN(n183) );
  AND2_X1 U79 ( .A1(b[5]), .A2(n203), .ZN(n184) );
  OR2_X1 U80 ( .A1(n182), .A2(n202), .ZN(y[4]) );
  OR2_X1 U81 ( .A1(n201), .A2(b[4]), .ZN(n181) );
  AND2_X1 U82 ( .A1(b[4]), .A2(n201), .ZN(n182) );
  OR2_X1 U83 ( .A1(n180), .A2(n200), .ZN(y[3]) );
  OR2_X1 U84 ( .A1(n199), .A2(b[3]), .ZN(n179) );
  AND2_X1 U85 ( .A1(b[3]), .A2(n199), .ZN(n180) );
  OR2_X1 U86 ( .A1(n178), .A2(n256), .ZN(y[31]) );
  OR2_X1 U87 ( .A1(n255), .A2(b[31]), .ZN(n177) );
  AND2_X1 U88 ( .A1(b[31]), .A2(n255), .ZN(n178) );
  OR2_X1 U89 ( .A1(n176), .A2(n254), .ZN(y[30]) );
  OR2_X1 U90 ( .A1(n253), .A2(b[30]), .ZN(n175) );
  AND2_X1 U91 ( .A1(b[30]), .A2(n253), .ZN(n176) );
  OR2_X1 U92 ( .A1(n174), .A2(n198), .ZN(y[2]) );
  OR2_X1 U93 ( .A1(n197), .A2(b[2]), .ZN(n173) );
  AND2_X1 U94 ( .A1(b[2]), .A2(n197), .ZN(n174) );
  OR2_X1 U95 ( .A1(n172), .A2(n252), .ZN(y[29]) );
  OR2_X1 U96 ( .A1(n251), .A2(b[29]), .ZN(n171) );
  AND2_X1 U97 ( .A1(b[29]), .A2(n251), .ZN(n172) );
  OR2_X1 U98 ( .A1(n170), .A2(n250), .ZN(y[28]) );
  OR2_X1 U99 ( .A1(n249), .A2(b[28]), .ZN(n169) );
  AND2_X1 U100 ( .A1(b[28]), .A2(n249), .ZN(n170) );
  OR2_X1 U101 ( .A1(n168), .A2(n248), .ZN(y[27]) );
  OR2_X1 U102 ( .A1(n247), .A2(b[27]), .ZN(n167) );
  AND2_X1 U103 ( .A1(b[27]), .A2(n247), .ZN(n168) );
  OR2_X1 U104 ( .A1(n166), .A2(n246), .ZN(y[26]) );
  OR2_X1 U105 ( .A1(n245), .A2(b[26]), .ZN(n165) );
  AND2_X1 U106 ( .A1(b[26]), .A2(n245), .ZN(n166) );
  OR2_X1 U107 ( .A1(n164), .A2(n244), .ZN(y[25]) );
  OR2_X1 U108 ( .A1(n243), .A2(b[25]), .ZN(n163) );
  AND2_X1 U109 ( .A1(b[25]), .A2(n243), .ZN(n164) );
  OR2_X1 U110 ( .A1(n162), .A2(n242), .ZN(y[24]) );
  OR2_X1 U111 ( .A1(n241), .A2(b[24]), .ZN(n161) );
  AND2_X1 U112 ( .A1(b[24]), .A2(n241), .ZN(n162) );
  OR2_X1 U113 ( .A1(n160), .A2(n240), .ZN(y[23]) );
  OR2_X1 U114 ( .A1(n239), .A2(b[23]), .ZN(n159) );
  AND2_X1 U115 ( .A1(b[23]), .A2(n239), .ZN(n160) );
  OR2_X1 U116 ( .A1(n158), .A2(n238), .ZN(y[22]) );
  OR2_X1 U117 ( .A1(n237), .A2(b[22]), .ZN(n157) );
  AND2_X1 U118 ( .A1(b[22]), .A2(n237), .ZN(n158) );
  OR2_X1 U119 ( .A1(n156), .A2(n236), .ZN(y[21]) );
  OR2_X1 U120 ( .A1(n235), .A2(b[21]), .ZN(n155) );
  AND2_X1 U121 ( .A1(b[21]), .A2(n235), .ZN(n156) );
  OR2_X1 U122 ( .A1(n154), .A2(n234), .ZN(y[20]) );
  OR2_X1 U123 ( .A1(n233), .A2(b[20]), .ZN(n153) );
  AND2_X1 U124 ( .A1(b[20]), .A2(n233), .ZN(n154) );
  OR2_X1 U125 ( .A1(n152), .A2(n196), .ZN(y[1]) );
  OR2_X1 U126 ( .A1(n195), .A2(b[1]), .ZN(n151) );
  AND2_X1 U127 ( .A1(b[1]), .A2(n195), .ZN(n152) );
  OR2_X1 U128 ( .A1(n150), .A2(n232), .ZN(y[19]) );
  OR2_X1 U129 ( .A1(n231), .A2(b[19]), .ZN(n149) );
  AND2_X1 U130 ( .A1(b[19]), .A2(n231), .ZN(n150) );
  OR2_X1 U131 ( .A1(n148), .A2(n230), .ZN(y[18]) );
  OR2_X1 U132 ( .A1(n229), .A2(b[18]), .ZN(n147) );
  AND2_X1 U133 ( .A1(b[18]), .A2(n229), .ZN(n148) );
  OR2_X1 U134 ( .A1(n146), .A2(n228), .ZN(y[17]) );
  OR2_X1 U135 ( .A1(n227), .A2(b[17]), .ZN(n145) );
  AND2_X1 U136 ( .A1(b[17]), .A2(n227), .ZN(n146) );
  OR2_X1 U137 ( .A1(n144), .A2(n226), .ZN(y[16]) );
  OR2_X1 U138 ( .A1(n225), .A2(b[16]), .ZN(n143) );
  AND2_X1 U139 ( .A1(b[16]), .A2(n225), .ZN(n144) );
  OR2_X1 U140 ( .A1(n142), .A2(n224), .ZN(y[15]) );
  OR2_X1 U141 ( .A1(n223), .A2(b[15]), .ZN(n141) );
  AND2_X1 U142 ( .A1(b[15]), .A2(n223), .ZN(n142) );
  OR2_X1 U143 ( .A1(n140), .A2(n222), .ZN(y[14]) );
  OR2_X1 U144 ( .A1(n221), .A2(b[14]), .ZN(n139) );
  AND2_X1 U145 ( .A1(b[14]), .A2(n221), .ZN(n140) );
  OR2_X1 U146 ( .A1(n138), .A2(n220), .ZN(y[13]) );
  OR2_X1 U147 ( .A1(n219), .A2(b[13]), .ZN(n137) );
  AND2_X1 U148 ( .A1(b[13]), .A2(n219), .ZN(n138) );
  OR2_X1 U149 ( .A1(n136), .A2(n218), .ZN(y[12]) );
  OR2_X1 U150 ( .A1(n217), .A2(b[12]), .ZN(n135) );
  AND2_X1 U151 ( .A1(b[12]), .A2(n217), .ZN(n136) );
  OR2_X1 U152 ( .A1(n134), .A2(n216), .ZN(y[11]) );
  OR2_X1 U153 ( .A1(n215), .A2(b[11]), .ZN(n133) );
  AND2_X1 U154 ( .A1(b[11]), .A2(n215), .ZN(n134) );
  OR2_X1 U155 ( .A1(n132), .A2(n214), .ZN(y[10]) );
  OR2_X1 U156 ( .A1(n213), .A2(b[10]), .ZN(n131) );
  AND2_X1 U157 ( .A1(b[10]), .A2(n213), .ZN(n132) );
  OR2_X1 U158 ( .A1(n130), .A2(n194), .ZN(y[0]) );
  OR2_X1 U159 ( .A1(n193), .A2(b[0]), .ZN(n129) );
  AND2_X1 U160 ( .A1(b[0]), .A2(n193), .ZN(n130) );
endmodule


module wordXor_3 ( a, b, y );
  input [31:0] a;
  input [31:0] b;
  //input_done

  output [31:0] y;
  //output_done

  wire   n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256;
  //wire_done

  INV_X1 U1 ( .A(n177), .ZN(n256) );
  INV_X1 U2 ( .A(a[31]), .ZN(n255) );
  INV_X1 U3 ( .A(n175), .ZN(n254) );
  INV_X1 U4 ( .A(a[30]), .ZN(n253) );
  INV_X1 U5 ( .A(n171), .ZN(n252) );
  INV_X1 U6 ( .A(a[29]), .ZN(n251) );
  INV_X1 U7 ( .A(n169), .ZN(n250) );
  INV_X1 U8 ( .A(a[28]), .ZN(n249) );
  INV_X1 U9 ( .A(n167), .ZN(n248) );
  INV_X1 U10 ( .A(a[27]), .ZN(n247) );
  INV_X1 U11 ( .A(n165), .ZN(n246) );
  INV_X1 U12 ( .A(a[26]), .ZN(n245) );
  INV_X1 U13 ( .A(n163), .ZN(n244) );
  INV_X1 U14 ( .A(a[25]), .ZN(n243) );
  INV_X1 U15 ( .A(n161), .ZN(n242) );
  INV_X1 U16 ( .A(a[24]), .ZN(n241) );
  INV_X1 U17 ( .A(n159), .ZN(n240) );
  INV_X1 U18 ( .A(a[23]), .ZN(n239) );
  INV_X1 U19 ( .A(n157), .ZN(n238) );
  INV_X1 U20 ( .A(a[22]), .ZN(n237) );
  INV_X1 U21 ( .A(n155), .ZN(n236) );
  INV_X1 U22 ( .A(a[21]), .ZN(n235) );
  INV_X1 U23 ( .A(n153), .ZN(n234) );
  INV_X1 U24 ( .A(a[20]), .ZN(n233) );
  INV_X1 U25 ( .A(n149), .ZN(n232) );
  INV_X1 U26 ( .A(a[19]), .ZN(n231) );
  INV_X1 U27 ( .A(n147), .ZN(n230) );
  INV_X1 U28 ( .A(a[18]), .ZN(n229) );
  INV_X1 U29 ( .A(n145), .ZN(n228) );
  INV_X1 U30 ( .A(a[17]), .ZN(n227) );
  INV_X1 U31 ( .A(n143), .ZN(n226) );
  INV_X1 U32 ( .A(a[16]), .ZN(n225) );
  INV_X1 U33 ( .A(n141), .ZN(n224) );
  INV_X1 U34 ( .A(a[15]), .ZN(n223) );
  INV_X1 U35 ( .A(n139), .ZN(n222) );
  INV_X1 U36 ( .A(a[14]), .ZN(n221) );
  INV_X1 U37 ( .A(n137), .ZN(n220) );
  INV_X1 U38 ( .A(a[13]), .ZN(n219) );
  INV_X1 U39 ( .A(n135), .ZN(n218) );
  INV_X1 U40 ( .A(a[12]), .ZN(n217) );
  INV_X1 U41 ( .A(n133), .ZN(n216) );
  INV_X1 U42 ( .A(a[11]), .ZN(n215) );
  INV_X1 U43 ( .A(n131), .ZN(n214) );
  INV_X1 U44 ( .A(a[10]), .ZN(n213) );
  INV_X1 U45 ( .A(n191), .ZN(n212) );
  INV_X1 U46 ( .A(a[9]), .ZN(n211) );
  INV_X1 U47 ( .A(n189), .ZN(n210) );
  INV_X1 U48 ( .A(a[8]), .ZN(n209) );
  INV_X1 U49 ( .A(n187), .ZN(n208) );
  INV_X1 U50 ( .A(a[7]), .ZN(n207) );
  INV_X1 U51 ( .A(n185), .ZN(n206) );
  INV_X1 U52 ( .A(a[6]), .ZN(n205) );
  INV_X1 U53 ( .A(n183), .ZN(n204) );
  INV_X1 U54 ( .A(a[5]), .ZN(n203) );
  INV_X1 U55 ( .A(n181), .ZN(n202) );
  INV_X1 U56 ( .A(a[4]), .ZN(n201) );
  INV_X1 U57 ( .A(n179), .ZN(n200) );
  INV_X1 U58 ( .A(a[3]), .ZN(n199) );
  INV_X1 U59 ( .A(n173), .ZN(n198) );
  INV_X1 U60 ( .A(a[2]), .ZN(n197) );
  INV_X1 U61 ( .A(n151), .ZN(n196) );
  INV_X1 U62 ( .A(a[1]), .ZN(n195) );
  INV_X1 U63 ( .A(n129), .ZN(n194) );
  INV_X1 U64 ( .A(a[0]), .ZN(n193) );
  OR2_X1 U65 ( .A1(n192), .A2(n212), .ZN(y[9]) );
  OR2_X1 U66 ( .A1(n211), .A2(b[9]), .ZN(n191) );
  AND2_X1 U67 ( .A1(b[9]), .A2(n211), .ZN(n192) );
  OR2_X1 U68 ( .A1(n190), .A2(n210), .ZN(y[8]) );
  OR2_X1 U69 ( .A1(n209), .A2(b[8]), .ZN(n189) );
  AND2_X1 U70 ( .A1(b[8]), .A2(n209), .ZN(n190) );
  OR2_X1 U71 ( .A1(n188), .A2(n208), .ZN(y[7]) );
  OR2_X1 U72 ( .A1(n207), .A2(b[7]), .ZN(n187) );
  AND2_X1 U73 ( .A1(b[7]), .A2(n207), .ZN(n188) );
  OR2_X1 U74 ( .A1(n186), .A2(n206), .ZN(y[6]) );
  OR2_X1 U75 ( .A1(n205), .A2(b[6]), .ZN(n185) );
  AND2_X1 U76 ( .A1(b[6]), .A2(n205), .ZN(n186) );
  OR2_X1 U77 ( .A1(n184), .A2(n204), .ZN(y[5]) );
  OR2_X1 U78 ( .A1(n203), .A2(b[5]), .ZN(n183) );
  AND2_X1 U79 ( .A1(b[5]), .A2(n203), .ZN(n184) );
  OR2_X1 U80 ( .A1(n182), .A2(n202), .ZN(y[4]) );
  OR2_X1 U81 ( .A1(n201), .A2(b[4]), .ZN(n181) );
  AND2_X1 U82 ( .A1(b[4]), .A2(n201), .ZN(n182) );
  OR2_X1 U83 ( .A1(n180), .A2(n200), .ZN(y[3]) );
  OR2_X1 U84 ( .A1(n199), .A2(b[3]), .ZN(n179) );
  AND2_X1 U85 ( .A1(b[3]), .A2(n199), .ZN(n180) );
  OR2_X1 U86 ( .A1(n178), .A2(n256), .ZN(y[31]) );
  OR2_X1 U87 ( .A1(n255), .A2(b[31]), .ZN(n177) );
  AND2_X1 U88 ( .A1(b[31]), .A2(n255), .ZN(n178) );
  OR2_X1 U89 ( .A1(n176), .A2(n254), .ZN(y[30]) );
  OR2_X1 U90 ( .A1(n253), .A2(b[30]), .ZN(n175) );
  AND2_X1 U91 ( .A1(b[30]), .A2(n253), .ZN(n176) );
  OR2_X1 U92 ( .A1(n174), .A2(n198), .ZN(y[2]) );
  OR2_X1 U93 ( .A1(n197), .A2(b[2]), .ZN(n173) );
  AND2_X1 U94 ( .A1(b[2]), .A2(n197), .ZN(n174) );
  OR2_X1 U95 ( .A1(n172), .A2(n252), .ZN(y[29]) );
  OR2_X1 U96 ( .A1(n251), .A2(b[29]), .ZN(n171) );
  AND2_X1 U97 ( .A1(b[29]), .A2(n251), .ZN(n172) );
  OR2_X1 U98 ( .A1(n170), .A2(n250), .ZN(y[28]) );
  OR2_X1 U99 ( .A1(n249), .A2(b[28]), .ZN(n169) );
  AND2_X1 U100 ( .A1(b[28]), .A2(n249), .ZN(n170) );
  OR2_X1 U101 ( .A1(n168), .A2(n248), .ZN(y[27]) );
  OR2_X1 U102 ( .A1(n247), .A2(b[27]), .ZN(n167) );
  AND2_X1 U103 ( .A1(b[27]), .A2(n247), .ZN(n168) );
  OR2_X1 U104 ( .A1(n166), .A2(n246), .ZN(y[26]) );
  OR2_X1 U105 ( .A1(n245), .A2(b[26]), .ZN(n165) );
  AND2_X1 U106 ( .A1(b[26]), .A2(n245), .ZN(n166) );
  OR2_X1 U107 ( .A1(n164), .A2(n244), .ZN(y[25]) );
  OR2_X1 U108 ( .A1(n243), .A2(b[25]), .ZN(n163) );
  AND2_X1 U109 ( .A1(b[25]), .A2(n243), .ZN(n164) );
  OR2_X1 U110 ( .A1(n162), .A2(n242), .ZN(y[24]) );
  OR2_X1 U111 ( .A1(n241), .A2(b[24]), .ZN(n161) );
  AND2_X1 U112 ( .A1(b[24]), .A2(n241), .ZN(n162) );
  OR2_X1 U113 ( .A1(n160), .A2(n240), .ZN(y[23]) );
  OR2_X1 U114 ( .A1(n239), .A2(b[23]), .ZN(n159) );
  AND2_X1 U115 ( .A1(b[23]), .A2(n239), .ZN(n160) );
  OR2_X1 U116 ( .A1(n158), .A2(n238), .ZN(y[22]) );
  OR2_X1 U117 ( .A1(n237), .A2(b[22]), .ZN(n157) );
  AND2_X1 U118 ( .A1(b[22]), .A2(n237), .ZN(n158) );
  OR2_X1 U119 ( .A1(n156), .A2(n236), .ZN(y[21]) );
  OR2_X1 U120 ( .A1(n235), .A2(b[21]), .ZN(n155) );
  AND2_X1 U121 ( .A1(b[21]), .A2(n235), .ZN(n156) );
  OR2_X1 U122 ( .A1(n154), .A2(n234), .ZN(y[20]) );
  OR2_X1 U123 ( .A1(n233), .A2(b[20]), .ZN(n153) );
  AND2_X1 U124 ( .A1(b[20]), .A2(n233), .ZN(n154) );
  OR2_X1 U125 ( .A1(n152), .A2(n196), .ZN(y[1]) );
  OR2_X1 U126 ( .A1(n195), .A2(b[1]), .ZN(n151) );
  AND2_X1 U127 ( .A1(b[1]), .A2(n195), .ZN(n152) );
  OR2_X1 U128 ( .A1(n150), .A2(n232), .ZN(y[19]) );
  OR2_X1 U129 ( .A1(n231), .A2(b[19]), .ZN(n149) );
  AND2_X1 U130 ( .A1(b[19]), .A2(n231), .ZN(n150) );
  OR2_X1 U131 ( .A1(n148), .A2(n230), .ZN(y[18]) );
  OR2_X1 U132 ( .A1(n229), .A2(b[18]), .ZN(n147) );
  AND2_X1 U133 ( .A1(b[18]), .A2(n229), .ZN(n148) );
  OR2_X1 U134 ( .A1(n146), .A2(n228), .ZN(y[17]) );
  OR2_X1 U135 ( .A1(n227), .A2(b[17]), .ZN(n145) );
  AND2_X1 U136 ( .A1(b[17]), .A2(n227), .ZN(n146) );
  OR2_X1 U137 ( .A1(n144), .A2(n226), .ZN(y[16]) );
  OR2_X1 U138 ( .A1(n225), .A2(b[16]), .ZN(n143) );
  AND2_X1 U139 ( .A1(b[16]), .A2(n225), .ZN(n144) );
  OR2_X1 U140 ( .A1(n142), .A2(n224), .ZN(y[15]) );
  OR2_X1 U141 ( .A1(n223), .A2(b[15]), .ZN(n141) );
  AND2_X1 U142 ( .A1(b[15]), .A2(n223), .ZN(n142) );
  OR2_X1 U143 ( .A1(n140), .A2(n222), .ZN(y[14]) );
  OR2_X1 U144 ( .A1(n221), .A2(b[14]), .ZN(n139) );
  AND2_X1 U145 ( .A1(b[14]), .A2(n221), .ZN(n140) );
  OR2_X1 U146 ( .A1(n138), .A2(n220), .ZN(y[13]) );
  OR2_X1 U147 ( .A1(n219), .A2(b[13]), .ZN(n137) );
  AND2_X1 U148 ( .A1(b[13]), .A2(n219), .ZN(n138) );
  OR2_X1 U149 ( .A1(n136), .A2(n218), .ZN(y[12]) );
  OR2_X1 U150 ( .A1(n217), .A2(b[12]), .ZN(n135) );
  AND2_X1 U151 ( .A1(b[12]), .A2(n217), .ZN(n136) );
  OR2_X1 U152 ( .A1(n134), .A2(n216), .ZN(y[11]) );
  OR2_X1 U153 ( .A1(n215), .A2(b[11]), .ZN(n133) );
  AND2_X1 U154 ( .A1(b[11]), .A2(n215), .ZN(n134) );
  OR2_X1 U155 ( .A1(n132), .A2(n214), .ZN(y[10]) );
  OR2_X1 U156 ( .A1(n213), .A2(b[10]), .ZN(n131) );
  AND2_X1 U157 ( .A1(b[10]), .A2(n213), .ZN(n132) );
  OR2_X1 U158 ( .A1(n130), .A2(n194), .ZN(y[0]) );
  OR2_X1 U159 ( .A1(n193), .A2(b[0]), .ZN(n129) );
  AND2_X1 U160 ( .A1(b[0]), .A2(n193), .ZN(n130) );
endmodule


module keyExpansion ( key_in, clk, firstRound, round_const, key_out );
  input [127:0] key_in;
  input [7:0] round_const;
  input clk, firstRound;
  //input_done

  output [127:0] key_out;
  //output_done
  

  wire   [127:0] key_reg;
  wire   [127:0] key;
  wire   [31:0] w3_g;
  //wire_done

  mux128_1 keyMux ( .a(key_reg), .b(key_in), .sel(firstRound), .y(key) );
  gFunction gw3 ( .in(key[31:0]), .rc(round_const), .out(w3_g) );
  wordXor_0 x0 ( .a(key[127:96]), .b(w3_g), .y(key_out[127:96]) );
  wordXor_3 x1 ( .a(key[95:64]), .b(key_out[127:96]), .y(key_out[95:64]) );
  wordXor_2 x2 ( .a(key[63:32]), .b(key_out[95:64]), .y(key_out[63:32]) );
  wordXor_1 x3 ( .a(key[31:0]), .b(key_out[63:32]), .y(key_out[31:0]) );
  DFF_X1 \key_reg_reg[0]  ( .D(key_out[0]), .CK(clk), .Q(key_reg[0]) );
  DFF_X1 \key_reg_reg[96]  ( .D(key_out[96]), .CK(clk), .Q(key_reg[96]) );
  DFF_X1 \key_reg_reg[97]  ( .D(key_out[97]), .CK(clk), .Q(key_reg[97]) );
  DFF_X1 \key_reg_reg[98]  ( .D(key_out[98]), .CK(clk), .Q(key_reg[98]) );
  DFF_X1 \key_reg_reg[99]  ( .D(key_out[99]), .CK(clk), .Q(key_reg[99]) );
  DFF_X1 \key_reg_reg[100]  ( .D(key_out[100]), .CK(clk), .Q(key_reg[100]) );
  DFF_X1 \key_reg_reg[101]  ( .D(key_out[101]), .CK(clk), .Q(key_reg[101]) );
  DFF_X1 \key_reg_reg[102]  ( .D(key_out[102]), .CK(clk), .Q(key_reg[102]) );
  DFF_X1 \key_reg_reg[103]  ( .D(key_out[103]), .CK(clk), .Q(key_reg[103]) );
  DFF_X1 \key_reg_reg[104]  ( .D(key_out[104]), .CK(clk), .Q(key_reg[104]) );
  DFF_X1 \key_reg_reg[105]  ( .D(key_out[105]), .CK(clk), .Q(key_reg[105]) );
  DFF_X1 \key_reg_reg[106]  ( .D(key_out[106]), .CK(clk), .Q(key_reg[106]) );
  DFF_X1 \key_reg_reg[107]  ( .D(key_out[107]), .CK(clk), .Q(key_reg[107]) );
  DFF_X1 \key_reg_reg[108]  ( .D(key_out[108]), .CK(clk), .Q(key_reg[108]) );
  DFF_X1 \key_reg_reg[109]  ( .D(key_out[109]), .CK(clk), .Q(key_reg[109]) );
  DFF_X1 \key_reg_reg[110]  ( .D(key_out[110]), .CK(clk), .Q(key_reg[110]) );
  DFF_X1 \key_reg_reg[111]  ( .D(key_out[111]), .CK(clk), .Q(key_reg[111]) );
  DFF_X1 \key_reg_reg[112]  ( .D(key_out[112]), .CK(clk), .Q(key_reg[112]) );
  DFF_X1 \key_reg_reg[113]  ( .D(key_out[113]), .CK(clk), .Q(key_reg[113]) );
  DFF_X1 \key_reg_reg[114]  ( .D(key_out[114]), .CK(clk), .Q(key_reg[114]) );
  DFF_X1 \key_reg_reg[115]  ( .D(key_out[115]), .CK(clk), .Q(key_reg[115]) );
  DFF_X1 \key_reg_reg[116]  ( .D(key_out[116]), .CK(clk), .Q(key_reg[116]) );
  DFF_X1 \key_reg_reg[117]  ( .D(key_out[117]), .CK(clk), .Q(key_reg[117]) );
  DFF_X1 \key_reg_reg[118]  ( .D(key_out[118]), .CK(clk), .Q(key_reg[118]) );
  DFF_X1 \key_reg_reg[119]  ( .D(key_out[119]), .CK(clk), .Q(key_reg[119]) );
  DFF_X1 \key_reg_reg[120]  ( .D(key_out[120]), .CK(clk), .Q(key_reg[120]) );
  DFF_X1 \key_reg_reg[121]  ( .D(key_out[121]), .CK(clk), .Q(key_reg[121]) );
  DFF_X1 \key_reg_reg[122]  ( .D(key_out[122]), .CK(clk), .Q(key_reg[122]) );
  DFF_X1 \key_reg_reg[123]  ( .D(key_out[123]), .CK(clk), .Q(key_reg[123]) );
  DFF_X1 \key_reg_reg[124]  ( .D(key_out[124]), .CK(clk), .Q(key_reg[124]) );
  DFF_X1 \key_reg_reg[125]  ( .D(key_out[125]), .CK(clk), .Q(key_reg[125]) );
  DFF_X1 \key_reg_reg[126]  ( .D(key_out[126]), .CK(clk), .Q(key_reg[126]) );
  DFF_X1 \key_reg_reg[127]  ( .D(key_out[127]), .CK(clk), .Q(key_reg[127]) );
  DFF_X1 \key_reg_reg[64]  ( .D(key_out[64]), .CK(clk), .Q(key_reg[64]) );
  DFF_X1 \key_reg_reg[65]  ( .D(key_out[65]), .CK(clk), .Q(key_reg[65]) );
  DFF_X1 \key_reg_reg[66]  ( .D(key_out[66]), .CK(clk), .Q(key_reg[66]) );
  DFF_X1 \key_reg_reg[67]  ( .D(key_out[67]), .CK(clk), .Q(key_reg[67]) );
  DFF_X1 \key_reg_reg[68]  ( .D(key_out[68]), .CK(clk), .Q(key_reg[68]) );
  DFF_X1 \key_reg_reg[69]  ( .D(key_out[69]), .CK(clk), .Q(key_reg[69]) );
  DFF_X1 \key_reg_reg[70]  ( .D(key_out[70]), .CK(clk), .Q(key_reg[70]) );
  DFF_X1 \key_reg_reg[71]  ( .D(key_out[71]), .CK(clk), .Q(key_reg[71]) );
  DFF_X1 \key_reg_reg[72]  ( .D(key_out[72]), .CK(clk), .Q(key_reg[72]) );
  DFF_X1 \key_reg_reg[73]  ( .D(key_out[73]), .CK(clk), .Q(key_reg[73]) );
  DFF_X1 \key_reg_reg[74]  ( .D(key_out[74]), .CK(clk), .Q(key_reg[74]) );
  DFF_X1 \key_reg_reg[75]  ( .D(key_out[75]), .CK(clk), .Q(key_reg[75]) );
  DFF_X1 \key_reg_reg[76]  ( .D(key_out[76]), .CK(clk), .Q(key_reg[76]) );
  DFF_X1 \key_reg_reg[77]  ( .D(key_out[77]), .CK(clk), .Q(key_reg[77]) );
  DFF_X1 \key_reg_reg[78]  ( .D(key_out[78]), .CK(clk), .Q(key_reg[78]) );
  DFF_X1 \key_reg_reg[79]  ( .D(key_out[79]), .CK(clk), .Q(key_reg[79]) );
  DFF_X1 \key_reg_reg[80]  ( .D(key_out[80]), .CK(clk), .Q(key_reg[80]) );
  DFF_X1 \key_reg_reg[81]  ( .D(key_out[81]), .CK(clk), .Q(key_reg[81]) );
  DFF_X1 \key_reg_reg[82]  ( .D(key_out[82]), .CK(clk), .Q(key_reg[82]) );
  DFF_X1 \key_reg_reg[83]  ( .D(key_out[83]), .CK(clk), .Q(key_reg[83]) );
  DFF_X1 \key_reg_reg[84]  ( .D(key_out[84]), .CK(clk), .Q(key_reg[84]) );
  DFF_X1 \key_reg_reg[85]  ( .D(key_out[85]), .CK(clk), .Q(key_reg[85]) );
  DFF_X1 \key_reg_reg[86]  ( .D(key_out[86]), .CK(clk), .Q(key_reg[86]) );
  DFF_X1 \key_reg_reg[87]  ( .D(key_out[87]), .CK(clk), .Q(key_reg[87]) );
  DFF_X1 \key_reg_reg[88]  ( .D(key_out[88]), .CK(clk), .Q(key_reg[88]) );
  DFF_X1 \key_reg_reg[89]  ( .D(key_out[89]), .CK(clk), .Q(key_reg[89]) );
  DFF_X1 \key_reg_reg[90]  ( .D(key_out[90]), .CK(clk), .Q(key_reg[90]) );
  DFF_X1 \key_reg_reg[91]  ( .D(key_out[91]), .CK(clk), .Q(key_reg[91]) );
  DFF_X1 \key_reg_reg[92]  ( .D(key_out[92]), .CK(clk), .Q(key_reg[92]) );
  DFF_X1 \key_reg_reg[93]  ( .D(key_out[93]), .CK(clk), .Q(key_reg[93]) );
  DFF_X1 \key_reg_reg[94]  ( .D(key_out[94]), .CK(clk), .Q(key_reg[94]) );
  DFF_X1 \key_reg_reg[95]  ( .D(key_out[95]), .CK(clk), .Q(key_reg[95]) );
  DFF_X1 \key_reg_reg[32]  ( .D(key_out[32]), .CK(clk), .Q(key_reg[32]) );
  DFF_X1 \key_reg_reg[33]  ( .D(key_out[33]), .CK(clk), .Q(key_reg[33]) );
  DFF_X1 \key_reg_reg[34]  ( .D(key_out[34]), .CK(clk), .Q(key_reg[34]) );
  DFF_X1 \key_reg_reg[35]  ( .D(key_out[35]), .CK(clk), .Q(key_reg[35]) );
  DFF_X1 \key_reg_reg[36]  ( .D(key_out[36]), .CK(clk), .Q(key_reg[36]) );
  DFF_X1 \key_reg_reg[37]  ( .D(key_out[37]), .CK(clk), .Q(key_reg[37]) );
  DFF_X1 \key_reg_reg[38]  ( .D(key_out[38]), .CK(clk), .Q(key_reg[38]) );
  DFF_X1 \key_reg_reg[39]  ( .D(key_out[39]), .CK(clk), .Q(key_reg[39]) );
  DFF_X1 \key_reg_reg[40]  ( .D(key_out[40]), .CK(clk), .Q(key_reg[40]) );
  DFF_X1 \key_reg_reg[41]  ( .D(key_out[41]), .CK(clk), .Q(key_reg[41]) );
  DFF_X1 \key_reg_reg[42]  ( .D(key_out[42]), .CK(clk), .Q(key_reg[42]) );
  DFF_X1 \key_reg_reg[43]  ( .D(key_out[43]), .CK(clk), .Q(key_reg[43]) );
  DFF_X1 \key_reg_reg[44]  ( .D(key_out[44]), .CK(clk), .Q(key_reg[44]) );
  DFF_X1 \key_reg_reg[45]  ( .D(key_out[45]), .CK(clk), .Q(key_reg[45]) );
  DFF_X1 \key_reg_reg[46]  ( .D(key_out[46]), .CK(clk), .Q(key_reg[46]) );
  DFF_X1 \key_reg_reg[47]  ( .D(key_out[47]), .CK(clk), .Q(key_reg[47]) );
  DFF_X1 \key_reg_reg[48]  ( .D(key_out[48]), .CK(clk), .Q(key_reg[48]) );
  DFF_X1 \key_reg_reg[49]  ( .D(key_out[49]), .CK(clk), .Q(key_reg[49]) );
  DFF_X1 \key_reg_reg[50]  ( .D(key_out[50]), .CK(clk), .Q(key_reg[50]) );
  DFF_X1 \key_reg_reg[51]  ( .D(key_out[51]), .CK(clk), .Q(key_reg[51]) );
  DFF_X1 \key_reg_reg[52]  ( .D(key_out[52]), .CK(clk), .Q(key_reg[52]) );
  DFF_X1 \key_reg_reg[53]  ( .D(key_out[53]), .CK(clk), .Q(key_reg[53]) );
  DFF_X1 \key_reg_reg[54]  ( .D(key_out[54]), .CK(clk), .Q(key_reg[54]) );
  DFF_X1 \key_reg_reg[55]  ( .D(key_out[55]), .CK(clk), .Q(key_reg[55]) );
  DFF_X1 \key_reg_reg[56]  ( .D(key_out[56]), .CK(clk), .Q(key_reg[56]) );
  DFF_X1 \key_reg_reg[57]  ( .D(key_out[57]), .CK(clk), .Q(key_reg[57]) );
  DFF_X1 \key_reg_reg[58]  ( .D(key_out[58]), .CK(clk), .Q(key_reg[58]) );
  DFF_X1 \key_reg_reg[59]  ( .D(key_out[59]), .CK(clk), .Q(key_reg[59]) );
  DFF_X1 \key_reg_reg[60]  ( .D(key_out[60]), .CK(clk), .Q(key_reg[60]) );
  DFF_X1 \key_reg_reg[61]  ( .D(key_out[61]), .CK(clk), .Q(key_reg[61]) );
  DFF_X1 \key_reg_reg[62]  ( .D(key_out[62]), .CK(clk), .Q(key_reg[62]) );
  DFF_X1 \key_reg_reg[63]  ( .D(key_out[63]), .CK(clk), .Q(key_reg[63]) );
  DFF_X1 \key_reg_reg[1]  ( .D(key_out[1]), .CK(clk), .Q(key_reg[1]) );
  DFF_X1 \key_reg_reg[2]  ( .D(key_out[2]), .CK(clk), .Q(key_reg[2]) );
  DFF_X1 \key_reg_reg[3]  ( .D(key_out[3]), .CK(clk), .Q(key_reg[3]) );
  DFF_X1 \key_reg_reg[4]  ( .D(key_out[4]), .CK(clk), .Q(key_reg[4]) );
  DFF_X1 \key_reg_reg[5]  ( .D(key_out[5]), .CK(clk), .Q(key_reg[5]) );
  DFF_X1 \key_reg_reg[6]  ( .D(key_out[6]), .CK(clk), .Q(key_reg[6]) );
  DFF_X1 \key_reg_reg[7]  ( .D(key_out[7]), .CK(clk), .Q(key_reg[7]) );
  DFF_X1 \key_reg_reg[8]  ( .D(key_out[8]), .CK(clk), .Q(key_reg[8]) );
  DFF_X1 \key_reg_reg[9]  ( .D(key_out[9]), .CK(clk), .Q(key_reg[9]) );
  DFF_X1 \key_reg_reg[10]  ( .D(key_out[10]), .CK(clk), .Q(key_reg[10]) );
  DFF_X1 \key_reg_reg[11]  ( .D(key_out[11]), .CK(clk), .Q(key_reg[11]) );
  DFF_X1 \key_reg_reg[12]  ( .D(key_out[12]), .CK(clk), .Q(key_reg[12]) );
  DFF_X1 \key_reg_reg[13]  ( .D(key_out[13]), .CK(clk), .Q(key_reg[13]) );
  DFF_X1 \key_reg_reg[14]  ( .D(key_out[14]), .CK(clk), .Q(key_reg[14]) );
  DFF_X1 \key_reg_reg[15]  ( .D(key_out[15]), .CK(clk), .Q(key_reg[15]) );
  DFF_X1 \key_reg_reg[16]  ( .D(key_out[16]), .CK(clk), .Q(key_reg[16]) );
  DFF_X1 \key_reg_reg[17]  ( .D(key_out[17]), .CK(clk), .Q(key_reg[17]) );
  DFF_X1 \key_reg_reg[18]  ( .D(key_out[18]), .CK(clk), .Q(key_reg[18]) );
  DFF_X1 \key_reg_reg[19]  ( .D(key_out[19]), .CK(clk), .Q(key_reg[19]) );
  DFF_X1 \key_reg_reg[20]  ( .D(key_out[20]), .CK(clk), .Q(key_reg[20]) );
  DFF_X1 \key_reg_reg[21]  ( .D(key_out[21]), .CK(clk), .Q(key_reg[21]) );
  DFF_X1 \key_reg_reg[22]  ( .D(key_out[22]), .CK(clk), .Q(key_reg[22]) );
  DFF_X1 \key_reg_reg[23]  ( .D(key_out[23]), .CK(clk), .Q(key_reg[23]) );
  DFF_X1 \key_reg_reg[24]  ( .D(key_out[24]), .CK(clk), .Q(key_reg[24]) );
  DFF_X1 \key_reg_reg[25]  ( .D(key_out[25]), .CK(clk), .Q(key_reg[25]) );
  DFF_X1 \key_reg_reg[26]  ( .D(key_out[26]), .CK(clk), .Q(key_reg[26]) );
  DFF_X1 \key_reg_reg[27]  ( .D(key_out[27]), .CK(clk), .Q(key_reg[27]) );
  DFF_X1 \key_reg_reg[28]  ( .D(key_out[28]), .CK(clk), .Q(key_reg[28]) );
  DFF_X1 \key_reg_reg[29]  ( .D(key_out[29]), .CK(clk), .Q(key_reg[29]) );
  DFF_X1 \key_reg_reg[30]  ( .D(key_out[30]), .CK(clk), .Q(key_reg[30]) );
  DFF_X1 \key_reg_reg[31]  ( .D(key_out[31]), .CK(clk), .Q(key_reg[31]) );
endmodule


module addKey ( data, key, out );
  input [127:0] data;
  input [127:0] key;
  //input_done

  output [127:0] out;
  //output_done

  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512;
  //wire_done

  INV_X1 U1 ( .A(n452), .ZN(n1) );
  INV_X1 U2 ( .A(data[127]), .ZN(n2) );
  INV_X1 U3 ( .A(n454), .ZN(n3) );
  INV_X1 U4 ( .A(data[126]), .ZN(n4) );
  INV_X1 U5 ( .A(n456), .ZN(n5) );
  INV_X1 U6 ( .A(data[125]), .ZN(n6) );
  INV_X1 U7 ( .A(n458), .ZN(n7) );
  INV_X1 U8 ( .A(data[124]), .ZN(n8) );
  INV_X1 U9 ( .A(n460), .ZN(n9) );
  INV_X1 U10 ( .A(data[123]), .ZN(n10) );
  INV_X1 U11 ( .A(n462), .ZN(n11) );
  INV_X1 U12 ( .A(data[122]), .ZN(n12) );
  INV_X1 U13 ( .A(n464), .ZN(n13) );
  INV_X1 U14 ( .A(data[121]), .ZN(n14) );
  INV_X1 U15 ( .A(n466), .ZN(n15) );
  INV_X1 U16 ( .A(data[120]), .ZN(n16) );
  INV_X1 U17 ( .A(n470), .ZN(n17) );
  INV_X1 U18 ( .A(data[119]), .ZN(n18) );
  INV_X1 U19 ( .A(n472), .ZN(n19) );
  INV_X1 U20 ( .A(data[118]), .ZN(n20) );
  INV_X1 U21 ( .A(n474), .ZN(n21) );
  INV_X1 U22 ( .A(data[117]), .ZN(n22) );
  INV_X1 U23 ( .A(n476), .ZN(n23) );
  INV_X1 U24 ( .A(data[116]), .ZN(n24) );
  INV_X1 U25 ( .A(n478), .ZN(n25) );
  INV_X1 U26 ( .A(data[115]), .ZN(n26) );
  INV_X1 U27 ( .A(n480), .ZN(n27) );
  INV_X1 U28 ( .A(data[114]), .ZN(n28) );
  INV_X1 U29 ( .A(n482), .ZN(n29) );
  INV_X1 U30 ( .A(data[113]), .ZN(n30) );
  INV_X1 U31 ( .A(n484), .ZN(n31) );
  INV_X1 U32 ( .A(data[112]), .ZN(n32) );
  INV_X1 U33 ( .A(n486), .ZN(n33) );
  INV_X1 U34 ( .A(data[111]), .ZN(n34) );
  INV_X1 U35 ( .A(n488), .ZN(n35) );
  INV_X1 U36 ( .A(data[110]), .ZN(n36) );
  INV_X1 U37 ( .A(n492), .ZN(n37) );
  INV_X1 U38 ( .A(data[109]), .ZN(n38) );
  INV_X1 U39 ( .A(n494), .ZN(n39) );
  INV_X1 U40 ( .A(data[108]), .ZN(n40) );
  INV_X1 U41 ( .A(n496), .ZN(n41) );
  INV_X1 U42 ( .A(data[107]), .ZN(n42) );
  INV_X1 U43 ( .A(n498), .ZN(n43) );
  INV_X1 U44 ( .A(data[106]), .ZN(n44) );
  INV_X1 U45 ( .A(n500), .ZN(n45) );
  INV_X1 U46 ( .A(data[105]), .ZN(n46) );
  INV_X1 U47 ( .A(n502), .ZN(n47) );
  INV_X1 U48 ( .A(data[104]), .ZN(n48) );
  INV_X1 U49 ( .A(n504), .ZN(n49) );
  INV_X1 U50 ( .A(data[103]), .ZN(n50) );
  INV_X1 U51 ( .A(n506), .ZN(n51) );
  INV_X1 U52 ( .A(data[102]), .ZN(n52) );
  INV_X1 U53 ( .A(n508), .ZN(n53) );
  INV_X1 U54 ( .A(data[101]), .ZN(n54) );
  INV_X1 U55 ( .A(n510), .ZN(n55) );
  INV_X1 U56 ( .A(data[100]), .ZN(n56) );
  INV_X1 U57 ( .A(n260), .ZN(n57) );
  INV_X1 U58 ( .A(data[99]), .ZN(n58) );
  INV_X1 U59 ( .A(n262), .ZN(n59) );
  INV_X1 U60 ( .A(data[98]), .ZN(n60) );
  INV_X1 U61 ( .A(n264), .ZN(n61) );
  INV_X1 U62 ( .A(data[97]), .ZN(n62) );
  INV_X1 U63 ( .A(n266), .ZN(n63) );
  INV_X1 U64 ( .A(data[96]), .ZN(n64) );
  INV_X1 U65 ( .A(n268), .ZN(n65) );
  INV_X1 U66 ( .A(data[95]), .ZN(n66) );
  INV_X1 U67 ( .A(n270), .ZN(n67) );
  INV_X1 U68 ( .A(data[94]), .ZN(n68) );
  INV_X1 U69 ( .A(n272), .ZN(n69) );
  INV_X1 U70 ( .A(data[93]), .ZN(n70) );
  INV_X1 U71 ( .A(n274), .ZN(n71) );
  INV_X1 U72 ( .A(data[92]), .ZN(n72) );
  INV_X1 U73 ( .A(n276), .ZN(n73) );
  INV_X1 U74 ( .A(data[91]), .ZN(n74) );
  INV_X1 U75 ( .A(n278), .ZN(n75) );
  INV_X1 U76 ( .A(data[90]), .ZN(n76) );
  INV_X1 U77 ( .A(n282), .ZN(n77) );
  INV_X1 U78 ( .A(data[89]), .ZN(n78) );
  INV_X1 U79 ( .A(n284), .ZN(n79) );
  INV_X1 U80 ( .A(data[88]), .ZN(n80) );
  INV_X1 U81 ( .A(n286), .ZN(n81) );
  INV_X1 U82 ( .A(data[87]), .ZN(n82) );
  INV_X1 U83 ( .A(n288), .ZN(n83) );
  INV_X1 U84 ( .A(data[86]), .ZN(n84) );
  INV_X1 U85 ( .A(n290), .ZN(n85) );
  INV_X1 U86 ( .A(data[85]), .ZN(n86) );
  INV_X1 U87 ( .A(n292), .ZN(n87) );
  INV_X1 U88 ( .A(data[84]), .ZN(n88) );
  INV_X1 U89 ( .A(n294), .ZN(n89) );
  INV_X1 U90 ( .A(data[83]), .ZN(n90) );
  INV_X1 U91 ( .A(n296), .ZN(n91) );
  INV_X1 U92 ( .A(data[82]), .ZN(n92) );
  INV_X1 U93 ( .A(n298), .ZN(n93) );
  INV_X1 U94 ( .A(data[81]), .ZN(n94) );
  INV_X1 U95 ( .A(n300), .ZN(n95) );
  INV_X1 U96 ( .A(data[80]), .ZN(n96) );
  INV_X1 U97 ( .A(n304), .ZN(n97) );
  INV_X1 U98 ( .A(data[79]), .ZN(n98) );
  INV_X1 U99 ( .A(n306), .ZN(n99) );
  INV_X1 U100 ( .A(data[78]), .ZN(n100) );
  INV_X1 U101 ( .A(n308), .ZN(n101) );
  INV_X1 U102 ( .A(data[77]), .ZN(n102) );
  INV_X1 U103 ( .A(n310), .ZN(n103) );
  INV_X1 U104 ( .A(data[76]), .ZN(n104) );
  INV_X1 U105 ( .A(n312), .ZN(n105) );
  INV_X1 U106 ( .A(data[75]), .ZN(n106) );
  INV_X1 U107 ( .A(n314), .ZN(n107) );
  INV_X1 U108 ( .A(data[74]), .ZN(n108) );
  INV_X1 U109 ( .A(n316), .ZN(n109) );
  INV_X1 U110 ( .A(data[73]), .ZN(n110) );
  INV_X1 U111 ( .A(n318), .ZN(n111) );
  INV_X1 U112 ( .A(data[72]), .ZN(n112) );
  INV_X1 U113 ( .A(n320), .ZN(n113) );
  INV_X1 U114 ( .A(data[71]), .ZN(n114) );
  INV_X1 U115 ( .A(n322), .ZN(n115) );
  INV_X1 U116 ( .A(data[70]), .ZN(n116) );
  INV_X1 U117 ( .A(n326), .ZN(n117) );
  INV_X1 U118 ( .A(data[69]), .ZN(n118) );
  INV_X1 U119 ( .A(n328), .ZN(n119) );
  INV_X1 U120 ( .A(data[68]), .ZN(n120) );
  INV_X1 U121 ( .A(n330), .ZN(n121) );
  INV_X1 U122 ( .A(data[67]), .ZN(n122) );
  INV_X1 U123 ( .A(n332), .ZN(n123) );
  INV_X1 U124 ( .A(data[66]), .ZN(n124) );
  INV_X1 U125 ( .A(n334), .ZN(n125) );
  INV_X1 U126 ( .A(data[65]), .ZN(n126) );
  INV_X1 U127 ( .A(n336), .ZN(n127) );
  INV_X1 U128 ( .A(data[64]), .ZN(n128) );
  INV_X1 U129 ( .A(n338), .ZN(n129) );
  INV_X1 U130 ( .A(data[63]), .ZN(n130) );
  INV_X1 U131 ( .A(n340), .ZN(n131) );
  INV_X1 U132 ( .A(data[62]), .ZN(n132) );
  INV_X1 U133 ( .A(n342), .ZN(n133) );
  INV_X1 U134 ( .A(data[61]), .ZN(n134) );
  INV_X1 U135 ( .A(n344), .ZN(n135) );
  INV_X1 U136 ( .A(data[60]), .ZN(n136) );
  INV_X1 U137 ( .A(n348), .ZN(n137) );
  INV_X1 U138 ( .A(data[59]), .ZN(n138) );
  INV_X1 U139 ( .A(n350), .ZN(n139) );
  INV_X1 U140 ( .A(data[58]), .ZN(n140) );
  INV_X1 U141 ( .A(n352), .ZN(n141) );
  INV_X1 U142 ( .A(data[57]), .ZN(n142) );
  INV_X1 U143 ( .A(n354), .ZN(n143) );
  INV_X1 U144 ( .A(data[56]), .ZN(n144) );
  INV_X1 U145 ( .A(n356), .ZN(n145) );
  INV_X1 U146 ( .A(data[55]), .ZN(n146) );
  INV_X1 U147 ( .A(n358), .ZN(n147) );
  INV_X1 U148 ( .A(data[54]), .ZN(n148) );
  INV_X1 U149 ( .A(n360), .ZN(n149) );
  INV_X1 U150 ( .A(data[53]), .ZN(n150) );
  INV_X1 U151 ( .A(n362), .ZN(n151) );
  INV_X1 U152 ( .A(data[52]), .ZN(n152) );
  INV_X1 U153 ( .A(n364), .ZN(n153) );
  INV_X1 U154 ( .A(data[51]), .ZN(n154) );
  INV_X1 U155 ( .A(n366), .ZN(n155) );
  INV_X1 U156 ( .A(data[50]), .ZN(n156) );
  INV_X1 U157 ( .A(n370), .ZN(n157) );
  INV_X1 U158 ( .A(data[49]), .ZN(n158) );
  INV_X1 U159 ( .A(n372), .ZN(n159) );
  INV_X1 U160 ( .A(data[48]), .ZN(n160) );
  INV_X1 U161 ( .A(n374), .ZN(n161) );
  INV_X1 U162 ( .A(data[47]), .ZN(n162) );
  INV_X1 U163 ( .A(n376), .ZN(n163) );
  INV_X1 U164 ( .A(data[46]), .ZN(n164) );
  INV_X1 U165 ( .A(n378), .ZN(n165) );
  INV_X1 U166 ( .A(data[45]), .ZN(n166) );
  INV_X1 U167 ( .A(n380), .ZN(n167) );
  INV_X1 U168 ( .A(data[44]), .ZN(n168) );
  INV_X1 U169 ( .A(n382), .ZN(n169) );
  INV_X1 U170 ( .A(data[43]), .ZN(n170) );
  INV_X1 U171 ( .A(n384), .ZN(n171) );
  INV_X1 U172 ( .A(data[42]), .ZN(n172) );
  INV_X1 U173 ( .A(n386), .ZN(n173) );
  INV_X1 U174 ( .A(data[41]), .ZN(n174) );
  INV_X1 U175 ( .A(n388), .ZN(n175) );
  INV_X1 U176 ( .A(data[40]), .ZN(n176) );
  INV_X1 U177 ( .A(n392), .ZN(n177) );
  INV_X1 U178 ( .A(data[39]), .ZN(n178) );
  INV_X1 U179 ( .A(n394), .ZN(n179) );
  INV_X1 U180 ( .A(data[38]), .ZN(n180) );
  INV_X1 U181 ( .A(n396), .ZN(n181) );
  INV_X1 U182 ( .A(data[37]), .ZN(n182) );
  INV_X1 U183 ( .A(n398), .ZN(n183) );
  INV_X1 U184 ( .A(data[36]), .ZN(n184) );
  INV_X1 U185 ( .A(n400), .ZN(n185) );
  INV_X1 U186 ( .A(data[35]), .ZN(n186) );
  INV_X1 U187 ( .A(n402), .ZN(n187) );
  INV_X1 U188 ( .A(data[34]), .ZN(n188) );
  INV_X1 U189 ( .A(n404), .ZN(n189) );
  INV_X1 U190 ( .A(data[33]), .ZN(n190) );
  INV_X1 U191 ( .A(n406), .ZN(n191) );
  INV_X1 U192 ( .A(data[32]), .ZN(n192) );
  INV_X1 U193 ( .A(n408), .ZN(n193) );
  INV_X1 U194 ( .A(data[31]), .ZN(n194) );
  INV_X1 U195 ( .A(n410), .ZN(n195) );
  INV_X1 U196 ( .A(data[30]), .ZN(n196) );
  INV_X1 U197 ( .A(n414), .ZN(n197) );
  INV_X1 U198 ( .A(data[29]), .ZN(n198) );
  INV_X1 U199 ( .A(n416), .ZN(n199) );
  INV_X1 U200 ( .A(data[28]), .ZN(n200) );
  INV_X1 U201 ( .A(n418), .ZN(n201) );
  INV_X1 U202 ( .A(data[27]), .ZN(n202) );
  INV_X1 U203 ( .A(n420), .ZN(n203) );
  INV_X1 U204 ( .A(data[26]), .ZN(n204) );
  INV_X1 U205 ( .A(n422), .ZN(n205) );
  INV_X1 U206 ( .A(data[25]), .ZN(n206) );
  INV_X1 U207 ( .A(n424), .ZN(n207) );
  INV_X1 U208 ( .A(data[24]), .ZN(n208) );
  INV_X1 U209 ( .A(n426), .ZN(n209) );
  INV_X1 U210 ( .A(data[23]), .ZN(n210) );
  INV_X1 U211 ( .A(n428), .ZN(n211) );
  INV_X1 U212 ( .A(data[22]), .ZN(n212) );
  INV_X1 U213 ( .A(n430), .ZN(n213) );
  INV_X1 U214 ( .A(data[21]), .ZN(n214) );
  INV_X1 U215 ( .A(n432), .ZN(n215) );
  INV_X1 U216 ( .A(data[20]), .ZN(n216) );
  INV_X1 U217 ( .A(n436), .ZN(n217) );
  INV_X1 U218 ( .A(data[19]), .ZN(n218) );
  INV_X1 U219 ( .A(n438), .ZN(n219) );
  INV_X1 U220 ( .A(data[18]), .ZN(n220) );
  INV_X1 U221 ( .A(n440), .ZN(n221) );
  INV_X1 U222 ( .A(data[17]), .ZN(n222) );
  INV_X1 U223 ( .A(n442), .ZN(n223) );
  INV_X1 U224 ( .A(data[16]), .ZN(n224) );
  INV_X1 U225 ( .A(n444), .ZN(n225) );
  INV_X1 U226 ( .A(data[15]), .ZN(n226) );
  INV_X1 U227 ( .A(n446), .ZN(n227) );
  INV_X1 U228 ( .A(data[14]), .ZN(n228) );
  INV_X1 U229 ( .A(n448), .ZN(n229) );
  INV_X1 U230 ( .A(data[13]), .ZN(n230) );
  INV_X1 U231 ( .A(n450), .ZN(n231) );
  INV_X1 U232 ( .A(data[12]), .ZN(n232) );
  INV_X1 U233 ( .A(n468), .ZN(n233) );
  INV_X1 U234 ( .A(data[11]), .ZN(n234) );
  INV_X1 U235 ( .A(n490), .ZN(n235) );
  INV_X1 U236 ( .A(data[10]), .ZN(n236) );
  INV_X1 U237 ( .A(n258), .ZN(n237) );
  INV_X1 U238 ( .A(data[9]), .ZN(n238) );
  INV_X1 U239 ( .A(n280), .ZN(n239) );
  INV_X1 U240 ( .A(data[8]), .ZN(n240) );
  INV_X1 U241 ( .A(n302), .ZN(n241) );
  INV_X1 U242 ( .A(data[7]), .ZN(n242) );
  INV_X1 U243 ( .A(n324), .ZN(n243) );
  INV_X1 U244 ( .A(data[6]), .ZN(n244) );
  INV_X1 U245 ( .A(n346), .ZN(n245) );
  INV_X1 U246 ( .A(data[5]), .ZN(n246) );
  INV_X1 U247 ( .A(n368), .ZN(n247) );
  INV_X1 U248 ( .A(data[4]), .ZN(n248) );
  INV_X1 U249 ( .A(n390), .ZN(n249) );
  INV_X1 U250 ( .A(data[3]), .ZN(n250) );
  INV_X1 U251 ( .A(n412), .ZN(n251) );
  INV_X1 U252 ( .A(data[2]), .ZN(n252) );
  INV_X1 U253 ( .A(n434), .ZN(n253) );
  INV_X1 U254 ( .A(data[1]), .ZN(n254) );
  INV_X1 U255 ( .A(n512), .ZN(n255) );
  INV_X1 U256 ( .A(data[0]), .ZN(n256) );
  OR2_X1 U257 ( .A1(n257), .A2(n237), .ZN(out[9]) );
  OR2_X1 U258 ( .A1(n238), .A2(key[9]), .ZN(n258) );
  AND2_X1 U259 ( .A1(key[9]), .A2(n238), .ZN(n257) );
  OR2_X1 U260 ( .A1(n259), .A2(n57), .ZN(out[99]) );
  OR2_X1 U261 ( .A1(n58), .A2(key[99]), .ZN(n260) );
  AND2_X1 U262 ( .A1(key[99]), .A2(n58), .ZN(n259) );
  OR2_X1 U263 ( .A1(n261), .A2(n59), .ZN(out[98]) );
  OR2_X1 U264 ( .A1(n60), .A2(key[98]), .ZN(n262) );
  AND2_X1 U265 ( .A1(key[98]), .A2(n60), .ZN(n261) );
  OR2_X1 U266 ( .A1(n263), .A2(n61), .ZN(out[97]) );
  OR2_X1 U267 ( .A1(n62), .A2(key[97]), .ZN(n264) );
  AND2_X1 U268 ( .A1(key[97]), .A2(n62), .ZN(n263) );
  OR2_X1 U269 ( .A1(n265), .A2(n63), .ZN(out[96]) );
  OR2_X1 U270 ( .A1(n64), .A2(key[96]), .ZN(n266) );
  AND2_X1 U271 ( .A1(key[96]), .A2(n64), .ZN(n265) );
  OR2_X1 U272 ( .A1(n267), .A2(n65), .ZN(out[95]) );
  OR2_X1 U273 ( .A1(n66), .A2(key[95]), .ZN(n268) );
  AND2_X1 U274 ( .A1(key[95]), .A2(n66), .ZN(n267) );
  OR2_X1 U275 ( .A1(n269), .A2(n67), .ZN(out[94]) );
  OR2_X1 U276 ( .A1(n68), .A2(key[94]), .ZN(n270) );
  AND2_X1 U277 ( .A1(key[94]), .A2(n68), .ZN(n269) );
  OR2_X1 U278 ( .A1(n271), .A2(n69), .ZN(out[93]) );
  OR2_X1 U279 ( .A1(n70), .A2(key[93]), .ZN(n272) );
  AND2_X1 U280 ( .A1(key[93]), .A2(n70), .ZN(n271) );
  OR2_X1 U281 ( .A1(n273), .A2(n71), .ZN(out[92]) );
  OR2_X1 U282 ( .A1(n72), .A2(key[92]), .ZN(n274) );
  AND2_X1 U283 ( .A1(key[92]), .A2(n72), .ZN(n273) );
  OR2_X1 U284 ( .A1(n275), .A2(n73), .ZN(out[91]) );
  OR2_X1 U285 ( .A1(n74), .A2(key[91]), .ZN(n276) );
  AND2_X1 U286 ( .A1(key[91]), .A2(n74), .ZN(n275) );
  OR2_X1 U287 ( .A1(n277), .A2(n75), .ZN(out[90]) );
  OR2_X1 U288 ( .A1(n76), .A2(key[90]), .ZN(n278) );
  AND2_X1 U289 ( .A1(key[90]), .A2(n76), .ZN(n277) );
  OR2_X1 U290 ( .A1(n279), .A2(n239), .ZN(out[8]) );
  OR2_X1 U291 ( .A1(n240), .A2(key[8]), .ZN(n280) );
  AND2_X1 U292 ( .A1(key[8]), .A2(n240), .ZN(n279) );
  OR2_X1 U293 ( .A1(n281), .A2(n77), .ZN(out[89]) );
  OR2_X1 U294 ( .A1(n78), .A2(key[89]), .ZN(n282) );
  AND2_X1 U295 ( .A1(key[89]), .A2(n78), .ZN(n281) );
  OR2_X1 U296 ( .A1(n283), .A2(n79), .ZN(out[88]) );
  OR2_X1 U297 ( .A1(n80), .A2(key[88]), .ZN(n284) );
  AND2_X1 U298 ( .A1(key[88]), .A2(n80), .ZN(n283) );
  OR2_X1 U299 ( .A1(n285), .A2(n81), .ZN(out[87]) );
  OR2_X1 U300 ( .A1(n82), .A2(key[87]), .ZN(n286) );
  AND2_X1 U301 ( .A1(key[87]), .A2(n82), .ZN(n285) );
  OR2_X1 U302 ( .A1(n287), .A2(n83), .ZN(out[86]) );
  OR2_X1 U303 ( .A1(n84), .A2(key[86]), .ZN(n288) );
  AND2_X1 U304 ( .A1(key[86]), .A2(n84), .ZN(n287) );
  OR2_X1 U305 ( .A1(n289), .A2(n85), .ZN(out[85]) );
  OR2_X1 U306 ( .A1(n86), .A2(key[85]), .ZN(n290) );
  AND2_X1 U307 ( .A1(key[85]), .A2(n86), .ZN(n289) );
  OR2_X1 U308 ( .A1(n291), .A2(n87), .ZN(out[84]) );
  OR2_X1 U309 ( .A1(n88), .A2(key[84]), .ZN(n292) );
  AND2_X1 U310 ( .A1(key[84]), .A2(n88), .ZN(n291) );
  OR2_X1 U311 ( .A1(n293), .A2(n89), .ZN(out[83]) );
  OR2_X1 U312 ( .A1(n90), .A2(key[83]), .ZN(n294) );
  AND2_X1 U313 ( .A1(key[83]), .A2(n90), .ZN(n293) );
  OR2_X1 U314 ( .A1(n295), .A2(n91), .ZN(out[82]) );
  OR2_X1 U315 ( .A1(n92), .A2(key[82]), .ZN(n296) );
  AND2_X1 U316 ( .A1(key[82]), .A2(n92), .ZN(n295) );
  OR2_X1 U317 ( .A1(n297), .A2(n93), .ZN(out[81]) );
  OR2_X1 U318 ( .A1(n94), .A2(key[81]), .ZN(n298) );
  AND2_X1 U319 ( .A1(key[81]), .A2(n94), .ZN(n297) );
  OR2_X1 U320 ( .A1(n299), .A2(n95), .ZN(out[80]) );
  OR2_X1 U321 ( .A1(n96), .A2(key[80]), .ZN(n300) );
  AND2_X1 U322 ( .A1(key[80]), .A2(n96), .ZN(n299) );
  OR2_X1 U323 ( .A1(n301), .A2(n241), .ZN(out[7]) );
  OR2_X1 U324 ( .A1(n242), .A2(key[7]), .ZN(n302) );
  AND2_X1 U325 ( .A1(key[7]), .A2(n242), .ZN(n301) );
  OR2_X1 U326 ( .A1(n303), .A2(n97), .ZN(out[79]) );
  OR2_X1 U327 ( .A1(n98), .A2(key[79]), .ZN(n304) );
  AND2_X1 U328 ( .A1(key[79]), .A2(n98), .ZN(n303) );
  OR2_X1 U329 ( .A1(n305), .A2(n99), .ZN(out[78]) );
  OR2_X1 U330 ( .A1(n100), .A2(key[78]), .ZN(n306) );
  AND2_X1 U331 ( .A1(key[78]), .A2(n100), .ZN(n305) );
  OR2_X1 U332 ( .A1(n307), .A2(n101), .ZN(out[77]) );
  OR2_X1 U333 ( .A1(n102), .A2(key[77]), .ZN(n308) );
  AND2_X1 U334 ( .A1(key[77]), .A2(n102), .ZN(n307) );
  OR2_X1 U335 ( .A1(n309), .A2(n103), .ZN(out[76]) );
  OR2_X1 U336 ( .A1(n104), .A2(key[76]), .ZN(n310) );
  AND2_X1 U337 ( .A1(key[76]), .A2(n104), .ZN(n309) );
  OR2_X1 U338 ( .A1(n311), .A2(n105), .ZN(out[75]) );
  OR2_X1 U339 ( .A1(n106), .A2(key[75]), .ZN(n312) );
  AND2_X1 U340 ( .A1(key[75]), .A2(n106), .ZN(n311) );
  OR2_X1 U341 ( .A1(n313), .A2(n107), .ZN(out[74]) );
  OR2_X1 U342 ( .A1(n108), .A2(key[74]), .ZN(n314) );
  AND2_X1 U343 ( .A1(key[74]), .A2(n108), .ZN(n313) );
  OR2_X1 U344 ( .A1(n315), .A2(n109), .ZN(out[73]) );
  OR2_X1 U345 ( .A1(n110), .A2(key[73]), .ZN(n316) );
  AND2_X1 U346 ( .A1(key[73]), .A2(n110), .ZN(n315) );
  OR2_X1 U347 ( .A1(n317), .A2(n111), .ZN(out[72]) );
  OR2_X1 U348 ( .A1(n112), .A2(key[72]), .ZN(n318) );
  AND2_X1 U349 ( .A1(key[72]), .A2(n112), .ZN(n317) );
  OR2_X1 U350 ( .A1(n319), .A2(n113), .ZN(out[71]) );
  OR2_X1 U351 ( .A1(n114), .A2(key[71]), .ZN(n320) );
  AND2_X1 U352 ( .A1(key[71]), .A2(n114), .ZN(n319) );
  OR2_X1 U353 ( .A1(n321), .A2(n115), .ZN(out[70]) );
  OR2_X1 U354 ( .A1(n116), .A2(key[70]), .ZN(n322) );
  AND2_X1 U355 ( .A1(key[70]), .A2(n116), .ZN(n321) );
  OR2_X1 U356 ( .A1(n323), .A2(n243), .ZN(out[6]) );
  OR2_X1 U357 ( .A1(n244), .A2(key[6]), .ZN(n324) );
  AND2_X1 U358 ( .A1(key[6]), .A2(n244), .ZN(n323) );
  OR2_X1 U359 ( .A1(n325), .A2(n117), .ZN(out[69]) );
  OR2_X1 U360 ( .A1(n118), .A2(key[69]), .ZN(n326) );
  AND2_X1 U361 ( .A1(key[69]), .A2(n118), .ZN(n325) );
  OR2_X1 U362 ( .A1(n327), .A2(n119), .ZN(out[68]) );
  OR2_X1 U363 ( .A1(n120), .A2(key[68]), .ZN(n328) );
  AND2_X1 U364 ( .A1(key[68]), .A2(n120), .ZN(n327) );
  OR2_X1 U365 ( .A1(n329), .A2(n121), .ZN(out[67]) );
  OR2_X1 U366 ( .A1(n122), .A2(key[67]), .ZN(n330) );
  AND2_X1 U367 ( .A1(key[67]), .A2(n122), .ZN(n329) );
  OR2_X1 U368 ( .A1(n331), .A2(n123), .ZN(out[66]) );
  OR2_X1 U369 ( .A1(n124), .A2(key[66]), .ZN(n332) );
  AND2_X1 U370 ( .A1(key[66]), .A2(n124), .ZN(n331) );
  OR2_X1 U371 ( .A1(n333), .A2(n125), .ZN(out[65]) );
  OR2_X1 U372 ( .A1(n126), .A2(key[65]), .ZN(n334) );
  AND2_X1 U373 ( .A1(key[65]), .A2(n126), .ZN(n333) );
  OR2_X1 U374 ( .A1(n335), .A2(n127), .ZN(out[64]) );
  OR2_X1 U375 ( .A1(n128), .A2(key[64]), .ZN(n336) );
  AND2_X1 U376 ( .A1(key[64]), .A2(n128), .ZN(n335) );
  OR2_X1 U377 ( .A1(n337), .A2(n129), .ZN(out[63]) );
  OR2_X1 U378 ( .A1(n130), .A2(key[63]), .ZN(n338) );
  AND2_X1 U379 ( .A1(key[63]), .A2(n130), .ZN(n337) );
  OR2_X1 U380 ( .A1(n339), .A2(n131), .ZN(out[62]) );
  OR2_X1 U381 ( .A1(n132), .A2(key[62]), .ZN(n340) );
  AND2_X1 U382 ( .A1(key[62]), .A2(n132), .ZN(n339) );
  OR2_X1 U383 ( .A1(n341), .A2(n133), .ZN(out[61]) );
  OR2_X1 U384 ( .A1(n134), .A2(key[61]), .ZN(n342) );
  AND2_X1 U385 ( .A1(key[61]), .A2(n134), .ZN(n341) );
  OR2_X1 U386 ( .A1(n343), .A2(n135), .ZN(out[60]) );
  OR2_X1 U387 ( .A1(n136), .A2(key[60]), .ZN(n344) );
  AND2_X1 U388 ( .A1(key[60]), .A2(n136), .ZN(n343) );
  OR2_X1 U389 ( .A1(n345), .A2(n245), .ZN(out[5]) );
  OR2_X1 U390 ( .A1(n246), .A2(key[5]), .ZN(n346) );
  AND2_X1 U391 ( .A1(key[5]), .A2(n246), .ZN(n345) );
  OR2_X1 U392 ( .A1(n347), .A2(n137), .ZN(out[59]) );
  OR2_X1 U393 ( .A1(n138), .A2(key[59]), .ZN(n348) );
  AND2_X1 U394 ( .A1(key[59]), .A2(n138), .ZN(n347) );
  OR2_X1 U395 ( .A1(n349), .A2(n139), .ZN(out[58]) );
  OR2_X1 U396 ( .A1(n140), .A2(key[58]), .ZN(n350) );
  AND2_X1 U397 ( .A1(key[58]), .A2(n140), .ZN(n349) );
  OR2_X1 U398 ( .A1(n351), .A2(n141), .ZN(out[57]) );
  OR2_X1 U399 ( .A1(n142), .A2(key[57]), .ZN(n352) );
  AND2_X1 U400 ( .A1(key[57]), .A2(n142), .ZN(n351) );
  OR2_X1 U401 ( .A1(n353), .A2(n143), .ZN(out[56]) );
  OR2_X1 U402 ( .A1(n144), .A2(key[56]), .ZN(n354) );
  AND2_X1 U403 ( .A1(key[56]), .A2(n144), .ZN(n353) );
  OR2_X1 U404 ( .A1(n355), .A2(n145), .ZN(out[55]) );
  OR2_X1 U405 ( .A1(n146), .A2(key[55]), .ZN(n356) );
  AND2_X1 U406 ( .A1(key[55]), .A2(n146), .ZN(n355) );
  OR2_X1 U407 ( .A1(n357), .A2(n147), .ZN(out[54]) );
  OR2_X1 U408 ( .A1(n148), .A2(key[54]), .ZN(n358) );
  AND2_X1 U409 ( .A1(key[54]), .A2(n148), .ZN(n357) );
  OR2_X1 U410 ( .A1(n359), .A2(n149), .ZN(out[53]) );
  OR2_X1 U411 ( .A1(n150), .A2(key[53]), .ZN(n360) );
  AND2_X1 U412 ( .A1(key[53]), .A2(n150), .ZN(n359) );
  OR2_X1 U413 ( .A1(n361), .A2(n151), .ZN(out[52]) );
  OR2_X1 U414 ( .A1(n152), .A2(key[52]), .ZN(n362) );
  AND2_X1 U415 ( .A1(key[52]), .A2(n152), .ZN(n361) );
  OR2_X1 U416 ( .A1(n363), .A2(n153), .ZN(out[51]) );
  OR2_X1 U417 ( .A1(n154), .A2(key[51]), .ZN(n364) );
  AND2_X1 U418 ( .A1(key[51]), .A2(n154), .ZN(n363) );
  OR2_X1 U419 ( .A1(n365), .A2(n155), .ZN(out[50]) );
  OR2_X1 U420 ( .A1(n156), .A2(key[50]), .ZN(n366) );
  AND2_X1 U421 ( .A1(key[50]), .A2(n156), .ZN(n365) );
  OR2_X1 U422 ( .A1(n367), .A2(n247), .ZN(out[4]) );
  OR2_X1 U423 ( .A1(n248), .A2(key[4]), .ZN(n368) );
  AND2_X1 U424 ( .A1(key[4]), .A2(n248), .ZN(n367) );
  OR2_X1 U425 ( .A1(n369), .A2(n157), .ZN(out[49]) );
  OR2_X1 U426 ( .A1(n158), .A2(key[49]), .ZN(n370) );
  AND2_X1 U427 ( .A1(key[49]), .A2(n158), .ZN(n369) );
  OR2_X1 U428 ( .A1(n371), .A2(n159), .ZN(out[48]) );
  OR2_X1 U429 ( .A1(n160), .A2(key[48]), .ZN(n372) );
  AND2_X1 U430 ( .A1(key[48]), .A2(n160), .ZN(n371) );
  OR2_X1 U431 ( .A1(n373), .A2(n161), .ZN(out[47]) );
  OR2_X1 U432 ( .A1(n162), .A2(key[47]), .ZN(n374) );
  AND2_X1 U433 ( .A1(key[47]), .A2(n162), .ZN(n373) );
  OR2_X1 U434 ( .A1(n375), .A2(n163), .ZN(out[46]) );
  OR2_X1 U435 ( .A1(n164), .A2(key[46]), .ZN(n376) );
  AND2_X1 U436 ( .A1(key[46]), .A2(n164), .ZN(n375) );
  OR2_X1 U437 ( .A1(n377), .A2(n165), .ZN(out[45]) );
  OR2_X1 U438 ( .A1(n166), .A2(key[45]), .ZN(n378) );
  AND2_X1 U439 ( .A1(key[45]), .A2(n166), .ZN(n377) );
  OR2_X1 U440 ( .A1(n379), .A2(n167), .ZN(out[44]) );
  OR2_X1 U441 ( .A1(n168), .A2(key[44]), .ZN(n380) );
  AND2_X1 U442 ( .A1(key[44]), .A2(n168), .ZN(n379) );
  OR2_X1 U443 ( .A1(n381), .A2(n169), .ZN(out[43]) );
  OR2_X1 U444 ( .A1(n170), .A2(key[43]), .ZN(n382) );
  AND2_X1 U445 ( .A1(key[43]), .A2(n170), .ZN(n381) );
  OR2_X1 U446 ( .A1(n383), .A2(n171), .ZN(out[42]) );
  OR2_X1 U447 ( .A1(n172), .A2(key[42]), .ZN(n384) );
  AND2_X1 U448 ( .A1(key[42]), .A2(n172), .ZN(n383) );
  OR2_X1 U449 ( .A1(n385), .A2(n173), .ZN(out[41]) );
  OR2_X1 U450 ( .A1(n174), .A2(key[41]), .ZN(n386) );
  AND2_X1 U451 ( .A1(key[41]), .A2(n174), .ZN(n385) );
  OR2_X1 U452 ( .A1(n387), .A2(n175), .ZN(out[40]) );
  OR2_X1 U453 ( .A1(n176), .A2(key[40]), .ZN(n388) );
  AND2_X1 U454 ( .A1(key[40]), .A2(n176), .ZN(n387) );
  OR2_X1 U455 ( .A1(n389), .A2(n249), .ZN(out[3]) );
  OR2_X1 U456 ( .A1(n250), .A2(key[3]), .ZN(n390) );
  AND2_X1 U457 ( .A1(key[3]), .A2(n250), .ZN(n389) );
  OR2_X1 U458 ( .A1(n391), .A2(n177), .ZN(out[39]) );
  OR2_X1 U459 ( .A1(n178), .A2(key[39]), .ZN(n392) );
  AND2_X1 U460 ( .A1(key[39]), .A2(n178), .ZN(n391) );
  OR2_X1 U461 ( .A1(n393), .A2(n179), .ZN(out[38]) );
  OR2_X1 U462 ( .A1(n180), .A2(key[38]), .ZN(n394) );
  AND2_X1 U463 ( .A1(key[38]), .A2(n180), .ZN(n393) );
  OR2_X1 U464 ( .A1(n395), .A2(n181), .ZN(out[37]) );
  OR2_X1 U465 ( .A1(n182), .A2(key[37]), .ZN(n396) );
  AND2_X1 U466 ( .A1(key[37]), .A2(n182), .ZN(n395) );
  OR2_X1 U467 ( .A1(n397), .A2(n183), .ZN(out[36]) );
  OR2_X1 U468 ( .A1(n184), .A2(key[36]), .ZN(n398) );
  AND2_X1 U469 ( .A1(key[36]), .A2(n184), .ZN(n397) );
  OR2_X1 U470 ( .A1(n399), .A2(n185), .ZN(out[35]) );
  OR2_X1 U471 ( .A1(n186), .A2(key[35]), .ZN(n400) );
  AND2_X1 U472 ( .A1(key[35]), .A2(n186), .ZN(n399) );
  OR2_X1 U473 ( .A1(n401), .A2(n187), .ZN(out[34]) );
  OR2_X1 U474 ( .A1(n188), .A2(key[34]), .ZN(n402) );
  AND2_X1 U475 ( .A1(key[34]), .A2(n188), .ZN(n401) );
  OR2_X1 U476 ( .A1(n403), .A2(n189), .ZN(out[33]) );
  OR2_X1 U477 ( .A1(n190), .A2(key[33]), .ZN(n404) );
  AND2_X1 U478 ( .A1(key[33]), .A2(n190), .ZN(n403) );
  OR2_X1 U479 ( .A1(n405), .A2(n191), .ZN(out[32]) );
  OR2_X1 U480 ( .A1(n192), .A2(key[32]), .ZN(n406) );
  AND2_X1 U481 ( .A1(key[32]), .A2(n192), .ZN(n405) );
  OR2_X1 U482 ( .A1(n407), .A2(n193), .ZN(out[31]) );
  OR2_X1 U483 ( .A1(n194), .A2(key[31]), .ZN(n408) );
  AND2_X1 U484 ( .A1(key[31]), .A2(n194), .ZN(n407) );
  OR2_X1 U485 ( .A1(n409), .A2(n195), .ZN(out[30]) );
  OR2_X1 U486 ( .A1(n196), .A2(key[30]), .ZN(n410) );
  AND2_X1 U487 ( .A1(key[30]), .A2(n196), .ZN(n409) );
  OR2_X1 U488 ( .A1(n411), .A2(n251), .ZN(out[2]) );
  OR2_X1 U489 ( .A1(n252), .A2(key[2]), .ZN(n412) );
  AND2_X1 U490 ( .A1(key[2]), .A2(n252), .ZN(n411) );
  OR2_X1 U491 ( .A1(n413), .A2(n197), .ZN(out[29]) );
  OR2_X1 U492 ( .A1(n198), .A2(key[29]), .ZN(n414) );
  AND2_X1 U493 ( .A1(key[29]), .A2(n198), .ZN(n413) );
  OR2_X1 U494 ( .A1(n415), .A2(n199), .ZN(out[28]) );
  OR2_X1 U495 ( .A1(n200), .A2(key[28]), .ZN(n416) );
  AND2_X1 U496 ( .A1(key[28]), .A2(n200), .ZN(n415) );
  OR2_X1 U497 ( .A1(n417), .A2(n201), .ZN(out[27]) );
  OR2_X1 U498 ( .A1(n202), .A2(key[27]), .ZN(n418) );
  AND2_X1 U499 ( .A1(key[27]), .A2(n202), .ZN(n417) );
  OR2_X1 U500 ( .A1(n419), .A2(n203), .ZN(out[26]) );
  OR2_X1 U501 ( .A1(n204), .A2(key[26]), .ZN(n420) );
  AND2_X1 U502 ( .A1(key[26]), .A2(n204), .ZN(n419) );
  OR2_X1 U503 ( .A1(n421), .A2(n205), .ZN(out[25]) );
  OR2_X1 U504 ( .A1(n206), .A2(key[25]), .ZN(n422) );
  AND2_X1 U505 ( .A1(key[25]), .A2(n206), .ZN(n421) );
  OR2_X1 U506 ( .A1(n423), .A2(n207), .ZN(out[24]) );
  OR2_X1 U507 ( .A1(n208), .A2(key[24]), .ZN(n424) );
  AND2_X1 U508 ( .A1(key[24]), .A2(n208), .ZN(n423) );
  OR2_X1 U509 ( .A1(n425), .A2(n209), .ZN(out[23]) );
  OR2_X1 U510 ( .A1(n210), .A2(key[23]), .ZN(n426) );
  AND2_X1 U511 ( .A1(key[23]), .A2(n210), .ZN(n425) );
  OR2_X1 U512 ( .A1(n427), .A2(n211), .ZN(out[22]) );
  OR2_X1 U513 ( .A1(n212), .A2(key[22]), .ZN(n428) );
  AND2_X1 U514 ( .A1(key[22]), .A2(n212), .ZN(n427) );
  OR2_X1 U515 ( .A1(n429), .A2(n213), .ZN(out[21]) );
  OR2_X1 U516 ( .A1(n214), .A2(key[21]), .ZN(n430) );
  AND2_X1 U517 ( .A1(key[21]), .A2(n214), .ZN(n429) );
  OR2_X1 U518 ( .A1(n431), .A2(n215), .ZN(out[20]) );
  OR2_X1 U519 ( .A1(n216), .A2(key[20]), .ZN(n432) );
  AND2_X1 U520 ( .A1(key[20]), .A2(n216), .ZN(n431) );
  OR2_X1 U521 ( .A1(n433), .A2(n253), .ZN(out[1]) );
  OR2_X1 U522 ( .A1(n254), .A2(key[1]), .ZN(n434) );
  AND2_X1 U523 ( .A1(key[1]), .A2(n254), .ZN(n433) );
  OR2_X1 U524 ( .A1(n435), .A2(n217), .ZN(out[19]) );
  OR2_X1 U525 ( .A1(n218), .A2(key[19]), .ZN(n436) );
  AND2_X1 U526 ( .A1(key[19]), .A2(n218), .ZN(n435) );
  OR2_X1 U527 ( .A1(n437), .A2(n219), .ZN(out[18]) );
  OR2_X1 U528 ( .A1(n220), .A2(key[18]), .ZN(n438) );
  AND2_X1 U529 ( .A1(key[18]), .A2(n220), .ZN(n437) );
  OR2_X1 U530 ( .A1(n439), .A2(n221), .ZN(out[17]) );
  OR2_X1 U531 ( .A1(n222), .A2(key[17]), .ZN(n440) );
  AND2_X1 U532 ( .A1(key[17]), .A2(n222), .ZN(n439) );
  OR2_X1 U533 ( .A1(n441), .A2(n223), .ZN(out[16]) );
  OR2_X1 U534 ( .A1(n224), .A2(key[16]), .ZN(n442) );
  AND2_X1 U535 ( .A1(key[16]), .A2(n224), .ZN(n441) );
  OR2_X1 U536 ( .A1(n443), .A2(n225), .ZN(out[15]) );
  OR2_X1 U537 ( .A1(n226), .A2(key[15]), .ZN(n444) );
  AND2_X1 U538 ( .A1(key[15]), .A2(n226), .ZN(n443) );
  OR2_X1 U539 ( .A1(n445), .A2(n227), .ZN(out[14]) );
  OR2_X1 U540 ( .A1(n228), .A2(key[14]), .ZN(n446) );
  AND2_X1 U541 ( .A1(key[14]), .A2(n228), .ZN(n445) );
  OR2_X1 U542 ( .A1(n447), .A2(n229), .ZN(out[13]) );
  OR2_X1 U543 ( .A1(n230), .A2(key[13]), .ZN(n448) );
  AND2_X1 U544 ( .A1(key[13]), .A2(n230), .ZN(n447) );
  OR2_X1 U545 ( .A1(n449), .A2(n231), .ZN(out[12]) );
  OR2_X1 U546 ( .A1(n232), .A2(key[12]), .ZN(n450) );
  AND2_X1 U547 ( .A1(key[12]), .A2(n232), .ZN(n449) );
  OR2_X1 U548 ( .A1(n451), .A2(n1), .ZN(out[127]) );
  OR2_X1 U549 ( .A1(n2), .A2(key[127]), .ZN(n452) );
  AND2_X1 U550 ( .A1(key[127]), .A2(n2), .ZN(n451) );
  OR2_X1 U551 ( .A1(n453), .A2(n3), .ZN(out[126]) );
  OR2_X1 U552 ( .A1(n4), .A2(key[126]), .ZN(n454) );
  AND2_X1 U553 ( .A1(key[126]), .A2(n4), .ZN(n453) );
  OR2_X1 U554 ( .A1(n455), .A2(n5), .ZN(out[125]) );
  OR2_X1 U555 ( .A1(n6), .A2(key[125]), .ZN(n456) );
  AND2_X1 U556 ( .A1(key[125]), .A2(n6), .ZN(n455) );
  OR2_X1 U557 ( .A1(n457), .A2(n7), .ZN(out[124]) );
  OR2_X1 U558 ( .A1(n8), .A2(key[124]), .ZN(n458) );
  AND2_X1 U559 ( .A1(key[124]), .A2(n8), .ZN(n457) );
  OR2_X1 U560 ( .A1(n459), .A2(n9), .ZN(out[123]) );
  OR2_X1 U561 ( .A1(n10), .A2(key[123]), .ZN(n460) );
  AND2_X1 U562 ( .A1(key[123]), .A2(n10), .ZN(n459) );
  OR2_X1 U563 ( .A1(n461), .A2(n11), .ZN(out[122]) );
  OR2_X1 U564 ( .A1(n12), .A2(key[122]), .ZN(n462) );
  AND2_X1 U565 ( .A1(key[122]), .A2(n12), .ZN(n461) );
  OR2_X1 U566 ( .A1(n463), .A2(n13), .ZN(out[121]) );
  OR2_X1 U567 ( .A1(n14), .A2(key[121]), .ZN(n464) );
  AND2_X1 U568 ( .A1(key[121]), .A2(n14), .ZN(n463) );
  OR2_X1 U569 ( .A1(n465), .A2(n15), .ZN(out[120]) );
  OR2_X1 U570 ( .A1(n16), .A2(key[120]), .ZN(n466) );
  AND2_X1 U571 ( .A1(key[120]), .A2(n16), .ZN(n465) );
  OR2_X1 U572 ( .A1(n467), .A2(n233), .ZN(out[11]) );
  OR2_X1 U573 ( .A1(n234), .A2(key[11]), .ZN(n468) );
  AND2_X1 U574 ( .A1(key[11]), .A2(n234), .ZN(n467) );
  OR2_X1 U575 ( .A1(n469), .A2(n17), .ZN(out[119]) );
  OR2_X1 U576 ( .A1(n18), .A2(key[119]), .ZN(n470) );
  AND2_X1 U577 ( .A1(key[119]), .A2(n18), .ZN(n469) );
  OR2_X1 U578 ( .A1(n471), .A2(n19), .ZN(out[118]) );
  OR2_X1 U579 ( .A1(n20), .A2(key[118]), .ZN(n472) );
  AND2_X1 U580 ( .A1(key[118]), .A2(n20), .ZN(n471) );
  OR2_X1 U581 ( .A1(n473), .A2(n21), .ZN(out[117]) );
  OR2_X1 U582 ( .A1(n22), .A2(key[117]), .ZN(n474) );
  AND2_X1 U583 ( .A1(key[117]), .A2(n22), .ZN(n473) );
  OR2_X1 U584 ( .A1(n475), .A2(n23), .ZN(out[116]) );
  OR2_X1 U585 ( .A1(n24), .A2(key[116]), .ZN(n476) );
  AND2_X1 U586 ( .A1(key[116]), .A2(n24), .ZN(n475) );
  OR2_X1 U587 ( .A1(n477), .A2(n25), .ZN(out[115]) );
  OR2_X1 U588 ( .A1(n26), .A2(key[115]), .ZN(n478) );
  AND2_X1 U589 ( .A1(key[115]), .A2(n26), .ZN(n477) );
  OR2_X1 U590 ( .A1(n479), .A2(n27), .ZN(out[114]) );
  OR2_X1 U591 ( .A1(n28), .A2(key[114]), .ZN(n480) );
  AND2_X1 U592 ( .A1(key[114]), .A2(n28), .ZN(n479) );
  OR2_X1 U593 ( .A1(n481), .A2(n29), .ZN(out[113]) );
  OR2_X1 U594 ( .A1(n30), .A2(key[113]), .ZN(n482) );
  AND2_X1 U595 ( .A1(key[113]), .A2(n30), .ZN(n481) );
  OR2_X1 U596 ( .A1(n483), .A2(n31), .ZN(out[112]) );
  OR2_X1 U597 ( .A1(n32), .A2(key[112]), .ZN(n484) );
  AND2_X1 U598 ( .A1(key[112]), .A2(n32), .ZN(n483) );
  OR2_X1 U599 ( .A1(n485), .A2(n33), .ZN(out[111]) );
  OR2_X1 U600 ( .A1(n34), .A2(key[111]), .ZN(n486) );
  AND2_X1 U601 ( .A1(key[111]), .A2(n34), .ZN(n485) );
  OR2_X1 U602 ( .A1(n487), .A2(n35), .ZN(out[110]) );
  OR2_X1 U603 ( .A1(n36), .A2(key[110]), .ZN(n488) );
  AND2_X1 U604 ( .A1(key[110]), .A2(n36), .ZN(n487) );
  OR2_X1 U605 ( .A1(n489), .A2(n235), .ZN(out[10]) );
  OR2_X1 U606 ( .A1(n236), .A2(key[10]), .ZN(n490) );
  AND2_X1 U607 ( .A1(key[10]), .A2(n236), .ZN(n489) );
  OR2_X1 U608 ( .A1(n491), .A2(n37), .ZN(out[109]) );
  OR2_X1 U609 ( .A1(n38), .A2(key[109]), .ZN(n492) );
  AND2_X1 U610 ( .A1(key[109]), .A2(n38), .ZN(n491) );
  OR2_X1 U611 ( .A1(n493), .A2(n39), .ZN(out[108]) );
  OR2_X1 U612 ( .A1(n40), .A2(key[108]), .ZN(n494) );
  AND2_X1 U613 ( .A1(key[108]), .A2(n40), .ZN(n493) );
  OR2_X1 U614 ( .A1(n495), .A2(n41), .ZN(out[107]) );
  OR2_X1 U615 ( .A1(n42), .A2(key[107]), .ZN(n496) );
  AND2_X1 U616 ( .A1(key[107]), .A2(n42), .ZN(n495) );
  OR2_X1 U617 ( .A1(n497), .A2(n43), .ZN(out[106]) );
  OR2_X1 U618 ( .A1(n44), .A2(key[106]), .ZN(n498) );
  AND2_X1 U619 ( .A1(key[106]), .A2(n44), .ZN(n497) );
  OR2_X1 U620 ( .A1(n499), .A2(n45), .ZN(out[105]) );
  OR2_X1 U621 ( .A1(n46), .A2(key[105]), .ZN(n500) );
  AND2_X1 U622 ( .A1(key[105]), .A2(n46), .ZN(n499) );
  OR2_X1 U623 ( .A1(n501), .A2(n47), .ZN(out[104]) );
  OR2_X1 U624 ( .A1(n48), .A2(key[104]), .ZN(n502) );
  AND2_X1 U625 ( .A1(key[104]), .A2(n48), .ZN(n501) );
  OR2_X1 U626 ( .A1(n503), .A2(n49), .ZN(out[103]) );
  OR2_X1 U627 ( .A1(n50), .A2(key[103]), .ZN(n504) );
  AND2_X1 U628 ( .A1(key[103]), .A2(n50), .ZN(n503) );
  OR2_X1 U629 ( .A1(n505), .A2(n51), .ZN(out[102]) );
  OR2_X1 U630 ( .A1(n52), .A2(key[102]), .ZN(n506) );
  AND2_X1 U631 ( .A1(key[102]), .A2(n52), .ZN(n505) );
  OR2_X1 U632 ( .A1(n507), .A2(n53), .ZN(out[101]) );
  OR2_X1 U633 ( .A1(n54), .A2(key[101]), .ZN(n508) );
  AND2_X1 U634 ( .A1(key[101]), .A2(n54), .ZN(n507) );
  OR2_X1 U635 ( .A1(n509), .A2(n55), .ZN(out[100]) );
  OR2_X1 U636 ( .A1(n56), .A2(key[100]), .ZN(n510) );
  AND2_X1 U637 ( .A1(key[100]), .A2(n56), .ZN(n509) );
  OR2_X1 U638 ( .A1(n511), .A2(n255), .ZN(out[0]) );
  OR2_X1 U639 ( .A1(n256), .A2(key[0]), .ZN(n512) );
  AND2_X1 U640 ( .A1(key[0]), .A2(n256), .ZN(n511) );
endmodule


module CD2_17 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_18 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done

  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_19 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done

  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_20 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD4_9 ( a, b, y );
  input [3:0] a;
  input [3:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  //input_done

  output [15:0] y;
  reg [15:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]);
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]);
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]);
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]);
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]);
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]);
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]);
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]);
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]);
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]);
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]);
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]);
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]);
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]);
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]);
endmodule




module CD4_10 ( a, b, y );
  input [3:0] a;
  input [3:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  //input_done

  output [15:0] y;
  reg [15:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]);
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]);
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]);
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]);
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]);
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]);
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]);
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]);
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]);
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]);
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]);
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]);
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]);
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]);
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]);
endmodule




module CD16_5 ( a, b, y );
  input [15:0] a;
  input [15:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign abar[8] = ~a[8];
  assign abar[9] = ~a[9];
  assign abar[10] = ~a[10];
  assign abar[11] = ~a[11];
  assign abar[12] = ~a[12];
  assign abar[13] = ~a[13];
  assign abar[14] = ~a[14];
  assign abar[15] = ~a[15];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign bbar[8] = ~b[8];
  assign bbar[9] = ~b[9];
  assign bbar[10] = ~b[10];
  assign bbar[11] = ~b[11];
  assign bbar[12] = ~b[12];
  assign bbar[13] = ~b[13];
  assign bbar[14] = ~b[14];
  assign bbar[15] = ~b[15];
  //input_done

  output [255:0] y;
  reg [255:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[9]), .A2(a[0]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[9]), .A2(abar[0]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[3]), .A2(a[6]), .ZN(y[99]) );
  OR2_X1 U2bar ( .A1(bbar[3]), .A2(abar[6]), .ZN(ybar[99]);
  AND2_X1 U3 ( .A1(b[2]), .A2(a[6]), .ZN(y[98]) );
  OR2_X1 U3bar ( .A1(bbar[2]), .A2(abar[6]), .ZN(ybar[98]);
  AND2_X1 U4 ( .A1(b[1]), .A2(a[6]), .ZN(y[97]) );
  OR2_X1 U4bar ( .A1(bbar[1]), .A2(abar[6]), .ZN(ybar[97]);
  AND2_X1 U5 ( .A1(b[0]), .A2(a[6]), .ZN(y[96]) );
  OR2_X1 U5bar ( .A1(bbar[0]), .A2(abar[6]), .ZN(ybar[96]);
  AND2_X1 U6 ( .A1(b[15]), .A2(a[5]), .ZN(y[95]) );
  OR2_X1 U6bar ( .A1(bbar[15]), .A2(abar[5]), .ZN(ybar[95]);
  AND2_X1 U7 ( .A1(b[14]), .A2(a[5]), .ZN(y[94]) );
  OR2_X1 U7bar ( .A1(bbar[14]), .A2(abar[5]), .ZN(ybar[94]);
  AND2_X1 U8 ( .A1(b[13]), .A2(a[5]), .ZN(y[93]) );
  OR2_X1 U8bar ( .A1(bbar[13]), .A2(abar[5]), .ZN(ybar[93]);
  AND2_X1 U9 ( .A1(b[12]), .A2(a[5]), .ZN(y[92]) );
  OR2_X1 U9bar ( .A1(bbar[12]), .A2(abar[5]), .ZN(ybar[92]);
  AND2_X1 U10 ( .A1(b[11]), .A2(a[5]), .ZN(y[91]) );
  OR2_X1 U10bar ( .A1(bbar[11]), .A2(abar[5]), .ZN(ybar[91]);
  AND2_X1 U11 ( .A1(b[10]), .A2(a[5]), .ZN(y[90]) );
  OR2_X1 U11bar ( .A1(bbar[10]), .A2(abar[5]), .ZN(ybar[90]);
  AND2_X1 U12 ( .A1(b[8]), .A2(a[0]), .ZN(y[8]) );
  OR2_X1 U12bar ( .A1(bbar[8]), .A2(abar[0]), .ZN(ybar[8]);
  AND2_X1 U13 ( .A1(a[5]), .A2(b[9]), .ZN(y[89]) );
  OR2_X1 U13bar ( .A1(abar[5]), .A2(bbar[9]), .ZN(ybar[89]);
  AND2_X1 U14 ( .A1(b[8]), .A2(a[5]), .ZN(y[88]) );
  OR2_X1 U14bar ( .A1(bbar[8]), .A2(abar[5]), .ZN(ybar[88]);
  AND2_X1 U15 ( .A1(b[7]), .A2(a[5]), .ZN(y[87]) );
  OR2_X1 U15bar ( .A1(bbar[7]), .A2(abar[5]), .ZN(ybar[87]);
  AND2_X1 U16 ( .A1(b[6]), .A2(a[5]), .ZN(y[86]) );
  OR2_X1 U16bar ( .A1(bbar[6]), .A2(abar[5]), .ZN(ybar[86]);
  AND2_X1 U17 ( .A1(b[5]), .A2(a[5]), .ZN(y[85]) );
  OR2_X1 U17bar ( .A1(bbar[5]), .A2(abar[5]), .ZN(ybar[85]);
  AND2_X1 U18 ( .A1(b[4]), .A2(a[5]), .ZN(y[84]) );
  OR2_X1 U18bar ( .A1(bbar[4]), .A2(abar[5]), .ZN(ybar[84]);
  AND2_X1 U19 ( .A1(a[5]), .A2(b[3]), .ZN(y[83]) );
  OR2_X1 U19bar ( .A1(abar[5]), .A2(bbar[3]), .ZN(ybar[83]);
  AND2_X1 U20 ( .A1(a[5]), .A2(b[2]), .ZN(y[82]) );
  OR2_X1 U20bar ( .A1(abar[5]), .A2(bbar[2]), .ZN(ybar[82]);
  AND2_X1 U21 ( .A1(a[5]), .A2(b[1]), .ZN(y[81]) );
  OR2_X1 U21bar ( .A1(abar[5]), .A2(bbar[1]), .ZN(ybar[81]);
  AND2_X1 U22 ( .A1(a[5]), .A2(b[0]), .ZN(y[80]) );
  OR2_X1 U22bar ( .A1(abar[5]), .A2(bbar[0]), .ZN(ybar[80]);
  AND2_X1 U23 ( .A1(b[7]), .A2(a[0]), .ZN(y[7]) );
  OR2_X1 U23bar ( .A1(bbar[7]), .A2(abar[0]), .ZN(ybar[7]);
  AND2_X1 U24 ( .A1(a[4]), .A2(b[15]), .ZN(y[79]) );
  OR2_X1 U24bar ( .A1(abar[4]), .A2(bbar[15]), .ZN(ybar[79]);
  AND2_X1 U25 ( .A1(a[4]), .A2(b[14]), .ZN(y[78]) );
  OR2_X1 U25bar ( .A1(abar[4]), .A2(bbar[14]), .ZN(ybar[78]);
  AND2_X1 U26 ( .A1(a[4]), .A2(b[13]), .ZN(y[77]) );
  OR2_X1 U26bar ( .A1(abar[4]), .A2(bbar[13]), .ZN(ybar[77]);
  AND2_X1 U27 ( .A1(a[4]), .A2(b[12]), .ZN(y[76]) );
  OR2_X1 U27bar ( .A1(abar[4]), .A2(bbar[12]), .ZN(ybar[76]);
  AND2_X1 U28 ( .A1(a[4]), .A2(b[11]), .ZN(y[75]) );
  OR2_X1 U28bar ( .A1(abar[4]), .A2(bbar[11]), .ZN(ybar[75]);
  AND2_X1 U29 ( .A1(a[4]), .A2(b[10]), .ZN(y[74]) );
  OR2_X1 U29bar ( .A1(abar[4]), .A2(bbar[10]), .ZN(ybar[74]);
  AND2_X1 U30 ( .A1(a[4]), .A2(b[9]), .ZN(y[73]) );
  OR2_X1 U30bar ( .A1(abar[4]), .A2(bbar[9]), .ZN(ybar[73]);
  AND2_X1 U31 ( .A1(a[4]), .A2(b[8]), .ZN(y[72]) );
  OR2_X1 U31bar ( .A1(abar[4]), .A2(bbar[8]), .ZN(ybar[72]);
  AND2_X1 U32 ( .A1(a[4]), .A2(b[7]), .ZN(y[71]) );
  OR2_X1 U32bar ( .A1(abar[4]), .A2(bbar[7]), .ZN(ybar[71]);
  AND2_X1 U33 ( .A1(a[4]), .A2(b[6]), .ZN(y[70]) );
  OR2_X1 U33bar ( .A1(abar[4]), .A2(bbar[6]), .ZN(ybar[70]);
  AND2_X1 U34 ( .A1(b[6]), .A2(a[0]), .ZN(y[6]) );
  OR2_X1 U34bar ( .A1(bbar[6]), .A2(abar[0]), .ZN(ybar[6]);
  AND2_X1 U35 ( .A1(a[4]), .A2(b[5]), .ZN(y[69]) );
  OR2_X1 U35bar ( .A1(abar[4]), .A2(bbar[5]), .ZN(ybar[69]);
  AND2_X1 U36 ( .A1(a[4]), .A2(b[4]), .ZN(y[68]) );
  OR2_X1 U36bar ( .A1(abar[4]), .A2(bbar[4]), .ZN(ybar[68]);
  AND2_X1 U37 ( .A1(a[4]), .A2(b[3]), .ZN(y[67]) );
  OR2_X1 U37bar ( .A1(abar[4]), .A2(bbar[3]), .ZN(ybar[67]);
  AND2_X1 U38 ( .A1(a[4]), .A2(b[2]), .ZN(y[66]) );
  OR2_X1 U38bar ( .A1(abar[4]), .A2(bbar[2]), .ZN(ybar[66]);
  AND2_X1 U39 ( .A1(a[4]), .A2(b[1]), .ZN(y[65]) );
  OR2_X1 U39bar ( .A1(abar[4]), .A2(bbar[1]), .ZN(ybar[65]);
  AND2_X1 U40 ( .A1(a[4]), .A2(b[0]), .ZN(y[64]) );
  OR2_X1 U40bar ( .A1(abar[4]), .A2(bbar[0]), .ZN(ybar[64]);
  AND2_X1 U41 ( .A1(a[3]), .A2(b[15]), .ZN(y[63]) );
  OR2_X1 U41bar ( .A1(abar[3]), .A2(bbar[15]), .ZN(ybar[63]);
  AND2_X1 U42 ( .A1(a[3]), .A2(b[14]), .ZN(y[62]) );
  OR2_X1 U42bar ( .A1(abar[3]), .A2(bbar[14]), .ZN(ybar[62]);
  AND2_X1 U43 ( .A1(a[3]), .A2(b[13]), .ZN(y[61]) );
  OR2_X1 U43bar ( .A1(abar[3]), .A2(bbar[13]), .ZN(ybar[61]);
  AND2_X1 U44 ( .A1(a[3]), .A2(b[12]), .ZN(y[60]) );
  OR2_X1 U44bar ( .A1(abar[3]), .A2(bbar[12]), .ZN(ybar[60]);
  AND2_X1 U45 ( .A1(b[5]), .A2(a[0]), .ZN(y[5]) );
  OR2_X1 U45bar ( .A1(bbar[5]), .A2(abar[0]), .ZN(ybar[5]);
  AND2_X1 U46 ( .A1(a[3]), .A2(b[11]), .ZN(y[59]) );
  OR2_X1 U46bar ( .A1(abar[3]), .A2(bbar[11]), .ZN(ybar[59]);
  AND2_X1 U47 ( .A1(a[3]), .A2(b[10]), .ZN(y[58]) );
  OR2_X1 U47bar ( .A1(abar[3]), .A2(bbar[10]), .ZN(ybar[58]);
  AND2_X1 U48 ( .A1(a[3]), .A2(b[9]), .ZN(y[57]) );
  OR2_X1 U48bar ( .A1(abar[3]), .A2(bbar[9]), .ZN(ybar[57]);
  AND2_X1 U49 ( .A1(a[3]), .A2(b[8]), .ZN(y[56]) );
  OR2_X1 U49bar ( .A1(abar[3]), .A2(bbar[8]), .ZN(ybar[56]);
  AND2_X1 U50 ( .A1(a[3]), .A2(b[7]), .ZN(y[55]) );
  OR2_X1 U50bar ( .A1(abar[3]), .A2(bbar[7]), .ZN(ybar[55]);
  AND2_X1 U51 ( .A1(a[3]), .A2(b[6]), .ZN(y[54]) );
  OR2_X1 U51bar ( .A1(abar[3]), .A2(bbar[6]), .ZN(ybar[54]);
  AND2_X1 U52 ( .A1(a[3]), .A2(b[5]), .ZN(y[53]) );
  OR2_X1 U52bar ( .A1(abar[3]), .A2(bbar[5]), .ZN(ybar[53]);
  AND2_X1 U53 ( .A1(a[3]), .A2(b[4]), .ZN(y[52]) );
  OR2_X1 U53bar ( .A1(abar[3]), .A2(bbar[4]), .ZN(ybar[52]);
  AND2_X1 U54 ( .A1(a[3]), .A2(b[3]), .ZN(y[51]) );
  OR2_X1 U54bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[51]);
  AND2_X1 U55 ( .A1(a[3]), .A2(b[2]), .ZN(y[50]) );
  OR2_X1 U55bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[50]);
  AND2_X1 U56 ( .A1(b[4]), .A2(a[0]), .ZN(y[4]) );
  OR2_X1 U56bar ( .A1(bbar[4]), .A2(abar[0]), .ZN(ybar[4]);
  AND2_X1 U57 ( .A1(a[3]), .A2(b[1]), .ZN(y[49]) );
  OR2_X1 U57bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[49]);
  AND2_X1 U58 ( .A1(a[3]), .A2(b[0]), .ZN(y[48]) );
  OR2_X1 U58bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[48]);
  AND2_X1 U59 ( .A1(a[2]), .A2(b[15]), .ZN(y[47]) );
  OR2_X1 U59bar ( .A1(abar[2]), .A2(bbar[15]), .ZN(ybar[47]);
  AND2_X1 U60 ( .A1(a[2]), .A2(b[14]), .ZN(y[46]) );
  OR2_X1 U60bar ( .A1(abar[2]), .A2(bbar[14]), .ZN(ybar[46]);
  AND2_X1 U61 ( .A1(a[2]), .A2(b[13]), .ZN(y[45]) );
  OR2_X1 U61bar ( .A1(abar[2]), .A2(bbar[13]), .ZN(ybar[45]);
  AND2_X1 U62 ( .A1(a[2]), .A2(b[12]), .ZN(y[44]) );
  OR2_X1 U62bar ( .A1(abar[2]), .A2(bbar[12]), .ZN(ybar[44]);
  AND2_X1 U63 ( .A1(a[2]), .A2(b[11]), .ZN(y[43]) );
  OR2_X1 U63bar ( .A1(abar[2]), .A2(bbar[11]), .ZN(ybar[43]);
  AND2_X1 U64 ( .A1(a[2]), .A2(b[10]), .ZN(y[42]) );
  OR2_X1 U64bar ( .A1(abar[2]), .A2(bbar[10]), .ZN(ybar[42]);
  AND2_X1 U65 ( .A1(a[2]), .A2(b[9]), .ZN(y[41]) );
  OR2_X1 U65bar ( .A1(abar[2]), .A2(bbar[9]), .ZN(ybar[41]);
  AND2_X1 U66 ( .A1(a[2]), .A2(b[8]), .ZN(y[40]) );
  OR2_X1 U66bar ( .A1(abar[2]), .A2(bbar[8]), .ZN(ybar[40]);
  AND2_X1 U67 ( .A1(b[3]), .A2(a[0]), .ZN(y[3]) );
  OR2_X1 U67bar ( .A1(bbar[3]), .A2(abar[0]), .ZN(ybar[3]);
  AND2_X1 U68 ( .A1(a[2]), .A2(b[7]), .ZN(y[39]) );
  OR2_X1 U68bar ( .A1(abar[2]), .A2(bbar[7]), .ZN(ybar[39]);
  AND2_X1 U69 ( .A1(a[2]), .A2(b[6]), .ZN(y[38]) );
  OR2_X1 U69bar ( .A1(abar[2]), .A2(bbar[6]), .ZN(ybar[38]);
  AND2_X1 U70 ( .A1(a[2]), .A2(b[5]), .ZN(y[37]) );
  OR2_X1 U70bar ( .A1(abar[2]), .A2(bbar[5]), .ZN(ybar[37]);
  AND2_X1 U71 ( .A1(a[2]), .A2(b[4]), .ZN(y[36]) );
  OR2_X1 U71bar ( .A1(abar[2]), .A2(bbar[4]), .ZN(ybar[36]);
  AND2_X1 U72 ( .A1(a[2]), .A2(b[3]), .ZN(y[35]) );
  OR2_X1 U72bar ( .A1(abar[2]), .A2(bbar[3]), .ZN(ybar[35]);
  AND2_X1 U73 ( .A1(a[2]), .A2(b[2]), .ZN(y[34]) );
  OR2_X1 U73bar ( .A1(abar[2]), .A2(bbar[2]), .ZN(ybar[34]);
  AND2_X1 U74 ( .A1(a[2]), .A2(b[1]), .ZN(y[33]) );
  OR2_X1 U74bar ( .A1(abar[2]), .A2(bbar[1]), .ZN(ybar[33]);
  AND2_X1 U75 ( .A1(a[2]), .A2(b[0]), .ZN(y[32]) );
  OR2_X1 U75bar ( .A1(abar[2]), .A2(bbar[0]), .ZN(ybar[32]);
  AND2_X1 U76 ( .A1(a[1]), .A2(b[15]), .ZN(y[31]) );
  OR2_X1 U76bar ( .A1(abar[1]), .A2(bbar[15]), .ZN(ybar[31]);
  AND2_X1 U77 ( .A1(a[1]), .A2(b[14]), .ZN(y[30]) );
  OR2_X1 U77bar ( .A1(abar[1]), .A2(bbar[14]), .ZN(ybar[30]);
  AND2_X1 U78 ( .A1(b[2]), .A2(a[0]), .ZN(y[2]) );
  OR2_X1 U78bar ( .A1(bbar[2]), .A2(abar[0]), .ZN(ybar[2]);
  AND2_X1 U79 ( .A1(a[1]), .A2(b[13]), .ZN(y[29]) );
  OR2_X1 U79bar ( .A1(abar[1]), .A2(bbar[13]), .ZN(ybar[29]);
  AND2_X1 U80 ( .A1(a[1]), .A2(b[12]), .ZN(y[28]) );
  OR2_X1 U80bar ( .A1(abar[1]), .A2(bbar[12]), .ZN(ybar[28]);
  AND2_X1 U81 ( .A1(a[1]), .A2(b[11]), .ZN(y[27]) );
  OR2_X1 U81bar ( .A1(abar[1]), .A2(bbar[11]), .ZN(ybar[27]);
  AND2_X1 U82 ( .A1(a[1]), .A2(b[10]), .ZN(y[26]) );
  OR2_X1 U82bar ( .A1(abar[1]), .A2(bbar[10]), .ZN(ybar[26]);
  AND2_X1 U83 ( .A1(a[1]), .A2(b[9]), .ZN(y[25]) );
  OR2_X1 U83bar ( .A1(abar[1]), .A2(bbar[9]), .ZN(ybar[25]);
  AND2_X1 U84 ( .A1(a[15]), .A2(b[15]), .ZN(y[255]) );
  OR2_X1 U84bar ( .A1(abar[15]), .A2(bbar[15]), .ZN(ybar[255]);
  AND2_X1 U85 ( .A1(a[15]), .A2(b[14]), .ZN(y[254]) );
  OR2_X1 U85bar ( .A1(abar[15]), .A2(bbar[14]), .ZN(ybar[254]);
  AND2_X1 U86 ( .A1(a[15]), .A2(b[13]), .ZN(y[253]) );
  OR2_X1 U86bar ( .A1(abar[15]), .A2(bbar[13]), .ZN(ybar[253]);
  AND2_X1 U87 ( .A1(a[15]), .A2(b[12]), .ZN(y[252]) );
  OR2_X1 U87bar ( .A1(abar[15]), .A2(bbar[12]), .ZN(ybar[252]);
  AND2_X1 U88 ( .A1(a[15]), .A2(b[11]), .ZN(y[251]) );
  OR2_X1 U88bar ( .A1(abar[15]), .A2(bbar[11]), .ZN(ybar[251]);
  AND2_X1 U89 ( .A1(a[15]), .A2(b[10]), .ZN(y[250]) );
  OR2_X1 U89bar ( .A1(abar[15]), .A2(bbar[10]), .ZN(ybar[250]);
  AND2_X1 U90 ( .A1(a[1]), .A2(b[8]), .ZN(y[24]) );
  OR2_X1 U90bar ( .A1(abar[1]), .A2(bbar[8]), .ZN(ybar[24]);
  AND2_X1 U91 ( .A1(a[15]), .A2(b[9]), .ZN(y[249]) );
  OR2_X1 U91bar ( .A1(abar[15]), .A2(bbar[9]), .ZN(ybar[249]);
  AND2_X1 U92 ( .A1(a[15]), .A2(b[8]), .ZN(y[248]) );
  OR2_X1 U92bar ( .A1(abar[15]), .A2(bbar[8]), .ZN(ybar[248]);
  AND2_X1 U93 ( .A1(a[15]), .A2(b[7]), .ZN(y[247]) );
  OR2_X1 U93bar ( .A1(abar[15]), .A2(bbar[7]), .ZN(ybar[247]);
  AND2_X1 U94 ( .A1(a[15]), .A2(b[6]), .ZN(y[246]) );
  OR2_X1 U94bar ( .A1(abar[15]), .A2(bbar[6]), .ZN(ybar[246]);
  AND2_X1 U95 ( .A1(a[15]), .A2(b[5]), .ZN(y[245]) );
  OR2_X1 U95bar ( .A1(abar[15]), .A2(bbar[5]), .ZN(ybar[245]);
  AND2_X1 U96 ( .A1(a[15]), .A2(b[4]), .ZN(y[244]) );
  OR2_X1 U96bar ( .A1(abar[15]), .A2(bbar[4]), .ZN(ybar[244]);
  AND2_X1 U97 ( .A1(a[15]), .A2(b[3]), .ZN(y[243]) );
  OR2_X1 U97bar ( .A1(abar[15]), .A2(bbar[3]), .ZN(ybar[243]);
  AND2_X1 U98 ( .A1(a[15]), .A2(b[2]), .ZN(y[242]) );
  OR2_X1 U98bar ( .A1(abar[15]), .A2(bbar[2]), .ZN(ybar[242]);
  AND2_X1 U99 ( .A1(a[15]), .A2(b[1]), .ZN(y[241]) );
  OR2_X1 U99bar ( .A1(abar[15]), .A2(bbar[1]), .ZN(ybar[241]);
  AND2_X1 U100 ( .A1(a[15]), .A2(b[0]), .ZN(y[240]) );
  OR2_X1 U100bar ( .A1(abar[15]), .A2(bbar[0]), .ZN(ybar[240]);
  AND2_X1 U101 ( .A1(a[1]), .A2(b[7]), .ZN(y[23]) );
  OR2_X1 U101bar ( .A1(abar[1]), .A2(bbar[7]), .ZN(ybar[23]);
  AND2_X1 U102 ( .A1(a[14]), .A2(b[15]), .ZN(y[239]) );
  OR2_X1 U102bar ( .A1(abar[14]), .A2(bbar[15]), .ZN(ybar[239]);
  AND2_X1 U103 ( .A1(a[14]), .A2(b[14]), .ZN(y[238]) );
  OR2_X1 U103bar ( .A1(abar[14]), .A2(bbar[14]), .ZN(ybar[238]);
  AND2_X1 U104 ( .A1(a[14]), .A2(b[13]), .ZN(y[237]) );
  OR2_X1 U104bar ( .A1(abar[14]), .A2(bbar[13]), .ZN(ybar[237]);
  AND2_X1 U105 ( .A1(a[14]), .A2(b[12]), .ZN(y[236]) );
  OR2_X1 U105bar ( .A1(abar[14]), .A2(bbar[12]), .ZN(ybar[236]);
  AND2_X1 U106 ( .A1(a[14]), .A2(b[11]), .ZN(y[235]) );
  OR2_X1 U106bar ( .A1(abar[14]), .A2(bbar[11]), .ZN(ybar[235]);
  AND2_X1 U107 ( .A1(a[14]), .A2(b[10]), .ZN(y[234]) );
  OR2_X1 U107bar ( .A1(abar[14]), .A2(bbar[10]), .ZN(ybar[234]);
  AND2_X1 U108 ( .A1(a[14]), .A2(b[9]), .ZN(y[233]) );
  OR2_X1 U108bar ( .A1(abar[14]), .A2(bbar[9]), .ZN(ybar[233]);
  AND2_X1 U109 ( .A1(a[14]), .A2(b[8]), .ZN(y[232]) );
  OR2_X1 U109bar ( .A1(abar[14]), .A2(bbar[8]), .ZN(ybar[232]);
  AND2_X1 U110 ( .A1(a[14]), .A2(b[7]), .ZN(y[231]) );
  OR2_X1 U110bar ( .A1(abar[14]), .A2(bbar[7]), .ZN(ybar[231]);
  AND2_X1 U111 ( .A1(a[14]), .A2(b[6]), .ZN(y[230]) );
  OR2_X1 U111bar ( .A1(abar[14]), .A2(bbar[6]), .ZN(ybar[230]);
  AND2_X1 U112 ( .A1(a[1]), .A2(b[6]), .ZN(y[22]) );
  OR2_X1 U112bar ( .A1(abar[1]), .A2(bbar[6]), .ZN(ybar[22]);
  AND2_X1 U113 ( .A1(a[14]), .A2(b[5]), .ZN(y[229]) );
  OR2_X1 U113bar ( .A1(abar[14]), .A2(bbar[5]), .ZN(ybar[229]);
  AND2_X1 U114 ( .A1(a[14]), .A2(b[4]), .ZN(y[228]) );
  OR2_X1 U114bar ( .A1(abar[14]), .A2(bbar[4]), .ZN(ybar[228]);
  AND2_X1 U115 ( .A1(a[14]), .A2(b[3]), .ZN(y[227]) );
  OR2_X1 U115bar ( .A1(abar[14]), .A2(bbar[3]), .ZN(ybar[227]);
  AND2_X1 U116 ( .A1(a[14]), .A2(b[2]), .ZN(y[226]) );
  OR2_X1 U116bar ( .A1(abar[14]), .A2(bbar[2]), .ZN(ybar[226]);
  AND2_X1 U117 ( .A1(a[14]), .A2(b[1]), .ZN(y[225]) );
  OR2_X1 U117bar ( .A1(abar[14]), .A2(bbar[1]), .ZN(ybar[225]);
  AND2_X1 U118 ( .A1(a[14]), .A2(b[0]), .ZN(y[224]) );
  OR2_X1 U118bar ( .A1(abar[14]), .A2(bbar[0]), .ZN(ybar[224]);
  AND2_X1 U119 ( .A1(a[13]), .A2(b[15]), .ZN(y[223]) );
  OR2_X1 U119bar ( .A1(abar[13]), .A2(bbar[15]), .ZN(ybar[223]);
  AND2_X1 U120 ( .A1(a[13]), .A2(b[14]), .ZN(y[222]) );
  OR2_X1 U120bar ( .A1(abar[13]), .A2(bbar[14]), .ZN(ybar[222]);
  AND2_X1 U121 ( .A1(a[13]), .A2(b[13]), .ZN(y[221]) );
  OR2_X1 U121bar ( .A1(abar[13]), .A2(bbar[13]), .ZN(ybar[221]);
  AND2_X1 U122 ( .A1(a[13]), .A2(b[12]), .ZN(y[220]) );
  OR2_X1 U122bar ( .A1(abar[13]), .A2(bbar[12]), .ZN(ybar[220]);
  AND2_X1 U123 ( .A1(a[1]), .A2(b[5]), .ZN(y[21]) );
  OR2_X1 U123bar ( .A1(abar[1]), .A2(bbar[5]), .ZN(ybar[21]);
  AND2_X1 U124 ( .A1(a[13]), .A2(b[11]), .ZN(y[219]) );
  OR2_X1 U124bar ( .A1(abar[13]), .A2(bbar[11]), .ZN(ybar[219]);
  AND2_X1 U125 ( .A1(a[13]), .A2(b[10]), .ZN(y[218]) );
  OR2_X1 U125bar ( .A1(abar[13]), .A2(bbar[10]), .ZN(ybar[218]);
  AND2_X1 U126 ( .A1(a[13]), .A2(b[9]), .ZN(y[217]) );
  OR2_X1 U126bar ( .A1(abar[13]), .A2(bbar[9]), .ZN(ybar[217]);
  AND2_X1 U127 ( .A1(a[13]), .A2(b[8]), .ZN(y[216]) );
  OR2_X1 U127bar ( .A1(abar[13]), .A2(bbar[8]), .ZN(ybar[216]);
  AND2_X1 U128 ( .A1(a[13]), .A2(b[7]), .ZN(y[215]) );
  OR2_X1 U128bar ( .A1(abar[13]), .A2(bbar[7]), .ZN(ybar[215]);
  AND2_X1 U129 ( .A1(a[13]), .A2(b[6]), .ZN(y[214]) );
  OR2_X1 U129bar ( .A1(abar[13]), .A2(bbar[6]), .ZN(ybar[214]);
  AND2_X1 U130 ( .A1(a[13]), .A2(b[5]), .ZN(y[213]) );
  OR2_X1 U130bar ( .A1(abar[13]), .A2(bbar[5]), .ZN(ybar[213]);
  AND2_X1 U131 ( .A1(a[13]), .A2(b[4]), .ZN(y[212]) );
  OR2_X1 U131bar ( .A1(abar[13]), .A2(bbar[4]), .ZN(ybar[212]);
  AND2_X1 U132 ( .A1(a[13]), .A2(b[3]), .ZN(y[211]) );
  OR2_X1 U132bar ( .A1(abar[13]), .A2(bbar[3]), .ZN(ybar[211]);
  AND2_X1 U133 ( .A1(a[13]), .A2(b[2]), .ZN(y[210]) );
  OR2_X1 U133bar ( .A1(abar[13]), .A2(bbar[2]), .ZN(ybar[210]);
  AND2_X1 U134 ( .A1(a[1]), .A2(b[4]), .ZN(y[20]) );
  OR2_X1 U134bar ( .A1(abar[1]), .A2(bbar[4]), .ZN(ybar[20]);
  AND2_X1 U135 ( .A1(a[13]), .A2(b[1]), .ZN(y[209]) );
  OR2_X1 U135bar ( .A1(abar[13]), .A2(bbar[1]), .ZN(ybar[209]);
  AND2_X1 U136 ( .A1(a[13]), .A2(b[0]), .ZN(y[208]) );
  OR2_X1 U136bar ( .A1(abar[13]), .A2(bbar[0]), .ZN(ybar[208]);
  AND2_X1 U137 ( .A1(a[12]), .A2(b[15]), .ZN(y[207]) );
  OR2_X1 U137bar ( .A1(abar[12]), .A2(bbar[15]), .ZN(ybar[207]);
  AND2_X1 U138 ( .A1(a[12]), .A2(b[14]), .ZN(y[206]) );
  OR2_X1 U138bar ( .A1(abar[12]), .A2(bbar[14]), .ZN(ybar[206]);
  AND2_X1 U139 ( .A1(a[12]), .A2(b[13]), .ZN(y[205]) );
  OR2_X1 U139bar ( .A1(abar[12]), .A2(bbar[13]), .ZN(ybar[205]);
  AND2_X1 U140 ( .A1(a[12]), .A2(b[12]), .ZN(y[204]) );
  OR2_X1 U140bar ( .A1(abar[12]), .A2(bbar[12]), .ZN(ybar[204]);
  AND2_X1 U141 ( .A1(a[12]), .A2(b[11]), .ZN(y[203]) );
  OR2_X1 U141bar ( .A1(abar[12]), .A2(bbar[11]), .ZN(ybar[203]);
  AND2_X1 U142 ( .A1(a[12]), .A2(b[10]), .ZN(y[202]) );
  OR2_X1 U142bar ( .A1(abar[12]), .A2(bbar[10]), .ZN(ybar[202]);
  AND2_X1 U143 ( .A1(a[12]), .A2(b[9]), .ZN(y[201]) );
  OR2_X1 U143bar ( .A1(abar[12]), .A2(bbar[9]), .ZN(ybar[201]);
  AND2_X1 U144 ( .A1(a[12]), .A2(b[8]), .ZN(y[200]) );
  OR2_X1 U144bar ( .A1(abar[12]), .A2(bbar[8]), .ZN(ybar[200]);
  AND2_X1 U145 ( .A1(b[1]), .A2(a[0]), .ZN(y[1]) );
  OR2_X1 U145bar ( .A1(bbar[1]), .A2(abar[0]), .ZN(ybar[1]);
  AND2_X1 U146 ( .A1(a[1]), .A2(b[3]), .ZN(y[19]) );
  OR2_X1 U146bar ( .A1(abar[1]), .A2(bbar[3]), .ZN(ybar[19]);
  AND2_X1 U147 ( .A1(a[12]), .A2(b[7]), .ZN(y[199]) );
  OR2_X1 U147bar ( .A1(abar[12]), .A2(bbar[7]), .ZN(ybar[199]);
  AND2_X1 U148 ( .A1(a[12]), .A2(b[6]), .ZN(y[198]) );
  OR2_X1 U148bar ( .A1(abar[12]), .A2(bbar[6]), .ZN(ybar[198]);
  AND2_X1 U149 ( .A1(a[12]), .A2(b[5]), .ZN(y[197]) );
  OR2_X1 U149bar ( .A1(abar[12]), .A2(bbar[5]), .ZN(ybar[197]);
  AND2_X1 U150 ( .A1(a[12]), .A2(b[4]), .ZN(y[196]) );
  OR2_X1 U150bar ( .A1(abar[12]), .A2(bbar[4]), .ZN(ybar[196]);
  AND2_X1 U151 ( .A1(a[12]), .A2(b[3]), .ZN(y[195]) );
  OR2_X1 U151bar ( .A1(abar[12]), .A2(bbar[3]), .ZN(ybar[195]);
  AND2_X1 U152 ( .A1(a[12]), .A2(b[2]), .ZN(y[194]) );
  OR2_X1 U152bar ( .A1(abar[12]), .A2(bbar[2]), .ZN(ybar[194]);
  AND2_X1 U153 ( .A1(a[12]), .A2(b[1]), .ZN(y[193]) );
  OR2_X1 U153bar ( .A1(abar[12]), .A2(bbar[1]), .ZN(ybar[193]);
  AND2_X1 U154 ( .A1(a[12]), .A2(b[0]), .ZN(y[192]) );
  OR2_X1 U154bar ( .A1(abar[12]), .A2(bbar[0]), .ZN(ybar[192]);
  AND2_X1 U155 ( .A1(a[11]), .A2(b[15]), .ZN(y[191]) );
  OR2_X1 U155bar ( .A1(abar[11]), .A2(bbar[15]), .ZN(ybar[191]);
  AND2_X1 U156 ( .A1(a[11]), .A2(b[14]), .ZN(y[190]) );
  OR2_X1 U156bar ( .A1(abar[11]), .A2(bbar[14]), .ZN(ybar[190]);
  AND2_X1 U157 ( .A1(a[1]), .A2(b[2]), .ZN(y[18]) );
  OR2_X1 U157bar ( .A1(abar[1]), .A2(bbar[2]), .ZN(ybar[18]);
  AND2_X1 U158 ( .A1(a[11]), .A2(b[13]), .ZN(y[189]) );
  OR2_X1 U158bar ( .A1(abar[11]), .A2(bbar[13]), .ZN(ybar[189]);
  AND2_X1 U159 ( .A1(a[11]), .A2(b[12]), .ZN(y[188]) );
  OR2_X1 U159bar ( .A1(abar[11]), .A2(bbar[12]), .ZN(ybar[188]);
  AND2_X1 U160 ( .A1(a[11]), .A2(b[11]), .ZN(y[187]) );
  OR2_X1 U160bar ( .A1(abar[11]), .A2(bbar[11]), .ZN(ybar[187]);
  AND2_X1 U161 ( .A1(a[11]), .A2(b[10]), .ZN(y[186]) );
  OR2_X1 U161bar ( .A1(abar[11]), .A2(bbar[10]), .ZN(ybar[186]);
  AND2_X1 U162 ( .A1(a[11]), .A2(b[9]), .ZN(y[185]) );
  OR2_X1 U162bar ( .A1(abar[11]), .A2(bbar[9]), .ZN(ybar[185]);
  AND2_X1 U163 ( .A1(a[11]), .A2(b[8]), .ZN(y[184]) );
  OR2_X1 U163bar ( .A1(abar[11]), .A2(bbar[8]), .ZN(ybar[184]);
  AND2_X1 U164 ( .A1(a[11]), .A2(b[7]), .ZN(y[183]) );
  OR2_X1 U164bar ( .A1(abar[11]), .A2(bbar[7]), .ZN(ybar[183]);
  AND2_X1 U165 ( .A1(a[11]), .A2(b[6]), .ZN(y[182]) );
  OR2_X1 U165bar ( .A1(abar[11]), .A2(bbar[6]), .ZN(ybar[182]);
  AND2_X1 U166 ( .A1(a[11]), .A2(b[5]), .ZN(y[181]) );
  OR2_X1 U166bar ( .A1(abar[11]), .A2(bbar[5]), .ZN(ybar[181]);
  AND2_X1 U167 ( .A1(a[11]), .A2(b[4]), .ZN(y[180]) );
  OR2_X1 U167bar ( .A1(abar[11]), .A2(bbar[4]), .ZN(ybar[180]);
  AND2_X1 U168 ( .A1(a[1]), .A2(b[1]), .ZN(y[17]) );
  OR2_X1 U168bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[17]);
  AND2_X1 U169 ( .A1(a[11]), .A2(b[3]), .ZN(y[179]) );
  OR2_X1 U169bar ( .A1(abar[11]), .A2(bbar[3]), .ZN(ybar[179]);
  AND2_X1 U170 ( .A1(a[11]), .A2(b[2]), .ZN(y[178]) );
  OR2_X1 U170bar ( .A1(abar[11]), .A2(bbar[2]), .ZN(ybar[178]);
  AND2_X1 U171 ( .A1(a[11]), .A2(b[1]), .ZN(y[177]) );
  OR2_X1 U171bar ( .A1(abar[11]), .A2(bbar[1]), .ZN(ybar[177]);
  AND2_X1 U172 ( .A1(a[11]), .A2(b[0]), .ZN(y[176]) );
  OR2_X1 U172bar ( .A1(abar[11]), .A2(bbar[0]), .ZN(ybar[176]);
  AND2_X1 U173 ( .A1(a[10]), .A2(b[15]), .ZN(y[175]) );
  OR2_X1 U173bar ( .A1(abar[10]), .A2(bbar[15]), .ZN(ybar[175]);
  AND2_X1 U174 ( .A1(a[10]), .A2(b[14]), .ZN(y[174]) );
  OR2_X1 U174bar ( .A1(abar[10]), .A2(bbar[14]), .ZN(ybar[174]);
  AND2_X1 U175 ( .A1(a[10]), .A2(b[13]), .ZN(y[173]) );
  OR2_X1 U175bar ( .A1(abar[10]), .A2(bbar[13]), .ZN(ybar[173]);
  AND2_X1 U176 ( .A1(a[10]), .A2(b[12]), .ZN(y[172]) );
  OR2_X1 U176bar ( .A1(abar[10]), .A2(bbar[12]), .ZN(ybar[172]);
  AND2_X1 U177 ( .A1(a[10]), .A2(b[11]), .ZN(y[171]) );
  OR2_X1 U177bar ( .A1(abar[10]), .A2(bbar[11]), .ZN(ybar[171]);
  AND2_X1 U178 ( .A1(a[10]), .A2(b[10]), .ZN(y[170]) );
  OR2_X1 U178bar ( .A1(abar[10]), .A2(bbar[10]), .ZN(ybar[170]);
  AND2_X1 U179 ( .A1(a[1]), .A2(b[0]), .ZN(y[16]) );
  OR2_X1 U179bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[16]);
  AND2_X1 U180 ( .A1(a[10]), .A2(b[9]), .ZN(y[169]) );
  OR2_X1 U180bar ( .A1(abar[10]), .A2(bbar[9]), .ZN(ybar[169]);
  AND2_X1 U181 ( .A1(a[10]), .A2(b[8]), .ZN(y[168]) );
  OR2_X1 U181bar ( .A1(abar[10]), .A2(bbar[8]), .ZN(ybar[168]);
  AND2_X1 U182 ( .A1(a[10]), .A2(b[7]), .ZN(y[167]) );
  OR2_X1 U182bar ( .A1(abar[10]), .A2(bbar[7]), .ZN(ybar[167]);
  AND2_X1 U183 ( .A1(a[10]), .A2(b[6]), .ZN(y[166]) );
  OR2_X1 U183bar ( .A1(abar[10]), .A2(bbar[6]), .ZN(ybar[166]);
  AND2_X1 U184 ( .A1(a[10]), .A2(b[5]), .ZN(y[165]) );
  OR2_X1 U184bar ( .A1(abar[10]), .A2(bbar[5]), .ZN(ybar[165]);
  AND2_X1 U185 ( .A1(a[10]), .A2(b[4]), .ZN(y[164]) );
  OR2_X1 U185bar ( .A1(abar[10]), .A2(bbar[4]), .ZN(ybar[164]);
  AND2_X1 U186 ( .A1(a[10]), .A2(b[3]), .ZN(y[163]) );
  OR2_X1 U186bar ( .A1(abar[10]), .A2(bbar[3]), .ZN(ybar[163]);
  AND2_X1 U187 ( .A1(a[10]), .A2(b[2]), .ZN(y[162]) );
  OR2_X1 U187bar ( .A1(abar[10]), .A2(bbar[2]), .ZN(ybar[162]);
  AND2_X1 U188 ( .A1(a[10]), .A2(b[1]), .ZN(y[161]) );
  OR2_X1 U188bar ( .A1(abar[10]), .A2(bbar[1]), .ZN(ybar[161]);
  AND2_X1 U189 ( .A1(a[10]), .A2(b[0]), .ZN(y[160]) );
  OR2_X1 U189bar ( .A1(abar[10]), .A2(bbar[0]), .ZN(ybar[160]);
  AND2_X1 U190 ( .A1(b[15]), .A2(a[0]), .ZN(y[15]) );
  OR2_X1 U190bar ( .A1(bbar[15]), .A2(abar[0]), .ZN(ybar[15]);
  AND2_X1 U191 ( .A1(a[9]), .A2(b[15]), .ZN(y[159]) );
  OR2_X1 U191bar ( .A1(abar[9]), .A2(bbar[15]), .ZN(ybar[159]);
  AND2_X1 U192 ( .A1(a[9]), .A2(b[14]), .ZN(y[158]) );
  OR2_X1 U192bar ( .A1(abar[9]), .A2(bbar[14]), .ZN(ybar[158]);
  AND2_X1 U193 ( .A1(a[9]), .A2(b[13]), .ZN(y[157]) );
  OR2_X1 U193bar ( .A1(abar[9]), .A2(bbar[13]), .ZN(ybar[157]);
  AND2_X1 U194 ( .A1(a[9]), .A2(b[12]), .ZN(y[156]) );
  OR2_X1 U194bar ( .A1(abar[9]), .A2(bbar[12]), .ZN(ybar[156]);
  AND2_X1 U195 ( .A1(a[9]), .A2(b[11]), .ZN(y[155]) );
  OR2_X1 U195bar ( .A1(abar[9]), .A2(bbar[11]), .ZN(ybar[155]);
  AND2_X1 U196 ( .A1(a[9]), .A2(b[10]), .ZN(y[154]) );
  OR2_X1 U196bar ( .A1(abar[9]), .A2(bbar[10]), .ZN(ybar[154]);
  AND2_X1 U197 ( .A1(a[9]), .A2(b[9]), .ZN(y[153]) );
  OR2_X1 U197bar ( .A1(abar[9]), .A2(bbar[9]), .ZN(ybar[153]);
  AND2_X1 U198 ( .A1(a[9]), .A2(b[8]), .ZN(y[152]) );
  OR2_X1 U198bar ( .A1(abar[9]), .A2(bbar[8]), .ZN(ybar[152]);
  AND2_X1 U199 ( .A1(a[9]), .A2(b[7]), .ZN(y[151]) );
  OR2_X1 U199bar ( .A1(abar[9]), .A2(bbar[7]), .ZN(ybar[151]);
  AND2_X1 U200 ( .A1(a[9]), .A2(b[6]), .ZN(y[150]) );
  OR2_X1 U200bar ( .A1(abar[9]), .A2(bbar[6]), .ZN(ybar[150]);
  AND2_X1 U201 ( .A1(b[14]), .A2(a[0]), .ZN(y[14]) );
  OR2_X1 U201bar ( .A1(bbar[14]), .A2(abar[0]), .ZN(ybar[14]);
  AND2_X1 U202 ( .A1(a[9]), .A2(b[5]), .ZN(y[149]) );
  OR2_X1 U202bar ( .A1(abar[9]), .A2(bbar[5]), .ZN(ybar[149]);
  AND2_X1 U203 ( .A1(a[9]), .A2(b[4]), .ZN(y[148]) );
  OR2_X1 U203bar ( .A1(abar[9]), .A2(bbar[4]), .ZN(ybar[148]);
  AND2_X1 U204 ( .A1(a[9]), .A2(b[3]), .ZN(y[147]) );
  OR2_X1 U204bar ( .A1(abar[9]), .A2(bbar[3]), .ZN(ybar[147]);
  AND2_X1 U205 ( .A1(a[9]), .A2(b[2]), .ZN(y[146]) );
  OR2_X1 U205bar ( .A1(abar[9]), .A2(bbar[2]), .ZN(ybar[146]);
  AND2_X1 U206 ( .A1(a[9]), .A2(b[1]), .ZN(y[145]) );
  OR2_X1 U206bar ( .A1(abar[9]), .A2(bbar[1]), .ZN(ybar[145]);
  AND2_X1 U207 ( .A1(a[9]), .A2(b[0]), .ZN(y[144]) );
  OR2_X1 U207bar ( .A1(abar[9]), .A2(bbar[0]), .ZN(ybar[144]);
  AND2_X1 U208 ( .A1(a[8]), .A2(b[15]), .ZN(y[143]) );
  OR2_X1 U208bar ( .A1(abar[8]), .A2(bbar[15]), .ZN(ybar[143]);
  AND2_X1 U209 ( .A1(a[8]), .A2(b[14]), .ZN(y[142]) );
  OR2_X1 U209bar ( .A1(abar[8]), .A2(bbar[14]), .ZN(ybar[142]);
  AND2_X1 U210 ( .A1(a[8]), .A2(b[13]), .ZN(y[141]) );
  OR2_X1 U210bar ( .A1(abar[8]), .A2(bbar[13]), .ZN(ybar[141]);
  AND2_X1 U211 ( .A1(a[8]), .A2(b[12]), .ZN(y[140]) );
  OR2_X1 U211bar ( .A1(abar[8]), .A2(bbar[12]), .ZN(ybar[140]);
  AND2_X1 U212 ( .A1(b[13]), .A2(a[0]), .ZN(y[13]) );
  OR2_X1 U212bar ( .A1(bbar[13]), .A2(abar[0]), .ZN(ybar[13]);
  AND2_X1 U213 ( .A1(a[8]), .A2(b[11]), .ZN(y[139]) );
  OR2_X1 U213bar ( .A1(abar[8]), .A2(bbar[11]), .ZN(ybar[139]);
  AND2_X1 U214 ( .A1(a[8]), .A2(b[10]), .ZN(y[138]) );
  OR2_X1 U214bar ( .A1(abar[8]), .A2(bbar[10]), .ZN(ybar[138]);
  AND2_X1 U215 ( .A1(a[8]), .A2(b[9]), .ZN(y[137]) );
  OR2_X1 U215bar ( .A1(abar[8]), .A2(bbar[9]), .ZN(ybar[137]);
  AND2_X1 U216 ( .A1(a[8]), .A2(b[8]), .ZN(y[136]) );
  OR2_X1 U216bar ( .A1(abar[8]), .A2(bbar[8]), .ZN(ybar[136]);
  AND2_X1 U217 ( .A1(a[8]), .A2(b[7]), .ZN(y[135]) );
  OR2_X1 U217bar ( .A1(abar[8]), .A2(bbar[7]), .ZN(ybar[135]);
  AND2_X1 U218 ( .A1(a[8]), .A2(b[6]), .ZN(y[134]) );
  OR2_X1 U218bar ( .A1(abar[8]), .A2(bbar[6]), .ZN(ybar[134]);
  AND2_X1 U219 ( .A1(a[8]), .A2(b[5]), .ZN(y[133]) );
  OR2_X1 U219bar ( .A1(abar[8]), .A2(bbar[5]), .ZN(ybar[133]);
  AND2_X1 U220 ( .A1(a[8]), .A2(b[4]), .ZN(y[132]) );
  OR2_X1 U220bar ( .A1(abar[8]), .A2(bbar[4]), .ZN(ybar[132]);
  AND2_X1 U221 ( .A1(a[8]), .A2(b[3]), .ZN(y[131]) );
  OR2_X1 U221bar ( .A1(abar[8]), .A2(bbar[3]), .ZN(ybar[131]);
  AND2_X1 U222 ( .A1(a[8]), .A2(b[2]), .ZN(y[130]) );
  OR2_X1 U222bar ( .A1(abar[8]), .A2(bbar[2]), .ZN(ybar[130]);
  AND2_X1 U223 ( .A1(b[12]), .A2(a[0]), .ZN(y[12]) );
  OR2_X1 U223bar ( .A1(bbar[12]), .A2(abar[0]), .ZN(ybar[12]);
  AND2_X1 U224 ( .A1(a[8]), .A2(b[1]), .ZN(y[129]) );
  OR2_X1 U224bar ( .A1(abar[8]), .A2(bbar[1]), .ZN(ybar[129]);
  AND2_X1 U225 ( .A1(a[8]), .A2(b[0]), .ZN(y[128]) );
  OR2_X1 U225bar ( .A1(abar[8]), .A2(bbar[0]), .ZN(ybar[128]);
  AND2_X1 U226 ( .A1(a[7]), .A2(b[15]), .ZN(y[127]) );
  OR2_X1 U226bar ( .A1(abar[7]), .A2(bbar[15]), .ZN(ybar[127]);
  AND2_X1 U227 ( .A1(a[7]), .A2(b[14]), .ZN(y[126]) );
  OR2_X1 U227bar ( .A1(abar[7]), .A2(bbar[14]), .ZN(ybar[126]);
  AND2_X1 U228 ( .A1(a[7]), .A2(b[13]), .ZN(y[125]) );
  OR2_X1 U228bar ( .A1(abar[7]), .A2(bbar[13]), .ZN(ybar[125]);
  AND2_X1 U229 ( .A1(a[7]), .A2(b[12]), .ZN(y[124]) );
  OR2_X1 U229bar ( .A1(abar[7]), .A2(bbar[12]), .ZN(ybar[124]);
  AND2_X1 U230 ( .A1(a[7]), .A2(b[11]), .ZN(y[123]) );
  OR2_X1 U230bar ( .A1(abar[7]), .A2(bbar[11]), .ZN(ybar[123]);
  AND2_X1 U231 ( .A1(a[7]), .A2(b[10]), .ZN(y[122]) );
  OR2_X1 U231bar ( .A1(abar[7]), .A2(bbar[10]), .ZN(ybar[122]);
  AND2_X1 U232 ( .A1(a[7]), .A2(b[9]), .ZN(y[121]) );
  OR2_X1 U232bar ( .A1(abar[7]), .A2(bbar[9]), .ZN(ybar[121]);
  AND2_X1 U233 ( .A1(a[7]), .A2(b[8]), .ZN(y[120]) );
  OR2_X1 U233bar ( .A1(abar[7]), .A2(bbar[8]), .ZN(ybar[120]);
  AND2_X1 U234 ( .A1(b[11]), .A2(a[0]), .ZN(y[11]) );
  OR2_X1 U234bar ( .A1(bbar[11]), .A2(abar[0]), .ZN(ybar[11]);
  AND2_X1 U235 ( .A1(a[7]), .A2(b[7]), .ZN(y[119]) );
  OR2_X1 U235bar ( .A1(abar[7]), .A2(bbar[7]), .ZN(ybar[119]);
  AND2_X1 U236 ( .A1(a[7]), .A2(b[6]), .ZN(y[118]) );
  OR2_X1 U236bar ( .A1(abar[7]), .A2(bbar[6]), .ZN(ybar[118]);
  AND2_X1 U237 ( .A1(a[7]), .A2(b[5]), .ZN(y[117]) );
  OR2_X1 U237bar ( .A1(abar[7]), .A2(bbar[5]), .ZN(ybar[117]);
  AND2_X1 U238 ( .A1(a[7]), .A2(b[4]), .ZN(y[116]) );
  OR2_X1 U238bar ( .A1(abar[7]), .A2(bbar[4]), .ZN(ybar[116]);
  AND2_X1 U239 ( .A1(a[7]), .A2(b[3]), .ZN(y[115]) );
  OR2_X1 U239bar ( .A1(abar[7]), .A2(bbar[3]), .ZN(ybar[115]);
  AND2_X1 U240 ( .A1(a[7]), .A2(b[2]), .ZN(y[114]) );
  OR2_X1 U240bar ( .A1(abar[7]), .A2(bbar[2]), .ZN(ybar[114]);
  AND2_X1 U241 ( .A1(a[7]), .A2(b[1]), .ZN(y[113]) );
  OR2_X1 U241bar ( .A1(abar[7]), .A2(bbar[1]), .ZN(ybar[113]);
  AND2_X1 U242 ( .A1(a[7]), .A2(b[0]), .ZN(y[112]) );
  OR2_X1 U242bar ( .A1(abar[7]), .A2(bbar[0]), .ZN(ybar[112]);
  AND2_X1 U243 ( .A1(b[15]), .A2(a[6]), .ZN(y[111]) );
  OR2_X1 U243bar ( .A1(bbar[15]), .A2(abar[6]), .ZN(ybar[111]);
  AND2_X1 U244 ( .A1(b[14]), .A2(a[6]), .ZN(y[110]) );
  OR2_X1 U244bar ( .A1(bbar[14]), .A2(abar[6]), .ZN(ybar[110]);
  AND2_X1 U245 ( .A1(b[10]), .A2(a[0]), .ZN(y[10]) );
  OR2_X1 U245bar ( .A1(bbar[10]), .A2(abar[0]), .ZN(ybar[10]);
  AND2_X1 U246 ( .A1(b[13]), .A2(a[6]), .ZN(y[109]) );
  OR2_X1 U246bar ( .A1(bbar[13]), .A2(abar[6]), .ZN(ybar[109]);
  AND2_X1 U247 ( .A1(b[12]), .A2(a[6]), .ZN(y[108]) );
  OR2_X1 U247bar ( .A1(bbar[12]), .A2(abar[6]), .ZN(ybar[108]);
  AND2_X1 U248 ( .A1(b[11]), .A2(a[6]), .ZN(y[107]) );
  OR2_X1 U248bar ( .A1(bbar[11]), .A2(abar[6]), .ZN(ybar[107]);
  AND2_X1 U249 ( .A1(b[10]), .A2(a[6]), .ZN(y[106]) );
  OR2_X1 U249bar ( .A1(bbar[10]), .A2(abar[6]), .ZN(ybar[106]);
  AND2_X1 U250 ( .A1(a[6]), .A2(b[9]), .ZN(y[105]) );
  OR2_X1 U250bar ( .A1(abar[6]), .A2(bbar[9]), .ZN(ybar[105]);
  AND2_X1 U251 ( .A1(b[8]), .A2(a[6]), .ZN(y[104]) );
  OR2_X1 U251bar ( .A1(bbar[8]), .A2(abar[6]), .ZN(ybar[104]);
  AND2_X1 U252 ( .A1(b[7]), .A2(a[6]), .ZN(y[103]) );
  OR2_X1 U252bar ( .A1(bbar[7]), .A2(abar[6]), .ZN(ybar[103]);
  AND2_X1 U253 ( .A1(b[6]), .A2(a[6]), .ZN(y[102]) );
  OR2_X1 U253bar ( .A1(bbar[6]), .A2(abar[6]), .ZN(ybar[102]);
  AND2_X1 U254 ( .A1(b[5]), .A2(a[6]), .ZN(y[101]) );
  OR2_X1 U254bar ( .A1(bbar[5]), .A2(abar[6]), .ZN(ybar[101]);
  AND2_X1 U255 ( .A1(b[4]), .A2(a[6]), .ZN(y[100]) );
  OR2_X1 U255bar ( .A1(bbar[4]), .A2(abar[6]), .ZN(ybar[100]);
  AND2_X1 U256 ( .A1(b[0]), .A2(a[0]), .ZN(y[0]) );
  OR2_X1 U256bar ( .A1(bbar[0]), .A2(abar[0]), .ZN(ybar[0]);
endmodule




module decode_5 ( in, out );
  input [7:0] in;
  //input_done

  output [255:0] out;
  //output_done

  wire   [15:0] level1;
  wire   [31:0] level2;
  //wire_done

  CD2_20 cd_l1_1 ( .a(in[1]), .b(in[0]), .y(level1[3:0]) );
  CD2_19 cd_l1_2 ( .a(in[3]), .b(in[2]), .y(level1[7:4]) );
  CD2_18 cd_l1_3 ( .a(in[5]), .b(in[4]), .y(level1[11:8]) );
  CD2_17 cd_l1_4 ( .a(in[7]), .b(in[6]), .y(level1[15:12]) );
  CD4_10 cd_l2_1 ( .a(level1[7:4]), .b(level1[3:0]), .y(level2[15:0]) );
  CD4_9 cd_l2_2 ( .a(level1[15:12]), .b(level1[11:8]), .y(level2[31:16]) );
  CD16_5 cd_l3 ( .a(level2[31:16]), .b(level2[15:0]), .y(out) );
endmodule


module encode_5 ( in, out );
  input [255:0] in;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
  assign inbar[8] = ~in[8];
  assign inbar[9] = ~in[9];
  assign inbar[10] = ~in[10];
  assign inbar[11] = ~in[11];
  assign inbar[12] = ~in[12];
  assign inbar[13] = ~in[13];
  assign inbar[14] = ~in[14];
  assign inbar[15] = ~in[15];
  assign inbar[16] = ~in[16];
  assign inbar[17] = ~in[17];
  assign inbar[18] = ~in[18];
  assign inbar[19] = ~in[19];
  assign inbar[20] = ~in[20];
  assign inbar[21] = ~in[21];
  assign inbar[22] = ~in[22];
  assign inbar[23] = ~in[23];
  assign inbar[24] = ~in[24];
  assign inbar[25] = ~in[25];
  assign inbar[26] = ~in[26];
  assign inbar[27] = ~in[27];
  assign inbar[28] = ~in[28];
  assign inbar[29] = ~in[29];
  assign inbar[30] = ~in[30];
  assign inbar[31] = ~in[31];
  assign inbar[32] = ~in[32];
  assign inbar[33] = ~in[33];
  assign inbar[34] = ~in[34];
  assign inbar[35] = ~in[35];
  assign inbar[36] = ~in[36];
  assign inbar[37] = ~in[37];
  assign inbar[38] = ~in[38];
  assign inbar[39] = ~in[39];
  assign inbar[40] = ~in[40];
  assign inbar[41] = ~in[41];
  assign inbar[42] = ~in[42];
  assign inbar[43] = ~in[43];
  assign inbar[44] = ~in[44];
  assign inbar[45] = ~in[45];
  assign inbar[46] = ~in[46];
  assign inbar[47] = ~in[47];
  assign inbar[48] = ~in[48];
  assign inbar[49] = ~in[49];
  assign inbar[50] = ~in[50];
  assign inbar[51] = ~in[51];
  assign inbar[52] = ~in[52];
  assign inbar[53] = ~in[53];
  assign inbar[54] = ~in[54];
  assign inbar[55] = ~in[55];
  assign inbar[56] = ~in[56];
  assign inbar[57] = ~in[57];
  assign inbar[58] = ~in[58];
  assign inbar[59] = ~in[59];
  assign inbar[60] = ~in[60];
  assign inbar[61] = ~in[61];
  assign inbar[62] = ~in[62];
  assign inbar[63] = ~in[63];
  assign inbar[64] = ~in[64];
  assign inbar[65] = ~in[65];
  assign inbar[66] = ~in[66];
  assign inbar[67] = ~in[67];
  assign inbar[68] = ~in[68];
  assign inbar[69] = ~in[69];
  assign inbar[70] = ~in[70];
  assign inbar[71] = ~in[71];
  assign inbar[72] = ~in[72];
  assign inbar[73] = ~in[73];
  assign inbar[74] = ~in[74];
  assign inbar[75] = ~in[75];
  assign inbar[76] = ~in[76];
  assign inbar[77] = ~in[77];
  assign inbar[78] = ~in[78];
  assign inbar[79] = ~in[79];
  assign inbar[80] = ~in[80];
  assign inbar[81] = ~in[81];
  assign inbar[82] = ~in[82];
  assign inbar[83] = ~in[83];
  assign inbar[84] = ~in[84];
  assign inbar[85] = ~in[85];
  assign inbar[86] = ~in[86];
  assign inbar[87] = ~in[87];
  assign inbar[88] = ~in[88];
  assign inbar[89] = ~in[89];
  assign inbar[90] = ~in[90];
  assign inbar[91] = ~in[91];
  assign inbar[92] = ~in[92];
  assign inbar[93] = ~in[93];
  assign inbar[94] = ~in[94];
  assign inbar[95] = ~in[95];
  assign inbar[96] = ~in[96];
  assign inbar[97] = ~in[97];
  assign inbar[98] = ~in[98];
  assign inbar[99] = ~in[99];
  assign inbar[100] = ~in[100];
  assign inbar[101] = ~in[101];
  assign inbar[102] = ~in[102];
  assign inbar[103] = ~in[103];
  assign inbar[104] = ~in[104];
  assign inbar[105] = ~in[105];
  assign inbar[106] = ~in[106];
  assign inbar[107] = ~in[107];
  assign inbar[108] = ~in[108];
  assign inbar[109] = ~in[109];
  assign inbar[110] = ~in[110];
  assign inbar[111] = ~in[111];
  assign inbar[112] = ~in[112];
  assign inbar[113] = ~in[113];
  assign inbar[114] = ~in[114];
  assign inbar[115] = ~in[115];
  assign inbar[116] = ~in[116];
  assign inbar[117] = ~in[117];
  assign inbar[118] = ~in[118];
  assign inbar[119] = ~in[119];
  assign inbar[120] = ~in[120];
  assign inbar[121] = ~in[121];
  assign inbar[122] = ~in[122];
  assign inbar[123] = ~in[123];
  assign inbar[124] = ~in[124];
  assign inbar[125] = ~in[125];
  assign inbar[126] = ~in[126];
  assign inbar[127] = ~in[127];
  assign inbar[128] = ~in[128];
  assign inbar[129] = ~in[129];
  assign inbar[130] = ~in[130];
  assign inbar[131] = ~in[131];
  assign inbar[132] = ~in[132];
  assign inbar[133] = ~in[133];
  assign inbar[134] = ~in[134];
  assign inbar[135] = ~in[135];
  assign inbar[136] = ~in[136];
  assign inbar[137] = ~in[137];
  assign inbar[138] = ~in[138];
  assign inbar[139] = ~in[139];
  assign inbar[140] = ~in[140];
  assign inbar[141] = ~in[141];
  assign inbar[142] = ~in[142];
  assign inbar[143] = ~in[143];
  assign inbar[144] = ~in[144];
  assign inbar[145] = ~in[145];
  assign inbar[146] = ~in[146];
  assign inbar[147] = ~in[147];
  assign inbar[148] = ~in[148];
  assign inbar[149] = ~in[149];
  assign inbar[150] = ~in[150];
  assign inbar[151] = ~in[151];
  assign inbar[152] = ~in[152];
  assign inbar[153] = ~in[153];
  assign inbar[154] = ~in[154];
  assign inbar[155] = ~in[155];
  assign inbar[156] = ~in[156];
  assign inbar[157] = ~in[157];
  assign inbar[158] = ~in[158];
  assign inbar[159] = ~in[159];
  assign inbar[160] = ~in[160];
  assign inbar[161] = ~in[161];
  assign inbar[162] = ~in[162];
  assign inbar[163] = ~in[163];
  assign inbar[164] = ~in[164];
  assign inbar[165] = ~in[165];
  assign inbar[166] = ~in[166];
  assign inbar[167] = ~in[167];
  assign inbar[168] = ~in[168];
  assign inbar[169] = ~in[169];
  assign inbar[170] = ~in[170];
  assign inbar[171] = ~in[171];
  assign inbar[172] = ~in[172];
  assign inbar[173] = ~in[173];
  assign inbar[174] = ~in[174];
  assign inbar[175] = ~in[175];
  assign inbar[176] = ~in[176];
  assign inbar[177] = ~in[177];
  assign inbar[178] = ~in[178];
  assign inbar[179] = ~in[179];
  assign inbar[180] = ~in[180];
  assign inbar[181] = ~in[181];
  assign inbar[182] = ~in[182];
  assign inbar[183] = ~in[183];
  assign inbar[184] = ~in[184];
  assign inbar[185] = ~in[185];
  assign inbar[186] = ~in[186];
  assign inbar[187] = ~in[187];
  assign inbar[188] = ~in[188];
  assign inbar[189] = ~in[189];
  assign inbar[190] = ~in[190];
  assign inbar[191] = ~in[191];
  assign inbar[192] = ~in[192];
  assign inbar[193] = ~in[193];
  assign inbar[194] = ~in[194];
  assign inbar[195] = ~in[195];
  assign inbar[196] = ~in[196];
  assign inbar[197] = ~in[197];
  assign inbar[198] = ~in[198];
  assign inbar[199] = ~in[199];
  assign inbar[200] = ~in[200];
  assign inbar[201] = ~in[201];
  assign inbar[202] = ~in[202];
  assign inbar[203] = ~in[203];
  assign inbar[204] = ~in[204];
  assign inbar[205] = ~in[205];
  assign inbar[206] = ~in[206];
  assign inbar[207] = ~in[207];
  assign inbar[208] = ~in[208];
  assign inbar[209] = ~in[209];
  assign inbar[210] = ~in[210];
  assign inbar[211] = ~in[211];
  assign inbar[212] = ~in[212];
  assign inbar[213] = ~in[213];
  assign inbar[214] = ~in[214];
  assign inbar[215] = ~in[215];
  assign inbar[216] = ~in[216];
  assign inbar[217] = ~in[217];
  assign inbar[218] = ~in[218];
  assign inbar[219] = ~in[219];
  assign inbar[220] = ~in[220];
  assign inbar[221] = ~in[221];
  assign inbar[222] = ~in[222];
  assign inbar[223] = ~in[223];
  assign inbar[224] = ~in[224];
  assign inbar[225] = ~in[225];
  assign inbar[226] = ~in[226];
  assign inbar[227] = ~in[227];
  assign inbar[228] = ~in[228];
  assign inbar[229] = ~in[229];
  assign inbar[230] = ~in[230];
  assign inbar[231] = ~in[231];
  assign inbar[232] = ~in[232];
  assign inbar[233] = ~in[233];
  assign inbar[234] = ~in[234];
  assign inbar[235] = ~in[235];
  assign inbar[236] = ~in[236];
  assign inbar[237] = ~in[237];
  assign inbar[238] = ~in[238];
  assign inbar[239] = ~in[239];
  assign inbar[240] = ~in[240];
  assign inbar[241] = ~in[241];
  assign inbar[242] = ~in[242];
  assign inbar[243] = ~in[243];
  assign inbar[244] = ~in[244];
  assign inbar[245] = ~in[245];
  assign inbar[246] = ~in[246];
  assign inbar[247] = ~in[247];
  assign inbar[248] = ~in[248];
  assign inbar[249] = ~in[249];
  assign inbar[250] = ~in[250];
  assign inbar[251] = ~in[251];
  assign inbar[252] = ~in[252];
  assign inbar[253] = ~in[253];
  assign inbar[254] = ~in[254];
  assign inbar[255] = ~in[255];
  //input_done

  output [7:0] out;
  reg [7:0] outbar;
  //output_done

  wire   in_81, in_80, in_79, in_78, in_77, in_76, in_75, in_74, in_73, in_72,
         in_71, in_70, in_69, in_68, in_67, in_66, in_65, in_64, in_63, in_62,
         in_61, in_60, in_59, in_58, in_57, in_56, in_55, in_54, in_53, in_52,
         in_51, in_50, in_49, in_48, in_47, in_46, in_45, in_44, in_43, in_42,
         in_41, in_40, in_39, in_38, in_37, in_36, in_35, in_34, in_33, in_32,
         in_31, in_30, in_29, in_28, in_27, in_26, in_25, in_24, in_23, in_22,
         in_21, in_20, in_19, in_18, in_17, in_16, in_15, in_14, in_13, in_12,
         in_11, in_10, in_9, in_8, in_7, in_6, in_5, in_4, in_3, in_2, in_1,
         in_0, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972;
  wire in_81bar, in_80bar, in_79bar, in_78bar, in_77bar, in_76bar, in_75bar, in_74bar, in_73bar, in_72bar, in_71bar, in_70bar, in_69bar, in_68bar, in_67bar, in_66bar, in_65bar, in_64bar, in_63bar, in_62bar, in_61bar, in_60bar, in_59bar, in_58bar, in_57bar, in_56bar, in_55bar, in_54bar, in_53bar, in_52bar, in_51bar, in_50bar, in_49bar, in_48bar, in_47bar, in_46bar, in_45bar, in_44bar, in_43bar, in_42bar, in_41bar, in_40bar, in_39bar, in_38bar, in_37bar, in_36bar, in_35bar, in_34bar, in_33bar, in_32bar, in_31bar, in_30bar, in_29bar, in_28bar, in_27bar, in_26bar, in_25bar, in_24bar, in_23bar, in_22bar, in_21bar, in_20bar, in_19bar, in_18bar, in_17bar, in_16bar, in_15bar, in_14bar, in_13bar, in_12bar, in_11bar, in_10bar, in_9bar, in_8bar, in_7bar, in_6bar, in_5bar, in_4bar, in_3bar, in_2bar, in_1bar, in_0bar, n487bar, n488bar, n489bar, n490bar, n491bar, n492bar, n493bar, n494bar, n495bar, n496bar, n497bar, n498bar, n499bar, n500bar, n501bar, n502bar, n503bar, n504bar, n505bar, n506bar, n507bar, n508bar, n509bar, n510bar, n511bar, n512bar, n513bar, n514bar, n515bar, n516bar, n517bar, n518bar, n519bar, n520bar, n521bar, n522bar, n523bar, n524bar, n525bar, n526bar, n527bar, n528bar, n529bar, n530bar, n531bar, n532bar, n533bar, n534bar, n535bar, n536bar, n537bar, n538bar, n539bar, n540bar, n541bar, n542bar, n543bar, n544bar, n545bar, n546bar, n547bar, n548bar, n549bar, n550bar, n551bar, n552bar, n553bar, n554bar, n555bar, n556bar, n557bar, n558bar, n559bar, n560bar, n561bar, n562bar, n563bar, n564bar, n565bar, n566bar, n567bar, n568bar, n569bar, n570bar, n571bar, n572bar, n573bar, n574bar, n575bar, n576bar, n577bar, n578bar, n579bar, n580bar, n581bar, n582bar, n583bar, n584bar, n585bar, n586bar, n587bar, n588bar, n589bar, n590bar, n591bar, n592bar, n593bar, n594bar, n595bar, n596bar, n597bar, n598bar, n599bar, n600bar, n601bar, n602bar, n603bar, n604bar, n605bar, n606bar, n607bar, n608bar, n609bar, n610bar, n611bar, n612bar, n613bar, n614bar, n615bar, n616bar, n617bar, n618bar, n619bar, n620bar, n621bar, n622bar, n623bar, n624bar, n625bar, n626bar, n627bar, n628bar, n629bar, n630bar, n631bar, n632bar, n633bar, n634bar, n635bar, n636bar, n637bar, n638bar, n639bar, n640bar, n641bar, n642bar, n643bar, n644bar, n645bar, n646bar, n647bar, n648bar, n649bar, n650bar, n651bar, n652bar, n653bar, n654bar, n655bar, n656bar, n657bar, n658bar, n659bar, n660bar, n661bar, n662bar, n663bar, n664bar, n665bar, n666bar, n667bar, n668bar, n669bar, n670bar, n671bar, n672bar, n673bar, n674bar, n675bar, n676bar, n677bar, n678bar, n679bar, n680bar, n681bar, n682bar, n683bar, n684bar, n685bar, n686bar, n687bar, n688bar, n689bar, n690bar, n691bar, n692bar, n693bar, n694bar, n695bar, n696bar, n697bar, n698bar, n699bar, n700bar, n701bar, n702bar, n703bar, n704bar, n705bar, n706bar, n707bar, n708bar, n709bar, n710bar, n711bar, n712bar, n713bar, n714bar, n715bar, n716bar, n717bar, n718bar, n719bar, n720bar, n721bar, n722bar, n723bar, n724bar, n725bar, n726bar, n727bar, n728bar, n729bar, n730bar, n731bar, n732bar, n733bar, n734bar, n735bar, n736bar, n737bar, n738bar, n739bar, n740bar, n741bar, n742bar, n743bar, n744bar, n745bar, n746bar, n747bar, n748bar, n749bar, n750bar, n751bar, n752bar, n753bar, n754bar, n755bar, n756bar, n757bar, n758bar, n759bar, n760bar, n761bar, n762bar, n763bar, n764bar, n765bar, n766bar, n767bar, n768bar, n769bar, n770bar, n771bar, n772bar, n773bar, n774bar, n775bar, n776bar, n777bar, n778bar, n779bar, n780bar, n781bar, n782bar, n783bar, n784bar, n785bar, n786bar, n787bar, n788bar, n789bar, n790bar, n791bar, n792bar, n793bar, n794bar, n795bar, n796bar, n797bar, n798bar, n799bar, n800bar, n801bar, n802bar, n803bar, n804bar, n805bar, n806bar, n807bar, n808bar, n809bar, n810bar, n811bar, n812bar, n813bar, n814bar, n815bar, n816bar, n817bar, n818bar, n819bar, n820bar, n821bar, n822bar, n823bar, n824bar, n825bar, n826bar, n827bar, n828bar, n829bar, n830bar, n831bar, n832bar, n833bar, n834bar, n835bar, n836bar, n837bar, n838bar, n839bar, n840bar, n841bar, n842bar, n843bar, n844bar, n845bar, n846bar, n847bar, n848bar, n849bar, n850bar, n851bar, n852bar, n853bar, n854bar, n855bar, n856bar, n857bar, n858bar, n859bar, n860bar, n861bar, n862bar, n863bar, n864bar, n865bar, n866bar, n867bar, n868bar, n869bar, n870bar, n871bar, n872bar, n873bar, n874bar, n875bar, n876bar, n877bar, n878bar, n879bar, n880bar, n881bar, n882bar, n883bar, n884bar, n885bar, n886bar, n887bar, n888bar, n889bar, n890bar, n891bar, n892bar, n893bar, n894bar, n895bar, n896bar, n897bar, n898bar, n899bar, n900bar, n901bar, n902bar, n903bar, n904bar, n905bar, n906bar, n907bar, n908bar, n909bar, n910bar, n911bar, n912bar, n913bar, n914bar, n915bar, n916bar, n917bar, n918bar, n919bar, n920bar, n921bar, n922bar, n923bar, n924bar, n925bar, n926bar, n927bar, n928bar, n929bar, n930bar, n931bar, n932bar, n933bar, n934bar, n935bar, n936bar, n937bar, n938bar, n939bar, n940bar, n941bar, n942bar, n943bar, n944bar, n945bar, n946bar, n947bar, n948bar, n949bar, n950bar, n951bar, n952bar, n953bar, n954bar, n955bar, n956bar, n957bar, n958bar, n959bar, n960bar, n961bar, n962bar, n963bar, n964bar, n965bar, n966bar, n967bar, n968bar, n969bar, n970bar, n971bar, n972bar;
  //wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];

  OR2_X1 U1 ( .A1(n972), .A2(n971), .ZN(out[7]) );
  AND2_X1 U1bar ( .A1(n972bar), .A2(n971bar), .ZN(outbar[7]);
  OR2_X1 U2 ( .A1(n970), .A2(n969), .ZN(n971) );
  AND2_X1 U2bar ( .A1(n970bar), .A2(n969bar), .ZN(n971bar);
  OR2_X1 U3 ( .A1(n968), .A2(n967), .ZN(n969) );
  AND2_X1 U3bar ( .A1(n968bar), .A2(n967bar), .ZN(n969bar);
  OR2_X1 U4 ( .A1(n966), .A2(n965), .ZN(n967) );
  AND2_X1 U4bar ( .A1(n966bar), .A2(n965bar), .ZN(n967bar);
  OR2_X1 U5 ( .A1(n964), .A2(n963), .ZN(n968) );
  AND2_X1 U5bar ( .A1(n964bar), .A2(n963bar), .ZN(n968bar);
  OR2_X1 U6 ( .A1(in[116]), .A2(n962), .ZN(n963) );
  AND2_X1 U6bar ( .A1(inbar[116]), .A2(n962bar), .ZN(n963bar);
  OR2_X1 U7 ( .A1(n961), .A2(n960), .ZN(n970) );
  AND2_X1 U7bar ( .A1(n961bar), .A2(n960bar), .ZN(n970bar);
  OR2_X1 U8 ( .A1(in[150]), .A2(in[127]), .ZN(n960) );
  AND2_X1 U8bar ( .A1(inbar[150]), .A2(inbar[127]), .ZN(n960bar);
  OR2_X1 U9 ( .A1(in[160]), .A2(n959), .ZN(n961) );
  AND2_X1 U9bar ( .A1(inbar[160]), .A2(n959bar), .ZN(n961bar);
  OR2_X1 U10 ( .A1(in[252]), .A2(in[168]), .ZN(n959) );
  AND2_X1 U10bar ( .A1(inbar[252]), .A2(inbar[168]), .ZN(n959bar);
  OR2_X1 U11 ( .A1(n958), .A2(n957), .ZN(n972) );
  AND2_X1 U11bar ( .A1(n958bar), .A2(n957bar), .ZN(n972bar);
  OR2_X1 U12 ( .A1(n956), .A2(n955), .ZN(n957) );
  AND2_X1 U12bar ( .A1(n956bar), .A2(n955bar), .ZN(n957bar);
  OR2_X1 U13 ( .A1(in_17), .A2(in[96]), .ZN(n955) );
  AND2_X1 U13bar ( .A1(in_17bar), .A2(inbar[96]), .ZN(n955bar);
  OR2_X1 U14 ( .A1(in_23), .A2(n954), .ZN(n956) );
  AND2_X1 U14bar ( .A1(in_23bar), .A2(n954bar), .ZN(n956bar);
  OR2_X1 U15 ( .A1(in_31), .A2(in_26), .ZN(n954) );
  AND2_X1 U15bar ( .A1(in_31bar), .A2(in_26bar), .ZN(n954bar);
  OR2_X1 U16 ( .A1(n953), .A2(n952), .ZN(n958) );
  AND2_X1 U16bar ( .A1(n953bar), .A2(n952bar), .ZN(n958bar);
  OR2_X1 U17 ( .A1(in_58), .A2(in_4), .ZN(n952) );
  AND2_X1 U17bar ( .A1(in_58bar), .A2(in_4bar), .ZN(n952bar);
  OR2_X1 U18 ( .A1(in_59), .A2(n951), .ZN(n953) );
  AND2_X1 U18bar ( .A1(in_59bar), .A2(n951bar), .ZN(n953bar);
  OR2_X1 U19 ( .A1(in_71), .A2(in_62), .ZN(n951) );
  AND2_X1 U19bar ( .A1(in_71bar), .A2(in_62bar), .ZN(n951bar);
  OR2_X1 U20 ( .A1(n950), .A2(n949), .ZN(out[6]) );
  AND2_X1 U20bar ( .A1(n950bar), .A2(n949bar), .ZN(outbar[6]);
  OR2_X1 U21 ( .A1(n948), .A2(n947), .ZN(n949) );
  AND2_X1 U21bar ( .A1(n948bar), .A2(n947bar), .ZN(n949bar);
  OR2_X1 U22 ( .A1(n946), .A2(n945), .ZN(n947) );
  AND2_X1 U22bar ( .A1(n946bar), .A2(n945bar), .ZN(n947bar);
  OR2_X1 U23 ( .A1(n944), .A2(n943), .ZN(n945) );
  AND2_X1 U23bar ( .A1(n944bar), .A2(n943bar), .ZN(n945bar);
  OR2_X1 U24 ( .A1(n942), .A2(n941), .ZN(n946) );
  AND2_X1 U24bar ( .A1(n942bar), .A2(n941bar), .ZN(n946bar);
  OR2_X1 U25 ( .A1(in[101]), .A2(n940), .ZN(n941) );
  AND2_X1 U25bar ( .A1(inbar[101]), .A2(n940bar), .ZN(n941bar);
  OR2_X1 U26 ( .A1(n939), .A2(n938), .ZN(n948) );
  AND2_X1 U26bar ( .A1(n939bar), .A2(n938bar), .ZN(n948bar);
  OR2_X1 U27 ( .A1(in[114]), .A2(in[104]), .ZN(n938) );
  AND2_X1 U27bar ( .A1(inbar[114]), .A2(inbar[104]), .ZN(n938bar);
  OR2_X1 U28 ( .A1(in[128]), .A2(n937), .ZN(n939) );
  AND2_X1 U28bar ( .A1(inbar[128]), .A2(n937bar), .ZN(n939bar);
  OR2_X1 U29 ( .A1(in[136]), .A2(in[134]), .ZN(n937) );
  AND2_X1 U29bar ( .A1(inbar[136]), .A2(inbar[134]), .ZN(n937bar);
  OR2_X1 U30 ( .A1(n936), .A2(n935), .ZN(n950) );
  AND2_X1 U30bar ( .A1(n936bar), .A2(n935bar), .ZN(n950bar);
  OR2_X1 U31 ( .A1(n934), .A2(n933), .ZN(n935) );
  AND2_X1 U31bar ( .A1(n934bar), .A2(n933bar), .ZN(n935bar);
  OR2_X1 U32 ( .A1(in[177]), .A2(in[164]), .ZN(n933) );
  AND2_X1 U32bar ( .A1(inbar[177]), .A2(inbar[164]), .ZN(n933bar);
  OR2_X1 U33 ( .A1(in[212]), .A2(n932), .ZN(n934) );
  AND2_X1 U33bar ( .A1(inbar[212]), .A2(n932bar), .ZN(n934bar);
  OR2_X1 U34 ( .A1(in[248]), .A2(in[221]), .ZN(n932) );
  AND2_X1 U34bar ( .A1(inbar[248]), .A2(inbar[221]), .ZN(n932bar);
  OR2_X1 U35 ( .A1(n931), .A2(n930), .ZN(n936) );
  AND2_X1 U35bar ( .A1(n931bar), .A2(n930bar), .ZN(n936bar);
  OR2_X1 U36 ( .A1(in_18), .A2(in[93]), .ZN(n930) );
  AND2_X1 U36bar ( .A1(in_18bar), .A2(inbar[93]), .ZN(n930bar);
  OR2_X1 U37 ( .A1(in_31), .A2(n929), .ZN(n931) );
  AND2_X1 U37bar ( .A1(in_31bar), .A2(n929bar), .ZN(n931bar);
  OR2_X1 U38 ( .A1(in_7), .A2(in_39), .ZN(n929) );
  AND2_X1 U38bar ( .A1(in_7bar), .A2(in_39bar), .ZN(n929bar);
  OR2_X1 U39 ( .A1(n928), .A2(n927), .ZN(out[5]) );
  AND2_X1 U39bar ( .A1(n928bar), .A2(n927bar), .ZN(outbar[5]);
  OR2_X1 U40 ( .A1(n926), .A2(n925), .ZN(n927) );
  AND2_X1 U40bar ( .A1(n926bar), .A2(n925bar), .ZN(n927bar);
  OR2_X1 U41 ( .A1(n924), .A2(n923), .ZN(n925) );
  AND2_X1 U41bar ( .A1(n924bar), .A2(n923bar), .ZN(n925bar);
  OR2_X1 U42 ( .A1(n922), .A2(n921), .ZN(n923) );
  AND2_X1 U42bar ( .A1(n922bar), .A2(n921bar), .ZN(n923bar);
  OR2_X1 U43 ( .A1(n940), .A2(n920), .ZN(n924) );
  AND2_X1 U43bar ( .A1(n940bar), .A2(n920bar), .ZN(n924bar);
  OR2_X1 U44 ( .A1(in[111]), .A2(n919), .ZN(n920) );
  AND2_X1 U44bar ( .A1(inbar[111]), .A2(n919bar), .ZN(n920bar);
  OR2_X1 U45 ( .A1(n918), .A2(n917), .ZN(n940) );
  AND2_X1 U45bar ( .A1(n918bar), .A2(n917bar), .ZN(n940bar);
  OR2_X1 U46 ( .A1(n916), .A2(n915), .ZN(n917) );
  AND2_X1 U46bar ( .A1(n916bar), .A2(n915bar), .ZN(n917bar);
  OR2_X1 U47 ( .A1(n914), .A2(n913), .ZN(n915) );
  AND2_X1 U47bar ( .A1(n914bar), .A2(n913bar), .ZN(n915bar);
  OR2_X1 U48 ( .A1(in[140]), .A2(in[131]), .ZN(n913) );
  AND2_X1 U48bar ( .A1(inbar[140]), .A2(inbar[131]), .ZN(n913bar);
  OR2_X1 U49 ( .A1(in[160]), .A2(in[144]), .ZN(n914) );
  AND2_X1 U49bar ( .A1(inbar[160]), .A2(inbar[144]), .ZN(n914bar);
  OR2_X1 U50 ( .A1(n912), .A2(n911), .ZN(n916) );
  AND2_X1 U50bar ( .A1(n912bar), .A2(n911bar), .ZN(n916bar);
  OR2_X1 U51 ( .A1(in[179]), .A2(in[174]), .ZN(n911) );
  AND2_X1 U51bar ( .A1(inbar[179]), .A2(inbar[174]), .ZN(n911bar);
  OR2_X1 U52 ( .A1(in[188]), .A2(in[184]), .ZN(n912) );
  AND2_X1 U52bar ( .A1(inbar[188]), .A2(inbar[184]), .ZN(n912bar);
  OR2_X1 U53 ( .A1(n910), .A2(n909), .ZN(n918) );
  AND2_X1 U53bar ( .A1(n910bar), .A2(n909bar), .ZN(n918bar);
  OR2_X1 U54 ( .A1(n908), .A2(n907), .ZN(n909) );
  AND2_X1 U54bar ( .A1(n908bar), .A2(n907bar), .ZN(n909bar);
  OR2_X1 U55 ( .A1(in[216]), .A2(in[200]), .ZN(n907) );
  AND2_X1 U55bar ( .A1(inbar[216]), .A2(inbar[200]), .ZN(n907bar);
  OR2_X1 U56 ( .A1(in[228]), .A2(in[224]), .ZN(n908) );
  AND2_X1 U56bar ( .A1(inbar[228]), .A2(inbar[224]), .ZN(n908bar);
  OR2_X1 U57 ( .A1(n906), .A2(n905), .ZN(n910) );
  AND2_X1 U57bar ( .A1(n906bar), .A2(n905bar), .ZN(n910bar);
  OR2_X1 U58 ( .A1(in[247]), .A2(in[235]), .ZN(n905) );
  AND2_X1 U58bar ( .A1(inbar[247]), .A2(inbar[235]), .ZN(n905bar);
  OR2_X1 U59 ( .A1(in_42), .A2(in[83]), .ZN(n906) );
  AND2_X1 U59bar ( .A1(in_42bar), .A2(inbar[83]), .ZN(n906bar);
  OR2_X1 U60 ( .A1(n904), .A2(n903), .ZN(n926) );
  AND2_X1 U60bar ( .A1(n904bar), .A2(n903bar), .ZN(n926bar);
  OR2_X1 U61 ( .A1(in[166]), .A2(in[123]), .ZN(n903) );
  AND2_X1 U61bar ( .A1(inbar[166]), .A2(inbar[123]), .ZN(n903bar);
  OR2_X1 U62 ( .A1(in[170]), .A2(n902), .ZN(n904) );
  AND2_X1 U62bar ( .A1(inbar[170]), .A2(n902bar), .ZN(n904bar);
  OR2_X1 U63 ( .A1(in[194]), .A2(in[183]), .ZN(n902) );
  AND2_X1 U63bar ( .A1(inbar[194]), .A2(inbar[183]), .ZN(n902bar);
  OR2_X1 U64 ( .A1(n901), .A2(n900), .ZN(n928) );
  AND2_X1 U64bar ( .A1(n901bar), .A2(n900bar), .ZN(n928bar);
  OR2_X1 U65 ( .A1(n899), .A2(n898), .ZN(n900) );
  AND2_X1 U65bar ( .A1(n899bar), .A2(n898bar), .ZN(n900bar);
  OR2_X1 U66 ( .A1(in[241]), .A2(in[238]), .ZN(n898) );
  AND2_X1 U66bar ( .A1(inbar[241]), .A2(inbar[238]), .ZN(n898bar);
  OR2_X1 U67 ( .A1(in[250]), .A2(n897), .ZN(n899) );
  AND2_X1 U67bar ( .A1(inbar[250]), .A2(n897bar), .ZN(n899bar);
  OR2_X1 U68 ( .A1(in_24), .A2(in[84]), .ZN(n897) );
  AND2_X1 U68bar ( .A1(in_24bar), .A2(inbar[84]), .ZN(n897bar);
  OR2_X1 U69 ( .A1(n896), .A2(n895), .ZN(n901) );
  AND2_X1 U69bar ( .A1(n896bar), .A2(n895bar), .ZN(n901bar);
  OR2_X1 U70 ( .A1(in_41), .A2(in_29), .ZN(n895) );
  AND2_X1 U70bar ( .A1(in_41bar), .A2(in_29bar), .ZN(n895bar);
  OR2_X1 U71 ( .A1(in_66), .A2(n894), .ZN(n896) );
  AND2_X1 U71bar ( .A1(in_66bar), .A2(n894bar), .ZN(n896bar);
  OR2_X1 U72 ( .A1(in_76), .A2(in_71), .ZN(n894) );
  AND2_X1 U72bar ( .A1(in_76bar), .A2(in_71bar), .ZN(n894bar);
  OR2_X1 U73 ( .A1(n893), .A2(n892), .ZN(out[4]) );
  AND2_X1 U73bar ( .A1(n893bar), .A2(n892bar), .ZN(outbar[4]);
  OR2_X1 U74 ( .A1(n891), .A2(n890), .ZN(n892) );
  AND2_X1 U74bar ( .A1(n891bar), .A2(n890bar), .ZN(n892bar);
  OR2_X1 U75 ( .A1(n889), .A2(n888), .ZN(n890) );
  AND2_X1 U75bar ( .A1(n889bar), .A2(n888bar), .ZN(n890bar);
  OR2_X1 U76 ( .A1(n922), .A2(n887), .ZN(n888) );
  AND2_X1 U76bar ( .A1(n922bar), .A2(n887bar), .ZN(n888bar);
  OR2_X1 U77 ( .A1(n886), .A2(n885), .ZN(n922) );
  AND2_X1 U77bar ( .A1(n886bar), .A2(n885bar), .ZN(n922bar);
  OR2_X1 U78 ( .A1(n884), .A2(n883), .ZN(n885) );
  AND2_X1 U78bar ( .A1(n884bar), .A2(n883bar), .ZN(n885bar);
  OR2_X1 U79 ( .A1(n882), .A2(n881), .ZN(n883) );
  AND2_X1 U79bar ( .A1(n882bar), .A2(n881bar), .ZN(n883bar);
  OR2_X1 U80 ( .A1(in[118]), .A2(in[109]), .ZN(n881) );
  AND2_X1 U80bar ( .A1(inbar[118]), .A2(inbar[109]), .ZN(n881bar);
  OR2_X1 U81 ( .A1(in[139]), .A2(in[120]), .ZN(n882) );
  AND2_X1 U81bar ( .A1(inbar[139]), .A2(inbar[120]), .ZN(n882bar);
  OR2_X1 U82 ( .A1(n880), .A2(n879), .ZN(n884) );
  AND2_X1 U82bar ( .A1(n880bar), .A2(n879bar), .ZN(n884bar);
  OR2_X1 U83 ( .A1(in[198]), .A2(in[154]), .ZN(n879) );
  AND2_X1 U83bar ( .A1(inbar[198]), .A2(inbar[154]), .ZN(n879bar);
  OR2_X1 U84 ( .A1(in[210]), .A2(in[205]), .ZN(n880) );
  AND2_X1 U84bar ( .A1(inbar[210]), .A2(inbar[205]), .ZN(n880bar);
  OR2_X1 U85 ( .A1(n878), .A2(n877), .ZN(n886) );
  AND2_X1 U85bar ( .A1(n878bar), .A2(n877bar), .ZN(n886bar);
  OR2_X1 U86 ( .A1(n876), .A2(n875), .ZN(n877) );
  AND2_X1 U86bar ( .A1(n876bar), .A2(n875bar), .ZN(n877bar);
  OR2_X1 U87 ( .A1(in[219]), .A2(in[217]), .ZN(n875) );
  AND2_X1 U87bar ( .A1(inbar[219]), .A2(inbar[217]), .ZN(n875bar);
  OR2_X1 U88 ( .A1(in[86]), .A2(in[252]), .ZN(n876) );
  AND2_X1 U88bar ( .A1(inbar[86]), .A2(inbar[252]), .ZN(n876bar);
  OR2_X1 U89 ( .A1(n874), .A2(n873), .ZN(n878) );
  AND2_X1 U89bar ( .A1(n874bar), .A2(n873bar), .ZN(n878bar);
  OR2_X1 U90 ( .A1(in_40), .A2(in[91]), .ZN(n873) );
  AND2_X1 U90bar ( .A1(in_40bar), .A2(inbar[91]), .ZN(n873bar);
  OR2_X1 U91 ( .A1(in_8), .A2(in_46), .ZN(n874) );
  AND2_X1 U91bar ( .A1(in_8bar), .A2(in_46bar), .ZN(n874bar);
  OR2_X1 U92 ( .A1(n872), .A2(n871), .ZN(n889) );
  AND2_X1 U92bar ( .A1(n872bar), .A2(n871bar), .ZN(n889bar);
  OR2_X1 U93 ( .A1(in[117]), .A2(n943), .ZN(n871) );
  AND2_X1 U93bar ( .A1(inbar[117]), .A2(n943bar), .ZN(n871bar);
  OR2_X1 U94 ( .A1(n870), .A2(n869), .ZN(n943) );
  AND2_X1 U94bar ( .A1(n870bar), .A2(n869bar), .ZN(n943bar);
  OR2_X1 U95 ( .A1(n868), .A2(n867), .ZN(n869) );
  AND2_X1 U95bar ( .A1(n868bar), .A2(n867bar), .ZN(n869bar);
  OR2_X1 U96 ( .A1(n866), .A2(n865), .ZN(n867) );
  AND2_X1 U96bar ( .A1(n866bar), .A2(n865bar), .ZN(n867bar);
  OR2_X1 U97 ( .A1(n864), .A2(n863), .ZN(n865) );
  AND2_X1 U97bar ( .A1(n864bar), .A2(n863bar), .ZN(n865bar);
  OR2_X1 U98 ( .A1(in[108]), .A2(n919), .ZN(n866) );
  AND2_X1 U98bar ( .A1(inbar[108]), .A2(n919bar), .ZN(n866bar);
  OR2_X1 U99 ( .A1(n862), .A2(n861), .ZN(n919) );
  AND2_X1 U99bar ( .A1(n862bar), .A2(n861bar), .ZN(n919bar);
  OR2_X1 U100 ( .A1(n860), .A2(n859), .ZN(n861) );
  AND2_X1 U100bar ( .A1(n860bar), .A2(n859bar), .ZN(n861bar);
  OR2_X1 U101 ( .A1(n858), .A2(n857), .ZN(n859) );
  AND2_X1 U101bar ( .A1(n858bar), .A2(n857bar), .ZN(n859bar);
  OR2_X1 U102 ( .A1(in[119]), .A2(in[105]), .ZN(n857) );
  AND2_X1 U102bar ( .A1(inbar[119]), .A2(inbar[105]), .ZN(n857bar);
  OR2_X1 U103 ( .A1(in[186]), .A2(in[175]), .ZN(n858) );
  AND2_X1 U103bar ( .A1(inbar[186]), .A2(inbar[175]), .ZN(n858bar);
  OR2_X1 U104 ( .A1(n856), .A2(n855), .ZN(n860) );
  AND2_X1 U104bar ( .A1(n856bar), .A2(n855bar), .ZN(n860bar);
  OR2_X1 U105 ( .A1(in[202]), .A2(in[193]), .ZN(n855) );
  AND2_X1 U105bar ( .A1(inbar[202]), .A2(inbar[193]), .ZN(n855bar);
  OR2_X1 U106 ( .A1(in[225]), .A2(in[208]), .ZN(n856) );
  AND2_X1 U106bar ( .A1(inbar[225]), .A2(inbar[208]), .ZN(n856bar);
  OR2_X1 U107 ( .A1(n854), .A2(n853), .ZN(n862) );
  AND2_X1 U107bar ( .A1(n854bar), .A2(n853bar), .ZN(n862bar);
  OR2_X1 U108 ( .A1(n852), .A2(n851), .ZN(n853) );
  AND2_X1 U108bar ( .A1(n852bar), .A2(n851bar), .ZN(n853bar);
  OR2_X1 U109 ( .A1(in_1), .A2(in[85]), .ZN(n851) );
  AND2_X1 U109bar ( .A1(in_1bar), .A2(inbar[85]), .ZN(n851bar);
  OR2_X1 U110 ( .A1(in_23), .A2(in_19), .ZN(n852) );
  AND2_X1 U110bar ( .A1(in_23bar), .A2(in_19bar), .ZN(n852bar);
  OR2_X1 U111 ( .A1(n850), .A2(n849), .ZN(n854) );
  AND2_X1 U111bar ( .A1(n850bar), .A2(n849bar), .ZN(n854bar);
  OR2_X1 U112 ( .A1(in_43), .A2(in_33), .ZN(n849) );
  AND2_X1 U112bar ( .A1(in_43bar), .A2(in_33bar), .ZN(n849bar);
  OR2_X1 U113 ( .A1(in_63), .A2(in_44), .ZN(n850) );
  AND2_X1 U113bar ( .A1(in_63bar), .A2(in_44bar), .ZN(n850bar);
  OR2_X1 U114 ( .A1(n848), .A2(n847), .ZN(n868) );
  AND2_X1 U114bar ( .A1(n848bar), .A2(n847bar), .ZN(n868bar);
  OR2_X1 U115 ( .A1(in[141]), .A2(in[112]), .ZN(n847) );
  AND2_X1 U115bar ( .A1(inbar[141]), .A2(inbar[112]), .ZN(n847bar);
  OR2_X1 U116 ( .A1(in[147]), .A2(n846), .ZN(n848) );
  AND2_X1 U116bar ( .A1(inbar[147]), .A2(n846bar), .ZN(n848bar);
  OR2_X1 U117 ( .A1(in[181]), .A2(in[167]), .ZN(n846) );
  AND2_X1 U117bar ( .A1(inbar[181]), .A2(inbar[167]), .ZN(n846bar);
  OR2_X1 U118 ( .A1(n845), .A2(n844), .ZN(n870) );
  AND2_X1 U118bar ( .A1(n845bar), .A2(n844bar), .ZN(n870bar);
  OR2_X1 U119 ( .A1(n843), .A2(n842), .ZN(n844) );
  AND2_X1 U119bar ( .A1(n843bar), .A2(n842bar), .ZN(n844bar);
  OR2_X1 U120 ( .A1(in[229]), .A2(in[201]), .ZN(n842) );
  AND2_X1 U120bar ( .A1(inbar[229]), .A2(inbar[201]), .ZN(n842bar);
  OR2_X1 U121 ( .A1(in[237]), .A2(n841), .ZN(n843) );
  AND2_X1 U121bar ( .A1(inbar[237]), .A2(n841bar), .ZN(n843bar);
  OR2_X1 U122 ( .A1(in[94]), .A2(in[253]), .ZN(n841) );
  AND2_X1 U122bar ( .A1(inbar[94]), .A2(inbar[253]), .ZN(n841bar);
  OR2_X1 U123 ( .A1(n840), .A2(n839), .ZN(n845) );
  AND2_X1 U123bar ( .A1(n840bar), .A2(n839bar), .ZN(n845bar);
  OR2_X1 U124 ( .A1(in_21), .A2(in[96]), .ZN(n839) );
  AND2_X1 U124bar ( .A1(in_21bar), .A2(inbar[96]), .ZN(n839bar);
  OR2_X1 U125 ( .A1(in_25), .A2(n838), .ZN(n840) );
  AND2_X1 U125bar ( .A1(in_25bar), .A2(n838bar), .ZN(n840bar);
  OR2_X1 U126 ( .A1(in_81), .A2(in_45), .ZN(n838) );
  AND2_X1 U126bar ( .A1(in_81bar), .A2(in_45bar), .ZN(n838bar);
  OR2_X1 U127 ( .A1(n837), .A2(n836), .ZN(n891) );
  AND2_X1 U127bar ( .A1(n837bar), .A2(n836bar), .ZN(n891bar);
  OR2_X1 U128 ( .A1(in[142]), .A2(in[124]), .ZN(n836) );
  AND2_X1 U128bar ( .A1(inbar[142]), .A2(inbar[124]), .ZN(n836bar);
  OR2_X1 U129 ( .A1(in[150]), .A2(n835), .ZN(n837) );
  AND2_X1 U129bar ( .A1(inbar[150]), .A2(n835bar), .ZN(n837bar);
  OR2_X1 U130 ( .A1(in[172]), .A2(in[155]), .ZN(n835) );
  AND2_X1 U130bar ( .A1(inbar[172]), .A2(inbar[155]), .ZN(n835bar);
  OR2_X1 U131 ( .A1(n834), .A2(n833), .ZN(n893) );
  AND2_X1 U131bar ( .A1(n834bar), .A2(n833bar), .ZN(n893bar);
  OR2_X1 U132 ( .A1(n832), .A2(n831), .ZN(n833) );
  AND2_X1 U132bar ( .A1(n832bar), .A2(n831bar), .ZN(n833bar);
  OR2_X1 U133 ( .A1(in[196]), .A2(in[173]), .ZN(n831) );
  AND2_X1 U133bar ( .A1(inbar[196]), .A2(inbar[173]), .ZN(n831bar);
  OR2_X1 U134 ( .A1(in[222]), .A2(n830), .ZN(n832) );
  AND2_X1 U134bar ( .A1(inbar[222]), .A2(n830bar), .ZN(n832bar);
  OR2_X1 U135 ( .A1(in[227]), .A2(in[226]), .ZN(n830) );
  AND2_X1 U135bar ( .A1(inbar[227]), .A2(inbar[226]), .ZN(n830bar);
  OR2_X1 U136 ( .A1(n829), .A2(n828), .ZN(n834) );
  AND2_X1 U136bar ( .A1(n829bar), .A2(n828bar), .ZN(n834bar);
  OR2_X1 U137 ( .A1(in[249]), .A2(in[231]), .ZN(n828) );
  AND2_X1 U137bar ( .A1(inbar[249]), .A2(inbar[231]), .ZN(n828bar);
  OR2_X1 U138 ( .A1(in_28), .A2(n827), .ZN(n829) );
  AND2_X1 U138bar ( .A1(in_28bar), .A2(n827bar), .ZN(n829bar);
  OR2_X1 U139 ( .A1(in_52), .A2(in_47), .ZN(n827) );
  AND2_X1 U139bar ( .A1(in_52bar), .A2(in_47bar), .ZN(n827bar);
  OR2_X1 U140 ( .A1(n826), .A2(n825), .ZN(out[3]) );
  AND2_X1 U140bar ( .A1(n826bar), .A2(n825bar), .ZN(outbar[3]);
  OR2_X1 U141 ( .A1(n824), .A2(n823), .ZN(n825) );
  AND2_X1 U141bar ( .A1(n824bar), .A2(n823bar), .ZN(n825bar);
  OR2_X1 U142 ( .A1(n822), .A2(n821), .ZN(n823) );
  AND2_X1 U142bar ( .A1(n822bar), .A2(n821bar), .ZN(n823bar);
  OR2_X1 U143 ( .A1(n820), .A2(n819), .ZN(n821) );
  AND2_X1 U143bar ( .A1(n820bar), .A2(n819bar), .ZN(n821bar);
  OR2_X1 U144 ( .A1(n964), .A2(n818), .ZN(n822) );
  AND2_X1 U144bar ( .A1(n964bar), .A2(n818bar), .ZN(n822bar);
  OR2_X1 U145 ( .A1(in[118]), .A2(n817), .ZN(n818) );
  AND2_X1 U145bar ( .A1(inbar[118]), .A2(n817bar), .ZN(n818bar);
  OR2_X1 U146 ( .A1(n816), .A2(n815), .ZN(n964) );
  AND2_X1 U146bar ( .A1(n816bar), .A2(n815bar), .ZN(n964bar);
  OR2_X1 U147 ( .A1(n814), .A2(n813), .ZN(n815) );
  AND2_X1 U147bar ( .A1(n814bar), .A2(n813bar), .ZN(n815bar);
  OR2_X1 U148 ( .A1(n812), .A2(n811), .ZN(n813) );
  AND2_X1 U148bar ( .A1(n812bar), .A2(n811bar), .ZN(n813bar);
  OR2_X1 U149 ( .A1(in[122]), .A2(in[111]), .ZN(n811) );
  AND2_X1 U149bar ( .A1(inbar[122]), .A2(inbar[111]), .ZN(n811bar);
  OR2_X1 U150 ( .A1(in[154]), .A2(in[151]), .ZN(n812) );
  AND2_X1 U150bar ( .A1(inbar[154]), .A2(inbar[151]), .ZN(n812bar);
  OR2_X1 U151 ( .A1(n810), .A2(n809), .ZN(n814) );
  AND2_X1 U151bar ( .A1(n810bar), .A2(n809bar), .ZN(n814bar);
  OR2_X1 U152 ( .A1(in[187]), .A2(in[177]), .ZN(n809) );
  AND2_X1 U152bar ( .A1(inbar[187]), .A2(inbar[177]), .ZN(n809bar);
  OR2_X1 U153 ( .A1(in[200]), .A2(in[192]), .ZN(n810) );
  AND2_X1 U153bar ( .A1(inbar[200]), .A2(inbar[192]), .ZN(n810bar);
  OR2_X1 U154 ( .A1(n808), .A2(n807), .ZN(n816) );
  AND2_X1 U154bar ( .A1(n808bar), .A2(n807bar), .ZN(n816bar);
  OR2_X1 U155 ( .A1(n806), .A2(n805), .ZN(n807) );
  AND2_X1 U155bar ( .A1(n806bar), .A2(n805bar), .ZN(n807bar);
  OR2_X1 U156 ( .A1(in[225]), .A2(in[207]), .ZN(n805) );
  AND2_X1 U156bar ( .A1(inbar[225]), .A2(inbar[207]), .ZN(n805bar);
  OR2_X1 U157 ( .A1(in[98]), .A2(in[226]), .ZN(n806) );
  AND2_X1 U157bar ( .A1(inbar[98]), .A2(inbar[226]), .ZN(n806bar);
  OR2_X1 U158 ( .A1(n804), .A2(n803), .ZN(n808) );
  AND2_X1 U158bar ( .A1(n804bar), .A2(n803bar), .ZN(n808bar);
  OR2_X1 U159 ( .A1(in_20), .A2(in_16), .ZN(n803) );
  AND2_X1 U159bar ( .A1(in_20bar), .A2(in_16bar), .ZN(n803bar);
  OR2_X1 U160 ( .A1(in_55), .A2(in_45), .ZN(n804) );
  AND2_X1 U160bar ( .A1(in_55bar), .A2(in_45bar), .ZN(n804bar);
  OR2_X1 U161 ( .A1(n802), .A2(n801), .ZN(n824) );
  AND2_X1 U161bar ( .A1(n802bar), .A2(n801bar), .ZN(n824bar);
  OR2_X1 U162 ( .A1(in[162]), .A2(in[149]), .ZN(n801) );
  AND2_X1 U162bar ( .A1(inbar[162]), .A2(inbar[149]), .ZN(n801bar);
  OR2_X1 U163 ( .A1(in[163]), .A2(n800), .ZN(n802) );
  AND2_X1 U163bar ( .A1(inbar[163]), .A2(n800bar), .ZN(n802bar);
  OR2_X1 U164 ( .A1(in[191]), .A2(in[189]), .ZN(n800) );
  AND2_X1 U164bar ( .A1(inbar[191]), .A2(inbar[189]), .ZN(n800bar);
  OR2_X1 U165 ( .A1(n799), .A2(n798), .ZN(n826) );
  AND2_X1 U165bar ( .A1(n799bar), .A2(n798bar), .ZN(n826bar);
  OR2_X1 U166 ( .A1(n797), .A2(n796), .ZN(n798) );
  AND2_X1 U166bar ( .A1(n797bar), .A2(n796bar), .ZN(n798bar);
  OR2_X1 U167 ( .A1(in[212]), .A2(in[193]), .ZN(n796) );
  AND2_X1 U167bar ( .A1(inbar[212]), .A2(inbar[193]), .ZN(n796bar);
  OR2_X1 U168 ( .A1(in[238]), .A2(n795), .ZN(n797) );
  AND2_X1 U168bar ( .A1(inbar[238]), .A2(n795bar), .ZN(n797bar);
  OR2_X1 U169 ( .A1(in[88]), .A2(in[247]), .ZN(n795) );
  AND2_X1 U169bar ( .A1(inbar[88]), .A2(inbar[247]), .ZN(n795bar);
  OR2_X1 U170 ( .A1(n794), .A2(n793), .ZN(n799) );
  AND2_X1 U170bar ( .A1(n794bar), .A2(n793bar), .ZN(n799bar);
  OR2_X1 U171 ( .A1(in[94]), .A2(in[92]), .ZN(n793) );
  AND2_X1 U171bar ( .A1(inbar[94]), .A2(inbar[92]), .ZN(n793bar);
  OR2_X1 U172 ( .A1(in_52), .A2(n792), .ZN(n794) );
  AND2_X1 U172bar ( .A1(in_52bar), .A2(n792bar), .ZN(n794bar);
  OR2_X1 U173 ( .A1(in_70), .A2(in_67), .ZN(n792) );
  AND2_X1 U173bar ( .A1(in_70bar), .A2(in_67bar), .ZN(n792bar);
  OR2_X1 U174 ( .A1(n791), .A2(n790), .ZN(out[2]) );
  AND2_X1 U174bar ( .A1(n791bar), .A2(n790bar), .ZN(outbar[2]);
  OR2_X1 U175 ( .A1(n789), .A2(n788), .ZN(n790) );
  AND2_X1 U175bar ( .A1(n789bar), .A2(n788bar), .ZN(n790bar);
  OR2_X1 U176 ( .A1(n787), .A2(n786), .ZN(n788) );
  AND2_X1 U176bar ( .A1(n787bar), .A2(n786bar), .ZN(n788bar);
  OR2_X1 U177 ( .A1(n819), .A2(n785), .ZN(n786) );
  AND2_X1 U177bar ( .A1(n819bar), .A2(n785bar), .ZN(n786bar);
  OR2_X1 U178 ( .A1(n784), .A2(n783), .ZN(n819) );
  AND2_X1 U178bar ( .A1(n784bar), .A2(n783bar), .ZN(n819bar);
  OR2_X1 U179 ( .A1(n782), .A2(n781), .ZN(n783) );
  AND2_X1 U179bar ( .A1(n782bar), .A2(n781bar), .ZN(n783bar);
  OR2_X1 U180 ( .A1(n780), .A2(n779), .ZN(n781) );
  AND2_X1 U180bar ( .A1(n780bar), .A2(n779bar), .ZN(n781bar);
  OR2_X1 U181 ( .A1(n962), .A2(n778), .ZN(n779) );
  AND2_X1 U181bar ( .A1(n962bar), .A2(n778bar), .ZN(n779bar);
  OR2_X1 U182 ( .A1(n777), .A2(n776), .ZN(n962) );
  AND2_X1 U182bar ( .A1(n777bar), .A2(n776bar), .ZN(n962bar);
  OR2_X1 U183 ( .A1(n775), .A2(n774), .ZN(n776) );
  AND2_X1 U183bar ( .A1(n775bar), .A2(n774bar), .ZN(n776bar);
  OR2_X1 U184 ( .A1(n773), .A2(n772), .ZN(n774) );
  AND2_X1 U184bar ( .A1(n773bar), .A2(n772bar), .ZN(n774bar);
  OR2_X1 U185 ( .A1(in[131]), .A2(in[120]), .ZN(n772) );
  AND2_X1 U185bar ( .A1(inbar[131]), .A2(inbar[120]), .ZN(n772bar);
  OR2_X1 U186 ( .A1(in[153]), .A2(in[147]), .ZN(n773) );
  AND2_X1 U186bar ( .A1(inbar[153]), .A2(inbar[147]), .ZN(n773bar);
  OR2_X1 U187 ( .A1(n771), .A2(n770), .ZN(n775) );
  AND2_X1 U187bar ( .A1(n771bar), .A2(n770bar), .ZN(n775bar);
  OR2_X1 U188 ( .A1(in[170]), .A2(in[156]), .ZN(n770) );
  AND2_X1 U188bar ( .A1(inbar[170]), .A2(inbar[156]), .ZN(n770bar);
  OR2_X1 U189 ( .A1(in[223]), .A2(in[190]), .ZN(n771) );
  AND2_X1 U189bar ( .A1(inbar[223]), .A2(inbar[190]), .ZN(n771bar);
  OR2_X1 U190 ( .A1(n769), .A2(n768), .ZN(n777) );
  AND2_X1 U190bar ( .A1(n769bar), .A2(n768bar), .ZN(n777bar);
  OR2_X1 U191 ( .A1(n767), .A2(n766), .ZN(n768) );
  AND2_X1 U191bar ( .A1(n767bar), .A2(n766bar), .ZN(n768bar);
  OR2_X1 U192 ( .A1(in[236]), .A2(in[230]), .ZN(n766) );
  AND2_X1 U192bar ( .A1(inbar[236]), .A2(inbar[230]), .ZN(n766bar);
  OR2_X1 U193 ( .A1(in[85]), .A2(in[240]), .ZN(n767) );
  AND2_X1 U193bar ( .A1(inbar[85]), .A2(inbar[240]), .ZN(n767bar);
  OR2_X1 U194 ( .A1(n765), .A2(n764), .ZN(n769) );
  AND2_X1 U194bar ( .A1(n765bar), .A2(n764bar), .ZN(n769bar);
  OR2_X1 U195 ( .A1(in_12), .A2(in[90]), .ZN(n764) );
  AND2_X1 U195bar ( .A1(in_12bar), .A2(inbar[90]), .ZN(n764bar);
  OR2_X1 U196 ( .A1(in_39), .A2(in_28), .ZN(n765) );
  AND2_X1 U196bar ( .A1(in_39bar), .A2(in_28bar), .ZN(n765bar);
  OR2_X1 U197 ( .A1(in[109]), .A2(n763), .ZN(n780) );
  AND2_X1 U197bar ( .A1(inbar[109]), .A2(n763bar), .ZN(n780bar);
  OR2_X1 U198 ( .A1(n762), .A2(n761), .ZN(n782) );
  AND2_X1 U198bar ( .A1(n762bar), .A2(n761bar), .ZN(n782bar);
  OR2_X1 U199 ( .A1(in[138]), .A2(in[129]), .ZN(n761) );
  AND2_X1 U199bar ( .A1(inbar[138]), .A2(inbar[129]), .ZN(n761bar);
  OR2_X1 U200 ( .A1(in[157]), .A2(n760), .ZN(n762) );
  AND2_X1 U200bar ( .A1(inbar[157]), .A2(n760bar), .ZN(n762bar);
  OR2_X1 U201 ( .A1(in[182]), .A2(in[167]), .ZN(n760) );
  AND2_X1 U201bar ( .A1(inbar[182]), .A2(inbar[167]), .ZN(n760bar);
  OR2_X1 U202 ( .A1(n759), .A2(n758), .ZN(n784) );
  AND2_X1 U202bar ( .A1(n759bar), .A2(n758bar), .ZN(n784bar);
  OR2_X1 U203 ( .A1(n757), .A2(n756), .ZN(n758) );
  AND2_X1 U203bar ( .A1(n757bar), .A2(n756bar), .ZN(n758bar);
  OR2_X1 U204 ( .A1(in[195]), .A2(in[184]), .ZN(n756) );
  AND2_X1 U204bar ( .A1(inbar[195]), .A2(inbar[184]), .ZN(n756bar);
  OR2_X1 U205 ( .A1(in[196]), .A2(n755), .ZN(n757) );
  AND2_X1 U205bar ( .A1(inbar[196]), .A2(n755bar), .ZN(n757bar);
  OR2_X1 U206 ( .A1(in[215]), .A2(in[209]), .ZN(n755) );
  AND2_X1 U206bar ( .A1(inbar[215]), .A2(inbar[209]), .ZN(n755bar);
  OR2_X1 U207 ( .A1(n754), .A2(n753), .ZN(n759) );
  AND2_X1 U207bar ( .A1(n754bar), .A2(n753bar), .ZN(n759bar);
  OR2_X1 U208 ( .A1(in[93]), .A2(in[233]), .ZN(n753) );
  AND2_X1 U208bar ( .A1(inbar[93]), .A2(inbar[233]), .ZN(n753bar);
  OR2_X1 U209 ( .A1(in_1), .A2(n752), .ZN(n754) );
  AND2_X1 U209bar ( .A1(in_1bar), .A2(n752bar), .ZN(n754bar);
  OR2_X1 U210 ( .A1(in_69), .A2(in_66), .ZN(n752) );
  AND2_X1 U210bar ( .A1(in_69bar), .A2(in_66bar), .ZN(n752bar);
  OR2_X1 U211 ( .A1(n966), .A2(n751), .ZN(n787) );
  AND2_X1 U211bar ( .A1(n966bar), .A2(n751bar), .ZN(n787bar);
  OR2_X1 U212 ( .A1(in[134]), .A2(n750), .ZN(n751) );
  AND2_X1 U212bar ( .A1(inbar[134]), .A2(n750bar), .ZN(n751bar);
  OR2_X1 U213 ( .A1(n749), .A2(n748), .ZN(n966) );
  AND2_X1 U213bar ( .A1(n749bar), .A2(n748bar), .ZN(n966bar);
  OR2_X1 U214 ( .A1(n747), .A2(n746), .ZN(n748) );
  AND2_X1 U214bar ( .A1(n747bar), .A2(n746bar), .ZN(n748bar);
  OR2_X1 U215 ( .A1(n745), .A2(n744), .ZN(n746) );
  AND2_X1 U215bar ( .A1(n745bar), .A2(n744bar), .ZN(n746bar);
  OR2_X1 U216 ( .A1(in[136]), .A2(in[121]), .ZN(n744) );
  AND2_X1 U216bar ( .A1(inbar[136]), .A2(inbar[121]), .ZN(n744bar);
  OR2_X1 U217 ( .A1(in[186]), .A2(in[174]), .ZN(n745) );
  AND2_X1 U217bar ( .A1(inbar[186]), .A2(inbar[174]), .ZN(n745bar);
  OR2_X1 U218 ( .A1(n743), .A2(n742), .ZN(n747) );
  AND2_X1 U218bar ( .A1(n743bar), .A2(n742bar), .ZN(n747bar);
  OR2_X1 U219 ( .A1(in[198]), .A2(in[197]), .ZN(n742) );
  AND2_X1 U219bar ( .A1(inbar[198]), .A2(inbar[197]), .ZN(n742bar);
  OR2_X1 U220 ( .A1(in[214]), .A2(in[199]), .ZN(n743) );
  AND2_X1 U220bar ( .A1(inbar[214]), .A2(inbar[199]), .ZN(n743bar);
  OR2_X1 U221 ( .A1(n741), .A2(n740), .ZN(n749) );
  AND2_X1 U221bar ( .A1(n741bar), .A2(n740bar), .ZN(n749bar);
  OR2_X1 U222 ( .A1(n739), .A2(n738), .ZN(n740) );
  AND2_X1 U222bar ( .A1(n739bar), .A2(n738bar), .ZN(n740bar);
  OR2_X1 U223 ( .A1(in[231]), .A2(in[220]), .ZN(n738) );
  AND2_X1 U223bar ( .A1(inbar[231]), .A2(inbar[220]), .ZN(n738bar);
  OR2_X1 U224 ( .A1(in_25), .A2(in[245]), .ZN(n739) );
  AND2_X1 U224bar ( .A1(in_25bar), .A2(inbar[245]), .ZN(n739bar);
  OR2_X1 U225 ( .A1(n737), .A2(n736), .ZN(n741) );
  AND2_X1 U225bar ( .A1(n737bar), .A2(n736bar), .ZN(n741bar);
  OR2_X1 U226 ( .A1(in_53), .A2(in_29), .ZN(n736) );
  AND2_X1 U226bar ( .A1(in_53bar), .A2(in_29bar), .ZN(n736bar);
  OR2_X1 U227 ( .A1(in_79), .A2(in_74), .ZN(n737) );
  AND2_X1 U227bar ( .A1(in_79bar), .A2(in_74bar), .ZN(n737bar);
  OR2_X1 U228 ( .A1(n735), .A2(n734), .ZN(n789) );
  AND2_X1 U228bar ( .A1(n735bar), .A2(n734bar), .ZN(n789bar);
  OR2_X1 U229 ( .A1(in[152]), .A2(in[140]), .ZN(n734) );
  AND2_X1 U229bar ( .A1(inbar[152]), .A2(inbar[140]), .ZN(n734bar);
  OR2_X1 U230 ( .A1(in[155]), .A2(n733), .ZN(n735) );
  AND2_X1 U230bar ( .A1(inbar[155]), .A2(n733bar), .ZN(n735bar);
  OR2_X1 U231 ( .A1(in[166]), .A2(in[165]), .ZN(n733) );
  AND2_X1 U231bar ( .A1(inbar[166]), .A2(inbar[165]), .ZN(n733bar);
  OR2_X1 U232 ( .A1(n732), .A2(n731), .ZN(n791) );
  AND2_X1 U232bar ( .A1(n732bar), .A2(n731bar), .ZN(n791bar);
  OR2_X1 U233 ( .A1(n730), .A2(n729), .ZN(n731) );
  AND2_X1 U233bar ( .A1(n730bar), .A2(n729bar), .ZN(n731bar);
  OR2_X1 U234 ( .A1(in[202]), .A2(in[185]), .ZN(n729) );
  AND2_X1 U234bar ( .A1(inbar[202]), .A2(inbar[185]), .ZN(n729bar);
  OR2_X1 U235 ( .A1(in[211]), .A2(n728), .ZN(n730) );
  AND2_X1 U235bar ( .A1(inbar[211]), .A2(n728bar), .ZN(n730bar);
  OR2_X1 U236 ( .A1(in[255]), .A2(in[253]), .ZN(n728) );
  AND2_X1 U236bar ( .A1(inbar[255]), .A2(inbar[253]), .ZN(n728bar);
  OR2_X1 U237 ( .A1(n727), .A2(n726), .ZN(n732) );
  AND2_X1 U237bar ( .A1(n727bar), .A2(n726bar), .ZN(n732bar);
  OR2_X1 U238 ( .A1(in_35), .A2(in_15), .ZN(n726) );
  AND2_X1 U238bar ( .A1(in_35bar), .A2(in_15bar), .ZN(n726bar);
  OR2_X1 U239 ( .A1(in_36), .A2(n725), .ZN(n727) );
  AND2_X1 U239bar ( .A1(in_36bar), .A2(n725bar), .ZN(n727bar);
  OR2_X1 U240 ( .A1(in_48), .A2(in_40), .ZN(n725) );
  AND2_X1 U240bar ( .A1(in_48bar), .A2(in_40bar), .ZN(n725bar);
  OR2_X1 U241 ( .A1(n724), .A2(n723), .ZN(out[1]) );
  AND2_X1 U241bar ( .A1(n724bar), .A2(n723bar), .ZN(outbar[1]);
  OR2_X1 U242 ( .A1(n722), .A2(n721), .ZN(n723) );
  AND2_X1 U242bar ( .A1(n722bar), .A2(n721bar), .ZN(n723bar);
  OR2_X1 U243 ( .A1(n720), .A2(n719), .ZN(n721) );
  AND2_X1 U243bar ( .A1(n720bar), .A2(n719bar), .ZN(n721bar);
  OR2_X1 U244 ( .A1(n921), .A2(n887), .ZN(n719) );
  AND2_X1 U244bar ( .A1(n921bar), .A2(n887bar), .ZN(n719bar);
  OR2_X1 U245 ( .A1(n718), .A2(n717), .ZN(n887) );
  AND2_X1 U245bar ( .A1(n718bar), .A2(n717bar), .ZN(n887bar);
  OR2_X1 U246 ( .A1(n716), .A2(n715), .ZN(n717) );
  AND2_X1 U246bar ( .A1(n716bar), .A2(n715bar), .ZN(n717bar);
  OR2_X1 U247 ( .A1(n714), .A2(n713), .ZN(n715) );
  AND2_X1 U247bar ( .A1(n714bar), .A2(n713bar), .ZN(n715bar);
  OR2_X1 U248 ( .A1(in[116]), .A2(in[110]), .ZN(n713) );
  AND2_X1 U248bar ( .A1(inbar[116]), .A2(inbar[110]), .ZN(n713bar);
  OR2_X1 U249 ( .A1(in[133]), .A2(in[130]), .ZN(n714) );
  AND2_X1 U249bar ( .A1(inbar[133]), .A2(inbar[130]), .ZN(n714bar);
  OR2_X1 U250 ( .A1(n712), .A2(n711), .ZN(n716) );
  AND2_X1 U250bar ( .A1(n712bar), .A2(n711bar), .ZN(n716bar);
  OR2_X1 U251 ( .A1(in[203]), .A2(in[135]), .ZN(n711) );
  AND2_X1 U251bar ( .A1(inbar[203]), .A2(inbar[135]), .ZN(n711bar);
  OR2_X1 U252 ( .A1(in[232]), .A2(in[223]), .ZN(n712) );
  AND2_X1 U252bar ( .A1(inbar[232]), .A2(inbar[223]), .ZN(n712bar);
  OR2_X1 U253 ( .A1(n710), .A2(n709), .ZN(n718) );
  AND2_X1 U253bar ( .A1(n710bar), .A2(n709bar), .ZN(n718bar);
  OR2_X1 U254 ( .A1(n708), .A2(n707), .ZN(n709) );
  AND2_X1 U254bar ( .A1(n708bar), .A2(n707bar), .ZN(n709bar);
  OR2_X1 U255 ( .A1(in[255]), .A2(in[233]), .ZN(n707) );
  AND2_X1 U255bar ( .A1(inbar[255]), .A2(inbar[233]), .ZN(n707bar);
  OR2_X1 U256 ( .A1(in_53), .A2(in_34), .ZN(n708) );
  AND2_X1 U256bar ( .A1(in_53bar), .A2(in_34bar), .ZN(n708bar);
  OR2_X1 U257 ( .A1(n706), .A2(n705), .ZN(n710) );
  AND2_X1 U257bar ( .A1(n706bar), .A2(n705bar), .ZN(n710bar);
  OR2_X1 U258 ( .A1(in_57), .A2(in_55), .ZN(n705) );
  AND2_X1 U258bar ( .A1(in_57bar), .A2(in_55bar), .ZN(n705bar);
  OR2_X1 U259 ( .A1(in_68), .A2(in_67), .ZN(n706) );
  AND2_X1 U259bar ( .A1(in_68bar), .A2(in_67bar), .ZN(n706bar);
  OR2_X1 U260 ( .A1(n704), .A2(n703), .ZN(n921) );
  AND2_X1 U260bar ( .A1(n704bar), .A2(n703bar), .ZN(n921bar);
  OR2_X1 U261 ( .A1(n702), .A2(n701), .ZN(n703) );
  AND2_X1 U261bar ( .A1(n702bar), .A2(n701bar), .ZN(n703bar);
  OR2_X1 U262 ( .A1(n700), .A2(n699), .ZN(n701) );
  AND2_X1 U262bar ( .A1(n700bar), .A2(n699bar), .ZN(n701bar);
  OR2_X1 U263 ( .A1(n944), .A2(n872), .ZN(n699) );
  AND2_X1 U263bar ( .A1(n944bar), .A2(n872bar), .ZN(n699bar);
  OR2_X1 U264 ( .A1(n698), .A2(n697), .ZN(n872) );
  AND2_X1 U264bar ( .A1(n698bar), .A2(n697bar), .ZN(n872bar);
  OR2_X1 U265 ( .A1(n696), .A2(n695), .ZN(n697) );
  AND2_X1 U265bar ( .A1(n696bar), .A2(n695bar), .ZN(n697bar);
  OR2_X1 U266 ( .A1(n694), .A2(n693), .ZN(n695) );
  AND2_X1 U266bar ( .A1(n694bar), .A2(n693bar), .ZN(n695bar);
  OR2_X1 U267 ( .A1(in[121]), .A2(in[102]), .ZN(n693) );
  AND2_X1 U267bar ( .A1(inbar[121]), .A2(inbar[102]), .ZN(n693bar);
  OR2_X1 U268 ( .A1(in[162]), .A2(in[161]), .ZN(n694) );
  AND2_X1 U268bar ( .A1(inbar[162]), .A2(inbar[161]), .ZN(n694bar);
  OR2_X1 U269 ( .A1(n692), .A2(n691), .ZN(n696) );
  AND2_X1 U269bar ( .A1(n692bar), .A2(n691bar), .ZN(n696bar);
  OR2_X1 U270 ( .A1(in[192]), .A2(in[178]), .ZN(n691) );
  AND2_X1 U270bar ( .A1(inbar[192]), .A2(inbar[178]), .ZN(n691bar);
  OR2_X1 U271 ( .A1(in[244]), .A2(in[209]), .ZN(n692) );
  AND2_X1 U271bar ( .A1(inbar[244]), .A2(inbar[209]), .ZN(n692bar);
  OR2_X1 U272 ( .A1(n690), .A2(n689), .ZN(n698) );
  AND2_X1 U272bar ( .A1(n690bar), .A2(n689bar), .ZN(n698bar);
  OR2_X1 U273 ( .A1(n688), .A2(n687), .ZN(n689) );
  AND2_X1 U273bar ( .A1(n688bar), .A2(n687bar), .ZN(n689bar);
  OR2_X1 U274 ( .A1(in[90]), .A2(in[254]), .ZN(n687) );
  AND2_X1 U274bar ( .A1(inbar[90]), .A2(inbar[254]), .ZN(n687bar);
  OR2_X1 U275 ( .A1(in_36), .A2(in_32), .ZN(n688) );
  AND2_X1 U275bar ( .A1(in_36bar), .A2(in_32bar), .ZN(n688bar);
  OR2_X1 U276 ( .A1(n686), .A2(n685), .ZN(n690) );
  AND2_X1 U276bar ( .A1(n686bar), .A2(n685bar), .ZN(n690bar);
  OR2_X1 U277 ( .A1(in_62), .A2(in_37), .ZN(n685) );
  AND2_X1 U277bar ( .A1(in_62bar), .A2(in_37bar), .ZN(n685bar);
  OR2_X1 U278 ( .A1(in_75), .A2(in_73), .ZN(n686) );
  AND2_X1 U278bar ( .A1(in_75bar), .A2(in_73bar), .ZN(n686bar);
  OR2_X1 U279 ( .A1(n684), .A2(n683), .ZN(n944) );
  AND2_X1 U279bar ( .A1(n684bar), .A2(n683bar), .ZN(n944bar);
  OR2_X1 U280 ( .A1(n682), .A2(n681), .ZN(n683) );
  AND2_X1 U280bar ( .A1(n682bar), .A2(n681bar), .ZN(n683bar);
  OR2_X1 U281 ( .A1(n680), .A2(n679), .ZN(n681) );
  AND2_X1 U281bar ( .A1(n680bar), .A2(n679bar), .ZN(n681bar);
  OR2_X1 U282 ( .A1(in[171]), .A2(in[153]), .ZN(n679) );
  AND2_X1 U282bar ( .A1(inbar[171]), .A2(inbar[153]), .ZN(n679bar);
  OR2_X1 U283 ( .A1(in[187]), .A2(in[176]), .ZN(n680) );
  AND2_X1 U283bar ( .A1(inbar[187]), .A2(inbar[176]), .ZN(n680bar);
  OR2_X1 U284 ( .A1(n678), .A2(n677), .ZN(n682) );
  AND2_X1 U284bar ( .A1(n678bar), .A2(n677bar), .ZN(n682bar);
  OR2_X1 U285 ( .A1(in[245]), .A2(in[211]), .ZN(n677) );
  AND2_X1 U285bar ( .A1(inbar[245]), .A2(inbar[211]), .ZN(n677bar);
  OR2_X1 U286 ( .A1(in[97]), .A2(in[88]), .ZN(n678) );
  AND2_X1 U286bar ( .A1(inbar[97]), .A2(inbar[88]), .ZN(n678bar);
  OR2_X1 U287 ( .A1(n676), .A2(n675), .ZN(n684) );
  AND2_X1 U287bar ( .A1(n676bar), .A2(n675bar), .ZN(n684bar);
  OR2_X1 U288 ( .A1(n674), .A2(n673), .ZN(n675) );
  AND2_X1 U288bar ( .A1(n674bar), .A2(n673bar), .ZN(n675bar);
  OR2_X1 U289 ( .A1(in_10), .A2(in_0), .ZN(n673) );
  AND2_X1 U289bar ( .A1(in_10bar), .A2(in_0bar), .ZN(n673bar);
  OR2_X1 U290 ( .A1(in_59), .A2(in_5), .ZN(n674) );
  AND2_X1 U290bar ( .A1(in_59bar), .A2(in_5bar), .ZN(n674bar);
  OR2_X1 U291 ( .A1(n672), .A2(n671), .ZN(n676) );
  AND2_X1 U291bar ( .A1(n672bar), .A2(n671bar), .ZN(n676bar);
  OR2_X1 U292 ( .A1(in_60), .A2(in_6), .ZN(n671) );
  AND2_X1 U292bar ( .A1(in_60bar), .A2(in_6bar), .ZN(n671bar);
  OR2_X1 U293 ( .A1(in_77), .A2(in_69), .ZN(n672) );
  AND2_X1 U293bar ( .A1(in_77bar), .A2(in_69bar), .ZN(n672bar);
  OR2_X1 U294 ( .A1(in[113]), .A2(n864), .ZN(n700) );
  AND2_X1 U294bar ( .A1(inbar[113]), .A2(n864bar), .ZN(n700bar);
  OR2_X1 U295 ( .A1(n670), .A2(n669), .ZN(n864) );
  AND2_X1 U295bar ( .A1(n670bar), .A2(n669bar), .ZN(n864bar);
  OR2_X1 U296 ( .A1(n668), .A2(n667), .ZN(n669) );
  AND2_X1 U296bar ( .A1(n668bar), .A2(n667bar), .ZN(n669bar);
  OR2_X1 U297 ( .A1(n666), .A2(n665), .ZN(n667) );
  AND2_X1 U297bar ( .A1(n666bar), .A2(n665bar), .ZN(n667bar);
  OR2_X1 U298 ( .A1(in[125]), .A2(in[107]), .ZN(n665) );
  AND2_X1 U298bar ( .A1(inbar[125]), .A2(inbar[107]), .ZN(n665bar);
  OR2_X1 U299 ( .A1(in[138]), .A2(in[126]), .ZN(n666) );
  AND2_X1 U299bar ( .A1(inbar[138]), .A2(inbar[126]), .ZN(n666bar);
  OR2_X1 U300 ( .A1(n664), .A2(n663), .ZN(n668) );
  AND2_X1 U300bar ( .A1(n664bar), .A2(n663bar), .ZN(n668bar);
  OR2_X1 U301 ( .A1(in[189]), .A2(in[143]), .ZN(n663) );
  AND2_X1 U301bar ( .A1(inbar[189]), .A2(inbar[143]), .ZN(n663bar);
  OR2_X1 U302 ( .A1(in[99]), .A2(in[214]), .ZN(n664) );
  AND2_X1 U302bar ( .A1(inbar[99]), .A2(inbar[214]), .ZN(n664bar);
  OR2_X1 U303 ( .A1(n662), .A2(n661), .ZN(n670) );
  AND2_X1 U303bar ( .A1(n662bar), .A2(n661bar), .ZN(n670bar);
  OR2_X1 U304 ( .A1(n660), .A2(n659), .ZN(n661) );
  AND2_X1 U304bar ( .A1(n660bar), .A2(n659bar), .ZN(n661bar);
  OR2_X1 U305 ( .A1(in_15), .A2(in_12), .ZN(n659) );
  AND2_X1 U305bar ( .A1(in_15bar), .A2(in_12bar), .ZN(n659bar);
  OR2_X1 U306 ( .A1(in_20), .A2(in_2), .ZN(n660) );
  AND2_X1 U306bar ( .A1(in_20bar), .A2(in_2bar), .ZN(n660bar);
  OR2_X1 U307 ( .A1(n658), .A2(n657), .ZN(n662) );
  AND2_X1 U307bar ( .A1(n658bar), .A2(n657bar), .ZN(n662bar);
  OR2_X1 U308 ( .A1(in_30), .A2(in_3), .ZN(n657) );
  AND2_X1 U308bar ( .A1(in_30bar), .A2(in_3bar), .ZN(n657bar);
  OR2_X1 U309 ( .A1(in_4), .A2(in_38), .ZN(n658) );
  AND2_X1 U309bar ( .A1(in_4bar), .A2(in_38bar), .ZN(n658bar);
  OR2_X1 U310 ( .A1(n656), .A2(n655), .ZN(n702) );
  AND2_X1 U310bar ( .A1(n656bar), .A2(n655bar), .ZN(n702bar);
  OR2_X1 U311 ( .A1(in[148]), .A2(in[137]), .ZN(n655) );
  AND2_X1 U311bar ( .A1(inbar[148]), .A2(inbar[137]), .ZN(n655bar);
  OR2_X1 U312 ( .A1(in[149]), .A2(n654), .ZN(n656) );
  AND2_X1 U312bar ( .A1(inbar[149]), .A2(n654bar), .ZN(n656bar);
  OR2_X1 U313 ( .A1(in[195]), .A2(in[190]), .ZN(n654) );
  AND2_X1 U313bar ( .A1(inbar[195]), .A2(inbar[190]), .ZN(n654bar);
  OR2_X1 U314 ( .A1(n653), .A2(n652), .ZN(n704) );
  AND2_X1 U314bar ( .A1(n653bar), .A2(n652bar), .ZN(n704bar);
  OR2_X1 U315 ( .A1(n651), .A2(n650), .ZN(n652) );
  AND2_X1 U315bar ( .A1(n651bar), .A2(n650bar), .ZN(n652bar);
  OR2_X1 U316 ( .A1(in[98]), .A2(in[197]), .ZN(n650) );
  AND2_X1 U316bar ( .A1(inbar[98]), .A2(inbar[197]), .ZN(n650bar);
  OR2_X1 U317 ( .A1(in_11), .A2(n649), .ZN(n651) );
  AND2_X1 U317bar ( .A1(in_11bar), .A2(n649bar), .ZN(n651bar);
  OR2_X1 U318 ( .A1(in_26), .A2(in_14), .ZN(n649) );
  AND2_X1 U318bar ( .A1(in_26bar), .A2(in_14bar), .ZN(n649bar);
  OR2_X1 U319 ( .A1(n648), .A2(n647), .ZN(n653) );
  AND2_X1 U319bar ( .A1(n648bar), .A2(n647bar), .ZN(n653bar);
  OR2_X1 U320 ( .A1(in_35), .A2(in_27), .ZN(n647) );
  AND2_X1 U320bar ( .A1(in_35bar), .A2(in_27bar), .ZN(n647bar);
  OR2_X1 U321 ( .A1(in_50), .A2(n646), .ZN(n648) );
  AND2_X1 U321bar ( .A1(in_50bar), .A2(n646bar), .ZN(n648bar);
  OR2_X1 U322 ( .A1(in_78), .A2(in_61), .ZN(n646) );
  AND2_X1 U322bar ( .A1(in_78bar), .A2(in_61bar), .ZN(n646bar);
  OR2_X1 U323 ( .A1(n942), .A2(n645), .ZN(n720) );
  AND2_X1 U323bar ( .A1(n942bar), .A2(n645bar), .ZN(n720bar);
  OR2_X1 U324 ( .A1(in[106]), .A2(n863), .ZN(n645) );
  AND2_X1 U324bar ( .A1(inbar[106]), .A2(n863bar), .ZN(n645bar);
  OR2_X1 U325 ( .A1(n644), .A2(n643), .ZN(n863) );
  AND2_X1 U325bar ( .A1(n644bar), .A2(n643bar), .ZN(n863bar);
  OR2_X1 U326 ( .A1(n642), .A2(n641), .ZN(n643) );
  AND2_X1 U326bar ( .A1(n642bar), .A2(n641bar), .ZN(n643bar);
  OR2_X1 U327 ( .A1(n640), .A2(n639), .ZN(n641) );
  AND2_X1 U327bar ( .A1(n640bar), .A2(n639bar), .ZN(n641bar);
  OR2_X1 U328 ( .A1(in[127]), .A2(in[122]), .ZN(n639) );
  AND2_X1 U328bar ( .A1(inbar[127]), .A2(inbar[122]), .ZN(n639bar);
  OR2_X1 U329 ( .A1(in[156]), .A2(in[132]), .ZN(n640) );
  AND2_X1 U329bar ( .A1(inbar[156]), .A2(inbar[132]), .ZN(n640bar);
  OR2_X1 U330 ( .A1(n638), .A2(n637), .ZN(n642) );
  AND2_X1 U330bar ( .A1(n638bar), .A2(n637bar), .ZN(n642bar);
  OR2_X1 U331 ( .A1(in[159]), .A2(in[157]), .ZN(n637) );
  AND2_X1 U331bar ( .A1(inbar[159]), .A2(inbar[157]), .ZN(n637bar);
  OR2_X1 U332 ( .A1(in[185]), .A2(in[169]), .ZN(n638) );
  AND2_X1 U332bar ( .A1(inbar[185]), .A2(inbar[169]), .ZN(n638bar);
  OR2_X1 U333 ( .A1(n636), .A2(n635), .ZN(n644) );
  AND2_X1 U333bar ( .A1(n636bar), .A2(n635bar), .ZN(n644bar);
  OR2_X1 U334 ( .A1(n634), .A2(n633), .ZN(n635) );
  AND2_X1 U334bar ( .A1(n634bar), .A2(n633bar), .ZN(n635bar);
  OR2_X1 U335 ( .A1(in[239]), .A2(in[218]), .ZN(n633) );
  AND2_X1 U335bar ( .A1(inbar[239]), .A2(inbar[218]), .ZN(n633bar);
  OR2_X1 U336 ( .A1(in_13), .A2(in[87]), .ZN(n634) );
  AND2_X1 U336bar ( .A1(in_13bar), .A2(inbar[87]), .ZN(n634bar);
  OR2_X1 U337 ( .A1(n632), .A2(n631), .ZN(n636) );
  AND2_X1 U337bar ( .A1(n632bar), .A2(n631bar), .ZN(n636bar);
  OR2_X1 U338 ( .A1(in_72), .A2(in_70), .ZN(n631) );
  AND2_X1 U338bar ( .A1(in_72bar), .A2(in_70bar), .ZN(n631bar);
  OR2_X1 U339 ( .A1(in_80), .A2(in_74), .ZN(n632) );
  AND2_X1 U339bar ( .A1(in_80bar), .A2(in_74bar), .ZN(n632bar);
  OR2_X1 U340 ( .A1(n630), .A2(n629), .ZN(n942) );
  AND2_X1 U340bar ( .A1(n630bar), .A2(n629bar), .ZN(n942bar);
  OR2_X1 U341 ( .A1(n628), .A2(n627), .ZN(n629) );
  AND2_X1 U341bar ( .A1(n628bar), .A2(n627bar), .ZN(n629bar);
  OR2_X1 U342 ( .A1(n626), .A2(n625), .ZN(n627) );
  AND2_X1 U342bar ( .A1(n626bar), .A2(n625bar), .ZN(n627bar);
  OR2_X1 U343 ( .A1(in[146]), .A2(in[100]), .ZN(n625) );
  AND2_X1 U343bar ( .A1(inbar[146]), .A2(inbar[100]), .ZN(n625bar);
  OR2_X1 U344 ( .A1(in[168]), .A2(in[152]), .ZN(n626) );
  AND2_X1 U344bar ( .A1(inbar[168]), .A2(inbar[152]), .ZN(n626bar);
  OR2_X1 U345 ( .A1(n624), .A2(n623), .ZN(n628) );
  AND2_X1 U345bar ( .A1(n624bar), .A2(n623bar), .ZN(n628bar);
  OR2_X1 U346 ( .A1(in[199]), .A2(in[182]), .ZN(n623) );
  AND2_X1 U346bar ( .A1(inbar[199]), .A2(inbar[182]), .ZN(n623bar);
  OR2_X1 U347 ( .A1(in[236]), .A2(in[204]), .ZN(n624) );
  AND2_X1 U347bar ( .A1(inbar[236]), .A2(inbar[204]), .ZN(n624bar);
  OR2_X1 U348 ( .A1(n622), .A2(n621), .ZN(n630) );
  AND2_X1 U348bar ( .A1(n622bar), .A2(n621bar), .ZN(n630bar);
  OR2_X1 U349 ( .A1(n620), .A2(n619), .ZN(n621) );
  AND2_X1 U349bar ( .A1(n620bar), .A2(n619bar), .ZN(n621bar);
  OR2_X1 U350 ( .A1(in[89]), .A2(in[246]), .ZN(n619) );
  AND2_X1 U350bar ( .A1(inbar[89]), .A2(inbar[246]), .ZN(n619bar);
  OR2_X1 U351 ( .A1(in[95]), .A2(in[92]), .ZN(n620) );
  AND2_X1 U351bar ( .A1(inbar[95]), .A2(inbar[92]), .ZN(n620bar);
  OR2_X1 U352 ( .A1(n618), .A2(n617), .ZN(n622) );
  AND2_X1 U352bar ( .A1(n618bar), .A2(n617bar), .ZN(n622bar);
  OR2_X1 U353 ( .A1(in_22), .A2(in_16), .ZN(n617) );
  AND2_X1 U353bar ( .A1(in_22bar), .A2(in_16bar), .ZN(n617bar);
  OR2_X1 U354 ( .A1(in_51), .A2(in_49), .ZN(n618) );
  AND2_X1 U354bar ( .A1(in_51bar), .A2(in_49bar), .ZN(n618bar);
  OR2_X1 U355 ( .A1(n616), .A2(n615), .ZN(n722) );
  AND2_X1 U355bar ( .A1(n616bar), .A2(n615bar), .ZN(n722bar);
  OR2_X1 U356 ( .A1(in[158]), .A2(in[115]), .ZN(n615) );
  AND2_X1 U356bar ( .A1(inbar[158]), .A2(inbar[115]), .ZN(n615bar);
  OR2_X1 U357 ( .A1(in[163]), .A2(n614), .ZN(n616) );
  AND2_X1 U357bar ( .A1(inbar[163]), .A2(n614bar), .ZN(n616bar);
  OR2_X1 U358 ( .A1(in[206]), .A2(in[165]), .ZN(n614) );
  AND2_X1 U358bar ( .A1(inbar[206]), .A2(inbar[165]), .ZN(n614bar);
  OR2_X1 U359 ( .A1(n613), .A2(n612), .ZN(n724) );
  AND2_X1 U359bar ( .A1(n613bar), .A2(n612bar), .ZN(n724bar);
  OR2_X1 U360 ( .A1(n611), .A2(n610), .ZN(n612) );
  AND2_X1 U360bar ( .A1(n611bar), .A2(n610bar), .ZN(n612bar);
  OR2_X1 U361 ( .A1(in[213]), .A2(in[207]), .ZN(n610) );
  AND2_X1 U361bar ( .A1(inbar[213]), .A2(inbar[207]), .ZN(n610bar);
  OR2_X1 U362 ( .A1(in[215]), .A2(n609), .ZN(n611) );
  AND2_X1 U362bar ( .A1(inbar[215]), .A2(n609bar), .ZN(n611bar);
  OR2_X1 U363 ( .A1(in[230]), .A2(in[220]), .ZN(n609) );
  AND2_X1 U363bar ( .A1(inbar[230]), .A2(inbar[220]), .ZN(n609bar);
  OR2_X1 U364 ( .A1(n608), .A2(n607), .ZN(n613) );
  AND2_X1 U364bar ( .A1(n608bar), .A2(n607bar), .ZN(n613bar);
  OR2_X1 U365 ( .A1(in[251]), .A2(in[234]), .ZN(n607) );
  AND2_X1 U365bar ( .A1(inbar[251]), .A2(inbar[234]), .ZN(n607bar);
  OR2_X1 U366 ( .A1(in_17), .A2(n606), .ZN(n608) );
  AND2_X1 U366bar ( .A1(in_17bar), .A2(n606bar), .ZN(n608bar);
  OR2_X1 U367 ( .A1(in_65), .A2(in_56), .ZN(n606) );
  AND2_X1 U367bar ( .A1(in_65bar), .A2(in_56bar), .ZN(n606bar);
  OR2_X1 U368 ( .A1(n605), .A2(n604), .ZN(out[0]) );
  AND2_X1 U368bar ( .A1(n605bar), .A2(n604bar), .ZN(outbar[0]);
  OR2_X1 U369 ( .A1(n603), .A2(n602), .ZN(n604) );
  AND2_X1 U369bar ( .A1(n603bar), .A2(n602bar), .ZN(n604bar);
  OR2_X1 U370 ( .A1(n601), .A2(n600), .ZN(n602) );
  AND2_X1 U370bar ( .A1(n601bar), .A2(n600bar), .ZN(n602bar);
  OR2_X1 U371 ( .A1(n820), .A2(n785), .ZN(n600) );
  AND2_X1 U371bar ( .A1(n820bar), .A2(n785bar), .ZN(n600bar);
  OR2_X1 U372 ( .A1(n599), .A2(n598), .ZN(n785) );
  AND2_X1 U372bar ( .A1(n599bar), .A2(n598bar), .ZN(n785bar);
  OR2_X1 U373 ( .A1(n597), .A2(n596), .ZN(n598) );
  AND2_X1 U373bar ( .A1(n597bar), .A2(n596bar), .ZN(n598bar);
  OR2_X1 U374 ( .A1(n595), .A2(n594), .ZN(n596) );
  AND2_X1 U374bar ( .A1(n595bar), .A2(n594bar), .ZN(n596bar);
  OR2_X1 U375 ( .A1(in[135]), .A2(in[104]), .ZN(n594) );
  AND2_X1 U375bar ( .A1(inbar[135]), .A2(inbar[104]), .ZN(n594bar);
  OR2_X1 U376 ( .A1(in[188]), .A2(in[178]), .ZN(n595) );
  AND2_X1 U376bar ( .A1(inbar[188]), .A2(inbar[178]), .ZN(n595bar);
  OR2_X1 U377 ( .A1(n593), .A2(n592), .ZN(n597) );
  AND2_X1 U377bar ( .A1(n593bar), .A2(n592bar), .ZN(n597bar);
  OR2_X1 U378 ( .A1(in[217]), .A2(in[194]), .ZN(n592) );
  AND2_X1 U378bar ( .A1(inbar[217]), .A2(inbar[194]), .ZN(n592bar);
  OR2_X1 U379 ( .A1(in[237]), .A2(in[218]), .ZN(n593) );
  AND2_X1 U379bar ( .A1(inbar[237]), .A2(inbar[218]), .ZN(n593bar);
  OR2_X1 U380 ( .A1(n591), .A2(n590), .ZN(n599) );
  AND2_X1 U380bar ( .A1(n591bar), .A2(n590bar), .ZN(n599bar);
  OR2_X1 U381 ( .A1(n589), .A2(n588), .ZN(n590) );
  AND2_X1 U381bar ( .A1(n589bar), .A2(n588bar), .ZN(n590bar);
  OR2_X1 U382 ( .A1(in_2), .A2(in_10), .ZN(n588) );
  AND2_X1 U382bar ( .A1(in_2bar), .A2(in_10bar), .ZN(n588bar);
  OR2_X1 U383 ( .A1(in_47), .A2(in_22), .ZN(n589) );
  AND2_X1 U383bar ( .A1(in_47bar), .A2(in_22bar), .ZN(n589bar);
  OR2_X1 U384 ( .A1(n587), .A2(n586), .ZN(n591) );
  AND2_X1 U384bar ( .A1(n587bar), .A2(n586bar), .ZN(n591bar);
  OR2_X1 U385 ( .A1(in_56), .A2(in_54), .ZN(n586) );
  AND2_X1 U385bar ( .A1(in_56bar), .A2(in_54bar), .ZN(n586bar);
  OR2_X1 U386 ( .A1(in_63), .A2(in_61), .ZN(n587) );
  AND2_X1 U386bar ( .A1(in_63bar), .A2(in_61bar), .ZN(n587bar);
  OR2_X1 U387 ( .A1(n585), .A2(n584), .ZN(n820) );
  AND2_X1 U387bar ( .A1(n585bar), .A2(n584bar), .ZN(n820bar);
  OR2_X1 U388 ( .A1(n583), .A2(n582), .ZN(n584) );
  AND2_X1 U388bar ( .A1(n583bar), .A2(n582bar), .ZN(n584bar);
  OR2_X1 U389 ( .A1(n581), .A2(n580), .ZN(n582) );
  AND2_X1 U389bar ( .A1(n581bar), .A2(n580bar), .ZN(n582bar);
  OR2_X1 U390 ( .A1(in[158]), .A2(in[142]), .ZN(n580) );
  AND2_X1 U390bar ( .A1(inbar[158]), .A2(inbar[142]), .ZN(n580bar);
  OR2_X1 U391 ( .A1(in[175]), .A2(in[164]), .ZN(n581) );
  AND2_X1 U391bar ( .A1(inbar[175]), .A2(inbar[164]), .ZN(n581bar);
  OR2_X1 U392 ( .A1(n579), .A2(n578), .ZN(n583) );
  AND2_X1 U392bar ( .A1(n579bar), .A2(n578bar), .ZN(n583bar);
  OR2_X1 U393 ( .A1(in[228]), .A2(in[204]), .ZN(n578) );
  AND2_X1 U393bar ( .A1(inbar[228]), .A2(inbar[204]), .ZN(n578bar);
  OR2_X1 U394 ( .A1(in[91]), .A2(in[87]), .ZN(n579) );
  AND2_X1 U394bar ( .A1(inbar[91]), .A2(inbar[87]), .ZN(n579bar);
  OR2_X1 U395 ( .A1(n577), .A2(n576), .ZN(n585) );
  AND2_X1 U395bar ( .A1(n577bar), .A2(n576bar), .ZN(n585bar);
  OR2_X1 U396 ( .A1(n575), .A2(n574), .ZN(n576) );
  AND2_X1 U396bar ( .A1(n575bar), .A2(n574bar), .ZN(n576bar);
  OR2_X1 U397 ( .A1(in_21), .A2(in_11), .ZN(n574) );
  AND2_X1 U397bar ( .A1(in_21bar), .A2(in_11bar), .ZN(n574bar);
  OR2_X1 U398 ( .A1(in_5), .A2(in_3), .ZN(n575) );
  AND2_X1 U398bar ( .A1(in_5bar), .A2(in_3bar), .ZN(n575bar);
  OR2_X1 U399 ( .A1(n573), .A2(n572), .ZN(n577) );
  AND2_X1 U399bar ( .A1(n573bar), .A2(n572bar), .ZN(n577bar);
  OR2_X1 U400 ( .A1(in_68), .A2(in_64), .ZN(n572) );
  AND2_X1 U400bar ( .A1(in_68bar), .A2(in_64bar), .ZN(n572bar);
  OR2_X1 U401 ( .A1(in_76), .A2(in_73), .ZN(n573) );
  AND2_X1 U401bar ( .A1(in_76bar), .A2(in_73bar), .ZN(n573bar);
  OR2_X1 U402 ( .A1(n778), .A2(n571), .ZN(n601) );
  AND2_X1 U402bar ( .A1(n778bar), .A2(n571bar), .ZN(n601bar);
  OR2_X1 U403 ( .A1(in[100]), .A2(n965), .ZN(n571) );
  AND2_X1 U403bar ( .A1(inbar[100]), .A2(n965bar), .ZN(n571bar);
  OR2_X1 U404 ( .A1(n570), .A2(n569), .ZN(n965) );
  AND2_X1 U404bar ( .A1(n570bar), .A2(n569bar), .ZN(n965bar);
  OR2_X1 U405 ( .A1(n568), .A2(n567), .ZN(n569) );
  AND2_X1 U405bar ( .A1(n568bar), .A2(n567bar), .ZN(n569bar);
  OR2_X1 U406 ( .A1(n566), .A2(n565), .ZN(n567) );
  AND2_X1 U406bar ( .A1(n566bar), .A2(n565bar), .ZN(n567bar);
  OR2_X1 U407 ( .A1(n817), .A2(n750), .ZN(n565) );
  AND2_X1 U407bar ( .A1(n817bar), .A2(n750bar), .ZN(n565bar);
  OR2_X1 U408 ( .A1(n564), .A2(n563), .ZN(n750) );
  AND2_X1 U408bar ( .A1(n564bar), .A2(n563bar), .ZN(n750bar);
  OR2_X1 U409 ( .A1(n562), .A2(n561), .ZN(n563) );
  AND2_X1 U409bar ( .A1(n562bar), .A2(n561bar), .ZN(n563bar);
  OR2_X1 U410 ( .A1(n560), .A2(n559), .ZN(n561) );
  AND2_X1 U410bar ( .A1(n560bar), .A2(n559bar), .ZN(n561bar);
  OR2_X1 U411 ( .A1(in[119]), .A2(in[103]), .ZN(n559) );
  AND2_X1 U411bar ( .A1(inbar[119]), .A2(inbar[103]), .ZN(n559bar);
  OR2_X1 U412 ( .A1(in[137]), .A2(in[133]), .ZN(n560) );
  AND2_X1 U412bar ( .A1(inbar[137]), .A2(inbar[133]), .ZN(n560bar);
  OR2_X1 U413 ( .A1(n558), .A2(n557), .ZN(n562) );
  AND2_X1 U413bar ( .A1(n558bar), .A2(n557bar), .ZN(n562bar);
  OR2_X1 U414 ( .A1(in[176]), .A2(in[173]), .ZN(n557) );
  AND2_X1 U414bar ( .A1(inbar[176]), .A2(inbar[173]), .ZN(n557bar);
  OR2_X1 U415 ( .A1(in[210]), .A2(in[181]), .ZN(n558) );
  AND2_X1 U415bar ( .A1(inbar[210]), .A2(inbar[181]), .ZN(n558bar);
  OR2_X1 U416 ( .A1(n556), .A2(n555), .ZN(n564) );
  AND2_X1 U416bar ( .A1(n556bar), .A2(n555bar), .ZN(n564bar);
  OR2_X1 U417 ( .A1(n554), .A2(n553), .ZN(n555) );
  AND2_X1 U417bar ( .A1(n554bar), .A2(n553bar), .ZN(n555bar);
  OR2_X1 U418 ( .A1(in_13), .A2(in[234]), .ZN(n553) );
  AND2_X1 U418bar ( .A1(in_13bar), .A2(inbar[234]), .ZN(n553bar);
  OR2_X1 U419 ( .A1(in_38), .A2(in_32), .ZN(n554) );
  AND2_X1 U419bar ( .A1(in_38bar), .A2(in_32bar), .ZN(n554bar);
  OR2_X1 U420 ( .A1(n552), .A2(n551), .ZN(n556) );
  AND2_X1 U420bar ( .A1(n552bar), .A2(n551bar), .ZN(n556bar);
  OR2_X1 U421 ( .A1(in_42), .A2(in_41), .ZN(n551) );
  AND2_X1 U421bar ( .A1(in_42bar), .A2(in_41bar), .ZN(n551bar);
  OR2_X1 U422 ( .A1(in_7), .A2(in_49), .ZN(n552) );
  AND2_X1 U422bar ( .A1(in_7bar), .A2(in_49bar), .ZN(n552bar);
  OR2_X1 U423 ( .A1(n550), .A2(n549), .ZN(n817) );
  AND2_X1 U423bar ( .A1(n550bar), .A2(n549bar), .ZN(n817bar);
  OR2_X1 U424 ( .A1(n548), .A2(n547), .ZN(n549) );
  AND2_X1 U424bar ( .A1(n548bar), .A2(n547bar), .ZN(n549bar);
  OR2_X1 U425 ( .A1(n546), .A2(n545), .ZN(n547) );
  AND2_X1 U425bar ( .A1(n546bar), .A2(n545bar), .ZN(n547bar);
  OR2_X1 U426 ( .A1(in[159]), .A2(in[105]), .ZN(n545) );
  AND2_X1 U426bar ( .A1(inbar[159]), .A2(inbar[105]), .ZN(n545bar);
  OR2_X1 U427 ( .A1(in[206]), .A2(in[183]), .ZN(n546) );
  AND2_X1 U427bar ( .A1(inbar[206]), .A2(inbar[183]), .ZN(n546bar);
  OR2_X1 U428 ( .A1(n544), .A2(n543), .ZN(n548) );
  AND2_X1 U428bar ( .A1(n544bar), .A2(n543bar), .ZN(n548bar);
  OR2_X1 U429 ( .A1(in[229]), .A2(in[219]), .ZN(n543) );
  AND2_X1 U429bar ( .A1(inbar[229]), .A2(inbar[219]), .ZN(n543bar);
  OR2_X1 U430 ( .A1(in[235]), .A2(in[232]), .ZN(n544) );
  AND2_X1 U430bar ( .A1(inbar[235]), .A2(inbar[232]), .ZN(n544bar);
  OR2_X1 U431 ( .A1(n542), .A2(n541), .ZN(n550) );
  AND2_X1 U431bar ( .A1(n542bar), .A2(n541bar), .ZN(n550bar);
  OR2_X1 U432 ( .A1(n540), .A2(n539), .ZN(n541) );
  AND2_X1 U432bar ( .A1(n540bar), .A2(n539bar), .ZN(n541bar);
  OR2_X1 U433 ( .A1(in[249]), .A2(in[242]), .ZN(n539) );
  AND2_X1 U433bar ( .A1(inbar[249]), .A2(inbar[242]), .ZN(n539bar);
  OR2_X1 U434 ( .A1(in[89]), .A2(in[254]), .ZN(n540) );
  AND2_X1 U434bar ( .A1(inbar[89]), .A2(inbar[254]), .ZN(n540bar);
  OR2_X1 U435 ( .A1(n538), .A2(n537), .ZN(n542) );
  AND2_X1 U435bar ( .A1(n538bar), .A2(n537bar), .ZN(n542bar);
  OR2_X1 U436 ( .A1(in_14), .A2(in[99]), .ZN(n537) );
  AND2_X1 U436bar ( .A1(in_14bar), .A2(inbar[99]), .ZN(n537bar);
  OR2_X1 U437 ( .A1(in_60), .A2(in_18), .ZN(n538) );
  AND2_X1 U437bar ( .A1(in_60bar), .A2(in_18bar), .ZN(n538bar);
  OR2_X1 U438 ( .A1(in[113]), .A2(n763), .ZN(n566) );
  AND2_X1 U438bar ( .A1(inbar[113]), .A2(n763bar), .ZN(n566bar);
  OR2_X1 U439 ( .A1(n536), .A2(n535), .ZN(n763) );
  AND2_X1 U439bar ( .A1(n536bar), .A2(n535bar), .ZN(n763bar);
  OR2_X1 U440 ( .A1(n534), .A2(n533), .ZN(n535) );
  AND2_X1 U440bar ( .A1(n534bar), .A2(n533bar), .ZN(n535bar);
  OR2_X1 U441 ( .A1(n532), .A2(n531), .ZN(n533) );
  AND2_X1 U441bar ( .A1(n532bar), .A2(n531bar), .ZN(n533bar);
  OR2_X1 U442 ( .A1(in[115]), .A2(in[110]), .ZN(n531) );
  AND2_X1 U442bar ( .A1(inbar[115]), .A2(inbar[110]), .ZN(n531bar);
  OR2_X1 U443 ( .A1(in[125]), .A2(in[117]), .ZN(n532) );
  AND2_X1 U443bar ( .A1(inbar[125]), .A2(inbar[117]), .ZN(n532bar);
  OR2_X1 U444 ( .A1(n530), .A2(n529), .ZN(n534) );
  AND2_X1 U444bar ( .A1(n530bar), .A2(n529bar), .ZN(n534bar);
  OR2_X1 U445 ( .A1(in[180]), .A2(in[128]), .ZN(n529) );
  AND2_X1 U445bar ( .A1(inbar[180]), .A2(inbar[128]), .ZN(n529bar);
  OR2_X1 U446 ( .A1(in[205]), .A2(in[201]), .ZN(n530) );
  AND2_X1 U446bar ( .A1(inbar[205]), .A2(inbar[201]), .ZN(n530bar);
  OR2_X1 U447 ( .A1(n528), .A2(n527), .ZN(n536) );
  AND2_X1 U447bar ( .A1(n528bar), .A2(n527bar), .ZN(n536bar);
  OR2_X1 U448 ( .A1(n526), .A2(n525), .ZN(n527) );
  AND2_X1 U448bar ( .A1(n526bar), .A2(n525bar), .ZN(n527bar);
  OR2_X1 U449 ( .A1(in[244]), .A2(in[239]), .ZN(n525) );
  AND2_X1 U449bar ( .A1(inbar[244]), .A2(inbar[239]), .ZN(n525bar);
  OR2_X1 U450 ( .A1(in[95]), .A2(in[83]), .ZN(n526) );
  AND2_X1 U450bar ( .A1(inbar[95]), .A2(inbar[83]), .ZN(n526bar);
  OR2_X1 U451 ( .A1(n524), .A2(n523), .ZN(n528) );
  AND2_X1 U451bar ( .A1(n524bar), .A2(n523bar), .ZN(n528bar);
  OR2_X1 U452 ( .A1(in_24), .A2(in[97]), .ZN(n523) );
  AND2_X1 U452bar ( .A1(in_24bar), .A2(inbar[97]), .ZN(n523bar);
  OR2_X1 U453 ( .A1(in_33), .A2(in_27), .ZN(n524) );
  AND2_X1 U453bar ( .A1(in_33bar), .A2(in_27bar), .ZN(n524bar);
  OR2_X1 U454 ( .A1(n522), .A2(n521), .ZN(n568) );
  AND2_X1 U454bar ( .A1(n522bar), .A2(n521bar), .ZN(n568bar);
  OR2_X1 U455 ( .A1(in[145]), .A2(in[126]), .ZN(n521) );
  AND2_X1 U455bar ( .A1(inbar[145]), .A2(inbar[126]), .ZN(n521bar);
  OR2_X1 U456 ( .A1(in[169]), .A2(n520), .ZN(n522) );
  AND2_X1 U456bar ( .A1(inbar[169]), .A2(n520bar), .ZN(n522bar);
  OR2_X1 U457 ( .A1(in[221]), .A2(in[172]), .ZN(n520) );
  AND2_X1 U457bar ( .A1(inbar[221]), .A2(inbar[172]), .ZN(n520bar);
  OR2_X1 U458 ( .A1(n519), .A2(n518), .ZN(n570) );
  AND2_X1 U458bar ( .A1(n519bar), .A2(n518bar), .ZN(n570bar);
  OR2_X1 U459 ( .A1(n517), .A2(n516), .ZN(n518) );
  AND2_X1 U459bar ( .A1(n517bar), .A2(n516bar), .ZN(n518bar);
  OR2_X1 U460 ( .A1(in[241]), .A2(in[224]), .ZN(n516) );
  AND2_X1 U460bar ( .A1(inbar[241]), .A2(inbar[224]), .ZN(n516bar);
  OR2_X1 U461 ( .A1(in[86]), .A2(n515), .ZN(n517) );
  AND2_X1 U461bar ( .A1(inbar[86]), .A2(n515bar), .ZN(n517bar);
  OR2_X1 U462 ( .A1(in_43), .A2(in_34), .ZN(n515) );
  AND2_X1 U462bar ( .A1(in_43bar), .A2(in_34bar), .ZN(n515bar);
  OR2_X1 U463 ( .A1(n514), .A2(n513), .ZN(n519) );
  AND2_X1 U463bar ( .A1(n514bar), .A2(n513bar), .ZN(n519bar);
  OR2_X1 U464 ( .A1(in_65), .A2(in_51), .ZN(n513) );
  AND2_X1 U464bar ( .A1(in_65bar), .A2(in_51bar), .ZN(n513bar);
  OR2_X1 U465 ( .A1(in_75), .A2(n512), .ZN(n514) );
  AND2_X1 U465bar ( .A1(in_75bar), .A2(n512bar), .ZN(n514bar);
  OR2_X1 U466 ( .A1(in_81), .A2(in_77), .ZN(n512) );
  AND2_X1 U466bar ( .A1(in_81bar), .A2(in_77bar), .ZN(n512bar);
  OR2_X1 U467 ( .A1(n511), .A2(n510), .ZN(n778) );
  AND2_X1 U467bar ( .A1(n511bar), .A2(n510bar), .ZN(n778bar);
  OR2_X1 U468 ( .A1(n509), .A2(n508), .ZN(n510) );
  AND2_X1 U468bar ( .A1(n509bar), .A2(n508bar), .ZN(n510bar);
  OR2_X1 U469 ( .A1(n507), .A2(n506), .ZN(n508) );
  AND2_X1 U469bar ( .A1(n507bar), .A2(n506bar), .ZN(n508bar);
  OR2_X1 U470 ( .A1(in[107]), .A2(in[101]), .ZN(n506) );
  AND2_X1 U470bar ( .A1(inbar[107]), .A2(inbar[101]), .ZN(n506bar);
  OR2_X1 U471 ( .A1(in[139]), .A2(in[132]), .ZN(n507) );
  AND2_X1 U471bar ( .A1(inbar[139]), .A2(inbar[132]), .ZN(n507bar);
  OR2_X1 U472 ( .A1(n505), .A2(n504), .ZN(n509) );
  AND2_X1 U472bar ( .A1(n505bar), .A2(n504bar), .ZN(n509bar);
  OR2_X1 U473 ( .A1(in[146]), .A2(in[141]), .ZN(n504) );
  AND2_X1 U473bar ( .A1(inbar[146]), .A2(inbar[141]), .ZN(n504bar);
  OR2_X1 U474 ( .A1(in[203]), .A2(in[179]), .ZN(n505) );
  AND2_X1 U474bar ( .A1(inbar[203]), .A2(inbar[179]), .ZN(n505bar);
  OR2_X1 U475 ( .A1(n503), .A2(n502), .ZN(n511) );
  AND2_X1 U475bar ( .A1(n503bar), .A2(n502bar), .ZN(n511bar);
  OR2_X1 U476 ( .A1(n501), .A2(n500), .ZN(n502) );
  AND2_X1 U476bar ( .A1(n501bar), .A2(n500bar), .ZN(n502bar);
  OR2_X1 U477 ( .A1(in[243]), .A2(in[222]), .ZN(n500) );
  AND2_X1 U477bar ( .A1(inbar[243]), .A2(inbar[222]), .ZN(n500bar);
  OR2_X1 U478 ( .A1(in[251]), .A2(in[250]), .ZN(n501) );
  AND2_X1 U478bar ( .A1(inbar[251]), .A2(inbar[250]), .ZN(n501bar);
  OR2_X1 U479 ( .A1(n499), .A2(n498), .ZN(n503) );
  AND2_X1 U479bar ( .A1(n499bar), .A2(n498bar), .ZN(n503bar);
  OR2_X1 U480 ( .A1(in_37), .A2(in_19), .ZN(n498) );
  AND2_X1 U480bar ( .A1(in_37bar), .A2(in_19bar), .ZN(n498bar);
  OR2_X1 U481 ( .A1(in_78), .A2(in_6), .ZN(n499) );
  AND2_X1 U481bar ( .A1(in_78bar), .A2(in_6bar), .ZN(n499bar);
  OR2_X1 U482 ( .A1(n497), .A2(n496), .ZN(n603) );
  AND2_X1 U482bar ( .A1(n497bar), .A2(n496bar), .ZN(n603bar);
  OR2_X1 U483 ( .A1(in[112]), .A2(in[102]), .ZN(n496) );
  AND2_X1 U483bar ( .A1(inbar[112]), .A2(inbar[102]), .ZN(n496bar);
  OR2_X1 U484 ( .A1(in[123]), .A2(n495), .ZN(n497) );
  AND2_X1 U484bar ( .A1(inbar[123]), .A2(n495bar), .ZN(n497bar);
  OR2_X1 U485 ( .A1(in[143]), .A2(in[130]), .ZN(n495) );
  AND2_X1 U485bar ( .A1(inbar[143]), .A2(inbar[130]), .ZN(n495bar);
  OR2_X1 U486 ( .A1(n494), .A2(n493), .ZN(n605) );
  AND2_X1 U486bar ( .A1(n494bar), .A2(n493bar), .ZN(n605bar);
  OR2_X1 U487 ( .A1(n492), .A2(n491), .ZN(n493) );
  AND2_X1 U487bar ( .A1(n492bar), .A2(n491bar), .ZN(n493bar);
  OR2_X1 U488 ( .A1(in[216]), .A2(in[213]), .ZN(n491) );
  AND2_X1 U488bar ( .A1(inbar[216]), .A2(inbar[213]), .ZN(n491bar);
  OR2_X1 U489 ( .A1(in[227]), .A2(n490), .ZN(n492) );
  AND2_X1 U489bar ( .A1(inbar[227]), .A2(n490bar), .ZN(n492bar);
  OR2_X1 U490 ( .A1(in_0), .A2(in[248]), .ZN(n490) );
  AND2_X1 U490bar ( .A1(in_0bar), .A2(inbar[248]), .ZN(n490bar);
  OR2_X1 U491 ( .A1(n489), .A2(n488), .ZN(n494) );
  AND2_X1 U491bar ( .A1(n489bar), .A2(n488bar), .ZN(n494bar);
  OR2_X1 U492 ( .A1(in_46), .A2(in_44), .ZN(n488) );
  AND2_X1 U492bar ( .A1(in_46bar), .A2(in_44bar), .ZN(n488bar);
  OR2_X1 U493 ( .A1(in_50), .A2(n487), .ZN(n489) );
  AND2_X1 U493bar ( .A1(in_50bar), .A2(n487bar), .ZN(n489bar);
  OR2_X1 U494 ( .A1(in_9), .A2(in_80), .ZN(n487) );
  AND2_X1 U494bar ( .A1(in_9bar), .A2(in_80bar), .ZN(n487bar);
endmodule




module sBox_5 ( in, out );
  input [7:0] in;
  //input_done

  output [7:0] out;
  //output_done

  wire   [255:0] decodeOut;
  //wire_done

  decode_5 dec ( .in(in), .out(decodeOut) );
  encode_5 enc ( .in(decodeOut), .out(out) );
endmodule


module CD2_21 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_22 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
 
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_23 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_24 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD4_11 ( a, b, y );
  input [3:0] a;
  input [3:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  //input_done

  output [15:0] y;
  reg [15:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]);
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]);
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]);
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]);
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]);
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]);
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]);
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]);
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]);
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]);
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]);
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]);
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]);
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]);
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]);
endmodule




module CD4_12 ( a, b, y );
  input [3:0] a;
  input [3:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  //input_done

  output [15:0] y;
  reg [15:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]);
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]);
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]);
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]);
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]);
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]);
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]);
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]);
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]);
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]);
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]);
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]);
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]);
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]);
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]);
endmodule




module CD16_6 ( a, b, y );
  input [15:0] a;
  input [15:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign abar[8] = ~a[8];
  assign abar[9] = ~a[9];
  assign abar[10] = ~a[10];
  assign abar[11] = ~a[11];
  assign abar[12] = ~a[12];
  assign abar[13] = ~a[13];
  assign abar[14] = ~a[14];
  assign abar[15] = ~a[15];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign bbar[8] = ~b[8];
  assign bbar[9] = ~b[9];
  assign bbar[10] = ~b[10];
  assign bbar[11] = ~b[11];
  assign bbar[12] = ~b[12];
  assign bbar[13] = ~b[13];
  assign bbar[14] = ~b[14];
  assign bbar[15] = ~b[15];
  //input_done

  output [255:0] y;
  reg [255:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[9]), .A2(a[0]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[9]), .A2(abar[0]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[3]), .A2(a[6]), .ZN(y[99]) );
  OR2_X1 U2bar ( .A1(bbar[3]), .A2(abar[6]), .ZN(ybar[99]);
  AND2_X1 U3 ( .A1(b[2]), .A2(a[6]), .ZN(y[98]) );
  OR2_X1 U3bar ( .A1(bbar[2]), .A2(abar[6]), .ZN(ybar[98]);
  AND2_X1 U4 ( .A1(b[1]), .A2(a[6]), .ZN(y[97]) );
  OR2_X1 U4bar ( .A1(bbar[1]), .A2(abar[6]), .ZN(ybar[97]);
  AND2_X1 U5 ( .A1(b[0]), .A2(a[6]), .ZN(y[96]) );
  OR2_X1 U5bar ( .A1(bbar[0]), .A2(abar[6]), .ZN(ybar[96]);
  AND2_X1 U6 ( .A1(b[15]), .A2(a[5]), .ZN(y[95]) );
  OR2_X1 U6bar ( .A1(bbar[15]), .A2(abar[5]), .ZN(ybar[95]);
  AND2_X1 U7 ( .A1(b[14]), .A2(a[5]), .ZN(y[94]) );
  OR2_X1 U7bar ( .A1(bbar[14]), .A2(abar[5]), .ZN(ybar[94]);
  AND2_X1 U8 ( .A1(b[13]), .A2(a[5]), .ZN(y[93]) );
  OR2_X1 U8bar ( .A1(bbar[13]), .A2(abar[5]), .ZN(ybar[93]);
  AND2_X1 U9 ( .A1(b[12]), .A2(a[5]), .ZN(y[92]) );
  OR2_X1 U9bar ( .A1(bbar[12]), .A2(abar[5]), .ZN(ybar[92]);
  AND2_X1 U10 ( .A1(b[11]), .A2(a[5]), .ZN(y[91]) );
  OR2_X1 U10bar ( .A1(bbar[11]), .A2(abar[5]), .ZN(ybar[91]);
  AND2_X1 U11 ( .A1(b[10]), .A2(a[5]), .ZN(y[90]) );
  OR2_X1 U11bar ( .A1(bbar[10]), .A2(abar[5]), .ZN(ybar[90]);
  AND2_X1 U12 ( .A1(b[8]), .A2(a[0]), .ZN(y[8]) );
  OR2_X1 U12bar ( .A1(bbar[8]), .A2(abar[0]), .ZN(ybar[8]);
  AND2_X1 U13 ( .A1(a[5]), .A2(b[9]), .ZN(y[89]) );
  OR2_X1 U13bar ( .A1(abar[5]), .A2(bbar[9]), .ZN(ybar[89]);
  AND2_X1 U14 ( .A1(b[8]), .A2(a[5]), .ZN(y[88]) );
  OR2_X1 U14bar ( .A1(bbar[8]), .A2(abar[5]), .ZN(ybar[88]);
  AND2_X1 U15 ( .A1(b[7]), .A2(a[5]), .ZN(y[87]) );
  OR2_X1 U15bar ( .A1(bbar[7]), .A2(abar[5]), .ZN(ybar[87]);
  AND2_X1 U16 ( .A1(b[6]), .A2(a[5]), .ZN(y[86]) );
  OR2_X1 U16bar ( .A1(bbar[6]), .A2(abar[5]), .ZN(ybar[86]);
  AND2_X1 U17 ( .A1(b[5]), .A2(a[5]), .ZN(y[85]) );
  OR2_X1 U17bar ( .A1(bbar[5]), .A2(abar[5]), .ZN(ybar[85]);
  AND2_X1 U18 ( .A1(b[4]), .A2(a[5]), .ZN(y[84]) );
  OR2_X1 U18bar ( .A1(bbar[4]), .A2(abar[5]), .ZN(ybar[84]);
  AND2_X1 U19 ( .A1(a[5]), .A2(b[3]), .ZN(y[83]) );
  OR2_X1 U19bar ( .A1(abar[5]), .A2(bbar[3]), .ZN(ybar[83]);
  AND2_X1 U20 ( .A1(a[5]), .A2(b[2]), .ZN(y[82]) );
  OR2_X1 U20bar ( .A1(abar[5]), .A2(bbar[2]), .ZN(ybar[82]);
  AND2_X1 U21 ( .A1(a[5]), .A2(b[1]), .ZN(y[81]) );
  OR2_X1 U21bar ( .A1(abar[5]), .A2(bbar[1]), .ZN(ybar[81]);
  AND2_X1 U22 ( .A1(a[5]), .A2(b[0]), .ZN(y[80]) );
  OR2_X1 U22bar ( .A1(abar[5]), .A2(bbar[0]), .ZN(ybar[80]);
  AND2_X1 U23 ( .A1(b[7]), .A2(a[0]), .ZN(y[7]) );
  OR2_X1 U23bar ( .A1(bbar[7]), .A2(abar[0]), .ZN(ybar[7]);
  AND2_X1 U24 ( .A1(a[4]), .A2(b[15]), .ZN(y[79]) );
  OR2_X1 U24bar ( .A1(abar[4]), .A2(bbar[15]), .ZN(ybar[79]);
  AND2_X1 U25 ( .A1(a[4]), .A2(b[14]), .ZN(y[78]) );
  OR2_X1 U25bar ( .A1(abar[4]), .A2(bbar[14]), .ZN(ybar[78]);
  AND2_X1 U26 ( .A1(a[4]), .A2(b[13]), .ZN(y[77]) );
  OR2_X1 U26bar ( .A1(abar[4]), .A2(bbar[13]), .ZN(ybar[77]);
  AND2_X1 U27 ( .A1(a[4]), .A2(b[12]), .ZN(y[76]) );
  OR2_X1 U27bar ( .A1(abar[4]), .A2(bbar[12]), .ZN(ybar[76]);
  AND2_X1 U28 ( .A1(a[4]), .A2(b[11]), .ZN(y[75]) );
  OR2_X1 U28bar ( .A1(abar[4]), .A2(bbar[11]), .ZN(ybar[75]);
  AND2_X1 U29 ( .A1(a[4]), .A2(b[10]), .ZN(y[74]) );
  OR2_X1 U29bar ( .A1(abar[4]), .A2(bbar[10]), .ZN(ybar[74]);
  AND2_X1 U30 ( .A1(a[4]), .A2(b[9]), .ZN(y[73]) );
  OR2_X1 U30bar ( .A1(abar[4]), .A2(bbar[9]), .ZN(ybar[73]);
  AND2_X1 U31 ( .A1(a[4]), .A2(b[8]), .ZN(y[72]) );
  OR2_X1 U31bar ( .A1(abar[4]), .A2(bbar[8]), .ZN(ybar[72]);
  AND2_X1 U32 ( .A1(a[4]), .A2(b[7]), .ZN(y[71]) );
  OR2_X1 U32bar ( .A1(abar[4]), .A2(bbar[7]), .ZN(ybar[71]);
  AND2_X1 U33 ( .A1(a[4]), .A2(b[6]), .ZN(y[70]) );
  OR2_X1 U33bar ( .A1(abar[4]), .A2(bbar[6]), .ZN(ybar[70]);
  AND2_X1 U34 ( .A1(b[6]), .A2(a[0]), .ZN(y[6]) );
  OR2_X1 U34bar ( .A1(bbar[6]), .A2(abar[0]), .ZN(ybar[6]);
  AND2_X1 U35 ( .A1(a[4]), .A2(b[5]), .ZN(y[69]) );
  OR2_X1 U35bar ( .A1(abar[4]), .A2(bbar[5]), .ZN(ybar[69]);
  AND2_X1 U36 ( .A1(a[4]), .A2(b[4]), .ZN(y[68]) );
  OR2_X1 U36bar ( .A1(abar[4]), .A2(bbar[4]), .ZN(ybar[68]);
  AND2_X1 U37 ( .A1(a[4]), .A2(b[3]), .ZN(y[67]) );
  OR2_X1 U37bar ( .A1(abar[4]), .A2(bbar[3]), .ZN(ybar[67]);
  AND2_X1 U38 ( .A1(a[4]), .A2(b[2]), .ZN(y[66]) );
  OR2_X1 U38bar ( .A1(abar[4]), .A2(bbar[2]), .ZN(ybar[66]);
  AND2_X1 U39 ( .A1(a[4]), .A2(b[1]), .ZN(y[65]) );
  OR2_X1 U39bar ( .A1(abar[4]), .A2(bbar[1]), .ZN(ybar[65]);
  AND2_X1 U40 ( .A1(a[4]), .A2(b[0]), .ZN(y[64]) );
  OR2_X1 U40bar ( .A1(abar[4]), .A2(bbar[0]), .ZN(ybar[64]);
  AND2_X1 U41 ( .A1(a[3]), .A2(b[15]), .ZN(y[63]) );
  OR2_X1 U41bar ( .A1(abar[3]), .A2(bbar[15]), .ZN(ybar[63]);
  AND2_X1 U42 ( .A1(a[3]), .A2(b[14]), .ZN(y[62]) );
  OR2_X1 U42bar ( .A1(abar[3]), .A2(bbar[14]), .ZN(ybar[62]);
  AND2_X1 U43 ( .A1(a[3]), .A2(b[13]), .ZN(y[61]) );
  OR2_X1 U43bar ( .A1(abar[3]), .A2(bbar[13]), .ZN(ybar[61]);
  AND2_X1 U44 ( .A1(a[3]), .A2(b[12]), .ZN(y[60]) );
  OR2_X1 U44bar ( .A1(abar[3]), .A2(bbar[12]), .ZN(ybar[60]);
  AND2_X1 U45 ( .A1(b[5]), .A2(a[0]), .ZN(y[5]) );
  OR2_X1 U45bar ( .A1(bbar[5]), .A2(abar[0]), .ZN(ybar[5]);
  AND2_X1 U46 ( .A1(a[3]), .A2(b[11]), .ZN(y[59]) );
  OR2_X1 U46bar ( .A1(abar[3]), .A2(bbar[11]), .ZN(ybar[59]);
  AND2_X1 U47 ( .A1(a[3]), .A2(b[10]), .ZN(y[58]) );
  OR2_X1 U47bar ( .A1(abar[3]), .A2(bbar[10]), .ZN(ybar[58]);
  AND2_X1 U48 ( .A1(a[3]), .A2(b[9]), .ZN(y[57]) );
  OR2_X1 U48bar ( .A1(abar[3]), .A2(bbar[9]), .ZN(ybar[57]);
  AND2_X1 U49 ( .A1(a[3]), .A2(b[8]), .ZN(y[56]) );
  OR2_X1 U49bar ( .A1(abar[3]), .A2(bbar[8]), .ZN(ybar[56]);
  AND2_X1 U50 ( .A1(a[3]), .A2(b[7]), .ZN(y[55]) );
  OR2_X1 U50bar ( .A1(abar[3]), .A2(bbar[7]), .ZN(ybar[55]);
  AND2_X1 U51 ( .A1(a[3]), .A2(b[6]), .ZN(y[54]) );
  OR2_X1 U51bar ( .A1(abar[3]), .A2(bbar[6]), .ZN(ybar[54]);
  AND2_X1 U52 ( .A1(a[3]), .A2(b[5]), .ZN(y[53]) );
  OR2_X1 U52bar ( .A1(abar[3]), .A2(bbar[5]), .ZN(ybar[53]);
  AND2_X1 U53 ( .A1(a[3]), .A2(b[4]), .ZN(y[52]) );
  OR2_X1 U53bar ( .A1(abar[3]), .A2(bbar[4]), .ZN(ybar[52]);
  AND2_X1 U54 ( .A1(a[3]), .A2(b[3]), .ZN(y[51]) );
  OR2_X1 U54bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[51]);
  AND2_X1 U55 ( .A1(a[3]), .A2(b[2]), .ZN(y[50]) );
  OR2_X1 U55bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[50]);
  AND2_X1 U56 ( .A1(b[4]), .A2(a[0]), .ZN(y[4]) );
  OR2_X1 U56bar ( .A1(bbar[4]), .A2(abar[0]), .ZN(ybar[4]);
  AND2_X1 U57 ( .A1(a[3]), .A2(b[1]), .ZN(y[49]) );
  OR2_X1 U57bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[49]);
  AND2_X1 U58 ( .A1(a[3]), .A2(b[0]), .ZN(y[48]) );
  OR2_X1 U58bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[48]);
  AND2_X1 U59 ( .A1(a[2]), .A2(b[15]), .ZN(y[47]) );
  OR2_X1 U59bar ( .A1(abar[2]), .A2(bbar[15]), .ZN(ybar[47]);
  AND2_X1 U60 ( .A1(a[2]), .A2(b[14]), .ZN(y[46]) );
  OR2_X1 U60bar ( .A1(abar[2]), .A2(bbar[14]), .ZN(ybar[46]);
  AND2_X1 U61 ( .A1(a[2]), .A2(b[13]), .ZN(y[45]) );
  OR2_X1 U61bar ( .A1(abar[2]), .A2(bbar[13]), .ZN(ybar[45]);
  AND2_X1 U62 ( .A1(a[2]), .A2(b[12]), .ZN(y[44]) );
  OR2_X1 U62bar ( .A1(abar[2]), .A2(bbar[12]), .ZN(ybar[44]);
  AND2_X1 U63 ( .A1(a[2]), .A2(b[11]), .ZN(y[43]) );
  OR2_X1 U63bar ( .A1(abar[2]), .A2(bbar[11]), .ZN(ybar[43]);
  AND2_X1 U64 ( .A1(a[2]), .A2(b[10]), .ZN(y[42]) );
  OR2_X1 U64bar ( .A1(abar[2]), .A2(bbar[10]), .ZN(ybar[42]);
  AND2_X1 U65 ( .A1(a[2]), .A2(b[9]), .ZN(y[41]) );
  OR2_X1 U65bar ( .A1(abar[2]), .A2(bbar[9]), .ZN(ybar[41]);
  AND2_X1 U66 ( .A1(a[2]), .A2(b[8]), .ZN(y[40]) );
  OR2_X1 U66bar ( .A1(abar[2]), .A2(bbar[8]), .ZN(ybar[40]);
  AND2_X1 U67 ( .A1(b[3]), .A2(a[0]), .ZN(y[3]) );
  OR2_X1 U67bar ( .A1(bbar[3]), .A2(abar[0]), .ZN(ybar[3]);
  AND2_X1 U68 ( .A1(a[2]), .A2(b[7]), .ZN(y[39]) );
  OR2_X1 U68bar ( .A1(abar[2]), .A2(bbar[7]), .ZN(ybar[39]);
  AND2_X1 U69 ( .A1(a[2]), .A2(b[6]), .ZN(y[38]) );
  OR2_X1 U69bar ( .A1(abar[2]), .A2(bbar[6]), .ZN(ybar[38]);
  AND2_X1 U70 ( .A1(a[2]), .A2(b[5]), .ZN(y[37]) );
  OR2_X1 U70bar ( .A1(abar[2]), .A2(bbar[5]), .ZN(ybar[37]);
  AND2_X1 U71 ( .A1(a[2]), .A2(b[4]), .ZN(y[36]) );
  OR2_X1 U71bar ( .A1(abar[2]), .A2(bbar[4]), .ZN(ybar[36]);
  AND2_X1 U72 ( .A1(a[2]), .A2(b[3]), .ZN(y[35]) );
  OR2_X1 U72bar ( .A1(abar[2]), .A2(bbar[3]), .ZN(ybar[35]);
  AND2_X1 U73 ( .A1(a[2]), .A2(b[2]), .ZN(y[34]) );
  OR2_X1 U73bar ( .A1(abar[2]), .A2(bbar[2]), .ZN(ybar[34]);
  AND2_X1 U74 ( .A1(a[2]), .A2(b[1]), .ZN(y[33]) );
  OR2_X1 U74bar ( .A1(abar[2]), .A2(bbar[1]), .ZN(ybar[33]);
  AND2_X1 U75 ( .A1(a[2]), .A2(b[0]), .ZN(y[32]) );
  OR2_X1 U75bar ( .A1(abar[2]), .A2(bbar[0]), .ZN(ybar[32]);
  AND2_X1 U76 ( .A1(a[1]), .A2(b[15]), .ZN(y[31]) );
  OR2_X1 U76bar ( .A1(abar[1]), .A2(bbar[15]), .ZN(ybar[31]);
  AND2_X1 U77 ( .A1(a[1]), .A2(b[14]), .ZN(y[30]) );
  OR2_X1 U77bar ( .A1(abar[1]), .A2(bbar[14]), .ZN(ybar[30]);
  AND2_X1 U78 ( .A1(b[2]), .A2(a[0]), .ZN(y[2]) );
  OR2_X1 U78bar ( .A1(bbar[2]), .A2(abar[0]), .ZN(ybar[2]);
  AND2_X1 U79 ( .A1(a[1]), .A2(b[13]), .ZN(y[29]) );
  OR2_X1 U79bar ( .A1(abar[1]), .A2(bbar[13]), .ZN(ybar[29]);
  AND2_X1 U80 ( .A1(a[1]), .A2(b[12]), .ZN(y[28]) );
  OR2_X1 U80bar ( .A1(abar[1]), .A2(bbar[12]), .ZN(ybar[28]);
  AND2_X1 U81 ( .A1(a[1]), .A2(b[11]), .ZN(y[27]) );
  OR2_X1 U81bar ( .A1(abar[1]), .A2(bbar[11]), .ZN(ybar[27]);
  AND2_X1 U82 ( .A1(a[1]), .A2(b[10]), .ZN(y[26]) );
  OR2_X1 U82bar ( .A1(abar[1]), .A2(bbar[10]), .ZN(ybar[26]);
  AND2_X1 U83 ( .A1(a[1]), .A2(b[9]), .ZN(y[25]) );
  OR2_X1 U83bar ( .A1(abar[1]), .A2(bbar[9]), .ZN(ybar[25]);
  AND2_X1 U84 ( .A1(a[15]), .A2(b[15]), .ZN(y[255]) );
  OR2_X1 U84bar ( .A1(abar[15]), .A2(bbar[15]), .ZN(ybar[255]);
  AND2_X1 U85 ( .A1(a[15]), .A2(b[14]), .ZN(y[254]) );
  OR2_X1 U85bar ( .A1(abar[15]), .A2(bbar[14]), .ZN(ybar[254]);
  AND2_X1 U86 ( .A1(a[15]), .A2(b[13]), .ZN(y[253]) );
  OR2_X1 U86bar ( .A1(abar[15]), .A2(bbar[13]), .ZN(ybar[253]);
  AND2_X1 U87 ( .A1(a[15]), .A2(b[12]), .ZN(y[252]) );
  OR2_X1 U87bar ( .A1(abar[15]), .A2(bbar[12]), .ZN(ybar[252]);
  AND2_X1 U88 ( .A1(a[15]), .A2(b[11]), .ZN(y[251]) );
  OR2_X1 U88bar ( .A1(abar[15]), .A2(bbar[11]), .ZN(ybar[251]);
  AND2_X1 U89 ( .A1(a[15]), .A2(b[10]), .ZN(y[250]) );
  OR2_X1 U89bar ( .A1(abar[15]), .A2(bbar[10]), .ZN(ybar[250]);
  AND2_X1 U90 ( .A1(a[1]), .A2(b[8]), .ZN(y[24]) );
  OR2_X1 U90bar ( .A1(abar[1]), .A2(bbar[8]), .ZN(ybar[24]);
  AND2_X1 U91 ( .A1(a[15]), .A2(b[9]), .ZN(y[249]) );
  OR2_X1 U91bar ( .A1(abar[15]), .A2(bbar[9]), .ZN(ybar[249]);
  AND2_X1 U92 ( .A1(a[15]), .A2(b[8]), .ZN(y[248]) );
  OR2_X1 U92bar ( .A1(abar[15]), .A2(bbar[8]), .ZN(ybar[248]);
  AND2_X1 U93 ( .A1(a[15]), .A2(b[7]), .ZN(y[247]) );
  OR2_X1 U93bar ( .A1(abar[15]), .A2(bbar[7]), .ZN(ybar[247]);
  AND2_X1 U94 ( .A1(a[15]), .A2(b[6]), .ZN(y[246]) );
  OR2_X1 U94bar ( .A1(abar[15]), .A2(bbar[6]), .ZN(ybar[246]);
  AND2_X1 U95 ( .A1(a[15]), .A2(b[5]), .ZN(y[245]) );
  OR2_X1 U95bar ( .A1(abar[15]), .A2(bbar[5]), .ZN(ybar[245]);
  AND2_X1 U96 ( .A1(a[15]), .A2(b[4]), .ZN(y[244]) );
  OR2_X1 U96bar ( .A1(abar[15]), .A2(bbar[4]), .ZN(ybar[244]);
  AND2_X1 U97 ( .A1(a[15]), .A2(b[3]), .ZN(y[243]) );
  OR2_X1 U97bar ( .A1(abar[15]), .A2(bbar[3]), .ZN(ybar[243]);
  AND2_X1 U98 ( .A1(a[15]), .A2(b[2]), .ZN(y[242]) );
  OR2_X1 U98bar ( .A1(abar[15]), .A2(bbar[2]), .ZN(ybar[242]);
  AND2_X1 U99 ( .A1(a[15]), .A2(b[1]), .ZN(y[241]) );
  OR2_X1 U99bar ( .A1(abar[15]), .A2(bbar[1]), .ZN(ybar[241]);
  AND2_X1 U100 ( .A1(a[15]), .A2(b[0]), .ZN(y[240]) );
  OR2_X1 U100bar ( .A1(abar[15]), .A2(bbar[0]), .ZN(ybar[240]);
  AND2_X1 U101 ( .A1(a[1]), .A2(b[7]), .ZN(y[23]) );
  OR2_X1 U101bar ( .A1(abar[1]), .A2(bbar[7]), .ZN(ybar[23]);
  AND2_X1 U102 ( .A1(a[14]), .A2(b[15]), .ZN(y[239]) );
  OR2_X1 U102bar ( .A1(abar[14]), .A2(bbar[15]), .ZN(ybar[239]);
  AND2_X1 U103 ( .A1(a[14]), .A2(b[14]), .ZN(y[238]) );
  OR2_X1 U103bar ( .A1(abar[14]), .A2(bbar[14]), .ZN(ybar[238]);
  AND2_X1 U104 ( .A1(a[14]), .A2(b[13]), .ZN(y[237]) );
  OR2_X1 U104bar ( .A1(abar[14]), .A2(bbar[13]), .ZN(ybar[237]);
  AND2_X1 U105 ( .A1(a[14]), .A2(b[12]), .ZN(y[236]) );
  OR2_X1 U105bar ( .A1(abar[14]), .A2(bbar[12]), .ZN(ybar[236]);
  AND2_X1 U106 ( .A1(a[14]), .A2(b[11]), .ZN(y[235]) );
  OR2_X1 U106bar ( .A1(abar[14]), .A2(bbar[11]), .ZN(ybar[235]);
  AND2_X1 U107 ( .A1(a[14]), .A2(b[10]), .ZN(y[234]) );
  OR2_X1 U107bar ( .A1(abar[14]), .A2(bbar[10]), .ZN(ybar[234]);
  AND2_X1 U108 ( .A1(a[14]), .A2(b[9]), .ZN(y[233]) );
  OR2_X1 U108bar ( .A1(abar[14]), .A2(bbar[9]), .ZN(ybar[233]);
  AND2_X1 U109 ( .A1(a[14]), .A2(b[8]), .ZN(y[232]) );
  OR2_X1 U109bar ( .A1(abar[14]), .A2(bbar[8]), .ZN(ybar[232]);
  AND2_X1 U110 ( .A1(a[14]), .A2(b[7]), .ZN(y[231]) );
  OR2_X1 U110bar ( .A1(abar[14]), .A2(bbar[7]), .ZN(ybar[231]);
  AND2_X1 U111 ( .A1(a[14]), .A2(b[6]), .ZN(y[230]) );
  OR2_X1 U111bar ( .A1(abar[14]), .A2(bbar[6]), .ZN(ybar[230]);
  AND2_X1 U112 ( .A1(a[1]), .A2(b[6]), .ZN(y[22]) );
  OR2_X1 U112bar ( .A1(abar[1]), .A2(bbar[6]), .ZN(ybar[22]);
  AND2_X1 U113 ( .A1(a[14]), .A2(b[5]), .ZN(y[229]) );
  OR2_X1 U113bar ( .A1(abar[14]), .A2(bbar[5]), .ZN(ybar[229]);
  AND2_X1 U114 ( .A1(a[14]), .A2(b[4]), .ZN(y[228]) );
  OR2_X1 U114bar ( .A1(abar[14]), .A2(bbar[4]), .ZN(ybar[228]);
  AND2_X1 U115 ( .A1(a[14]), .A2(b[3]), .ZN(y[227]) );
  OR2_X1 U115bar ( .A1(abar[14]), .A2(bbar[3]), .ZN(ybar[227]);
  AND2_X1 U116 ( .A1(a[14]), .A2(b[2]), .ZN(y[226]) );
  OR2_X1 U116bar ( .A1(abar[14]), .A2(bbar[2]), .ZN(ybar[226]);
  AND2_X1 U117 ( .A1(a[14]), .A2(b[1]), .ZN(y[225]) );
  OR2_X1 U117bar ( .A1(abar[14]), .A2(bbar[1]), .ZN(ybar[225]);
  AND2_X1 U118 ( .A1(a[14]), .A2(b[0]), .ZN(y[224]) );
  OR2_X1 U118bar ( .A1(abar[14]), .A2(bbar[0]), .ZN(ybar[224]);
  AND2_X1 U119 ( .A1(a[13]), .A2(b[15]), .ZN(y[223]) );
  OR2_X1 U119bar ( .A1(abar[13]), .A2(bbar[15]), .ZN(ybar[223]);
  AND2_X1 U120 ( .A1(a[13]), .A2(b[14]), .ZN(y[222]) );
  OR2_X1 U120bar ( .A1(abar[13]), .A2(bbar[14]), .ZN(ybar[222]);
  AND2_X1 U121 ( .A1(a[13]), .A2(b[13]), .ZN(y[221]) );
  OR2_X1 U121bar ( .A1(abar[13]), .A2(bbar[13]), .ZN(ybar[221]);
  AND2_X1 U122 ( .A1(a[13]), .A2(b[12]), .ZN(y[220]) );
  OR2_X1 U122bar ( .A1(abar[13]), .A2(bbar[12]), .ZN(ybar[220]);
  AND2_X1 U123 ( .A1(a[1]), .A2(b[5]), .ZN(y[21]) );
  OR2_X1 U123bar ( .A1(abar[1]), .A2(bbar[5]), .ZN(ybar[21]);
  AND2_X1 U124 ( .A1(a[13]), .A2(b[11]), .ZN(y[219]) );
  OR2_X1 U124bar ( .A1(abar[13]), .A2(bbar[11]), .ZN(ybar[219]);
  AND2_X1 U125 ( .A1(a[13]), .A2(b[10]), .ZN(y[218]) );
  OR2_X1 U125bar ( .A1(abar[13]), .A2(bbar[10]), .ZN(ybar[218]);
  AND2_X1 U126 ( .A1(a[13]), .A2(b[9]), .ZN(y[217]) );
  OR2_X1 U126bar ( .A1(abar[13]), .A2(bbar[9]), .ZN(ybar[217]);
  AND2_X1 U127 ( .A1(a[13]), .A2(b[8]), .ZN(y[216]) );
  OR2_X1 U127bar ( .A1(abar[13]), .A2(bbar[8]), .ZN(ybar[216]);
  AND2_X1 U128 ( .A1(a[13]), .A2(b[7]), .ZN(y[215]) );
  OR2_X1 U128bar ( .A1(abar[13]), .A2(bbar[7]), .ZN(ybar[215]);
  AND2_X1 U129 ( .A1(a[13]), .A2(b[6]), .ZN(y[214]) );
  OR2_X1 U129bar ( .A1(abar[13]), .A2(bbar[6]), .ZN(ybar[214]);
  AND2_X1 U130 ( .A1(a[13]), .A2(b[5]), .ZN(y[213]) );
  OR2_X1 U130bar ( .A1(abar[13]), .A2(bbar[5]), .ZN(ybar[213]);
  AND2_X1 U131 ( .A1(a[13]), .A2(b[4]), .ZN(y[212]) );
  OR2_X1 U131bar ( .A1(abar[13]), .A2(bbar[4]), .ZN(ybar[212]);
  AND2_X1 U132 ( .A1(a[13]), .A2(b[3]), .ZN(y[211]) );
  OR2_X1 U132bar ( .A1(abar[13]), .A2(bbar[3]), .ZN(ybar[211]);
  AND2_X1 U133 ( .A1(a[13]), .A2(b[2]), .ZN(y[210]) );
  OR2_X1 U133bar ( .A1(abar[13]), .A2(bbar[2]), .ZN(ybar[210]);
  AND2_X1 U134 ( .A1(a[1]), .A2(b[4]), .ZN(y[20]) );
  OR2_X1 U134bar ( .A1(abar[1]), .A2(bbar[4]), .ZN(ybar[20]);
  AND2_X1 U135 ( .A1(a[13]), .A2(b[1]), .ZN(y[209]) );
  OR2_X1 U135bar ( .A1(abar[13]), .A2(bbar[1]), .ZN(ybar[209]);
  AND2_X1 U136 ( .A1(a[13]), .A2(b[0]), .ZN(y[208]) );
  OR2_X1 U136bar ( .A1(abar[13]), .A2(bbar[0]), .ZN(ybar[208]);
  AND2_X1 U137 ( .A1(a[12]), .A2(b[15]), .ZN(y[207]) );
  OR2_X1 U137bar ( .A1(abar[12]), .A2(bbar[15]), .ZN(ybar[207]);
  AND2_X1 U138 ( .A1(a[12]), .A2(b[14]), .ZN(y[206]) );
  OR2_X1 U138bar ( .A1(abar[12]), .A2(bbar[14]), .ZN(ybar[206]);
  AND2_X1 U139 ( .A1(a[12]), .A2(b[13]), .ZN(y[205]) );
  OR2_X1 U139bar ( .A1(abar[12]), .A2(bbar[13]), .ZN(ybar[205]);
  AND2_X1 U140 ( .A1(a[12]), .A2(b[12]), .ZN(y[204]) );
  OR2_X1 U140bar ( .A1(abar[12]), .A2(bbar[12]), .ZN(ybar[204]);
  AND2_X1 U141 ( .A1(a[12]), .A2(b[11]), .ZN(y[203]) );
  OR2_X1 U141bar ( .A1(abar[12]), .A2(bbar[11]), .ZN(ybar[203]);
  AND2_X1 U142 ( .A1(a[12]), .A2(b[10]), .ZN(y[202]) );
  OR2_X1 U142bar ( .A1(abar[12]), .A2(bbar[10]), .ZN(ybar[202]);
  AND2_X1 U143 ( .A1(a[12]), .A2(b[9]), .ZN(y[201]) );
  OR2_X1 U143bar ( .A1(abar[12]), .A2(bbar[9]), .ZN(ybar[201]);
  AND2_X1 U144 ( .A1(a[12]), .A2(b[8]), .ZN(y[200]) );
  OR2_X1 U144bar ( .A1(abar[12]), .A2(bbar[8]), .ZN(ybar[200]);
  AND2_X1 U145 ( .A1(b[1]), .A2(a[0]), .ZN(y[1]) );
  OR2_X1 U145bar ( .A1(bbar[1]), .A2(abar[0]), .ZN(ybar[1]);
  AND2_X1 U146 ( .A1(a[1]), .A2(b[3]), .ZN(y[19]) );
  OR2_X1 U146bar ( .A1(abar[1]), .A2(bbar[3]), .ZN(ybar[19]);
  AND2_X1 U147 ( .A1(a[12]), .A2(b[7]), .ZN(y[199]) );
  OR2_X1 U147bar ( .A1(abar[12]), .A2(bbar[7]), .ZN(ybar[199]);
  AND2_X1 U148 ( .A1(a[12]), .A2(b[6]), .ZN(y[198]) );
  OR2_X1 U148bar ( .A1(abar[12]), .A2(bbar[6]), .ZN(ybar[198]);
  AND2_X1 U149 ( .A1(a[12]), .A2(b[5]), .ZN(y[197]) );
  OR2_X1 U149bar ( .A1(abar[12]), .A2(bbar[5]), .ZN(ybar[197]);
  AND2_X1 U150 ( .A1(a[12]), .A2(b[4]), .ZN(y[196]) );
  OR2_X1 U150bar ( .A1(abar[12]), .A2(bbar[4]), .ZN(ybar[196]);
  AND2_X1 U151 ( .A1(a[12]), .A2(b[3]), .ZN(y[195]) );
  OR2_X1 U151bar ( .A1(abar[12]), .A2(bbar[3]), .ZN(ybar[195]);
  AND2_X1 U152 ( .A1(a[12]), .A2(b[2]), .ZN(y[194]) );
  OR2_X1 U152bar ( .A1(abar[12]), .A2(bbar[2]), .ZN(ybar[194]);
  AND2_X1 U153 ( .A1(a[12]), .A2(b[1]), .ZN(y[193]) );
  OR2_X1 U153bar ( .A1(abar[12]), .A2(bbar[1]), .ZN(ybar[193]);
  AND2_X1 U154 ( .A1(a[12]), .A2(b[0]), .ZN(y[192]) );
  OR2_X1 U154bar ( .A1(abar[12]), .A2(bbar[0]), .ZN(ybar[192]);
  AND2_X1 U155 ( .A1(a[11]), .A2(b[15]), .ZN(y[191]) );
  OR2_X1 U155bar ( .A1(abar[11]), .A2(bbar[15]), .ZN(ybar[191]);
  AND2_X1 U156 ( .A1(a[11]), .A2(b[14]), .ZN(y[190]) );
  OR2_X1 U156bar ( .A1(abar[11]), .A2(bbar[14]), .ZN(ybar[190]);
  AND2_X1 U157 ( .A1(a[1]), .A2(b[2]), .ZN(y[18]) );
  OR2_X1 U157bar ( .A1(abar[1]), .A2(bbar[2]), .ZN(ybar[18]);
  AND2_X1 U158 ( .A1(a[11]), .A2(b[13]), .ZN(y[189]) );
  OR2_X1 U158bar ( .A1(abar[11]), .A2(bbar[13]), .ZN(ybar[189]);
  AND2_X1 U159 ( .A1(a[11]), .A2(b[12]), .ZN(y[188]) );
  OR2_X1 U159bar ( .A1(abar[11]), .A2(bbar[12]), .ZN(ybar[188]);
  AND2_X1 U160 ( .A1(a[11]), .A2(b[11]), .ZN(y[187]) );
  OR2_X1 U160bar ( .A1(abar[11]), .A2(bbar[11]), .ZN(ybar[187]);
  AND2_X1 U161 ( .A1(a[11]), .A2(b[10]), .ZN(y[186]) );
  OR2_X1 U161bar ( .A1(abar[11]), .A2(bbar[10]), .ZN(ybar[186]);
  AND2_X1 U162 ( .A1(a[11]), .A2(b[9]), .ZN(y[185]) );
  OR2_X1 U162bar ( .A1(abar[11]), .A2(bbar[9]), .ZN(ybar[185]);
  AND2_X1 U163 ( .A1(a[11]), .A2(b[8]), .ZN(y[184]) );
  OR2_X1 U163bar ( .A1(abar[11]), .A2(bbar[8]), .ZN(ybar[184]);
  AND2_X1 U164 ( .A1(a[11]), .A2(b[7]), .ZN(y[183]) );
  OR2_X1 U164bar ( .A1(abar[11]), .A2(bbar[7]), .ZN(ybar[183]);
  AND2_X1 U165 ( .A1(a[11]), .A2(b[6]), .ZN(y[182]) );
  OR2_X1 U165bar ( .A1(abar[11]), .A2(bbar[6]), .ZN(ybar[182]);
  AND2_X1 U166 ( .A1(a[11]), .A2(b[5]), .ZN(y[181]) );
  OR2_X1 U166bar ( .A1(abar[11]), .A2(bbar[5]), .ZN(ybar[181]);
  AND2_X1 U167 ( .A1(a[11]), .A2(b[4]), .ZN(y[180]) );
  OR2_X1 U167bar ( .A1(abar[11]), .A2(bbar[4]), .ZN(ybar[180]);
  AND2_X1 U168 ( .A1(a[1]), .A2(b[1]), .ZN(y[17]) );
  OR2_X1 U168bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[17]);
  AND2_X1 U169 ( .A1(a[11]), .A2(b[3]), .ZN(y[179]) );
  OR2_X1 U169bar ( .A1(abar[11]), .A2(bbar[3]), .ZN(ybar[179]);
  AND2_X1 U170 ( .A1(a[11]), .A2(b[2]), .ZN(y[178]) );
  OR2_X1 U170bar ( .A1(abar[11]), .A2(bbar[2]), .ZN(ybar[178]);
  AND2_X1 U171 ( .A1(a[11]), .A2(b[1]), .ZN(y[177]) );
  OR2_X1 U171bar ( .A1(abar[11]), .A2(bbar[1]), .ZN(ybar[177]);
  AND2_X1 U172 ( .A1(a[11]), .A2(b[0]), .ZN(y[176]) );
  OR2_X1 U172bar ( .A1(abar[11]), .A2(bbar[0]), .ZN(ybar[176]);
  AND2_X1 U173 ( .A1(a[10]), .A2(b[15]), .ZN(y[175]) );
  OR2_X1 U173bar ( .A1(abar[10]), .A2(bbar[15]), .ZN(ybar[175]);
  AND2_X1 U174 ( .A1(a[10]), .A2(b[14]), .ZN(y[174]) );
  OR2_X1 U174bar ( .A1(abar[10]), .A2(bbar[14]), .ZN(ybar[174]);
  AND2_X1 U175 ( .A1(a[10]), .A2(b[13]), .ZN(y[173]) );
  OR2_X1 U175bar ( .A1(abar[10]), .A2(bbar[13]), .ZN(ybar[173]);
  AND2_X1 U176 ( .A1(a[10]), .A2(b[12]), .ZN(y[172]) );
  OR2_X1 U176bar ( .A1(abar[10]), .A2(bbar[12]), .ZN(ybar[172]);
  AND2_X1 U177 ( .A1(a[10]), .A2(b[11]), .ZN(y[171]) );
  OR2_X1 U177bar ( .A1(abar[10]), .A2(bbar[11]), .ZN(ybar[171]);
  AND2_X1 U178 ( .A1(a[10]), .A2(b[10]), .ZN(y[170]) );
  OR2_X1 U178bar ( .A1(abar[10]), .A2(bbar[10]), .ZN(ybar[170]);
  AND2_X1 U179 ( .A1(a[1]), .A2(b[0]), .ZN(y[16]) );
  OR2_X1 U179bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[16]);
  AND2_X1 U180 ( .A1(a[10]), .A2(b[9]), .ZN(y[169]) );
  OR2_X1 U180bar ( .A1(abar[10]), .A2(bbar[9]), .ZN(ybar[169]);
  AND2_X1 U181 ( .A1(a[10]), .A2(b[8]), .ZN(y[168]) );
  OR2_X1 U181bar ( .A1(abar[10]), .A2(bbar[8]), .ZN(ybar[168]);
  AND2_X1 U182 ( .A1(a[10]), .A2(b[7]), .ZN(y[167]) );
  OR2_X1 U182bar ( .A1(abar[10]), .A2(bbar[7]), .ZN(ybar[167]);
  AND2_X1 U183 ( .A1(a[10]), .A2(b[6]), .ZN(y[166]) );
  OR2_X1 U183bar ( .A1(abar[10]), .A2(bbar[6]), .ZN(ybar[166]);
  AND2_X1 U184 ( .A1(a[10]), .A2(b[5]), .ZN(y[165]) );
  OR2_X1 U184bar ( .A1(abar[10]), .A2(bbar[5]), .ZN(ybar[165]);
  AND2_X1 U185 ( .A1(a[10]), .A2(b[4]), .ZN(y[164]) );
  OR2_X1 U185bar ( .A1(abar[10]), .A2(bbar[4]), .ZN(ybar[164]);
  AND2_X1 U186 ( .A1(a[10]), .A2(b[3]), .ZN(y[163]) );
  OR2_X1 U186bar ( .A1(abar[10]), .A2(bbar[3]), .ZN(ybar[163]);
  AND2_X1 U187 ( .A1(a[10]), .A2(b[2]), .ZN(y[162]) );
  OR2_X1 U187bar ( .A1(abar[10]), .A2(bbar[2]), .ZN(ybar[162]);
  AND2_X1 U188 ( .A1(a[10]), .A2(b[1]), .ZN(y[161]) );
  OR2_X1 U188bar ( .A1(abar[10]), .A2(bbar[1]), .ZN(ybar[161]);
  AND2_X1 U189 ( .A1(a[10]), .A2(b[0]), .ZN(y[160]) );
  OR2_X1 U189bar ( .A1(abar[10]), .A2(bbar[0]), .ZN(ybar[160]);
  AND2_X1 U190 ( .A1(b[15]), .A2(a[0]), .ZN(y[15]) );
  OR2_X1 U190bar ( .A1(bbar[15]), .A2(abar[0]), .ZN(ybar[15]);
  AND2_X1 U191 ( .A1(a[9]), .A2(b[15]), .ZN(y[159]) );
  OR2_X1 U191bar ( .A1(abar[9]), .A2(bbar[15]), .ZN(ybar[159]);
  AND2_X1 U192 ( .A1(a[9]), .A2(b[14]), .ZN(y[158]) );
  OR2_X1 U192bar ( .A1(abar[9]), .A2(bbar[14]), .ZN(ybar[158]);
  AND2_X1 U193 ( .A1(a[9]), .A2(b[13]), .ZN(y[157]) );
  OR2_X1 U193bar ( .A1(abar[9]), .A2(bbar[13]), .ZN(ybar[157]);
  AND2_X1 U194 ( .A1(a[9]), .A2(b[12]), .ZN(y[156]) );
  OR2_X1 U194bar ( .A1(abar[9]), .A2(bbar[12]), .ZN(ybar[156]);
  AND2_X1 U195 ( .A1(a[9]), .A2(b[11]), .ZN(y[155]) );
  OR2_X1 U195bar ( .A1(abar[9]), .A2(bbar[11]), .ZN(ybar[155]);
  AND2_X1 U196 ( .A1(a[9]), .A2(b[10]), .ZN(y[154]) );
  OR2_X1 U196bar ( .A1(abar[9]), .A2(bbar[10]), .ZN(ybar[154]);
  AND2_X1 U197 ( .A1(a[9]), .A2(b[9]), .ZN(y[153]) );
  OR2_X1 U197bar ( .A1(abar[9]), .A2(bbar[9]), .ZN(ybar[153]);
  AND2_X1 U198 ( .A1(a[9]), .A2(b[8]), .ZN(y[152]) );
  OR2_X1 U198bar ( .A1(abar[9]), .A2(bbar[8]), .ZN(ybar[152]);
  AND2_X1 U199 ( .A1(a[9]), .A2(b[7]), .ZN(y[151]) );
  OR2_X1 U199bar ( .A1(abar[9]), .A2(bbar[7]), .ZN(ybar[151]);
  AND2_X1 U200 ( .A1(a[9]), .A2(b[6]), .ZN(y[150]) );
  OR2_X1 U200bar ( .A1(abar[9]), .A2(bbar[6]), .ZN(ybar[150]);
  AND2_X1 U201 ( .A1(b[14]), .A2(a[0]), .ZN(y[14]) );
  OR2_X1 U201bar ( .A1(bbar[14]), .A2(abar[0]), .ZN(ybar[14]);
  AND2_X1 U202 ( .A1(a[9]), .A2(b[5]), .ZN(y[149]) );
  OR2_X1 U202bar ( .A1(abar[9]), .A2(bbar[5]), .ZN(ybar[149]);
  AND2_X1 U203 ( .A1(a[9]), .A2(b[4]), .ZN(y[148]) );
  OR2_X1 U203bar ( .A1(abar[9]), .A2(bbar[4]), .ZN(ybar[148]);
  AND2_X1 U204 ( .A1(a[9]), .A2(b[3]), .ZN(y[147]) );
  OR2_X1 U204bar ( .A1(abar[9]), .A2(bbar[3]), .ZN(ybar[147]);
  AND2_X1 U205 ( .A1(a[9]), .A2(b[2]), .ZN(y[146]) );
  OR2_X1 U205bar ( .A1(abar[9]), .A2(bbar[2]), .ZN(ybar[146]);
  AND2_X1 U206 ( .A1(a[9]), .A2(b[1]), .ZN(y[145]) );
  OR2_X1 U206bar ( .A1(abar[9]), .A2(bbar[1]), .ZN(ybar[145]);
  AND2_X1 U207 ( .A1(a[9]), .A2(b[0]), .ZN(y[144]) );
  OR2_X1 U207bar ( .A1(abar[9]), .A2(bbar[0]), .ZN(ybar[144]);
  AND2_X1 U208 ( .A1(a[8]), .A2(b[15]), .ZN(y[143]) );
  OR2_X1 U208bar ( .A1(abar[8]), .A2(bbar[15]), .ZN(ybar[143]);
  AND2_X1 U209 ( .A1(a[8]), .A2(b[14]), .ZN(y[142]) );
  OR2_X1 U209bar ( .A1(abar[8]), .A2(bbar[14]), .ZN(ybar[142]);
  AND2_X1 U210 ( .A1(a[8]), .A2(b[13]), .ZN(y[141]) );
  OR2_X1 U210bar ( .A1(abar[8]), .A2(bbar[13]), .ZN(ybar[141]);
  AND2_X1 U211 ( .A1(a[8]), .A2(b[12]), .ZN(y[140]) );
  OR2_X1 U211bar ( .A1(abar[8]), .A2(bbar[12]), .ZN(ybar[140]);
  AND2_X1 U212 ( .A1(b[13]), .A2(a[0]), .ZN(y[13]) );
  OR2_X1 U212bar ( .A1(bbar[13]), .A2(abar[0]), .ZN(ybar[13]);
  AND2_X1 U213 ( .A1(a[8]), .A2(b[11]), .ZN(y[139]) );
  OR2_X1 U213bar ( .A1(abar[8]), .A2(bbar[11]), .ZN(ybar[139]);
  AND2_X1 U214 ( .A1(a[8]), .A2(b[10]), .ZN(y[138]) );
  OR2_X1 U214bar ( .A1(abar[8]), .A2(bbar[10]), .ZN(ybar[138]);
  AND2_X1 U215 ( .A1(a[8]), .A2(b[9]), .ZN(y[137]) );
  OR2_X1 U215bar ( .A1(abar[8]), .A2(bbar[9]), .ZN(ybar[137]);
  AND2_X1 U216 ( .A1(a[8]), .A2(b[8]), .ZN(y[136]) );
  OR2_X1 U216bar ( .A1(abar[8]), .A2(bbar[8]), .ZN(ybar[136]);
  AND2_X1 U217 ( .A1(a[8]), .A2(b[7]), .ZN(y[135]) );
  OR2_X1 U217bar ( .A1(abar[8]), .A2(bbar[7]), .ZN(ybar[135]);
  AND2_X1 U218 ( .A1(a[8]), .A2(b[6]), .ZN(y[134]) );
  OR2_X1 U218bar ( .A1(abar[8]), .A2(bbar[6]), .ZN(ybar[134]);
  AND2_X1 U219 ( .A1(a[8]), .A2(b[5]), .ZN(y[133]) );
  OR2_X1 U219bar ( .A1(abar[8]), .A2(bbar[5]), .ZN(ybar[133]);
  AND2_X1 U220 ( .A1(a[8]), .A2(b[4]), .ZN(y[132]) );
  OR2_X1 U220bar ( .A1(abar[8]), .A2(bbar[4]), .ZN(ybar[132]);
  AND2_X1 U221 ( .A1(a[8]), .A2(b[3]), .ZN(y[131]) );
  OR2_X1 U221bar ( .A1(abar[8]), .A2(bbar[3]), .ZN(ybar[131]);
  AND2_X1 U222 ( .A1(a[8]), .A2(b[2]), .ZN(y[130]) );
  OR2_X1 U222bar ( .A1(abar[8]), .A2(bbar[2]), .ZN(ybar[130]);
  AND2_X1 U223 ( .A1(b[12]), .A2(a[0]), .ZN(y[12]) );
  OR2_X1 U223bar ( .A1(bbar[12]), .A2(abar[0]), .ZN(ybar[12]);
  AND2_X1 U224 ( .A1(a[8]), .A2(b[1]), .ZN(y[129]) );
  OR2_X1 U224bar ( .A1(abar[8]), .A2(bbar[1]), .ZN(ybar[129]);
  AND2_X1 U225 ( .A1(a[8]), .A2(b[0]), .ZN(y[128]) );
  OR2_X1 U225bar ( .A1(abar[8]), .A2(bbar[0]), .ZN(ybar[128]);
  AND2_X1 U226 ( .A1(a[7]), .A2(b[15]), .ZN(y[127]) );
  OR2_X1 U226bar ( .A1(abar[7]), .A2(bbar[15]), .ZN(ybar[127]);
  AND2_X1 U227 ( .A1(a[7]), .A2(b[14]), .ZN(y[126]) );
  OR2_X1 U227bar ( .A1(abar[7]), .A2(bbar[14]), .ZN(ybar[126]);
  AND2_X1 U228 ( .A1(a[7]), .A2(b[13]), .ZN(y[125]) );
  OR2_X1 U228bar ( .A1(abar[7]), .A2(bbar[13]), .ZN(ybar[125]);
  AND2_X1 U229 ( .A1(a[7]), .A2(b[12]), .ZN(y[124]) );
  OR2_X1 U229bar ( .A1(abar[7]), .A2(bbar[12]), .ZN(ybar[124]);
  AND2_X1 U230 ( .A1(a[7]), .A2(b[11]), .ZN(y[123]) );
  OR2_X1 U230bar ( .A1(abar[7]), .A2(bbar[11]), .ZN(ybar[123]);
  AND2_X1 U231 ( .A1(a[7]), .A2(b[10]), .ZN(y[122]) );
  OR2_X1 U231bar ( .A1(abar[7]), .A2(bbar[10]), .ZN(ybar[122]);
  AND2_X1 U232 ( .A1(a[7]), .A2(b[9]), .ZN(y[121]) );
  OR2_X1 U232bar ( .A1(abar[7]), .A2(bbar[9]), .ZN(ybar[121]);
  AND2_X1 U233 ( .A1(a[7]), .A2(b[8]), .ZN(y[120]) );
  OR2_X1 U233bar ( .A1(abar[7]), .A2(bbar[8]), .ZN(ybar[120]);
  AND2_X1 U234 ( .A1(b[11]), .A2(a[0]), .ZN(y[11]) );
  OR2_X1 U234bar ( .A1(bbar[11]), .A2(abar[0]), .ZN(ybar[11]);
  AND2_X1 U235 ( .A1(a[7]), .A2(b[7]), .ZN(y[119]) );
  OR2_X1 U235bar ( .A1(abar[7]), .A2(bbar[7]), .ZN(ybar[119]);
  AND2_X1 U236 ( .A1(a[7]), .A2(b[6]), .ZN(y[118]) );
  OR2_X1 U236bar ( .A1(abar[7]), .A2(bbar[6]), .ZN(ybar[118]);
  AND2_X1 U237 ( .A1(a[7]), .A2(b[5]), .ZN(y[117]) );
  OR2_X1 U237bar ( .A1(abar[7]), .A2(bbar[5]), .ZN(ybar[117]);
  AND2_X1 U238 ( .A1(a[7]), .A2(b[4]), .ZN(y[116]) );
  OR2_X1 U238bar ( .A1(abar[7]), .A2(bbar[4]), .ZN(ybar[116]);
  AND2_X1 U239 ( .A1(a[7]), .A2(b[3]), .ZN(y[115]) );
  OR2_X1 U239bar ( .A1(abar[7]), .A2(bbar[3]), .ZN(ybar[115]);
  AND2_X1 U240 ( .A1(a[7]), .A2(b[2]), .ZN(y[114]) );
  OR2_X1 U240bar ( .A1(abar[7]), .A2(bbar[2]), .ZN(ybar[114]);
  AND2_X1 U241 ( .A1(a[7]), .A2(b[1]), .ZN(y[113]) );
  OR2_X1 U241bar ( .A1(abar[7]), .A2(bbar[1]), .ZN(ybar[113]);
  AND2_X1 U242 ( .A1(a[7]), .A2(b[0]), .ZN(y[112]) );
  OR2_X1 U242bar ( .A1(abar[7]), .A2(bbar[0]), .ZN(ybar[112]);
  AND2_X1 U243 ( .A1(b[15]), .A2(a[6]), .ZN(y[111]) );
  OR2_X1 U243bar ( .A1(bbar[15]), .A2(abar[6]), .ZN(ybar[111]);
  AND2_X1 U244 ( .A1(b[14]), .A2(a[6]), .ZN(y[110]) );
  OR2_X1 U244bar ( .A1(bbar[14]), .A2(abar[6]), .ZN(ybar[110]);
  AND2_X1 U245 ( .A1(b[10]), .A2(a[0]), .ZN(y[10]) );
  OR2_X1 U245bar ( .A1(bbar[10]), .A2(abar[0]), .ZN(ybar[10]);
  AND2_X1 U246 ( .A1(b[13]), .A2(a[6]), .ZN(y[109]) );
  OR2_X1 U246bar ( .A1(bbar[13]), .A2(abar[6]), .ZN(ybar[109]);
  AND2_X1 U247 ( .A1(b[12]), .A2(a[6]), .ZN(y[108]) );
  OR2_X1 U247bar ( .A1(bbar[12]), .A2(abar[6]), .ZN(ybar[108]);
  AND2_X1 U248 ( .A1(b[11]), .A2(a[6]), .ZN(y[107]) );
  OR2_X1 U248bar ( .A1(bbar[11]), .A2(abar[6]), .ZN(ybar[107]);
  AND2_X1 U249 ( .A1(b[10]), .A2(a[6]), .ZN(y[106]) );
  OR2_X1 U249bar ( .A1(bbar[10]), .A2(abar[6]), .ZN(ybar[106]);
  AND2_X1 U250 ( .A1(a[6]), .A2(b[9]), .ZN(y[105]) );
  OR2_X1 U250bar ( .A1(abar[6]), .A2(bbar[9]), .ZN(ybar[105]);
  AND2_X1 U251 ( .A1(b[8]), .A2(a[6]), .ZN(y[104]) );
  OR2_X1 U251bar ( .A1(bbar[8]), .A2(abar[6]), .ZN(ybar[104]);
  AND2_X1 U252 ( .A1(b[7]), .A2(a[6]), .ZN(y[103]) );
  OR2_X1 U252bar ( .A1(bbar[7]), .A2(abar[6]), .ZN(ybar[103]);
  AND2_X1 U253 ( .A1(b[6]), .A2(a[6]), .ZN(y[102]) );
  OR2_X1 U253bar ( .A1(bbar[6]), .A2(abar[6]), .ZN(ybar[102]);
  AND2_X1 U254 ( .A1(b[5]), .A2(a[6]), .ZN(y[101]) );
  OR2_X1 U254bar ( .A1(bbar[5]), .A2(abar[6]), .ZN(ybar[101]);
  AND2_X1 U255 ( .A1(b[4]), .A2(a[6]), .ZN(y[100]) );
  OR2_X1 U255bar ( .A1(bbar[4]), .A2(abar[6]), .ZN(ybar[100]);
  AND2_X1 U256 ( .A1(b[0]), .A2(a[0]), .ZN(y[0]) );
  OR2_X1 U256bar ( .A1(bbar[0]), .A2(abar[0]), .ZN(ybar[0]);
endmodule




module decode_6 ( in, out );
  input [7:0] in;
  //input_done

  output [255:0] out;
  //output_done

  wire   [15:0] level1;
  wire   [31:0] level2;
  //wire_done

  CD2_24 cd_l1_1 ( .a(in[1]), .b(in[0]), .y(level1[3:0]) );
  CD2_23 cd_l1_2 ( .a(in[3]), .b(in[2]), .y(level1[7:4]) );
  CD2_22 cd_l1_3 ( .a(in[5]), .b(in[4]), .y(level1[11:8]) );
  CD2_21 cd_l1_4 ( .a(in[7]), .b(in[6]), .y(level1[15:12]) );
  CD4_12 cd_l2_1 ( .a(level1[7:4]), .b(level1[3:0]), .y(level2[15:0]) );
  CD4_11 cd_l2_2 ( .a(level1[15:12]), .b(level1[11:8]), .y(level2[31:16]) );
  CD16_6 cd_l3 ( .a(level2[31:16]), .b(level2[15:0]), .y(out) );
endmodule


module encode_6 ( in, out );
  input [255:0] in;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
  assign inbar[8] = ~in[8];
  assign inbar[9] = ~in[9];
  assign inbar[10] = ~in[10];
  assign inbar[11] = ~in[11];
  assign inbar[12] = ~in[12];
  assign inbar[13] = ~in[13];
  assign inbar[14] = ~in[14];
  assign inbar[15] = ~in[15];
  assign inbar[16] = ~in[16];
  assign inbar[17] = ~in[17];
  assign inbar[18] = ~in[18];
  assign inbar[19] = ~in[19];
  assign inbar[20] = ~in[20];
  assign inbar[21] = ~in[21];
  assign inbar[22] = ~in[22];
  assign inbar[23] = ~in[23];
  assign inbar[24] = ~in[24];
  assign inbar[25] = ~in[25];
  assign inbar[26] = ~in[26];
  assign inbar[27] = ~in[27];
  assign inbar[28] = ~in[28];
  assign inbar[29] = ~in[29];
  assign inbar[30] = ~in[30];
  assign inbar[31] = ~in[31];
  assign inbar[32] = ~in[32];
  assign inbar[33] = ~in[33];
  assign inbar[34] = ~in[34];
  assign inbar[35] = ~in[35];
  assign inbar[36] = ~in[36];
  assign inbar[37] = ~in[37];
  assign inbar[38] = ~in[38];
  assign inbar[39] = ~in[39];
  assign inbar[40] = ~in[40];
  assign inbar[41] = ~in[41];
  assign inbar[42] = ~in[42];
  assign inbar[43] = ~in[43];
  assign inbar[44] = ~in[44];
  assign inbar[45] = ~in[45];
  assign inbar[46] = ~in[46];
  assign inbar[47] = ~in[47];
  assign inbar[48] = ~in[48];
  assign inbar[49] = ~in[49];
  assign inbar[50] = ~in[50];
  assign inbar[51] = ~in[51];
  assign inbar[52] = ~in[52];
  assign inbar[53] = ~in[53];
  assign inbar[54] = ~in[54];
  assign inbar[55] = ~in[55];
  assign inbar[56] = ~in[56];
  assign inbar[57] = ~in[57];
  assign inbar[58] = ~in[58];
  assign inbar[59] = ~in[59];
  assign inbar[60] = ~in[60];
  assign inbar[61] = ~in[61];
  assign inbar[62] = ~in[62];
  assign inbar[63] = ~in[63];
  assign inbar[64] = ~in[64];
  assign inbar[65] = ~in[65];
  assign inbar[66] = ~in[66];
  assign inbar[67] = ~in[67];
  assign inbar[68] = ~in[68];
  assign inbar[69] = ~in[69];
  assign inbar[70] = ~in[70];
  assign inbar[71] = ~in[71];
  assign inbar[72] = ~in[72];
  assign inbar[73] = ~in[73];
  assign inbar[74] = ~in[74];
  assign inbar[75] = ~in[75];
  assign inbar[76] = ~in[76];
  assign inbar[77] = ~in[77];
  assign inbar[78] = ~in[78];
  assign inbar[79] = ~in[79];
  assign inbar[80] = ~in[80];
  assign inbar[81] = ~in[81];
  assign inbar[82] = ~in[82];
  assign inbar[83] = ~in[83];
  assign inbar[84] = ~in[84];
  assign inbar[85] = ~in[85];
  assign inbar[86] = ~in[86];
  assign inbar[87] = ~in[87];
  assign inbar[88] = ~in[88];
  assign inbar[89] = ~in[89];
  assign inbar[90] = ~in[90];
  assign inbar[91] = ~in[91];
  assign inbar[92] = ~in[92];
  assign inbar[93] = ~in[93];
  assign inbar[94] = ~in[94];
  assign inbar[95] = ~in[95];
  assign inbar[96] = ~in[96];
  assign inbar[97] = ~in[97];
  assign inbar[98] = ~in[98];
  assign inbar[99] = ~in[99];
  assign inbar[100] = ~in[100];
  assign inbar[101] = ~in[101];
  assign inbar[102] = ~in[102];
  assign inbar[103] = ~in[103];
  assign inbar[104] = ~in[104];
  assign inbar[105] = ~in[105];
  assign inbar[106] = ~in[106];
  assign inbar[107] = ~in[107];
  assign inbar[108] = ~in[108];
  assign inbar[109] = ~in[109];
  assign inbar[110] = ~in[110];
  assign inbar[111] = ~in[111];
  assign inbar[112] = ~in[112];
  assign inbar[113] = ~in[113];
  assign inbar[114] = ~in[114];
  assign inbar[115] = ~in[115];
  assign inbar[116] = ~in[116];
  assign inbar[117] = ~in[117];
  assign inbar[118] = ~in[118];
  assign inbar[119] = ~in[119];
  assign inbar[120] = ~in[120];
  assign inbar[121] = ~in[121];
  assign inbar[122] = ~in[122];
  assign inbar[123] = ~in[123];
  assign inbar[124] = ~in[124];
  assign inbar[125] = ~in[125];
  assign inbar[126] = ~in[126];
  assign inbar[127] = ~in[127];
  assign inbar[128] = ~in[128];
  assign inbar[129] = ~in[129];
  assign inbar[130] = ~in[130];
  assign inbar[131] = ~in[131];
  assign inbar[132] = ~in[132];
  assign inbar[133] = ~in[133];
  assign inbar[134] = ~in[134];
  assign inbar[135] = ~in[135];
  assign inbar[136] = ~in[136];
  assign inbar[137] = ~in[137];
  assign inbar[138] = ~in[138];
  assign inbar[139] = ~in[139];
  assign inbar[140] = ~in[140];
  assign inbar[141] = ~in[141];
  assign inbar[142] = ~in[142];
  assign inbar[143] = ~in[143];
  assign inbar[144] = ~in[144];
  assign inbar[145] = ~in[145];
  assign inbar[146] = ~in[146];
  assign inbar[147] = ~in[147];
  assign inbar[148] = ~in[148];
  assign inbar[149] = ~in[149];
  assign inbar[150] = ~in[150];
  assign inbar[151] = ~in[151];
  assign inbar[152] = ~in[152];
  assign inbar[153] = ~in[153];
  assign inbar[154] = ~in[154];
  assign inbar[155] = ~in[155];
  assign inbar[156] = ~in[156];
  assign inbar[157] = ~in[157];
  assign inbar[158] = ~in[158];
  assign inbar[159] = ~in[159];
  assign inbar[160] = ~in[160];
  assign inbar[161] = ~in[161];
  assign inbar[162] = ~in[162];
  assign inbar[163] = ~in[163];
  assign inbar[164] = ~in[164];
  assign inbar[165] = ~in[165];
  assign inbar[166] = ~in[166];
  assign inbar[167] = ~in[167];
  assign inbar[168] = ~in[168];
  assign inbar[169] = ~in[169];
  assign inbar[170] = ~in[170];
  assign inbar[171] = ~in[171];
  assign inbar[172] = ~in[172];
  assign inbar[173] = ~in[173];
  assign inbar[174] = ~in[174];
  assign inbar[175] = ~in[175];
  assign inbar[176] = ~in[176];
  assign inbar[177] = ~in[177];
  assign inbar[178] = ~in[178];
  assign inbar[179] = ~in[179];
  assign inbar[180] = ~in[180];
  assign inbar[181] = ~in[181];
  assign inbar[182] = ~in[182];
  assign inbar[183] = ~in[183];
  assign inbar[184] = ~in[184];
  assign inbar[185] = ~in[185];
  assign inbar[186] = ~in[186];
  assign inbar[187] = ~in[187];
  assign inbar[188] = ~in[188];
  assign inbar[189] = ~in[189];
  assign inbar[190] = ~in[190];
  assign inbar[191] = ~in[191];
  assign inbar[192] = ~in[192];
  assign inbar[193] = ~in[193];
  assign inbar[194] = ~in[194];
  assign inbar[195] = ~in[195];
  assign inbar[196] = ~in[196];
  assign inbar[197] = ~in[197];
  assign inbar[198] = ~in[198];
  assign inbar[199] = ~in[199];
  assign inbar[200] = ~in[200];
  assign inbar[201] = ~in[201];
  assign inbar[202] = ~in[202];
  assign inbar[203] = ~in[203];
  assign inbar[204] = ~in[204];
  assign inbar[205] = ~in[205];
  assign inbar[206] = ~in[206];
  assign inbar[207] = ~in[207];
  assign inbar[208] = ~in[208];
  assign inbar[209] = ~in[209];
  assign inbar[210] = ~in[210];
  assign inbar[211] = ~in[211];
  assign inbar[212] = ~in[212];
  assign inbar[213] = ~in[213];
  assign inbar[214] = ~in[214];
  assign inbar[215] = ~in[215];
  assign inbar[216] = ~in[216];
  assign inbar[217] = ~in[217];
  assign inbar[218] = ~in[218];
  assign inbar[219] = ~in[219];
  assign inbar[220] = ~in[220];
  assign inbar[221] = ~in[221];
  assign inbar[222] = ~in[222];
  assign inbar[223] = ~in[223];
  assign inbar[224] = ~in[224];
  assign inbar[225] = ~in[225];
  assign inbar[226] = ~in[226];
  assign inbar[227] = ~in[227];
  assign inbar[228] = ~in[228];
  assign inbar[229] = ~in[229];
  assign inbar[230] = ~in[230];
  assign inbar[231] = ~in[231];
  assign inbar[232] = ~in[232];
  assign inbar[233] = ~in[233];
  assign inbar[234] = ~in[234];
  assign inbar[235] = ~in[235];
  assign inbar[236] = ~in[236];
  assign inbar[237] = ~in[237];
  assign inbar[238] = ~in[238];
  assign inbar[239] = ~in[239];
  assign inbar[240] = ~in[240];
  assign inbar[241] = ~in[241];
  assign inbar[242] = ~in[242];
  assign inbar[243] = ~in[243];
  assign inbar[244] = ~in[244];
  assign inbar[245] = ~in[245];
  assign inbar[246] = ~in[246];
  assign inbar[247] = ~in[247];
  assign inbar[248] = ~in[248];
  assign inbar[249] = ~in[249];
  assign inbar[250] = ~in[250];
  assign inbar[251] = ~in[251];
  assign inbar[252] = ~in[252];
  assign inbar[253] = ~in[253];
  assign inbar[254] = ~in[254];
  assign inbar[255] = ~in[255];
  //input_done

  output [7:0] out;
  reg [7:0] outbar;
  //output_done

  wire   in_81, in_80, in_79, in_78, in_77, in_76, in_75, in_74, in_73, in_72,
         in_71, in_70, in_69, in_68, in_67, in_66, in_65, in_64, in_63, in_62,
         in_61, in_60, in_59, in_58, in_57, in_56, in_55, in_54, in_53, in_52,
         in_51, in_50, in_49, in_48, in_47, in_46, in_45, in_44, in_43, in_42,
         in_41, in_40, in_39, in_38, in_37, in_36, in_35, in_34, in_33, in_32,
         in_31, in_30, in_29, in_28, in_27, in_26, in_25, in_24, in_23, in_22,
         in_21, in_20, in_19, in_18, in_17, in_16, in_15, in_14, in_13, in_12,
         in_11, in_10, in_9, in_8, in_7, in_6, in_5, in_4, in_3, in_2, in_1,
         in_0, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972;
  wire in_81bar, in_80bar, in_79bar, in_78bar, in_77bar, in_76bar, in_75bar, in_74bar, in_73bar, in_72bar, in_71bar, in_70bar, in_69bar, in_68bar, in_67bar, in_66bar, in_65bar, in_64bar, in_63bar, in_62bar, in_61bar, in_60bar, in_59bar, in_58bar, in_57bar, in_56bar, in_55bar, in_54bar, in_53bar, in_52bar, in_51bar, in_50bar, in_49bar, in_48bar, in_47bar, in_46bar, in_45bar, in_44bar, in_43bar, in_42bar, in_41bar, in_40bar, in_39bar, in_38bar, in_37bar, in_36bar, in_35bar, in_34bar, in_33bar, in_32bar, in_31bar, in_30bar, in_29bar, in_28bar, in_27bar, in_26bar, in_25bar, in_24bar, in_23bar, in_22bar, in_21bar, in_20bar, in_19bar, in_18bar, in_17bar, in_16bar, in_15bar, in_14bar, in_13bar, in_12bar, in_11bar, in_10bar, in_9bar, in_8bar, in_7bar, in_6bar, in_5bar, in_4bar, in_3bar, in_2bar, in_1bar, in_0bar, n487bar, n488bar, n489bar, n490bar, n491bar, n492bar, n493bar, n494bar, n495bar, n496bar, n497bar, n498bar, n499bar, n500bar, n501bar, n502bar, n503bar, n504bar, n505bar, n506bar, n507bar, n508bar, n509bar, n510bar, n511bar, n512bar, n513bar, n514bar, n515bar, n516bar, n517bar, n518bar, n519bar, n520bar, n521bar, n522bar, n523bar, n524bar, n525bar, n526bar, n527bar, n528bar, n529bar, n530bar, n531bar, n532bar, n533bar, n534bar, n535bar, n536bar, n537bar, n538bar, n539bar, n540bar, n541bar, n542bar, n543bar, n544bar, n545bar, n546bar, n547bar, n548bar, n549bar, n550bar, n551bar, n552bar, n553bar, n554bar, n555bar, n556bar, n557bar, n558bar, n559bar, n560bar, n561bar, n562bar, n563bar, n564bar, n565bar, n566bar, n567bar, n568bar, n569bar, n570bar, n571bar, n572bar, n573bar, n574bar, n575bar, n576bar, n577bar, n578bar, n579bar, n580bar, n581bar, n582bar, n583bar, n584bar, n585bar, n586bar, n587bar, n588bar, n589bar, n590bar, n591bar, n592bar, n593bar, n594bar, n595bar, n596bar, n597bar, n598bar, n599bar, n600bar, n601bar, n602bar, n603bar, n604bar, n605bar, n606bar, n607bar, n608bar, n609bar, n610bar, n611bar, n612bar, n613bar, n614bar, n615bar, n616bar, n617bar, n618bar, n619bar, n620bar, n621bar, n622bar, n623bar, n624bar, n625bar, n626bar, n627bar, n628bar, n629bar, n630bar, n631bar, n632bar, n633bar, n634bar, n635bar, n636bar, n637bar, n638bar, n639bar, n640bar, n641bar, n642bar, n643bar, n644bar, n645bar, n646bar, n647bar, n648bar, n649bar, n650bar, n651bar, n652bar, n653bar, n654bar, n655bar, n656bar, n657bar, n658bar, n659bar, n660bar, n661bar, n662bar, n663bar, n664bar, n665bar, n666bar, n667bar, n668bar, n669bar, n670bar, n671bar, n672bar, n673bar, n674bar, n675bar, n676bar, n677bar, n678bar, n679bar, n680bar, n681bar, n682bar, n683bar, n684bar, n685bar, n686bar, n687bar, n688bar, n689bar, n690bar, n691bar, n692bar, n693bar, n694bar, n695bar, n696bar, n697bar, n698bar, n699bar, n700bar, n701bar, n702bar, n703bar, n704bar, n705bar, n706bar, n707bar, n708bar, n709bar, n710bar, n711bar, n712bar, n713bar, n714bar, n715bar, n716bar, n717bar, n718bar, n719bar, n720bar, n721bar, n722bar, n723bar, n724bar, n725bar, n726bar, n727bar, n728bar, n729bar, n730bar, n731bar, n732bar, n733bar, n734bar, n735bar, n736bar, n737bar, n738bar, n739bar, n740bar, n741bar, n742bar, n743bar, n744bar, n745bar, n746bar, n747bar, n748bar, n749bar, n750bar, n751bar, n752bar, n753bar, n754bar, n755bar, n756bar, n757bar, n758bar, n759bar, n760bar, n761bar, n762bar, n763bar, n764bar, n765bar, n766bar, n767bar, n768bar, n769bar, n770bar, n771bar, n772bar, n773bar, n774bar, n775bar, n776bar, n777bar, n778bar, n779bar, n780bar, n781bar, n782bar, n783bar, n784bar, n785bar, n786bar, n787bar, n788bar, n789bar, n790bar, n791bar, n792bar, n793bar, n794bar, n795bar, n796bar, n797bar, n798bar, n799bar, n800bar, n801bar, n802bar, n803bar, n804bar, n805bar, n806bar, n807bar, n808bar, n809bar, n810bar, n811bar, n812bar, n813bar, n814bar, n815bar, n816bar, n817bar, n818bar, n819bar, n820bar, n821bar, n822bar, n823bar, n824bar, n825bar, n826bar, n827bar, n828bar, n829bar, n830bar, n831bar, n832bar, n833bar, n834bar, n835bar, n836bar, n837bar, n838bar, n839bar, n840bar, n841bar, n842bar, n843bar, n844bar, n845bar, n846bar, n847bar, n848bar, n849bar, n850bar, n851bar, n852bar, n853bar, n854bar, n855bar, n856bar, n857bar, n858bar, n859bar, n860bar, n861bar, n862bar, n863bar, n864bar, n865bar, n866bar, n867bar, n868bar, n869bar, n870bar, n871bar, n872bar, n873bar, n874bar, n875bar, n876bar, n877bar, n878bar, n879bar, n880bar, n881bar, n882bar, n883bar, n884bar, n885bar, n886bar, n887bar, n888bar, n889bar, n890bar, n891bar, n892bar, n893bar, n894bar, n895bar, n896bar, n897bar, n898bar, n899bar, n900bar, n901bar, n902bar, n903bar, n904bar, n905bar, n906bar, n907bar, n908bar, n909bar, n910bar, n911bar, n912bar, n913bar, n914bar, n915bar, n916bar, n917bar, n918bar, n919bar, n920bar, n921bar, n922bar, n923bar, n924bar, n925bar, n926bar, n927bar, n928bar, n929bar, n930bar, n931bar, n932bar, n933bar, n934bar, n935bar, n936bar, n937bar, n938bar, n939bar, n940bar, n941bar, n942bar, n943bar, n944bar, n945bar, n946bar, n947bar, n948bar, n949bar, n950bar, n951bar, n952bar, n953bar, n954bar, n955bar, n956bar, n957bar, n958bar, n959bar, n960bar, n961bar, n962bar, n963bar, n964bar, n965bar, n966bar, n967bar, n968bar, n969bar, n970bar, n971bar, n972bar;
  //wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];

  OR2_X1 U1 ( .A1(n972), .A2(n971), .ZN(out[7]) );
  AND2_X1 U1bar ( .A1(n972bar), .A2(n971bar), .ZN(outbar[7]);
  OR2_X1 U2 ( .A1(n970), .A2(n969), .ZN(n971) );
  AND2_X1 U2bar ( .A1(n970bar), .A2(n969bar), .ZN(n971bar);
  OR2_X1 U3 ( .A1(n968), .A2(n967), .ZN(n969) );
  AND2_X1 U3bar ( .A1(n968bar), .A2(n967bar), .ZN(n969bar);
  OR2_X1 U4 ( .A1(n966), .A2(n965), .ZN(n967) );
  AND2_X1 U4bar ( .A1(n966bar), .A2(n965bar), .ZN(n967bar);
  OR2_X1 U5 ( .A1(n964), .A2(n963), .ZN(n968) );
  AND2_X1 U5bar ( .A1(n964bar), .A2(n963bar), .ZN(n968bar);
  OR2_X1 U6 ( .A1(in[116]), .A2(n962), .ZN(n963) );
  AND2_X1 U6bar ( .A1(inbar[116]), .A2(n962bar), .ZN(n963bar);
  OR2_X1 U7 ( .A1(n961), .A2(n960), .ZN(n970) );
  AND2_X1 U7bar ( .A1(n961bar), .A2(n960bar), .ZN(n970bar);
  OR2_X1 U8 ( .A1(in[150]), .A2(in[127]), .ZN(n960) );
  AND2_X1 U8bar ( .A1(inbar[150]), .A2(inbar[127]), .ZN(n960bar);
  OR2_X1 U9 ( .A1(in[160]), .A2(n959), .ZN(n961) );
  AND2_X1 U9bar ( .A1(inbar[160]), .A2(n959bar), .ZN(n961bar);
  OR2_X1 U10 ( .A1(in[252]), .A2(in[168]), .ZN(n959) );
  AND2_X1 U10bar ( .A1(inbar[252]), .A2(inbar[168]), .ZN(n959bar);
  OR2_X1 U11 ( .A1(n958), .A2(n957), .ZN(n972) );
  AND2_X1 U11bar ( .A1(n958bar), .A2(n957bar), .ZN(n972bar);
  OR2_X1 U12 ( .A1(n956), .A2(n955), .ZN(n957) );
  AND2_X1 U12bar ( .A1(n956bar), .A2(n955bar), .ZN(n957bar);
  OR2_X1 U13 ( .A1(in_17), .A2(in[96]), .ZN(n955) );
  AND2_X1 U13bar ( .A1(in_17bar), .A2(inbar[96]), .ZN(n955bar);
  OR2_X1 U14 ( .A1(in_23), .A2(n954), .ZN(n956) );
  AND2_X1 U14bar ( .A1(in_23bar), .A2(n954bar), .ZN(n956bar);
  OR2_X1 U15 ( .A1(in_31), .A2(in_26), .ZN(n954) );
  AND2_X1 U15bar ( .A1(in_31bar), .A2(in_26bar), .ZN(n954bar);
  OR2_X1 U16 ( .A1(n953), .A2(n952), .ZN(n958) );
  AND2_X1 U16bar ( .A1(n953bar), .A2(n952bar), .ZN(n958bar);
  OR2_X1 U17 ( .A1(in_58), .A2(in_4), .ZN(n952) );
  AND2_X1 U17bar ( .A1(in_58bar), .A2(in_4bar), .ZN(n952bar);
  OR2_X1 U18 ( .A1(in_59), .A2(n951), .ZN(n953) );
  AND2_X1 U18bar ( .A1(in_59bar), .A2(n951bar), .ZN(n953bar);
  OR2_X1 U19 ( .A1(in_71), .A2(in_62), .ZN(n951) );
  AND2_X1 U19bar ( .A1(in_71bar), .A2(in_62bar), .ZN(n951bar);
  OR2_X1 U20 ( .A1(n950), .A2(n949), .ZN(out[6]) );
  AND2_X1 U20bar ( .A1(n950bar), .A2(n949bar), .ZN(outbar[6]);
  OR2_X1 U21 ( .A1(n948), .A2(n947), .ZN(n949) );
  AND2_X1 U21bar ( .A1(n948bar), .A2(n947bar), .ZN(n949bar);
  OR2_X1 U22 ( .A1(n946), .A2(n945), .ZN(n947) );
  AND2_X1 U22bar ( .A1(n946bar), .A2(n945bar), .ZN(n947bar);
  OR2_X1 U23 ( .A1(n944), .A2(n943), .ZN(n945) );
  AND2_X1 U23bar ( .A1(n944bar), .A2(n943bar), .ZN(n945bar);
  OR2_X1 U24 ( .A1(n942), .A2(n941), .ZN(n946) );
  AND2_X1 U24bar ( .A1(n942bar), .A2(n941bar), .ZN(n946bar);
  OR2_X1 U25 ( .A1(in[101]), .A2(n940), .ZN(n941) );
  AND2_X1 U25bar ( .A1(inbar[101]), .A2(n940bar), .ZN(n941bar);
  OR2_X1 U26 ( .A1(n939), .A2(n938), .ZN(n948) );
  AND2_X1 U26bar ( .A1(n939bar), .A2(n938bar), .ZN(n948bar);
  OR2_X1 U27 ( .A1(in[114]), .A2(in[104]), .ZN(n938) );
  AND2_X1 U27bar ( .A1(inbar[114]), .A2(inbar[104]), .ZN(n938bar);
  OR2_X1 U28 ( .A1(in[128]), .A2(n937), .ZN(n939) );
  AND2_X1 U28bar ( .A1(inbar[128]), .A2(n937bar), .ZN(n939bar);
  OR2_X1 U29 ( .A1(in[136]), .A2(in[134]), .ZN(n937) );
  AND2_X1 U29bar ( .A1(inbar[136]), .A2(inbar[134]), .ZN(n937bar);
  OR2_X1 U30 ( .A1(n936), .A2(n935), .ZN(n950) );
  AND2_X1 U30bar ( .A1(n936bar), .A2(n935bar), .ZN(n950bar);
  OR2_X1 U31 ( .A1(n934), .A2(n933), .ZN(n935) );
  AND2_X1 U31bar ( .A1(n934bar), .A2(n933bar), .ZN(n935bar);
  OR2_X1 U32 ( .A1(in[177]), .A2(in[164]), .ZN(n933) );
  AND2_X1 U32bar ( .A1(inbar[177]), .A2(inbar[164]), .ZN(n933bar);
  OR2_X1 U33 ( .A1(in[212]), .A2(n932), .ZN(n934) );
  AND2_X1 U33bar ( .A1(inbar[212]), .A2(n932bar), .ZN(n934bar);
  OR2_X1 U34 ( .A1(in[248]), .A2(in[221]), .ZN(n932) );
  AND2_X1 U34bar ( .A1(inbar[248]), .A2(inbar[221]), .ZN(n932bar);
  OR2_X1 U35 ( .A1(n931), .A2(n930), .ZN(n936) );
  AND2_X1 U35bar ( .A1(n931bar), .A2(n930bar), .ZN(n936bar);
  OR2_X1 U36 ( .A1(in_18), .A2(in[93]), .ZN(n930) );
  AND2_X1 U36bar ( .A1(in_18bar), .A2(inbar[93]), .ZN(n930bar);
  OR2_X1 U37 ( .A1(in_31), .A2(n929), .ZN(n931) );
  AND2_X1 U37bar ( .A1(in_31bar), .A2(n929bar), .ZN(n931bar);
  OR2_X1 U38 ( .A1(in_7), .A2(in_39), .ZN(n929) );
  AND2_X1 U38bar ( .A1(in_7bar), .A2(in_39bar), .ZN(n929bar);
  OR2_X1 U39 ( .A1(n928), .A2(n927), .ZN(out[5]) );
  AND2_X1 U39bar ( .A1(n928bar), .A2(n927bar), .ZN(outbar[5]);
  OR2_X1 U40 ( .A1(n926), .A2(n925), .ZN(n927) );
  AND2_X1 U40bar ( .A1(n926bar), .A2(n925bar), .ZN(n927bar);
  OR2_X1 U41 ( .A1(n924), .A2(n923), .ZN(n925) );
  AND2_X1 U41bar ( .A1(n924bar), .A2(n923bar), .ZN(n925bar);
  OR2_X1 U42 ( .A1(n922), .A2(n921), .ZN(n923) );
  AND2_X1 U42bar ( .A1(n922bar), .A2(n921bar), .ZN(n923bar);
  OR2_X1 U43 ( .A1(n940), .A2(n920), .ZN(n924) );
  AND2_X1 U43bar ( .A1(n940bar), .A2(n920bar), .ZN(n924bar);
  OR2_X1 U44 ( .A1(in[111]), .A2(n919), .ZN(n920) );
  AND2_X1 U44bar ( .A1(inbar[111]), .A2(n919bar), .ZN(n920bar);
  OR2_X1 U45 ( .A1(n918), .A2(n917), .ZN(n940) );
  AND2_X1 U45bar ( .A1(n918bar), .A2(n917bar), .ZN(n940bar);
  OR2_X1 U46 ( .A1(n916), .A2(n915), .ZN(n917) );
  AND2_X1 U46bar ( .A1(n916bar), .A2(n915bar), .ZN(n917bar);
  OR2_X1 U47 ( .A1(n914), .A2(n913), .ZN(n915) );
  AND2_X1 U47bar ( .A1(n914bar), .A2(n913bar), .ZN(n915bar);
  OR2_X1 U48 ( .A1(in[140]), .A2(in[131]), .ZN(n913) );
  AND2_X1 U48bar ( .A1(inbar[140]), .A2(inbar[131]), .ZN(n913bar);
  OR2_X1 U49 ( .A1(in[160]), .A2(in[144]), .ZN(n914) );
  AND2_X1 U49bar ( .A1(inbar[160]), .A2(inbar[144]), .ZN(n914bar);
  OR2_X1 U50 ( .A1(n912), .A2(n911), .ZN(n916) );
  AND2_X1 U50bar ( .A1(n912bar), .A2(n911bar), .ZN(n916bar);
  OR2_X1 U51 ( .A1(in[179]), .A2(in[174]), .ZN(n911) );
  AND2_X1 U51bar ( .A1(inbar[179]), .A2(inbar[174]), .ZN(n911bar);
  OR2_X1 U52 ( .A1(in[188]), .A2(in[184]), .ZN(n912) );
  AND2_X1 U52bar ( .A1(inbar[188]), .A2(inbar[184]), .ZN(n912bar);
  OR2_X1 U53 ( .A1(n910), .A2(n909), .ZN(n918) );
  AND2_X1 U53bar ( .A1(n910bar), .A2(n909bar), .ZN(n918bar);
  OR2_X1 U54 ( .A1(n908), .A2(n907), .ZN(n909) );
  AND2_X1 U54bar ( .A1(n908bar), .A2(n907bar), .ZN(n909bar);
  OR2_X1 U55 ( .A1(in[216]), .A2(in[200]), .ZN(n907) );
  AND2_X1 U55bar ( .A1(inbar[216]), .A2(inbar[200]), .ZN(n907bar);
  OR2_X1 U56 ( .A1(in[228]), .A2(in[224]), .ZN(n908) );
  AND2_X1 U56bar ( .A1(inbar[228]), .A2(inbar[224]), .ZN(n908bar);
  OR2_X1 U57 ( .A1(n906), .A2(n905), .ZN(n910) );
  AND2_X1 U57bar ( .A1(n906bar), .A2(n905bar), .ZN(n910bar);
  OR2_X1 U58 ( .A1(in[247]), .A2(in[235]), .ZN(n905) );
  AND2_X1 U58bar ( .A1(inbar[247]), .A2(inbar[235]), .ZN(n905bar);
  OR2_X1 U59 ( .A1(in_42), .A2(in[83]), .ZN(n906) );
  AND2_X1 U59bar ( .A1(in_42bar), .A2(inbar[83]), .ZN(n906bar);
  OR2_X1 U60 ( .A1(n904), .A2(n903), .ZN(n926) );
  AND2_X1 U60bar ( .A1(n904bar), .A2(n903bar), .ZN(n926bar);
  OR2_X1 U61 ( .A1(in[166]), .A2(in[123]), .ZN(n903) );
  AND2_X1 U61bar ( .A1(inbar[166]), .A2(inbar[123]), .ZN(n903bar);
  OR2_X1 U62 ( .A1(in[170]), .A2(n902), .ZN(n904) );
  AND2_X1 U62bar ( .A1(inbar[170]), .A2(n902bar), .ZN(n904bar);
  OR2_X1 U63 ( .A1(in[194]), .A2(in[183]), .ZN(n902) );
  AND2_X1 U63bar ( .A1(inbar[194]), .A2(inbar[183]), .ZN(n902bar);
  OR2_X1 U64 ( .A1(n901), .A2(n900), .ZN(n928) );
  AND2_X1 U64bar ( .A1(n901bar), .A2(n900bar), .ZN(n928bar);
  OR2_X1 U65 ( .A1(n899), .A2(n898), .ZN(n900) );
  AND2_X1 U65bar ( .A1(n899bar), .A2(n898bar), .ZN(n900bar);
  OR2_X1 U66 ( .A1(in[241]), .A2(in[238]), .ZN(n898) );
  AND2_X1 U66bar ( .A1(inbar[241]), .A2(inbar[238]), .ZN(n898bar);
  OR2_X1 U67 ( .A1(in[250]), .A2(n897), .ZN(n899) );
  AND2_X1 U67bar ( .A1(inbar[250]), .A2(n897bar), .ZN(n899bar);
  OR2_X1 U68 ( .A1(in_24), .A2(in[84]), .ZN(n897) );
  AND2_X1 U68bar ( .A1(in_24bar), .A2(inbar[84]), .ZN(n897bar);
  OR2_X1 U69 ( .A1(n896), .A2(n895), .ZN(n901) );
  AND2_X1 U69bar ( .A1(n896bar), .A2(n895bar), .ZN(n901bar);
  OR2_X1 U70 ( .A1(in_41), .A2(in_29), .ZN(n895) );
  AND2_X1 U70bar ( .A1(in_41bar), .A2(in_29bar), .ZN(n895bar);
  OR2_X1 U71 ( .A1(in_66), .A2(n894), .ZN(n896) );
  AND2_X1 U71bar ( .A1(in_66bar), .A2(n894bar), .ZN(n896bar);
  OR2_X1 U72 ( .A1(in_76), .A2(in_71), .ZN(n894) );
  AND2_X1 U72bar ( .A1(in_76bar), .A2(in_71bar), .ZN(n894bar);
  OR2_X1 U73 ( .A1(n893), .A2(n892), .ZN(out[4]) );
  AND2_X1 U73bar ( .A1(n893bar), .A2(n892bar), .ZN(outbar[4]);
  OR2_X1 U74 ( .A1(n891), .A2(n890), .ZN(n892) );
  AND2_X1 U74bar ( .A1(n891bar), .A2(n890bar), .ZN(n892bar);
  OR2_X1 U75 ( .A1(n889), .A2(n888), .ZN(n890) );
  AND2_X1 U75bar ( .A1(n889bar), .A2(n888bar), .ZN(n890bar);
  OR2_X1 U76 ( .A1(n922), .A2(n887), .ZN(n888) );
  AND2_X1 U76bar ( .A1(n922bar), .A2(n887bar), .ZN(n888bar);
  OR2_X1 U77 ( .A1(n886), .A2(n885), .ZN(n922) );
  AND2_X1 U77bar ( .A1(n886bar), .A2(n885bar), .ZN(n922bar);
  OR2_X1 U78 ( .A1(n884), .A2(n883), .ZN(n885) );
  AND2_X1 U78bar ( .A1(n884bar), .A2(n883bar), .ZN(n885bar);
  OR2_X1 U79 ( .A1(n882), .A2(n881), .ZN(n883) );
  AND2_X1 U79bar ( .A1(n882bar), .A2(n881bar), .ZN(n883bar);
  OR2_X1 U80 ( .A1(in[118]), .A2(in[109]), .ZN(n881) );
  AND2_X1 U80bar ( .A1(inbar[118]), .A2(inbar[109]), .ZN(n881bar);
  OR2_X1 U81 ( .A1(in[139]), .A2(in[120]), .ZN(n882) );
  AND2_X1 U81bar ( .A1(inbar[139]), .A2(inbar[120]), .ZN(n882bar);
  OR2_X1 U82 ( .A1(n880), .A2(n879), .ZN(n884) );
  AND2_X1 U82bar ( .A1(n880bar), .A2(n879bar), .ZN(n884bar);
  OR2_X1 U83 ( .A1(in[198]), .A2(in[154]), .ZN(n879) );
  AND2_X1 U83bar ( .A1(inbar[198]), .A2(inbar[154]), .ZN(n879bar);
  OR2_X1 U84 ( .A1(in[210]), .A2(in[205]), .ZN(n880) );
  AND2_X1 U84bar ( .A1(inbar[210]), .A2(inbar[205]), .ZN(n880bar);
  OR2_X1 U85 ( .A1(n878), .A2(n877), .ZN(n886) );
  AND2_X1 U85bar ( .A1(n878bar), .A2(n877bar), .ZN(n886bar);
  OR2_X1 U86 ( .A1(n876), .A2(n875), .ZN(n877) );
  AND2_X1 U86bar ( .A1(n876bar), .A2(n875bar), .ZN(n877bar);
  OR2_X1 U87 ( .A1(in[219]), .A2(in[217]), .ZN(n875) );
  AND2_X1 U87bar ( .A1(inbar[219]), .A2(inbar[217]), .ZN(n875bar);
  OR2_X1 U88 ( .A1(in[86]), .A2(in[252]), .ZN(n876) );
  AND2_X1 U88bar ( .A1(inbar[86]), .A2(inbar[252]), .ZN(n876bar);
  OR2_X1 U89 ( .A1(n874), .A2(n873), .ZN(n878) );
  AND2_X1 U89bar ( .A1(n874bar), .A2(n873bar), .ZN(n878bar);
  OR2_X1 U90 ( .A1(in_40), .A2(in[91]), .ZN(n873) );
  AND2_X1 U90bar ( .A1(in_40bar), .A2(inbar[91]), .ZN(n873bar);
  OR2_X1 U91 ( .A1(in_8), .A2(in_46), .ZN(n874) );
  AND2_X1 U91bar ( .A1(in_8bar), .A2(in_46bar), .ZN(n874bar);
  OR2_X1 U92 ( .A1(n872), .A2(n871), .ZN(n889) );
  AND2_X1 U92bar ( .A1(n872bar), .A2(n871bar), .ZN(n889bar);
  OR2_X1 U93 ( .A1(in[117]), .A2(n943), .ZN(n871) );
  AND2_X1 U93bar ( .A1(inbar[117]), .A2(n943bar), .ZN(n871bar);
  OR2_X1 U94 ( .A1(n870), .A2(n869), .ZN(n943) );
  AND2_X1 U94bar ( .A1(n870bar), .A2(n869bar), .ZN(n943bar);
  OR2_X1 U95 ( .A1(n868), .A2(n867), .ZN(n869) );
  AND2_X1 U95bar ( .A1(n868bar), .A2(n867bar), .ZN(n869bar);
  OR2_X1 U96 ( .A1(n866), .A2(n865), .ZN(n867) );
  AND2_X1 U96bar ( .A1(n866bar), .A2(n865bar), .ZN(n867bar);
  OR2_X1 U97 ( .A1(n864), .A2(n863), .ZN(n865) );
  AND2_X1 U97bar ( .A1(n864bar), .A2(n863bar), .ZN(n865bar);
  OR2_X1 U98 ( .A1(in[108]), .A2(n919), .ZN(n866) );
  AND2_X1 U98bar ( .A1(inbar[108]), .A2(n919bar), .ZN(n866bar);
  OR2_X1 U99 ( .A1(n862), .A2(n861), .ZN(n919) );
  AND2_X1 U99bar ( .A1(n862bar), .A2(n861bar), .ZN(n919bar);
  OR2_X1 U100 ( .A1(n860), .A2(n859), .ZN(n861) );
  AND2_X1 U100bar ( .A1(n860bar), .A2(n859bar), .ZN(n861bar);
  OR2_X1 U101 ( .A1(n858), .A2(n857), .ZN(n859) );
  AND2_X1 U101bar ( .A1(n858bar), .A2(n857bar), .ZN(n859bar);
  OR2_X1 U102 ( .A1(in[119]), .A2(in[105]), .ZN(n857) );
  AND2_X1 U102bar ( .A1(inbar[119]), .A2(inbar[105]), .ZN(n857bar);
  OR2_X1 U103 ( .A1(in[186]), .A2(in[175]), .ZN(n858) );
  AND2_X1 U103bar ( .A1(inbar[186]), .A2(inbar[175]), .ZN(n858bar);
  OR2_X1 U104 ( .A1(n856), .A2(n855), .ZN(n860) );
  AND2_X1 U104bar ( .A1(n856bar), .A2(n855bar), .ZN(n860bar);
  OR2_X1 U105 ( .A1(in[202]), .A2(in[193]), .ZN(n855) );
  AND2_X1 U105bar ( .A1(inbar[202]), .A2(inbar[193]), .ZN(n855bar);
  OR2_X1 U106 ( .A1(in[225]), .A2(in[208]), .ZN(n856) );
  AND2_X1 U106bar ( .A1(inbar[225]), .A2(inbar[208]), .ZN(n856bar);
  OR2_X1 U107 ( .A1(n854), .A2(n853), .ZN(n862) );
  AND2_X1 U107bar ( .A1(n854bar), .A2(n853bar), .ZN(n862bar);
  OR2_X1 U108 ( .A1(n852), .A2(n851), .ZN(n853) );
  AND2_X1 U108bar ( .A1(n852bar), .A2(n851bar), .ZN(n853bar);
  OR2_X1 U109 ( .A1(in_1), .A2(in[85]), .ZN(n851) );
  AND2_X1 U109bar ( .A1(in_1bar), .A2(inbar[85]), .ZN(n851bar);
  OR2_X1 U110 ( .A1(in_23), .A2(in_19), .ZN(n852) );
  AND2_X1 U110bar ( .A1(in_23bar), .A2(in_19bar), .ZN(n852bar);
  OR2_X1 U111 ( .A1(n850), .A2(n849), .ZN(n854) );
  AND2_X1 U111bar ( .A1(n850bar), .A2(n849bar), .ZN(n854bar);
  OR2_X1 U112 ( .A1(in_43), .A2(in_33), .ZN(n849) );
  AND2_X1 U112bar ( .A1(in_43bar), .A2(in_33bar), .ZN(n849bar);
  OR2_X1 U113 ( .A1(in_63), .A2(in_44), .ZN(n850) );
  AND2_X1 U113bar ( .A1(in_63bar), .A2(in_44bar), .ZN(n850bar);
  OR2_X1 U114 ( .A1(n848), .A2(n847), .ZN(n868) );
  AND2_X1 U114bar ( .A1(n848bar), .A2(n847bar), .ZN(n868bar);
  OR2_X1 U115 ( .A1(in[141]), .A2(in[112]), .ZN(n847) );
  AND2_X1 U115bar ( .A1(inbar[141]), .A2(inbar[112]), .ZN(n847bar);
  OR2_X1 U116 ( .A1(in[147]), .A2(n846), .ZN(n848) );
  AND2_X1 U116bar ( .A1(inbar[147]), .A2(n846bar), .ZN(n848bar);
  OR2_X1 U117 ( .A1(in[181]), .A2(in[167]), .ZN(n846) );
  AND2_X1 U117bar ( .A1(inbar[181]), .A2(inbar[167]), .ZN(n846bar);
  OR2_X1 U118 ( .A1(n845), .A2(n844), .ZN(n870) );
  AND2_X1 U118bar ( .A1(n845bar), .A2(n844bar), .ZN(n870bar);
  OR2_X1 U119 ( .A1(n843), .A2(n842), .ZN(n844) );
  AND2_X1 U119bar ( .A1(n843bar), .A2(n842bar), .ZN(n844bar);
  OR2_X1 U120 ( .A1(in[229]), .A2(in[201]), .ZN(n842) );
  AND2_X1 U120bar ( .A1(inbar[229]), .A2(inbar[201]), .ZN(n842bar);
  OR2_X1 U121 ( .A1(in[237]), .A2(n841), .ZN(n843) );
  AND2_X1 U121bar ( .A1(inbar[237]), .A2(n841bar), .ZN(n843bar);
  OR2_X1 U122 ( .A1(in[94]), .A2(in[253]), .ZN(n841) );
  AND2_X1 U122bar ( .A1(inbar[94]), .A2(inbar[253]), .ZN(n841bar);
  OR2_X1 U123 ( .A1(n840), .A2(n839), .ZN(n845) );
  AND2_X1 U123bar ( .A1(n840bar), .A2(n839bar), .ZN(n845bar);
  OR2_X1 U124 ( .A1(in_21), .A2(in[96]), .ZN(n839) );
  AND2_X1 U124bar ( .A1(in_21bar), .A2(inbar[96]), .ZN(n839bar);
  OR2_X1 U125 ( .A1(in_25), .A2(n838), .ZN(n840) );
  AND2_X1 U125bar ( .A1(in_25bar), .A2(n838bar), .ZN(n840bar);
  OR2_X1 U126 ( .A1(in_81), .A2(in_45), .ZN(n838) );
  AND2_X1 U126bar ( .A1(in_81bar), .A2(in_45bar), .ZN(n838bar);
  OR2_X1 U127 ( .A1(n837), .A2(n836), .ZN(n891) );
  AND2_X1 U127bar ( .A1(n837bar), .A2(n836bar), .ZN(n891bar);
  OR2_X1 U128 ( .A1(in[142]), .A2(in[124]), .ZN(n836) );
  AND2_X1 U128bar ( .A1(inbar[142]), .A2(inbar[124]), .ZN(n836bar);
  OR2_X1 U129 ( .A1(in[150]), .A2(n835), .ZN(n837) );
  AND2_X1 U129bar ( .A1(inbar[150]), .A2(n835bar), .ZN(n837bar);
  OR2_X1 U130 ( .A1(in[172]), .A2(in[155]), .ZN(n835) );
  AND2_X1 U130bar ( .A1(inbar[172]), .A2(inbar[155]), .ZN(n835bar);
  OR2_X1 U131 ( .A1(n834), .A2(n833), .ZN(n893) );
  AND2_X1 U131bar ( .A1(n834bar), .A2(n833bar), .ZN(n893bar);
  OR2_X1 U132 ( .A1(n832), .A2(n831), .ZN(n833) );
  AND2_X1 U132bar ( .A1(n832bar), .A2(n831bar), .ZN(n833bar);
  OR2_X1 U133 ( .A1(in[196]), .A2(in[173]), .ZN(n831) );
  AND2_X1 U133bar ( .A1(inbar[196]), .A2(inbar[173]), .ZN(n831bar);
  OR2_X1 U134 ( .A1(in[222]), .A2(n830), .ZN(n832) );
  AND2_X1 U134bar ( .A1(inbar[222]), .A2(n830bar), .ZN(n832bar);
  OR2_X1 U135 ( .A1(in[227]), .A2(in[226]), .ZN(n830) );
  AND2_X1 U135bar ( .A1(inbar[227]), .A2(inbar[226]), .ZN(n830bar);
  OR2_X1 U136 ( .A1(n829), .A2(n828), .ZN(n834) );
  AND2_X1 U136bar ( .A1(n829bar), .A2(n828bar), .ZN(n834bar);
  OR2_X1 U137 ( .A1(in[249]), .A2(in[231]), .ZN(n828) );
  AND2_X1 U137bar ( .A1(inbar[249]), .A2(inbar[231]), .ZN(n828bar);
  OR2_X1 U138 ( .A1(in_28), .A2(n827), .ZN(n829) );
  AND2_X1 U138bar ( .A1(in_28bar), .A2(n827bar), .ZN(n829bar);
  OR2_X1 U139 ( .A1(in_52), .A2(in_47), .ZN(n827) );
  AND2_X1 U139bar ( .A1(in_52bar), .A2(in_47bar), .ZN(n827bar);
  OR2_X1 U140 ( .A1(n826), .A2(n825), .ZN(out[3]) );
  AND2_X1 U140bar ( .A1(n826bar), .A2(n825bar), .ZN(outbar[3]);
  OR2_X1 U141 ( .A1(n824), .A2(n823), .ZN(n825) );
  AND2_X1 U141bar ( .A1(n824bar), .A2(n823bar), .ZN(n825bar);
  OR2_X1 U142 ( .A1(n822), .A2(n821), .ZN(n823) );
  AND2_X1 U142bar ( .A1(n822bar), .A2(n821bar), .ZN(n823bar);
  OR2_X1 U143 ( .A1(n820), .A2(n819), .ZN(n821) );
  AND2_X1 U143bar ( .A1(n820bar), .A2(n819bar), .ZN(n821bar);
  OR2_X1 U144 ( .A1(n964), .A2(n818), .ZN(n822) );
  AND2_X1 U144bar ( .A1(n964bar), .A2(n818bar), .ZN(n822bar);
  OR2_X1 U145 ( .A1(in[118]), .A2(n817), .ZN(n818) );
  AND2_X1 U145bar ( .A1(inbar[118]), .A2(n817bar), .ZN(n818bar);
  OR2_X1 U146 ( .A1(n816), .A2(n815), .ZN(n964) );
  AND2_X1 U146bar ( .A1(n816bar), .A2(n815bar), .ZN(n964bar);
  OR2_X1 U147 ( .A1(n814), .A2(n813), .ZN(n815) );
  AND2_X1 U147bar ( .A1(n814bar), .A2(n813bar), .ZN(n815bar);
  OR2_X1 U148 ( .A1(n812), .A2(n811), .ZN(n813) );
  AND2_X1 U148bar ( .A1(n812bar), .A2(n811bar), .ZN(n813bar);
  OR2_X1 U149 ( .A1(in[122]), .A2(in[111]), .ZN(n811) );
  AND2_X1 U149bar ( .A1(inbar[122]), .A2(inbar[111]), .ZN(n811bar);
  OR2_X1 U150 ( .A1(in[154]), .A2(in[151]), .ZN(n812) );
  AND2_X1 U150bar ( .A1(inbar[154]), .A2(inbar[151]), .ZN(n812bar);
  OR2_X1 U151 ( .A1(n810), .A2(n809), .ZN(n814) );
  AND2_X1 U151bar ( .A1(n810bar), .A2(n809bar), .ZN(n814bar);
  OR2_X1 U152 ( .A1(in[187]), .A2(in[177]), .ZN(n809) );
  AND2_X1 U152bar ( .A1(inbar[187]), .A2(inbar[177]), .ZN(n809bar);
  OR2_X1 U153 ( .A1(in[200]), .A2(in[192]), .ZN(n810) );
  AND2_X1 U153bar ( .A1(inbar[200]), .A2(inbar[192]), .ZN(n810bar);
  OR2_X1 U154 ( .A1(n808), .A2(n807), .ZN(n816) );
  AND2_X1 U154bar ( .A1(n808bar), .A2(n807bar), .ZN(n816bar);
  OR2_X1 U155 ( .A1(n806), .A2(n805), .ZN(n807) );
  AND2_X1 U155bar ( .A1(n806bar), .A2(n805bar), .ZN(n807bar);
  OR2_X1 U156 ( .A1(in[225]), .A2(in[207]), .ZN(n805) );
  AND2_X1 U156bar ( .A1(inbar[225]), .A2(inbar[207]), .ZN(n805bar);
  OR2_X1 U157 ( .A1(in[98]), .A2(in[226]), .ZN(n806) );
  AND2_X1 U157bar ( .A1(inbar[98]), .A2(inbar[226]), .ZN(n806bar);
  OR2_X1 U158 ( .A1(n804), .A2(n803), .ZN(n808) );
  AND2_X1 U158bar ( .A1(n804bar), .A2(n803bar), .ZN(n808bar);
  OR2_X1 U159 ( .A1(in_20), .A2(in_16), .ZN(n803) );
  AND2_X1 U159bar ( .A1(in_20bar), .A2(in_16bar), .ZN(n803bar);
  OR2_X1 U160 ( .A1(in_55), .A2(in_45), .ZN(n804) );
  AND2_X1 U160bar ( .A1(in_55bar), .A2(in_45bar), .ZN(n804bar);
  OR2_X1 U161 ( .A1(n802), .A2(n801), .ZN(n824) );
  AND2_X1 U161bar ( .A1(n802bar), .A2(n801bar), .ZN(n824bar);
  OR2_X1 U162 ( .A1(in[162]), .A2(in[149]), .ZN(n801) );
  AND2_X1 U162bar ( .A1(inbar[162]), .A2(inbar[149]), .ZN(n801bar);
  OR2_X1 U163 ( .A1(in[163]), .A2(n800), .ZN(n802) );
  AND2_X1 U163bar ( .A1(inbar[163]), .A2(n800bar), .ZN(n802bar);
  OR2_X1 U164 ( .A1(in[191]), .A2(in[189]), .ZN(n800) );
  AND2_X1 U164bar ( .A1(inbar[191]), .A2(inbar[189]), .ZN(n800bar);
  OR2_X1 U165 ( .A1(n799), .A2(n798), .ZN(n826) );
  AND2_X1 U165bar ( .A1(n799bar), .A2(n798bar), .ZN(n826bar);
  OR2_X1 U166 ( .A1(n797), .A2(n796), .ZN(n798) );
  AND2_X1 U166bar ( .A1(n797bar), .A2(n796bar), .ZN(n798bar);
  OR2_X1 U167 ( .A1(in[212]), .A2(in[193]), .ZN(n796) );
  AND2_X1 U167bar ( .A1(inbar[212]), .A2(inbar[193]), .ZN(n796bar);
  OR2_X1 U168 ( .A1(in[238]), .A2(n795), .ZN(n797) );
  AND2_X1 U168bar ( .A1(inbar[238]), .A2(n795bar), .ZN(n797bar);
  OR2_X1 U169 ( .A1(in[88]), .A2(in[247]), .ZN(n795) );
  AND2_X1 U169bar ( .A1(inbar[88]), .A2(inbar[247]), .ZN(n795bar);
  OR2_X1 U170 ( .A1(n794), .A2(n793), .ZN(n799) );
  AND2_X1 U170bar ( .A1(n794bar), .A2(n793bar), .ZN(n799bar);
  OR2_X1 U171 ( .A1(in[94]), .A2(in[92]), .ZN(n793) );
  AND2_X1 U171bar ( .A1(inbar[94]), .A2(inbar[92]), .ZN(n793bar);
  OR2_X1 U172 ( .A1(in_52), .A2(n792), .ZN(n794) );
  AND2_X1 U172bar ( .A1(in_52bar), .A2(n792bar), .ZN(n794bar);
  OR2_X1 U173 ( .A1(in_70), .A2(in_67), .ZN(n792) );
  AND2_X1 U173bar ( .A1(in_70bar), .A2(in_67bar), .ZN(n792bar);
  OR2_X1 U174 ( .A1(n791), .A2(n790), .ZN(out[2]) );
  AND2_X1 U174bar ( .A1(n791bar), .A2(n790bar), .ZN(outbar[2]);
  OR2_X1 U175 ( .A1(n789), .A2(n788), .ZN(n790) );
  AND2_X1 U175bar ( .A1(n789bar), .A2(n788bar), .ZN(n790bar);
  OR2_X1 U176 ( .A1(n787), .A2(n786), .ZN(n788) );
  AND2_X1 U176bar ( .A1(n787bar), .A2(n786bar), .ZN(n788bar);
  OR2_X1 U177 ( .A1(n819), .A2(n785), .ZN(n786) );
  AND2_X1 U177bar ( .A1(n819bar), .A2(n785bar), .ZN(n786bar);
  OR2_X1 U178 ( .A1(n784), .A2(n783), .ZN(n819) );
  AND2_X1 U178bar ( .A1(n784bar), .A2(n783bar), .ZN(n819bar);
  OR2_X1 U179 ( .A1(n782), .A2(n781), .ZN(n783) );
  AND2_X1 U179bar ( .A1(n782bar), .A2(n781bar), .ZN(n783bar);
  OR2_X1 U180 ( .A1(n780), .A2(n779), .ZN(n781) );
  AND2_X1 U180bar ( .A1(n780bar), .A2(n779bar), .ZN(n781bar);
  OR2_X1 U181 ( .A1(n962), .A2(n778), .ZN(n779) );
  AND2_X1 U181bar ( .A1(n962bar), .A2(n778bar), .ZN(n779bar);
  OR2_X1 U182 ( .A1(n777), .A2(n776), .ZN(n962) );
  AND2_X1 U182bar ( .A1(n777bar), .A2(n776bar), .ZN(n962bar);
  OR2_X1 U183 ( .A1(n775), .A2(n774), .ZN(n776) );
  AND2_X1 U183bar ( .A1(n775bar), .A2(n774bar), .ZN(n776bar);
  OR2_X1 U184 ( .A1(n773), .A2(n772), .ZN(n774) );
  AND2_X1 U184bar ( .A1(n773bar), .A2(n772bar), .ZN(n774bar);
  OR2_X1 U185 ( .A1(in[131]), .A2(in[120]), .ZN(n772) );
  AND2_X1 U185bar ( .A1(inbar[131]), .A2(inbar[120]), .ZN(n772bar);
  OR2_X1 U186 ( .A1(in[153]), .A2(in[147]), .ZN(n773) );
  AND2_X1 U186bar ( .A1(inbar[153]), .A2(inbar[147]), .ZN(n773bar);
  OR2_X1 U187 ( .A1(n771), .A2(n770), .ZN(n775) );
  AND2_X1 U187bar ( .A1(n771bar), .A2(n770bar), .ZN(n775bar);
  OR2_X1 U188 ( .A1(in[170]), .A2(in[156]), .ZN(n770) );
  AND2_X1 U188bar ( .A1(inbar[170]), .A2(inbar[156]), .ZN(n770bar);
  OR2_X1 U189 ( .A1(in[223]), .A2(in[190]), .ZN(n771) );
  AND2_X1 U189bar ( .A1(inbar[223]), .A2(inbar[190]), .ZN(n771bar);
  OR2_X1 U190 ( .A1(n769), .A2(n768), .ZN(n777) );
  AND2_X1 U190bar ( .A1(n769bar), .A2(n768bar), .ZN(n777bar);
  OR2_X1 U191 ( .A1(n767), .A2(n766), .ZN(n768) );
  AND2_X1 U191bar ( .A1(n767bar), .A2(n766bar), .ZN(n768bar);
  OR2_X1 U192 ( .A1(in[236]), .A2(in[230]), .ZN(n766) );
  AND2_X1 U192bar ( .A1(inbar[236]), .A2(inbar[230]), .ZN(n766bar);
  OR2_X1 U193 ( .A1(in[85]), .A2(in[240]), .ZN(n767) );
  AND2_X1 U193bar ( .A1(inbar[85]), .A2(inbar[240]), .ZN(n767bar);
  OR2_X1 U194 ( .A1(n765), .A2(n764), .ZN(n769) );
  AND2_X1 U194bar ( .A1(n765bar), .A2(n764bar), .ZN(n769bar);
  OR2_X1 U195 ( .A1(in_12), .A2(in[90]), .ZN(n764) );
  AND2_X1 U195bar ( .A1(in_12bar), .A2(inbar[90]), .ZN(n764bar);
  OR2_X1 U196 ( .A1(in_39), .A2(in_28), .ZN(n765) );
  AND2_X1 U196bar ( .A1(in_39bar), .A2(in_28bar), .ZN(n765bar);
  OR2_X1 U197 ( .A1(in[109]), .A2(n763), .ZN(n780) );
  AND2_X1 U197bar ( .A1(inbar[109]), .A2(n763bar), .ZN(n780bar);
  OR2_X1 U198 ( .A1(n762), .A2(n761), .ZN(n782) );
  AND2_X1 U198bar ( .A1(n762bar), .A2(n761bar), .ZN(n782bar);
  OR2_X1 U199 ( .A1(in[138]), .A2(in[129]), .ZN(n761) );
  AND2_X1 U199bar ( .A1(inbar[138]), .A2(inbar[129]), .ZN(n761bar);
  OR2_X1 U200 ( .A1(in[157]), .A2(n760), .ZN(n762) );
  AND2_X1 U200bar ( .A1(inbar[157]), .A2(n760bar), .ZN(n762bar);
  OR2_X1 U201 ( .A1(in[182]), .A2(in[167]), .ZN(n760) );
  AND2_X1 U201bar ( .A1(inbar[182]), .A2(inbar[167]), .ZN(n760bar);
  OR2_X1 U202 ( .A1(n759), .A2(n758), .ZN(n784) );
  AND2_X1 U202bar ( .A1(n759bar), .A2(n758bar), .ZN(n784bar);
  OR2_X1 U203 ( .A1(n757), .A2(n756), .ZN(n758) );
  AND2_X1 U203bar ( .A1(n757bar), .A2(n756bar), .ZN(n758bar);
  OR2_X1 U204 ( .A1(in[195]), .A2(in[184]), .ZN(n756) );
  AND2_X1 U204bar ( .A1(inbar[195]), .A2(inbar[184]), .ZN(n756bar);
  OR2_X1 U205 ( .A1(in[196]), .A2(n755), .ZN(n757) );
  AND2_X1 U205bar ( .A1(inbar[196]), .A2(n755bar), .ZN(n757bar);
  OR2_X1 U206 ( .A1(in[215]), .A2(in[209]), .ZN(n755) );
  AND2_X1 U206bar ( .A1(inbar[215]), .A2(inbar[209]), .ZN(n755bar);
  OR2_X1 U207 ( .A1(n754), .A2(n753), .ZN(n759) );
  AND2_X1 U207bar ( .A1(n754bar), .A2(n753bar), .ZN(n759bar);
  OR2_X1 U208 ( .A1(in[93]), .A2(in[233]), .ZN(n753) );
  AND2_X1 U208bar ( .A1(inbar[93]), .A2(inbar[233]), .ZN(n753bar);
  OR2_X1 U209 ( .A1(in_1), .A2(n752), .ZN(n754) );
  AND2_X1 U209bar ( .A1(in_1bar), .A2(n752bar), .ZN(n754bar);
  OR2_X1 U210 ( .A1(in_69), .A2(in_66), .ZN(n752) );
  AND2_X1 U210bar ( .A1(in_69bar), .A2(in_66bar), .ZN(n752bar);
  OR2_X1 U211 ( .A1(n966), .A2(n751), .ZN(n787) );
  AND2_X1 U211bar ( .A1(n966bar), .A2(n751bar), .ZN(n787bar);
  OR2_X1 U212 ( .A1(in[134]), .A2(n750), .ZN(n751) );
  AND2_X1 U212bar ( .A1(inbar[134]), .A2(n750bar), .ZN(n751bar);
  OR2_X1 U213 ( .A1(n749), .A2(n748), .ZN(n966) );
  AND2_X1 U213bar ( .A1(n749bar), .A2(n748bar), .ZN(n966bar);
  OR2_X1 U214 ( .A1(n747), .A2(n746), .ZN(n748) );
  AND2_X1 U214bar ( .A1(n747bar), .A2(n746bar), .ZN(n748bar);
  OR2_X1 U215 ( .A1(n745), .A2(n744), .ZN(n746) );
  AND2_X1 U215bar ( .A1(n745bar), .A2(n744bar), .ZN(n746bar);
  OR2_X1 U216 ( .A1(in[136]), .A2(in[121]), .ZN(n744) );
  AND2_X1 U216bar ( .A1(inbar[136]), .A2(inbar[121]), .ZN(n744bar);
  OR2_X1 U217 ( .A1(in[186]), .A2(in[174]), .ZN(n745) );
  AND2_X1 U217bar ( .A1(inbar[186]), .A2(inbar[174]), .ZN(n745bar);
  OR2_X1 U218 ( .A1(n743), .A2(n742), .ZN(n747) );
  AND2_X1 U218bar ( .A1(n743bar), .A2(n742bar), .ZN(n747bar);
  OR2_X1 U219 ( .A1(in[198]), .A2(in[197]), .ZN(n742) );
  AND2_X1 U219bar ( .A1(inbar[198]), .A2(inbar[197]), .ZN(n742bar);
  OR2_X1 U220 ( .A1(in[214]), .A2(in[199]), .ZN(n743) );
  AND2_X1 U220bar ( .A1(inbar[214]), .A2(inbar[199]), .ZN(n743bar);
  OR2_X1 U221 ( .A1(n741), .A2(n740), .ZN(n749) );
  AND2_X1 U221bar ( .A1(n741bar), .A2(n740bar), .ZN(n749bar);
  OR2_X1 U222 ( .A1(n739), .A2(n738), .ZN(n740) );
  AND2_X1 U222bar ( .A1(n739bar), .A2(n738bar), .ZN(n740bar);
  OR2_X1 U223 ( .A1(in[231]), .A2(in[220]), .ZN(n738) );
  AND2_X1 U223bar ( .A1(inbar[231]), .A2(inbar[220]), .ZN(n738bar);
  OR2_X1 U224 ( .A1(in_25), .A2(in[245]), .ZN(n739) );
  AND2_X1 U224bar ( .A1(in_25bar), .A2(inbar[245]), .ZN(n739bar);
  OR2_X1 U225 ( .A1(n737), .A2(n736), .ZN(n741) );
  AND2_X1 U225bar ( .A1(n737bar), .A2(n736bar), .ZN(n741bar);
  OR2_X1 U226 ( .A1(in_53), .A2(in_29), .ZN(n736) );
  AND2_X1 U226bar ( .A1(in_53bar), .A2(in_29bar), .ZN(n736bar);
  OR2_X1 U227 ( .A1(in_79), .A2(in_74), .ZN(n737) );
  AND2_X1 U227bar ( .A1(in_79bar), .A2(in_74bar), .ZN(n737bar);
  OR2_X1 U228 ( .A1(n735), .A2(n734), .ZN(n789) );
  AND2_X1 U228bar ( .A1(n735bar), .A2(n734bar), .ZN(n789bar);
  OR2_X1 U229 ( .A1(in[152]), .A2(in[140]), .ZN(n734) );
  AND2_X1 U229bar ( .A1(inbar[152]), .A2(inbar[140]), .ZN(n734bar);
  OR2_X1 U230 ( .A1(in[155]), .A2(n733), .ZN(n735) );
  AND2_X1 U230bar ( .A1(inbar[155]), .A2(n733bar), .ZN(n735bar);
  OR2_X1 U231 ( .A1(in[166]), .A2(in[165]), .ZN(n733) );
  AND2_X1 U231bar ( .A1(inbar[166]), .A2(inbar[165]), .ZN(n733bar);
  OR2_X1 U232 ( .A1(n732), .A2(n731), .ZN(n791) );
  AND2_X1 U232bar ( .A1(n732bar), .A2(n731bar), .ZN(n791bar);
  OR2_X1 U233 ( .A1(n730), .A2(n729), .ZN(n731) );
  AND2_X1 U233bar ( .A1(n730bar), .A2(n729bar), .ZN(n731bar);
  OR2_X1 U234 ( .A1(in[202]), .A2(in[185]), .ZN(n729) );
  AND2_X1 U234bar ( .A1(inbar[202]), .A2(inbar[185]), .ZN(n729bar);
  OR2_X1 U235 ( .A1(in[211]), .A2(n728), .ZN(n730) );
  AND2_X1 U235bar ( .A1(inbar[211]), .A2(n728bar), .ZN(n730bar);
  OR2_X1 U236 ( .A1(in[255]), .A2(in[253]), .ZN(n728) );
  AND2_X1 U236bar ( .A1(inbar[255]), .A2(inbar[253]), .ZN(n728bar);
  OR2_X1 U237 ( .A1(n727), .A2(n726), .ZN(n732) );
  AND2_X1 U237bar ( .A1(n727bar), .A2(n726bar), .ZN(n732bar);
  OR2_X1 U238 ( .A1(in_35), .A2(in_15), .ZN(n726) );
  AND2_X1 U238bar ( .A1(in_35bar), .A2(in_15bar), .ZN(n726bar);
  OR2_X1 U239 ( .A1(in_36), .A2(n725), .ZN(n727) );
  AND2_X1 U239bar ( .A1(in_36bar), .A2(n725bar), .ZN(n727bar);
  OR2_X1 U240 ( .A1(in_48), .A2(in_40), .ZN(n725) );
  AND2_X1 U240bar ( .A1(in_48bar), .A2(in_40bar), .ZN(n725bar);
  OR2_X1 U241 ( .A1(n724), .A2(n723), .ZN(out[1]) );
  AND2_X1 U241bar ( .A1(n724bar), .A2(n723bar), .ZN(outbar[1]);
  OR2_X1 U242 ( .A1(n722), .A2(n721), .ZN(n723) );
  AND2_X1 U242bar ( .A1(n722bar), .A2(n721bar), .ZN(n723bar);
  OR2_X1 U243 ( .A1(n720), .A2(n719), .ZN(n721) );
  AND2_X1 U243bar ( .A1(n720bar), .A2(n719bar), .ZN(n721bar);
  OR2_X1 U244 ( .A1(n921), .A2(n887), .ZN(n719) );
  AND2_X1 U244bar ( .A1(n921bar), .A2(n887bar), .ZN(n719bar);
  OR2_X1 U245 ( .A1(n718), .A2(n717), .ZN(n887) );
  AND2_X1 U245bar ( .A1(n718bar), .A2(n717bar), .ZN(n887bar);
  OR2_X1 U246 ( .A1(n716), .A2(n715), .ZN(n717) );
  AND2_X1 U246bar ( .A1(n716bar), .A2(n715bar), .ZN(n717bar);
  OR2_X1 U247 ( .A1(n714), .A2(n713), .ZN(n715) );
  AND2_X1 U247bar ( .A1(n714bar), .A2(n713bar), .ZN(n715bar);
  OR2_X1 U248 ( .A1(in[116]), .A2(in[110]), .ZN(n713) );
  AND2_X1 U248bar ( .A1(inbar[116]), .A2(inbar[110]), .ZN(n713bar);
  OR2_X1 U249 ( .A1(in[133]), .A2(in[130]), .ZN(n714) );
  AND2_X1 U249bar ( .A1(inbar[133]), .A2(inbar[130]), .ZN(n714bar);
  OR2_X1 U250 ( .A1(n712), .A2(n711), .ZN(n716) );
  AND2_X1 U250bar ( .A1(n712bar), .A2(n711bar), .ZN(n716bar);
  OR2_X1 U251 ( .A1(in[203]), .A2(in[135]), .ZN(n711) );
  AND2_X1 U251bar ( .A1(inbar[203]), .A2(inbar[135]), .ZN(n711bar);
  OR2_X1 U252 ( .A1(in[232]), .A2(in[223]), .ZN(n712) );
  AND2_X1 U252bar ( .A1(inbar[232]), .A2(inbar[223]), .ZN(n712bar);
  OR2_X1 U253 ( .A1(n710), .A2(n709), .ZN(n718) );
  AND2_X1 U253bar ( .A1(n710bar), .A2(n709bar), .ZN(n718bar);
  OR2_X1 U254 ( .A1(n708), .A2(n707), .ZN(n709) );
  AND2_X1 U254bar ( .A1(n708bar), .A2(n707bar), .ZN(n709bar);
  OR2_X1 U255 ( .A1(in[255]), .A2(in[233]), .ZN(n707) );
  AND2_X1 U255bar ( .A1(inbar[255]), .A2(inbar[233]), .ZN(n707bar);
  OR2_X1 U256 ( .A1(in_53), .A2(in_34), .ZN(n708) );
  AND2_X1 U256bar ( .A1(in_53bar), .A2(in_34bar), .ZN(n708bar);
  OR2_X1 U257 ( .A1(n706), .A2(n705), .ZN(n710) );
  AND2_X1 U257bar ( .A1(n706bar), .A2(n705bar), .ZN(n710bar);
  OR2_X1 U258 ( .A1(in_57), .A2(in_55), .ZN(n705) );
  AND2_X1 U258bar ( .A1(in_57bar), .A2(in_55bar), .ZN(n705bar);
  OR2_X1 U259 ( .A1(in_68), .A2(in_67), .ZN(n706) );
  AND2_X1 U259bar ( .A1(in_68bar), .A2(in_67bar), .ZN(n706bar);
  OR2_X1 U260 ( .A1(n704), .A2(n703), .ZN(n921) );
  AND2_X1 U260bar ( .A1(n704bar), .A2(n703bar), .ZN(n921bar);
  OR2_X1 U261 ( .A1(n702), .A2(n701), .ZN(n703) );
  AND2_X1 U261bar ( .A1(n702bar), .A2(n701bar), .ZN(n703bar);
  OR2_X1 U262 ( .A1(n700), .A2(n699), .ZN(n701) );
  AND2_X1 U262bar ( .A1(n700bar), .A2(n699bar), .ZN(n701bar);
  OR2_X1 U263 ( .A1(n944), .A2(n872), .ZN(n699) );
  AND2_X1 U263bar ( .A1(n944bar), .A2(n872bar), .ZN(n699bar);
  OR2_X1 U264 ( .A1(n698), .A2(n697), .ZN(n872) );
  AND2_X1 U264bar ( .A1(n698bar), .A2(n697bar), .ZN(n872bar);
  OR2_X1 U265 ( .A1(n696), .A2(n695), .ZN(n697) );
  AND2_X1 U265bar ( .A1(n696bar), .A2(n695bar), .ZN(n697bar);
  OR2_X1 U266 ( .A1(n694), .A2(n693), .ZN(n695) );
  AND2_X1 U266bar ( .A1(n694bar), .A2(n693bar), .ZN(n695bar);
  OR2_X1 U267 ( .A1(in[121]), .A2(in[102]), .ZN(n693) );
  AND2_X1 U267bar ( .A1(inbar[121]), .A2(inbar[102]), .ZN(n693bar);
  OR2_X1 U268 ( .A1(in[162]), .A2(in[161]), .ZN(n694) );
  AND2_X1 U268bar ( .A1(inbar[162]), .A2(inbar[161]), .ZN(n694bar);
  OR2_X1 U269 ( .A1(n692), .A2(n691), .ZN(n696) );
  AND2_X1 U269bar ( .A1(n692bar), .A2(n691bar), .ZN(n696bar);
  OR2_X1 U270 ( .A1(in[192]), .A2(in[178]), .ZN(n691) );
  AND2_X1 U270bar ( .A1(inbar[192]), .A2(inbar[178]), .ZN(n691bar);
  OR2_X1 U271 ( .A1(in[244]), .A2(in[209]), .ZN(n692) );
  AND2_X1 U271bar ( .A1(inbar[244]), .A2(inbar[209]), .ZN(n692bar);
  OR2_X1 U272 ( .A1(n690), .A2(n689), .ZN(n698) );
  AND2_X1 U272bar ( .A1(n690bar), .A2(n689bar), .ZN(n698bar);
  OR2_X1 U273 ( .A1(n688), .A2(n687), .ZN(n689) );
  AND2_X1 U273bar ( .A1(n688bar), .A2(n687bar), .ZN(n689bar);
  OR2_X1 U274 ( .A1(in[90]), .A2(in[254]), .ZN(n687) );
  AND2_X1 U274bar ( .A1(inbar[90]), .A2(inbar[254]), .ZN(n687bar);
  OR2_X1 U275 ( .A1(in_36), .A2(in_32), .ZN(n688) );
  AND2_X1 U275bar ( .A1(in_36bar), .A2(in_32bar), .ZN(n688bar);
  OR2_X1 U276 ( .A1(n686), .A2(n685), .ZN(n690) );
  AND2_X1 U276bar ( .A1(n686bar), .A2(n685bar), .ZN(n690bar);
  OR2_X1 U277 ( .A1(in_62), .A2(in_37), .ZN(n685) );
  AND2_X1 U277bar ( .A1(in_62bar), .A2(in_37bar), .ZN(n685bar);
  OR2_X1 U278 ( .A1(in_75), .A2(in_73), .ZN(n686) );
  AND2_X1 U278bar ( .A1(in_75bar), .A2(in_73bar), .ZN(n686bar);
  OR2_X1 U279 ( .A1(n684), .A2(n683), .ZN(n944) );
  AND2_X1 U279bar ( .A1(n684bar), .A2(n683bar), .ZN(n944bar);
  OR2_X1 U280 ( .A1(n682), .A2(n681), .ZN(n683) );
  AND2_X1 U280bar ( .A1(n682bar), .A2(n681bar), .ZN(n683bar);
  OR2_X1 U281 ( .A1(n680), .A2(n679), .ZN(n681) );
  AND2_X1 U281bar ( .A1(n680bar), .A2(n679bar), .ZN(n681bar);
  OR2_X1 U282 ( .A1(in[171]), .A2(in[153]), .ZN(n679) );
  AND2_X1 U282bar ( .A1(inbar[171]), .A2(inbar[153]), .ZN(n679bar);
  OR2_X1 U283 ( .A1(in[187]), .A2(in[176]), .ZN(n680) );
  AND2_X1 U283bar ( .A1(inbar[187]), .A2(inbar[176]), .ZN(n680bar);
  OR2_X1 U284 ( .A1(n678), .A2(n677), .ZN(n682) );
  AND2_X1 U284bar ( .A1(n678bar), .A2(n677bar), .ZN(n682bar);
  OR2_X1 U285 ( .A1(in[245]), .A2(in[211]), .ZN(n677) );
  AND2_X1 U285bar ( .A1(inbar[245]), .A2(inbar[211]), .ZN(n677bar);
  OR2_X1 U286 ( .A1(in[97]), .A2(in[88]), .ZN(n678) );
  AND2_X1 U286bar ( .A1(inbar[97]), .A2(inbar[88]), .ZN(n678bar);
  OR2_X1 U287 ( .A1(n676), .A2(n675), .ZN(n684) );
  AND2_X1 U287bar ( .A1(n676bar), .A2(n675bar), .ZN(n684bar);
  OR2_X1 U288 ( .A1(n674), .A2(n673), .ZN(n675) );
  AND2_X1 U288bar ( .A1(n674bar), .A2(n673bar), .ZN(n675bar);
  OR2_X1 U289 ( .A1(in_10), .A2(in_0), .ZN(n673) );
  AND2_X1 U289bar ( .A1(in_10bar), .A2(in_0bar), .ZN(n673bar);
  OR2_X1 U290 ( .A1(in_59), .A2(in_5), .ZN(n674) );
  AND2_X1 U290bar ( .A1(in_59bar), .A2(in_5bar), .ZN(n674bar);
  OR2_X1 U291 ( .A1(n672), .A2(n671), .ZN(n676) );
  AND2_X1 U291bar ( .A1(n672bar), .A2(n671bar), .ZN(n676bar);
  OR2_X1 U292 ( .A1(in_60), .A2(in_6), .ZN(n671) );
  AND2_X1 U292bar ( .A1(in_60bar), .A2(in_6bar), .ZN(n671bar);
  OR2_X1 U293 ( .A1(in_77), .A2(in_69), .ZN(n672) );
  AND2_X1 U293bar ( .A1(in_77bar), .A2(in_69bar), .ZN(n672bar);
  OR2_X1 U294 ( .A1(in[113]), .A2(n864), .ZN(n700) );
  AND2_X1 U294bar ( .A1(inbar[113]), .A2(n864bar), .ZN(n700bar);
  OR2_X1 U295 ( .A1(n670), .A2(n669), .ZN(n864) );
  AND2_X1 U295bar ( .A1(n670bar), .A2(n669bar), .ZN(n864bar);
  OR2_X1 U296 ( .A1(n668), .A2(n667), .ZN(n669) );
  AND2_X1 U296bar ( .A1(n668bar), .A2(n667bar), .ZN(n669bar);
  OR2_X1 U297 ( .A1(n666), .A2(n665), .ZN(n667) );
  AND2_X1 U297bar ( .A1(n666bar), .A2(n665bar), .ZN(n667bar);
  OR2_X1 U298 ( .A1(in[125]), .A2(in[107]), .ZN(n665) );
  AND2_X1 U298bar ( .A1(inbar[125]), .A2(inbar[107]), .ZN(n665bar);
  OR2_X1 U299 ( .A1(in[138]), .A2(in[126]), .ZN(n666) );
  AND2_X1 U299bar ( .A1(inbar[138]), .A2(inbar[126]), .ZN(n666bar);
  OR2_X1 U300 ( .A1(n664), .A2(n663), .ZN(n668) );
  AND2_X1 U300bar ( .A1(n664bar), .A2(n663bar), .ZN(n668bar);
  OR2_X1 U301 ( .A1(in[189]), .A2(in[143]), .ZN(n663) );
  AND2_X1 U301bar ( .A1(inbar[189]), .A2(inbar[143]), .ZN(n663bar);
  OR2_X1 U302 ( .A1(in[99]), .A2(in[214]), .ZN(n664) );
  AND2_X1 U302bar ( .A1(inbar[99]), .A2(inbar[214]), .ZN(n664bar);
  OR2_X1 U303 ( .A1(n662), .A2(n661), .ZN(n670) );
  AND2_X1 U303bar ( .A1(n662bar), .A2(n661bar), .ZN(n670bar);
  OR2_X1 U304 ( .A1(n660), .A2(n659), .ZN(n661) );
  AND2_X1 U304bar ( .A1(n660bar), .A2(n659bar), .ZN(n661bar);
  OR2_X1 U305 ( .A1(in_15), .A2(in_12), .ZN(n659) );
  AND2_X1 U305bar ( .A1(in_15bar), .A2(in_12bar), .ZN(n659bar);
  OR2_X1 U306 ( .A1(in_20), .A2(in_2), .ZN(n660) );
  AND2_X1 U306bar ( .A1(in_20bar), .A2(in_2bar), .ZN(n660bar);
  OR2_X1 U307 ( .A1(n658), .A2(n657), .ZN(n662) );
  AND2_X1 U307bar ( .A1(n658bar), .A2(n657bar), .ZN(n662bar);
  OR2_X1 U308 ( .A1(in_30), .A2(in_3), .ZN(n657) );
  AND2_X1 U308bar ( .A1(in_30bar), .A2(in_3bar), .ZN(n657bar);
  OR2_X1 U309 ( .A1(in_4), .A2(in_38), .ZN(n658) );
  AND2_X1 U309bar ( .A1(in_4bar), .A2(in_38bar), .ZN(n658bar);
  OR2_X1 U310 ( .A1(n656), .A2(n655), .ZN(n702) );
  AND2_X1 U310bar ( .A1(n656bar), .A2(n655bar), .ZN(n702bar);
  OR2_X1 U311 ( .A1(in[148]), .A2(in[137]), .ZN(n655) );
  AND2_X1 U311bar ( .A1(inbar[148]), .A2(inbar[137]), .ZN(n655bar);
  OR2_X1 U312 ( .A1(in[149]), .A2(n654), .ZN(n656) );
  AND2_X1 U312bar ( .A1(inbar[149]), .A2(n654bar), .ZN(n656bar);
  OR2_X1 U313 ( .A1(in[195]), .A2(in[190]), .ZN(n654) );
  AND2_X1 U313bar ( .A1(inbar[195]), .A2(inbar[190]), .ZN(n654bar);
  OR2_X1 U314 ( .A1(n653), .A2(n652), .ZN(n704) );
  AND2_X1 U314bar ( .A1(n653bar), .A2(n652bar), .ZN(n704bar);
  OR2_X1 U315 ( .A1(n651), .A2(n650), .ZN(n652) );
  AND2_X1 U315bar ( .A1(n651bar), .A2(n650bar), .ZN(n652bar);
  OR2_X1 U316 ( .A1(in[98]), .A2(in[197]), .ZN(n650) );
  AND2_X1 U316bar ( .A1(inbar[98]), .A2(inbar[197]), .ZN(n650bar);
  OR2_X1 U317 ( .A1(in_11), .A2(n649), .ZN(n651) );
  AND2_X1 U317bar ( .A1(in_11bar), .A2(n649bar), .ZN(n651bar);
  OR2_X1 U318 ( .A1(in_26), .A2(in_14), .ZN(n649) );
  AND2_X1 U318bar ( .A1(in_26bar), .A2(in_14bar), .ZN(n649bar);
  OR2_X1 U319 ( .A1(n648), .A2(n647), .ZN(n653) );
  AND2_X1 U319bar ( .A1(n648bar), .A2(n647bar), .ZN(n653bar);
  OR2_X1 U320 ( .A1(in_35), .A2(in_27), .ZN(n647) );
  AND2_X1 U320bar ( .A1(in_35bar), .A2(in_27bar), .ZN(n647bar);
  OR2_X1 U321 ( .A1(in_50), .A2(n646), .ZN(n648) );
  AND2_X1 U321bar ( .A1(in_50bar), .A2(n646bar), .ZN(n648bar);
  OR2_X1 U322 ( .A1(in_78), .A2(in_61), .ZN(n646) );
  AND2_X1 U322bar ( .A1(in_78bar), .A2(in_61bar), .ZN(n646bar);
  OR2_X1 U323 ( .A1(n942), .A2(n645), .ZN(n720) );
  AND2_X1 U323bar ( .A1(n942bar), .A2(n645bar), .ZN(n720bar);
  OR2_X1 U324 ( .A1(in[106]), .A2(n863), .ZN(n645) );
  AND2_X1 U324bar ( .A1(inbar[106]), .A2(n863bar), .ZN(n645bar);
  OR2_X1 U325 ( .A1(n644), .A2(n643), .ZN(n863) );
  AND2_X1 U325bar ( .A1(n644bar), .A2(n643bar), .ZN(n863bar);
  OR2_X1 U326 ( .A1(n642), .A2(n641), .ZN(n643) );
  AND2_X1 U326bar ( .A1(n642bar), .A2(n641bar), .ZN(n643bar);
  OR2_X1 U327 ( .A1(n640), .A2(n639), .ZN(n641) );
  AND2_X1 U327bar ( .A1(n640bar), .A2(n639bar), .ZN(n641bar);
  OR2_X1 U328 ( .A1(in[127]), .A2(in[122]), .ZN(n639) );
  AND2_X1 U328bar ( .A1(inbar[127]), .A2(inbar[122]), .ZN(n639bar);
  OR2_X1 U329 ( .A1(in[156]), .A2(in[132]), .ZN(n640) );
  AND2_X1 U329bar ( .A1(inbar[156]), .A2(inbar[132]), .ZN(n640bar);
  OR2_X1 U330 ( .A1(n638), .A2(n637), .ZN(n642) );
  AND2_X1 U330bar ( .A1(n638bar), .A2(n637bar), .ZN(n642bar);
  OR2_X1 U331 ( .A1(in[159]), .A2(in[157]), .ZN(n637) );
  AND2_X1 U331bar ( .A1(inbar[159]), .A2(inbar[157]), .ZN(n637bar);
  OR2_X1 U332 ( .A1(in[185]), .A2(in[169]), .ZN(n638) );
  AND2_X1 U332bar ( .A1(inbar[185]), .A2(inbar[169]), .ZN(n638bar);
  OR2_X1 U333 ( .A1(n636), .A2(n635), .ZN(n644) );
  AND2_X1 U333bar ( .A1(n636bar), .A2(n635bar), .ZN(n644bar);
  OR2_X1 U334 ( .A1(n634), .A2(n633), .ZN(n635) );
  AND2_X1 U334bar ( .A1(n634bar), .A2(n633bar), .ZN(n635bar);
  OR2_X1 U335 ( .A1(in[239]), .A2(in[218]), .ZN(n633) );
  AND2_X1 U335bar ( .A1(inbar[239]), .A2(inbar[218]), .ZN(n633bar);
  OR2_X1 U336 ( .A1(in_13), .A2(in[87]), .ZN(n634) );
  AND2_X1 U336bar ( .A1(in_13bar), .A2(inbar[87]), .ZN(n634bar);
  OR2_X1 U337 ( .A1(n632), .A2(n631), .ZN(n636) );
  AND2_X1 U337bar ( .A1(n632bar), .A2(n631bar), .ZN(n636bar);
  OR2_X1 U338 ( .A1(in_72), .A2(in_70), .ZN(n631) );
  AND2_X1 U338bar ( .A1(in_72bar), .A2(in_70bar), .ZN(n631bar);
  OR2_X1 U339 ( .A1(in_80), .A2(in_74), .ZN(n632) );
  AND2_X1 U339bar ( .A1(in_80bar), .A2(in_74bar), .ZN(n632bar);
  OR2_X1 U340 ( .A1(n630), .A2(n629), .ZN(n942) );
  AND2_X1 U340bar ( .A1(n630bar), .A2(n629bar), .ZN(n942bar);
  OR2_X1 U341 ( .A1(n628), .A2(n627), .ZN(n629) );
  AND2_X1 U341bar ( .A1(n628bar), .A2(n627bar), .ZN(n629bar);
  OR2_X1 U342 ( .A1(n626), .A2(n625), .ZN(n627) );
  AND2_X1 U342bar ( .A1(n626bar), .A2(n625bar), .ZN(n627bar);
  OR2_X1 U343 ( .A1(in[146]), .A2(in[100]), .ZN(n625) );
  AND2_X1 U343bar ( .A1(inbar[146]), .A2(inbar[100]), .ZN(n625bar);
  OR2_X1 U344 ( .A1(in[168]), .A2(in[152]), .ZN(n626) );
  AND2_X1 U344bar ( .A1(inbar[168]), .A2(inbar[152]), .ZN(n626bar);
  OR2_X1 U345 ( .A1(n624), .A2(n623), .ZN(n628) );
  AND2_X1 U345bar ( .A1(n624bar), .A2(n623bar), .ZN(n628bar);
  OR2_X1 U346 ( .A1(in[199]), .A2(in[182]), .ZN(n623) );
  AND2_X1 U346bar ( .A1(inbar[199]), .A2(inbar[182]), .ZN(n623bar);
  OR2_X1 U347 ( .A1(in[236]), .A2(in[204]), .ZN(n624) );
  AND2_X1 U347bar ( .A1(inbar[236]), .A2(inbar[204]), .ZN(n624bar);
  OR2_X1 U348 ( .A1(n622), .A2(n621), .ZN(n630) );
  AND2_X1 U348bar ( .A1(n622bar), .A2(n621bar), .ZN(n630bar);
  OR2_X1 U349 ( .A1(n620), .A2(n619), .ZN(n621) );
  AND2_X1 U349bar ( .A1(n620bar), .A2(n619bar), .ZN(n621bar);
  OR2_X1 U350 ( .A1(in[89]), .A2(in[246]), .ZN(n619) );
  AND2_X1 U350bar ( .A1(inbar[89]), .A2(inbar[246]), .ZN(n619bar);
  OR2_X1 U351 ( .A1(in[95]), .A2(in[92]), .ZN(n620) );
  AND2_X1 U351bar ( .A1(inbar[95]), .A2(inbar[92]), .ZN(n620bar);
  OR2_X1 U352 ( .A1(n618), .A2(n617), .ZN(n622) );
  AND2_X1 U352bar ( .A1(n618bar), .A2(n617bar), .ZN(n622bar);
  OR2_X1 U353 ( .A1(in_22), .A2(in_16), .ZN(n617) );
  AND2_X1 U353bar ( .A1(in_22bar), .A2(in_16bar), .ZN(n617bar);
  OR2_X1 U354 ( .A1(in_51), .A2(in_49), .ZN(n618) );
  AND2_X1 U354bar ( .A1(in_51bar), .A2(in_49bar), .ZN(n618bar);
  OR2_X1 U355 ( .A1(n616), .A2(n615), .ZN(n722) );
  AND2_X1 U355bar ( .A1(n616bar), .A2(n615bar), .ZN(n722bar);
  OR2_X1 U356 ( .A1(in[158]), .A2(in[115]), .ZN(n615) );
  AND2_X1 U356bar ( .A1(inbar[158]), .A2(inbar[115]), .ZN(n615bar);
  OR2_X1 U357 ( .A1(in[163]), .A2(n614), .ZN(n616) );
  AND2_X1 U357bar ( .A1(inbar[163]), .A2(n614bar), .ZN(n616bar);
  OR2_X1 U358 ( .A1(in[206]), .A2(in[165]), .ZN(n614) );
  AND2_X1 U358bar ( .A1(inbar[206]), .A2(inbar[165]), .ZN(n614bar);
  OR2_X1 U359 ( .A1(n613), .A2(n612), .ZN(n724) );
  AND2_X1 U359bar ( .A1(n613bar), .A2(n612bar), .ZN(n724bar);
  OR2_X1 U360 ( .A1(n611), .A2(n610), .ZN(n612) );
  AND2_X1 U360bar ( .A1(n611bar), .A2(n610bar), .ZN(n612bar);
  OR2_X1 U361 ( .A1(in[213]), .A2(in[207]), .ZN(n610) );
  AND2_X1 U361bar ( .A1(inbar[213]), .A2(inbar[207]), .ZN(n610bar);
  OR2_X1 U362 ( .A1(in[215]), .A2(n609), .ZN(n611) );
  AND2_X1 U362bar ( .A1(inbar[215]), .A2(n609bar), .ZN(n611bar);
  OR2_X1 U363 ( .A1(in[230]), .A2(in[220]), .ZN(n609) );
  AND2_X1 U363bar ( .A1(inbar[230]), .A2(inbar[220]), .ZN(n609bar);
  OR2_X1 U364 ( .A1(n608), .A2(n607), .ZN(n613) );
  AND2_X1 U364bar ( .A1(n608bar), .A2(n607bar), .ZN(n613bar);
  OR2_X1 U365 ( .A1(in[251]), .A2(in[234]), .ZN(n607) );
  AND2_X1 U365bar ( .A1(inbar[251]), .A2(inbar[234]), .ZN(n607bar);
  OR2_X1 U366 ( .A1(in_17), .A2(n606), .ZN(n608) );
  AND2_X1 U366bar ( .A1(in_17bar), .A2(n606bar), .ZN(n608bar);
  OR2_X1 U367 ( .A1(in_65), .A2(in_56), .ZN(n606) );
  AND2_X1 U367bar ( .A1(in_65bar), .A2(in_56bar), .ZN(n606bar);
  OR2_X1 U368 ( .A1(n605), .A2(n604), .ZN(out[0]) );
  AND2_X1 U368bar ( .A1(n605bar), .A2(n604bar), .ZN(outbar[0]);
  OR2_X1 U369 ( .A1(n603), .A2(n602), .ZN(n604) );
  AND2_X1 U369bar ( .A1(n603bar), .A2(n602bar), .ZN(n604bar);
  OR2_X1 U370 ( .A1(n601), .A2(n600), .ZN(n602) );
  AND2_X1 U370bar ( .A1(n601bar), .A2(n600bar), .ZN(n602bar);
  OR2_X1 U371 ( .A1(n820), .A2(n785), .ZN(n600) );
  AND2_X1 U371bar ( .A1(n820bar), .A2(n785bar), .ZN(n600bar);
  OR2_X1 U372 ( .A1(n599), .A2(n598), .ZN(n785) );
  AND2_X1 U372bar ( .A1(n599bar), .A2(n598bar), .ZN(n785bar);
  OR2_X1 U373 ( .A1(n597), .A2(n596), .ZN(n598) );
  AND2_X1 U373bar ( .A1(n597bar), .A2(n596bar), .ZN(n598bar);
  OR2_X1 U374 ( .A1(n595), .A2(n594), .ZN(n596) );
  AND2_X1 U374bar ( .A1(n595bar), .A2(n594bar), .ZN(n596bar);
  OR2_X1 U375 ( .A1(in[135]), .A2(in[104]), .ZN(n594) );
  AND2_X1 U375bar ( .A1(inbar[135]), .A2(inbar[104]), .ZN(n594bar);
  OR2_X1 U376 ( .A1(in[188]), .A2(in[178]), .ZN(n595) );
  AND2_X1 U376bar ( .A1(inbar[188]), .A2(inbar[178]), .ZN(n595bar);
  OR2_X1 U377 ( .A1(n593), .A2(n592), .ZN(n597) );
  AND2_X1 U377bar ( .A1(n593bar), .A2(n592bar), .ZN(n597bar);
  OR2_X1 U378 ( .A1(in[217]), .A2(in[194]), .ZN(n592) );
  AND2_X1 U378bar ( .A1(inbar[217]), .A2(inbar[194]), .ZN(n592bar);
  OR2_X1 U379 ( .A1(in[237]), .A2(in[218]), .ZN(n593) );
  AND2_X1 U379bar ( .A1(inbar[237]), .A2(inbar[218]), .ZN(n593bar);
  OR2_X1 U380 ( .A1(n591), .A2(n590), .ZN(n599) );
  AND2_X1 U380bar ( .A1(n591bar), .A2(n590bar), .ZN(n599bar);
  OR2_X1 U381 ( .A1(n589), .A2(n588), .ZN(n590) );
  AND2_X1 U381bar ( .A1(n589bar), .A2(n588bar), .ZN(n590bar);
  OR2_X1 U382 ( .A1(in_2), .A2(in_10), .ZN(n588) );
  AND2_X1 U382bar ( .A1(in_2bar), .A2(in_10bar), .ZN(n588bar);
  OR2_X1 U383 ( .A1(in_47), .A2(in_22), .ZN(n589) );
  AND2_X1 U383bar ( .A1(in_47bar), .A2(in_22bar), .ZN(n589bar);
  OR2_X1 U384 ( .A1(n587), .A2(n586), .ZN(n591) );
  AND2_X1 U384bar ( .A1(n587bar), .A2(n586bar), .ZN(n591bar);
  OR2_X1 U385 ( .A1(in_56), .A2(in_54), .ZN(n586) );
  AND2_X1 U385bar ( .A1(in_56bar), .A2(in_54bar), .ZN(n586bar);
  OR2_X1 U386 ( .A1(in_63), .A2(in_61), .ZN(n587) );
  AND2_X1 U386bar ( .A1(in_63bar), .A2(in_61bar), .ZN(n587bar);
  OR2_X1 U387 ( .A1(n585), .A2(n584), .ZN(n820) );
  AND2_X1 U387bar ( .A1(n585bar), .A2(n584bar), .ZN(n820bar);
  OR2_X1 U388 ( .A1(n583), .A2(n582), .ZN(n584) );
  AND2_X1 U388bar ( .A1(n583bar), .A2(n582bar), .ZN(n584bar);
  OR2_X1 U389 ( .A1(n581), .A2(n580), .ZN(n582) );
  AND2_X1 U389bar ( .A1(n581bar), .A2(n580bar), .ZN(n582bar);
  OR2_X1 U390 ( .A1(in[158]), .A2(in[142]), .ZN(n580) );
  AND2_X1 U390bar ( .A1(inbar[158]), .A2(inbar[142]), .ZN(n580bar);
  OR2_X1 U391 ( .A1(in[175]), .A2(in[164]), .ZN(n581) );
  AND2_X1 U391bar ( .A1(inbar[175]), .A2(inbar[164]), .ZN(n581bar);
  OR2_X1 U392 ( .A1(n579), .A2(n578), .ZN(n583) );
  AND2_X1 U392bar ( .A1(n579bar), .A2(n578bar), .ZN(n583bar);
  OR2_X1 U393 ( .A1(in[228]), .A2(in[204]), .ZN(n578) );
  AND2_X1 U393bar ( .A1(inbar[228]), .A2(inbar[204]), .ZN(n578bar);
  OR2_X1 U394 ( .A1(in[91]), .A2(in[87]), .ZN(n579) );
  AND2_X1 U394bar ( .A1(inbar[91]), .A2(inbar[87]), .ZN(n579bar);
  OR2_X1 U395 ( .A1(n577), .A2(n576), .ZN(n585) );
  AND2_X1 U395bar ( .A1(n577bar), .A2(n576bar), .ZN(n585bar);
  OR2_X1 U396 ( .A1(n575), .A2(n574), .ZN(n576) );
  AND2_X1 U396bar ( .A1(n575bar), .A2(n574bar), .ZN(n576bar);
  OR2_X1 U397 ( .A1(in_21), .A2(in_11), .ZN(n574) );
  AND2_X1 U397bar ( .A1(in_21bar), .A2(in_11bar), .ZN(n574bar);
  OR2_X1 U398 ( .A1(in_5), .A2(in_3), .ZN(n575) );
  AND2_X1 U398bar ( .A1(in_5bar), .A2(in_3bar), .ZN(n575bar);
  OR2_X1 U399 ( .A1(n573), .A2(n572), .ZN(n577) );
  AND2_X1 U399bar ( .A1(n573bar), .A2(n572bar), .ZN(n577bar);
  OR2_X1 U400 ( .A1(in_68), .A2(in_64), .ZN(n572) );
  AND2_X1 U400bar ( .A1(in_68bar), .A2(in_64bar), .ZN(n572bar);
  OR2_X1 U401 ( .A1(in_76), .A2(in_73), .ZN(n573) );
  AND2_X1 U401bar ( .A1(in_76bar), .A2(in_73bar), .ZN(n573bar);
  OR2_X1 U402 ( .A1(n778), .A2(n571), .ZN(n601) );
  AND2_X1 U402bar ( .A1(n778bar), .A2(n571bar), .ZN(n601bar);
  OR2_X1 U403 ( .A1(in[100]), .A2(n965), .ZN(n571) );
  AND2_X1 U403bar ( .A1(inbar[100]), .A2(n965bar), .ZN(n571bar);
  OR2_X1 U404 ( .A1(n570), .A2(n569), .ZN(n965) );
  AND2_X1 U404bar ( .A1(n570bar), .A2(n569bar), .ZN(n965bar);
  OR2_X1 U405 ( .A1(n568), .A2(n567), .ZN(n569) );
  AND2_X1 U405bar ( .A1(n568bar), .A2(n567bar), .ZN(n569bar);
  OR2_X1 U406 ( .A1(n566), .A2(n565), .ZN(n567) );
  AND2_X1 U406bar ( .A1(n566bar), .A2(n565bar), .ZN(n567bar);
  OR2_X1 U407 ( .A1(n817), .A2(n750), .ZN(n565) );
  AND2_X1 U407bar ( .A1(n817bar), .A2(n750bar), .ZN(n565bar);
  OR2_X1 U408 ( .A1(n564), .A2(n563), .ZN(n750) );
  AND2_X1 U408bar ( .A1(n564bar), .A2(n563bar), .ZN(n750bar);
  OR2_X1 U409 ( .A1(n562), .A2(n561), .ZN(n563) );
  AND2_X1 U409bar ( .A1(n562bar), .A2(n561bar), .ZN(n563bar);
  OR2_X1 U410 ( .A1(n560), .A2(n559), .ZN(n561) );
  AND2_X1 U410bar ( .A1(n560bar), .A2(n559bar), .ZN(n561bar);
  OR2_X1 U411 ( .A1(in[119]), .A2(in[103]), .ZN(n559) );
  AND2_X1 U411bar ( .A1(inbar[119]), .A2(inbar[103]), .ZN(n559bar);
  OR2_X1 U412 ( .A1(in[137]), .A2(in[133]), .ZN(n560) );
  AND2_X1 U412bar ( .A1(inbar[137]), .A2(inbar[133]), .ZN(n560bar);
  OR2_X1 U413 ( .A1(n558), .A2(n557), .ZN(n562) );
  AND2_X1 U413bar ( .A1(n558bar), .A2(n557bar), .ZN(n562bar);
  OR2_X1 U414 ( .A1(in[176]), .A2(in[173]), .ZN(n557) );
  AND2_X1 U414bar ( .A1(inbar[176]), .A2(inbar[173]), .ZN(n557bar);
  OR2_X1 U415 ( .A1(in[210]), .A2(in[181]), .ZN(n558) );
  AND2_X1 U415bar ( .A1(inbar[210]), .A2(inbar[181]), .ZN(n558bar);
  OR2_X1 U416 ( .A1(n556), .A2(n555), .ZN(n564) );
  AND2_X1 U416bar ( .A1(n556bar), .A2(n555bar), .ZN(n564bar);
  OR2_X1 U417 ( .A1(n554), .A2(n553), .ZN(n555) );
  AND2_X1 U417bar ( .A1(n554bar), .A2(n553bar), .ZN(n555bar);
  OR2_X1 U418 ( .A1(in_13), .A2(in[234]), .ZN(n553) );
  AND2_X1 U418bar ( .A1(in_13bar), .A2(inbar[234]), .ZN(n553bar);
  OR2_X1 U419 ( .A1(in_38), .A2(in_32), .ZN(n554) );
  AND2_X1 U419bar ( .A1(in_38bar), .A2(in_32bar), .ZN(n554bar);
  OR2_X1 U420 ( .A1(n552), .A2(n551), .ZN(n556) );
  AND2_X1 U420bar ( .A1(n552bar), .A2(n551bar), .ZN(n556bar);
  OR2_X1 U421 ( .A1(in_42), .A2(in_41), .ZN(n551) );
  AND2_X1 U421bar ( .A1(in_42bar), .A2(in_41bar), .ZN(n551bar);
  OR2_X1 U422 ( .A1(in_7), .A2(in_49), .ZN(n552) );
  AND2_X1 U422bar ( .A1(in_7bar), .A2(in_49bar), .ZN(n552bar);
  OR2_X1 U423 ( .A1(n550), .A2(n549), .ZN(n817) );
  AND2_X1 U423bar ( .A1(n550bar), .A2(n549bar), .ZN(n817bar);
  OR2_X1 U424 ( .A1(n548), .A2(n547), .ZN(n549) );
  AND2_X1 U424bar ( .A1(n548bar), .A2(n547bar), .ZN(n549bar);
  OR2_X1 U425 ( .A1(n546), .A2(n545), .ZN(n547) );
  AND2_X1 U425bar ( .A1(n546bar), .A2(n545bar), .ZN(n547bar);
  OR2_X1 U426 ( .A1(in[159]), .A2(in[105]), .ZN(n545) );
  AND2_X1 U426bar ( .A1(inbar[159]), .A2(inbar[105]), .ZN(n545bar);
  OR2_X1 U427 ( .A1(in[206]), .A2(in[183]), .ZN(n546) );
  AND2_X1 U427bar ( .A1(inbar[206]), .A2(inbar[183]), .ZN(n546bar);
  OR2_X1 U428 ( .A1(n544), .A2(n543), .ZN(n548) );
  AND2_X1 U428bar ( .A1(n544bar), .A2(n543bar), .ZN(n548bar);
  OR2_X1 U429 ( .A1(in[229]), .A2(in[219]), .ZN(n543) );
  AND2_X1 U429bar ( .A1(inbar[229]), .A2(inbar[219]), .ZN(n543bar);
  OR2_X1 U430 ( .A1(in[235]), .A2(in[232]), .ZN(n544) );
  AND2_X1 U430bar ( .A1(inbar[235]), .A2(inbar[232]), .ZN(n544bar);
  OR2_X1 U431 ( .A1(n542), .A2(n541), .ZN(n550) );
  AND2_X1 U431bar ( .A1(n542bar), .A2(n541bar), .ZN(n550bar);
  OR2_X1 U432 ( .A1(n540), .A2(n539), .ZN(n541) );
  AND2_X1 U432bar ( .A1(n540bar), .A2(n539bar), .ZN(n541bar);
  OR2_X1 U433 ( .A1(in[249]), .A2(in[242]), .ZN(n539) );
  AND2_X1 U433bar ( .A1(inbar[249]), .A2(inbar[242]), .ZN(n539bar);
  OR2_X1 U434 ( .A1(in[89]), .A2(in[254]), .ZN(n540) );
  AND2_X1 U434bar ( .A1(inbar[89]), .A2(inbar[254]), .ZN(n540bar);
  OR2_X1 U435 ( .A1(n538), .A2(n537), .ZN(n542) );
  AND2_X1 U435bar ( .A1(n538bar), .A2(n537bar), .ZN(n542bar);
  OR2_X1 U436 ( .A1(in_14), .A2(in[99]), .ZN(n537) );
  AND2_X1 U436bar ( .A1(in_14bar), .A2(inbar[99]), .ZN(n537bar);
  OR2_X1 U437 ( .A1(in_60), .A2(in_18), .ZN(n538) );
  AND2_X1 U437bar ( .A1(in_60bar), .A2(in_18bar), .ZN(n538bar);
  OR2_X1 U438 ( .A1(in[113]), .A2(n763), .ZN(n566) );
  AND2_X1 U438bar ( .A1(inbar[113]), .A2(n763bar), .ZN(n566bar);
  OR2_X1 U439 ( .A1(n536), .A2(n535), .ZN(n763) );
  AND2_X1 U439bar ( .A1(n536bar), .A2(n535bar), .ZN(n763bar);
  OR2_X1 U440 ( .A1(n534), .A2(n533), .ZN(n535) );
  AND2_X1 U440bar ( .A1(n534bar), .A2(n533bar), .ZN(n535bar);
  OR2_X1 U441 ( .A1(n532), .A2(n531), .ZN(n533) );
  AND2_X1 U441bar ( .A1(n532bar), .A2(n531bar), .ZN(n533bar);
  OR2_X1 U442 ( .A1(in[115]), .A2(in[110]), .ZN(n531) );
  AND2_X1 U442bar ( .A1(inbar[115]), .A2(inbar[110]), .ZN(n531bar);
  OR2_X1 U443 ( .A1(in[125]), .A2(in[117]), .ZN(n532) );
  AND2_X1 U443bar ( .A1(inbar[125]), .A2(inbar[117]), .ZN(n532bar);
  OR2_X1 U444 ( .A1(n530), .A2(n529), .ZN(n534) );
  AND2_X1 U444bar ( .A1(n530bar), .A2(n529bar), .ZN(n534bar);
  OR2_X1 U445 ( .A1(in[180]), .A2(in[128]), .ZN(n529) );
  AND2_X1 U445bar ( .A1(inbar[180]), .A2(inbar[128]), .ZN(n529bar);
  OR2_X1 U446 ( .A1(in[205]), .A2(in[201]), .ZN(n530) );
  AND2_X1 U446bar ( .A1(inbar[205]), .A2(inbar[201]), .ZN(n530bar);
  OR2_X1 U447 ( .A1(n528), .A2(n527), .ZN(n536) );
  AND2_X1 U447bar ( .A1(n528bar), .A2(n527bar), .ZN(n536bar);
  OR2_X1 U448 ( .A1(n526), .A2(n525), .ZN(n527) );
  AND2_X1 U448bar ( .A1(n526bar), .A2(n525bar), .ZN(n527bar);
  OR2_X1 U449 ( .A1(in[244]), .A2(in[239]), .ZN(n525) );
  AND2_X1 U449bar ( .A1(inbar[244]), .A2(inbar[239]), .ZN(n525bar);
  OR2_X1 U450 ( .A1(in[95]), .A2(in[83]), .ZN(n526) );
  AND2_X1 U450bar ( .A1(inbar[95]), .A2(inbar[83]), .ZN(n526bar);
  OR2_X1 U451 ( .A1(n524), .A2(n523), .ZN(n528) );
  AND2_X1 U451bar ( .A1(n524bar), .A2(n523bar), .ZN(n528bar);
  OR2_X1 U452 ( .A1(in_24), .A2(in[97]), .ZN(n523) );
  AND2_X1 U452bar ( .A1(in_24bar), .A2(inbar[97]), .ZN(n523bar);
  OR2_X1 U453 ( .A1(in_33), .A2(in_27), .ZN(n524) );
  AND2_X1 U453bar ( .A1(in_33bar), .A2(in_27bar), .ZN(n524bar);
  OR2_X1 U454 ( .A1(n522), .A2(n521), .ZN(n568) );
  AND2_X1 U454bar ( .A1(n522bar), .A2(n521bar), .ZN(n568bar);
  OR2_X1 U455 ( .A1(in[145]), .A2(in[126]), .ZN(n521) );
  AND2_X1 U455bar ( .A1(inbar[145]), .A2(inbar[126]), .ZN(n521bar);
  OR2_X1 U456 ( .A1(in[169]), .A2(n520), .ZN(n522) );
  AND2_X1 U456bar ( .A1(inbar[169]), .A2(n520bar), .ZN(n522bar);
  OR2_X1 U457 ( .A1(in[221]), .A2(in[172]), .ZN(n520) );
  AND2_X1 U457bar ( .A1(inbar[221]), .A2(inbar[172]), .ZN(n520bar);
  OR2_X1 U458 ( .A1(n519), .A2(n518), .ZN(n570) );
  AND2_X1 U458bar ( .A1(n519bar), .A2(n518bar), .ZN(n570bar);
  OR2_X1 U459 ( .A1(n517), .A2(n516), .ZN(n518) );
  AND2_X1 U459bar ( .A1(n517bar), .A2(n516bar), .ZN(n518bar);
  OR2_X1 U460 ( .A1(in[241]), .A2(in[224]), .ZN(n516) );
  AND2_X1 U460bar ( .A1(inbar[241]), .A2(inbar[224]), .ZN(n516bar);
  OR2_X1 U461 ( .A1(in[86]), .A2(n515), .ZN(n517) );
  AND2_X1 U461bar ( .A1(inbar[86]), .A2(n515bar), .ZN(n517bar);
  OR2_X1 U462 ( .A1(in_43), .A2(in_34), .ZN(n515) );
  AND2_X1 U462bar ( .A1(in_43bar), .A2(in_34bar), .ZN(n515bar);
  OR2_X1 U463 ( .A1(n514), .A2(n513), .ZN(n519) );
  AND2_X1 U463bar ( .A1(n514bar), .A2(n513bar), .ZN(n519bar);
  OR2_X1 U464 ( .A1(in_65), .A2(in_51), .ZN(n513) );
  AND2_X1 U464bar ( .A1(in_65bar), .A2(in_51bar), .ZN(n513bar);
  OR2_X1 U465 ( .A1(in_75), .A2(n512), .ZN(n514) );
  AND2_X1 U465bar ( .A1(in_75bar), .A2(n512bar), .ZN(n514bar);
  OR2_X1 U466 ( .A1(in_81), .A2(in_77), .ZN(n512) );
  AND2_X1 U466bar ( .A1(in_81bar), .A2(in_77bar), .ZN(n512bar);
  OR2_X1 U467 ( .A1(n511), .A2(n510), .ZN(n778) );
  AND2_X1 U467bar ( .A1(n511bar), .A2(n510bar), .ZN(n778bar);
  OR2_X1 U468 ( .A1(n509), .A2(n508), .ZN(n510) );
  AND2_X1 U468bar ( .A1(n509bar), .A2(n508bar), .ZN(n510bar);
  OR2_X1 U469 ( .A1(n507), .A2(n506), .ZN(n508) );
  AND2_X1 U469bar ( .A1(n507bar), .A2(n506bar), .ZN(n508bar);
  OR2_X1 U470 ( .A1(in[107]), .A2(in[101]), .ZN(n506) );
  AND2_X1 U470bar ( .A1(inbar[107]), .A2(inbar[101]), .ZN(n506bar);
  OR2_X1 U471 ( .A1(in[139]), .A2(in[132]), .ZN(n507) );
  AND2_X1 U471bar ( .A1(inbar[139]), .A2(inbar[132]), .ZN(n507bar);
  OR2_X1 U472 ( .A1(n505), .A2(n504), .ZN(n509) );
  AND2_X1 U472bar ( .A1(n505bar), .A2(n504bar), .ZN(n509bar);
  OR2_X1 U473 ( .A1(in[146]), .A2(in[141]), .ZN(n504) );
  AND2_X1 U473bar ( .A1(inbar[146]), .A2(inbar[141]), .ZN(n504bar);
  OR2_X1 U474 ( .A1(in[203]), .A2(in[179]), .ZN(n505) );
  AND2_X1 U474bar ( .A1(inbar[203]), .A2(inbar[179]), .ZN(n505bar);
  OR2_X1 U475 ( .A1(n503), .A2(n502), .ZN(n511) );
  AND2_X1 U475bar ( .A1(n503bar), .A2(n502bar), .ZN(n511bar);
  OR2_X1 U476 ( .A1(n501), .A2(n500), .ZN(n502) );
  AND2_X1 U476bar ( .A1(n501bar), .A2(n500bar), .ZN(n502bar);
  OR2_X1 U477 ( .A1(in[243]), .A2(in[222]), .ZN(n500) );
  AND2_X1 U477bar ( .A1(inbar[243]), .A2(inbar[222]), .ZN(n500bar);
  OR2_X1 U478 ( .A1(in[251]), .A2(in[250]), .ZN(n501) );
  AND2_X1 U478bar ( .A1(inbar[251]), .A2(inbar[250]), .ZN(n501bar);
  OR2_X1 U479 ( .A1(n499), .A2(n498), .ZN(n503) );
  AND2_X1 U479bar ( .A1(n499bar), .A2(n498bar), .ZN(n503bar);
  OR2_X1 U480 ( .A1(in_37), .A2(in_19), .ZN(n498) );
  AND2_X1 U480bar ( .A1(in_37bar), .A2(in_19bar), .ZN(n498bar);
  OR2_X1 U481 ( .A1(in_78), .A2(in_6), .ZN(n499) );
  AND2_X1 U481bar ( .A1(in_78bar), .A2(in_6bar), .ZN(n499bar);
  OR2_X1 U482 ( .A1(n497), .A2(n496), .ZN(n603) );
  AND2_X1 U482bar ( .A1(n497bar), .A2(n496bar), .ZN(n603bar);
  OR2_X1 U483 ( .A1(in[112]), .A2(in[102]), .ZN(n496) );
  AND2_X1 U483bar ( .A1(inbar[112]), .A2(inbar[102]), .ZN(n496bar);
  OR2_X1 U484 ( .A1(in[123]), .A2(n495), .ZN(n497) );
  AND2_X1 U484bar ( .A1(inbar[123]), .A2(n495bar), .ZN(n497bar);
  OR2_X1 U485 ( .A1(in[143]), .A2(in[130]), .ZN(n495) );
  AND2_X1 U485bar ( .A1(inbar[143]), .A2(inbar[130]), .ZN(n495bar);
  OR2_X1 U486 ( .A1(n494), .A2(n493), .ZN(n605) );
  AND2_X1 U486bar ( .A1(n494bar), .A2(n493bar), .ZN(n605bar);
  OR2_X1 U487 ( .A1(n492), .A2(n491), .ZN(n493) );
  AND2_X1 U487bar ( .A1(n492bar), .A2(n491bar), .ZN(n493bar);
  OR2_X1 U488 ( .A1(in[216]), .A2(in[213]), .ZN(n491) );
  AND2_X1 U488bar ( .A1(inbar[216]), .A2(inbar[213]), .ZN(n491bar);
  OR2_X1 U489 ( .A1(in[227]), .A2(n490), .ZN(n492) );
  AND2_X1 U489bar ( .A1(inbar[227]), .A2(n490bar), .ZN(n492bar);
  OR2_X1 U490 ( .A1(in_0), .A2(in[248]), .ZN(n490) );
  AND2_X1 U490bar ( .A1(in_0bar), .A2(inbar[248]), .ZN(n490bar);
  OR2_X1 U491 ( .A1(n489), .A2(n488), .ZN(n494) );
  AND2_X1 U491bar ( .A1(n489bar), .A2(n488bar), .ZN(n494bar);
  OR2_X1 U492 ( .A1(in_46), .A2(in_44), .ZN(n488) );
  AND2_X1 U492bar ( .A1(in_46bar), .A2(in_44bar), .ZN(n488bar);
  OR2_X1 U493 ( .A1(in_50), .A2(n487), .ZN(n489) );
  AND2_X1 U493bar ( .A1(in_50bar), .A2(n487bar), .ZN(n489bar);
  OR2_X1 U494 ( .A1(in_9), .A2(in_80), .ZN(n487) );
  AND2_X1 U494bar ( .A1(in_9bar), .A2(in_80bar), .ZN(n487bar);
endmodule




module sBox_6 ( in, out );
  input [7:0] in;
  //input_done

  output [7:0] out;
  //output_done

  wire   [255:0] decodeOut;
  //wire_done

  decode_6 dec ( .in(in), .out(decodeOut) );
  encode_6 enc ( .in(decodeOut), .out(out) );
endmodule


module CD2_25 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_26 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_27 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_28 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD4_13 ( a, b, y );
  input [3:0] a;
  input [3:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  //input_done

  output [15:0] y;
  reg [15:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]);
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]);
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]);
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]);
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]);
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]);
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]);
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]);
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]);
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]);
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]);
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]);
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]);
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]);
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]);
endmodule




module CD4_14 ( a, b, y );
  input [3:0] a;
  input [3:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  //input_done

  output [15:0] y;
  reg [15:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]);
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]);
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]);
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]);
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]);
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]);
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]);
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]);
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]);
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]);
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]);
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]);
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]);
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]);
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]);
endmodule




module CD16_7 ( a, b, y );
  input [15:0] a;
  input [15:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign abar[8] = ~a[8];
  assign abar[9] = ~a[9];
  assign abar[10] = ~a[10];
  assign abar[11] = ~a[11];
  assign abar[12] = ~a[12];
  assign abar[13] = ~a[13];
  assign abar[14] = ~a[14];
  assign abar[15] = ~a[15];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign bbar[8] = ~b[8];
  assign bbar[9] = ~b[9];
  assign bbar[10] = ~b[10];
  assign bbar[11] = ~b[11];
  assign bbar[12] = ~b[12];
  assign bbar[13] = ~b[13];
  assign bbar[14] = ~b[14];
  assign bbar[15] = ~b[15];
  //input_done

  output [255:0] y;
  reg [255:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[9]), .A2(a[0]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[9]), .A2(abar[0]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[3]), .A2(a[6]), .ZN(y[99]) );
  OR2_X1 U2bar ( .A1(bbar[3]), .A2(abar[6]), .ZN(ybar[99]);
  AND2_X1 U3 ( .A1(b[2]), .A2(a[6]), .ZN(y[98]) );
  OR2_X1 U3bar ( .A1(bbar[2]), .A2(abar[6]), .ZN(ybar[98]);
  AND2_X1 U4 ( .A1(b[1]), .A2(a[6]), .ZN(y[97]) );
  OR2_X1 U4bar ( .A1(bbar[1]), .A2(abar[6]), .ZN(ybar[97]);
  AND2_X1 U5 ( .A1(b[0]), .A2(a[6]), .ZN(y[96]) );
  OR2_X1 U5bar ( .A1(bbar[0]), .A2(abar[6]), .ZN(ybar[96]);
  AND2_X1 U6 ( .A1(b[15]), .A2(a[5]), .ZN(y[95]) );
  OR2_X1 U6bar ( .A1(bbar[15]), .A2(abar[5]), .ZN(ybar[95]);
  AND2_X1 U7 ( .A1(b[14]), .A2(a[5]), .ZN(y[94]) );
  OR2_X1 U7bar ( .A1(bbar[14]), .A2(abar[5]), .ZN(ybar[94]);
  AND2_X1 U8 ( .A1(b[13]), .A2(a[5]), .ZN(y[93]) );
  OR2_X1 U8bar ( .A1(bbar[13]), .A2(abar[5]), .ZN(ybar[93]);
  AND2_X1 U9 ( .A1(b[12]), .A2(a[5]), .ZN(y[92]) );
  OR2_X1 U9bar ( .A1(bbar[12]), .A2(abar[5]), .ZN(ybar[92]);
  AND2_X1 U10 ( .A1(b[11]), .A2(a[5]), .ZN(y[91]) );
  OR2_X1 U10bar ( .A1(bbar[11]), .A2(abar[5]), .ZN(ybar[91]);
  AND2_X1 U11 ( .A1(b[10]), .A2(a[5]), .ZN(y[90]) );
  OR2_X1 U11bar ( .A1(bbar[10]), .A2(abar[5]), .ZN(ybar[90]);
  AND2_X1 U12 ( .A1(b[8]), .A2(a[0]), .ZN(y[8]) );
  OR2_X1 U12bar ( .A1(bbar[8]), .A2(abar[0]), .ZN(ybar[8]);
  AND2_X1 U13 ( .A1(a[5]), .A2(b[9]), .ZN(y[89]) );
  OR2_X1 U13bar ( .A1(abar[5]), .A2(bbar[9]), .ZN(ybar[89]);
  AND2_X1 U14 ( .A1(b[8]), .A2(a[5]), .ZN(y[88]) );
  OR2_X1 U14bar ( .A1(bbar[8]), .A2(abar[5]), .ZN(ybar[88]);
  AND2_X1 U15 ( .A1(b[7]), .A2(a[5]), .ZN(y[87]) );
  OR2_X1 U15bar ( .A1(bbar[7]), .A2(abar[5]), .ZN(ybar[87]);
  AND2_X1 U16 ( .A1(b[6]), .A2(a[5]), .ZN(y[86]) );
  OR2_X1 U16bar ( .A1(bbar[6]), .A2(abar[5]), .ZN(ybar[86]);
  AND2_X1 U17 ( .A1(b[5]), .A2(a[5]), .ZN(y[85]) );
  OR2_X1 U17bar ( .A1(bbar[5]), .A2(abar[5]), .ZN(ybar[85]);
  AND2_X1 U18 ( .A1(b[4]), .A2(a[5]), .ZN(y[84]) );
  OR2_X1 U18bar ( .A1(bbar[4]), .A2(abar[5]), .ZN(ybar[84]);
  AND2_X1 U19 ( .A1(a[5]), .A2(b[3]), .ZN(y[83]) );
  OR2_X1 U19bar ( .A1(abar[5]), .A2(bbar[3]), .ZN(ybar[83]);
  AND2_X1 U20 ( .A1(a[5]), .A2(b[2]), .ZN(y[82]) );
  OR2_X1 U20bar ( .A1(abar[5]), .A2(bbar[2]), .ZN(ybar[82]);
  AND2_X1 U21 ( .A1(a[5]), .A2(b[1]), .ZN(y[81]) );
  OR2_X1 U21bar ( .A1(abar[5]), .A2(bbar[1]), .ZN(ybar[81]);
  AND2_X1 U22 ( .A1(a[5]), .A2(b[0]), .ZN(y[80]) );
  OR2_X1 U22bar ( .A1(abar[5]), .A2(bbar[0]), .ZN(ybar[80]);
  AND2_X1 U23 ( .A1(b[7]), .A2(a[0]), .ZN(y[7]) );
  OR2_X1 U23bar ( .A1(bbar[7]), .A2(abar[0]), .ZN(ybar[7]);
  AND2_X1 U24 ( .A1(a[4]), .A2(b[15]), .ZN(y[79]) );
  OR2_X1 U24bar ( .A1(abar[4]), .A2(bbar[15]), .ZN(ybar[79]);
  AND2_X1 U25 ( .A1(a[4]), .A2(b[14]), .ZN(y[78]) );
  OR2_X1 U25bar ( .A1(abar[4]), .A2(bbar[14]), .ZN(ybar[78]);
  AND2_X1 U26 ( .A1(a[4]), .A2(b[13]), .ZN(y[77]) );
  OR2_X1 U26bar ( .A1(abar[4]), .A2(bbar[13]), .ZN(ybar[77]);
  AND2_X1 U27 ( .A1(a[4]), .A2(b[12]), .ZN(y[76]) );
  OR2_X1 U27bar ( .A1(abar[4]), .A2(bbar[12]), .ZN(ybar[76]);
  AND2_X1 U28 ( .A1(a[4]), .A2(b[11]), .ZN(y[75]) );
  OR2_X1 U28bar ( .A1(abar[4]), .A2(bbar[11]), .ZN(ybar[75]);
  AND2_X1 U29 ( .A1(a[4]), .A2(b[10]), .ZN(y[74]) );
  OR2_X1 U29bar ( .A1(abar[4]), .A2(bbar[10]), .ZN(ybar[74]);
  AND2_X1 U30 ( .A1(a[4]), .A2(b[9]), .ZN(y[73]) );
  OR2_X1 U30bar ( .A1(abar[4]), .A2(bbar[9]), .ZN(ybar[73]);
  AND2_X1 U31 ( .A1(a[4]), .A2(b[8]), .ZN(y[72]) );
  OR2_X1 U31bar ( .A1(abar[4]), .A2(bbar[8]), .ZN(ybar[72]);
  AND2_X1 U32 ( .A1(a[4]), .A2(b[7]), .ZN(y[71]) );
  OR2_X1 U32bar ( .A1(abar[4]), .A2(bbar[7]), .ZN(ybar[71]);
  AND2_X1 U33 ( .A1(a[4]), .A2(b[6]), .ZN(y[70]) );
  OR2_X1 U33bar ( .A1(abar[4]), .A2(bbar[6]), .ZN(ybar[70]);
  AND2_X1 U34 ( .A1(b[6]), .A2(a[0]), .ZN(y[6]) );
  OR2_X1 U34bar ( .A1(bbar[6]), .A2(abar[0]), .ZN(ybar[6]);
  AND2_X1 U35 ( .A1(a[4]), .A2(b[5]), .ZN(y[69]) );
  OR2_X1 U35bar ( .A1(abar[4]), .A2(bbar[5]), .ZN(ybar[69]);
  AND2_X1 U36 ( .A1(a[4]), .A2(b[4]), .ZN(y[68]) );
  OR2_X1 U36bar ( .A1(abar[4]), .A2(bbar[4]), .ZN(ybar[68]);
  AND2_X1 U37 ( .A1(a[4]), .A2(b[3]), .ZN(y[67]) );
  OR2_X1 U37bar ( .A1(abar[4]), .A2(bbar[3]), .ZN(ybar[67]);
  AND2_X1 U38 ( .A1(a[4]), .A2(b[2]), .ZN(y[66]) );
  OR2_X1 U38bar ( .A1(abar[4]), .A2(bbar[2]), .ZN(ybar[66]);
  AND2_X1 U39 ( .A1(a[4]), .A2(b[1]), .ZN(y[65]) );
  OR2_X1 U39bar ( .A1(abar[4]), .A2(bbar[1]), .ZN(ybar[65]);
  AND2_X1 U40 ( .A1(a[4]), .A2(b[0]), .ZN(y[64]) );
  OR2_X1 U40bar ( .A1(abar[4]), .A2(bbar[0]), .ZN(ybar[64]);
  AND2_X1 U41 ( .A1(a[3]), .A2(b[15]), .ZN(y[63]) );
  OR2_X1 U41bar ( .A1(abar[3]), .A2(bbar[15]), .ZN(ybar[63]);
  AND2_X1 U42 ( .A1(a[3]), .A2(b[14]), .ZN(y[62]) );
  OR2_X1 U42bar ( .A1(abar[3]), .A2(bbar[14]), .ZN(ybar[62]);
  AND2_X1 U43 ( .A1(a[3]), .A2(b[13]), .ZN(y[61]) );
  OR2_X1 U43bar ( .A1(abar[3]), .A2(bbar[13]), .ZN(ybar[61]);
  AND2_X1 U44 ( .A1(a[3]), .A2(b[12]), .ZN(y[60]) );
  OR2_X1 U44bar ( .A1(abar[3]), .A2(bbar[12]), .ZN(ybar[60]);
  AND2_X1 U45 ( .A1(b[5]), .A2(a[0]), .ZN(y[5]) );
  OR2_X1 U45bar ( .A1(bbar[5]), .A2(abar[0]), .ZN(ybar[5]);
  AND2_X1 U46 ( .A1(a[3]), .A2(b[11]), .ZN(y[59]) );
  OR2_X1 U46bar ( .A1(abar[3]), .A2(bbar[11]), .ZN(ybar[59]);
  AND2_X1 U47 ( .A1(a[3]), .A2(b[10]), .ZN(y[58]) );
  OR2_X1 U47bar ( .A1(abar[3]), .A2(bbar[10]), .ZN(ybar[58]);
  AND2_X1 U48 ( .A1(a[3]), .A2(b[9]), .ZN(y[57]) );
  OR2_X1 U48bar ( .A1(abar[3]), .A2(bbar[9]), .ZN(ybar[57]);
  AND2_X1 U49 ( .A1(a[3]), .A2(b[8]), .ZN(y[56]) );
  OR2_X1 U49bar ( .A1(abar[3]), .A2(bbar[8]), .ZN(ybar[56]);
  AND2_X1 U50 ( .A1(a[3]), .A2(b[7]), .ZN(y[55]) );
  OR2_X1 U50bar ( .A1(abar[3]), .A2(bbar[7]), .ZN(ybar[55]);
  AND2_X1 U51 ( .A1(a[3]), .A2(b[6]), .ZN(y[54]) );
  OR2_X1 U51bar ( .A1(abar[3]), .A2(bbar[6]), .ZN(ybar[54]);
  AND2_X1 U52 ( .A1(a[3]), .A2(b[5]), .ZN(y[53]) );
  OR2_X1 U52bar ( .A1(abar[3]), .A2(bbar[5]), .ZN(ybar[53]);
  AND2_X1 U53 ( .A1(a[3]), .A2(b[4]), .ZN(y[52]) );
  OR2_X1 U53bar ( .A1(abar[3]), .A2(bbar[4]), .ZN(ybar[52]);
  AND2_X1 U54 ( .A1(a[3]), .A2(b[3]), .ZN(y[51]) );
  OR2_X1 U54bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[51]);
  AND2_X1 U55 ( .A1(a[3]), .A2(b[2]), .ZN(y[50]) );
  OR2_X1 U55bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[50]);
  AND2_X1 U56 ( .A1(b[4]), .A2(a[0]), .ZN(y[4]) );
  OR2_X1 U56bar ( .A1(bbar[4]), .A2(abar[0]), .ZN(ybar[4]);
  AND2_X1 U57 ( .A1(a[3]), .A2(b[1]), .ZN(y[49]) );
  OR2_X1 U57bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[49]);
  AND2_X1 U58 ( .A1(a[3]), .A2(b[0]), .ZN(y[48]) );
  OR2_X1 U58bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[48]);
  AND2_X1 U59 ( .A1(a[2]), .A2(b[15]), .ZN(y[47]) );
  OR2_X1 U59bar ( .A1(abar[2]), .A2(bbar[15]), .ZN(ybar[47]);
  AND2_X1 U60 ( .A1(a[2]), .A2(b[14]), .ZN(y[46]) );
  OR2_X1 U60bar ( .A1(abar[2]), .A2(bbar[14]), .ZN(ybar[46]);
  AND2_X1 U61 ( .A1(a[2]), .A2(b[13]), .ZN(y[45]) );
  OR2_X1 U61bar ( .A1(abar[2]), .A2(bbar[13]), .ZN(ybar[45]);
  AND2_X1 U62 ( .A1(a[2]), .A2(b[12]), .ZN(y[44]) );
  OR2_X1 U62bar ( .A1(abar[2]), .A2(bbar[12]), .ZN(ybar[44]);
  AND2_X1 U63 ( .A1(a[2]), .A2(b[11]), .ZN(y[43]) );
  OR2_X1 U63bar ( .A1(abar[2]), .A2(bbar[11]), .ZN(ybar[43]);
  AND2_X1 U64 ( .A1(a[2]), .A2(b[10]), .ZN(y[42]) );
  OR2_X1 U64bar ( .A1(abar[2]), .A2(bbar[10]), .ZN(ybar[42]);
  AND2_X1 U65 ( .A1(a[2]), .A2(b[9]), .ZN(y[41]) );
  OR2_X1 U65bar ( .A1(abar[2]), .A2(bbar[9]), .ZN(ybar[41]);
  AND2_X1 U66 ( .A1(a[2]), .A2(b[8]), .ZN(y[40]) );
  OR2_X1 U66bar ( .A1(abar[2]), .A2(bbar[8]), .ZN(ybar[40]);
  AND2_X1 U67 ( .A1(b[3]), .A2(a[0]), .ZN(y[3]) );
  OR2_X1 U67bar ( .A1(bbar[3]), .A2(abar[0]), .ZN(ybar[3]);
  AND2_X1 U68 ( .A1(a[2]), .A2(b[7]), .ZN(y[39]) );
  OR2_X1 U68bar ( .A1(abar[2]), .A2(bbar[7]), .ZN(ybar[39]);
  AND2_X1 U69 ( .A1(a[2]), .A2(b[6]), .ZN(y[38]) );
  OR2_X1 U69bar ( .A1(abar[2]), .A2(bbar[6]), .ZN(ybar[38]);
  AND2_X1 U70 ( .A1(a[2]), .A2(b[5]), .ZN(y[37]) );
  OR2_X1 U70bar ( .A1(abar[2]), .A2(bbar[5]), .ZN(ybar[37]);
  AND2_X1 U71 ( .A1(a[2]), .A2(b[4]), .ZN(y[36]) );
  OR2_X1 U71bar ( .A1(abar[2]), .A2(bbar[4]), .ZN(ybar[36]);
  AND2_X1 U72 ( .A1(a[2]), .A2(b[3]), .ZN(y[35]) );
  OR2_X1 U72bar ( .A1(abar[2]), .A2(bbar[3]), .ZN(ybar[35]);
  AND2_X1 U73 ( .A1(a[2]), .A2(b[2]), .ZN(y[34]) );
  OR2_X1 U73bar ( .A1(abar[2]), .A2(bbar[2]), .ZN(ybar[34]);
  AND2_X1 U74 ( .A1(a[2]), .A2(b[1]), .ZN(y[33]) );
  OR2_X1 U74bar ( .A1(abar[2]), .A2(bbar[1]), .ZN(ybar[33]);
  AND2_X1 U75 ( .A1(a[2]), .A2(b[0]), .ZN(y[32]) );
  OR2_X1 U75bar ( .A1(abar[2]), .A2(bbar[0]), .ZN(ybar[32]);
  AND2_X1 U76 ( .A1(a[1]), .A2(b[15]), .ZN(y[31]) );
  OR2_X1 U76bar ( .A1(abar[1]), .A2(bbar[15]), .ZN(ybar[31]);
  AND2_X1 U77 ( .A1(a[1]), .A2(b[14]), .ZN(y[30]) );
  OR2_X1 U77bar ( .A1(abar[1]), .A2(bbar[14]), .ZN(ybar[30]);
  AND2_X1 U78 ( .A1(b[2]), .A2(a[0]), .ZN(y[2]) );
  OR2_X1 U78bar ( .A1(bbar[2]), .A2(abar[0]), .ZN(ybar[2]);
  AND2_X1 U79 ( .A1(a[1]), .A2(b[13]), .ZN(y[29]) );
  OR2_X1 U79bar ( .A1(abar[1]), .A2(bbar[13]), .ZN(ybar[29]);
  AND2_X1 U80 ( .A1(a[1]), .A2(b[12]), .ZN(y[28]) );
  OR2_X1 U80bar ( .A1(abar[1]), .A2(bbar[12]), .ZN(ybar[28]);
  AND2_X1 U81 ( .A1(a[1]), .A2(b[11]), .ZN(y[27]) );
  OR2_X1 U81bar ( .A1(abar[1]), .A2(bbar[11]), .ZN(ybar[27]);
  AND2_X1 U82 ( .A1(a[1]), .A2(b[10]), .ZN(y[26]) );
  OR2_X1 U82bar ( .A1(abar[1]), .A2(bbar[10]), .ZN(ybar[26]);
  AND2_X1 U83 ( .A1(a[1]), .A2(b[9]), .ZN(y[25]) );
  OR2_X1 U83bar ( .A1(abar[1]), .A2(bbar[9]), .ZN(ybar[25]);
  AND2_X1 U84 ( .A1(a[15]), .A2(b[15]), .ZN(y[255]) );
  OR2_X1 U84bar ( .A1(abar[15]), .A2(bbar[15]), .ZN(ybar[255]);
  AND2_X1 U85 ( .A1(a[15]), .A2(b[14]), .ZN(y[254]) );
  OR2_X1 U85bar ( .A1(abar[15]), .A2(bbar[14]), .ZN(ybar[254]);
  AND2_X1 U86 ( .A1(a[15]), .A2(b[13]), .ZN(y[253]) );
  OR2_X1 U86bar ( .A1(abar[15]), .A2(bbar[13]), .ZN(ybar[253]);
  AND2_X1 U87 ( .A1(a[15]), .A2(b[12]), .ZN(y[252]) );
  OR2_X1 U87bar ( .A1(abar[15]), .A2(bbar[12]), .ZN(ybar[252]);
  AND2_X1 U88 ( .A1(a[15]), .A2(b[11]), .ZN(y[251]) );
  OR2_X1 U88bar ( .A1(abar[15]), .A2(bbar[11]), .ZN(ybar[251]);
  AND2_X1 U89 ( .A1(a[15]), .A2(b[10]), .ZN(y[250]) );
  OR2_X1 U89bar ( .A1(abar[15]), .A2(bbar[10]), .ZN(ybar[250]);
  AND2_X1 U90 ( .A1(a[1]), .A2(b[8]), .ZN(y[24]) );
  OR2_X1 U90bar ( .A1(abar[1]), .A2(bbar[8]), .ZN(ybar[24]);
  AND2_X1 U91 ( .A1(a[15]), .A2(b[9]), .ZN(y[249]) );
  OR2_X1 U91bar ( .A1(abar[15]), .A2(bbar[9]), .ZN(ybar[249]);
  AND2_X1 U92 ( .A1(a[15]), .A2(b[8]), .ZN(y[248]) );
  OR2_X1 U92bar ( .A1(abar[15]), .A2(bbar[8]), .ZN(ybar[248]);
  AND2_X1 U93 ( .A1(a[15]), .A2(b[7]), .ZN(y[247]) );
  OR2_X1 U93bar ( .A1(abar[15]), .A2(bbar[7]), .ZN(ybar[247]);
  AND2_X1 U94 ( .A1(a[15]), .A2(b[6]), .ZN(y[246]) );
  OR2_X1 U94bar ( .A1(abar[15]), .A2(bbar[6]), .ZN(ybar[246]);
  AND2_X1 U95 ( .A1(a[15]), .A2(b[5]), .ZN(y[245]) );
  OR2_X1 U95bar ( .A1(abar[15]), .A2(bbar[5]), .ZN(ybar[245]);
  AND2_X1 U96 ( .A1(a[15]), .A2(b[4]), .ZN(y[244]) );
  OR2_X1 U96bar ( .A1(abar[15]), .A2(bbar[4]), .ZN(ybar[244]);
  AND2_X1 U97 ( .A1(a[15]), .A2(b[3]), .ZN(y[243]) );
  OR2_X1 U97bar ( .A1(abar[15]), .A2(bbar[3]), .ZN(ybar[243]);
  AND2_X1 U98 ( .A1(a[15]), .A2(b[2]), .ZN(y[242]) );
  OR2_X1 U98bar ( .A1(abar[15]), .A2(bbar[2]), .ZN(ybar[242]);
  AND2_X1 U99 ( .A1(a[15]), .A2(b[1]), .ZN(y[241]) );
  OR2_X1 U99bar ( .A1(abar[15]), .A2(bbar[1]), .ZN(ybar[241]);
  AND2_X1 U100 ( .A1(a[15]), .A2(b[0]), .ZN(y[240]) );
  OR2_X1 U100bar ( .A1(abar[15]), .A2(bbar[0]), .ZN(ybar[240]);
  AND2_X1 U101 ( .A1(a[1]), .A2(b[7]), .ZN(y[23]) );
  OR2_X1 U101bar ( .A1(abar[1]), .A2(bbar[7]), .ZN(ybar[23]);
  AND2_X1 U102 ( .A1(a[14]), .A2(b[15]), .ZN(y[239]) );
  OR2_X1 U102bar ( .A1(abar[14]), .A2(bbar[15]), .ZN(ybar[239]);
  AND2_X1 U103 ( .A1(a[14]), .A2(b[14]), .ZN(y[238]) );
  OR2_X1 U103bar ( .A1(abar[14]), .A2(bbar[14]), .ZN(ybar[238]);
  AND2_X1 U104 ( .A1(a[14]), .A2(b[13]), .ZN(y[237]) );
  OR2_X1 U104bar ( .A1(abar[14]), .A2(bbar[13]), .ZN(ybar[237]);
  AND2_X1 U105 ( .A1(a[14]), .A2(b[12]), .ZN(y[236]) );
  OR2_X1 U105bar ( .A1(abar[14]), .A2(bbar[12]), .ZN(ybar[236]);
  AND2_X1 U106 ( .A1(a[14]), .A2(b[11]), .ZN(y[235]) );
  OR2_X1 U106bar ( .A1(abar[14]), .A2(bbar[11]), .ZN(ybar[235]);
  AND2_X1 U107 ( .A1(a[14]), .A2(b[10]), .ZN(y[234]) );
  OR2_X1 U107bar ( .A1(abar[14]), .A2(bbar[10]), .ZN(ybar[234]);
  AND2_X1 U108 ( .A1(a[14]), .A2(b[9]), .ZN(y[233]) );
  OR2_X1 U108bar ( .A1(abar[14]), .A2(bbar[9]), .ZN(ybar[233]);
  AND2_X1 U109 ( .A1(a[14]), .A2(b[8]), .ZN(y[232]) );
  OR2_X1 U109bar ( .A1(abar[14]), .A2(bbar[8]), .ZN(ybar[232]);
  AND2_X1 U110 ( .A1(a[14]), .A2(b[7]), .ZN(y[231]) );
  OR2_X1 U110bar ( .A1(abar[14]), .A2(bbar[7]), .ZN(ybar[231]);
  AND2_X1 U111 ( .A1(a[14]), .A2(b[6]), .ZN(y[230]) );
  OR2_X1 U111bar ( .A1(abar[14]), .A2(bbar[6]), .ZN(ybar[230]);
  AND2_X1 U112 ( .A1(a[1]), .A2(b[6]), .ZN(y[22]) );
  OR2_X1 U112bar ( .A1(abar[1]), .A2(bbar[6]), .ZN(ybar[22]);
  AND2_X1 U113 ( .A1(a[14]), .A2(b[5]), .ZN(y[229]) );
  OR2_X1 U113bar ( .A1(abar[14]), .A2(bbar[5]), .ZN(ybar[229]);
  AND2_X1 U114 ( .A1(a[14]), .A2(b[4]), .ZN(y[228]) );
  OR2_X1 U114bar ( .A1(abar[14]), .A2(bbar[4]), .ZN(ybar[228]);
  AND2_X1 U115 ( .A1(a[14]), .A2(b[3]), .ZN(y[227]) );
  OR2_X1 U115bar ( .A1(abar[14]), .A2(bbar[3]), .ZN(ybar[227]);
  AND2_X1 U116 ( .A1(a[14]), .A2(b[2]), .ZN(y[226]) );
  OR2_X1 U116bar ( .A1(abar[14]), .A2(bbar[2]), .ZN(ybar[226]);
  AND2_X1 U117 ( .A1(a[14]), .A2(b[1]), .ZN(y[225]) );
  OR2_X1 U117bar ( .A1(abar[14]), .A2(bbar[1]), .ZN(ybar[225]);
  AND2_X1 U118 ( .A1(a[14]), .A2(b[0]), .ZN(y[224]) );
  OR2_X1 U118bar ( .A1(abar[14]), .A2(bbar[0]), .ZN(ybar[224]);
  AND2_X1 U119 ( .A1(a[13]), .A2(b[15]), .ZN(y[223]) );
  OR2_X1 U119bar ( .A1(abar[13]), .A2(bbar[15]), .ZN(ybar[223]);
  AND2_X1 U120 ( .A1(a[13]), .A2(b[14]), .ZN(y[222]) );
  OR2_X1 U120bar ( .A1(abar[13]), .A2(bbar[14]), .ZN(ybar[222]);
  AND2_X1 U121 ( .A1(a[13]), .A2(b[13]), .ZN(y[221]) );
  OR2_X1 U121bar ( .A1(abar[13]), .A2(bbar[13]), .ZN(ybar[221]);
  AND2_X1 U122 ( .A1(a[13]), .A2(b[12]), .ZN(y[220]) );
  OR2_X1 U122bar ( .A1(abar[13]), .A2(bbar[12]), .ZN(ybar[220]);
  AND2_X1 U123 ( .A1(a[1]), .A2(b[5]), .ZN(y[21]) );
  OR2_X1 U123bar ( .A1(abar[1]), .A2(bbar[5]), .ZN(ybar[21]);
  AND2_X1 U124 ( .A1(a[13]), .A2(b[11]), .ZN(y[219]) );
  OR2_X1 U124bar ( .A1(abar[13]), .A2(bbar[11]), .ZN(ybar[219]);
  AND2_X1 U125 ( .A1(a[13]), .A2(b[10]), .ZN(y[218]) );
  OR2_X1 U125bar ( .A1(abar[13]), .A2(bbar[10]), .ZN(ybar[218]);
  AND2_X1 U126 ( .A1(a[13]), .A2(b[9]), .ZN(y[217]) );
  OR2_X1 U126bar ( .A1(abar[13]), .A2(bbar[9]), .ZN(ybar[217]);
  AND2_X1 U127 ( .A1(a[13]), .A2(b[8]), .ZN(y[216]) );
  OR2_X1 U127bar ( .A1(abar[13]), .A2(bbar[8]), .ZN(ybar[216]);
  AND2_X1 U128 ( .A1(a[13]), .A2(b[7]), .ZN(y[215]) );
  OR2_X1 U128bar ( .A1(abar[13]), .A2(bbar[7]), .ZN(ybar[215]);
  AND2_X1 U129 ( .A1(a[13]), .A2(b[6]), .ZN(y[214]) );
  OR2_X1 U129bar ( .A1(abar[13]), .A2(bbar[6]), .ZN(ybar[214]);
  AND2_X1 U130 ( .A1(a[13]), .A2(b[5]), .ZN(y[213]) );
  OR2_X1 U130bar ( .A1(abar[13]), .A2(bbar[5]), .ZN(ybar[213]);
  AND2_X1 U131 ( .A1(a[13]), .A2(b[4]), .ZN(y[212]) );
  OR2_X1 U131bar ( .A1(abar[13]), .A2(bbar[4]), .ZN(ybar[212]);
  AND2_X1 U132 ( .A1(a[13]), .A2(b[3]), .ZN(y[211]) );
  OR2_X1 U132bar ( .A1(abar[13]), .A2(bbar[3]), .ZN(ybar[211]);
  AND2_X1 U133 ( .A1(a[13]), .A2(b[2]), .ZN(y[210]) );
  OR2_X1 U133bar ( .A1(abar[13]), .A2(bbar[2]), .ZN(ybar[210]);
  AND2_X1 U134 ( .A1(a[1]), .A2(b[4]), .ZN(y[20]) );
  OR2_X1 U134bar ( .A1(abar[1]), .A2(bbar[4]), .ZN(ybar[20]);
  AND2_X1 U135 ( .A1(a[13]), .A2(b[1]), .ZN(y[209]) );
  OR2_X1 U135bar ( .A1(abar[13]), .A2(bbar[1]), .ZN(ybar[209]);
  AND2_X1 U136 ( .A1(a[13]), .A2(b[0]), .ZN(y[208]) );
  OR2_X1 U136bar ( .A1(abar[13]), .A2(bbar[0]), .ZN(ybar[208]);
  AND2_X1 U137 ( .A1(a[12]), .A2(b[15]), .ZN(y[207]) );
  OR2_X1 U137bar ( .A1(abar[12]), .A2(bbar[15]), .ZN(ybar[207]);
  AND2_X1 U138 ( .A1(a[12]), .A2(b[14]), .ZN(y[206]) );
  OR2_X1 U138bar ( .A1(abar[12]), .A2(bbar[14]), .ZN(ybar[206]);
  AND2_X1 U139 ( .A1(a[12]), .A2(b[13]), .ZN(y[205]) );
  OR2_X1 U139bar ( .A1(abar[12]), .A2(bbar[13]), .ZN(ybar[205]);
  AND2_X1 U140 ( .A1(a[12]), .A2(b[12]), .ZN(y[204]) );
  OR2_X1 U140bar ( .A1(abar[12]), .A2(bbar[12]), .ZN(ybar[204]);
  AND2_X1 U141 ( .A1(a[12]), .A2(b[11]), .ZN(y[203]) );
  OR2_X1 U141bar ( .A1(abar[12]), .A2(bbar[11]), .ZN(ybar[203]);
  AND2_X1 U142 ( .A1(a[12]), .A2(b[10]), .ZN(y[202]) );
  OR2_X1 U142bar ( .A1(abar[12]), .A2(bbar[10]), .ZN(ybar[202]);
  AND2_X1 U143 ( .A1(a[12]), .A2(b[9]), .ZN(y[201]) );
  OR2_X1 U143bar ( .A1(abar[12]), .A2(bbar[9]), .ZN(ybar[201]);
  AND2_X1 U144 ( .A1(a[12]), .A2(b[8]), .ZN(y[200]) );
  OR2_X1 U144bar ( .A1(abar[12]), .A2(bbar[8]), .ZN(ybar[200]);
  AND2_X1 U145 ( .A1(b[1]), .A2(a[0]), .ZN(y[1]) );
  OR2_X1 U145bar ( .A1(bbar[1]), .A2(abar[0]), .ZN(ybar[1]);
  AND2_X1 U146 ( .A1(a[1]), .A2(b[3]), .ZN(y[19]) );
  OR2_X1 U146bar ( .A1(abar[1]), .A2(bbar[3]), .ZN(ybar[19]);
  AND2_X1 U147 ( .A1(a[12]), .A2(b[7]), .ZN(y[199]) );
  OR2_X1 U147bar ( .A1(abar[12]), .A2(bbar[7]), .ZN(ybar[199]);
  AND2_X1 U148 ( .A1(a[12]), .A2(b[6]), .ZN(y[198]) );
  OR2_X1 U148bar ( .A1(abar[12]), .A2(bbar[6]), .ZN(ybar[198]);
  AND2_X1 U149 ( .A1(a[12]), .A2(b[5]), .ZN(y[197]) );
  OR2_X1 U149bar ( .A1(abar[12]), .A2(bbar[5]), .ZN(ybar[197]);
  AND2_X1 U150 ( .A1(a[12]), .A2(b[4]), .ZN(y[196]) );
  OR2_X1 U150bar ( .A1(abar[12]), .A2(bbar[4]), .ZN(ybar[196]);
  AND2_X1 U151 ( .A1(a[12]), .A2(b[3]), .ZN(y[195]) );
  OR2_X1 U151bar ( .A1(abar[12]), .A2(bbar[3]), .ZN(ybar[195]);
  AND2_X1 U152 ( .A1(a[12]), .A2(b[2]), .ZN(y[194]) );
  OR2_X1 U152bar ( .A1(abar[12]), .A2(bbar[2]), .ZN(ybar[194]);
  AND2_X1 U153 ( .A1(a[12]), .A2(b[1]), .ZN(y[193]) );
  OR2_X1 U153bar ( .A1(abar[12]), .A2(bbar[1]), .ZN(ybar[193]);
  AND2_X1 U154 ( .A1(a[12]), .A2(b[0]), .ZN(y[192]) );
  OR2_X1 U154bar ( .A1(abar[12]), .A2(bbar[0]), .ZN(ybar[192]);
  AND2_X1 U155 ( .A1(a[11]), .A2(b[15]), .ZN(y[191]) );
  OR2_X1 U155bar ( .A1(abar[11]), .A2(bbar[15]), .ZN(ybar[191]);
  AND2_X1 U156 ( .A1(a[11]), .A2(b[14]), .ZN(y[190]) );
  OR2_X1 U156bar ( .A1(abar[11]), .A2(bbar[14]), .ZN(ybar[190]);
  AND2_X1 U157 ( .A1(a[1]), .A2(b[2]), .ZN(y[18]) );
  OR2_X1 U157bar ( .A1(abar[1]), .A2(bbar[2]), .ZN(ybar[18]);
  AND2_X1 U158 ( .A1(a[11]), .A2(b[13]), .ZN(y[189]) );
  OR2_X1 U158bar ( .A1(abar[11]), .A2(bbar[13]), .ZN(ybar[189]);
  AND2_X1 U159 ( .A1(a[11]), .A2(b[12]), .ZN(y[188]) );
  OR2_X1 U159bar ( .A1(abar[11]), .A2(bbar[12]), .ZN(ybar[188]);
  AND2_X1 U160 ( .A1(a[11]), .A2(b[11]), .ZN(y[187]) );
  OR2_X1 U160bar ( .A1(abar[11]), .A2(bbar[11]), .ZN(ybar[187]);
  AND2_X1 U161 ( .A1(a[11]), .A2(b[10]), .ZN(y[186]) );
  OR2_X1 U161bar ( .A1(abar[11]), .A2(bbar[10]), .ZN(ybar[186]);
  AND2_X1 U162 ( .A1(a[11]), .A2(b[9]), .ZN(y[185]) );
  OR2_X1 U162bar ( .A1(abar[11]), .A2(bbar[9]), .ZN(ybar[185]);
  AND2_X1 U163 ( .A1(a[11]), .A2(b[8]), .ZN(y[184]) );
  OR2_X1 U163bar ( .A1(abar[11]), .A2(bbar[8]), .ZN(ybar[184]);
  AND2_X1 U164 ( .A1(a[11]), .A2(b[7]), .ZN(y[183]) );
  OR2_X1 U164bar ( .A1(abar[11]), .A2(bbar[7]), .ZN(ybar[183]);
  AND2_X1 U165 ( .A1(a[11]), .A2(b[6]), .ZN(y[182]) );
  OR2_X1 U165bar ( .A1(abar[11]), .A2(bbar[6]), .ZN(ybar[182]);
  AND2_X1 U166 ( .A1(a[11]), .A2(b[5]), .ZN(y[181]) );
  OR2_X1 U166bar ( .A1(abar[11]), .A2(bbar[5]), .ZN(ybar[181]);
  AND2_X1 U167 ( .A1(a[11]), .A2(b[4]), .ZN(y[180]) );
  OR2_X1 U167bar ( .A1(abar[11]), .A2(bbar[4]), .ZN(ybar[180]);
  AND2_X1 U168 ( .A1(a[1]), .A2(b[1]), .ZN(y[17]) );
  OR2_X1 U168bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[17]);
  AND2_X1 U169 ( .A1(a[11]), .A2(b[3]), .ZN(y[179]) );
  OR2_X1 U169bar ( .A1(abar[11]), .A2(bbar[3]), .ZN(ybar[179]);
  AND2_X1 U170 ( .A1(a[11]), .A2(b[2]), .ZN(y[178]) );
  OR2_X1 U170bar ( .A1(abar[11]), .A2(bbar[2]), .ZN(ybar[178]);
  AND2_X1 U171 ( .A1(a[11]), .A2(b[1]), .ZN(y[177]) );
  OR2_X1 U171bar ( .A1(abar[11]), .A2(bbar[1]), .ZN(ybar[177]);
  AND2_X1 U172 ( .A1(a[11]), .A2(b[0]), .ZN(y[176]) );
  OR2_X1 U172bar ( .A1(abar[11]), .A2(bbar[0]), .ZN(ybar[176]);
  AND2_X1 U173 ( .A1(a[10]), .A2(b[15]), .ZN(y[175]) );
  OR2_X1 U173bar ( .A1(abar[10]), .A2(bbar[15]), .ZN(ybar[175]);
  AND2_X1 U174 ( .A1(a[10]), .A2(b[14]), .ZN(y[174]) );
  OR2_X1 U174bar ( .A1(abar[10]), .A2(bbar[14]), .ZN(ybar[174]);
  AND2_X1 U175 ( .A1(a[10]), .A2(b[13]), .ZN(y[173]) );
  OR2_X1 U175bar ( .A1(abar[10]), .A2(bbar[13]), .ZN(ybar[173]);
  AND2_X1 U176 ( .A1(a[10]), .A2(b[12]), .ZN(y[172]) );
  OR2_X1 U176bar ( .A1(abar[10]), .A2(bbar[12]), .ZN(ybar[172]);
  AND2_X1 U177 ( .A1(a[10]), .A2(b[11]), .ZN(y[171]) );
  OR2_X1 U177bar ( .A1(abar[10]), .A2(bbar[11]), .ZN(ybar[171]);
  AND2_X1 U178 ( .A1(a[10]), .A2(b[10]), .ZN(y[170]) );
  OR2_X1 U178bar ( .A1(abar[10]), .A2(bbar[10]), .ZN(ybar[170]);
  AND2_X1 U179 ( .A1(a[1]), .A2(b[0]), .ZN(y[16]) );
  OR2_X1 U179bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[16]);
  AND2_X1 U180 ( .A1(a[10]), .A2(b[9]), .ZN(y[169]) );
  OR2_X1 U180bar ( .A1(abar[10]), .A2(bbar[9]), .ZN(ybar[169]);
  AND2_X1 U181 ( .A1(a[10]), .A2(b[8]), .ZN(y[168]) );
  OR2_X1 U181bar ( .A1(abar[10]), .A2(bbar[8]), .ZN(ybar[168]);
  AND2_X1 U182 ( .A1(a[10]), .A2(b[7]), .ZN(y[167]) );
  OR2_X1 U182bar ( .A1(abar[10]), .A2(bbar[7]), .ZN(ybar[167]);
  AND2_X1 U183 ( .A1(a[10]), .A2(b[6]), .ZN(y[166]) );
  OR2_X1 U183bar ( .A1(abar[10]), .A2(bbar[6]), .ZN(ybar[166]);
  AND2_X1 U184 ( .A1(a[10]), .A2(b[5]), .ZN(y[165]) );
  OR2_X1 U184bar ( .A1(abar[10]), .A2(bbar[5]), .ZN(ybar[165]);
  AND2_X1 U185 ( .A1(a[10]), .A2(b[4]), .ZN(y[164]) );
  OR2_X1 U185bar ( .A1(abar[10]), .A2(bbar[4]), .ZN(ybar[164]);
  AND2_X1 U186 ( .A1(a[10]), .A2(b[3]), .ZN(y[163]) );
  OR2_X1 U186bar ( .A1(abar[10]), .A2(bbar[3]), .ZN(ybar[163]);
  AND2_X1 U187 ( .A1(a[10]), .A2(b[2]), .ZN(y[162]) );
  OR2_X1 U187bar ( .A1(abar[10]), .A2(bbar[2]), .ZN(ybar[162]);
  AND2_X1 U188 ( .A1(a[10]), .A2(b[1]), .ZN(y[161]) );
  OR2_X1 U188bar ( .A1(abar[10]), .A2(bbar[1]), .ZN(ybar[161]);
  AND2_X1 U189 ( .A1(a[10]), .A2(b[0]), .ZN(y[160]) );
  OR2_X1 U189bar ( .A1(abar[10]), .A2(bbar[0]), .ZN(ybar[160]);
  AND2_X1 U190 ( .A1(b[15]), .A2(a[0]), .ZN(y[15]) );
  OR2_X1 U190bar ( .A1(bbar[15]), .A2(abar[0]), .ZN(ybar[15]);
  AND2_X1 U191 ( .A1(a[9]), .A2(b[15]), .ZN(y[159]) );
  OR2_X1 U191bar ( .A1(abar[9]), .A2(bbar[15]), .ZN(ybar[159]);
  AND2_X1 U192 ( .A1(a[9]), .A2(b[14]), .ZN(y[158]) );
  OR2_X1 U192bar ( .A1(abar[9]), .A2(bbar[14]), .ZN(ybar[158]);
  AND2_X1 U193 ( .A1(a[9]), .A2(b[13]), .ZN(y[157]) );
  OR2_X1 U193bar ( .A1(abar[9]), .A2(bbar[13]), .ZN(ybar[157]);
  AND2_X1 U194 ( .A1(a[9]), .A2(b[12]), .ZN(y[156]) );
  OR2_X1 U194bar ( .A1(abar[9]), .A2(bbar[12]), .ZN(ybar[156]);
  AND2_X1 U195 ( .A1(a[9]), .A2(b[11]), .ZN(y[155]) );
  OR2_X1 U195bar ( .A1(abar[9]), .A2(bbar[11]), .ZN(ybar[155]);
  AND2_X1 U196 ( .A1(a[9]), .A2(b[10]), .ZN(y[154]) );
  OR2_X1 U196bar ( .A1(abar[9]), .A2(bbar[10]), .ZN(ybar[154]);
  AND2_X1 U197 ( .A1(a[9]), .A2(b[9]), .ZN(y[153]) );
  OR2_X1 U197bar ( .A1(abar[9]), .A2(bbar[9]), .ZN(ybar[153]);
  AND2_X1 U198 ( .A1(a[9]), .A2(b[8]), .ZN(y[152]) );
  OR2_X1 U198bar ( .A1(abar[9]), .A2(bbar[8]), .ZN(ybar[152]);
  AND2_X1 U199 ( .A1(a[9]), .A2(b[7]), .ZN(y[151]) );
  OR2_X1 U199bar ( .A1(abar[9]), .A2(bbar[7]), .ZN(ybar[151]);
  AND2_X1 U200 ( .A1(a[9]), .A2(b[6]), .ZN(y[150]) );
  OR2_X1 U200bar ( .A1(abar[9]), .A2(bbar[6]), .ZN(ybar[150]);
  AND2_X1 U201 ( .A1(b[14]), .A2(a[0]), .ZN(y[14]) );
  OR2_X1 U201bar ( .A1(bbar[14]), .A2(abar[0]), .ZN(ybar[14]);
  AND2_X1 U202 ( .A1(a[9]), .A2(b[5]), .ZN(y[149]) );
  OR2_X1 U202bar ( .A1(abar[9]), .A2(bbar[5]), .ZN(ybar[149]);
  AND2_X1 U203 ( .A1(a[9]), .A2(b[4]), .ZN(y[148]) );
  OR2_X1 U203bar ( .A1(abar[9]), .A2(bbar[4]), .ZN(ybar[148]);
  AND2_X1 U204 ( .A1(a[9]), .A2(b[3]), .ZN(y[147]) );
  OR2_X1 U204bar ( .A1(abar[9]), .A2(bbar[3]), .ZN(ybar[147]);
  AND2_X1 U205 ( .A1(a[9]), .A2(b[2]), .ZN(y[146]) );
  OR2_X1 U205bar ( .A1(abar[9]), .A2(bbar[2]), .ZN(ybar[146]);
  AND2_X1 U206 ( .A1(a[9]), .A2(b[1]), .ZN(y[145]) );
  OR2_X1 U206bar ( .A1(abar[9]), .A2(bbar[1]), .ZN(ybar[145]);
  AND2_X1 U207 ( .A1(a[9]), .A2(b[0]), .ZN(y[144]) );
  OR2_X1 U207bar ( .A1(abar[9]), .A2(bbar[0]), .ZN(ybar[144]);
  AND2_X1 U208 ( .A1(a[8]), .A2(b[15]), .ZN(y[143]) );
  OR2_X1 U208bar ( .A1(abar[8]), .A2(bbar[15]), .ZN(ybar[143]);
  AND2_X1 U209 ( .A1(a[8]), .A2(b[14]), .ZN(y[142]) );
  OR2_X1 U209bar ( .A1(abar[8]), .A2(bbar[14]), .ZN(ybar[142]);
  AND2_X1 U210 ( .A1(a[8]), .A2(b[13]), .ZN(y[141]) );
  OR2_X1 U210bar ( .A1(abar[8]), .A2(bbar[13]), .ZN(ybar[141]);
  AND2_X1 U211 ( .A1(a[8]), .A2(b[12]), .ZN(y[140]) );
  OR2_X1 U211bar ( .A1(abar[8]), .A2(bbar[12]), .ZN(ybar[140]);
  AND2_X1 U212 ( .A1(b[13]), .A2(a[0]), .ZN(y[13]) );
  OR2_X1 U212bar ( .A1(bbar[13]), .A2(abar[0]), .ZN(ybar[13]);
  AND2_X1 U213 ( .A1(a[8]), .A2(b[11]), .ZN(y[139]) );
  OR2_X1 U213bar ( .A1(abar[8]), .A2(bbar[11]), .ZN(ybar[139]);
  AND2_X1 U214 ( .A1(a[8]), .A2(b[10]), .ZN(y[138]) );
  OR2_X1 U214bar ( .A1(abar[8]), .A2(bbar[10]), .ZN(ybar[138]);
  AND2_X1 U215 ( .A1(a[8]), .A2(b[9]), .ZN(y[137]) );
  OR2_X1 U215bar ( .A1(abar[8]), .A2(bbar[9]), .ZN(ybar[137]);
  AND2_X1 U216 ( .A1(a[8]), .A2(b[8]), .ZN(y[136]) );
  OR2_X1 U216bar ( .A1(abar[8]), .A2(bbar[8]), .ZN(ybar[136]);
  AND2_X1 U217 ( .A1(a[8]), .A2(b[7]), .ZN(y[135]) );
  OR2_X1 U217bar ( .A1(abar[8]), .A2(bbar[7]), .ZN(ybar[135]);
  AND2_X1 U218 ( .A1(a[8]), .A2(b[6]), .ZN(y[134]) );
  OR2_X1 U218bar ( .A1(abar[8]), .A2(bbar[6]), .ZN(ybar[134]);
  AND2_X1 U219 ( .A1(a[8]), .A2(b[5]), .ZN(y[133]) );
  OR2_X1 U219bar ( .A1(abar[8]), .A2(bbar[5]), .ZN(ybar[133]);
  AND2_X1 U220 ( .A1(a[8]), .A2(b[4]), .ZN(y[132]) );
  OR2_X1 U220bar ( .A1(abar[8]), .A2(bbar[4]), .ZN(ybar[132]);
  AND2_X1 U221 ( .A1(a[8]), .A2(b[3]), .ZN(y[131]) );
  OR2_X1 U221bar ( .A1(abar[8]), .A2(bbar[3]), .ZN(ybar[131]);
  AND2_X1 U222 ( .A1(a[8]), .A2(b[2]), .ZN(y[130]) );
  OR2_X1 U222bar ( .A1(abar[8]), .A2(bbar[2]), .ZN(ybar[130]);
  AND2_X1 U223 ( .A1(b[12]), .A2(a[0]), .ZN(y[12]) );
  OR2_X1 U223bar ( .A1(bbar[12]), .A2(abar[0]), .ZN(ybar[12]);
  AND2_X1 U224 ( .A1(a[8]), .A2(b[1]), .ZN(y[129]) );
  OR2_X1 U224bar ( .A1(abar[8]), .A2(bbar[1]), .ZN(ybar[129]);
  AND2_X1 U225 ( .A1(a[8]), .A2(b[0]), .ZN(y[128]) );
  OR2_X1 U225bar ( .A1(abar[8]), .A2(bbar[0]), .ZN(ybar[128]);
  AND2_X1 U226 ( .A1(a[7]), .A2(b[15]), .ZN(y[127]) );
  OR2_X1 U226bar ( .A1(abar[7]), .A2(bbar[15]), .ZN(ybar[127]);
  AND2_X1 U227 ( .A1(a[7]), .A2(b[14]), .ZN(y[126]) );
  OR2_X1 U227bar ( .A1(abar[7]), .A2(bbar[14]), .ZN(ybar[126]);
  AND2_X1 U228 ( .A1(a[7]), .A2(b[13]), .ZN(y[125]) );
  OR2_X1 U228bar ( .A1(abar[7]), .A2(bbar[13]), .ZN(ybar[125]);
  AND2_X1 U229 ( .A1(a[7]), .A2(b[12]), .ZN(y[124]) );
  OR2_X1 U229bar ( .A1(abar[7]), .A2(bbar[12]), .ZN(ybar[124]);
  AND2_X1 U230 ( .A1(a[7]), .A2(b[11]), .ZN(y[123]) );
  OR2_X1 U230bar ( .A1(abar[7]), .A2(bbar[11]), .ZN(ybar[123]);
  AND2_X1 U231 ( .A1(a[7]), .A2(b[10]), .ZN(y[122]) );
  OR2_X1 U231bar ( .A1(abar[7]), .A2(bbar[10]), .ZN(ybar[122]);
  AND2_X1 U232 ( .A1(a[7]), .A2(b[9]), .ZN(y[121]) );
  OR2_X1 U232bar ( .A1(abar[7]), .A2(bbar[9]), .ZN(ybar[121]);
  AND2_X1 U233 ( .A1(a[7]), .A2(b[8]), .ZN(y[120]) );
  OR2_X1 U233bar ( .A1(abar[7]), .A2(bbar[8]), .ZN(ybar[120]);
  AND2_X1 U234 ( .A1(b[11]), .A2(a[0]), .ZN(y[11]) );
  OR2_X1 U234bar ( .A1(bbar[11]), .A2(abar[0]), .ZN(ybar[11]);
  AND2_X1 U235 ( .A1(a[7]), .A2(b[7]), .ZN(y[119]) );
  OR2_X1 U235bar ( .A1(abar[7]), .A2(bbar[7]), .ZN(ybar[119]);
  AND2_X1 U236 ( .A1(a[7]), .A2(b[6]), .ZN(y[118]) );
  OR2_X1 U236bar ( .A1(abar[7]), .A2(bbar[6]), .ZN(ybar[118]);
  AND2_X1 U237 ( .A1(a[7]), .A2(b[5]), .ZN(y[117]) );
  OR2_X1 U237bar ( .A1(abar[7]), .A2(bbar[5]), .ZN(ybar[117]);
  AND2_X1 U238 ( .A1(a[7]), .A2(b[4]), .ZN(y[116]) );
  OR2_X1 U238bar ( .A1(abar[7]), .A2(bbar[4]), .ZN(ybar[116]);
  AND2_X1 U239 ( .A1(a[7]), .A2(b[3]), .ZN(y[115]) );
  OR2_X1 U239bar ( .A1(abar[7]), .A2(bbar[3]), .ZN(ybar[115]);
  AND2_X1 U240 ( .A1(a[7]), .A2(b[2]), .ZN(y[114]) );
  OR2_X1 U240bar ( .A1(abar[7]), .A2(bbar[2]), .ZN(ybar[114]);
  AND2_X1 U241 ( .A1(a[7]), .A2(b[1]), .ZN(y[113]) );
  OR2_X1 U241bar ( .A1(abar[7]), .A2(bbar[1]), .ZN(ybar[113]);
  AND2_X1 U242 ( .A1(a[7]), .A2(b[0]), .ZN(y[112]) );
  OR2_X1 U242bar ( .A1(abar[7]), .A2(bbar[0]), .ZN(ybar[112]);
  AND2_X1 U243 ( .A1(b[15]), .A2(a[6]), .ZN(y[111]) );
  OR2_X1 U243bar ( .A1(bbar[15]), .A2(abar[6]), .ZN(ybar[111]);
  AND2_X1 U244 ( .A1(b[14]), .A2(a[6]), .ZN(y[110]) );
  OR2_X1 U244bar ( .A1(bbar[14]), .A2(abar[6]), .ZN(ybar[110]);
  AND2_X1 U245 ( .A1(b[10]), .A2(a[0]), .ZN(y[10]) );
  OR2_X1 U245bar ( .A1(bbar[10]), .A2(abar[0]), .ZN(ybar[10]);
  AND2_X1 U246 ( .A1(b[13]), .A2(a[6]), .ZN(y[109]) );
  OR2_X1 U246bar ( .A1(bbar[13]), .A2(abar[6]), .ZN(ybar[109]);
  AND2_X1 U247 ( .A1(b[12]), .A2(a[6]), .ZN(y[108]) );
  OR2_X1 U247bar ( .A1(bbar[12]), .A2(abar[6]), .ZN(ybar[108]);
  AND2_X1 U248 ( .A1(b[11]), .A2(a[6]), .ZN(y[107]) );
  OR2_X1 U248bar ( .A1(bbar[11]), .A2(abar[6]), .ZN(ybar[107]);
  AND2_X1 U249 ( .A1(b[10]), .A2(a[6]), .ZN(y[106]) );
  OR2_X1 U249bar ( .A1(bbar[10]), .A2(abar[6]), .ZN(ybar[106]);
  AND2_X1 U250 ( .A1(a[6]), .A2(b[9]), .ZN(y[105]) );
  OR2_X1 U250bar ( .A1(abar[6]), .A2(bbar[9]), .ZN(ybar[105]);
  AND2_X1 U251 ( .A1(b[8]), .A2(a[6]), .ZN(y[104]) );
  OR2_X1 U251bar ( .A1(bbar[8]), .A2(abar[6]), .ZN(ybar[104]);
  AND2_X1 U252 ( .A1(b[7]), .A2(a[6]), .ZN(y[103]) );
  OR2_X1 U252bar ( .A1(bbar[7]), .A2(abar[6]), .ZN(ybar[103]);
  AND2_X1 U253 ( .A1(b[6]), .A2(a[6]), .ZN(y[102]) );
  OR2_X1 U253bar ( .A1(bbar[6]), .A2(abar[6]), .ZN(ybar[102]);
  AND2_X1 U254 ( .A1(b[5]), .A2(a[6]), .ZN(y[101]) );
  OR2_X1 U254bar ( .A1(bbar[5]), .A2(abar[6]), .ZN(ybar[101]);
  AND2_X1 U255 ( .A1(b[4]), .A2(a[6]), .ZN(y[100]) );
  OR2_X1 U255bar ( .A1(bbar[4]), .A2(abar[6]), .ZN(ybar[100]);
  AND2_X1 U256 ( .A1(b[0]), .A2(a[0]), .ZN(y[0]) );
  OR2_X1 U256bar ( .A1(bbar[0]), .A2(abar[0]), .ZN(ybar[0]);
endmodule




module decode_7 ( in, out );
  input [7:0] in;
  //input_done

  output [255:0] out;
  //output_done

  wire   [15:0] level1;
  wire   [31:0] level2;
  //wire_done

  CD2_28 cd_l1_1 ( .a(in[1]), .b(in[0]), .y(level1[3:0]) );
  CD2_27 cd_l1_2 ( .a(in[3]), .b(in[2]), .y(level1[7:4]) );
  CD2_26 cd_l1_3 ( .a(in[5]), .b(in[4]), .y(level1[11:8]) );
  CD2_25 cd_l1_4 ( .a(in[7]), .b(in[6]), .y(level1[15:12]) );
  CD4_14 cd_l2_1 ( .a(level1[7:4]), .b(level1[3:0]), .y(level2[15:0]) );
  CD4_13 cd_l2_2 ( .a(level1[15:12]), .b(level1[11:8]), .y(level2[31:16]) );
  CD16_7 cd_l3 ( .a(level2[31:16]), .b(level2[15:0]), .y(out) );
endmodule


module encode_7 ( in, out );
  input [255:0] in;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
  assign inbar[8] = ~in[8];
  assign inbar[9] = ~in[9];
  assign inbar[10] = ~in[10];
  assign inbar[11] = ~in[11];
  assign inbar[12] = ~in[12];
  assign inbar[13] = ~in[13];
  assign inbar[14] = ~in[14];
  assign inbar[15] = ~in[15];
  assign inbar[16] = ~in[16];
  assign inbar[17] = ~in[17];
  assign inbar[18] = ~in[18];
  assign inbar[19] = ~in[19];
  assign inbar[20] = ~in[20];
  assign inbar[21] = ~in[21];
  assign inbar[22] = ~in[22];
  assign inbar[23] = ~in[23];
  assign inbar[24] = ~in[24];
  assign inbar[25] = ~in[25];
  assign inbar[26] = ~in[26];
  assign inbar[27] = ~in[27];
  assign inbar[28] = ~in[28];
  assign inbar[29] = ~in[29];
  assign inbar[30] = ~in[30];
  assign inbar[31] = ~in[31];
  assign inbar[32] = ~in[32];
  assign inbar[33] = ~in[33];
  assign inbar[34] = ~in[34];
  assign inbar[35] = ~in[35];
  assign inbar[36] = ~in[36];
  assign inbar[37] = ~in[37];
  assign inbar[38] = ~in[38];
  assign inbar[39] = ~in[39];
  assign inbar[40] = ~in[40];
  assign inbar[41] = ~in[41];
  assign inbar[42] = ~in[42];
  assign inbar[43] = ~in[43];
  assign inbar[44] = ~in[44];
  assign inbar[45] = ~in[45];
  assign inbar[46] = ~in[46];
  assign inbar[47] = ~in[47];
  assign inbar[48] = ~in[48];
  assign inbar[49] = ~in[49];
  assign inbar[50] = ~in[50];
  assign inbar[51] = ~in[51];
  assign inbar[52] = ~in[52];
  assign inbar[53] = ~in[53];
  assign inbar[54] = ~in[54];
  assign inbar[55] = ~in[55];
  assign inbar[56] = ~in[56];
  assign inbar[57] = ~in[57];
  assign inbar[58] = ~in[58];
  assign inbar[59] = ~in[59];
  assign inbar[60] = ~in[60];
  assign inbar[61] = ~in[61];
  assign inbar[62] = ~in[62];
  assign inbar[63] = ~in[63];
  assign inbar[64] = ~in[64];
  assign inbar[65] = ~in[65];
  assign inbar[66] = ~in[66];
  assign inbar[67] = ~in[67];
  assign inbar[68] = ~in[68];
  assign inbar[69] = ~in[69];
  assign inbar[70] = ~in[70];
  assign inbar[71] = ~in[71];
  assign inbar[72] = ~in[72];
  assign inbar[73] = ~in[73];
  assign inbar[74] = ~in[74];
  assign inbar[75] = ~in[75];
  assign inbar[76] = ~in[76];
  assign inbar[77] = ~in[77];
  assign inbar[78] = ~in[78];
  assign inbar[79] = ~in[79];
  assign inbar[80] = ~in[80];
  assign inbar[81] = ~in[81];
  assign inbar[82] = ~in[82];
  assign inbar[83] = ~in[83];
  assign inbar[84] = ~in[84];
  assign inbar[85] = ~in[85];
  assign inbar[86] = ~in[86];
  assign inbar[87] = ~in[87];
  assign inbar[88] = ~in[88];
  assign inbar[89] = ~in[89];
  assign inbar[90] = ~in[90];
  assign inbar[91] = ~in[91];
  assign inbar[92] = ~in[92];
  assign inbar[93] = ~in[93];
  assign inbar[94] = ~in[94];
  assign inbar[95] = ~in[95];
  assign inbar[96] = ~in[96];
  assign inbar[97] = ~in[97];
  assign inbar[98] = ~in[98];
  assign inbar[99] = ~in[99];
  assign inbar[100] = ~in[100];
  assign inbar[101] = ~in[101];
  assign inbar[102] = ~in[102];
  assign inbar[103] = ~in[103];
  assign inbar[104] = ~in[104];
  assign inbar[105] = ~in[105];
  assign inbar[106] = ~in[106];
  assign inbar[107] = ~in[107];
  assign inbar[108] = ~in[108];
  assign inbar[109] = ~in[109];
  assign inbar[110] = ~in[110];
  assign inbar[111] = ~in[111];
  assign inbar[112] = ~in[112];
  assign inbar[113] = ~in[113];
  assign inbar[114] = ~in[114];
  assign inbar[115] = ~in[115];
  assign inbar[116] = ~in[116];
  assign inbar[117] = ~in[117];
  assign inbar[118] = ~in[118];
  assign inbar[119] = ~in[119];
  assign inbar[120] = ~in[120];
  assign inbar[121] = ~in[121];
  assign inbar[122] = ~in[122];
  assign inbar[123] = ~in[123];
  assign inbar[124] = ~in[124];
  assign inbar[125] = ~in[125];
  assign inbar[126] = ~in[126];
  assign inbar[127] = ~in[127];
  assign inbar[128] = ~in[128];
  assign inbar[129] = ~in[129];
  assign inbar[130] = ~in[130];
  assign inbar[131] = ~in[131];
  assign inbar[132] = ~in[132];
  assign inbar[133] = ~in[133];
  assign inbar[134] = ~in[134];
  assign inbar[135] = ~in[135];
  assign inbar[136] = ~in[136];
  assign inbar[137] = ~in[137];
  assign inbar[138] = ~in[138];
  assign inbar[139] = ~in[139];
  assign inbar[140] = ~in[140];
  assign inbar[141] = ~in[141];
  assign inbar[142] = ~in[142];
  assign inbar[143] = ~in[143];
  assign inbar[144] = ~in[144];
  assign inbar[145] = ~in[145];
  assign inbar[146] = ~in[146];
  assign inbar[147] = ~in[147];
  assign inbar[148] = ~in[148];
  assign inbar[149] = ~in[149];
  assign inbar[150] = ~in[150];
  assign inbar[151] = ~in[151];
  assign inbar[152] = ~in[152];
  assign inbar[153] = ~in[153];
  assign inbar[154] = ~in[154];
  assign inbar[155] = ~in[155];
  assign inbar[156] = ~in[156];
  assign inbar[157] = ~in[157];
  assign inbar[158] = ~in[158];
  assign inbar[159] = ~in[159];
  assign inbar[160] = ~in[160];
  assign inbar[161] = ~in[161];
  assign inbar[162] = ~in[162];
  assign inbar[163] = ~in[163];
  assign inbar[164] = ~in[164];
  assign inbar[165] = ~in[165];
  assign inbar[166] = ~in[166];
  assign inbar[167] = ~in[167];
  assign inbar[168] = ~in[168];
  assign inbar[169] = ~in[169];
  assign inbar[170] = ~in[170];
  assign inbar[171] = ~in[171];
  assign inbar[172] = ~in[172];
  assign inbar[173] = ~in[173];
  assign inbar[174] = ~in[174];
  assign inbar[175] = ~in[175];
  assign inbar[176] = ~in[176];
  assign inbar[177] = ~in[177];
  assign inbar[178] = ~in[178];
  assign inbar[179] = ~in[179];
  assign inbar[180] = ~in[180];
  assign inbar[181] = ~in[181];
  assign inbar[182] = ~in[182];
  assign inbar[183] = ~in[183];
  assign inbar[184] = ~in[184];
  assign inbar[185] = ~in[185];
  assign inbar[186] = ~in[186];
  assign inbar[187] = ~in[187];
  assign inbar[188] = ~in[188];
  assign inbar[189] = ~in[189];
  assign inbar[190] = ~in[190];
  assign inbar[191] = ~in[191];
  assign inbar[192] = ~in[192];
  assign inbar[193] = ~in[193];
  assign inbar[194] = ~in[194];
  assign inbar[195] = ~in[195];
  assign inbar[196] = ~in[196];
  assign inbar[197] = ~in[197];
  assign inbar[198] = ~in[198];
  assign inbar[199] = ~in[199];
  assign inbar[200] = ~in[200];
  assign inbar[201] = ~in[201];
  assign inbar[202] = ~in[202];
  assign inbar[203] = ~in[203];
  assign inbar[204] = ~in[204];
  assign inbar[205] = ~in[205];
  assign inbar[206] = ~in[206];
  assign inbar[207] = ~in[207];
  assign inbar[208] = ~in[208];
  assign inbar[209] = ~in[209];
  assign inbar[210] = ~in[210];
  assign inbar[211] = ~in[211];
  assign inbar[212] = ~in[212];
  assign inbar[213] = ~in[213];
  assign inbar[214] = ~in[214];
  assign inbar[215] = ~in[215];
  assign inbar[216] = ~in[216];
  assign inbar[217] = ~in[217];
  assign inbar[218] = ~in[218];
  assign inbar[219] = ~in[219];
  assign inbar[220] = ~in[220];
  assign inbar[221] = ~in[221];
  assign inbar[222] = ~in[222];
  assign inbar[223] = ~in[223];
  assign inbar[224] = ~in[224];
  assign inbar[225] = ~in[225];
  assign inbar[226] = ~in[226];
  assign inbar[227] = ~in[227];
  assign inbar[228] = ~in[228];
  assign inbar[229] = ~in[229];
  assign inbar[230] = ~in[230];
  assign inbar[231] = ~in[231];
  assign inbar[232] = ~in[232];
  assign inbar[233] = ~in[233];
  assign inbar[234] = ~in[234];
  assign inbar[235] = ~in[235];
  assign inbar[236] = ~in[236];
  assign inbar[237] = ~in[237];
  assign inbar[238] = ~in[238];
  assign inbar[239] = ~in[239];
  assign inbar[240] = ~in[240];
  assign inbar[241] = ~in[241];
  assign inbar[242] = ~in[242];
  assign inbar[243] = ~in[243];
  assign inbar[244] = ~in[244];
  assign inbar[245] = ~in[245];
  assign inbar[246] = ~in[246];
  assign inbar[247] = ~in[247];
  assign inbar[248] = ~in[248];
  assign inbar[249] = ~in[249];
  assign inbar[250] = ~in[250];
  assign inbar[251] = ~in[251];
  assign inbar[252] = ~in[252];
  assign inbar[253] = ~in[253];
  assign inbar[254] = ~in[254];
  assign inbar[255] = ~in[255];
  //input_done

  output [7:0] out;
  reg [7:0] outbar;
  //output_done

  wire   in_81, in_80, in_79, in_78, in_77, in_76, in_75, in_74, in_73, in_72,
         in_71, in_70, in_69, in_68, in_67, in_66, in_65, in_64, in_63, in_62,
         in_61, in_60, in_59, in_58, in_57, in_56, in_55, in_54, in_53, in_52,
         in_51, in_50, in_49, in_48, in_47, in_46, in_45, in_44, in_43, in_42,
         in_41, in_40, in_39, in_38, in_37, in_36, in_35, in_34, in_33, in_32,
         in_31, in_30, in_29, in_28, in_27, in_26, in_25, in_24, in_23, in_22,
         in_21, in_20, in_19, in_18, in_17, in_16, in_15, in_14, in_13, in_12,
         in_11, in_10, in_9, in_8, in_7, in_6, in_5, in_4, in_3, in_2, in_1,
         in_0, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972;
  wire in_81bar, in_80bar, in_79bar, in_78bar, in_77bar, in_76bar, in_75bar, in_74bar, in_73bar, in_72bar, in_71bar, in_70bar, in_69bar, in_68bar, in_67bar, in_66bar, in_65bar, in_64bar, in_63bar, in_62bar, in_61bar, in_60bar, in_59bar, in_58bar, in_57bar, in_56bar, in_55bar, in_54bar, in_53bar, in_52bar, in_51bar, in_50bar, in_49bar, in_48bar, in_47bar, in_46bar, in_45bar, in_44bar, in_43bar, in_42bar, in_41bar, in_40bar, in_39bar, in_38bar, in_37bar, in_36bar, in_35bar, in_34bar, in_33bar, in_32bar, in_31bar, in_30bar, in_29bar, in_28bar, in_27bar, in_26bar, in_25bar, in_24bar, in_23bar, in_22bar, in_21bar, in_20bar, in_19bar, in_18bar, in_17bar, in_16bar, in_15bar, in_14bar, in_13bar, in_12bar, in_11bar, in_10bar, in_9bar, in_8bar, in_7bar, in_6bar, in_5bar, in_4bar, in_3bar, in_2bar, in_1bar, in_0bar, n487bar, n488bar, n489bar, n490bar, n491bar, n492bar, n493bar, n494bar, n495bar, n496bar, n497bar, n498bar, n499bar, n500bar, n501bar, n502bar, n503bar, n504bar, n505bar, n506bar, n507bar, n508bar, n509bar, n510bar, n511bar, n512bar, n513bar, n514bar, n515bar, n516bar, n517bar, n518bar, n519bar, n520bar, n521bar, n522bar, n523bar, n524bar, n525bar, n526bar, n527bar, n528bar, n529bar, n530bar, n531bar, n532bar, n533bar, n534bar, n535bar, n536bar, n537bar, n538bar, n539bar, n540bar, n541bar, n542bar, n543bar, n544bar, n545bar, n546bar, n547bar, n548bar, n549bar, n550bar, n551bar, n552bar, n553bar, n554bar, n555bar, n556bar, n557bar, n558bar, n559bar, n560bar, n561bar, n562bar, n563bar, n564bar, n565bar, n566bar, n567bar, n568bar, n569bar, n570bar, n571bar, n572bar, n573bar, n574bar, n575bar, n576bar, n577bar, n578bar, n579bar, n580bar, n581bar, n582bar, n583bar, n584bar, n585bar, n586bar, n587bar, n588bar, n589bar, n590bar, n591bar, n592bar, n593bar, n594bar, n595bar, n596bar, n597bar, n598bar, n599bar, n600bar, n601bar, n602bar, n603bar, n604bar, n605bar, n606bar, n607bar, n608bar, n609bar, n610bar, n611bar, n612bar, n613bar, n614bar, n615bar, n616bar, n617bar, n618bar, n619bar, n620bar, n621bar, n622bar, n623bar, n624bar, n625bar, n626bar, n627bar, n628bar, n629bar, n630bar, n631bar, n632bar, n633bar, n634bar, n635bar, n636bar, n637bar, n638bar, n639bar, n640bar, n641bar, n642bar, n643bar, n644bar, n645bar, n646bar, n647bar, n648bar, n649bar, n650bar, n651bar, n652bar, n653bar, n654bar, n655bar, n656bar, n657bar, n658bar, n659bar, n660bar, n661bar, n662bar, n663bar, n664bar, n665bar, n666bar, n667bar, n668bar, n669bar, n670bar, n671bar, n672bar, n673bar, n674bar, n675bar, n676bar, n677bar, n678bar, n679bar, n680bar, n681bar, n682bar, n683bar, n684bar, n685bar, n686bar, n687bar, n688bar, n689bar, n690bar, n691bar, n692bar, n693bar, n694bar, n695bar, n696bar, n697bar, n698bar, n699bar, n700bar, n701bar, n702bar, n703bar, n704bar, n705bar, n706bar, n707bar, n708bar, n709bar, n710bar, n711bar, n712bar, n713bar, n714bar, n715bar, n716bar, n717bar, n718bar, n719bar, n720bar, n721bar, n722bar, n723bar, n724bar, n725bar, n726bar, n727bar, n728bar, n729bar, n730bar, n731bar, n732bar, n733bar, n734bar, n735bar, n736bar, n737bar, n738bar, n739bar, n740bar, n741bar, n742bar, n743bar, n744bar, n745bar, n746bar, n747bar, n748bar, n749bar, n750bar, n751bar, n752bar, n753bar, n754bar, n755bar, n756bar, n757bar, n758bar, n759bar, n760bar, n761bar, n762bar, n763bar, n764bar, n765bar, n766bar, n767bar, n768bar, n769bar, n770bar, n771bar, n772bar, n773bar, n774bar, n775bar, n776bar, n777bar, n778bar, n779bar, n780bar, n781bar, n782bar, n783bar, n784bar, n785bar, n786bar, n787bar, n788bar, n789bar, n790bar, n791bar, n792bar, n793bar, n794bar, n795bar, n796bar, n797bar, n798bar, n799bar, n800bar, n801bar, n802bar, n803bar, n804bar, n805bar, n806bar, n807bar, n808bar, n809bar, n810bar, n811bar, n812bar, n813bar, n814bar, n815bar, n816bar, n817bar, n818bar, n819bar, n820bar, n821bar, n822bar, n823bar, n824bar, n825bar, n826bar, n827bar, n828bar, n829bar, n830bar, n831bar, n832bar, n833bar, n834bar, n835bar, n836bar, n837bar, n838bar, n839bar, n840bar, n841bar, n842bar, n843bar, n844bar, n845bar, n846bar, n847bar, n848bar, n849bar, n850bar, n851bar, n852bar, n853bar, n854bar, n855bar, n856bar, n857bar, n858bar, n859bar, n860bar, n861bar, n862bar, n863bar, n864bar, n865bar, n866bar, n867bar, n868bar, n869bar, n870bar, n871bar, n872bar, n873bar, n874bar, n875bar, n876bar, n877bar, n878bar, n879bar, n880bar, n881bar, n882bar, n883bar, n884bar, n885bar, n886bar, n887bar, n888bar, n889bar, n890bar, n891bar, n892bar, n893bar, n894bar, n895bar, n896bar, n897bar, n898bar, n899bar, n900bar, n901bar, n902bar, n903bar, n904bar, n905bar, n906bar, n907bar, n908bar, n909bar, n910bar, n911bar, n912bar, n913bar, n914bar, n915bar, n916bar, n917bar, n918bar, n919bar, n920bar, n921bar, n922bar, n923bar, n924bar, n925bar, n926bar, n927bar, n928bar, n929bar, n930bar, n931bar, n932bar, n933bar, n934bar, n935bar, n936bar, n937bar, n938bar, n939bar, n940bar, n941bar, n942bar, n943bar, n944bar, n945bar, n946bar, n947bar, n948bar, n949bar, n950bar, n951bar, n952bar, n953bar, n954bar, n955bar, n956bar, n957bar, n958bar, n959bar, n960bar, n961bar, n962bar, n963bar, n964bar, n965bar, n966bar, n967bar, n968bar, n969bar, n970bar, n971bar, n972bar;
  //wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];

  OR2_X1 U1 ( .A1(n972), .A2(n971), .ZN(out[7]) );
  AND2_X1 U1bar ( .A1(n972bar), .A2(n971bar), .ZN(outbar[7]);
  OR2_X1 U2 ( .A1(n970), .A2(n969), .ZN(n971) );
  AND2_X1 U2bar ( .A1(n970bar), .A2(n969bar), .ZN(n971bar);
  OR2_X1 U3 ( .A1(n968), .A2(n967), .ZN(n969) );
  AND2_X1 U3bar ( .A1(n968bar), .A2(n967bar), .ZN(n969bar);
  OR2_X1 U4 ( .A1(n966), .A2(n965), .ZN(n967) );
  AND2_X1 U4bar ( .A1(n966bar), .A2(n965bar), .ZN(n967bar);
  OR2_X1 U5 ( .A1(n964), .A2(n963), .ZN(n968) );
  AND2_X1 U5bar ( .A1(n964bar), .A2(n963bar), .ZN(n968bar);
  OR2_X1 U6 ( .A1(in[116]), .A2(n962), .ZN(n963) );
  AND2_X1 U6bar ( .A1(inbar[116]), .A2(n962bar), .ZN(n963bar);
  OR2_X1 U7 ( .A1(n961), .A2(n960), .ZN(n970) );
  AND2_X1 U7bar ( .A1(n961bar), .A2(n960bar), .ZN(n970bar);
  OR2_X1 U8 ( .A1(in[150]), .A2(in[127]), .ZN(n960) );
  AND2_X1 U8bar ( .A1(inbar[150]), .A2(inbar[127]), .ZN(n960bar);
  OR2_X1 U9 ( .A1(in[160]), .A2(n959), .ZN(n961) );
  AND2_X1 U9bar ( .A1(inbar[160]), .A2(n959bar), .ZN(n961bar);
  OR2_X1 U10 ( .A1(in[252]), .A2(in[168]), .ZN(n959) );
  AND2_X1 U10bar ( .A1(inbar[252]), .A2(inbar[168]), .ZN(n959bar);
  OR2_X1 U11 ( .A1(n958), .A2(n957), .ZN(n972) );
  AND2_X1 U11bar ( .A1(n958bar), .A2(n957bar), .ZN(n972bar);
  OR2_X1 U12 ( .A1(n956), .A2(n955), .ZN(n957) );
  AND2_X1 U12bar ( .A1(n956bar), .A2(n955bar), .ZN(n957bar);
  OR2_X1 U13 ( .A1(in_17), .A2(in[96]), .ZN(n955) );
  AND2_X1 U13bar ( .A1(in_17bar), .A2(inbar[96]), .ZN(n955bar);
  OR2_X1 U14 ( .A1(in_23), .A2(n954), .ZN(n956) );
  AND2_X1 U14bar ( .A1(in_23bar), .A2(n954bar), .ZN(n956bar);
  OR2_X1 U15 ( .A1(in_31), .A2(in_26), .ZN(n954) );
  AND2_X1 U15bar ( .A1(in_31bar), .A2(in_26bar), .ZN(n954bar);
  OR2_X1 U16 ( .A1(n953), .A2(n952), .ZN(n958) );
  AND2_X1 U16bar ( .A1(n953bar), .A2(n952bar), .ZN(n958bar);
  OR2_X1 U17 ( .A1(in_58), .A2(in_4), .ZN(n952) );
  AND2_X1 U17bar ( .A1(in_58bar), .A2(in_4bar), .ZN(n952bar);
  OR2_X1 U18 ( .A1(in_59), .A2(n951), .ZN(n953) );
  AND2_X1 U18bar ( .A1(in_59bar), .A2(n951bar), .ZN(n953bar);
  OR2_X1 U19 ( .A1(in_71), .A2(in_62), .ZN(n951) );
  AND2_X1 U19bar ( .A1(in_71bar), .A2(in_62bar), .ZN(n951bar);
  OR2_X1 U20 ( .A1(n950), .A2(n949), .ZN(out[6]) );
  AND2_X1 U20bar ( .A1(n950bar), .A2(n949bar), .ZN(outbar[6]);
  OR2_X1 U21 ( .A1(n948), .A2(n947), .ZN(n949) );
  AND2_X1 U21bar ( .A1(n948bar), .A2(n947bar), .ZN(n949bar);
  OR2_X1 U22 ( .A1(n946), .A2(n945), .ZN(n947) );
  AND2_X1 U22bar ( .A1(n946bar), .A2(n945bar), .ZN(n947bar);
  OR2_X1 U23 ( .A1(n944), .A2(n943), .ZN(n945) );
  AND2_X1 U23bar ( .A1(n944bar), .A2(n943bar), .ZN(n945bar);
  OR2_X1 U24 ( .A1(n942), .A2(n941), .ZN(n946) );
  AND2_X1 U24bar ( .A1(n942bar), .A2(n941bar), .ZN(n946bar);
  OR2_X1 U25 ( .A1(in[101]), .A2(n940), .ZN(n941) );
  AND2_X1 U25bar ( .A1(inbar[101]), .A2(n940bar), .ZN(n941bar);
  OR2_X1 U26 ( .A1(n939), .A2(n938), .ZN(n948) );
  AND2_X1 U26bar ( .A1(n939bar), .A2(n938bar), .ZN(n948bar);
  OR2_X1 U27 ( .A1(in[114]), .A2(in[104]), .ZN(n938) );
  AND2_X1 U27bar ( .A1(inbar[114]), .A2(inbar[104]), .ZN(n938bar);
  OR2_X1 U28 ( .A1(in[128]), .A2(n937), .ZN(n939) );
  AND2_X1 U28bar ( .A1(inbar[128]), .A2(n937bar), .ZN(n939bar);
  OR2_X1 U29 ( .A1(in[136]), .A2(in[134]), .ZN(n937) );
  AND2_X1 U29bar ( .A1(inbar[136]), .A2(inbar[134]), .ZN(n937bar);
  OR2_X1 U30 ( .A1(n936), .A2(n935), .ZN(n950) );
  AND2_X1 U30bar ( .A1(n936bar), .A2(n935bar), .ZN(n950bar);
  OR2_X1 U31 ( .A1(n934), .A2(n933), .ZN(n935) );
  AND2_X1 U31bar ( .A1(n934bar), .A2(n933bar), .ZN(n935bar);
  OR2_X1 U32 ( .A1(in[177]), .A2(in[164]), .ZN(n933) );
  AND2_X1 U32bar ( .A1(inbar[177]), .A2(inbar[164]), .ZN(n933bar);
  OR2_X1 U33 ( .A1(in[212]), .A2(n932), .ZN(n934) );
  AND2_X1 U33bar ( .A1(inbar[212]), .A2(n932bar), .ZN(n934bar);
  OR2_X1 U34 ( .A1(in[248]), .A2(in[221]), .ZN(n932) );
  AND2_X1 U34bar ( .A1(inbar[248]), .A2(inbar[221]), .ZN(n932bar);
  OR2_X1 U35 ( .A1(n931), .A2(n930), .ZN(n936) );
  AND2_X1 U35bar ( .A1(n931bar), .A2(n930bar), .ZN(n936bar);
  OR2_X1 U36 ( .A1(in_18), .A2(in[93]), .ZN(n930) );
  AND2_X1 U36bar ( .A1(in_18bar), .A2(inbar[93]), .ZN(n930bar);
  OR2_X1 U37 ( .A1(in_31), .A2(n929), .ZN(n931) );
  AND2_X1 U37bar ( .A1(in_31bar), .A2(n929bar), .ZN(n931bar);
  OR2_X1 U38 ( .A1(in_7), .A2(in_39), .ZN(n929) );
  AND2_X1 U38bar ( .A1(in_7bar), .A2(in_39bar), .ZN(n929bar);
  OR2_X1 U39 ( .A1(n928), .A2(n927), .ZN(out[5]) );
  AND2_X1 U39bar ( .A1(n928bar), .A2(n927bar), .ZN(outbar[5]);
  OR2_X1 U40 ( .A1(n926), .A2(n925), .ZN(n927) );
  AND2_X1 U40bar ( .A1(n926bar), .A2(n925bar), .ZN(n927bar);
  OR2_X1 U41 ( .A1(n924), .A2(n923), .ZN(n925) );
  AND2_X1 U41bar ( .A1(n924bar), .A2(n923bar), .ZN(n925bar);
  OR2_X1 U42 ( .A1(n922), .A2(n921), .ZN(n923) );
  AND2_X1 U42bar ( .A1(n922bar), .A2(n921bar), .ZN(n923bar);
  OR2_X1 U43 ( .A1(n940), .A2(n920), .ZN(n924) );
  AND2_X1 U43bar ( .A1(n940bar), .A2(n920bar), .ZN(n924bar);
  OR2_X1 U44 ( .A1(in[111]), .A2(n919), .ZN(n920) );
  AND2_X1 U44bar ( .A1(inbar[111]), .A2(n919bar), .ZN(n920bar);
  OR2_X1 U45 ( .A1(n918), .A2(n917), .ZN(n940) );
  AND2_X1 U45bar ( .A1(n918bar), .A2(n917bar), .ZN(n940bar);
  OR2_X1 U46 ( .A1(n916), .A2(n915), .ZN(n917) );
  AND2_X1 U46bar ( .A1(n916bar), .A2(n915bar), .ZN(n917bar);
  OR2_X1 U47 ( .A1(n914), .A2(n913), .ZN(n915) );
  AND2_X1 U47bar ( .A1(n914bar), .A2(n913bar), .ZN(n915bar);
  OR2_X1 U48 ( .A1(in[140]), .A2(in[131]), .ZN(n913) );
  AND2_X1 U48bar ( .A1(inbar[140]), .A2(inbar[131]), .ZN(n913bar);
  OR2_X1 U49 ( .A1(in[160]), .A2(in[144]), .ZN(n914) );
  AND2_X1 U49bar ( .A1(inbar[160]), .A2(inbar[144]), .ZN(n914bar);
  OR2_X1 U50 ( .A1(n912), .A2(n911), .ZN(n916) );
  AND2_X1 U50bar ( .A1(n912bar), .A2(n911bar), .ZN(n916bar);
  OR2_X1 U51 ( .A1(in[179]), .A2(in[174]), .ZN(n911) );
  AND2_X1 U51bar ( .A1(inbar[179]), .A2(inbar[174]), .ZN(n911bar);
  OR2_X1 U52 ( .A1(in[188]), .A2(in[184]), .ZN(n912) );
  AND2_X1 U52bar ( .A1(inbar[188]), .A2(inbar[184]), .ZN(n912bar);
  OR2_X1 U53 ( .A1(n910), .A2(n909), .ZN(n918) );
  AND2_X1 U53bar ( .A1(n910bar), .A2(n909bar), .ZN(n918bar);
  OR2_X1 U54 ( .A1(n908), .A2(n907), .ZN(n909) );
  AND2_X1 U54bar ( .A1(n908bar), .A2(n907bar), .ZN(n909bar);
  OR2_X1 U55 ( .A1(in[216]), .A2(in[200]), .ZN(n907) );
  AND2_X1 U55bar ( .A1(inbar[216]), .A2(inbar[200]), .ZN(n907bar);
  OR2_X1 U56 ( .A1(in[228]), .A2(in[224]), .ZN(n908) );
  AND2_X1 U56bar ( .A1(inbar[228]), .A2(inbar[224]), .ZN(n908bar);
  OR2_X1 U57 ( .A1(n906), .A2(n905), .ZN(n910) );
  AND2_X1 U57bar ( .A1(n906bar), .A2(n905bar), .ZN(n910bar);
  OR2_X1 U58 ( .A1(in[247]), .A2(in[235]), .ZN(n905) );
  AND2_X1 U58bar ( .A1(inbar[247]), .A2(inbar[235]), .ZN(n905bar);
  OR2_X1 U59 ( .A1(in_42), .A2(in[83]), .ZN(n906) );
  AND2_X1 U59bar ( .A1(in_42bar), .A2(inbar[83]), .ZN(n906bar);
  OR2_X1 U60 ( .A1(n904), .A2(n903), .ZN(n926) );
  AND2_X1 U60bar ( .A1(n904bar), .A2(n903bar), .ZN(n926bar);
  OR2_X1 U61 ( .A1(in[166]), .A2(in[123]), .ZN(n903) );
  AND2_X1 U61bar ( .A1(inbar[166]), .A2(inbar[123]), .ZN(n903bar);
  OR2_X1 U62 ( .A1(in[170]), .A2(n902), .ZN(n904) );
  AND2_X1 U62bar ( .A1(inbar[170]), .A2(n902bar), .ZN(n904bar);
  OR2_X1 U63 ( .A1(in[194]), .A2(in[183]), .ZN(n902) );
  AND2_X1 U63bar ( .A1(inbar[194]), .A2(inbar[183]), .ZN(n902bar);
  OR2_X1 U64 ( .A1(n901), .A2(n900), .ZN(n928) );
  AND2_X1 U64bar ( .A1(n901bar), .A2(n900bar), .ZN(n928bar);
  OR2_X1 U65 ( .A1(n899), .A2(n898), .ZN(n900) );
  AND2_X1 U65bar ( .A1(n899bar), .A2(n898bar), .ZN(n900bar);
  OR2_X1 U66 ( .A1(in[241]), .A2(in[238]), .ZN(n898) );
  AND2_X1 U66bar ( .A1(inbar[241]), .A2(inbar[238]), .ZN(n898bar);
  OR2_X1 U67 ( .A1(in[250]), .A2(n897), .ZN(n899) );
  AND2_X1 U67bar ( .A1(inbar[250]), .A2(n897bar), .ZN(n899bar);
  OR2_X1 U68 ( .A1(in_24), .A2(in[84]), .ZN(n897) );
  AND2_X1 U68bar ( .A1(in_24bar), .A2(inbar[84]), .ZN(n897bar);
  OR2_X1 U69 ( .A1(n896), .A2(n895), .ZN(n901) );
  AND2_X1 U69bar ( .A1(n896bar), .A2(n895bar), .ZN(n901bar);
  OR2_X1 U70 ( .A1(in_41), .A2(in_29), .ZN(n895) );
  AND2_X1 U70bar ( .A1(in_41bar), .A2(in_29bar), .ZN(n895bar);
  OR2_X1 U71 ( .A1(in_66), .A2(n894), .ZN(n896) );
  AND2_X1 U71bar ( .A1(in_66bar), .A2(n894bar), .ZN(n896bar);
  OR2_X1 U72 ( .A1(in_76), .A2(in_71), .ZN(n894) );
  AND2_X1 U72bar ( .A1(in_76bar), .A2(in_71bar), .ZN(n894bar);
  OR2_X1 U73 ( .A1(n893), .A2(n892), .ZN(out[4]) );
  AND2_X1 U73bar ( .A1(n893bar), .A2(n892bar), .ZN(outbar[4]);
  OR2_X1 U74 ( .A1(n891), .A2(n890), .ZN(n892) );
  AND2_X1 U74bar ( .A1(n891bar), .A2(n890bar), .ZN(n892bar);
  OR2_X1 U75 ( .A1(n889), .A2(n888), .ZN(n890) );
  AND2_X1 U75bar ( .A1(n889bar), .A2(n888bar), .ZN(n890bar);
  OR2_X1 U76 ( .A1(n922), .A2(n887), .ZN(n888) );
  AND2_X1 U76bar ( .A1(n922bar), .A2(n887bar), .ZN(n888bar);
  OR2_X1 U77 ( .A1(n886), .A2(n885), .ZN(n922) );
  AND2_X1 U77bar ( .A1(n886bar), .A2(n885bar), .ZN(n922bar);
  OR2_X1 U78 ( .A1(n884), .A2(n883), .ZN(n885) );
  AND2_X1 U78bar ( .A1(n884bar), .A2(n883bar), .ZN(n885bar);
  OR2_X1 U79 ( .A1(n882), .A2(n881), .ZN(n883) );
  AND2_X1 U79bar ( .A1(n882bar), .A2(n881bar), .ZN(n883bar);
  OR2_X1 U80 ( .A1(in[118]), .A2(in[109]), .ZN(n881) );
  AND2_X1 U80bar ( .A1(inbar[118]), .A2(inbar[109]), .ZN(n881bar);
  OR2_X1 U81 ( .A1(in[139]), .A2(in[120]), .ZN(n882) );
  AND2_X1 U81bar ( .A1(inbar[139]), .A2(inbar[120]), .ZN(n882bar);
  OR2_X1 U82 ( .A1(n880), .A2(n879), .ZN(n884) );
  AND2_X1 U82bar ( .A1(n880bar), .A2(n879bar), .ZN(n884bar);
  OR2_X1 U83 ( .A1(in[198]), .A2(in[154]), .ZN(n879) );
  AND2_X1 U83bar ( .A1(inbar[198]), .A2(inbar[154]), .ZN(n879bar);
  OR2_X1 U84 ( .A1(in[210]), .A2(in[205]), .ZN(n880) );
  AND2_X1 U84bar ( .A1(inbar[210]), .A2(inbar[205]), .ZN(n880bar);
  OR2_X1 U85 ( .A1(n878), .A2(n877), .ZN(n886) );
  AND2_X1 U85bar ( .A1(n878bar), .A2(n877bar), .ZN(n886bar);
  OR2_X1 U86 ( .A1(n876), .A2(n875), .ZN(n877) );
  AND2_X1 U86bar ( .A1(n876bar), .A2(n875bar), .ZN(n877bar);
  OR2_X1 U87 ( .A1(in[219]), .A2(in[217]), .ZN(n875) );
  AND2_X1 U87bar ( .A1(inbar[219]), .A2(inbar[217]), .ZN(n875bar);
  OR2_X1 U88 ( .A1(in[86]), .A2(in[252]), .ZN(n876) );
  AND2_X1 U88bar ( .A1(inbar[86]), .A2(inbar[252]), .ZN(n876bar);
  OR2_X1 U89 ( .A1(n874), .A2(n873), .ZN(n878) );
  AND2_X1 U89bar ( .A1(n874bar), .A2(n873bar), .ZN(n878bar);
  OR2_X1 U90 ( .A1(in_40), .A2(in[91]), .ZN(n873) );
  AND2_X1 U90bar ( .A1(in_40bar), .A2(inbar[91]), .ZN(n873bar);
  OR2_X1 U91 ( .A1(in_8), .A2(in_46), .ZN(n874) );
  AND2_X1 U91bar ( .A1(in_8bar), .A2(in_46bar), .ZN(n874bar);
  OR2_X1 U92 ( .A1(n872), .A2(n871), .ZN(n889) );
  AND2_X1 U92bar ( .A1(n872bar), .A2(n871bar), .ZN(n889bar);
  OR2_X1 U93 ( .A1(in[117]), .A2(n943), .ZN(n871) );
  AND2_X1 U93bar ( .A1(inbar[117]), .A2(n943bar), .ZN(n871bar);
  OR2_X1 U94 ( .A1(n870), .A2(n869), .ZN(n943) );
  AND2_X1 U94bar ( .A1(n870bar), .A2(n869bar), .ZN(n943bar);
  OR2_X1 U95 ( .A1(n868), .A2(n867), .ZN(n869) );
  AND2_X1 U95bar ( .A1(n868bar), .A2(n867bar), .ZN(n869bar);
  OR2_X1 U96 ( .A1(n866), .A2(n865), .ZN(n867) );
  AND2_X1 U96bar ( .A1(n866bar), .A2(n865bar), .ZN(n867bar);
  OR2_X1 U97 ( .A1(n864), .A2(n863), .ZN(n865) );
  AND2_X1 U97bar ( .A1(n864bar), .A2(n863bar), .ZN(n865bar);
  OR2_X1 U98 ( .A1(in[108]), .A2(n919), .ZN(n866) );
  AND2_X1 U98bar ( .A1(inbar[108]), .A2(n919bar), .ZN(n866bar);
  OR2_X1 U99 ( .A1(n862), .A2(n861), .ZN(n919) );
  AND2_X1 U99bar ( .A1(n862bar), .A2(n861bar), .ZN(n919bar);
  OR2_X1 U100 ( .A1(n860), .A2(n859), .ZN(n861) );
  AND2_X1 U100bar ( .A1(n860bar), .A2(n859bar), .ZN(n861bar);
  OR2_X1 U101 ( .A1(n858), .A2(n857), .ZN(n859) );
  AND2_X1 U101bar ( .A1(n858bar), .A2(n857bar), .ZN(n859bar);
  OR2_X1 U102 ( .A1(in[119]), .A2(in[105]), .ZN(n857) );
  AND2_X1 U102bar ( .A1(inbar[119]), .A2(inbar[105]), .ZN(n857bar);
  OR2_X1 U103 ( .A1(in[186]), .A2(in[175]), .ZN(n858) );
  AND2_X1 U103bar ( .A1(inbar[186]), .A2(inbar[175]), .ZN(n858bar);
  OR2_X1 U104 ( .A1(n856), .A2(n855), .ZN(n860) );
  AND2_X1 U104bar ( .A1(n856bar), .A2(n855bar), .ZN(n860bar);
  OR2_X1 U105 ( .A1(in[202]), .A2(in[193]), .ZN(n855) );
  AND2_X1 U105bar ( .A1(inbar[202]), .A2(inbar[193]), .ZN(n855bar);
  OR2_X1 U106 ( .A1(in[225]), .A2(in[208]), .ZN(n856) );
  AND2_X1 U106bar ( .A1(inbar[225]), .A2(inbar[208]), .ZN(n856bar);
  OR2_X1 U107 ( .A1(n854), .A2(n853), .ZN(n862) );
  AND2_X1 U107bar ( .A1(n854bar), .A2(n853bar), .ZN(n862bar);
  OR2_X1 U108 ( .A1(n852), .A2(n851), .ZN(n853) );
  AND2_X1 U108bar ( .A1(n852bar), .A2(n851bar), .ZN(n853bar);
  OR2_X1 U109 ( .A1(in_1), .A2(in[85]), .ZN(n851) );
  AND2_X1 U109bar ( .A1(in_1bar), .A2(inbar[85]), .ZN(n851bar);
  OR2_X1 U110 ( .A1(in_23), .A2(in_19), .ZN(n852) );
  AND2_X1 U110bar ( .A1(in_23bar), .A2(in_19bar), .ZN(n852bar);
  OR2_X1 U111 ( .A1(n850), .A2(n849), .ZN(n854) );
  AND2_X1 U111bar ( .A1(n850bar), .A2(n849bar), .ZN(n854bar);
  OR2_X1 U112 ( .A1(in_43), .A2(in_33), .ZN(n849) );
  AND2_X1 U112bar ( .A1(in_43bar), .A2(in_33bar), .ZN(n849bar);
  OR2_X1 U113 ( .A1(in_63), .A2(in_44), .ZN(n850) );
  AND2_X1 U113bar ( .A1(in_63bar), .A2(in_44bar), .ZN(n850bar);
  OR2_X1 U114 ( .A1(n848), .A2(n847), .ZN(n868) );
  AND2_X1 U114bar ( .A1(n848bar), .A2(n847bar), .ZN(n868bar);
  OR2_X1 U115 ( .A1(in[141]), .A2(in[112]), .ZN(n847) );
  AND2_X1 U115bar ( .A1(inbar[141]), .A2(inbar[112]), .ZN(n847bar);
  OR2_X1 U116 ( .A1(in[147]), .A2(n846), .ZN(n848) );
  AND2_X1 U116bar ( .A1(inbar[147]), .A2(n846bar), .ZN(n848bar);
  OR2_X1 U117 ( .A1(in[181]), .A2(in[167]), .ZN(n846) );
  AND2_X1 U117bar ( .A1(inbar[181]), .A2(inbar[167]), .ZN(n846bar);
  OR2_X1 U118 ( .A1(n845), .A2(n844), .ZN(n870) );
  AND2_X1 U118bar ( .A1(n845bar), .A2(n844bar), .ZN(n870bar);
  OR2_X1 U119 ( .A1(n843), .A2(n842), .ZN(n844) );
  AND2_X1 U119bar ( .A1(n843bar), .A2(n842bar), .ZN(n844bar);
  OR2_X1 U120 ( .A1(in[229]), .A2(in[201]), .ZN(n842) );
  AND2_X1 U120bar ( .A1(inbar[229]), .A2(inbar[201]), .ZN(n842bar);
  OR2_X1 U121 ( .A1(in[237]), .A2(n841), .ZN(n843) );
  AND2_X1 U121bar ( .A1(inbar[237]), .A2(n841bar), .ZN(n843bar);
  OR2_X1 U122 ( .A1(in[94]), .A2(in[253]), .ZN(n841) );
  AND2_X1 U122bar ( .A1(inbar[94]), .A2(inbar[253]), .ZN(n841bar);
  OR2_X1 U123 ( .A1(n840), .A2(n839), .ZN(n845) );
  AND2_X1 U123bar ( .A1(n840bar), .A2(n839bar), .ZN(n845bar);
  OR2_X1 U124 ( .A1(in_21), .A2(in[96]), .ZN(n839) );
  AND2_X1 U124bar ( .A1(in_21bar), .A2(inbar[96]), .ZN(n839bar);
  OR2_X1 U125 ( .A1(in_25), .A2(n838), .ZN(n840) );
  AND2_X1 U125bar ( .A1(in_25bar), .A2(n838bar), .ZN(n840bar);
  OR2_X1 U126 ( .A1(in_81), .A2(in_45), .ZN(n838) );
  AND2_X1 U126bar ( .A1(in_81bar), .A2(in_45bar), .ZN(n838bar);
  OR2_X1 U127 ( .A1(n837), .A2(n836), .ZN(n891) );
  AND2_X1 U127bar ( .A1(n837bar), .A2(n836bar), .ZN(n891bar);
  OR2_X1 U128 ( .A1(in[142]), .A2(in[124]), .ZN(n836) );
  AND2_X1 U128bar ( .A1(inbar[142]), .A2(inbar[124]), .ZN(n836bar);
  OR2_X1 U129 ( .A1(in[150]), .A2(n835), .ZN(n837) );
  AND2_X1 U129bar ( .A1(inbar[150]), .A2(n835bar), .ZN(n837bar);
  OR2_X1 U130 ( .A1(in[172]), .A2(in[155]), .ZN(n835) );
  AND2_X1 U130bar ( .A1(inbar[172]), .A2(inbar[155]), .ZN(n835bar);
  OR2_X1 U131 ( .A1(n834), .A2(n833), .ZN(n893) );
  AND2_X1 U131bar ( .A1(n834bar), .A2(n833bar), .ZN(n893bar);
  OR2_X1 U132 ( .A1(n832), .A2(n831), .ZN(n833) );
  AND2_X1 U132bar ( .A1(n832bar), .A2(n831bar), .ZN(n833bar);
  OR2_X1 U133 ( .A1(in[196]), .A2(in[173]), .ZN(n831) );
  AND2_X1 U133bar ( .A1(inbar[196]), .A2(inbar[173]), .ZN(n831bar);
  OR2_X1 U134 ( .A1(in[222]), .A2(n830), .ZN(n832) );
  AND2_X1 U134bar ( .A1(inbar[222]), .A2(n830bar), .ZN(n832bar);
  OR2_X1 U135 ( .A1(in[227]), .A2(in[226]), .ZN(n830) );
  AND2_X1 U135bar ( .A1(inbar[227]), .A2(inbar[226]), .ZN(n830bar);
  OR2_X1 U136 ( .A1(n829), .A2(n828), .ZN(n834) );
  AND2_X1 U136bar ( .A1(n829bar), .A2(n828bar), .ZN(n834bar);
  OR2_X1 U137 ( .A1(in[249]), .A2(in[231]), .ZN(n828) );
  AND2_X1 U137bar ( .A1(inbar[249]), .A2(inbar[231]), .ZN(n828bar);
  OR2_X1 U138 ( .A1(in_28), .A2(n827), .ZN(n829) );
  AND2_X1 U138bar ( .A1(in_28bar), .A2(n827bar), .ZN(n829bar);
  OR2_X1 U139 ( .A1(in_52), .A2(in_47), .ZN(n827) );
  AND2_X1 U139bar ( .A1(in_52bar), .A2(in_47bar), .ZN(n827bar);
  OR2_X1 U140 ( .A1(n826), .A2(n825), .ZN(out[3]) );
  AND2_X1 U140bar ( .A1(n826bar), .A2(n825bar), .ZN(outbar[3]);
  OR2_X1 U141 ( .A1(n824), .A2(n823), .ZN(n825) );
  AND2_X1 U141bar ( .A1(n824bar), .A2(n823bar), .ZN(n825bar);
  OR2_X1 U142 ( .A1(n822), .A2(n821), .ZN(n823) );
  AND2_X1 U142bar ( .A1(n822bar), .A2(n821bar), .ZN(n823bar);
  OR2_X1 U143 ( .A1(n820), .A2(n819), .ZN(n821) );
  AND2_X1 U143bar ( .A1(n820bar), .A2(n819bar), .ZN(n821bar);
  OR2_X1 U144 ( .A1(n964), .A2(n818), .ZN(n822) );
  AND2_X1 U144bar ( .A1(n964bar), .A2(n818bar), .ZN(n822bar);
  OR2_X1 U145 ( .A1(in[118]), .A2(n817), .ZN(n818) );
  AND2_X1 U145bar ( .A1(inbar[118]), .A2(n817bar), .ZN(n818bar);
  OR2_X1 U146 ( .A1(n816), .A2(n815), .ZN(n964) );
  AND2_X1 U146bar ( .A1(n816bar), .A2(n815bar), .ZN(n964bar);
  OR2_X1 U147 ( .A1(n814), .A2(n813), .ZN(n815) );
  AND2_X1 U147bar ( .A1(n814bar), .A2(n813bar), .ZN(n815bar);
  OR2_X1 U148 ( .A1(n812), .A2(n811), .ZN(n813) );
  AND2_X1 U148bar ( .A1(n812bar), .A2(n811bar), .ZN(n813bar);
  OR2_X1 U149 ( .A1(in[122]), .A2(in[111]), .ZN(n811) );
  AND2_X1 U149bar ( .A1(inbar[122]), .A2(inbar[111]), .ZN(n811bar);
  OR2_X1 U150 ( .A1(in[154]), .A2(in[151]), .ZN(n812) );
  AND2_X1 U150bar ( .A1(inbar[154]), .A2(inbar[151]), .ZN(n812bar);
  OR2_X1 U151 ( .A1(n810), .A2(n809), .ZN(n814) );
  AND2_X1 U151bar ( .A1(n810bar), .A2(n809bar), .ZN(n814bar);
  OR2_X1 U152 ( .A1(in[187]), .A2(in[177]), .ZN(n809) );
  AND2_X1 U152bar ( .A1(inbar[187]), .A2(inbar[177]), .ZN(n809bar);
  OR2_X1 U153 ( .A1(in[200]), .A2(in[192]), .ZN(n810) );
  AND2_X1 U153bar ( .A1(inbar[200]), .A2(inbar[192]), .ZN(n810bar);
  OR2_X1 U154 ( .A1(n808), .A2(n807), .ZN(n816) );
  AND2_X1 U154bar ( .A1(n808bar), .A2(n807bar), .ZN(n816bar);
  OR2_X1 U155 ( .A1(n806), .A2(n805), .ZN(n807) );
  AND2_X1 U155bar ( .A1(n806bar), .A2(n805bar), .ZN(n807bar);
  OR2_X1 U156 ( .A1(in[225]), .A2(in[207]), .ZN(n805) );
  AND2_X1 U156bar ( .A1(inbar[225]), .A2(inbar[207]), .ZN(n805bar);
  OR2_X1 U157 ( .A1(in[98]), .A2(in[226]), .ZN(n806) );
  AND2_X1 U157bar ( .A1(inbar[98]), .A2(inbar[226]), .ZN(n806bar);
  OR2_X1 U158 ( .A1(n804), .A2(n803), .ZN(n808) );
  AND2_X1 U158bar ( .A1(n804bar), .A2(n803bar), .ZN(n808bar);
  OR2_X1 U159 ( .A1(in_20), .A2(in_16), .ZN(n803) );
  AND2_X1 U159bar ( .A1(in_20bar), .A2(in_16bar), .ZN(n803bar);
  OR2_X1 U160 ( .A1(in_55), .A2(in_45), .ZN(n804) );
  AND2_X1 U160bar ( .A1(in_55bar), .A2(in_45bar), .ZN(n804bar);
  OR2_X1 U161 ( .A1(n802), .A2(n801), .ZN(n824) );
  AND2_X1 U161bar ( .A1(n802bar), .A2(n801bar), .ZN(n824bar);
  OR2_X1 U162 ( .A1(in[162]), .A2(in[149]), .ZN(n801) );
  AND2_X1 U162bar ( .A1(inbar[162]), .A2(inbar[149]), .ZN(n801bar);
  OR2_X1 U163 ( .A1(in[163]), .A2(n800), .ZN(n802) );
  AND2_X1 U163bar ( .A1(inbar[163]), .A2(n800bar), .ZN(n802bar);
  OR2_X1 U164 ( .A1(in[191]), .A2(in[189]), .ZN(n800) );
  AND2_X1 U164bar ( .A1(inbar[191]), .A2(inbar[189]), .ZN(n800bar);
  OR2_X1 U165 ( .A1(n799), .A2(n798), .ZN(n826) );
  AND2_X1 U165bar ( .A1(n799bar), .A2(n798bar), .ZN(n826bar);
  OR2_X1 U166 ( .A1(n797), .A2(n796), .ZN(n798) );
  AND2_X1 U166bar ( .A1(n797bar), .A2(n796bar), .ZN(n798bar);
  OR2_X1 U167 ( .A1(in[212]), .A2(in[193]), .ZN(n796) );
  AND2_X1 U167bar ( .A1(inbar[212]), .A2(inbar[193]), .ZN(n796bar);
  OR2_X1 U168 ( .A1(in[238]), .A2(n795), .ZN(n797) );
  AND2_X1 U168bar ( .A1(inbar[238]), .A2(n795bar), .ZN(n797bar);
  OR2_X1 U169 ( .A1(in[88]), .A2(in[247]), .ZN(n795) );
  AND2_X1 U169bar ( .A1(inbar[88]), .A2(inbar[247]), .ZN(n795bar);
  OR2_X1 U170 ( .A1(n794), .A2(n793), .ZN(n799) );
  AND2_X1 U170bar ( .A1(n794bar), .A2(n793bar), .ZN(n799bar);
  OR2_X1 U171 ( .A1(in[94]), .A2(in[92]), .ZN(n793) );
  AND2_X1 U171bar ( .A1(inbar[94]), .A2(inbar[92]), .ZN(n793bar);
  OR2_X1 U172 ( .A1(in_52), .A2(n792), .ZN(n794) );
  AND2_X1 U172bar ( .A1(in_52bar), .A2(n792bar), .ZN(n794bar);
  OR2_X1 U173 ( .A1(in_70), .A2(in_67), .ZN(n792) );
  AND2_X1 U173bar ( .A1(in_70bar), .A2(in_67bar), .ZN(n792bar);
  OR2_X1 U174 ( .A1(n791), .A2(n790), .ZN(out[2]) );
  AND2_X1 U174bar ( .A1(n791bar), .A2(n790bar), .ZN(outbar[2]);
  OR2_X1 U175 ( .A1(n789), .A2(n788), .ZN(n790) );
  AND2_X1 U175bar ( .A1(n789bar), .A2(n788bar), .ZN(n790bar);
  OR2_X1 U176 ( .A1(n787), .A2(n786), .ZN(n788) );
  AND2_X1 U176bar ( .A1(n787bar), .A2(n786bar), .ZN(n788bar);
  OR2_X1 U177 ( .A1(n819), .A2(n785), .ZN(n786) );
  AND2_X1 U177bar ( .A1(n819bar), .A2(n785bar), .ZN(n786bar);
  OR2_X1 U178 ( .A1(n784), .A2(n783), .ZN(n819) );
  AND2_X1 U178bar ( .A1(n784bar), .A2(n783bar), .ZN(n819bar);
  OR2_X1 U179 ( .A1(n782), .A2(n781), .ZN(n783) );
  AND2_X1 U179bar ( .A1(n782bar), .A2(n781bar), .ZN(n783bar);
  OR2_X1 U180 ( .A1(n780), .A2(n779), .ZN(n781) );
  AND2_X1 U180bar ( .A1(n780bar), .A2(n779bar), .ZN(n781bar);
  OR2_X1 U181 ( .A1(n962), .A2(n778), .ZN(n779) );
  AND2_X1 U181bar ( .A1(n962bar), .A2(n778bar), .ZN(n779bar);
  OR2_X1 U182 ( .A1(n777), .A2(n776), .ZN(n962) );
  AND2_X1 U182bar ( .A1(n777bar), .A2(n776bar), .ZN(n962bar);
  OR2_X1 U183 ( .A1(n775), .A2(n774), .ZN(n776) );
  AND2_X1 U183bar ( .A1(n775bar), .A2(n774bar), .ZN(n776bar);
  OR2_X1 U184 ( .A1(n773), .A2(n772), .ZN(n774) );
  AND2_X1 U184bar ( .A1(n773bar), .A2(n772bar), .ZN(n774bar);
  OR2_X1 U185 ( .A1(in[131]), .A2(in[120]), .ZN(n772) );
  AND2_X1 U185bar ( .A1(inbar[131]), .A2(inbar[120]), .ZN(n772bar);
  OR2_X1 U186 ( .A1(in[153]), .A2(in[147]), .ZN(n773) );
  AND2_X1 U186bar ( .A1(inbar[153]), .A2(inbar[147]), .ZN(n773bar);
  OR2_X1 U187 ( .A1(n771), .A2(n770), .ZN(n775) );
  AND2_X1 U187bar ( .A1(n771bar), .A2(n770bar), .ZN(n775bar);
  OR2_X1 U188 ( .A1(in[170]), .A2(in[156]), .ZN(n770) );
  AND2_X1 U188bar ( .A1(inbar[170]), .A2(inbar[156]), .ZN(n770bar);
  OR2_X1 U189 ( .A1(in[223]), .A2(in[190]), .ZN(n771) );
  AND2_X1 U189bar ( .A1(inbar[223]), .A2(inbar[190]), .ZN(n771bar);
  OR2_X1 U190 ( .A1(n769), .A2(n768), .ZN(n777) );
  AND2_X1 U190bar ( .A1(n769bar), .A2(n768bar), .ZN(n777bar);
  OR2_X1 U191 ( .A1(n767), .A2(n766), .ZN(n768) );
  AND2_X1 U191bar ( .A1(n767bar), .A2(n766bar), .ZN(n768bar);
  OR2_X1 U192 ( .A1(in[236]), .A2(in[230]), .ZN(n766) );
  AND2_X1 U192bar ( .A1(inbar[236]), .A2(inbar[230]), .ZN(n766bar);
  OR2_X1 U193 ( .A1(in[85]), .A2(in[240]), .ZN(n767) );
  AND2_X1 U193bar ( .A1(inbar[85]), .A2(inbar[240]), .ZN(n767bar);
  OR2_X1 U194 ( .A1(n765), .A2(n764), .ZN(n769) );
  AND2_X1 U194bar ( .A1(n765bar), .A2(n764bar), .ZN(n769bar);
  OR2_X1 U195 ( .A1(in_12), .A2(in[90]), .ZN(n764) );
  AND2_X1 U195bar ( .A1(in_12bar), .A2(inbar[90]), .ZN(n764bar);
  OR2_X1 U196 ( .A1(in_39), .A2(in_28), .ZN(n765) );
  AND2_X1 U196bar ( .A1(in_39bar), .A2(in_28bar), .ZN(n765bar);
  OR2_X1 U197 ( .A1(in[109]), .A2(n763), .ZN(n780) );
  AND2_X1 U197bar ( .A1(inbar[109]), .A2(n763bar), .ZN(n780bar);
  OR2_X1 U198 ( .A1(n762), .A2(n761), .ZN(n782) );
  AND2_X1 U198bar ( .A1(n762bar), .A2(n761bar), .ZN(n782bar);
  OR2_X1 U199 ( .A1(in[138]), .A2(in[129]), .ZN(n761) );
  AND2_X1 U199bar ( .A1(inbar[138]), .A2(inbar[129]), .ZN(n761bar);
  OR2_X1 U200 ( .A1(in[157]), .A2(n760), .ZN(n762) );
  AND2_X1 U200bar ( .A1(inbar[157]), .A2(n760bar), .ZN(n762bar);
  OR2_X1 U201 ( .A1(in[182]), .A2(in[167]), .ZN(n760) );
  AND2_X1 U201bar ( .A1(inbar[182]), .A2(inbar[167]), .ZN(n760bar);
  OR2_X1 U202 ( .A1(n759), .A2(n758), .ZN(n784) );
  AND2_X1 U202bar ( .A1(n759bar), .A2(n758bar), .ZN(n784bar);
  OR2_X1 U203 ( .A1(n757), .A2(n756), .ZN(n758) );
  AND2_X1 U203bar ( .A1(n757bar), .A2(n756bar), .ZN(n758bar);
  OR2_X1 U204 ( .A1(in[195]), .A2(in[184]), .ZN(n756) );
  AND2_X1 U204bar ( .A1(inbar[195]), .A2(inbar[184]), .ZN(n756bar);
  OR2_X1 U205 ( .A1(in[196]), .A2(n755), .ZN(n757) );
  AND2_X1 U205bar ( .A1(inbar[196]), .A2(n755bar), .ZN(n757bar);
  OR2_X1 U206 ( .A1(in[215]), .A2(in[209]), .ZN(n755) );
  AND2_X1 U206bar ( .A1(inbar[215]), .A2(inbar[209]), .ZN(n755bar);
  OR2_X1 U207 ( .A1(n754), .A2(n753), .ZN(n759) );
  AND2_X1 U207bar ( .A1(n754bar), .A2(n753bar), .ZN(n759bar);
  OR2_X1 U208 ( .A1(in[93]), .A2(in[233]), .ZN(n753) );
  AND2_X1 U208bar ( .A1(inbar[93]), .A2(inbar[233]), .ZN(n753bar);
  OR2_X1 U209 ( .A1(in_1), .A2(n752), .ZN(n754) );
  AND2_X1 U209bar ( .A1(in_1bar), .A2(n752bar), .ZN(n754bar);
  OR2_X1 U210 ( .A1(in_69), .A2(in_66), .ZN(n752) );
  AND2_X1 U210bar ( .A1(in_69bar), .A2(in_66bar), .ZN(n752bar);
  OR2_X1 U211 ( .A1(n966), .A2(n751), .ZN(n787) );
  AND2_X1 U211bar ( .A1(n966bar), .A2(n751bar), .ZN(n787bar);
  OR2_X1 U212 ( .A1(in[134]), .A2(n750), .ZN(n751) );
  AND2_X1 U212bar ( .A1(inbar[134]), .A2(n750bar), .ZN(n751bar);
  OR2_X1 U213 ( .A1(n749), .A2(n748), .ZN(n966) );
  AND2_X1 U213bar ( .A1(n749bar), .A2(n748bar), .ZN(n966bar);
  OR2_X1 U214 ( .A1(n747), .A2(n746), .ZN(n748) );
  AND2_X1 U214bar ( .A1(n747bar), .A2(n746bar), .ZN(n748bar);
  OR2_X1 U215 ( .A1(n745), .A2(n744), .ZN(n746) );
  AND2_X1 U215bar ( .A1(n745bar), .A2(n744bar), .ZN(n746bar);
  OR2_X1 U216 ( .A1(in[136]), .A2(in[121]), .ZN(n744) );
  AND2_X1 U216bar ( .A1(inbar[136]), .A2(inbar[121]), .ZN(n744bar);
  OR2_X1 U217 ( .A1(in[186]), .A2(in[174]), .ZN(n745) );
  AND2_X1 U217bar ( .A1(inbar[186]), .A2(inbar[174]), .ZN(n745bar);
  OR2_X1 U218 ( .A1(n743), .A2(n742), .ZN(n747) );
  AND2_X1 U218bar ( .A1(n743bar), .A2(n742bar), .ZN(n747bar);
  OR2_X1 U219 ( .A1(in[198]), .A2(in[197]), .ZN(n742) );
  AND2_X1 U219bar ( .A1(inbar[198]), .A2(inbar[197]), .ZN(n742bar);
  OR2_X1 U220 ( .A1(in[214]), .A2(in[199]), .ZN(n743) );
  AND2_X1 U220bar ( .A1(inbar[214]), .A2(inbar[199]), .ZN(n743bar);
  OR2_X1 U221 ( .A1(n741), .A2(n740), .ZN(n749) );
  AND2_X1 U221bar ( .A1(n741bar), .A2(n740bar), .ZN(n749bar);
  OR2_X1 U222 ( .A1(n739), .A2(n738), .ZN(n740) );
  AND2_X1 U222bar ( .A1(n739bar), .A2(n738bar), .ZN(n740bar);
  OR2_X1 U223 ( .A1(in[231]), .A2(in[220]), .ZN(n738) );
  AND2_X1 U223bar ( .A1(inbar[231]), .A2(inbar[220]), .ZN(n738bar);
  OR2_X1 U224 ( .A1(in_25), .A2(in[245]), .ZN(n739) );
  AND2_X1 U224bar ( .A1(in_25bar), .A2(inbar[245]), .ZN(n739bar);
  OR2_X1 U225 ( .A1(n737), .A2(n736), .ZN(n741) );
  AND2_X1 U225bar ( .A1(n737bar), .A2(n736bar), .ZN(n741bar);
  OR2_X1 U226 ( .A1(in_53), .A2(in_29), .ZN(n736) );
  AND2_X1 U226bar ( .A1(in_53bar), .A2(in_29bar), .ZN(n736bar);
  OR2_X1 U227 ( .A1(in_79), .A2(in_74), .ZN(n737) );
  AND2_X1 U227bar ( .A1(in_79bar), .A2(in_74bar), .ZN(n737bar);
  OR2_X1 U228 ( .A1(n735), .A2(n734), .ZN(n789) );
  AND2_X1 U228bar ( .A1(n735bar), .A2(n734bar), .ZN(n789bar);
  OR2_X1 U229 ( .A1(in[152]), .A2(in[140]), .ZN(n734) );
  AND2_X1 U229bar ( .A1(inbar[152]), .A2(inbar[140]), .ZN(n734bar);
  OR2_X1 U230 ( .A1(in[155]), .A2(n733), .ZN(n735) );
  AND2_X1 U230bar ( .A1(inbar[155]), .A2(n733bar), .ZN(n735bar);
  OR2_X1 U231 ( .A1(in[166]), .A2(in[165]), .ZN(n733) );
  AND2_X1 U231bar ( .A1(inbar[166]), .A2(inbar[165]), .ZN(n733bar);
  OR2_X1 U232 ( .A1(n732), .A2(n731), .ZN(n791) );
  AND2_X1 U232bar ( .A1(n732bar), .A2(n731bar), .ZN(n791bar);
  OR2_X1 U233 ( .A1(n730), .A2(n729), .ZN(n731) );
  AND2_X1 U233bar ( .A1(n730bar), .A2(n729bar), .ZN(n731bar);
  OR2_X1 U234 ( .A1(in[202]), .A2(in[185]), .ZN(n729) );
  AND2_X1 U234bar ( .A1(inbar[202]), .A2(inbar[185]), .ZN(n729bar);
  OR2_X1 U235 ( .A1(in[211]), .A2(n728), .ZN(n730) );
  AND2_X1 U235bar ( .A1(inbar[211]), .A2(n728bar), .ZN(n730bar);
  OR2_X1 U236 ( .A1(in[255]), .A2(in[253]), .ZN(n728) );
  AND2_X1 U236bar ( .A1(inbar[255]), .A2(inbar[253]), .ZN(n728bar);
  OR2_X1 U237 ( .A1(n727), .A2(n726), .ZN(n732) );
  AND2_X1 U237bar ( .A1(n727bar), .A2(n726bar), .ZN(n732bar);
  OR2_X1 U238 ( .A1(in_35), .A2(in_15), .ZN(n726) );
  AND2_X1 U238bar ( .A1(in_35bar), .A2(in_15bar), .ZN(n726bar);
  OR2_X1 U239 ( .A1(in_36), .A2(n725), .ZN(n727) );
  AND2_X1 U239bar ( .A1(in_36bar), .A2(n725bar), .ZN(n727bar);
  OR2_X1 U240 ( .A1(in_48), .A2(in_40), .ZN(n725) );
  AND2_X1 U240bar ( .A1(in_48bar), .A2(in_40bar), .ZN(n725bar);
  OR2_X1 U241 ( .A1(n724), .A2(n723), .ZN(out[1]) );
  AND2_X1 U241bar ( .A1(n724bar), .A2(n723bar), .ZN(outbar[1]);
  OR2_X1 U242 ( .A1(n722), .A2(n721), .ZN(n723) );
  AND2_X1 U242bar ( .A1(n722bar), .A2(n721bar), .ZN(n723bar);
  OR2_X1 U243 ( .A1(n720), .A2(n719), .ZN(n721) );
  AND2_X1 U243bar ( .A1(n720bar), .A2(n719bar), .ZN(n721bar);
  OR2_X1 U244 ( .A1(n921), .A2(n887), .ZN(n719) );
  AND2_X1 U244bar ( .A1(n921bar), .A2(n887bar), .ZN(n719bar);
  OR2_X1 U245 ( .A1(n718), .A2(n717), .ZN(n887) );
  AND2_X1 U245bar ( .A1(n718bar), .A2(n717bar), .ZN(n887bar);
  OR2_X1 U246 ( .A1(n716), .A2(n715), .ZN(n717) );
  AND2_X1 U246bar ( .A1(n716bar), .A2(n715bar), .ZN(n717bar);
  OR2_X1 U247 ( .A1(n714), .A2(n713), .ZN(n715) );
  AND2_X1 U247bar ( .A1(n714bar), .A2(n713bar), .ZN(n715bar);
  OR2_X1 U248 ( .A1(in[116]), .A2(in[110]), .ZN(n713) );
  AND2_X1 U248bar ( .A1(inbar[116]), .A2(inbar[110]), .ZN(n713bar);
  OR2_X1 U249 ( .A1(in[133]), .A2(in[130]), .ZN(n714) );
  AND2_X1 U249bar ( .A1(inbar[133]), .A2(inbar[130]), .ZN(n714bar);
  OR2_X1 U250 ( .A1(n712), .A2(n711), .ZN(n716) );
  AND2_X1 U250bar ( .A1(n712bar), .A2(n711bar), .ZN(n716bar);
  OR2_X1 U251 ( .A1(in[203]), .A2(in[135]), .ZN(n711) );
  AND2_X1 U251bar ( .A1(inbar[203]), .A2(inbar[135]), .ZN(n711bar);
  OR2_X1 U252 ( .A1(in[232]), .A2(in[223]), .ZN(n712) );
  AND2_X1 U252bar ( .A1(inbar[232]), .A2(inbar[223]), .ZN(n712bar);
  OR2_X1 U253 ( .A1(n710), .A2(n709), .ZN(n718) );
  AND2_X1 U253bar ( .A1(n710bar), .A2(n709bar), .ZN(n718bar);
  OR2_X1 U254 ( .A1(n708), .A2(n707), .ZN(n709) );
  AND2_X1 U254bar ( .A1(n708bar), .A2(n707bar), .ZN(n709bar);
  OR2_X1 U255 ( .A1(in[255]), .A2(in[233]), .ZN(n707) );
  AND2_X1 U255bar ( .A1(inbar[255]), .A2(inbar[233]), .ZN(n707bar);
  OR2_X1 U256 ( .A1(in_53), .A2(in_34), .ZN(n708) );
  AND2_X1 U256bar ( .A1(in_53bar), .A2(in_34bar), .ZN(n708bar);
  OR2_X1 U257 ( .A1(n706), .A2(n705), .ZN(n710) );
  AND2_X1 U257bar ( .A1(n706bar), .A2(n705bar), .ZN(n710bar);
  OR2_X1 U258 ( .A1(in_57), .A2(in_55), .ZN(n705) );
  AND2_X1 U258bar ( .A1(in_57bar), .A2(in_55bar), .ZN(n705bar);
  OR2_X1 U259 ( .A1(in_68), .A2(in_67), .ZN(n706) );
  AND2_X1 U259bar ( .A1(in_68bar), .A2(in_67bar), .ZN(n706bar);
  OR2_X1 U260 ( .A1(n704), .A2(n703), .ZN(n921) );
  AND2_X1 U260bar ( .A1(n704bar), .A2(n703bar), .ZN(n921bar);
  OR2_X1 U261 ( .A1(n702), .A2(n701), .ZN(n703) );
  AND2_X1 U261bar ( .A1(n702bar), .A2(n701bar), .ZN(n703bar);
  OR2_X1 U262 ( .A1(n700), .A2(n699), .ZN(n701) );
  AND2_X1 U262bar ( .A1(n700bar), .A2(n699bar), .ZN(n701bar);
  OR2_X1 U263 ( .A1(n944), .A2(n872), .ZN(n699) );
  AND2_X1 U263bar ( .A1(n944bar), .A2(n872bar), .ZN(n699bar);
  OR2_X1 U264 ( .A1(n698), .A2(n697), .ZN(n872) );
  AND2_X1 U264bar ( .A1(n698bar), .A2(n697bar), .ZN(n872bar);
  OR2_X1 U265 ( .A1(n696), .A2(n695), .ZN(n697) );
  AND2_X1 U265bar ( .A1(n696bar), .A2(n695bar), .ZN(n697bar);
  OR2_X1 U266 ( .A1(n694), .A2(n693), .ZN(n695) );
  AND2_X1 U266bar ( .A1(n694bar), .A2(n693bar), .ZN(n695bar);
  OR2_X1 U267 ( .A1(in[121]), .A2(in[102]), .ZN(n693) );
  AND2_X1 U267bar ( .A1(inbar[121]), .A2(inbar[102]), .ZN(n693bar);
  OR2_X1 U268 ( .A1(in[162]), .A2(in[161]), .ZN(n694) );
  AND2_X1 U268bar ( .A1(inbar[162]), .A2(inbar[161]), .ZN(n694bar);
  OR2_X1 U269 ( .A1(n692), .A2(n691), .ZN(n696) );
  AND2_X1 U269bar ( .A1(n692bar), .A2(n691bar), .ZN(n696bar);
  OR2_X1 U270 ( .A1(in[192]), .A2(in[178]), .ZN(n691) );
  AND2_X1 U270bar ( .A1(inbar[192]), .A2(inbar[178]), .ZN(n691bar);
  OR2_X1 U271 ( .A1(in[244]), .A2(in[209]), .ZN(n692) );
  AND2_X1 U271bar ( .A1(inbar[244]), .A2(inbar[209]), .ZN(n692bar);
  OR2_X1 U272 ( .A1(n690), .A2(n689), .ZN(n698) );
  AND2_X1 U272bar ( .A1(n690bar), .A2(n689bar), .ZN(n698bar);
  OR2_X1 U273 ( .A1(n688), .A2(n687), .ZN(n689) );
  AND2_X1 U273bar ( .A1(n688bar), .A2(n687bar), .ZN(n689bar);
  OR2_X1 U274 ( .A1(in[90]), .A2(in[254]), .ZN(n687) );
  AND2_X1 U274bar ( .A1(inbar[90]), .A2(inbar[254]), .ZN(n687bar);
  OR2_X1 U275 ( .A1(in_36), .A2(in_32), .ZN(n688) );
  AND2_X1 U275bar ( .A1(in_36bar), .A2(in_32bar), .ZN(n688bar);
  OR2_X1 U276 ( .A1(n686), .A2(n685), .ZN(n690) );
  AND2_X1 U276bar ( .A1(n686bar), .A2(n685bar), .ZN(n690bar);
  OR2_X1 U277 ( .A1(in_62), .A2(in_37), .ZN(n685) );
  AND2_X1 U277bar ( .A1(in_62bar), .A2(in_37bar), .ZN(n685bar);
  OR2_X1 U278 ( .A1(in_75), .A2(in_73), .ZN(n686) );
  AND2_X1 U278bar ( .A1(in_75bar), .A2(in_73bar), .ZN(n686bar);
  OR2_X1 U279 ( .A1(n684), .A2(n683), .ZN(n944) );
  AND2_X1 U279bar ( .A1(n684bar), .A2(n683bar), .ZN(n944bar);
  OR2_X1 U280 ( .A1(n682), .A2(n681), .ZN(n683) );
  AND2_X1 U280bar ( .A1(n682bar), .A2(n681bar), .ZN(n683bar);
  OR2_X1 U281 ( .A1(n680), .A2(n679), .ZN(n681) );
  AND2_X1 U281bar ( .A1(n680bar), .A2(n679bar), .ZN(n681bar);
  OR2_X1 U282 ( .A1(in[171]), .A2(in[153]), .ZN(n679) );
  AND2_X1 U282bar ( .A1(inbar[171]), .A2(inbar[153]), .ZN(n679bar);
  OR2_X1 U283 ( .A1(in[187]), .A2(in[176]), .ZN(n680) );
  AND2_X1 U283bar ( .A1(inbar[187]), .A2(inbar[176]), .ZN(n680bar);
  OR2_X1 U284 ( .A1(n678), .A2(n677), .ZN(n682) );
  AND2_X1 U284bar ( .A1(n678bar), .A2(n677bar), .ZN(n682bar);
  OR2_X1 U285 ( .A1(in[245]), .A2(in[211]), .ZN(n677) );
  AND2_X1 U285bar ( .A1(inbar[245]), .A2(inbar[211]), .ZN(n677bar);
  OR2_X1 U286 ( .A1(in[97]), .A2(in[88]), .ZN(n678) );
  AND2_X1 U286bar ( .A1(inbar[97]), .A2(inbar[88]), .ZN(n678bar);
  OR2_X1 U287 ( .A1(n676), .A2(n675), .ZN(n684) );
  AND2_X1 U287bar ( .A1(n676bar), .A2(n675bar), .ZN(n684bar);
  OR2_X1 U288 ( .A1(n674), .A2(n673), .ZN(n675) );
  AND2_X1 U288bar ( .A1(n674bar), .A2(n673bar), .ZN(n675bar);
  OR2_X1 U289 ( .A1(in_10), .A2(in_0), .ZN(n673) );
  AND2_X1 U289bar ( .A1(in_10bar), .A2(in_0bar), .ZN(n673bar);
  OR2_X1 U290 ( .A1(in_59), .A2(in_5), .ZN(n674) );
  AND2_X1 U290bar ( .A1(in_59bar), .A2(in_5bar), .ZN(n674bar);
  OR2_X1 U291 ( .A1(n672), .A2(n671), .ZN(n676) );
  AND2_X1 U291bar ( .A1(n672bar), .A2(n671bar), .ZN(n676bar);
  OR2_X1 U292 ( .A1(in_60), .A2(in_6), .ZN(n671) );
  AND2_X1 U292bar ( .A1(in_60bar), .A2(in_6bar), .ZN(n671bar);
  OR2_X1 U293 ( .A1(in_77), .A2(in_69), .ZN(n672) );
  AND2_X1 U293bar ( .A1(in_77bar), .A2(in_69bar), .ZN(n672bar);
  OR2_X1 U294 ( .A1(in[113]), .A2(n864), .ZN(n700) );
  AND2_X1 U294bar ( .A1(inbar[113]), .A2(n864bar), .ZN(n700bar);
  OR2_X1 U295 ( .A1(n670), .A2(n669), .ZN(n864) );
  AND2_X1 U295bar ( .A1(n670bar), .A2(n669bar), .ZN(n864bar);
  OR2_X1 U296 ( .A1(n668), .A2(n667), .ZN(n669) );
  AND2_X1 U296bar ( .A1(n668bar), .A2(n667bar), .ZN(n669bar);
  OR2_X1 U297 ( .A1(n666), .A2(n665), .ZN(n667) );
  AND2_X1 U297bar ( .A1(n666bar), .A2(n665bar), .ZN(n667bar);
  OR2_X1 U298 ( .A1(in[125]), .A2(in[107]), .ZN(n665) );
  AND2_X1 U298bar ( .A1(inbar[125]), .A2(inbar[107]), .ZN(n665bar);
  OR2_X1 U299 ( .A1(in[138]), .A2(in[126]), .ZN(n666) );
  AND2_X1 U299bar ( .A1(inbar[138]), .A2(inbar[126]), .ZN(n666bar);
  OR2_X1 U300 ( .A1(n664), .A2(n663), .ZN(n668) );
  AND2_X1 U300bar ( .A1(n664bar), .A2(n663bar), .ZN(n668bar);
  OR2_X1 U301 ( .A1(in[189]), .A2(in[143]), .ZN(n663) );
  AND2_X1 U301bar ( .A1(inbar[189]), .A2(inbar[143]), .ZN(n663bar);
  OR2_X1 U302 ( .A1(in[99]), .A2(in[214]), .ZN(n664) );
  AND2_X1 U302bar ( .A1(inbar[99]), .A2(inbar[214]), .ZN(n664bar);
  OR2_X1 U303 ( .A1(n662), .A2(n661), .ZN(n670) );
  AND2_X1 U303bar ( .A1(n662bar), .A2(n661bar), .ZN(n670bar);
  OR2_X1 U304 ( .A1(n660), .A2(n659), .ZN(n661) );
  AND2_X1 U304bar ( .A1(n660bar), .A2(n659bar), .ZN(n661bar);
  OR2_X1 U305 ( .A1(in_15), .A2(in_12), .ZN(n659) );
  AND2_X1 U305bar ( .A1(in_15bar), .A2(in_12bar), .ZN(n659bar);
  OR2_X1 U306 ( .A1(in_20), .A2(in_2), .ZN(n660) );
  AND2_X1 U306bar ( .A1(in_20bar), .A2(in_2bar), .ZN(n660bar);
  OR2_X1 U307 ( .A1(n658), .A2(n657), .ZN(n662) );
  AND2_X1 U307bar ( .A1(n658bar), .A2(n657bar), .ZN(n662bar);
  OR2_X1 U308 ( .A1(in_30), .A2(in_3), .ZN(n657) );
  AND2_X1 U308bar ( .A1(in_30bar), .A2(in_3bar), .ZN(n657bar);
  OR2_X1 U309 ( .A1(in_4), .A2(in_38), .ZN(n658) );
  AND2_X1 U309bar ( .A1(in_4bar), .A2(in_38bar), .ZN(n658bar);
  OR2_X1 U310 ( .A1(n656), .A2(n655), .ZN(n702) );
  AND2_X1 U310bar ( .A1(n656bar), .A2(n655bar), .ZN(n702bar);
  OR2_X1 U311 ( .A1(in[148]), .A2(in[137]), .ZN(n655) );
  AND2_X1 U311bar ( .A1(inbar[148]), .A2(inbar[137]), .ZN(n655bar);
  OR2_X1 U312 ( .A1(in[149]), .A2(n654), .ZN(n656) );
  AND2_X1 U312bar ( .A1(inbar[149]), .A2(n654bar), .ZN(n656bar);
  OR2_X1 U313 ( .A1(in[195]), .A2(in[190]), .ZN(n654) );
  AND2_X1 U313bar ( .A1(inbar[195]), .A2(inbar[190]), .ZN(n654bar);
  OR2_X1 U314 ( .A1(n653), .A2(n652), .ZN(n704) );
  AND2_X1 U314bar ( .A1(n653bar), .A2(n652bar), .ZN(n704bar);
  OR2_X1 U315 ( .A1(n651), .A2(n650), .ZN(n652) );
  AND2_X1 U315bar ( .A1(n651bar), .A2(n650bar), .ZN(n652bar);
  OR2_X1 U316 ( .A1(in[98]), .A2(in[197]), .ZN(n650) );
  AND2_X1 U316bar ( .A1(inbar[98]), .A2(inbar[197]), .ZN(n650bar);
  OR2_X1 U317 ( .A1(in_11), .A2(n649), .ZN(n651) );
  AND2_X1 U317bar ( .A1(in_11bar), .A2(n649bar), .ZN(n651bar);
  OR2_X1 U318 ( .A1(in_26), .A2(in_14), .ZN(n649) );
  AND2_X1 U318bar ( .A1(in_26bar), .A2(in_14bar), .ZN(n649bar);
  OR2_X1 U319 ( .A1(n648), .A2(n647), .ZN(n653) );
  AND2_X1 U319bar ( .A1(n648bar), .A2(n647bar), .ZN(n653bar);
  OR2_X1 U320 ( .A1(in_35), .A2(in_27), .ZN(n647) );
  AND2_X1 U320bar ( .A1(in_35bar), .A2(in_27bar), .ZN(n647bar);
  OR2_X1 U321 ( .A1(in_50), .A2(n646), .ZN(n648) );
  AND2_X1 U321bar ( .A1(in_50bar), .A2(n646bar), .ZN(n648bar);
  OR2_X1 U322 ( .A1(in_78), .A2(in_61), .ZN(n646) );
  AND2_X1 U322bar ( .A1(in_78bar), .A2(in_61bar), .ZN(n646bar);
  OR2_X1 U323 ( .A1(n942), .A2(n645), .ZN(n720) );
  AND2_X1 U323bar ( .A1(n942bar), .A2(n645bar), .ZN(n720bar);
  OR2_X1 U324 ( .A1(in[106]), .A2(n863), .ZN(n645) );
  AND2_X1 U324bar ( .A1(inbar[106]), .A2(n863bar), .ZN(n645bar);
  OR2_X1 U325 ( .A1(n644), .A2(n643), .ZN(n863) );
  AND2_X1 U325bar ( .A1(n644bar), .A2(n643bar), .ZN(n863bar);
  OR2_X1 U326 ( .A1(n642), .A2(n641), .ZN(n643) );
  AND2_X1 U326bar ( .A1(n642bar), .A2(n641bar), .ZN(n643bar);
  OR2_X1 U327 ( .A1(n640), .A2(n639), .ZN(n641) );
  AND2_X1 U327bar ( .A1(n640bar), .A2(n639bar), .ZN(n641bar);
  OR2_X1 U328 ( .A1(in[127]), .A2(in[122]), .ZN(n639) );
  AND2_X1 U328bar ( .A1(inbar[127]), .A2(inbar[122]), .ZN(n639bar);
  OR2_X1 U329 ( .A1(in[156]), .A2(in[132]), .ZN(n640) );
  AND2_X1 U329bar ( .A1(inbar[156]), .A2(inbar[132]), .ZN(n640bar);
  OR2_X1 U330 ( .A1(n638), .A2(n637), .ZN(n642) );
  AND2_X1 U330bar ( .A1(n638bar), .A2(n637bar), .ZN(n642bar);
  OR2_X1 U331 ( .A1(in[159]), .A2(in[157]), .ZN(n637) );
  AND2_X1 U331bar ( .A1(inbar[159]), .A2(inbar[157]), .ZN(n637bar);
  OR2_X1 U332 ( .A1(in[185]), .A2(in[169]), .ZN(n638) );
  AND2_X1 U332bar ( .A1(inbar[185]), .A2(inbar[169]), .ZN(n638bar);
  OR2_X1 U333 ( .A1(n636), .A2(n635), .ZN(n644) );
  AND2_X1 U333bar ( .A1(n636bar), .A2(n635bar), .ZN(n644bar);
  OR2_X1 U334 ( .A1(n634), .A2(n633), .ZN(n635) );
  AND2_X1 U334bar ( .A1(n634bar), .A2(n633bar), .ZN(n635bar);
  OR2_X1 U335 ( .A1(in[239]), .A2(in[218]), .ZN(n633) );
  AND2_X1 U335bar ( .A1(inbar[239]), .A2(inbar[218]), .ZN(n633bar);
  OR2_X1 U336 ( .A1(in_13), .A2(in[87]), .ZN(n634) );
  AND2_X1 U336bar ( .A1(in_13bar), .A2(inbar[87]), .ZN(n634bar);
  OR2_X1 U337 ( .A1(n632), .A2(n631), .ZN(n636) );
  AND2_X1 U337bar ( .A1(n632bar), .A2(n631bar), .ZN(n636bar);
  OR2_X1 U338 ( .A1(in_72), .A2(in_70), .ZN(n631) );
  AND2_X1 U338bar ( .A1(in_72bar), .A2(in_70bar), .ZN(n631bar);
  OR2_X1 U339 ( .A1(in_80), .A2(in_74), .ZN(n632) );
  AND2_X1 U339bar ( .A1(in_80bar), .A2(in_74bar), .ZN(n632bar);
  OR2_X1 U340 ( .A1(n630), .A2(n629), .ZN(n942) );
  AND2_X1 U340bar ( .A1(n630bar), .A2(n629bar), .ZN(n942bar);
  OR2_X1 U341 ( .A1(n628), .A2(n627), .ZN(n629) );
  AND2_X1 U341bar ( .A1(n628bar), .A2(n627bar), .ZN(n629bar);
  OR2_X1 U342 ( .A1(n626), .A2(n625), .ZN(n627) );
  AND2_X1 U342bar ( .A1(n626bar), .A2(n625bar), .ZN(n627bar);
  OR2_X1 U343 ( .A1(in[146]), .A2(in[100]), .ZN(n625) );
  AND2_X1 U343bar ( .A1(inbar[146]), .A2(inbar[100]), .ZN(n625bar);
  OR2_X1 U344 ( .A1(in[168]), .A2(in[152]), .ZN(n626) );
  AND2_X1 U344bar ( .A1(inbar[168]), .A2(inbar[152]), .ZN(n626bar);
  OR2_X1 U345 ( .A1(n624), .A2(n623), .ZN(n628) );
  AND2_X1 U345bar ( .A1(n624bar), .A2(n623bar), .ZN(n628bar);
  OR2_X1 U346 ( .A1(in[199]), .A2(in[182]), .ZN(n623) );
  AND2_X1 U346bar ( .A1(inbar[199]), .A2(inbar[182]), .ZN(n623bar);
  OR2_X1 U347 ( .A1(in[236]), .A2(in[204]), .ZN(n624) );
  AND2_X1 U347bar ( .A1(inbar[236]), .A2(inbar[204]), .ZN(n624bar);
  OR2_X1 U348 ( .A1(n622), .A2(n621), .ZN(n630) );
  AND2_X1 U348bar ( .A1(n622bar), .A2(n621bar), .ZN(n630bar);
  OR2_X1 U349 ( .A1(n620), .A2(n619), .ZN(n621) );
  AND2_X1 U349bar ( .A1(n620bar), .A2(n619bar), .ZN(n621bar);
  OR2_X1 U350 ( .A1(in[89]), .A2(in[246]), .ZN(n619) );
  AND2_X1 U350bar ( .A1(inbar[89]), .A2(inbar[246]), .ZN(n619bar);
  OR2_X1 U351 ( .A1(in[95]), .A2(in[92]), .ZN(n620) );
  AND2_X1 U351bar ( .A1(inbar[95]), .A2(inbar[92]), .ZN(n620bar);
  OR2_X1 U352 ( .A1(n618), .A2(n617), .ZN(n622) );
  AND2_X1 U352bar ( .A1(n618bar), .A2(n617bar), .ZN(n622bar);
  OR2_X1 U353 ( .A1(in_22), .A2(in_16), .ZN(n617) );
  AND2_X1 U353bar ( .A1(in_22bar), .A2(in_16bar), .ZN(n617bar);
  OR2_X1 U354 ( .A1(in_51), .A2(in_49), .ZN(n618) );
  AND2_X1 U354bar ( .A1(in_51bar), .A2(in_49bar), .ZN(n618bar);
  OR2_X1 U355 ( .A1(n616), .A2(n615), .ZN(n722) );
  AND2_X1 U355bar ( .A1(n616bar), .A2(n615bar), .ZN(n722bar);
  OR2_X1 U356 ( .A1(in[158]), .A2(in[115]), .ZN(n615) );
  AND2_X1 U356bar ( .A1(inbar[158]), .A2(inbar[115]), .ZN(n615bar);
  OR2_X1 U357 ( .A1(in[163]), .A2(n614), .ZN(n616) );
  AND2_X1 U357bar ( .A1(inbar[163]), .A2(n614bar), .ZN(n616bar);
  OR2_X1 U358 ( .A1(in[206]), .A2(in[165]), .ZN(n614) );
  AND2_X1 U358bar ( .A1(inbar[206]), .A2(inbar[165]), .ZN(n614bar);
  OR2_X1 U359 ( .A1(n613), .A2(n612), .ZN(n724) );
  AND2_X1 U359bar ( .A1(n613bar), .A2(n612bar), .ZN(n724bar);
  OR2_X1 U360 ( .A1(n611), .A2(n610), .ZN(n612) );
  AND2_X1 U360bar ( .A1(n611bar), .A2(n610bar), .ZN(n612bar);
  OR2_X1 U361 ( .A1(in[213]), .A2(in[207]), .ZN(n610) );
  AND2_X1 U361bar ( .A1(inbar[213]), .A2(inbar[207]), .ZN(n610bar);
  OR2_X1 U362 ( .A1(in[215]), .A2(n609), .ZN(n611) );
  AND2_X1 U362bar ( .A1(inbar[215]), .A2(n609bar), .ZN(n611bar);
  OR2_X1 U363 ( .A1(in[230]), .A2(in[220]), .ZN(n609) );
  AND2_X1 U363bar ( .A1(inbar[230]), .A2(inbar[220]), .ZN(n609bar);
  OR2_X1 U364 ( .A1(n608), .A2(n607), .ZN(n613) );
  AND2_X1 U364bar ( .A1(n608bar), .A2(n607bar), .ZN(n613bar);
  OR2_X1 U365 ( .A1(in[251]), .A2(in[234]), .ZN(n607) );
  AND2_X1 U365bar ( .A1(inbar[251]), .A2(inbar[234]), .ZN(n607bar);
  OR2_X1 U366 ( .A1(in_17), .A2(n606), .ZN(n608) );
  AND2_X1 U366bar ( .A1(in_17bar), .A2(n606bar), .ZN(n608bar);
  OR2_X1 U367 ( .A1(in_65), .A2(in_56), .ZN(n606) );
  AND2_X1 U367bar ( .A1(in_65bar), .A2(in_56bar), .ZN(n606bar);
  OR2_X1 U368 ( .A1(n605), .A2(n604), .ZN(out[0]) );
  AND2_X1 U368bar ( .A1(n605bar), .A2(n604bar), .ZN(outbar[0]);
  OR2_X1 U369 ( .A1(n603), .A2(n602), .ZN(n604) );
  AND2_X1 U369bar ( .A1(n603bar), .A2(n602bar), .ZN(n604bar);
  OR2_X1 U370 ( .A1(n601), .A2(n600), .ZN(n602) );
  AND2_X1 U370bar ( .A1(n601bar), .A2(n600bar), .ZN(n602bar);
  OR2_X1 U371 ( .A1(n820), .A2(n785), .ZN(n600) );
  AND2_X1 U371bar ( .A1(n820bar), .A2(n785bar), .ZN(n600bar);
  OR2_X1 U372 ( .A1(n599), .A2(n598), .ZN(n785) );
  AND2_X1 U372bar ( .A1(n599bar), .A2(n598bar), .ZN(n785bar);
  OR2_X1 U373 ( .A1(n597), .A2(n596), .ZN(n598) );
  AND2_X1 U373bar ( .A1(n597bar), .A2(n596bar), .ZN(n598bar);
  OR2_X1 U374 ( .A1(n595), .A2(n594), .ZN(n596) );
  AND2_X1 U374bar ( .A1(n595bar), .A2(n594bar), .ZN(n596bar);
  OR2_X1 U375 ( .A1(in[135]), .A2(in[104]), .ZN(n594) );
  AND2_X1 U375bar ( .A1(inbar[135]), .A2(inbar[104]), .ZN(n594bar);
  OR2_X1 U376 ( .A1(in[188]), .A2(in[178]), .ZN(n595) );
  AND2_X1 U376bar ( .A1(inbar[188]), .A2(inbar[178]), .ZN(n595bar);
  OR2_X1 U377 ( .A1(n593), .A2(n592), .ZN(n597) );
  AND2_X1 U377bar ( .A1(n593bar), .A2(n592bar), .ZN(n597bar);
  OR2_X1 U378 ( .A1(in[217]), .A2(in[194]), .ZN(n592) );
  AND2_X1 U378bar ( .A1(inbar[217]), .A2(inbar[194]), .ZN(n592bar);
  OR2_X1 U379 ( .A1(in[237]), .A2(in[218]), .ZN(n593) );
  AND2_X1 U379bar ( .A1(inbar[237]), .A2(inbar[218]), .ZN(n593bar);
  OR2_X1 U380 ( .A1(n591), .A2(n590), .ZN(n599) );
  AND2_X1 U380bar ( .A1(n591bar), .A2(n590bar), .ZN(n599bar);
  OR2_X1 U381 ( .A1(n589), .A2(n588), .ZN(n590) );
  AND2_X1 U381bar ( .A1(n589bar), .A2(n588bar), .ZN(n590bar);
  OR2_X1 U382 ( .A1(in_2), .A2(in_10), .ZN(n588) );
  AND2_X1 U382bar ( .A1(in_2bar), .A2(in_10bar), .ZN(n588bar);
  OR2_X1 U383 ( .A1(in_47), .A2(in_22), .ZN(n589) );
  AND2_X1 U383bar ( .A1(in_47bar), .A2(in_22bar), .ZN(n589bar);
  OR2_X1 U384 ( .A1(n587), .A2(n586), .ZN(n591) );
  AND2_X1 U384bar ( .A1(n587bar), .A2(n586bar), .ZN(n591bar);
  OR2_X1 U385 ( .A1(in_56), .A2(in_54), .ZN(n586) );
  AND2_X1 U385bar ( .A1(in_56bar), .A2(in_54bar), .ZN(n586bar);
  OR2_X1 U386 ( .A1(in_63), .A2(in_61), .ZN(n587) );
  AND2_X1 U386bar ( .A1(in_63bar), .A2(in_61bar), .ZN(n587bar);
  OR2_X1 U387 ( .A1(n585), .A2(n584), .ZN(n820) );
  AND2_X1 U387bar ( .A1(n585bar), .A2(n584bar), .ZN(n820bar);
  OR2_X1 U388 ( .A1(n583), .A2(n582), .ZN(n584) );
  AND2_X1 U388bar ( .A1(n583bar), .A2(n582bar), .ZN(n584bar);
  OR2_X1 U389 ( .A1(n581), .A2(n580), .ZN(n582) );
  AND2_X1 U389bar ( .A1(n581bar), .A2(n580bar), .ZN(n582bar);
  OR2_X1 U390 ( .A1(in[158]), .A2(in[142]), .ZN(n580) );
  AND2_X1 U390bar ( .A1(inbar[158]), .A2(inbar[142]), .ZN(n580bar);
  OR2_X1 U391 ( .A1(in[175]), .A2(in[164]), .ZN(n581) );
  AND2_X1 U391bar ( .A1(inbar[175]), .A2(inbar[164]), .ZN(n581bar);
  OR2_X1 U392 ( .A1(n579), .A2(n578), .ZN(n583) );
  AND2_X1 U392bar ( .A1(n579bar), .A2(n578bar), .ZN(n583bar);
  OR2_X1 U393 ( .A1(in[228]), .A2(in[204]), .ZN(n578) );
  AND2_X1 U393bar ( .A1(inbar[228]), .A2(inbar[204]), .ZN(n578bar);
  OR2_X1 U394 ( .A1(in[91]), .A2(in[87]), .ZN(n579) );
  AND2_X1 U394bar ( .A1(inbar[91]), .A2(inbar[87]), .ZN(n579bar);
  OR2_X1 U395 ( .A1(n577), .A2(n576), .ZN(n585) );
  AND2_X1 U395bar ( .A1(n577bar), .A2(n576bar), .ZN(n585bar);
  OR2_X1 U396 ( .A1(n575), .A2(n574), .ZN(n576) );
  AND2_X1 U396bar ( .A1(n575bar), .A2(n574bar), .ZN(n576bar);
  OR2_X1 U397 ( .A1(in_21), .A2(in_11), .ZN(n574) );
  AND2_X1 U397bar ( .A1(in_21bar), .A2(in_11bar), .ZN(n574bar);
  OR2_X1 U398 ( .A1(in_5), .A2(in_3), .ZN(n575) );
  AND2_X1 U398bar ( .A1(in_5bar), .A2(in_3bar), .ZN(n575bar);
  OR2_X1 U399 ( .A1(n573), .A2(n572), .ZN(n577) );
  AND2_X1 U399bar ( .A1(n573bar), .A2(n572bar), .ZN(n577bar);
  OR2_X1 U400 ( .A1(in_68), .A2(in_64), .ZN(n572) );
  AND2_X1 U400bar ( .A1(in_68bar), .A2(in_64bar), .ZN(n572bar);
  OR2_X1 U401 ( .A1(in_76), .A2(in_73), .ZN(n573) );
  AND2_X1 U401bar ( .A1(in_76bar), .A2(in_73bar), .ZN(n573bar);
  OR2_X1 U402 ( .A1(n778), .A2(n571), .ZN(n601) );
  AND2_X1 U402bar ( .A1(n778bar), .A2(n571bar), .ZN(n601bar);
  OR2_X1 U403 ( .A1(in[100]), .A2(n965), .ZN(n571) );
  AND2_X1 U403bar ( .A1(inbar[100]), .A2(n965bar), .ZN(n571bar);
  OR2_X1 U404 ( .A1(n570), .A2(n569), .ZN(n965) );
  AND2_X1 U404bar ( .A1(n570bar), .A2(n569bar), .ZN(n965bar);
  OR2_X1 U405 ( .A1(n568), .A2(n567), .ZN(n569) );
  AND2_X1 U405bar ( .A1(n568bar), .A2(n567bar), .ZN(n569bar);
  OR2_X1 U406 ( .A1(n566), .A2(n565), .ZN(n567) );
  AND2_X1 U406bar ( .A1(n566bar), .A2(n565bar), .ZN(n567bar);
  OR2_X1 U407 ( .A1(n817), .A2(n750), .ZN(n565) );
  AND2_X1 U407bar ( .A1(n817bar), .A2(n750bar), .ZN(n565bar);
  OR2_X1 U408 ( .A1(n564), .A2(n563), .ZN(n750) );
  AND2_X1 U408bar ( .A1(n564bar), .A2(n563bar), .ZN(n750bar);
  OR2_X1 U409 ( .A1(n562), .A2(n561), .ZN(n563) );
  AND2_X1 U409bar ( .A1(n562bar), .A2(n561bar), .ZN(n563bar);
  OR2_X1 U410 ( .A1(n560), .A2(n559), .ZN(n561) );
  AND2_X1 U410bar ( .A1(n560bar), .A2(n559bar), .ZN(n561bar);
  OR2_X1 U411 ( .A1(in[119]), .A2(in[103]), .ZN(n559) );
  AND2_X1 U411bar ( .A1(inbar[119]), .A2(inbar[103]), .ZN(n559bar);
  OR2_X1 U412 ( .A1(in[137]), .A2(in[133]), .ZN(n560) );
  AND2_X1 U412bar ( .A1(inbar[137]), .A2(inbar[133]), .ZN(n560bar);
  OR2_X1 U413 ( .A1(n558), .A2(n557), .ZN(n562) );
  AND2_X1 U413bar ( .A1(n558bar), .A2(n557bar), .ZN(n562bar);
  OR2_X1 U414 ( .A1(in[176]), .A2(in[173]), .ZN(n557) );
  AND2_X1 U414bar ( .A1(inbar[176]), .A2(inbar[173]), .ZN(n557bar);
  OR2_X1 U415 ( .A1(in[210]), .A2(in[181]), .ZN(n558) );
  AND2_X1 U415bar ( .A1(inbar[210]), .A2(inbar[181]), .ZN(n558bar);
  OR2_X1 U416 ( .A1(n556), .A2(n555), .ZN(n564) );
  AND2_X1 U416bar ( .A1(n556bar), .A2(n555bar), .ZN(n564bar);
  OR2_X1 U417 ( .A1(n554), .A2(n553), .ZN(n555) );
  AND2_X1 U417bar ( .A1(n554bar), .A2(n553bar), .ZN(n555bar);
  OR2_X1 U418 ( .A1(in_13), .A2(in[234]), .ZN(n553) );
  AND2_X1 U418bar ( .A1(in_13bar), .A2(inbar[234]), .ZN(n553bar);
  OR2_X1 U419 ( .A1(in_38), .A2(in_32), .ZN(n554) );
  AND2_X1 U419bar ( .A1(in_38bar), .A2(in_32bar), .ZN(n554bar);
  OR2_X1 U420 ( .A1(n552), .A2(n551), .ZN(n556) );
  AND2_X1 U420bar ( .A1(n552bar), .A2(n551bar), .ZN(n556bar);
  OR2_X1 U421 ( .A1(in_42), .A2(in_41), .ZN(n551) );
  AND2_X1 U421bar ( .A1(in_42bar), .A2(in_41bar), .ZN(n551bar);
  OR2_X1 U422 ( .A1(in_7), .A2(in_49), .ZN(n552) );
  AND2_X1 U422bar ( .A1(in_7bar), .A2(in_49bar), .ZN(n552bar);
  OR2_X1 U423 ( .A1(n550), .A2(n549), .ZN(n817) );
  AND2_X1 U423bar ( .A1(n550bar), .A2(n549bar), .ZN(n817bar);
  OR2_X1 U424 ( .A1(n548), .A2(n547), .ZN(n549) );
  AND2_X1 U424bar ( .A1(n548bar), .A2(n547bar), .ZN(n549bar);
  OR2_X1 U425 ( .A1(n546), .A2(n545), .ZN(n547) );
  AND2_X1 U425bar ( .A1(n546bar), .A2(n545bar), .ZN(n547bar);
  OR2_X1 U426 ( .A1(in[159]), .A2(in[105]), .ZN(n545) );
  AND2_X1 U426bar ( .A1(inbar[159]), .A2(inbar[105]), .ZN(n545bar);
  OR2_X1 U427 ( .A1(in[206]), .A2(in[183]), .ZN(n546) );
  AND2_X1 U427bar ( .A1(inbar[206]), .A2(inbar[183]), .ZN(n546bar);
  OR2_X1 U428 ( .A1(n544), .A2(n543), .ZN(n548) );
  AND2_X1 U428bar ( .A1(n544bar), .A2(n543bar), .ZN(n548bar);
  OR2_X1 U429 ( .A1(in[229]), .A2(in[219]), .ZN(n543) );
  AND2_X1 U429bar ( .A1(inbar[229]), .A2(inbar[219]), .ZN(n543bar);
  OR2_X1 U430 ( .A1(in[235]), .A2(in[232]), .ZN(n544) );
  AND2_X1 U430bar ( .A1(inbar[235]), .A2(inbar[232]), .ZN(n544bar);
  OR2_X1 U431 ( .A1(n542), .A2(n541), .ZN(n550) );
  AND2_X1 U431bar ( .A1(n542bar), .A2(n541bar), .ZN(n550bar);
  OR2_X1 U432 ( .A1(n540), .A2(n539), .ZN(n541) );
  AND2_X1 U432bar ( .A1(n540bar), .A2(n539bar), .ZN(n541bar);
  OR2_X1 U433 ( .A1(in[249]), .A2(in[242]), .ZN(n539) );
  AND2_X1 U433bar ( .A1(inbar[249]), .A2(inbar[242]), .ZN(n539bar);
  OR2_X1 U434 ( .A1(in[89]), .A2(in[254]), .ZN(n540) );
  AND2_X1 U434bar ( .A1(inbar[89]), .A2(inbar[254]), .ZN(n540bar);
  OR2_X1 U435 ( .A1(n538), .A2(n537), .ZN(n542) );
  AND2_X1 U435bar ( .A1(n538bar), .A2(n537bar), .ZN(n542bar);
  OR2_X1 U436 ( .A1(in_14), .A2(in[99]), .ZN(n537) );
  AND2_X1 U436bar ( .A1(in_14bar), .A2(inbar[99]), .ZN(n537bar);
  OR2_X1 U437 ( .A1(in_60), .A2(in_18), .ZN(n538) );
  AND2_X1 U437bar ( .A1(in_60bar), .A2(in_18bar), .ZN(n538bar);
  OR2_X1 U438 ( .A1(in[113]), .A2(n763), .ZN(n566) );
  AND2_X1 U438bar ( .A1(inbar[113]), .A2(n763bar), .ZN(n566bar);
  OR2_X1 U439 ( .A1(n536), .A2(n535), .ZN(n763) );
  AND2_X1 U439bar ( .A1(n536bar), .A2(n535bar), .ZN(n763bar);
  OR2_X1 U440 ( .A1(n534), .A2(n533), .ZN(n535) );
  AND2_X1 U440bar ( .A1(n534bar), .A2(n533bar), .ZN(n535bar);
  OR2_X1 U441 ( .A1(n532), .A2(n531), .ZN(n533) );
  AND2_X1 U441bar ( .A1(n532bar), .A2(n531bar), .ZN(n533bar);
  OR2_X1 U442 ( .A1(in[115]), .A2(in[110]), .ZN(n531) );
  AND2_X1 U442bar ( .A1(inbar[115]), .A2(inbar[110]), .ZN(n531bar);
  OR2_X1 U443 ( .A1(in[125]), .A2(in[117]), .ZN(n532) );
  AND2_X1 U443bar ( .A1(inbar[125]), .A2(inbar[117]), .ZN(n532bar);
  OR2_X1 U444 ( .A1(n530), .A2(n529), .ZN(n534) );
  AND2_X1 U444bar ( .A1(n530bar), .A2(n529bar), .ZN(n534bar);
  OR2_X1 U445 ( .A1(in[180]), .A2(in[128]), .ZN(n529) );
  AND2_X1 U445bar ( .A1(inbar[180]), .A2(inbar[128]), .ZN(n529bar);
  OR2_X1 U446 ( .A1(in[205]), .A2(in[201]), .ZN(n530) );
  AND2_X1 U446bar ( .A1(inbar[205]), .A2(inbar[201]), .ZN(n530bar);
  OR2_X1 U447 ( .A1(n528), .A2(n527), .ZN(n536) );
  AND2_X1 U447bar ( .A1(n528bar), .A2(n527bar), .ZN(n536bar);
  OR2_X1 U448 ( .A1(n526), .A2(n525), .ZN(n527) );
  AND2_X1 U448bar ( .A1(n526bar), .A2(n525bar), .ZN(n527bar);
  OR2_X1 U449 ( .A1(in[244]), .A2(in[239]), .ZN(n525) );
  AND2_X1 U449bar ( .A1(inbar[244]), .A2(inbar[239]), .ZN(n525bar);
  OR2_X1 U450 ( .A1(in[95]), .A2(in[83]), .ZN(n526) );
  AND2_X1 U450bar ( .A1(inbar[95]), .A2(inbar[83]), .ZN(n526bar);
  OR2_X1 U451 ( .A1(n524), .A2(n523), .ZN(n528) );
  AND2_X1 U451bar ( .A1(n524bar), .A2(n523bar), .ZN(n528bar);
  OR2_X1 U452 ( .A1(in_24), .A2(in[97]), .ZN(n523) );
  AND2_X1 U452bar ( .A1(in_24bar), .A2(inbar[97]), .ZN(n523bar);
  OR2_X1 U453 ( .A1(in_33), .A2(in_27), .ZN(n524) );
  AND2_X1 U453bar ( .A1(in_33bar), .A2(in_27bar), .ZN(n524bar);
  OR2_X1 U454 ( .A1(n522), .A2(n521), .ZN(n568) );
  AND2_X1 U454bar ( .A1(n522bar), .A2(n521bar), .ZN(n568bar);
  OR2_X1 U455 ( .A1(in[145]), .A2(in[126]), .ZN(n521) );
  AND2_X1 U455bar ( .A1(inbar[145]), .A2(inbar[126]), .ZN(n521bar);
  OR2_X1 U456 ( .A1(in[169]), .A2(n520), .ZN(n522) );
  AND2_X1 U456bar ( .A1(inbar[169]), .A2(n520bar), .ZN(n522bar);
  OR2_X1 U457 ( .A1(in[221]), .A2(in[172]), .ZN(n520) );
  AND2_X1 U457bar ( .A1(inbar[221]), .A2(inbar[172]), .ZN(n520bar);
  OR2_X1 U458 ( .A1(n519), .A2(n518), .ZN(n570) );
  AND2_X1 U458bar ( .A1(n519bar), .A2(n518bar), .ZN(n570bar);
  OR2_X1 U459 ( .A1(n517), .A2(n516), .ZN(n518) );
  AND2_X1 U459bar ( .A1(n517bar), .A2(n516bar), .ZN(n518bar);
  OR2_X1 U460 ( .A1(in[241]), .A2(in[224]), .ZN(n516) );
  AND2_X1 U460bar ( .A1(inbar[241]), .A2(inbar[224]), .ZN(n516bar);
  OR2_X1 U461 ( .A1(in[86]), .A2(n515), .ZN(n517) );
  AND2_X1 U461bar ( .A1(inbar[86]), .A2(n515bar), .ZN(n517bar);
  OR2_X1 U462 ( .A1(in_43), .A2(in_34), .ZN(n515) );
  AND2_X1 U462bar ( .A1(in_43bar), .A2(in_34bar), .ZN(n515bar);
  OR2_X1 U463 ( .A1(n514), .A2(n513), .ZN(n519) );
  AND2_X1 U463bar ( .A1(n514bar), .A2(n513bar), .ZN(n519bar);
  OR2_X1 U464 ( .A1(in_65), .A2(in_51), .ZN(n513) );
  AND2_X1 U464bar ( .A1(in_65bar), .A2(in_51bar), .ZN(n513bar);
  OR2_X1 U465 ( .A1(in_75), .A2(n512), .ZN(n514) );
  AND2_X1 U465bar ( .A1(in_75bar), .A2(n512bar), .ZN(n514bar);
  OR2_X1 U466 ( .A1(in_81), .A2(in_77), .ZN(n512) );
  AND2_X1 U466bar ( .A1(in_81bar), .A2(in_77bar), .ZN(n512bar);
  OR2_X1 U467 ( .A1(n511), .A2(n510), .ZN(n778) );
  AND2_X1 U467bar ( .A1(n511bar), .A2(n510bar), .ZN(n778bar);
  OR2_X1 U468 ( .A1(n509), .A2(n508), .ZN(n510) );
  AND2_X1 U468bar ( .A1(n509bar), .A2(n508bar), .ZN(n510bar);
  OR2_X1 U469 ( .A1(n507), .A2(n506), .ZN(n508) );
  AND2_X1 U469bar ( .A1(n507bar), .A2(n506bar), .ZN(n508bar);
  OR2_X1 U470 ( .A1(in[107]), .A2(in[101]), .ZN(n506) );
  AND2_X1 U470bar ( .A1(inbar[107]), .A2(inbar[101]), .ZN(n506bar);
  OR2_X1 U471 ( .A1(in[139]), .A2(in[132]), .ZN(n507) );
  AND2_X1 U471bar ( .A1(inbar[139]), .A2(inbar[132]), .ZN(n507bar);
  OR2_X1 U472 ( .A1(n505), .A2(n504), .ZN(n509) );
  AND2_X1 U472bar ( .A1(n505bar), .A2(n504bar), .ZN(n509bar);
  OR2_X1 U473 ( .A1(in[146]), .A2(in[141]), .ZN(n504) );
  AND2_X1 U473bar ( .A1(inbar[146]), .A2(inbar[141]), .ZN(n504bar);
  OR2_X1 U474 ( .A1(in[203]), .A2(in[179]), .ZN(n505) );
  AND2_X1 U474bar ( .A1(inbar[203]), .A2(inbar[179]), .ZN(n505bar);
  OR2_X1 U475 ( .A1(n503), .A2(n502), .ZN(n511) );
  AND2_X1 U475bar ( .A1(n503bar), .A2(n502bar), .ZN(n511bar);
  OR2_X1 U476 ( .A1(n501), .A2(n500), .ZN(n502) );
  AND2_X1 U476bar ( .A1(n501bar), .A2(n500bar), .ZN(n502bar);
  OR2_X1 U477 ( .A1(in[243]), .A2(in[222]), .ZN(n500) );
  AND2_X1 U477bar ( .A1(inbar[243]), .A2(inbar[222]), .ZN(n500bar);
  OR2_X1 U478 ( .A1(in[251]), .A2(in[250]), .ZN(n501) );
  AND2_X1 U478bar ( .A1(inbar[251]), .A2(inbar[250]), .ZN(n501bar);
  OR2_X1 U479 ( .A1(n499), .A2(n498), .ZN(n503) );
  AND2_X1 U479bar ( .A1(n499bar), .A2(n498bar), .ZN(n503bar);
  OR2_X1 U480 ( .A1(in_37), .A2(in_19), .ZN(n498) );
  AND2_X1 U480bar ( .A1(in_37bar), .A2(in_19bar), .ZN(n498bar);
  OR2_X1 U481 ( .A1(in_78), .A2(in_6), .ZN(n499) );
  AND2_X1 U481bar ( .A1(in_78bar), .A2(in_6bar), .ZN(n499bar);
  OR2_X1 U482 ( .A1(n497), .A2(n496), .ZN(n603) );
  AND2_X1 U482bar ( .A1(n497bar), .A2(n496bar), .ZN(n603bar);
  OR2_X1 U483 ( .A1(in[112]), .A2(in[102]), .ZN(n496) );
  AND2_X1 U483bar ( .A1(inbar[112]), .A2(inbar[102]), .ZN(n496bar);
  OR2_X1 U484 ( .A1(in[123]), .A2(n495), .ZN(n497) );
  AND2_X1 U484bar ( .A1(inbar[123]), .A2(n495bar), .ZN(n497bar);
  OR2_X1 U485 ( .A1(in[143]), .A2(in[130]), .ZN(n495) );
  AND2_X1 U485bar ( .A1(inbar[143]), .A2(inbar[130]), .ZN(n495bar);
  OR2_X1 U486 ( .A1(n494), .A2(n493), .ZN(n605) );
  AND2_X1 U486bar ( .A1(n494bar), .A2(n493bar), .ZN(n605bar);
  OR2_X1 U487 ( .A1(n492), .A2(n491), .ZN(n493) );
  AND2_X1 U487bar ( .A1(n492bar), .A2(n491bar), .ZN(n493bar);
  OR2_X1 U488 ( .A1(in[216]), .A2(in[213]), .ZN(n491) );
  AND2_X1 U488bar ( .A1(inbar[216]), .A2(inbar[213]), .ZN(n491bar);
  OR2_X1 U489 ( .A1(in[227]), .A2(n490), .ZN(n492) );
  AND2_X1 U489bar ( .A1(inbar[227]), .A2(n490bar), .ZN(n492bar);
  OR2_X1 U490 ( .A1(in_0), .A2(in[248]), .ZN(n490) );
  AND2_X1 U490bar ( .A1(in_0bar), .A2(inbar[248]), .ZN(n490bar);
  OR2_X1 U491 ( .A1(n489), .A2(n488), .ZN(n494) );
  AND2_X1 U491bar ( .A1(n489bar), .A2(n488bar), .ZN(n494bar);
  OR2_X1 U492 ( .A1(in_46), .A2(in_44), .ZN(n488) );
  AND2_X1 U492bar ( .A1(in_46bar), .A2(in_44bar), .ZN(n488bar);
  OR2_X1 U493 ( .A1(in_50), .A2(n487), .ZN(n489) );
  AND2_X1 U493bar ( .A1(in_50bar), .A2(n487bar), .ZN(n489bar);
  OR2_X1 U494 ( .A1(in_9), .A2(in_80), .ZN(n487) );
  AND2_X1 U494bar ( .A1(in_9bar), .A2(in_80bar), .ZN(n487bar);
endmodule




module sBox_7 ( in, out );
  input [7:0] in;
  //input_done

  output [7:0] out;
  //output_done

  wire   [255:0] decodeOut;
  //wire_done

  decode_7 dec ( .in(in), .out(decodeOut) );
  encode_7 enc ( .in(decodeOut), .out(out) );
endmodule


module CD2_29 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_30 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_31 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_32 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD4_15 ( a, b, y );
  input [3:0] a;
  input [3:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  //input_done

  output [15:0] y;
  reg [15:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]);
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]);
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]);
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]);
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]);
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]);
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]);
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]);
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]);
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]);
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]);
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]);
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]);
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]);
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]);
endmodule




module CD4_16 ( a, b, y );
  input [3:0] a;
  input [3:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  //input_done

  output [15:0] y;
  reg [15:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]);
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]);
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]);
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]);
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]);
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]);
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]);
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]);
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]);
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]);
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]);
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]);
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]);
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]);
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]);
endmodule




module CD16_8 ( a, b, y );
  input [15:0] a;
  input [15:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign abar[8] = ~a[8];
  assign abar[9] = ~a[9];
  assign abar[10] = ~a[10];
  assign abar[11] = ~a[11];
  assign abar[12] = ~a[12];
  assign abar[13] = ~a[13];
  assign abar[14] = ~a[14];
  assign abar[15] = ~a[15];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign bbar[8] = ~b[8];
  assign bbar[9] = ~b[9];
  assign bbar[10] = ~b[10];
  assign bbar[11] = ~b[11];
  assign bbar[12] = ~b[12];
  assign bbar[13] = ~b[13];
  assign bbar[14] = ~b[14];
  assign bbar[15] = ~b[15];
  //input_done

  output [255:0] y;
  reg [255:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[9]), .A2(a[0]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[9]), .A2(abar[0]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[3]), .A2(a[6]), .ZN(y[99]) );
  OR2_X1 U2bar ( .A1(bbar[3]), .A2(abar[6]), .ZN(ybar[99]);
  AND2_X1 U3 ( .A1(b[2]), .A2(a[6]), .ZN(y[98]) );
  OR2_X1 U3bar ( .A1(bbar[2]), .A2(abar[6]), .ZN(ybar[98]);
  AND2_X1 U4 ( .A1(b[1]), .A2(a[6]), .ZN(y[97]) );
  OR2_X1 U4bar ( .A1(bbar[1]), .A2(abar[6]), .ZN(ybar[97]);
  AND2_X1 U5 ( .A1(b[0]), .A2(a[6]), .ZN(y[96]) );
  OR2_X1 U5bar ( .A1(bbar[0]), .A2(abar[6]), .ZN(ybar[96]);
  AND2_X1 U6 ( .A1(b[15]), .A2(a[5]), .ZN(y[95]) );
  OR2_X1 U6bar ( .A1(bbar[15]), .A2(abar[5]), .ZN(ybar[95]);
  AND2_X1 U7 ( .A1(b[14]), .A2(a[5]), .ZN(y[94]) );
  OR2_X1 U7bar ( .A1(bbar[14]), .A2(abar[5]), .ZN(ybar[94]);
  AND2_X1 U8 ( .A1(b[13]), .A2(a[5]), .ZN(y[93]) );
  OR2_X1 U8bar ( .A1(bbar[13]), .A2(abar[5]), .ZN(ybar[93]);
  AND2_X1 U9 ( .A1(b[12]), .A2(a[5]), .ZN(y[92]) );
  OR2_X1 U9bar ( .A1(bbar[12]), .A2(abar[5]), .ZN(ybar[92]);
  AND2_X1 U10 ( .A1(b[11]), .A2(a[5]), .ZN(y[91]) );
  OR2_X1 U10bar ( .A1(bbar[11]), .A2(abar[5]), .ZN(ybar[91]);
  AND2_X1 U11 ( .A1(b[10]), .A2(a[5]), .ZN(y[90]) );
  OR2_X1 U11bar ( .A1(bbar[10]), .A2(abar[5]), .ZN(ybar[90]);
  AND2_X1 U12 ( .A1(b[8]), .A2(a[0]), .ZN(y[8]) );
  OR2_X1 U12bar ( .A1(bbar[8]), .A2(abar[0]), .ZN(ybar[8]);
  AND2_X1 U13 ( .A1(a[5]), .A2(b[9]), .ZN(y[89]) );
  OR2_X1 U13bar ( .A1(abar[5]), .A2(bbar[9]), .ZN(ybar[89]);
  AND2_X1 U14 ( .A1(b[8]), .A2(a[5]), .ZN(y[88]) );
  OR2_X1 U14bar ( .A1(bbar[8]), .A2(abar[5]), .ZN(ybar[88]);
  AND2_X1 U15 ( .A1(b[7]), .A2(a[5]), .ZN(y[87]) );
  OR2_X1 U15bar ( .A1(bbar[7]), .A2(abar[5]), .ZN(ybar[87]);
  AND2_X1 U16 ( .A1(b[6]), .A2(a[5]), .ZN(y[86]) );
  OR2_X1 U16bar ( .A1(bbar[6]), .A2(abar[5]), .ZN(ybar[86]);
  AND2_X1 U17 ( .A1(b[5]), .A2(a[5]), .ZN(y[85]) );
  OR2_X1 U17bar ( .A1(bbar[5]), .A2(abar[5]), .ZN(ybar[85]);
  AND2_X1 U18 ( .A1(b[4]), .A2(a[5]), .ZN(y[84]) );
  OR2_X1 U18bar ( .A1(bbar[4]), .A2(abar[5]), .ZN(ybar[84]);
  AND2_X1 U19 ( .A1(a[5]), .A2(b[3]), .ZN(y[83]) );
  OR2_X1 U19bar ( .A1(abar[5]), .A2(bbar[3]), .ZN(ybar[83]);
  AND2_X1 U20 ( .A1(a[5]), .A2(b[2]), .ZN(y[82]) );
  OR2_X1 U20bar ( .A1(abar[5]), .A2(bbar[2]), .ZN(ybar[82]);
  AND2_X1 U21 ( .A1(a[5]), .A2(b[1]), .ZN(y[81]) );
  OR2_X1 U21bar ( .A1(abar[5]), .A2(bbar[1]), .ZN(ybar[81]);
  AND2_X1 U22 ( .A1(a[5]), .A2(b[0]), .ZN(y[80]) );
  OR2_X1 U22bar ( .A1(abar[5]), .A2(bbar[0]), .ZN(ybar[80]);
  AND2_X1 U23 ( .A1(b[7]), .A2(a[0]), .ZN(y[7]) );
  OR2_X1 U23bar ( .A1(bbar[7]), .A2(abar[0]), .ZN(ybar[7]);
  AND2_X1 U24 ( .A1(a[4]), .A2(b[15]), .ZN(y[79]) );
  OR2_X1 U24bar ( .A1(abar[4]), .A2(bbar[15]), .ZN(ybar[79]);
  AND2_X1 U25 ( .A1(a[4]), .A2(b[14]), .ZN(y[78]) );
  OR2_X1 U25bar ( .A1(abar[4]), .A2(bbar[14]), .ZN(ybar[78]);
  AND2_X1 U26 ( .A1(a[4]), .A2(b[13]), .ZN(y[77]) );
  OR2_X1 U26bar ( .A1(abar[4]), .A2(bbar[13]), .ZN(ybar[77]);
  AND2_X1 U27 ( .A1(a[4]), .A2(b[12]), .ZN(y[76]) );
  OR2_X1 U27bar ( .A1(abar[4]), .A2(bbar[12]), .ZN(ybar[76]);
  AND2_X1 U28 ( .A1(a[4]), .A2(b[11]), .ZN(y[75]) );
  OR2_X1 U28bar ( .A1(abar[4]), .A2(bbar[11]), .ZN(ybar[75]);
  AND2_X1 U29 ( .A1(a[4]), .A2(b[10]), .ZN(y[74]) );
  OR2_X1 U29bar ( .A1(abar[4]), .A2(bbar[10]), .ZN(ybar[74]);
  AND2_X1 U30 ( .A1(a[4]), .A2(b[9]), .ZN(y[73]) );
  OR2_X1 U30bar ( .A1(abar[4]), .A2(bbar[9]), .ZN(ybar[73]);
  AND2_X1 U31 ( .A1(a[4]), .A2(b[8]), .ZN(y[72]) );
  OR2_X1 U31bar ( .A1(abar[4]), .A2(bbar[8]), .ZN(ybar[72]);
  AND2_X1 U32 ( .A1(a[4]), .A2(b[7]), .ZN(y[71]) );
  OR2_X1 U32bar ( .A1(abar[4]), .A2(bbar[7]), .ZN(ybar[71]);
  AND2_X1 U33 ( .A1(a[4]), .A2(b[6]), .ZN(y[70]) );
  OR2_X1 U33bar ( .A1(abar[4]), .A2(bbar[6]), .ZN(ybar[70]);
  AND2_X1 U34 ( .A1(b[6]), .A2(a[0]), .ZN(y[6]) );
  OR2_X1 U34bar ( .A1(bbar[6]), .A2(abar[0]), .ZN(ybar[6]);
  AND2_X1 U35 ( .A1(a[4]), .A2(b[5]), .ZN(y[69]) );
  OR2_X1 U35bar ( .A1(abar[4]), .A2(bbar[5]), .ZN(ybar[69]);
  AND2_X1 U36 ( .A1(a[4]), .A2(b[4]), .ZN(y[68]) );
  OR2_X1 U36bar ( .A1(abar[4]), .A2(bbar[4]), .ZN(ybar[68]);
  AND2_X1 U37 ( .A1(a[4]), .A2(b[3]), .ZN(y[67]) );
  OR2_X1 U37bar ( .A1(abar[4]), .A2(bbar[3]), .ZN(ybar[67]);
  AND2_X1 U38 ( .A1(a[4]), .A2(b[2]), .ZN(y[66]) );
  OR2_X1 U38bar ( .A1(abar[4]), .A2(bbar[2]), .ZN(ybar[66]);
  AND2_X1 U39 ( .A1(a[4]), .A2(b[1]), .ZN(y[65]) );
  OR2_X1 U39bar ( .A1(abar[4]), .A2(bbar[1]), .ZN(ybar[65]);
  AND2_X1 U40 ( .A1(a[4]), .A2(b[0]), .ZN(y[64]) );
  OR2_X1 U40bar ( .A1(abar[4]), .A2(bbar[0]), .ZN(ybar[64]);
  AND2_X1 U41 ( .A1(a[3]), .A2(b[15]), .ZN(y[63]) );
  OR2_X1 U41bar ( .A1(abar[3]), .A2(bbar[15]), .ZN(ybar[63]);
  AND2_X1 U42 ( .A1(a[3]), .A2(b[14]), .ZN(y[62]) );
  OR2_X1 U42bar ( .A1(abar[3]), .A2(bbar[14]), .ZN(ybar[62]);
  AND2_X1 U43 ( .A1(a[3]), .A2(b[13]), .ZN(y[61]) );
  OR2_X1 U43bar ( .A1(abar[3]), .A2(bbar[13]), .ZN(ybar[61]);
  AND2_X1 U44 ( .A1(a[3]), .A2(b[12]), .ZN(y[60]) );
  OR2_X1 U44bar ( .A1(abar[3]), .A2(bbar[12]), .ZN(ybar[60]);
  AND2_X1 U45 ( .A1(b[5]), .A2(a[0]), .ZN(y[5]) );
  OR2_X1 U45bar ( .A1(bbar[5]), .A2(abar[0]), .ZN(ybar[5]);
  AND2_X1 U46 ( .A1(a[3]), .A2(b[11]), .ZN(y[59]) );
  OR2_X1 U46bar ( .A1(abar[3]), .A2(bbar[11]), .ZN(ybar[59]);
  AND2_X1 U47 ( .A1(a[3]), .A2(b[10]), .ZN(y[58]) );
  OR2_X1 U47bar ( .A1(abar[3]), .A2(bbar[10]), .ZN(ybar[58]);
  AND2_X1 U48 ( .A1(a[3]), .A2(b[9]), .ZN(y[57]) );
  OR2_X1 U48bar ( .A1(abar[3]), .A2(bbar[9]), .ZN(ybar[57]);
  AND2_X1 U49 ( .A1(a[3]), .A2(b[8]), .ZN(y[56]) );
  OR2_X1 U49bar ( .A1(abar[3]), .A2(bbar[8]), .ZN(ybar[56]);
  AND2_X1 U50 ( .A1(a[3]), .A2(b[7]), .ZN(y[55]) );
  OR2_X1 U50bar ( .A1(abar[3]), .A2(bbar[7]), .ZN(ybar[55]);
  AND2_X1 U51 ( .A1(a[3]), .A2(b[6]), .ZN(y[54]) );
  OR2_X1 U51bar ( .A1(abar[3]), .A2(bbar[6]), .ZN(ybar[54]);
  AND2_X1 U52 ( .A1(a[3]), .A2(b[5]), .ZN(y[53]) );
  OR2_X1 U52bar ( .A1(abar[3]), .A2(bbar[5]), .ZN(ybar[53]);
  AND2_X1 U53 ( .A1(a[3]), .A2(b[4]), .ZN(y[52]) );
  OR2_X1 U53bar ( .A1(abar[3]), .A2(bbar[4]), .ZN(ybar[52]);
  AND2_X1 U54 ( .A1(a[3]), .A2(b[3]), .ZN(y[51]) );
  OR2_X1 U54bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[51]);
  AND2_X1 U55 ( .A1(a[3]), .A2(b[2]), .ZN(y[50]) );
  OR2_X1 U55bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[50]);
  AND2_X1 U56 ( .A1(b[4]), .A2(a[0]), .ZN(y[4]) );
  OR2_X1 U56bar ( .A1(bbar[4]), .A2(abar[0]), .ZN(ybar[4]);
  AND2_X1 U57 ( .A1(a[3]), .A2(b[1]), .ZN(y[49]) );
  OR2_X1 U57bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[49]);
  AND2_X1 U58 ( .A1(a[3]), .A2(b[0]), .ZN(y[48]) );
  OR2_X1 U58bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[48]);
  AND2_X1 U59 ( .A1(a[2]), .A2(b[15]), .ZN(y[47]) );
  OR2_X1 U59bar ( .A1(abar[2]), .A2(bbar[15]), .ZN(ybar[47]);
  AND2_X1 U60 ( .A1(a[2]), .A2(b[14]), .ZN(y[46]) );
  OR2_X1 U60bar ( .A1(abar[2]), .A2(bbar[14]), .ZN(ybar[46]);
  AND2_X1 U61 ( .A1(a[2]), .A2(b[13]), .ZN(y[45]) );
  OR2_X1 U61bar ( .A1(abar[2]), .A2(bbar[13]), .ZN(ybar[45]);
  AND2_X1 U62 ( .A1(a[2]), .A2(b[12]), .ZN(y[44]) );
  OR2_X1 U62bar ( .A1(abar[2]), .A2(bbar[12]), .ZN(ybar[44]);
  AND2_X1 U63 ( .A1(a[2]), .A2(b[11]), .ZN(y[43]) );
  OR2_X1 U63bar ( .A1(abar[2]), .A2(bbar[11]), .ZN(ybar[43]);
  AND2_X1 U64 ( .A1(a[2]), .A2(b[10]), .ZN(y[42]) );
  OR2_X1 U64bar ( .A1(abar[2]), .A2(bbar[10]), .ZN(ybar[42]);
  AND2_X1 U65 ( .A1(a[2]), .A2(b[9]), .ZN(y[41]) );
  OR2_X1 U65bar ( .A1(abar[2]), .A2(bbar[9]), .ZN(ybar[41]);
  AND2_X1 U66 ( .A1(a[2]), .A2(b[8]), .ZN(y[40]) );
  OR2_X1 U66bar ( .A1(abar[2]), .A2(bbar[8]), .ZN(ybar[40]);
  AND2_X1 U67 ( .A1(b[3]), .A2(a[0]), .ZN(y[3]) );
  OR2_X1 U67bar ( .A1(bbar[3]), .A2(abar[0]), .ZN(ybar[3]);
  AND2_X1 U68 ( .A1(a[2]), .A2(b[7]), .ZN(y[39]) );
  OR2_X1 U68bar ( .A1(abar[2]), .A2(bbar[7]), .ZN(ybar[39]);
  AND2_X1 U69 ( .A1(a[2]), .A2(b[6]), .ZN(y[38]) );
  OR2_X1 U69bar ( .A1(abar[2]), .A2(bbar[6]), .ZN(ybar[38]);
  AND2_X1 U70 ( .A1(a[2]), .A2(b[5]), .ZN(y[37]) );
  OR2_X1 U70bar ( .A1(abar[2]), .A2(bbar[5]), .ZN(ybar[37]);
  AND2_X1 U71 ( .A1(a[2]), .A2(b[4]), .ZN(y[36]) );
  OR2_X1 U71bar ( .A1(abar[2]), .A2(bbar[4]), .ZN(ybar[36]);
  AND2_X1 U72 ( .A1(a[2]), .A2(b[3]), .ZN(y[35]) );
  OR2_X1 U72bar ( .A1(abar[2]), .A2(bbar[3]), .ZN(ybar[35]);
  AND2_X1 U73 ( .A1(a[2]), .A2(b[2]), .ZN(y[34]) );
  OR2_X1 U73bar ( .A1(abar[2]), .A2(bbar[2]), .ZN(ybar[34]);
  AND2_X1 U74 ( .A1(a[2]), .A2(b[1]), .ZN(y[33]) );
  OR2_X1 U74bar ( .A1(abar[2]), .A2(bbar[1]), .ZN(ybar[33]);
  AND2_X1 U75 ( .A1(a[2]), .A2(b[0]), .ZN(y[32]) );
  OR2_X1 U75bar ( .A1(abar[2]), .A2(bbar[0]), .ZN(ybar[32]);
  AND2_X1 U76 ( .A1(a[1]), .A2(b[15]), .ZN(y[31]) );
  OR2_X1 U76bar ( .A1(abar[1]), .A2(bbar[15]), .ZN(ybar[31]);
  AND2_X1 U77 ( .A1(a[1]), .A2(b[14]), .ZN(y[30]) );
  OR2_X1 U77bar ( .A1(abar[1]), .A2(bbar[14]), .ZN(ybar[30]);
  AND2_X1 U78 ( .A1(b[2]), .A2(a[0]), .ZN(y[2]) );
  OR2_X1 U78bar ( .A1(bbar[2]), .A2(abar[0]), .ZN(ybar[2]);
  AND2_X1 U79 ( .A1(a[1]), .A2(b[13]), .ZN(y[29]) );
  OR2_X1 U79bar ( .A1(abar[1]), .A2(bbar[13]), .ZN(ybar[29]);
  AND2_X1 U80 ( .A1(a[1]), .A2(b[12]), .ZN(y[28]) );
  OR2_X1 U80bar ( .A1(abar[1]), .A2(bbar[12]), .ZN(ybar[28]);
  AND2_X1 U81 ( .A1(a[1]), .A2(b[11]), .ZN(y[27]) );
  OR2_X1 U81bar ( .A1(abar[1]), .A2(bbar[11]), .ZN(ybar[27]);
  AND2_X1 U82 ( .A1(a[1]), .A2(b[10]), .ZN(y[26]) );
  OR2_X1 U82bar ( .A1(abar[1]), .A2(bbar[10]), .ZN(ybar[26]);
  AND2_X1 U83 ( .A1(a[1]), .A2(b[9]), .ZN(y[25]) );
  OR2_X1 U83bar ( .A1(abar[1]), .A2(bbar[9]), .ZN(ybar[25]);
  AND2_X1 U84 ( .A1(a[15]), .A2(b[15]), .ZN(y[255]) );
  OR2_X1 U84bar ( .A1(abar[15]), .A2(bbar[15]), .ZN(ybar[255]);
  AND2_X1 U85 ( .A1(a[15]), .A2(b[14]), .ZN(y[254]) );
  OR2_X1 U85bar ( .A1(abar[15]), .A2(bbar[14]), .ZN(ybar[254]);
  AND2_X1 U86 ( .A1(a[15]), .A2(b[13]), .ZN(y[253]) );
  OR2_X1 U86bar ( .A1(abar[15]), .A2(bbar[13]), .ZN(ybar[253]);
  AND2_X1 U87 ( .A1(a[15]), .A2(b[12]), .ZN(y[252]) );
  OR2_X1 U87bar ( .A1(abar[15]), .A2(bbar[12]), .ZN(ybar[252]);
  AND2_X1 U88 ( .A1(a[15]), .A2(b[11]), .ZN(y[251]) );
  OR2_X1 U88bar ( .A1(abar[15]), .A2(bbar[11]), .ZN(ybar[251]);
  AND2_X1 U89 ( .A1(a[15]), .A2(b[10]), .ZN(y[250]) );
  OR2_X1 U89bar ( .A1(abar[15]), .A2(bbar[10]), .ZN(ybar[250]);
  AND2_X1 U90 ( .A1(a[1]), .A2(b[8]), .ZN(y[24]) );
  OR2_X1 U90bar ( .A1(abar[1]), .A2(bbar[8]), .ZN(ybar[24]);
  AND2_X1 U91 ( .A1(a[15]), .A2(b[9]), .ZN(y[249]) );
  OR2_X1 U91bar ( .A1(abar[15]), .A2(bbar[9]), .ZN(ybar[249]);
  AND2_X1 U92 ( .A1(a[15]), .A2(b[8]), .ZN(y[248]) );
  OR2_X1 U92bar ( .A1(abar[15]), .A2(bbar[8]), .ZN(ybar[248]);
  AND2_X1 U93 ( .A1(a[15]), .A2(b[7]), .ZN(y[247]) );
  OR2_X1 U93bar ( .A1(abar[15]), .A2(bbar[7]), .ZN(ybar[247]);
  AND2_X1 U94 ( .A1(a[15]), .A2(b[6]), .ZN(y[246]) );
  OR2_X1 U94bar ( .A1(abar[15]), .A2(bbar[6]), .ZN(ybar[246]);
  AND2_X1 U95 ( .A1(a[15]), .A2(b[5]), .ZN(y[245]) );
  OR2_X1 U95bar ( .A1(abar[15]), .A2(bbar[5]), .ZN(ybar[245]);
  AND2_X1 U96 ( .A1(a[15]), .A2(b[4]), .ZN(y[244]) );
  OR2_X1 U96bar ( .A1(abar[15]), .A2(bbar[4]), .ZN(ybar[244]);
  AND2_X1 U97 ( .A1(a[15]), .A2(b[3]), .ZN(y[243]) );
  OR2_X1 U97bar ( .A1(abar[15]), .A2(bbar[3]), .ZN(ybar[243]);
  AND2_X1 U98 ( .A1(a[15]), .A2(b[2]), .ZN(y[242]) );
  OR2_X1 U98bar ( .A1(abar[15]), .A2(bbar[2]), .ZN(ybar[242]);
  AND2_X1 U99 ( .A1(a[15]), .A2(b[1]), .ZN(y[241]) );
  OR2_X1 U99bar ( .A1(abar[15]), .A2(bbar[1]), .ZN(ybar[241]);
  AND2_X1 U100 ( .A1(a[15]), .A2(b[0]), .ZN(y[240]) );
  OR2_X1 U100bar ( .A1(abar[15]), .A2(bbar[0]), .ZN(ybar[240]);
  AND2_X1 U101 ( .A1(a[1]), .A2(b[7]), .ZN(y[23]) );
  OR2_X1 U101bar ( .A1(abar[1]), .A2(bbar[7]), .ZN(ybar[23]);
  AND2_X1 U102 ( .A1(a[14]), .A2(b[15]), .ZN(y[239]) );
  OR2_X1 U102bar ( .A1(abar[14]), .A2(bbar[15]), .ZN(ybar[239]);
  AND2_X1 U103 ( .A1(a[14]), .A2(b[14]), .ZN(y[238]) );
  OR2_X1 U103bar ( .A1(abar[14]), .A2(bbar[14]), .ZN(ybar[238]);
  AND2_X1 U104 ( .A1(a[14]), .A2(b[13]), .ZN(y[237]) );
  OR2_X1 U104bar ( .A1(abar[14]), .A2(bbar[13]), .ZN(ybar[237]);
  AND2_X1 U105 ( .A1(a[14]), .A2(b[12]), .ZN(y[236]) );
  OR2_X1 U105bar ( .A1(abar[14]), .A2(bbar[12]), .ZN(ybar[236]);
  AND2_X1 U106 ( .A1(a[14]), .A2(b[11]), .ZN(y[235]) );
  OR2_X1 U106bar ( .A1(abar[14]), .A2(bbar[11]), .ZN(ybar[235]);
  AND2_X1 U107 ( .A1(a[14]), .A2(b[10]), .ZN(y[234]) );
  OR2_X1 U107bar ( .A1(abar[14]), .A2(bbar[10]), .ZN(ybar[234]);
  AND2_X1 U108 ( .A1(a[14]), .A2(b[9]), .ZN(y[233]) );
  OR2_X1 U108bar ( .A1(abar[14]), .A2(bbar[9]), .ZN(ybar[233]);
  AND2_X1 U109 ( .A1(a[14]), .A2(b[8]), .ZN(y[232]) );
  OR2_X1 U109bar ( .A1(abar[14]), .A2(bbar[8]), .ZN(ybar[232]);
  AND2_X1 U110 ( .A1(a[14]), .A2(b[7]), .ZN(y[231]) );
  OR2_X1 U110bar ( .A1(abar[14]), .A2(bbar[7]), .ZN(ybar[231]);
  AND2_X1 U111 ( .A1(a[14]), .A2(b[6]), .ZN(y[230]) );
  OR2_X1 U111bar ( .A1(abar[14]), .A2(bbar[6]), .ZN(ybar[230]);
  AND2_X1 U112 ( .A1(a[1]), .A2(b[6]), .ZN(y[22]) );
  OR2_X1 U112bar ( .A1(abar[1]), .A2(bbar[6]), .ZN(ybar[22]);
  AND2_X1 U113 ( .A1(a[14]), .A2(b[5]), .ZN(y[229]) );
  OR2_X1 U113bar ( .A1(abar[14]), .A2(bbar[5]), .ZN(ybar[229]);
  AND2_X1 U114 ( .A1(a[14]), .A2(b[4]), .ZN(y[228]) );
  OR2_X1 U114bar ( .A1(abar[14]), .A2(bbar[4]), .ZN(ybar[228]);
  AND2_X1 U115 ( .A1(a[14]), .A2(b[3]), .ZN(y[227]) );
  OR2_X1 U115bar ( .A1(abar[14]), .A2(bbar[3]), .ZN(ybar[227]);
  AND2_X1 U116 ( .A1(a[14]), .A2(b[2]), .ZN(y[226]) );
  OR2_X1 U116bar ( .A1(abar[14]), .A2(bbar[2]), .ZN(ybar[226]);
  AND2_X1 U117 ( .A1(a[14]), .A2(b[1]), .ZN(y[225]) );
  OR2_X1 U117bar ( .A1(abar[14]), .A2(bbar[1]), .ZN(ybar[225]);
  AND2_X1 U118 ( .A1(a[14]), .A2(b[0]), .ZN(y[224]) );
  OR2_X1 U118bar ( .A1(abar[14]), .A2(bbar[0]), .ZN(ybar[224]);
  AND2_X1 U119 ( .A1(a[13]), .A2(b[15]), .ZN(y[223]) );
  OR2_X1 U119bar ( .A1(abar[13]), .A2(bbar[15]), .ZN(ybar[223]);
  AND2_X1 U120 ( .A1(a[13]), .A2(b[14]), .ZN(y[222]) );
  OR2_X1 U120bar ( .A1(abar[13]), .A2(bbar[14]), .ZN(ybar[222]);
  AND2_X1 U121 ( .A1(a[13]), .A2(b[13]), .ZN(y[221]) );
  OR2_X1 U121bar ( .A1(abar[13]), .A2(bbar[13]), .ZN(ybar[221]);
  AND2_X1 U122 ( .A1(a[13]), .A2(b[12]), .ZN(y[220]) );
  OR2_X1 U122bar ( .A1(abar[13]), .A2(bbar[12]), .ZN(ybar[220]);
  AND2_X1 U123 ( .A1(a[1]), .A2(b[5]), .ZN(y[21]) );
  OR2_X1 U123bar ( .A1(abar[1]), .A2(bbar[5]), .ZN(ybar[21]);
  AND2_X1 U124 ( .A1(a[13]), .A2(b[11]), .ZN(y[219]) );
  OR2_X1 U124bar ( .A1(abar[13]), .A2(bbar[11]), .ZN(ybar[219]);
  AND2_X1 U125 ( .A1(a[13]), .A2(b[10]), .ZN(y[218]) );
  OR2_X1 U125bar ( .A1(abar[13]), .A2(bbar[10]), .ZN(ybar[218]);
  AND2_X1 U126 ( .A1(a[13]), .A2(b[9]), .ZN(y[217]) );
  OR2_X1 U126bar ( .A1(abar[13]), .A2(bbar[9]), .ZN(ybar[217]);
  AND2_X1 U127 ( .A1(a[13]), .A2(b[8]), .ZN(y[216]) );
  OR2_X1 U127bar ( .A1(abar[13]), .A2(bbar[8]), .ZN(ybar[216]);
  AND2_X1 U128 ( .A1(a[13]), .A2(b[7]), .ZN(y[215]) );
  OR2_X1 U128bar ( .A1(abar[13]), .A2(bbar[7]), .ZN(ybar[215]);
  AND2_X1 U129 ( .A1(a[13]), .A2(b[6]), .ZN(y[214]) );
  OR2_X1 U129bar ( .A1(abar[13]), .A2(bbar[6]), .ZN(ybar[214]);
  AND2_X1 U130 ( .A1(a[13]), .A2(b[5]), .ZN(y[213]) );
  OR2_X1 U130bar ( .A1(abar[13]), .A2(bbar[5]), .ZN(ybar[213]);
  AND2_X1 U131 ( .A1(a[13]), .A2(b[4]), .ZN(y[212]) );
  OR2_X1 U131bar ( .A1(abar[13]), .A2(bbar[4]), .ZN(ybar[212]);
  AND2_X1 U132 ( .A1(a[13]), .A2(b[3]), .ZN(y[211]) );
  OR2_X1 U132bar ( .A1(abar[13]), .A2(bbar[3]), .ZN(ybar[211]);
  AND2_X1 U133 ( .A1(a[13]), .A2(b[2]), .ZN(y[210]) );
  OR2_X1 U133bar ( .A1(abar[13]), .A2(bbar[2]), .ZN(ybar[210]);
  AND2_X1 U134 ( .A1(a[1]), .A2(b[4]), .ZN(y[20]) );
  OR2_X1 U134bar ( .A1(abar[1]), .A2(bbar[4]), .ZN(ybar[20]);
  AND2_X1 U135 ( .A1(a[13]), .A2(b[1]), .ZN(y[209]) );
  OR2_X1 U135bar ( .A1(abar[13]), .A2(bbar[1]), .ZN(ybar[209]);
  AND2_X1 U136 ( .A1(a[13]), .A2(b[0]), .ZN(y[208]) );
  OR2_X1 U136bar ( .A1(abar[13]), .A2(bbar[0]), .ZN(ybar[208]);
  AND2_X1 U137 ( .A1(a[12]), .A2(b[15]), .ZN(y[207]) );
  OR2_X1 U137bar ( .A1(abar[12]), .A2(bbar[15]), .ZN(ybar[207]);
  AND2_X1 U138 ( .A1(a[12]), .A2(b[14]), .ZN(y[206]) );
  OR2_X1 U138bar ( .A1(abar[12]), .A2(bbar[14]), .ZN(ybar[206]);
  AND2_X1 U139 ( .A1(a[12]), .A2(b[13]), .ZN(y[205]) );
  OR2_X1 U139bar ( .A1(abar[12]), .A2(bbar[13]), .ZN(ybar[205]);
  AND2_X1 U140 ( .A1(a[12]), .A2(b[12]), .ZN(y[204]) );
  OR2_X1 U140bar ( .A1(abar[12]), .A2(bbar[12]), .ZN(ybar[204]);
  AND2_X1 U141 ( .A1(a[12]), .A2(b[11]), .ZN(y[203]) );
  OR2_X1 U141bar ( .A1(abar[12]), .A2(bbar[11]), .ZN(ybar[203]);
  AND2_X1 U142 ( .A1(a[12]), .A2(b[10]), .ZN(y[202]) );
  OR2_X1 U142bar ( .A1(abar[12]), .A2(bbar[10]), .ZN(ybar[202]);
  AND2_X1 U143 ( .A1(a[12]), .A2(b[9]), .ZN(y[201]) );
  OR2_X1 U143bar ( .A1(abar[12]), .A2(bbar[9]), .ZN(ybar[201]);
  AND2_X1 U144 ( .A1(a[12]), .A2(b[8]), .ZN(y[200]) );
  OR2_X1 U144bar ( .A1(abar[12]), .A2(bbar[8]), .ZN(ybar[200]);
  AND2_X1 U145 ( .A1(b[1]), .A2(a[0]), .ZN(y[1]) );
  OR2_X1 U145bar ( .A1(bbar[1]), .A2(abar[0]), .ZN(ybar[1]);
  AND2_X1 U146 ( .A1(a[1]), .A2(b[3]), .ZN(y[19]) );
  OR2_X1 U146bar ( .A1(abar[1]), .A2(bbar[3]), .ZN(ybar[19]);
  AND2_X1 U147 ( .A1(a[12]), .A2(b[7]), .ZN(y[199]) );
  OR2_X1 U147bar ( .A1(abar[12]), .A2(bbar[7]), .ZN(ybar[199]);
  AND2_X1 U148 ( .A1(a[12]), .A2(b[6]), .ZN(y[198]) );
  OR2_X1 U148bar ( .A1(abar[12]), .A2(bbar[6]), .ZN(ybar[198]);
  AND2_X1 U149 ( .A1(a[12]), .A2(b[5]), .ZN(y[197]) );
  OR2_X1 U149bar ( .A1(abar[12]), .A2(bbar[5]), .ZN(ybar[197]);
  AND2_X1 U150 ( .A1(a[12]), .A2(b[4]), .ZN(y[196]) );
  OR2_X1 U150bar ( .A1(abar[12]), .A2(bbar[4]), .ZN(ybar[196]);
  AND2_X1 U151 ( .A1(a[12]), .A2(b[3]), .ZN(y[195]) );
  OR2_X1 U151bar ( .A1(abar[12]), .A2(bbar[3]), .ZN(ybar[195]);
  AND2_X1 U152 ( .A1(a[12]), .A2(b[2]), .ZN(y[194]) );
  OR2_X1 U152bar ( .A1(abar[12]), .A2(bbar[2]), .ZN(ybar[194]);
  AND2_X1 U153 ( .A1(a[12]), .A2(b[1]), .ZN(y[193]) );
  OR2_X1 U153bar ( .A1(abar[12]), .A2(bbar[1]), .ZN(ybar[193]);
  AND2_X1 U154 ( .A1(a[12]), .A2(b[0]), .ZN(y[192]) );
  OR2_X1 U154bar ( .A1(abar[12]), .A2(bbar[0]), .ZN(ybar[192]);
  AND2_X1 U155 ( .A1(a[11]), .A2(b[15]), .ZN(y[191]) );
  OR2_X1 U155bar ( .A1(abar[11]), .A2(bbar[15]), .ZN(ybar[191]);
  AND2_X1 U156 ( .A1(a[11]), .A2(b[14]), .ZN(y[190]) );
  OR2_X1 U156bar ( .A1(abar[11]), .A2(bbar[14]), .ZN(ybar[190]);
  AND2_X1 U157 ( .A1(a[1]), .A2(b[2]), .ZN(y[18]) );
  OR2_X1 U157bar ( .A1(abar[1]), .A2(bbar[2]), .ZN(ybar[18]);
  AND2_X1 U158 ( .A1(a[11]), .A2(b[13]), .ZN(y[189]) );
  OR2_X1 U158bar ( .A1(abar[11]), .A2(bbar[13]), .ZN(ybar[189]);
  AND2_X1 U159 ( .A1(a[11]), .A2(b[12]), .ZN(y[188]) );
  OR2_X1 U159bar ( .A1(abar[11]), .A2(bbar[12]), .ZN(ybar[188]);
  AND2_X1 U160 ( .A1(a[11]), .A2(b[11]), .ZN(y[187]) );
  OR2_X1 U160bar ( .A1(abar[11]), .A2(bbar[11]), .ZN(ybar[187]);
  AND2_X1 U161 ( .A1(a[11]), .A2(b[10]), .ZN(y[186]) );
  OR2_X1 U161bar ( .A1(abar[11]), .A2(bbar[10]), .ZN(ybar[186]);
  AND2_X1 U162 ( .A1(a[11]), .A2(b[9]), .ZN(y[185]) );
  OR2_X1 U162bar ( .A1(abar[11]), .A2(bbar[9]), .ZN(ybar[185]);
  AND2_X1 U163 ( .A1(a[11]), .A2(b[8]), .ZN(y[184]) );
  OR2_X1 U163bar ( .A1(abar[11]), .A2(bbar[8]), .ZN(ybar[184]);
  AND2_X1 U164 ( .A1(a[11]), .A2(b[7]), .ZN(y[183]) );
  OR2_X1 U164bar ( .A1(abar[11]), .A2(bbar[7]), .ZN(ybar[183]);
  AND2_X1 U165 ( .A1(a[11]), .A2(b[6]), .ZN(y[182]) );
  OR2_X1 U165bar ( .A1(abar[11]), .A2(bbar[6]), .ZN(ybar[182]);
  AND2_X1 U166 ( .A1(a[11]), .A2(b[5]), .ZN(y[181]) );
  OR2_X1 U166bar ( .A1(abar[11]), .A2(bbar[5]), .ZN(ybar[181]);
  AND2_X1 U167 ( .A1(a[11]), .A2(b[4]), .ZN(y[180]) );
  OR2_X1 U167bar ( .A1(abar[11]), .A2(bbar[4]), .ZN(ybar[180]);
  AND2_X1 U168 ( .A1(a[1]), .A2(b[1]), .ZN(y[17]) );
  OR2_X1 U168bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[17]);
  AND2_X1 U169 ( .A1(a[11]), .A2(b[3]), .ZN(y[179]) );
  OR2_X1 U169bar ( .A1(abar[11]), .A2(bbar[3]), .ZN(ybar[179]);
  AND2_X1 U170 ( .A1(a[11]), .A2(b[2]), .ZN(y[178]) );
  OR2_X1 U170bar ( .A1(abar[11]), .A2(bbar[2]), .ZN(ybar[178]);
  AND2_X1 U171 ( .A1(a[11]), .A2(b[1]), .ZN(y[177]) );
  OR2_X1 U171bar ( .A1(abar[11]), .A2(bbar[1]), .ZN(ybar[177]);
  AND2_X1 U172 ( .A1(a[11]), .A2(b[0]), .ZN(y[176]) );
  OR2_X1 U172bar ( .A1(abar[11]), .A2(bbar[0]), .ZN(ybar[176]);
  AND2_X1 U173 ( .A1(a[10]), .A2(b[15]), .ZN(y[175]) );
  OR2_X1 U173bar ( .A1(abar[10]), .A2(bbar[15]), .ZN(ybar[175]);
  AND2_X1 U174 ( .A1(a[10]), .A2(b[14]), .ZN(y[174]) );
  OR2_X1 U174bar ( .A1(abar[10]), .A2(bbar[14]), .ZN(ybar[174]);
  AND2_X1 U175 ( .A1(a[10]), .A2(b[13]), .ZN(y[173]) );
  OR2_X1 U175bar ( .A1(abar[10]), .A2(bbar[13]), .ZN(ybar[173]);
  AND2_X1 U176 ( .A1(a[10]), .A2(b[12]), .ZN(y[172]) );
  OR2_X1 U176bar ( .A1(abar[10]), .A2(bbar[12]), .ZN(ybar[172]);
  AND2_X1 U177 ( .A1(a[10]), .A2(b[11]), .ZN(y[171]) );
  OR2_X1 U177bar ( .A1(abar[10]), .A2(bbar[11]), .ZN(ybar[171]);
  AND2_X1 U178 ( .A1(a[10]), .A2(b[10]), .ZN(y[170]) );
  OR2_X1 U178bar ( .A1(abar[10]), .A2(bbar[10]), .ZN(ybar[170]);
  AND2_X1 U179 ( .A1(a[1]), .A2(b[0]), .ZN(y[16]) );
  OR2_X1 U179bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[16]);
  AND2_X1 U180 ( .A1(a[10]), .A2(b[9]), .ZN(y[169]) );
  OR2_X1 U180bar ( .A1(abar[10]), .A2(bbar[9]), .ZN(ybar[169]);
  AND2_X1 U181 ( .A1(a[10]), .A2(b[8]), .ZN(y[168]) );
  OR2_X1 U181bar ( .A1(abar[10]), .A2(bbar[8]), .ZN(ybar[168]);
  AND2_X1 U182 ( .A1(a[10]), .A2(b[7]), .ZN(y[167]) );
  OR2_X1 U182bar ( .A1(abar[10]), .A2(bbar[7]), .ZN(ybar[167]);
  AND2_X1 U183 ( .A1(a[10]), .A2(b[6]), .ZN(y[166]) );
  OR2_X1 U183bar ( .A1(abar[10]), .A2(bbar[6]), .ZN(ybar[166]);
  AND2_X1 U184 ( .A1(a[10]), .A2(b[5]), .ZN(y[165]) );
  OR2_X1 U184bar ( .A1(abar[10]), .A2(bbar[5]), .ZN(ybar[165]);
  AND2_X1 U185 ( .A1(a[10]), .A2(b[4]), .ZN(y[164]) );
  OR2_X1 U185bar ( .A1(abar[10]), .A2(bbar[4]), .ZN(ybar[164]);
  AND2_X1 U186 ( .A1(a[10]), .A2(b[3]), .ZN(y[163]) );
  OR2_X1 U186bar ( .A1(abar[10]), .A2(bbar[3]), .ZN(ybar[163]);
  AND2_X1 U187 ( .A1(a[10]), .A2(b[2]), .ZN(y[162]) );
  OR2_X1 U187bar ( .A1(abar[10]), .A2(bbar[2]), .ZN(ybar[162]);
  AND2_X1 U188 ( .A1(a[10]), .A2(b[1]), .ZN(y[161]) );
  OR2_X1 U188bar ( .A1(abar[10]), .A2(bbar[1]), .ZN(ybar[161]);
  AND2_X1 U189 ( .A1(a[10]), .A2(b[0]), .ZN(y[160]) );
  OR2_X1 U189bar ( .A1(abar[10]), .A2(bbar[0]), .ZN(ybar[160]);
  AND2_X1 U190 ( .A1(b[15]), .A2(a[0]), .ZN(y[15]) );
  OR2_X1 U190bar ( .A1(bbar[15]), .A2(abar[0]), .ZN(ybar[15]);
  AND2_X1 U191 ( .A1(a[9]), .A2(b[15]), .ZN(y[159]) );
  OR2_X1 U191bar ( .A1(abar[9]), .A2(bbar[15]), .ZN(ybar[159]);
  AND2_X1 U192 ( .A1(a[9]), .A2(b[14]), .ZN(y[158]) );
  OR2_X1 U192bar ( .A1(abar[9]), .A2(bbar[14]), .ZN(ybar[158]);
  AND2_X1 U193 ( .A1(a[9]), .A2(b[13]), .ZN(y[157]) );
  OR2_X1 U193bar ( .A1(abar[9]), .A2(bbar[13]), .ZN(ybar[157]);
  AND2_X1 U194 ( .A1(a[9]), .A2(b[12]), .ZN(y[156]) );
  OR2_X1 U194bar ( .A1(abar[9]), .A2(bbar[12]), .ZN(ybar[156]);
  AND2_X1 U195 ( .A1(a[9]), .A2(b[11]), .ZN(y[155]) );
  OR2_X1 U195bar ( .A1(abar[9]), .A2(bbar[11]), .ZN(ybar[155]);
  AND2_X1 U196 ( .A1(a[9]), .A2(b[10]), .ZN(y[154]) );
  OR2_X1 U196bar ( .A1(abar[9]), .A2(bbar[10]), .ZN(ybar[154]);
  AND2_X1 U197 ( .A1(a[9]), .A2(b[9]), .ZN(y[153]) );
  OR2_X1 U197bar ( .A1(abar[9]), .A2(bbar[9]), .ZN(ybar[153]);
  AND2_X1 U198 ( .A1(a[9]), .A2(b[8]), .ZN(y[152]) );
  OR2_X1 U198bar ( .A1(abar[9]), .A2(bbar[8]), .ZN(ybar[152]);
  AND2_X1 U199 ( .A1(a[9]), .A2(b[7]), .ZN(y[151]) );
  OR2_X1 U199bar ( .A1(abar[9]), .A2(bbar[7]), .ZN(ybar[151]);
  AND2_X1 U200 ( .A1(a[9]), .A2(b[6]), .ZN(y[150]) );
  OR2_X1 U200bar ( .A1(abar[9]), .A2(bbar[6]), .ZN(ybar[150]);
  AND2_X1 U201 ( .A1(b[14]), .A2(a[0]), .ZN(y[14]) );
  OR2_X1 U201bar ( .A1(bbar[14]), .A2(abar[0]), .ZN(ybar[14]);
  AND2_X1 U202 ( .A1(a[9]), .A2(b[5]), .ZN(y[149]) );
  OR2_X1 U202bar ( .A1(abar[9]), .A2(bbar[5]), .ZN(ybar[149]);
  AND2_X1 U203 ( .A1(a[9]), .A2(b[4]), .ZN(y[148]) );
  OR2_X1 U203bar ( .A1(abar[9]), .A2(bbar[4]), .ZN(ybar[148]);
  AND2_X1 U204 ( .A1(a[9]), .A2(b[3]), .ZN(y[147]) );
  OR2_X1 U204bar ( .A1(abar[9]), .A2(bbar[3]), .ZN(ybar[147]);
  AND2_X1 U205 ( .A1(a[9]), .A2(b[2]), .ZN(y[146]) );
  OR2_X1 U205bar ( .A1(abar[9]), .A2(bbar[2]), .ZN(ybar[146]);
  AND2_X1 U206 ( .A1(a[9]), .A2(b[1]), .ZN(y[145]) );
  OR2_X1 U206bar ( .A1(abar[9]), .A2(bbar[1]), .ZN(ybar[145]);
  AND2_X1 U207 ( .A1(a[9]), .A2(b[0]), .ZN(y[144]) );
  OR2_X1 U207bar ( .A1(abar[9]), .A2(bbar[0]), .ZN(ybar[144]);
  AND2_X1 U208 ( .A1(a[8]), .A2(b[15]), .ZN(y[143]) );
  OR2_X1 U208bar ( .A1(abar[8]), .A2(bbar[15]), .ZN(ybar[143]);
  AND2_X1 U209 ( .A1(a[8]), .A2(b[14]), .ZN(y[142]) );
  OR2_X1 U209bar ( .A1(abar[8]), .A2(bbar[14]), .ZN(ybar[142]);
  AND2_X1 U210 ( .A1(a[8]), .A2(b[13]), .ZN(y[141]) );
  OR2_X1 U210bar ( .A1(abar[8]), .A2(bbar[13]), .ZN(ybar[141]);
  AND2_X1 U211 ( .A1(a[8]), .A2(b[12]), .ZN(y[140]) );
  OR2_X1 U211bar ( .A1(abar[8]), .A2(bbar[12]), .ZN(ybar[140]);
  AND2_X1 U212 ( .A1(b[13]), .A2(a[0]), .ZN(y[13]) );
  OR2_X1 U212bar ( .A1(bbar[13]), .A2(abar[0]), .ZN(ybar[13]);
  AND2_X1 U213 ( .A1(a[8]), .A2(b[11]), .ZN(y[139]) );
  OR2_X1 U213bar ( .A1(abar[8]), .A2(bbar[11]), .ZN(ybar[139]);
  AND2_X1 U214 ( .A1(a[8]), .A2(b[10]), .ZN(y[138]) );
  OR2_X1 U214bar ( .A1(abar[8]), .A2(bbar[10]), .ZN(ybar[138]);
  AND2_X1 U215 ( .A1(a[8]), .A2(b[9]), .ZN(y[137]) );
  OR2_X1 U215bar ( .A1(abar[8]), .A2(bbar[9]), .ZN(ybar[137]);
  AND2_X1 U216 ( .A1(a[8]), .A2(b[8]), .ZN(y[136]) );
  OR2_X1 U216bar ( .A1(abar[8]), .A2(bbar[8]), .ZN(ybar[136]);
  AND2_X1 U217 ( .A1(a[8]), .A2(b[7]), .ZN(y[135]) );
  OR2_X1 U217bar ( .A1(abar[8]), .A2(bbar[7]), .ZN(ybar[135]);
  AND2_X1 U218 ( .A1(a[8]), .A2(b[6]), .ZN(y[134]) );
  OR2_X1 U218bar ( .A1(abar[8]), .A2(bbar[6]), .ZN(ybar[134]);
  AND2_X1 U219 ( .A1(a[8]), .A2(b[5]), .ZN(y[133]) );
  OR2_X1 U219bar ( .A1(abar[8]), .A2(bbar[5]), .ZN(ybar[133]);
  AND2_X1 U220 ( .A1(a[8]), .A2(b[4]), .ZN(y[132]) );
  OR2_X1 U220bar ( .A1(abar[8]), .A2(bbar[4]), .ZN(ybar[132]);
  AND2_X1 U221 ( .A1(a[8]), .A2(b[3]), .ZN(y[131]) );
  OR2_X1 U221bar ( .A1(abar[8]), .A2(bbar[3]), .ZN(ybar[131]);
  AND2_X1 U222 ( .A1(a[8]), .A2(b[2]), .ZN(y[130]) );
  OR2_X1 U222bar ( .A1(abar[8]), .A2(bbar[2]), .ZN(ybar[130]);
  AND2_X1 U223 ( .A1(b[12]), .A2(a[0]), .ZN(y[12]) );
  OR2_X1 U223bar ( .A1(bbar[12]), .A2(abar[0]), .ZN(ybar[12]);
  AND2_X1 U224 ( .A1(a[8]), .A2(b[1]), .ZN(y[129]) );
  OR2_X1 U224bar ( .A1(abar[8]), .A2(bbar[1]), .ZN(ybar[129]);
  AND2_X1 U225 ( .A1(a[8]), .A2(b[0]), .ZN(y[128]) );
  OR2_X1 U225bar ( .A1(abar[8]), .A2(bbar[0]), .ZN(ybar[128]);
  AND2_X1 U226 ( .A1(a[7]), .A2(b[15]), .ZN(y[127]) );
  OR2_X1 U226bar ( .A1(abar[7]), .A2(bbar[15]), .ZN(ybar[127]);
  AND2_X1 U227 ( .A1(a[7]), .A2(b[14]), .ZN(y[126]) );
  OR2_X1 U227bar ( .A1(abar[7]), .A2(bbar[14]), .ZN(ybar[126]);
  AND2_X1 U228 ( .A1(a[7]), .A2(b[13]), .ZN(y[125]) );
  OR2_X1 U228bar ( .A1(abar[7]), .A2(bbar[13]), .ZN(ybar[125]);
  AND2_X1 U229 ( .A1(a[7]), .A2(b[12]), .ZN(y[124]) );
  OR2_X1 U229bar ( .A1(abar[7]), .A2(bbar[12]), .ZN(ybar[124]);
  AND2_X1 U230 ( .A1(a[7]), .A2(b[11]), .ZN(y[123]) );
  OR2_X1 U230bar ( .A1(abar[7]), .A2(bbar[11]), .ZN(ybar[123]);
  AND2_X1 U231 ( .A1(a[7]), .A2(b[10]), .ZN(y[122]) );
  OR2_X1 U231bar ( .A1(abar[7]), .A2(bbar[10]), .ZN(ybar[122]);
  AND2_X1 U232 ( .A1(a[7]), .A2(b[9]), .ZN(y[121]) );
  OR2_X1 U232bar ( .A1(abar[7]), .A2(bbar[9]), .ZN(ybar[121]);
  AND2_X1 U233 ( .A1(a[7]), .A2(b[8]), .ZN(y[120]) );
  OR2_X1 U233bar ( .A1(abar[7]), .A2(bbar[8]), .ZN(ybar[120]);
  AND2_X1 U234 ( .A1(b[11]), .A2(a[0]), .ZN(y[11]) );
  OR2_X1 U234bar ( .A1(bbar[11]), .A2(abar[0]), .ZN(ybar[11]);
  AND2_X1 U235 ( .A1(a[7]), .A2(b[7]), .ZN(y[119]) );
  OR2_X1 U235bar ( .A1(abar[7]), .A2(bbar[7]), .ZN(ybar[119]);
  AND2_X1 U236 ( .A1(a[7]), .A2(b[6]), .ZN(y[118]) );
  OR2_X1 U236bar ( .A1(abar[7]), .A2(bbar[6]), .ZN(ybar[118]);
  AND2_X1 U237 ( .A1(a[7]), .A2(b[5]), .ZN(y[117]) );
  OR2_X1 U237bar ( .A1(abar[7]), .A2(bbar[5]), .ZN(ybar[117]);
  AND2_X1 U238 ( .A1(a[7]), .A2(b[4]), .ZN(y[116]) );
  OR2_X1 U238bar ( .A1(abar[7]), .A2(bbar[4]), .ZN(ybar[116]);
  AND2_X1 U239 ( .A1(a[7]), .A2(b[3]), .ZN(y[115]) );
  OR2_X1 U239bar ( .A1(abar[7]), .A2(bbar[3]), .ZN(ybar[115]);
  AND2_X1 U240 ( .A1(a[7]), .A2(b[2]), .ZN(y[114]) );
  OR2_X1 U240bar ( .A1(abar[7]), .A2(bbar[2]), .ZN(ybar[114]);
  AND2_X1 U241 ( .A1(a[7]), .A2(b[1]), .ZN(y[113]) );
  OR2_X1 U241bar ( .A1(abar[7]), .A2(bbar[1]), .ZN(ybar[113]);
  AND2_X1 U242 ( .A1(a[7]), .A2(b[0]), .ZN(y[112]) );
  OR2_X1 U242bar ( .A1(abar[7]), .A2(bbar[0]), .ZN(ybar[112]);
  AND2_X1 U243 ( .A1(b[15]), .A2(a[6]), .ZN(y[111]) );
  OR2_X1 U243bar ( .A1(bbar[15]), .A2(abar[6]), .ZN(ybar[111]);
  AND2_X1 U244 ( .A1(b[14]), .A2(a[6]), .ZN(y[110]) );
  OR2_X1 U244bar ( .A1(bbar[14]), .A2(abar[6]), .ZN(ybar[110]);
  AND2_X1 U245 ( .A1(b[10]), .A2(a[0]), .ZN(y[10]) );
  OR2_X1 U245bar ( .A1(bbar[10]), .A2(abar[0]), .ZN(ybar[10]);
  AND2_X1 U246 ( .A1(b[13]), .A2(a[6]), .ZN(y[109]) );
  OR2_X1 U246bar ( .A1(bbar[13]), .A2(abar[6]), .ZN(ybar[109]);
  AND2_X1 U247 ( .A1(b[12]), .A2(a[6]), .ZN(y[108]) );
  OR2_X1 U247bar ( .A1(bbar[12]), .A2(abar[6]), .ZN(ybar[108]);
  AND2_X1 U248 ( .A1(b[11]), .A2(a[6]), .ZN(y[107]) );
  OR2_X1 U248bar ( .A1(bbar[11]), .A2(abar[6]), .ZN(ybar[107]);
  AND2_X1 U249 ( .A1(b[10]), .A2(a[6]), .ZN(y[106]) );
  OR2_X1 U249bar ( .A1(bbar[10]), .A2(abar[6]), .ZN(ybar[106]);
  AND2_X1 U250 ( .A1(a[6]), .A2(b[9]), .ZN(y[105]) );
  OR2_X1 U250bar ( .A1(abar[6]), .A2(bbar[9]), .ZN(ybar[105]);
  AND2_X1 U251 ( .A1(b[8]), .A2(a[6]), .ZN(y[104]) );
  OR2_X1 U251bar ( .A1(bbar[8]), .A2(abar[6]), .ZN(ybar[104]);
  AND2_X1 U252 ( .A1(b[7]), .A2(a[6]), .ZN(y[103]) );
  OR2_X1 U252bar ( .A1(bbar[7]), .A2(abar[6]), .ZN(ybar[103]);
  AND2_X1 U253 ( .A1(b[6]), .A2(a[6]), .ZN(y[102]) );
  OR2_X1 U253bar ( .A1(bbar[6]), .A2(abar[6]), .ZN(ybar[102]);
  AND2_X1 U254 ( .A1(b[5]), .A2(a[6]), .ZN(y[101]) );
  OR2_X1 U254bar ( .A1(bbar[5]), .A2(abar[6]), .ZN(ybar[101]);
  AND2_X1 U255 ( .A1(b[4]), .A2(a[6]), .ZN(y[100]) );
  OR2_X1 U255bar ( .A1(bbar[4]), .A2(abar[6]), .ZN(ybar[100]);
  AND2_X1 U256 ( .A1(b[0]), .A2(a[0]), .ZN(y[0]) );
  OR2_X1 U256bar ( .A1(bbar[0]), .A2(abar[0]), .ZN(ybar[0]);
endmodule




module decode_8 ( in, out );
  input [7:0] in;
  //input_done

  output [255:0] out;
  //output_done

  wire   [15:0] level1;
  wire   [31:0] level2;
  //wire_done

  CD2_32 cd_l1_1 ( .a(in[1]), .b(in[0]), .y(level1[3:0]) );
  CD2_31 cd_l1_2 ( .a(in[3]), .b(in[2]), .y(level1[7:4]) );
  CD2_30 cd_l1_3 ( .a(in[5]), .b(in[4]), .y(level1[11:8]) );
  CD2_29 cd_l1_4 ( .a(in[7]), .b(in[6]), .y(level1[15:12]) );
  CD4_16 cd_l2_1 ( .a(level1[7:4]), .b(level1[3:0]), .y(level2[15:0]) );
  CD4_15 cd_l2_2 ( .a(level1[15:12]), .b(level1[11:8]), .y(level2[31:16]) );
  CD16_8 cd_l3 ( .a(level2[31:16]), .b(level2[15:0]), .y(out) );
endmodule


module encode_8 ( in, out );
  input [255:0] in;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
  assign inbar[8] = ~in[8];
  assign inbar[9] = ~in[9];
  assign inbar[10] = ~in[10];
  assign inbar[11] = ~in[11];
  assign inbar[12] = ~in[12];
  assign inbar[13] = ~in[13];
  assign inbar[14] = ~in[14];
  assign inbar[15] = ~in[15];
  assign inbar[16] = ~in[16];
  assign inbar[17] = ~in[17];
  assign inbar[18] = ~in[18];
  assign inbar[19] = ~in[19];
  assign inbar[20] = ~in[20];
  assign inbar[21] = ~in[21];
  assign inbar[22] = ~in[22];
  assign inbar[23] = ~in[23];
  assign inbar[24] = ~in[24];
  assign inbar[25] = ~in[25];
  assign inbar[26] = ~in[26];
  assign inbar[27] = ~in[27];
  assign inbar[28] = ~in[28];
  assign inbar[29] = ~in[29];
  assign inbar[30] = ~in[30];
  assign inbar[31] = ~in[31];
  assign inbar[32] = ~in[32];
  assign inbar[33] = ~in[33];
  assign inbar[34] = ~in[34];
  assign inbar[35] = ~in[35];
  assign inbar[36] = ~in[36];
  assign inbar[37] = ~in[37];
  assign inbar[38] = ~in[38];
  assign inbar[39] = ~in[39];
  assign inbar[40] = ~in[40];
  assign inbar[41] = ~in[41];
  assign inbar[42] = ~in[42];
  assign inbar[43] = ~in[43];
  assign inbar[44] = ~in[44];
  assign inbar[45] = ~in[45];
  assign inbar[46] = ~in[46];
  assign inbar[47] = ~in[47];
  assign inbar[48] = ~in[48];
  assign inbar[49] = ~in[49];
  assign inbar[50] = ~in[50];
  assign inbar[51] = ~in[51];
  assign inbar[52] = ~in[52];
  assign inbar[53] = ~in[53];
  assign inbar[54] = ~in[54];
  assign inbar[55] = ~in[55];
  assign inbar[56] = ~in[56];
  assign inbar[57] = ~in[57];
  assign inbar[58] = ~in[58];
  assign inbar[59] = ~in[59];
  assign inbar[60] = ~in[60];
  assign inbar[61] = ~in[61];
  assign inbar[62] = ~in[62];
  assign inbar[63] = ~in[63];
  assign inbar[64] = ~in[64];
  assign inbar[65] = ~in[65];
  assign inbar[66] = ~in[66];
  assign inbar[67] = ~in[67];
  assign inbar[68] = ~in[68];
  assign inbar[69] = ~in[69];
  assign inbar[70] = ~in[70];
  assign inbar[71] = ~in[71];
  assign inbar[72] = ~in[72];
  assign inbar[73] = ~in[73];
  assign inbar[74] = ~in[74];
  assign inbar[75] = ~in[75];
  assign inbar[76] = ~in[76];
  assign inbar[77] = ~in[77];
  assign inbar[78] = ~in[78];
  assign inbar[79] = ~in[79];
  assign inbar[80] = ~in[80];
  assign inbar[81] = ~in[81];
  assign inbar[82] = ~in[82];
  assign inbar[83] = ~in[83];
  assign inbar[84] = ~in[84];
  assign inbar[85] = ~in[85];
  assign inbar[86] = ~in[86];
  assign inbar[87] = ~in[87];
  assign inbar[88] = ~in[88];
  assign inbar[89] = ~in[89];
  assign inbar[90] = ~in[90];
  assign inbar[91] = ~in[91];
  assign inbar[92] = ~in[92];
  assign inbar[93] = ~in[93];
  assign inbar[94] = ~in[94];
  assign inbar[95] = ~in[95];
  assign inbar[96] = ~in[96];
  assign inbar[97] = ~in[97];
  assign inbar[98] = ~in[98];
  assign inbar[99] = ~in[99];
  assign inbar[100] = ~in[100];
  assign inbar[101] = ~in[101];
  assign inbar[102] = ~in[102];
  assign inbar[103] = ~in[103];
  assign inbar[104] = ~in[104];
  assign inbar[105] = ~in[105];
  assign inbar[106] = ~in[106];
  assign inbar[107] = ~in[107];
  assign inbar[108] = ~in[108];
  assign inbar[109] = ~in[109];
  assign inbar[110] = ~in[110];
  assign inbar[111] = ~in[111];
  assign inbar[112] = ~in[112];
  assign inbar[113] = ~in[113];
  assign inbar[114] = ~in[114];
  assign inbar[115] = ~in[115];
  assign inbar[116] = ~in[116];
  assign inbar[117] = ~in[117];
  assign inbar[118] = ~in[118];
  assign inbar[119] = ~in[119];
  assign inbar[120] = ~in[120];
  assign inbar[121] = ~in[121];
  assign inbar[122] = ~in[122];
  assign inbar[123] = ~in[123];
  assign inbar[124] = ~in[124];
  assign inbar[125] = ~in[125];
  assign inbar[126] = ~in[126];
  assign inbar[127] = ~in[127];
  assign inbar[128] = ~in[128];
  assign inbar[129] = ~in[129];
  assign inbar[130] = ~in[130];
  assign inbar[131] = ~in[131];
  assign inbar[132] = ~in[132];
  assign inbar[133] = ~in[133];
  assign inbar[134] = ~in[134];
  assign inbar[135] = ~in[135];
  assign inbar[136] = ~in[136];
  assign inbar[137] = ~in[137];
  assign inbar[138] = ~in[138];
  assign inbar[139] = ~in[139];
  assign inbar[140] = ~in[140];
  assign inbar[141] = ~in[141];
  assign inbar[142] = ~in[142];
  assign inbar[143] = ~in[143];
  assign inbar[144] = ~in[144];
  assign inbar[145] = ~in[145];
  assign inbar[146] = ~in[146];
  assign inbar[147] = ~in[147];
  assign inbar[148] = ~in[148];
  assign inbar[149] = ~in[149];
  assign inbar[150] = ~in[150];
  assign inbar[151] = ~in[151];
  assign inbar[152] = ~in[152];
  assign inbar[153] = ~in[153];
  assign inbar[154] = ~in[154];
  assign inbar[155] = ~in[155];
  assign inbar[156] = ~in[156];
  assign inbar[157] = ~in[157];
  assign inbar[158] = ~in[158];
  assign inbar[159] = ~in[159];
  assign inbar[160] = ~in[160];
  assign inbar[161] = ~in[161];
  assign inbar[162] = ~in[162];
  assign inbar[163] = ~in[163];
  assign inbar[164] = ~in[164];
  assign inbar[165] = ~in[165];
  assign inbar[166] = ~in[166];
  assign inbar[167] = ~in[167];
  assign inbar[168] = ~in[168];
  assign inbar[169] = ~in[169];
  assign inbar[170] = ~in[170];
  assign inbar[171] = ~in[171];
  assign inbar[172] = ~in[172];
  assign inbar[173] = ~in[173];
  assign inbar[174] = ~in[174];
  assign inbar[175] = ~in[175];
  assign inbar[176] = ~in[176];
  assign inbar[177] = ~in[177];
  assign inbar[178] = ~in[178];
  assign inbar[179] = ~in[179];
  assign inbar[180] = ~in[180];
  assign inbar[181] = ~in[181];
  assign inbar[182] = ~in[182];
  assign inbar[183] = ~in[183];
  assign inbar[184] = ~in[184];
  assign inbar[185] = ~in[185];
  assign inbar[186] = ~in[186];
  assign inbar[187] = ~in[187];
  assign inbar[188] = ~in[188];
  assign inbar[189] = ~in[189];
  assign inbar[190] = ~in[190];
  assign inbar[191] = ~in[191];
  assign inbar[192] = ~in[192];
  assign inbar[193] = ~in[193];
  assign inbar[194] = ~in[194];
  assign inbar[195] = ~in[195];
  assign inbar[196] = ~in[196];
  assign inbar[197] = ~in[197];
  assign inbar[198] = ~in[198];
  assign inbar[199] = ~in[199];
  assign inbar[200] = ~in[200];
  assign inbar[201] = ~in[201];
  assign inbar[202] = ~in[202];
  assign inbar[203] = ~in[203];
  assign inbar[204] = ~in[204];
  assign inbar[205] = ~in[205];
  assign inbar[206] = ~in[206];
  assign inbar[207] = ~in[207];
  assign inbar[208] = ~in[208];
  assign inbar[209] = ~in[209];
  assign inbar[210] = ~in[210];
  assign inbar[211] = ~in[211];
  assign inbar[212] = ~in[212];
  assign inbar[213] = ~in[213];
  assign inbar[214] = ~in[214];
  assign inbar[215] = ~in[215];
  assign inbar[216] = ~in[216];
  assign inbar[217] = ~in[217];
  assign inbar[218] = ~in[218];
  assign inbar[219] = ~in[219];
  assign inbar[220] = ~in[220];
  assign inbar[221] = ~in[221];
  assign inbar[222] = ~in[222];
  assign inbar[223] = ~in[223];
  assign inbar[224] = ~in[224];
  assign inbar[225] = ~in[225];
  assign inbar[226] = ~in[226];
  assign inbar[227] = ~in[227];
  assign inbar[228] = ~in[228];
  assign inbar[229] = ~in[229];
  assign inbar[230] = ~in[230];
  assign inbar[231] = ~in[231];
  assign inbar[232] = ~in[232];
  assign inbar[233] = ~in[233];
  assign inbar[234] = ~in[234];
  assign inbar[235] = ~in[235];
  assign inbar[236] = ~in[236];
  assign inbar[237] = ~in[237];
  assign inbar[238] = ~in[238];
  assign inbar[239] = ~in[239];
  assign inbar[240] = ~in[240];
  assign inbar[241] = ~in[241];
  assign inbar[242] = ~in[242];
  assign inbar[243] = ~in[243];
  assign inbar[244] = ~in[244];
  assign inbar[245] = ~in[245];
  assign inbar[246] = ~in[246];
  assign inbar[247] = ~in[247];
  assign inbar[248] = ~in[248];
  assign inbar[249] = ~in[249];
  assign inbar[250] = ~in[250];
  assign inbar[251] = ~in[251];
  assign inbar[252] = ~in[252];
  assign inbar[253] = ~in[253];
  assign inbar[254] = ~in[254];
  assign inbar[255] = ~in[255];
  //input_done

  output [7:0] out;
  reg [7:0] outbar;
  //output_done

  wire   in_81, in_80, in_79, in_78, in_77, in_76, in_75, in_74, in_73, in_72,
         in_71, in_70, in_69, in_68, in_67, in_66, in_65, in_64, in_63, in_62,
         in_61, in_60, in_59, in_58, in_57, in_56, in_55, in_54, in_53, in_52,
         in_51, in_50, in_49, in_48, in_47, in_46, in_45, in_44, in_43, in_42,
         in_41, in_40, in_39, in_38, in_37, in_36, in_35, in_34, in_33, in_32,
         in_31, in_30, in_29, in_28, in_27, in_26, in_25, in_24, in_23, in_22,
         in_21, in_20, in_19, in_18, in_17, in_16, in_15, in_14, in_13, in_12,
         in_11, in_10, in_9, in_8, in_7, in_6, in_5, in_4, in_3, in_2, in_1,
         in_0, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972;
  wire in_81bar, in_80bar, in_79bar, in_78bar, in_77bar, in_76bar, in_75bar, in_74bar, in_73bar, in_72bar, in_71bar, in_70bar, in_69bar, in_68bar, in_67bar, in_66bar, in_65bar, in_64bar, in_63bar, in_62bar, in_61bar, in_60bar, in_59bar, in_58bar, in_57bar, in_56bar, in_55bar, in_54bar, in_53bar, in_52bar, in_51bar, in_50bar, in_49bar, in_48bar, in_47bar, in_46bar, in_45bar, in_44bar, in_43bar, in_42bar, in_41bar, in_40bar, in_39bar, in_38bar, in_37bar, in_36bar, in_35bar, in_34bar, in_33bar, in_32bar, in_31bar, in_30bar, in_29bar, in_28bar, in_27bar, in_26bar, in_25bar, in_24bar, in_23bar, in_22bar, in_21bar, in_20bar, in_19bar, in_18bar, in_17bar, in_16bar, in_15bar, in_14bar, in_13bar, in_12bar, in_11bar, in_10bar, in_9bar, in_8bar, in_7bar, in_6bar, in_5bar, in_4bar, in_3bar, in_2bar, in_1bar, in_0bar, n487bar, n488bar, n489bar, n490bar, n491bar, n492bar, n493bar, n494bar, n495bar, n496bar, n497bar, n498bar, n499bar, n500bar, n501bar, n502bar, n503bar, n504bar, n505bar, n506bar, n507bar, n508bar, n509bar, n510bar, n511bar, n512bar, n513bar, n514bar, n515bar, n516bar, n517bar, n518bar, n519bar, n520bar, n521bar, n522bar, n523bar, n524bar, n525bar, n526bar, n527bar, n528bar, n529bar, n530bar, n531bar, n532bar, n533bar, n534bar, n535bar, n536bar, n537bar, n538bar, n539bar, n540bar, n541bar, n542bar, n543bar, n544bar, n545bar, n546bar, n547bar, n548bar, n549bar, n550bar, n551bar, n552bar, n553bar, n554bar, n555bar, n556bar, n557bar, n558bar, n559bar, n560bar, n561bar, n562bar, n563bar, n564bar, n565bar, n566bar, n567bar, n568bar, n569bar, n570bar, n571bar, n572bar, n573bar, n574bar, n575bar, n576bar, n577bar, n578bar, n579bar, n580bar, n581bar, n582bar, n583bar, n584bar, n585bar, n586bar, n587bar, n588bar, n589bar, n590bar, n591bar, n592bar, n593bar, n594bar, n595bar, n596bar, n597bar, n598bar, n599bar, n600bar, n601bar, n602bar, n603bar, n604bar, n605bar, n606bar, n607bar, n608bar, n609bar, n610bar, n611bar, n612bar, n613bar, n614bar, n615bar, n616bar, n617bar, n618bar, n619bar, n620bar, n621bar, n622bar, n623bar, n624bar, n625bar, n626bar, n627bar, n628bar, n629bar, n630bar, n631bar, n632bar, n633bar, n634bar, n635bar, n636bar, n637bar, n638bar, n639bar, n640bar, n641bar, n642bar, n643bar, n644bar, n645bar, n646bar, n647bar, n648bar, n649bar, n650bar, n651bar, n652bar, n653bar, n654bar, n655bar, n656bar, n657bar, n658bar, n659bar, n660bar, n661bar, n662bar, n663bar, n664bar, n665bar, n666bar, n667bar, n668bar, n669bar, n670bar, n671bar, n672bar, n673bar, n674bar, n675bar, n676bar, n677bar, n678bar, n679bar, n680bar, n681bar, n682bar, n683bar, n684bar, n685bar, n686bar, n687bar, n688bar, n689bar, n690bar, n691bar, n692bar, n693bar, n694bar, n695bar, n696bar, n697bar, n698bar, n699bar, n700bar, n701bar, n702bar, n703bar, n704bar, n705bar, n706bar, n707bar, n708bar, n709bar, n710bar, n711bar, n712bar, n713bar, n714bar, n715bar, n716bar, n717bar, n718bar, n719bar, n720bar, n721bar, n722bar, n723bar, n724bar, n725bar, n726bar, n727bar, n728bar, n729bar, n730bar, n731bar, n732bar, n733bar, n734bar, n735bar, n736bar, n737bar, n738bar, n739bar, n740bar, n741bar, n742bar, n743bar, n744bar, n745bar, n746bar, n747bar, n748bar, n749bar, n750bar, n751bar, n752bar, n753bar, n754bar, n755bar, n756bar, n757bar, n758bar, n759bar, n760bar, n761bar, n762bar, n763bar, n764bar, n765bar, n766bar, n767bar, n768bar, n769bar, n770bar, n771bar, n772bar, n773bar, n774bar, n775bar, n776bar, n777bar, n778bar, n779bar, n780bar, n781bar, n782bar, n783bar, n784bar, n785bar, n786bar, n787bar, n788bar, n789bar, n790bar, n791bar, n792bar, n793bar, n794bar, n795bar, n796bar, n797bar, n798bar, n799bar, n800bar, n801bar, n802bar, n803bar, n804bar, n805bar, n806bar, n807bar, n808bar, n809bar, n810bar, n811bar, n812bar, n813bar, n814bar, n815bar, n816bar, n817bar, n818bar, n819bar, n820bar, n821bar, n822bar, n823bar, n824bar, n825bar, n826bar, n827bar, n828bar, n829bar, n830bar, n831bar, n832bar, n833bar, n834bar, n835bar, n836bar, n837bar, n838bar, n839bar, n840bar, n841bar, n842bar, n843bar, n844bar, n845bar, n846bar, n847bar, n848bar, n849bar, n850bar, n851bar, n852bar, n853bar, n854bar, n855bar, n856bar, n857bar, n858bar, n859bar, n860bar, n861bar, n862bar, n863bar, n864bar, n865bar, n866bar, n867bar, n868bar, n869bar, n870bar, n871bar, n872bar, n873bar, n874bar, n875bar, n876bar, n877bar, n878bar, n879bar, n880bar, n881bar, n882bar, n883bar, n884bar, n885bar, n886bar, n887bar, n888bar, n889bar, n890bar, n891bar, n892bar, n893bar, n894bar, n895bar, n896bar, n897bar, n898bar, n899bar, n900bar, n901bar, n902bar, n903bar, n904bar, n905bar, n906bar, n907bar, n908bar, n909bar, n910bar, n911bar, n912bar, n913bar, n914bar, n915bar, n916bar, n917bar, n918bar, n919bar, n920bar, n921bar, n922bar, n923bar, n924bar, n925bar, n926bar, n927bar, n928bar, n929bar, n930bar, n931bar, n932bar, n933bar, n934bar, n935bar, n936bar, n937bar, n938bar, n939bar, n940bar, n941bar, n942bar, n943bar, n944bar, n945bar, n946bar, n947bar, n948bar, n949bar, n950bar, n951bar, n952bar, n953bar, n954bar, n955bar, n956bar, n957bar, n958bar, n959bar, n960bar, n961bar, n962bar, n963bar, n964bar, n965bar, n966bar, n967bar, n968bar, n969bar, n970bar, n971bar, n972bar;
  //wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];

  OR2_X1 U1 ( .A1(n972), .A2(n971), .ZN(out[7]) );
  AND2_X1 U1bar ( .A1(n972bar), .A2(n971bar), .ZN(outbar[7]);
  OR2_X1 U2 ( .A1(n970), .A2(n969), .ZN(n971) );
  AND2_X1 U2bar ( .A1(n970bar), .A2(n969bar), .ZN(n971bar);
  OR2_X1 U3 ( .A1(n968), .A2(n967), .ZN(n969) );
  AND2_X1 U3bar ( .A1(n968bar), .A2(n967bar), .ZN(n969bar);
  OR2_X1 U4 ( .A1(n966), .A2(n965), .ZN(n967) );
  AND2_X1 U4bar ( .A1(n966bar), .A2(n965bar), .ZN(n967bar);
  OR2_X1 U5 ( .A1(n964), .A2(n963), .ZN(n968) );
  AND2_X1 U5bar ( .A1(n964bar), .A2(n963bar), .ZN(n968bar);
  OR2_X1 U6 ( .A1(in[116]), .A2(n962), .ZN(n963) );
  AND2_X1 U6bar ( .A1(inbar[116]), .A2(n962bar), .ZN(n963bar);
  OR2_X1 U7 ( .A1(n961), .A2(n960), .ZN(n970) );
  AND2_X1 U7bar ( .A1(n961bar), .A2(n960bar), .ZN(n970bar);
  OR2_X1 U8 ( .A1(in[150]), .A2(in[127]), .ZN(n960) );
  AND2_X1 U8bar ( .A1(inbar[150]), .A2(inbar[127]), .ZN(n960bar);
  OR2_X1 U9 ( .A1(in[160]), .A2(n959), .ZN(n961) );
  AND2_X1 U9bar ( .A1(inbar[160]), .A2(n959bar), .ZN(n961bar);
  OR2_X1 U10 ( .A1(in[252]), .A2(in[168]), .ZN(n959) );
  AND2_X1 U10bar ( .A1(inbar[252]), .A2(inbar[168]), .ZN(n959bar);
  OR2_X1 U11 ( .A1(n958), .A2(n957), .ZN(n972) );
  AND2_X1 U11bar ( .A1(n958bar), .A2(n957bar), .ZN(n972bar);
  OR2_X1 U12 ( .A1(n956), .A2(n955), .ZN(n957) );
  AND2_X1 U12bar ( .A1(n956bar), .A2(n955bar), .ZN(n957bar);
  OR2_X1 U13 ( .A1(in_17), .A2(in[96]), .ZN(n955) );
  AND2_X1 U13bar ( .A1(in_17bar), .A2(inbar[96]), .ZN(n955bar);
  OR2_X1 U14 ( .A1(in_23), .A2(n954), .ZN(n956) );
  AND2_X1 U14bar ( .A1(in_23bar), .A2(n954bar), .ZN(n956bar);
  OR2_X1 U15 ( .A1(in_31), .A2(in_26), .ZN(n954) );
  AND2_X1 U15bar ( .A1(in_31bar), .A2(in_26bar), .ZN(n954bar);
  OR2_X1 U16 ( .A1(n953), .A2(n952), .ZN(n958) );
  AND2_X1 U16bar ( .A1(n953bar), .A2(n952bar), .ZN(n958bar);
  OR2_X1 U17 ( .A1(in_58), .A2(in_4), .ZN(n952) );
  AND2_X1 U17bar ( .A1(in_58bar), .A2(in_4bar), .ZN(n952bar);
  OR2_X1 U18 ( .A1(in_59), .A2(n951), .ZN(n953) );
  AND2_X1 U18bar ( .A1(in_59bar), .A2(n951bar), .ZN(n953bar);
  OR2_X1 U19 ( .A1(in_71), .A2(in_62), .ZN(n951) );
  AND2_X1 U19bar ( .A1(in_71bar), .A2(in_62bar), .ZN(n951bar);
  OR2_X1 U20 ( .A1(n950), .A2(n949), .ZN(out[6]) );
  AND2_X1 U20bar ( .A1(n950bar), .A2(n949bar), .ZN(outbar[6]);
  OR2_X1 U21 ( .A1(n948), .A2(n947), .ZN(n949) );
  AND2_X1 U21bar ( .A1(n948bar), .A2(n947bar), .ZN(n949bar);
  OR2_X1 U22 ( .A1(n946), .A2(n945), .ZN(n947) );
  AND2_X1 U22bar ( .A1(n946bar), .A2(n945bar), .ZN(n947bar);
  OR2_X1 U23 ( .A1(n944), .A2(n943), .ZN(n945) );
  AND2_X1 U23bar ( .A1(n944bar), .A2(n943bar), .ZN(n945bar);
  OR2_X1 U24 ( .A1(n942), .A2(n941), .ZN(n946) );
  AND2_X1 U24bar ( .A1(n942bar), .A2(n941bar), .ZN(n946bar);
  OR2_X1 U25 ( .A1(in[101]), .A2(n940), .ZN(n941) );
  AND2_X1 U25bar ( .A1(inbar[101]), .A2(n940bar), .ZN(n941bar);
  OR2_X1 U26 ( .A1(n939), .A2(n938), .ZN(n948) );
  AND2_X1 U26bar ( .A1(n939bar), .A2(n938bar), .ZN(n948bar);
  OR2_X1 U27 ( .A1(in[114]), .A2(in[104]), .ZN(n938) );
  AND2_X1 U27bar ( .A1(inbar[114]), .A2(inbar[104]), .ZN(n938bar);
  OR2_X1 U28 ( .A1(in[128]), .A2(n937), .ZN(n939) );
  AND2_X1 U28bar ( .A1(inbar[128]), .A2(n937bar), .ZN(n939bar);
  OR2_X1 U29 ( .A1(in[136]), .A2(in[134]), .ZN(n937) );
  AND2_X1 U29bar ( .A1(inbar[136]), .A2(inbar[134]), .ZN(n937bar);
  OR2_X1 U30 ( .A1(n936), .A2(n935), .ZN(n950) );
  AND2_X1 U30bar ( .A1(n936bar), .A2(n935bar), .ZN(n950bar);
  OR2_X1 U31 ( .A1(n934), .A2(n933), .ZN(n935) );
  AND2_X1 U31bar ( .A1(n934bar), .A2(n933bar), .ZN(n935bar);
  OR2_X1 U32 ( .A1(in[177]), .A2(in[164]), .ZN(n933) );
  AND2_X1 U32bar ( .A1(inbar[177]), .A2(inbar[164]), .ZN(n933bar);
  OR2_X1 U33 ( .A1(in[212]), .A2(n932), .ZN(n934) );
  AND2_X1 U33bar ( .A1(inbar[212]), .A2(n932bar), .ZN(n934bar);
  OR2_X1 U34 ( .A1(in[248]), .A2(in[221]), .ZN(n932) );
  AND2_X1 U34bar ( .A1(inbar[248]), .A2(inbar[221]), .ZN(n932bar);
  OR2_X1 U35 ( .A1(n931), .A2(n930), .ZN(n936) );
  AND2_X1 U35bar ( .A1(n931bar), .A2(n930bar), .ZN(n936bar);
  OR2_X1 U36 ( .A1(in_18), .A2(in[93]), .ZN(n930) );
  AND2_X1 U36bar ( .A1(in_18bar), .A2(inbar[93]), .ZN(n930bar);
  OR2_X1 U37 ( .A1(in_31), .A2(n929), .ZN(n931) );
  AND2_X1 U37bar ( .A1(in_31bar), .A2(n929bar), .ZN(n931bar);
  OR2_X1 U38 ( .A1(in_7), .A2(in_39), .ZN(n929) );
  AND2_X1 U38bar ( .A1(in_7bar), .A2(in_39bar), .ZN(n929bar);
  OR2_X1 U39 ( .A1(n928), .A2(n927), .ZN(out[5]) );
  AND2_X1 U39bar ( .A1(n928bar), .A2(n927bar), .ZN(outbar[5]);
  OR2_X1 U40 ( .A1(n926), .A2(n925), .ZN(n927) );
  AND2_X1 U40bar ( .A1(n926bar), .A2(n925bar), .ZN(n927bar);
  OR2_X1 U41 ( .A1(n924), .A2(n923), .ZN(n925) );
  AND2_X1 U41bar ( .A1(n924bar), .A2(n923bar), .ZN(n925bar);
  OR2_X1 U42 ( .A1(n922), .A2(n921), .ZN(n923) );
  AND2_X1 U42bar ( .A1(n922bar), .A2(n921bar), .ZN(n923bar);
  OR2_X1 U43 ( .A1(n940), .A2(n920), .ZN(n924) );
  AND2_X1 U43bar ( .A1(n940bar), .A2(n920bar), .ZN(n924bar);
  OR2_X1 U44 ( .A1(in[111]), .A2(n919), .ZN(n920) );
  AND2_X1 U44bar ( .A1(inbar[111]), .A2(n919bar), .ZN(n920bar);
  OR2_X1 U45 ( .A1(n918), .A2(n917), .ZN(n940) );
  AND2_X1 U45bar ( .A1(n918bar), .A2(n917bar), .ZN(n940bar);
  OR2_X1 U46 ( .A1(n916), .A2(n915), .ZN(n917) );
  AND2_X1 U46bar ( .A1(n916bar), .A2(n915bar), .ZN(n917bar);
  OR2_X1 U47 ( .A1(n914), .A2(n913), .ZN(n915) );
  AND2_X1 U47bar ( .A1(n914bar), .A2(n913bar), .ZN(n915bar);
  OR2_X1 U48 ( .A1(in[140]), .A2(in[131]), .ZN(n913) );
  AND2_X1 U48bar ( .A1(inbar[140]), .A2(inbar[131]), .ZN(n913bar);
  OR2_X1 U49 ( .A1(in[160]), .A2(in[144]), .ZN(n914) );
  AND2_X1 U49bar ( .A1(inbar[160]), .A2(inbar[144]), .ZN(n914bar);
  OR2_X1 U50 ( .A1(n912), .A2(n911), .ZN(n916) );
  AND2_X1 U50bar ( .A1(n912bar), .A2(n911bar), .ZN(n916bar);
  OR2_X1 U51 ( .A1(in[179]), .A2(in[174]), .ZN(n911) );
  AND2_X1 U51bar ( .A1(inbar[179]), .A2(inbar[174]), .ZN(n911bar);
  OR2_X1 U52 ( .A1(in[188]), .A2(in[184]), .ZN(n912) );
  AND2_X1 U52bar ( .A1(inbar[188]), .A2(inbar[184]), .ZN(n912bar);
  OR2_X1 U53 ( .A1(n910), .A2(n909), .ZN(n918) );
  AND2_X1 U53bar ( .A1(n910bar), .A2(n909bar), .ZN(n918bar);
  OR2_X1 U54 ( .A1(n908), .A2(n907), .ZN(n909) );
  AND2_X1 U54bar ( .A1(n908bar), .A2(n907bar), .ZN(n909bar);
  OR2_X1 U55 ( .A1(in[216]), .A2(in[200]), .ZN(n907) );
  AND2_X1 U55bar ( .A1(inbar[216]), .A2(inbar[200]), .ZN(n907bar);
  OR2_X1 U56 ( .A1(in[228]), .A2(in[224]), .ZN(n908) );
  AND2_X1 U56bar ( .A1(inbar[228]), .A2(inbar[224]), .ZN(n908bar);
  OR2_X1 U57 ( .A1(n906), .A2(n905), .ZN(n910) );
  AND2_X1 U57bar ( .A1(n906bar), .A2(n905bar), .ZN(n910bar);
  OR2_X1 U58 ( .A1(in[247]), .A2(in[235]), .ZN(n905) );
  AND2_X1 U58bar ( .A1(inbar[247]), .A2(inbar[235]), .ZN(n905bar);
  OR2_X1 U59 ( .A1(in_42), .A2(in[83]), .ZN(n906) );
  AND2_X1 U59bar ( .A1(in_42bar), .A2(inbar[83]), .ZN(n906bar);
  OR2_X1 U60 ( .A1(n904), .A2(n903), .ZN(n926) );
  AND2_X1 U60bar ( .A1(n904bar), .A2(n903bar), .ZN(n926bar);
  OR2_X1 U61 ( .A1(in[166]), .A2(in[123]), .ZN(n903) );
  AND2_X1 U61bar ( .A1(inbar[166]), .A2(inbar[123]), .ZN(n903bar);
  OR2_X1 U62 ( .A1(in[170]), .A2(n902), .ZN(n904) );
  AND2_X1 U62bar ( .A1(inbar[170]), .A2(n902bar), .ZN(n904bar);
  OR2_X1 U63 ( .A1(in[194]), .A2(in[183]), .ZN(n902) );
  AND2_X1 U63bar ( .A1(inbar[194]), .A2(inbar[183]), .ZN(n902bar);
  OR2_X1 U64 ( .A1(n901), .A2(n900), .ZN(n928) );
  AND2_X1 U64bar ( .A1(n901bar), .A2(n900bar), .ZN(n928bar);
  OR2_X1 U65 ( .A1(n899), .A2(n898), .ZN(n900) );
  AND2_X1 U65bar ( .A1(n899bar), .A2(n898bar), .ZN(n900bar);
  OR2_X1 U66 ( .A1(in[241]), .A2(in[238]), .ZN(n898) );
  AND2_X1 U66bar ( .A1(inbar[241]), .A2(inbar[238]), .ZN(n898bar);
  OR2_X1 U67 ( .A1(in[250]), .A2(n897), .ZN(n899) );
  AND2_X1 U67bar ( .A1(inbar[250]), .A2(n897bar), .ZN(n899bar);
  OR2_X1 U68 ( .A1(in_24), .A2(in[84]), .ZN(n897) );
  AND2_X1 U68bar ( .A1(in_24bar), .A2(inbar[84]), .ZN(n897bar);
  OR2_X1 U69 ( .A1(n896), .A2(n895), .ZN(n901) );
  AND2_X1 U69bar ( .A1(n896bar), .A2(n895bar), .ZN(n901bar);
  OR2_X1 U70 ( .A1(in_41), .A2(in_29), .ZN(n895) );
  AND2_X1 U70bar ( .A1(in_41bar), .A2(in_29bar), .ZN(n895bar);
  OR2_X1 U71 ( .A1(in_66), .A2(n894), .ZN(n896) );
  AND2_X1 U71bar ( .A1(in_66bar), .A2(n894bar), .ZN(n896bar);
  OR2_X1 U72 ( .A1(in_76), .A2(in_71), .ZN(n894) );
  AND2_X1 U72bar ( .A1(in_76bar), .A2(in_71bar), .ZN(n894bar);
  OR2_X1 U73 ( .A1(n893), .A2(n892), .ZN(out[4]) );
  AND2_X1 U73bar ( .A1(n893bar), .A2(n892bar), .ZN(outbar[4]);
  OR2_X1 U74 ( .A1(n891), .A2(n890), .ZN(n892) );
  AND2_X1 U74bar ( .A1(n891bar), .A2(n890bar), .ZN(n892bar);
  OR2_X1 U75 ( .A1(n889), .A2(n888), .ZN(n890) );
  AND2_X1 U75bar ( .A1(n889bar), .A2(n888bar), .ZN(n890bar);
  OR2_X1 U76 ( .A1(n922), .A2(n887), .ZN(n888) );
  AND2_X1 U76bar ( .A1(n922bar), .A2(n887bar), .ZN(n888bar);
  OR2_X1 U77 ( .A1(n886), .A2(n885), .ZN(n922) );
  AND2_X1 U77bar ( .A1(n886bar), .A2(n885bar), .ZN(n922bar);
  OR2_X1 U78 ( .A1(n884), .A2(n883), .ZN(n885) );
  AND2_X1 U78bar ( .A1(n884bar), .A2(n883bar), .ZN(n885bar);
  OR2_X1 U79 ( .A1(n882), .A2(n881), .ZN(n883) );
  AND2_X1 U79bar ( .A1(n882bar), .A2(n881bar), .ZN(n883bar);
  OR2_X1 U80 ( .A1(in[118]), .A2(in[109]), .ZN(n881) );
  AND2_X1 U80bar ( .A1(inbar[118]), .A2(inbar[109]), .ZN(n881bar);
  OR2_X1 U81 ( .A1(in[139]), .A2(in[120]), .ZN(n882) );
  AND2_X1 U81bar ( .A1(inbar[139]), .A2(inbar[120]), .ZN(n882bar);
  OR2_X1 U82 ( .A1(n880), .A2(n879), .ZN(n884) );
  AND2_X1 U82bar ( .A1(n880bar), .A2(n879bar), .ZN(n884bar);
  OR2_X1 U83 ( .A1(in[198]), .A2(in[154]), .ZN(n879) );
  AND2_X1 U83bar ( .A1(inbar[198]), .A2(inbar[154]), .ZN(n879bar);
  OR2_X1 U84 ( .A1(in[210]), .A2(in[205]), .ZN(n880) );
  AND2_X1 U84bar ( .A1(inbar[210]), .A2(inbar[205]), .ZN(n880bar);
  OR2_X1 U85 ( .A1(n878), .A2(n877), .ZN(n886) );
  AND2_X1 U85bar ( .A1(n878bar), .A2(n877bar), .ZN(n886bar);
  OR2_X1 U86 ( .A1(n876), .A2(n875), .ZN(n877) );
  AND2_X1 U86bar ( .A1(n876bar), .A2(n875bar), .ZN(n877bar);
  OR2_X1 U87 ( .A1(in[219]), .A2(in[217]), .ZN(n875) );
  AND2_X1 U87bar ( .A1(inbar[219]), .A2(inbar[217]), .ZN(n875bar);
  OR2_X1 U88 ( .A1(in[86]), .A2(in[252]), .ZN(n876) );
  AND2_X1 U88bar ( .A1(inbar[86]), .A2(inbar[252]), .ZN(n876bar);
  OR2_X1 U89 ( .A1(n874), .A2(n873), .ZN(n878) );
  AND2_X1 U89bar ( .A1(n874bar), .A2(n873bar), .ZN(n878bar);
  OR2_X1 U90 ( .A1(in_40), .A2(in[91]), .ZN(n873) );
  AND2_X1 U90bar ( .A1(in_40bar), .A2(inbar[91]), .ZN(n873bar);
  OR2_X1 U91 ( .A1(in_8), .A2(in_46), .ZN(n874) );
  AND2_X1 U91bar ( .A1(in_8bar), .A2(in_46bar), .ZN(n874bar);
  OR2_X1 U92 ( .A1(n872), .A2(n871), .ZN(n889) );
  AND2_X1 U92bar ( .A1(n872bar), .A2(n871bar), .ZN(n889bar);
  OR2_X1 U93 ( .A1(in[117]), .A2(n943), .ZN(n871) );
  AND2_X1 U93bar ( .A1(inbar[117]), .A2(n943bar), .ZN(n871bar);
  OR2_X1 U94 ( .A1(n870), .A2(n869), .ZN(n943) );
  AND2_X1 U94bar ( .A1(n870bar), .A2(n869bar), .ZN(n943bar);
  OR2_X1 U95 ( .A1(n868), .A2(n867), .ZN(n869) );
  AND2_X1 U95bar ( .A1(n868bar), .A2(n867bar), .ZN(n869bar);
  OR2_X1 U96 ( .A1(n866), .A2(n865), .ZN(n867) );
  AND2_X1 U96bar ( .A1(n866bar), .A2(n865bar), .ZN(n867bar);
  OR2_X1 U97 ( .A1(n864), .A2(n863), .ZN(n865) );
  AND2_X1 U97bar ( .A1(n864bar), .A2(n863bar), .ZN(n865bar);
  OR2_X1 U98 ( .A1(in[108]), .A2(n919), .ZN(n866) );
  AND2_X1 U98bar ( .A1(inbar[108]), .A2(n919bar), .ZN(n866bar);
  OR2_X1 U99 ( .A1(n862), .A2(n861), .ZN(n919) );
  AND2_X1 U99bar ( .A1(n862bar), .A2(n861bar), .ZN(n919bar);
  OR2_X1 U100 ( .A1(n860), .A2(n859), .ZN(n861) );
  AND2_X1 U100bar ( .A1(n860bar), .A2(n859bar), .ZN(n861bar);
  OR2_X1 U101 ( .A1(n858), .A2(n857), .ZN(n859) );
  AND2_X1 U101bar ( .A1(n858bar), .A2(n857bar), .ZN(n859bar);
  OR2_X1 U102 ( .A1(in[119]), .A2(in[105]), .ZN(n857) );
  AND2_X1 U102bar ( .A1(inbar[119]), .A2(inbar[105]), .ZN(n857bar);
  OR2_X1 U103 ( .A1(in[186]), .A2(in[175]), .ZN(n858) );
  AND2_X1 U103bar ( .A1(inbar[186]), .A2(inbar[175]), .ZN(n858bar);
  OR2_X1 U104 ( .A1(n856), .A2(n855), .ZN(n860) );
  AND2_X1 U104bar ( .A1(n856bar), .A2(n855bar), .ZN(n860bar);
  OR2_X1 U105 ( .A1(in[202]), .A2(in[193]), .ZN(n855) );
  AND2_X1 U105bar ( .A1(inbar[202]), .A2(inbar[193]), .ZN(n855bar);
  OR2_X1 U106 ( .A1(in[225]), .A2(in[208]), .ZN(n856) );
  AND2_X1 U106bar ( .A1(inbar[225]), .A2(inbar[208]), .ZN(n856bar);
  OR2_X1 U107 ( .A1(n854), .A2(n853), .ZN(n862) );
  AND2_X1 U107bar ( .A1(n854bar), .A2(n853bar), .ZN(n862bar);
  OR2_X1 U108 ( .A1(n852), .A2(n851), .ZN(n853) );
  AND2_X1 U108bar ( .A1(n852bar), .A2(n851bar), .ZN(n853bar);
  OR2_X1 U109 ( .A1(in_1), .A2(in[85]), .ZN(n851) );
  AND2_X1 U109bar ( .A1(in_1bar), .A2(inbar[85]), .ZN(n851bar);
  OR2_X1 U110 ( .A1(in_23), .A2(in_19), .ZN(n852) );
  AND2_X1 U110bar ( .A1(in_23bar), .A2(in_19bar), .ZN(n852bar);
  OR2_X1 U111 ( .A1(n850), .A2(n849), .ZN(n854) );
  AND2_X1 U111bar ( .A1(n850bar), .A2(n849bar), .ZN(n854bar);
  OR2_X1 U112 ( .A1(in_43), .A2(in_33), .ZN(n849) );
  AND2_X1 U112bar ( .A1(in_43bar), .A2(in_33bar), .ZN(n849bar);
  OR2_X1 U113 ( .A1(in_63), .A2(in_44), .ZN(n850) );
  AND2_X1 U113bar ( .A1(in_63bar), .A2(in_44bar), .ZN(n850bar);
  OR2_X1 U114 ( .A1(n848), .A2(n847), .ZN(n868) );
  AND2_X1 U114bar ( .A1(n848bar), .A2(n847bar), .ZN(n868bar);
  OR2_X1 U115 ( .A1(in[141]), .A2(in[112]), .ZN(n847) );
  AND2_X1 U115bar ( .A1(inbar[141]), .A2(inbar[112]), .ZN(n847bar);
  OR2_X1 U116 ( .A1(in[147]), .A2(n846), .ZN(n848) );
  AND2_X1 U116bar ( .A1(inbar[147]), .A2(n846bar), .ZN(n848bar);
  OR2_X1 U117 ( .A1(in[181]), .A2(in[167]), .ZN(n846) );
  AND2_X1 U117bar ( .A1(inbar[181]), .A2(inbar[167]), .ZN(n846bar);
  OR2_X1 U118 ( .A1(n845), .A2(n844), .ZN(n870) );
  AND2_X1 U118bar ( .A1(n845bar), .A2(n844bar), .ZN(n870bar);
  OR2_X1 U119 ( .A1(n843), .A2(n842), .ZN(n844) );
  AND2_X1 U119bar ( .A1(n843bar), .A2(n842bar), .ZN(n844bar);
  OR2_X1 U120 ( .A1(in[229]), .A2(in[201]), .ZN(n842) );
  AND2_X1 U120bar ( .A1(inbar[229]), .A2(inbar[201]), .ZN(n842bar);
  OR2_X1 U121 ( .A1(in[237]), .A2(n841), .ZN(n843) );
  AND2_X1 U121bar ( .A1(inbar[237]), .A2(n841bar), .ZN(n843bar);
  OR2_X1 U122 ( .A1(in[94]), .A2(in[253]), .ZN(n841) );
  AND2_X1 U122bar ( .A1(inbar[94]), .A2(inbar[253]), .ZN(n841bar);
  OR2_X1 U123 ( .A1(n840), .A2(n839), .ZN(n845) );
  AND2_X1 U123bar ( .A1(n840bar), .A2(n839bar), .ZN(n845bar);
  OR2_X1 U124 ( .A1(in_21), .A2(in[96]), .ZN(n839) );
  AND2_X1 U124bar ( .A1(in_21bar), .A2(inbar[96]), .ZN(n839bar);
  OR2_X1 U125 ( .A1(in_25), .A2(n838), .ZN(n840) );
  AND2_X1 U125bar ( .A1(in_25bar), .A2(n838bar), .ZN(n840bar);
  OR2_X1 U126 ( .A1(in_81), .A2(in_45), .ZN(n838) );
  AND2_X1 U126bar ( .A1(in_81bar), .A2(in_45bar), .ZN(n838bar);
  OR2_X1 U127 ( .A1(n837), .A2(n836), .ZN(n891) );
  AND2_X1 U127bar ( .A1(n837bar), .A2(n836bar), .ZN(n891bar);
  OR2_X1 U128 ( .A1(in[142]), .A2(in[124]), .ZN(n836) );
  AND2_X1 U128bar ( .A1(inbar[142]), .A2(inbar[124]), .ZN(n836bar);
  OR2_X1 U129 ( .A1(in[150]), .A2(n835), .ZN(n837) );
  AND2_X1 U129bar ( .A1(inbar[150]), .A2(n835bar), .ZN(n837bar);
  OR2_X1 U130 ( .A1(in[172]), .A2(in[155]), .ZN(n835) );
  AND2_X1 U130bar ( .A1(inbar[172]), .A2(inbar[155]), .ZN(n835bar);
  OR2_X1 U131 ( .A1(n834), .A2(n833), .ZN(n893) );
  AND2_X1 U131bar ( .A1(n834bar), .A2(n833bar), .ZN(n893bar);
  OR2_X1 U132 ( .A1(n832), .A2(n831), .ZN(n833) );
  AND2_X1 U132bar ( .A1(n832bar), .A2(n831bar), .ZN(n833bar);
  OR2_X1 U133 ( .A1(in[196]), .A2(in[173]), .ZN(n831) );
  AND2_X1 U133bar ( .A1(inbar[196]), .A2(inbar[173]), .ZN(n831bar);
  OR2_X1 U134 ( .A1(in[222]), .A2(n830), .ZN(n832) );
  AND2_X1 U134bar ( .A1(inbar[222]), .A2(n830bar), .ZN(n832bar);
  OR2_X1 U135 ( .A1(in[227]), .A2(in[226]), .ZN(n830) );
  AND2_X1 U135bar ( .A1(inbar[227]), .A2(inbar[226]), .ZN(n830bar);
  OR2_X1 U136 ( .A1(n829), .A2(n828), .ZN(n834) );
  AND2_X1 U136bar ( .A1(n829bar), .A2(n828bar), .ZN(n834bar);
  OR2_X1 U137 ( .A1(in[249]), .A2(in[231]), .ZN(n828) );
  AND2_X1 U137bar ( .A1(inbar[249]), .A2(inbar[231]), .ZN(n828bar);
  OR2_X1 U138 ( .A1(in_28), .A2(n827), .ZN(n829) );
  AND2_X1 U138bar ( .A1(in_28bar), .A2(n827bar), .ZN(n829bar);
  OR2_X1 U139 ( .A1(in_52), .A2(in_47), .ZN(n827) );
  AND2_X1 U139bar ( .A1(in_52bar), .A2(in_47bar), .ZN(n827bar);
  OR2_X1 U140 ( .A1(n826), .A2(n825), .ZN(out[3]) );
  AND2_X1 U140bar ( .A1(n826bar), .A2(n825bar), .ZN(outbar[3]);
  OR2_X1 U141 ( .A1(n824), .A2(n823), .ZN(n825) );
  AND2_X1 U141bar ( .A1(n824bar), .A2(n823bar), .ZN(n825bar);
  OR2_X1 U142 ( .A1(n822), .A2(n821), .ZN(n823) );
  AND2_X1 U142bar ( .A1(n822bar), .A2(n821bar), .ZN(n823bar);
  OR2_X1 U143 ( .A1(n820), .A2(n819), .ZN(n821) );
  AND2_X1 U143bar ( .A1(n820bar), .A2(n819bar), .ZN(n821bar);
  OR2_X1 U144 ( .A1(n964), .A2(n818), .ZN(n822) );
  AND2_X1 U144bar ( .A1(n964bar), .A2(n818bar), .ZN(n822bar);
  OR2_X1 U145 ( .A1(in[118]), .A2(n817), .ZN(n818) );
  AND2_X1 U145bar ( .A1(inbar[118]), .A2(n817bar), .ZN(n818bar);
  OR2_X1 U146 ( .A1(n816), .A2(n815), .ZN(n964) );
  AND2_X1 U146bar ( .A1(n816bar), .A2(n815bar), .ZN(n964bar);
  OR2_X1 U147 ( .A1(n814), .A2(n813), .ZN(n815) );
  AND2_X1 U147bar ( .A1(n814bar), .A2(n813bar), .ZN(n815bar);
  OR2_X1 U148 ( .A1(n812), .A2(n811), .ZN(n813) );
  AND2_X1 U148bar ( .A1(n812bar), .A2(n811bar), .ZN(n813bar);
  OR2_X1 U149 ( .A1(in[122]), .A2(in[111]), .ZN(n811) );
  AND2_X1 U149bar ( .A1(inbar[122]), .A2(inbar[111]), .ZN(n811bar);
  OR2_X1 U150 ( .A1(in[154]), .A2(in[151]), .ZN(n812) );
  AND2_X1 U150bar ( .A1(inbar[154]), .A2(inbar[151]), .ZN(n812bar);
  OR2_X1 U151 ( .A1(n810), .A2(n809), .ZN(n814) );
  AND2_X1 U151bar ( .A1(n810bar), .A2(n809bar), .ZN(n814bar);
  OR2_X1 U152 ( .A1(in[187]), .A2(in[177]), .ZN(n809) );
  AND2_X1 U152bar ( .A1(inbar[187]), .A2(inbar[177]), .ZN(n809bar);
  OR2_X1 U153 ( .A1(in[200]), .A2(in[192]), .ZN(n810) );
  AND2_X1 U153bar ( .A1(inbar[200]), .A2(inbar[192]), .ZN(n810bar);
  OR2_X1 U154 ( .A1(n808), .A2(n807), .ZN(n816) );
  AND2_X1 U154bar ( .A1(n808bar), .A2(n807bar), .ZN(n816bar);
  OR2_X1 U155 ( .A1(n806), .A2(n805), .ZN(n807) );
  AND2_X1 U155bar ( .A1(n806bar), .A2(n805bar), .ZN(n807bar);
  OR2_X1 U156 ( .A1(in[225]), .A2(in[207]), .ZN(n805) );
  AND2_X1 U156bar ( .A1(inbar[225]), .A2(inbar[207]), .ZN(n805bar);
  OR2_X1 U157 ( .A1(in[98]), .A2(in[226]), .ZN(n806) );
  AND2_X1 U157bar ( .A1(inbar[98]), .A2(inbar[226]), .ZN(n806bar);
  OR2_X1 U158 ( .A1(n804), .A2(n803), .ZN(n808) );
  AND2_X1 U158bar ( .A1(n804bar), .A2(n803bar), .ZN(n808bar);
  OR2_X1 U159 ( .A1(in_20), .A2(in_16), .ZN(n803) );
  AND2_X1 U159bar ( .A1(in_20bar), .A2(in_16bar), .ZN(n803bar);
  OR2_X1 U160 ( .A1(in_55), .A2(in_45), .ZN(n804) );
  AND2_X1 U160bar ( .A1(in_55bar), .A2(in_45bar), .ZN(n804bar);
  OR2_X1 U161 ( .A1(n802), .A2(n801), .ZN(n824) );
  AND2_X1 U161bar ( .A1(n802bar), .A2(n801bar), .ZN(n824bar);
  OR2_X1 U162 ( .A1(in[162]), .A2(in[149]), .ZN(n801) );
  AND2_X1 U162bar ( .A1(inbar[162]), .A2(inbar[149]), .ZN(n801bar);
  OR2_X1 U163 ( .A1(in[163]), .A2(n800), .ZN(n802) );
  AND2_X1 U163bar ( .A1(inbar[163]), .A2(n800bar), .ZN(n802bar);
  OR2_X1 U164 ( .A1(in[191]), .A2(in[189]), .ZN(n800) );
  AND2_X1 U164bar ( .A1(inbar[191]), .A2(inbar[189]), .ZN(n800bar);
  OR2_X1 U165 ( .A1(n799), .A2(n798), .ZN(n826) );
  AND2_X1 U165bar ( .A1(n799bar), .A2(n798bar), .ZN(n826bar);
  OR2_X1 U166 ( .A1(n797), .A2(n796), .ZN(n798) );
  AND2_X1 U166bar ( .A1(n797bar), .A2(n796bar), .ZN(n798bar);
  OR2_X1 U167 ( .A1(in[212]), .A2(in[193]), .ZN(n796) );
  AND2_X1 U167bar ( .A1(inbar[212]), .A2(inbar[193]), .ZN(n796bar);
  OR2_X1 U168 ( .A1(in[238]), .A2(n795), .ZN(n797) );
  AND2_X1 U168bar ( .A1(inbar[238]), .A2(n795bar), .ZN(n797bar);
  OR2_X1 U169 ( .A1(in[88]), .A2(in[247]), .ZN(n795) );
  AND2_X1 U169bar ( .A1(inbar[88]), .A2(inbar[247]), .ZN(n795bar);
  OR2_X1 U170 ( .A1(n794), .A2(n793), .ZN(n799) );
  AND2_X1 U170bar ( .A1(n794bar), .A2(n793bar), .ZN(n799bar);
  OR2_X1 U171 ( .A1(in[94]), .A2(in[92]), .ZN(n793) );
  AND2_X1 U171bar ( .A1(inbar[94]), .A2(inbar[92]), .ZN(n793bar);
  OR2_X1 U172 ( .A1(in_52), .A2(n792), .ZN(n794) );
  AND2_X1 U172bar ( .A1(in_52bar), .A2(n792bar), .ZN(n794bar);
  OR2_X1 U173 ( .A1(in_70), .A2(in_67), .ZN(n792) );
  AND2_X1 U173bar ( .A1(in_70bar), .A2(in_67bar), .ZN(n792bar);
  OR2_X1 U174 ( .A1(n791), .A2(n790), .ZN(out[2]) );
  AND2_X1 U174bar ( .A1(n791bar), .A2(n790bar), .ZN(outbar[2]);
  OR2_X1 U175 ( .A1(n789), .A2(n788), .ZN(n790) );
  AND2_X1 U175bar ( .A1(n789bar), .A2(n788bar), .ZN(n790bar);
  OR2_X1 U176 ( .A1(n787), .A2(n786), .ZN(n788) );
  AND2_X1 U176bar ( .A1(n787bar), .A2(n786bar), .ZN(n788bar);
  OR2_X1 U177 ( .A1(n819), .A2(n785), .ZN(n786) );
  AND2_X1 U177bar ( .A1(n819bar), .A2(n785bar), .ZN(n786bar);
  OR2_X1 U178 ( .A1(n784), .A2(n783), .ZN(n819) );
  AND2_X1 U178bar ( .A1(n784bar), .A2(n783bar), .ZN(n819bar);
  OR2_X1 U179 ( .A1(n782), .A2(n781), .ZN(n783) );
  AND2_X1 U179bar ( .A1(n782bar), .A2(n781bar), .ZN(n783bar);
  OR2_X1 U180 ( .A1(n780), .A2(n779), .ZN(n781) );
  AND2_X1 U180bar ( .A1(n780bar), .A2(n779bar), .ZN(n781bar);
  OR2_X1 U181 ( .A1(n962), .A2(n778), .ZN(n779) );
  AND2_X1 U181bar ( .A1(n962bar), .A2(n778bar), .ZN(n779bar);
  OR2_X1 U182 ( .A1(n777), .A2(n776), .ZN(n962) );
  AND2_X1 U182bar ( .A1(n777bar), .A2(n776bar), .ZN(n962bar);
  OR2_X1 U183 ( .A1(n775), .A2(n774), .ZN(n776) );
  AND2_X1 U183bar ( .A1(n775bar), .A2(n774bar), .ZN(n776bar);
  OR2_X1 U184 ( .A1(n773), .A2(n772), .ZN(n774) );
  AND2_X1 U184bar ( .A1(n773bar), .A2(n772bar), .ZN(n774bar);
  OR2_X1 U185 ( .A1(in[131]), .A2(in[120]), .ZN(n772) );
  AND2_X1 U185bar ( .A1(inbar[131]), .A2(inbar[120]), .ZN(n772bar);
  OR2_X1 U186 ( .A1(in[153]), .A2(in[147]), .ZN(n773) );
  AND2_X1 U186bar ( .A1(inbar[153]), .A2(inbar[147]), .ZN(n773bar);
  OR2_X1 U187 ( .A1(n771), .A2(n770), .ZN(n775) );
  AND2_X1 U187bar ( .A1(n771bar), .A2(n770bar), .ZN(n775bar);
  OR2_X1 U188 ( .A1(in[170]), .A2(in[156]), .ZN(n770) );
  AND2_X1 U188bar ( .A1(inbar[170]), .A2(inbar[156]), .ZN(n770bar);
  OR2_X1 U189 ( .A1(in[223]), .A2(in[190]), .ZN(n771) );
  AND2_X1 U189bar ( .A1(inbar[223]), .A2(inbar[190]), .ZN(n771bar);
  OR2_X1 U190 ( .A1(n769), .A2(n768), .ZN(n777) );
  AND2_X1 U190bar ( .A1(n769bar), .A2(n768bar), .ZN(n777bar);
  OR2_X1 U191 ( .A1(n767), .A2(n766), .ZN(n768) );
  AND2_X1 U191bar ( .A1(n767bar), .A2(n766bar), .ZN(n768bar);
  OR2_X1 U192 ( .A1(in[236]), .A2(in[230]), .ZN(n766) );
  AND2_X1 U192bar ( .A1(inbar[236]), .A2(inbar[230]), .ZN(n766bar);
  OR2_X1 U193 ( .A1(in[85]), .A2(in[240]), .ZN(n767) );
  AND2_X1 U193bar ( .A1(inbar[85]), .A2(inbar[240]), .ZN(n767bar);
  OR2_X1 U194 ( .A1(n765), .A2(n764), .ZN(n769) );
  AND2_X1 U194bar ( .A1(n765bar), .A2(n764bar), .ZN(n769bar);
  OR2_X1 U195 ( .A1(in_12), .A2(in[90]), .ZN(n764) );
  AND2_X1 U195bar ( .A1(in_12bar), .A2(inbar[90]), .ZN(n764bar);
  OR2_X1 U196 ( .A1(in_39), .A2(in_28), .ZN(n765) );
  AND2_X1 U196bar ( .A1(in_39bar), .A2(in_28bar), .ZN(n765bar);
  OR2_X1 U197 ( .A1(in[109]), .A2(n763), .ZN(n780) );
  AND2_X1 U197bar ( .A1(inbar[109]), .A2(n763bar), .ZN(n780bar);
  OR2_X1 U198 ( .A1(n762), .A2(n761), .ZN(n782) );
  AND2_X1 U198bar ( .A1(n762bar), .A2(n761bar), .ZN(n782bar);
  OR2_X1 U199 ( .A1(in[138]), .A2(in[129]), .ZN(n761) );
  AND2_X1 U199bar ( .A1(inbar[138]), .A2(inbar[129]), .ZN(n761bar);
  OR2_X1 U200 ( .A1(in[157]), .A2(n760), .ZN(n762) );
  AND2_X1 U200bar ( .A1(inbar[157]), .A2(n760bar), .ZN(n762bar);
  OR2_X1 U201 ( .A1(in[182]), .A2(in[167]), .ZN(n760) );
  AND2_X1 U201bar ( .A1(inbar[182]), .A2(inbar[167]), .ZN(n760bar);
  OR2_X1 U202 ( .A1(n759), .A2(n758), .ZN(n784) );
  AND2_X1 U202bar ( .A1(n759bar), .A2(n758bar), .ZN(n784bar);
  OR2_X1 U203 ( .A1(n757), .A2(n756), .ZN(n758) );
  AND2_X1 U203bar ( .A1(n757bar), .A2(n756bar), .ZN(n758bar);
  OR2_X1 U204 ( .A1(in[195]), .A2(in[184]), .ZN(n756) );
  AND2_X1 U204bar ( .A1(inbar[195]), .A2(inbar[184]), .ZN(n756bar);
  OR2_X1 U205 ( .A1(in[196]), .A2(n755), .ZN(n757) );
  AND2_X1 U205bar ( .A1(inbar[196]), .A2(n755bar), .ZN(n757bar);
  OR2_X1 U206 ( .A1(in[215]), .A2(in[209]), .ZN(n755) );
  AND2_X1 U206bar ( .A1(inbar[215]), .A2(inbar[209]), .ZN(n755bar);
  OR2_X1 U207 ( .A1(n754), .A2(n753), .ZN(n759) );
  AND2_X1 U207bar ( .A1(n754bar), .A2(n753bar), .ZN(n759bar);
  OR2_X1 U208 ( .A1(in[93]), .A2(in[233]), .ZN(n753) );
  AND2_X1 U208bar ( .A1(inbar[93]), .A2(inbar[233]), .ZN(n753bar);
  OR2_X1 U209 ( .A1(in_1), .A2(n752), .ZN(n754) );
  AND2_X1 U209bar ( .A1(in_1bar), .A2(n752bar), .ZN(n754bar);
  OR2_X1 U210 ( .A1(in_69), .A2(in_66), .ZN(n752) );
  AND2_X1 U210bar ( .A1(in_69bar), .A2(in_66bar), .ZN(n752bar);
  OR2_X1 U211 ( .A1(n966), .A2(n751), .ZN(n787) );
  AND2_X1 U211bar ( .A1(n966bar), .A2(n751bar), .ZN(n787bar);
  OR2_X1 U212 ( .A1(in[134]), .A2(n750), .ZN(n751) );
  AND2_X1 U212bar ( .A1(inbar[134]), .A2(n750bar), .ZN(n751bar);
  OR2_X1 U213 ( .A1(n749), .A2(n748), .ZN(n966) );
  AND2_X1 U213bar ( .A1(n749bar), .A2(n748bar), .ZN(n966bar);
  OR2_X1 U214 ( .A1(n747), .A2(n746), .ZN(n748) );
  AND2_X1 U214bar ( .A1(n747bar), .A2(n746bar), .ZN(n748bar);
  OR2_X1 U215 ( .A1(n745), .A2(n744), .ZN(n746) );
  AND2_X1 U215bar ( .A1(n745bar), .A2(n744bar), .ZN(n746bar);
  OR2_X1 U216 ( .A1(in[136]), .A2(in[121]), .ZN(n744) );
  AND2_X1 U216bar ( .A1(inbar[136]), .A2(inbar[121]), .ZN(n744bar);
  OR2_X1 U217 ( .A1(in[186]), .A2(in[174]), .ZN(n745) );
  AND2_X1 U217bar ( .A1(inbar[186]), .A2(inbar[174]), .ZN(n745bar);
  OR2_X1 U218 ( .A1(n743), .A2(n742), .ZN(n747) );
  AND2_X1 U218bar ( .A1(n743bar), .A2(n742bar), .ZN(n747bar);
  OR2_X1 U219 ( .A1(in[198]), .A2(in[197]), .ZN(n742) );
  AND2_X1 U219bar ( .A1(inbar[198]), .A2(inbar[197]), .ZN(n742bar);
  OR2_X1 U220 ( .A1(in[214]), .A2(in[199]), .ZN(n743) );
  AND2_X1 U220bar ( .A1(inbar[214]), .A2(inbar[199]), .ZN(n743bar);
  OR2_X1 U221 ( .A1(n741), .A2(n740), .ZN(n749) );
  AND2_X1 U221bar ( .A1(n741bar), .A2(n740bar), .ZN(n749bar);
  OR2_X1 U222 ( .A1(n739), .A2(n738), .ZN(n740) );
  AND2_X1 U222bar ( .A1(n739bar), .A2(n738bar), .ZN(n740bar);
  OR2_X1 U223 ( .A1(in[231]), .A2(in[220]), .ZN(n738) );
  AND2_X1 U223bar ( .A1(inbar[231]), .A2(inbar[220]), .ZN(n738bar);
  OR2_X1 U224 ( .A1(in_25), .A2(in[245]), .ZN(n739) );
  AND2_X1 U224bar ( .A1(in_25bar), .A2(inbar[245]), .ZN(n739bar);
  OR2_X1 U225 ( .A1(n737), .A2(n736), .ZN(n741) );
  AND2_X1 U225bar ( .A1(n737bar), .A2(n736bar), .ZN(n741bar);
  OR2_X1 U226 ( .A1(in_53), .A2(in_29), .ZN(n736) );
  AND2_X1 U226bar ( .A1(in_53bar), .A2(in_29bar), .ZN(n736bar);
  OR2_X1 U227 ( .A1(in_79), .A2(in_74), .ZN(n737) );
  AND2_X1 U227bar ( .A1(in_79bar), .A2(in_74bar), .ZN(n737bar);
  OR2_X1 U228 ( .A1(n735), .A2(n734), .ZN(n789) );
  AND2_X1 U228bar ( .A1(n735bar), .A2(n734bar), .ZN(n789bar);
  OR2_X1 U229 ( .A1(in[152]), .A2(in[140]), .ZN(n734) );
  AND2_X1 U229bar ( .A1(inbar[152]), .A2(inbar[140]), .ZN(n734bar);
  OR2_X1 U230 ( .A1(in[155]), .A2(n733), .ZN(n735) );
  AND2_X1 U230bar ( .A1(inbar[155]), .A2(n733bar), .ZN(n735bar);
  OR2_X1 U231 ( .A1(in[166]), .A2(in[165]), .ZN(n733) );
  AND2_X1 U231bar ( .A1(inbar[166]), .A2(inbar[165]), .ZN(n733bar);
  OR2_X1 U232 ( .A1(n732), .A2(n731), .ZN(n791) );
  AND2_X1 U232bar ( .A1(n732bar), .A2(n731bar), .ZN(n791bar);
  OR2_X1 U233 ( .A1(n730), .A2(n729), .ZN(n731) );
  AND2_X1 U233bar ( .A1(n730bar), .A2(n729bar), .ZN(n731bar);
  OR2_X1 U234 ( .A1(in[202]), .A2(in[185]), .ZN(n729) );
  AND2_X1 U234bar ( .A1(inbar[202]), .A2(inbar[185]), .ZN(n729bar);
  OR2_X1 U235 ( .A1(in[211]), .A2(n728), .ZN(n730) );
  AND2_X1 U235bar ( .A1(inbar[211]), .A2(n728bar), .ZN(n730bar);
  OR2_X1 U236 ( .A1(in[255]), .A2(in[253]), .ZN(n728) );
  AND2_X1 U236bar ( .A1(inbar[255]), .A2(inbar[253]), .ZN(n728bar);
  OR2_X1 U237 ( .A1(n727), .A2(n726), .ZN(n732) );
  AND2_X1 U237bar ( .A1(n727bar), .A2(n726bar), .ZN(n732bar);
  OR2_X1 U238 ( .A1(in_35), .A2(in_15), .ZN(n726) );
  AND2_X1 U238bar ( .A1(in_35bar), .A2(in_15bar), .ZN(n726bar);
  OR2_X1 U239 ( .A1(in_36), .A2(n725), .ZN(n727) );
  AND2_X1 U239bar ( .A1(in_36bar), .A2(n725bar), .ZN(n727bar);
  OR2_X1 U240 ( .A1(in_48), .A2(in_40), .ZN(n725) );
  AND2_X1 U240bar ( .A1(in_48bar), .A2(in_40bar), .ZN(n725bar);
  OR2_X1 U241 ( .A1(n724), .A2(n723), .ZN(out[1]) );
  AND2_X1 U241bar ( .A1(n724bar), .A2(n723bar), .ZN(outbar[1]);
  OR2_X1 U242 ( .A1(n722), .A2(n721), .ZN(n723) );
  AND2_X1 U242bar ( .A1(n722bar), .A2(n721bar), .ZN(n723bar);
  OR2_X1 U243 ( .A1(n720), .A2(n719), .ZN(n721) );
  AND2_X1 U243bar ( .A1(n720bar), .A2(n719bar), .ZN(n721bar);
  OR2_X1 U244 ( .A1(n921), .A2(n887), .ZN(n719) );
  AND2_X1 U244bar ( .A1(n921bar), .A2(n887bar), .ZN(n719bar);
  OR2_X1 U245 ( .A1(n718), .A2(n717), .ZN(n887) );
  AND2_X1 U245bar ( .A1(n718bar), .A2(n717bar), .ZN(n887bar);
  OR2_X1 U246 ( .A1(n716), .A2(n715), .ZN(n717) );
  AND2_X1 U246bar ( .A1(n716bar), .A2(n715bar), .ZN(n717bar);
  OR2_X1 U247 ( .A1(n714), .A2(n713), .ZN(n715) );
  AND2_X1 U247bar ( .A1(n714bar), .A2(n713bar), .ZN(n715bar);
  OR2_X1 U248 ( .A1(in[116]), .A2(in[110]), .ZN(n713) );
  AND2_X1 U248bar ( .A1(inbar[116]), .A2(inbar[110]), .ZN(n713bar);
  OR2_X1 U249 ( .A1(in[133]), .A2(in[130]), .ZN(n714) );
  AND2_X1 U249bar ( .A1(inbar[133]), .A2(inbar[130]), .ZN(n714bar);
  OR2_X1 U250 ( .A1(n712), .A2(n711), .ZN(n716) );
  AND2_X1 U250bar ( .A1(n712bar), .A2(n711bar), .ZN(n716bar);
  OR2_X1 U251 ( .A1(in[203]), .A2(in[135]), .ZN(n711) );
  AND2_X1 U251bar ( .A1(inbar[203]), .A2(inbar[135]), .ZN(n711bar);
  OR2_X1 U252 ( .A1(in[232]), .A2(in[223]), .ZN(n712) );
  AND2_X1 U252bar ( .A1(inbar[232]), .A2(inbar[223]), .ZN(n712bar);
  OR2_X1 U253 ( .A1(n710), .A2(n709), .ZN(n718) );
  AND2_X1 U253bar ( .A1(n710bar), .A2(n709bar), .ZN(n718bar);
  OR2_X1 U254 ( .A1(n708), .A2(n707), .ZN(n709) );
  AND2_X1 U254bar ( .A1(n708bar), .A2(n707bar), .ZN(n709bar);
  OR2_X1 U255 ( .A1(in[255]), .A2(in[233]), .ZN(n707) );
  AND2_X1 U255bar ( .A1(inbar[255]), .A2(inbar[233]), .ZN(n707bar);
  OR2_X1 U256 ( .A1(in_53), .A2(in_34), .ZN(n708) );
  AND2_X1 U256bar ( .A1(in_53bar), .A2(in_34bar), .ZN(n708bar);
  OR2_X1 U257 ( .A1(n706), .A2(n705), .ZN(n710) );
  AND2_X1 U257bar ( .A1(n706bar), .A2(n705bar), .ZN(n710bar);
  OR2_X1 U258 ( .A1(in_57), .A2(in_55), .ZN(n705) );
  AND2_X1 U258bar ( .A1(in_57bar), .A2(in_55bar), .ZN(n705bar);
  OR2_X1 U259 ( .A1(in_68), .A2(in_67), .ZN(n706) );
  AND2_X1 U259bar ( .A1(in_68bar), .A2(in_67bar), .ZN(n706bar);
  OR2_X1 U260 ( .A1(n704), .A2(n703), .ZN(n921) );
  AND2_X1 U260bar ( .A1(n704bar), .A2(n703bar), .ZN(n921bar);
  OR2_X1 U261 ( .A1(n702), .A2(n701), .ZN(n703) );
  AND2_X1 U261bar ( .A1(n702bar), .A2(n701bar), .ZN(n703bar);
  OR2_X1 U262 ( .A1(n700), .A2(n699), .ZN(n701) );
  AND2_X1 U262bar ( .A1(n700bar), .A2(n699bar), .ZN(n701bar);
  OR2_X1 U263 ( .A1(n944), .A2(n872), .ZN(n699) );
  AND2_X1 U263bar ( .A1(n944bar), .A2(n872bar), .ZN(n699bar);
  OR2_X1 U264 ( .A1(n698), .A2(n697), .ZN(n872) );
  AND2_X1 U264bar ( .A1(n698bar), .A2(n697bar), .ZN(n872bar);
  OR2_X1 U265 ( .A1(n696), .A2(n695), .ZN(n697) );
  AND2_X1 U265bar ( .A1(n696bar), .A2(n695bar), .ZN(n697bar);
  OR2_X1 U266 ( .A1(n694), .A2(n693), .ZN(n695) );
  AND2_X1 U266bar ( .A1(n694bar), .A2(n693bar), .ZN(n695bar);
  OR2_X1 U267 ( .A1(in[121]), .A2(in[102]), .ZN(n693) );
  AND2_X1 U267bar ( .A1(inbar[121]), .A2(inbar[102]), .ZN(n693bar);
  OR2_X1 U268 ( .A1(in[162]), .A2(in[161]), .ZN(n694) );
  AND2_X1 U268bar ( .A1(inbar[162]), .A2(inbar[161]), .ZN(n694bar);
  OR2_X1 U269 ( .A1(n692), .A2(n691), .ZN(n696) );
  AND2_X1 U269bar ( .A1(n692bar), .A2(n691bar), .ZN(n696bar);
  OR2_X1 U270 ( .A1(in[192]), .A2(in[178]), .ZN(n691) );
  AND2_X1 U270bar ( .A1(inbar[192]), .A2(inbar[178]), .ZN(n691bar);
  OR2_X1 U271 ( .A1(in[244]), .A2(in[209]), .ZN(n692) );
  AND2_X1 U271bar ( .A1(inbar[244]), .A2(inbar[209]), .ZN(n692bar);
  OR2_X1 U272 ( .A1(n690), .A2(n689), .ZN(n698) );
  AND2_X1 U272bar ( .A1(n690bar), .A2(n689bar), .ZN(n698bar);
  OR2_X1 U273 ( .A1(n688), .A2(n687), .ZN(n689) );
  AND2_X1 U273bar ( .A1(n688bar), .A2(n687bar), .ZN(n689bar);
  OR2_X1 U274 ( .A1(in[90]), .A2(in[254]), .ZN(n687) );
  AND2_X1 U274bar ( .A1(inbar[90]), .A2(inbar[254]), .ZN(n687bar);
  OR2_X1 U275 ( .A1(in_36), .A2(in_32), .ZN(n688) );
  AND2_X1 U275bar ( .A1(in_36bar), .A2(in_32bar), .ZN(n688bar);
  OR2_X1 U276 ( .A1(n686), .A2(n685), .ZN(n690) );
  AND2_X1 U276bar ( .A1(n686bar), .A2(n685bar), .ZN(n690bar);
  OR2_X1 U277 ( .A1(in_62), .A2(in_37), .ZN(n685) );
  AND2_X1 U277bar ( .A1(in_62bar), .A2(in_37bar), .ZN(n685bar);
  OR2_X1 U278 ( .A1(in_75), .A2(in_73), .ZN(n686) );
  AND2_X1 U278bar ( .A1(in_75bar), .A2(in_73bar), .ZN(n686bar);
  OR2_X1 U279 ( .A1(n684), .A2(n683), .ZN(n944) );
  AND2_X1 U279bar ( .A1(n684bar), .A2(n683bar), .ZN(n944bar);
  OR2_X1 U280 ( .A1(n682), .A2(n681), .ZN(n683) );
  AND2_X1 U280bar ( .A1(n682bar), .A2(n681bar), .ZN(n683bar);
  OR2_X1 U281 ( .A1(n680), .A2(n679), .ZN(n681) );
  AND2_X1 U281bar ( .A1(n680bar), .A2(n679bar), .ZN(n681bar);
  OR2_X1 U282 ( .A1(in[171]), .A2(in[153]), .ZN(n679) );
  AND2_X1 U282bar ( .A1(inbar[171]), .A2(inbar[153]), .ZN(n679bar);
  OR2_X1 U283 ( .A1(in[187]), .A2(in[176]), .ZN(n680) );
  AND2_X1 U283bar ( .A1(inbar[187]), .A2(inbar[176]), .ZN(n680bar);
  OR2_X1 U284 ( .A1(n678), .A2(n677), .ZN(n682) );
  AND2_X1 U284bar ( .A1(n678bar), .A2(n677bar), .ZN(n682bar);
  OR2_X1 U285 ( .A1(in[245]), .A2(in[211]), .ZN(n677) );
  AND2_X1 U285bar ( .A1(inbar[245]), .A2(inbar[211]), .ZN(n677bar);
  OR2_X1 U286 ( .A1(in[97]), .A2(in[88]), .ZN(n678) );
  AND2_X1 U286bar ( .A1(inbar[97]), .A2(inbar[88]), .ZN(n678bar);
  OR2_X1 U287 ( .A1(n676), .A2(n675), .ZN(n684) );
  AND2_X1 U287bar ( .A1(n676bar), .A2(n675bar), .ZN(n684bar);
  OR2_X1 U288 ( .A1(n674), .A2(n673), .ZN(n675) );
  AND2_X1 U288bar ( .A1(n674bar), .A2(n673bar), .ZN(n675bar);
  OR2_X1 U289 ( .A1(in_10), .A2(in_0), .ZN(n673) );
  AND2_X1 U289bar ( .A1(in_10bar), .A2(in_0bar), .ZN(n673bar);
  OR2_X1 U290 ( .A1(in_59), .A2(in_5), .ZN(n674) );
  AND2_X1 U290bar ( .A1(in_59bar), .A2(in_5bar), .ZN(n674bar);
  OR2_X1 U291 ( .A1(n672), .A2(n671), .ZN(n676) );
  AND2_X1 U291bar ( .A1(n672bar), .A2(n671bar), .ZN(n676bar);
  OR2_X1 U292 ( .A1(in_60), .A2(in_6), .ZN(n671) );
  AND2_X1 U292bar ( .A1(in_60bar), .A2(in_6bar), .ZN(n671bar);
  OR2_X1 U293 ( .A1(in_77), .A2(in_69), .ZN(n672) );
  AND2_X1 U293bar ( .A1(in_77bar), .A2(in_69bar), .ZN(n672bar);
  OR2_X1 U294 ( .A1(in[113]), .A2(n864), .ZN(n700) );
  AND2_X1 U294bar ( .A1(inbar[113]), .A2(n864bar), .ZN(n700bar);
  OR2_X1 U295 ( .A1(n670), .A2(n669), .ZN(n864) );
  AND2_X1 U295bar ( .A1(n670bar), .A2(n669bar), .ZN(n864bar);
  OR2_X1 U296 ( .A1(n668), .A2(n667), .ZN(n669) );
  AND2_X1 U296bar ( .A1(n668bar), .A2(n667bar), .ZN(n669bar);
  OR2_X1 U297 ( .A1(n666), .A2(n665), .ZN(n667) );
  AND2_X1 U297bar ( .A1(n666bar), .A2(n665bar), .ZN(n667bar);
  OR2_X1 U298 ( .A1(in[125]), .A2(in[107]), .ZN(n665) );
  AND2_X1 U298bar ( .A1(inbar[125]), .A2(inbar[107]), .ZN(n665bar);
  OR2_X1 U299 ( .A1(in[138]), .A2(in[126]), .ZN(n666) );
  AND2_X1 U299bar ( .A1(inbar[138]), .A2(inbar[126]), .ZN(n666bar);
  OR2_X1 U300 ( .A1(n664), .A2(n663), .ZN(n668) );
  AND2_X1 U300bar ( .A1(n664bar), .A2(n663bar), .ZN(n668bar);
  OR2_X1 U301 ( .A1(in[189]), .A2(in[143]), .ZN(n663) );
  AND2_X1 U301bar ( .A1(inbar[189]), .A2(inbar[143]), .ZN(n663bar);
  OR2_X1 U302 ( .A1(in[99]), .A2(in[214]), .ZN(n664) );
  AND2_X1 U302bar ( .A1(inbar[99]), .A2(inbar[214]), .ZN(n664bar);
  OR2_X1 U303 ( .A1(n662), .A2(n661), .ZN(n670) );
  AND2_X1 U303bar ( .A1(n662bar), .A2(n661bar), .ZN(n670bar);
  OR2_X1 U304 ( .A1(n660), .A2(n659), .ZN(n661) );
  AND2_X1 U304bar ( .A1(n660bar), .A2(n659bar), .ZN(n661bar);
  OR2_X1 U305 ( .A1(in_15), .A2(in_12), .ZN(n659) );
  AND2_X1 U305bar ( .A1(in_15bar), .A2(in_12bar), .ZN(n659bar);
  OR2_X1 U306 ( .A1(in_20), .A2(in_2), .ZN(n660) );
  AND2_X1 U306bar ( .A1(in_20bar), .A2(in_2bar), .ZN(n660bar);
  OR2_X1 U307 ( .A1(n658), .A2(n657), .ZN(n662) );
  AND2_X1 U307bar ( .A1(n658bar), .A2(n657bar), .ZN(n662bar);
  OR2_X1 U308 ( .A1(in_30), .A2(in_3), .ZN(n657) );
  AND2_X1 U308bar ( .A1(in_30bar), .A2(in_3bar), .ZN(n657bar);
  OR2_X1 U309 ( .A1(in_4), .A2(in_38), .ZN(n658) );
  AND2_X1 U309bar ( .A1(in_4bar), .A2(in_38bar), .ZN(n658bar);
  OR2_X1 U310 ( .A1(n656), .A2(n655), .ZN(n702) );
  AND2_X1 U310bar ( .A1(n656bar), .A2(n655bar), .ZN(n702bar);
  OR2_X1 U311 ( .A1(in[148]), .A2(in[137]), .ZN(n655) );
  AND2_X1 U311bar ( .A1(inbar[148]), .A2(inbar[137]), .ZN(n655bar);
  OR2_X1 U312 ( .A1(in[149]), .A2(n654), .ZN(n656) );
  AND2_X1 U312bar ( .A1(inbar[149]), .A2(n654bar), .ZN(n656bar);
  OR2_X1 U313 ( .A1(in[195]), .A2(in[190]), .ZN(n654) );
  AND2_X1 U313bar ( .A1(inbar[195]), .A2(inbar[190]), .ZN(n654bar);
  OR2_X1 U314 ( .A1(n653), .A2(n652), .ZN(n704) );
  AND2_X1 U314bar ( .A1(n653bar), .A2(n652bar), .ZN(n704bar);
  OR2_X1 U315 ( .A1(n651), .A2(n650), .ZN(n652) );
  AND2_X1 U315bar ( .A1(n651bar), .A2(n650bar), .ZN(n652bar);
  OR2_X1 U316 ( .A1(in[98]), .A2(in[197]), .ZN(n650) );
  AND2_X1 U316bar ( .A1(inbar[98]), .A2(inbar[197]), .ZN(n650bar);
  OR2_X1 U317 ( .A1(in_11), .A2(n649), .ZN(n651) );
  AND2_X1 U317bar ( .A1(in_11bar), .A2(n649bar), .ZN(n651bar);
  OR2_X1 U318 ( .A1(in_26), .A2(in_14), .ZN(n649) );
  AND2_X1 U318bar ( .A1(in_26bar), .A2(in_14bar), .ZN(n649bar);
  OR2_X1 U319 ( .A1(n648), .A2(n647), .ZN(n653) );
  AND2_X1 U319bar ( .A1(n648bar), .A2(n647bar), .ZN(n653bar);
  OR2_X1 U320 ( .A1(in_35), .A2(in_27), .ZN(n647) );
  AND2_X1 U320bar ( .A1(in_35bar), .A2(in_27bar), .ZN(n647bar);
  OR2_X1 U321 ( .A1(in_50), .A2(n646), .ZN(n648) );
  AND2_X1 U321bar ( .A1(in_50bar), .A2(n646bar), .ZN(n648bar);
  OR2_X1 U322 ( .A1(in_78), .A2(in_61), .ZN(n646) );
  AND2_X1 U322bar ( .A1(in_78bar), .A2(in_61bar), .ZN(n646bar);
  OR2_X1 U323 ( .A1(n942), .A2(n645), .ZN(n720) );
  AND2_X1 U323bar ( .A1(n942bar), .A2(n645bar), .ZN(n720bar);
  OR2_X1 U324 ( .A1(in[106]), .A2(n863), .ZN(n645) );
  AND2_X1 U324bar ( .A1(inbar[106]), .A2(n863bar), .ZN(n645bar);
  OR2_X1 U325 ( .A1(n644), .A2(n643), .ZN(n863) );
  AND2_X1 U325bar ( .A1(n644bar), .A2(n643bar), .ZN(n863bar);
  OR2_X1 U326 ( .A1(n642), .A2(n641), .ZN(n643) );
  AND2_X1 U326bar ( .A1(n642bar), .A2(n641bar), .ZN(n643bar);
  OR2_X1 U327 ( .A1(n640), .A2(n639), .ZN(n641) );
  AND2_X1 U327bar ( .A1(n640bar), .A2(n639bar), .ZN(n641bar);
  OR2_X1 U328 ( .A1(in[127]), .A2(in[122]), .ZN(n639) );
  AND2_X1 U328bar ( .A1(inbar[127]), .A2(inbar[122]), .ZN(n639bar);
  OR2_X1 U329 ( .A1(in[156]), .A2(in[132]), .ZN(n640) );
  AND2_X1 U329bar ( .A1(inbar[156]), .A2(inbar[132]), .ZN(n640bar);
  OR2_X1 U330 ( .A1(n638), .A2(n637), .ZN(n642) );
  AND2_X1 U330bar ( .A1(n638bar), .A2(n637bar), .ZN(n642bar);
  OR2_X1 U331 ( .A1(in[159]), .A2(in[157]), .ZN(n637) );
  AND2_X1 U331bar ( .A1(inbar[159]), .A2(inbar[157]), .ZN(n637bar);
  OR2_X1 U332 ( .A1(in[185]), .A2(in[169]), .ZN(n638) );
  AND2_X1 U332bar ( .A1(inbar[185]), .A2(inbar[169]), .ZN(n638bar);
  OR2_X1 U333 ( .A1(n636), .A2(n635), .ZN(n644) );
  AND2_X1 U333bar ( .A1(n636bar), .A2(n635bar), .ZN(n644bar);
  OR2_X1 U334 ( .A1(n634), .A2(n633), .ZN(n635) );
  AND2_X1 U334bar ( .A1(n634bar), .A2(n633bar), .ZN(n635bar);
  OR2_X1 U335 ( .A1(in[239]), .A2(in[218]), .ZN(n633) );
  AND2_X1 U335bar ( .A1(inbar[239]), .A2(inbar[218]), .ZN(n633bar);
  OR2_X1 U336 ( .A1(in_13), .A2(in[87]), .ZN(n634) );
  AND2_X1 U336bar ( .A1(in_13bar), .A2(inbar[87]), .ZN(n634bar);
  OR2_X1 U337 ( .A1(n632), .A2(n631), .ZN(n636) );
  AND2_X1 U337bar ( .A1(n632bar), .A2(n631bar), .ZN(n636bar);
  OR2_X1 U338 ( .A1(in_72), .A2(in_70), .ZN(n631) );
  AND2_X1 U338bar ( .A1(in_72bar), .A2(in_70bar), .ZN(n631bar);
  OR2_X1 U339 ( .A1(in_80), .A2(in_74), .ZN(n632) );
  AND2_X1 U339bar ( .A1(in_80bar), .A2(in_74bar), .ZN(n632bar);
  OR2_X1 U340 ( .A1(n630), .A2(n629), .ZN(n942) );
  AND2_X1 U340bar ( .A1(n630bar), .A2(n629bar), .ZN(n942bar);
  OR2_X1 U341 ( .A1(n628), .A2(n627), .ZN(n629) );
  AND2_X1 U341bar ( .A1(n628bar), .A2(n627bar), .ZN(n629bar);
  OR2_X1 U342 ( .A1(n626), .A2(n625), .ZN(n627) );
  AND2_X1 U342bar ( .A1(n626bar), .A2(n625bar), .ZN(n627bar);
  OR2_X1 U343 ( .A1(in[146]), .A2(in[100]), .ZN(n625) );
  AND2_X1 U343bar ( .A1(inbar[146]), .A2(inbar[100]), .ZN(n625bar);
  OR2_X1 U344 ( .A1(in[168]), .A2(in[152]), .ZN(n626) );
  AND2_X1 U344bar ( .A1(inbar[168]), .A2(inbar[152]), .ZN(n626bar);
  OR2_X1 U345 ( .A1(n624), .A2(n623), .ZN(n628) );
  AND2_X1 U345bar ( .A1(n624bar), .A2(n623bar), .ZN(n628bar);
  OR2_X1 U346 ( .A1(in[199]), .A2(in[182]), .ZN(n623) );
  AND2_X1 U346bar ( .A1(inbar[199]), .A2(inbar[182]), .ZN(n623bar);
  OR2_X1 U347 ( .A1(in[236]), .A2(in[204]), .ZN(n624) );
  AND2_X1 U347bar ( .A1(inbar[236]), .A2(inbar[204]), .ZN(n624bar);
  OR2_X1 U348 ( .A1(n622), .A2(n621), .ZN(n630) );
  AND2_X1 U348bar ( .A1(n622bar), .A2(n621bar), .ZN(n630bar);
  OR2_X1 U349 ( .A1(n620), .A2(n619), .ZN(n621) );
  AND2_X1 U349bar ( .A1(n620bar), .A2(n619bar), .ZN(n621bar);
  OR2_X1 U350 ( .A1(in[89]), .A2(in[246]), .ZN(n619) );
  AND2_X1 U350bar ( .A1(inbar[89]), .A2(inbar[246]), .ZN(n619bar);
  OR2_X1 U351 ( .A1(in[95]), .A2(in[92]), .ZN(n620) );
  AND2_X1 U351bar ( .A1(inbar[95]), .A2(inbar[92]), .ZN(n620bar);
  OR2_X1 U352 ( .A1(n618), .A2(n617), .ZN(n622) );
  AND2_X1 U352bar ( .A1(n618bar), .A2(n617bar), .ZN(n622bar);
  OR2_X1 U353 ( .A1(in_22), .A2(in_16), .ZN(n617) );
  AND2_X1 U353bar ( .A1(in_22bar), .A2(in_16bar), .ZN(n617bar);
  OR2_X1 U354 ( .A1(in_51), .A2(in_49), .ZN(n618) );
  AND2_X1 U354bar ( .A1(in_51bar), .A2(in_49bar), .ZN(n618bar);
  OR2_X1 U355 ( .A1(n616), .A2(n615), .ZN(n722) );
  AND2_X1 U355bar ( .A1(n616bar), .A2(n615bar), .ZN(n722bar);
  OR2_X1 U356 ( .A1(in[158]), .A2(in[115]), .ZN(n615) );
  AND2_X1 U356bar ( .A1(inbar[158]), .A2(inbar[115]), .ZN(n615bar);
  OR2_X1 U357 ( .A1(in[163]), .A2(n614), .ZN(n616) );
  AND2_X1 U357bar ( .A1(inbar[163]), .A2(n614bar), .ZN(n616bar);
  OR2_X1 U358 ( .A1(in[206]), .A2(in[165]), .ZN(n614) );
  AND2_X1 U358bar ( .A1(inbar[206]), .A2(inbar[165]), .ZN(n614bar);
  OR2_X1 U359 ( .A1(n613), .A2(n612), .ZN(n724) );
  AND2_X1 U359bar ( .A1(n613bar), .A2(n612bar), .ZN(n724bar);
  OR2_X1 U360 ( .A1(n611), .A2(n610), .ZN(n612) );
  AND2_X1 U360bar ( .A1(n611bar), .A2(n610bar), .ZN(n612bar);
  OR2_X1 U361 ( .A1(in[213]), .A2(in[207]), .ZN(n610) );
  AND2_X1 U361bar ( .A1(inbar[213]), .A2(inbar[207]), .ZN(n610bar);
  OR2_X1 U362 ( .A1(in[215]), .A2(n609), .ZN(n611) );
  AND2_X1 U362bar ( .A1(inbar[215]), .A2(n609bar), .ZN(n611bar);
  OR2_X1 U363 ( .A1(in[230]), .A2(in[220]), .ZN(n609) );
  AND2_X1 U363bar ( .A1(inbar[230]), .A2(inbar[220]), .ZN(n609bar);
  OR2_X1 U364 ( .A1(n608), .A2(n607), .ZN(n613) );
  AND2_X1 U364bar ( .A1(n608bar), .A2(n607bar), .ZN(n613bar);
  OR2_X1 U365 ( .A1(in[251]), .A2(in[234]), .ZN(n607) );
  AND2_X1 U365bar ( .A1(inbar[251]), .A2(inbar[234]), .ZN(n607bar);
  OR2_X1 U366 ( .A1(in_17), .A2(n606), .ZN(n608) );
  AND2_X1 U366bar ( .A1(in_17bar), .A2(n606bar), .ZN(n608bar);
  OR2_X1 U367 ( .A1(in_65), .A2(in_56), .ZN(n606) );
  AND2_X1 U367bar ( .A1(in_65bar), .A2(in_56bar), .ZN(n606bar);
  OR2_X1 U368 ( .A1(n605), .A2(n604), .ZN(out[0]) );
  AND2_X1 U368bar ( .A1(n605bar), .A2(n604bar), .ZN(outbar[0]);
  OR2_X1 U369 ( .A1(n603), .A2(n602), .ZN(n604) );
  AND2_X1 U369bar ( .A1(n603bar), .A2(n602bar), .ZN(n604bar);
  OR2_X1 U370 ( .A1(n601), .A2(n600), .ZN(n602) );
  AND2_X1 U370bar ( .A1(n601bar), .A2(n600bar), .ZN(n602bar);
  OR2_X1 U371 ( .A1(n820), .A2(n785), .ZN(n600) );
  AND2_X1 U371bar ( .A1(n820bar), .A2(n785bar), .ZN(n600bar);
  OR2_X1 U372 ( .A1(n599), .A2(n598), .ZN(n785) );
  AND2_X1 U372bar ( .A1(n599bar), .A2(n598bar), .ZN(n785bar);
  OR2_X1 U373 ( .A1(n597), .A2(n596), .ZN(n598) );
  AND2_X1 U373bar ( .A1(n597bar), .A2(n596bar), .ZN(n598bar);
  OR2_X1 U374 ( .A1(n595), .A2(n594), .ZN(n596) );
  AND2_X1 U374bar ( .A1(n595bar), .A2(n594bar), .ZN(n596bar);
  OR2_X1 U375 ( .A1(in[135]), .A2(in[104]), .ZN(n594) );
  AND2_X1 U375bar ( .A1(inbar[135]), .A2(inbar[104]), .ZN(n594bar);
  OR2_X1 U376 ( .A1(in[188]), .A2(in[178]), .ZN(n595) );
  AND2_X1 U376bar ( .A1(inbar[188]), .A2(inbar[178]), .ZN(n595bar);
  OR2_X1 U377 ( .A1(n593), .A2(n592), .ZN(n597) );
  AND2_X1 U377bar ( .A1(n593bar), .A2(n592bar), .ZN(n597bar);
  OR2_X1 U378 ( .A1(in[217]), .A2(in[194]), .ZN(n592) );
  AND2_X1 U378bar ( .A1(inbar[217]), .A2(inbar[194]), .ZN(n592bar);
  OR2_X1 U379 ( .A1(in[237]), .A2(in[218]), .ZN(n593) );
  AND2_X1 U379bar ( .A1(inbar[237]), .A2(inbar[218]), .ZN(n593bar);
  OR2_X1 U380 ( .A1(n591), .A2(n590), .ZN(n599) );
  AND2_X1 U380bar ( .A1(n591bar), .A2(n590bar), .ZN(n599bar);
  OR2_X1 U381 ( .A1(n589), .A2(n588), .ZN(n590) );
  AND2_X1 U381bar ( .A1(n589bar), .A2(n588bar), .ZN(n590bar);
  OR2_X1 U382 ( .A1(in_2), .A2(in_10), .ZN(n588) );
  AND2_X1 U382bar ( .A1(in_2bar), .A2(in_10bar), .ZN(n588bar);
  OR2_X1 U383 ( .A1(in_47), .A2(in_22), .ZN(n589) );
  AND2_X1 U383bar ( .A1(in_47bar), .A2(in_22bar), .ZN(n589bar);
  OR2_X1 U384 ( .A1(n587), .A2(n586), .ZN(n591) );
  AND2_X1 U384bar ( .A1(n587bar), .A2(n586bar), .ZN(n591bar);
  OR2_X1 U385 ( .A1(in_56), .A2(in_54), .ZN(n586) );
  AND2_X1 U385bar ( .A1(in_56bar), .A2(in_54bar), .ZN(n586bar);
  OR2_X1 U386 ( .A1(in_63), .A2(in_61), .ZN(n587) );
  AND2_X1 U386bar ( .A1(in_63bar), .A2(in_61bar), .ZN(n587bar);
  OR2_X1 U387 ( .A1(n585), .A2(n584), .ZN(n820) );
  AND2_X1 U387bar ( .A1(n585bar), .A2(n584bar), .ZN(n820bar);
  OR2_X1 U388 ( .A1(n583), .A2(n582), .ZN(n584) );
  AND2_X1 U388bar ( .A1(n583bar), .A2(n582bar), .ZN(n584bar);
  OR2_X1 U389 ( .A1(n581), .A2(n580), .ZN(n582) );
  AND2_X1 U389bar ( .A1(n581bar), .A2(n580bar), .ZN(n582bar);
  OR2_X1 U390 ( .A1(in[158]), .A2(in[142]), .ZN(n580) );
  AND2_X1 U390bar ( .A1(inbar[158]), .A2(inbar[142]), .ZN(n580bar);
  OR2_X1 U391 ( .A1(in[175]), .A2(in[164]), .ZN(n581) );
  AND2_X1 U391bar ( .A1(inbar[175]), .A2(inbar[164]), .ZN(n581bar);
  OR2_X1 U392 ( .A1(n579), .A2(n578), .ZN(n583) );
  AND2_X1 U392bar ( .A1(n579bar), .A2(n578bar), .ZN(n583bar);
  OR2_X1 U393 ( .A1(in[228]), .A2(in[204]), .ZN(n578) );
  AND2_X1 U393bar ( .A1(inbar[228]), .A2(inbar[204]), .ZN(n578bar);
  OR2_X1 U394 ( .A1(in[91]), .A2(in[87]), .ZN(n579) );
  AND2_X1 U394bar ( .A1(inbar[91]), .A2(inbar[87]), .ZN(n579bar);
  OR2_X1 U395 ( .A1(n577), .A2(n576), .ZN(n585) );
  AND2_X1 U395bar ( .A1(n577bar), .A2(n576bar), .ZN(n585bar);
  OR2_X1 U396 ( .A1(n575), .A2(n574), .ZN(n576) );
  AND2_X1 U396bar ( .A1(n575bar), .A2(n574bar), .ZN(n576bar);
  OR2_X1 U397 ( .A1(in_21), .A2(in_11), .ZN(n574) );
  AND2_X1 U397bar ( .A1(in_21bar), .A2(in_11bar), .ZN(n574bar);
  OR2_X1 U398 ( .A1(in_5), .A2(in_3), .ZN(n575) );
  AND2_X1 U398bar ( .A1(in_5bar), .A2(in_3bar), .ZN(n575bar);
  OR2_X1 U399 ( .A1(n573), .A2(n572), .ZN(n577) );
  AND2_X1 U399bar ( .A1(n573bar), .A2(n572bar), .ZN(n577bar);
  OR2_X1 U400 ( .A1(in_68), .A2(in_64), .ZN(n572) );
  AND2_X1 U400bar ( .A1(in_68bar), .A2(in_64bar), .ZN(n572bar);
  OR2_X1 U401 ( .A1(in_76), .A2(in_73), .ZN(n573) );
  AND2_X1 U401bar ( .A1(in_76bar), .A2(in_73bar), .ZN(n573bar);
  OR2_X1 U402 ( .A1(n778), .A2(n571), .ZN(n601) );
  AND2_X1 U402bar ( .A1(n778bar), .A2(n571bar), .ZN(n601bar);
  OR2_X1 U403 ( .A1(in[100]), .A2(n965), .ZN(n571) );
  AND2_X1 U403bar ( .A1(inbar[100]), .A2(n965bar), .ZN(n571bar);
  OR2_X1 U404 ( .A1(n570), .A2(n569), .ZN(n965) );
  AND2_X1 U404bar ( .A1(n570bar), .A2(n569bar), .ZN(n965bar);
  OR2_X1 U405 ( .A1(n568), .A2(n567), .ZN(n569) );
  AND2_X1 U405bar ( .A1(n568bar), .A2(n567bar), .ZN(n569bar);
  OR2_X1 U406 ( .A1(n566), .A2(n565), .ZN(n567) );
  AND2_X1 U406bar ( .A1(n566bar), .A2(n565bar), .ZN(n567bar);
  OR2_X1 U407 ( .A1(n817), .A2(n750), .ZN(n565) );
  AND2_X1 U407bar ( .A1(n817bar), .A2(n750bar), .ZN(n565bar);
  OR2_X1 U408 ( .A1(n564), .A2(n563), .ZN(n750) );
  AND2_X1 U408bar ( .A1(n564bar), .A2(n563bar), .ZN(n750bar);
  OR2_X1 U409 ( .A1(n562), .A2(n561), .ZN(n563) );
  AND2_X1 U409bar ( .A1(n562bar), .A2(n561bar), .ZN(n563bar);
  OR2_X1 U410 ( .A1(n560), .A2(n559), .ZN(n561) );
  AND2_X1 U410bar ( .A1(n560bar), .A2(n559bar), .ZN(n561bar);
  OR2_X1 U411 ( .A1(in[119]), .A2(in[103]), .ZN(n559) );
  AND2_X1 U411bar ( .A1(inbar[119]), .A2(inbar[103]), .ZN(n559bar);
  OR2_X1 U412 ( .A1(in[137]), .A2(in[133]), .ZN(n560) );
  AND2_X1 U412bar ( .A1(inbar[137]), .A2(inbar[133]), .ZN(n560bar);
  OR2_X1 U413 ( .A1(n558), .A2(n557), .ZN(n562) );
  AND2_X1 U413bar ( .A1(n558bar), .A2(n557bar), .ZN(n562bar);
  OR2_X1 U414 ( .A1(in[176]), .A2(in[173]), .ZN(n557) );
  AND2_X1 U414bar ( .A1(inbar[176]), .A2(inbar[173]), .ZN(n557bar);
  OR2_X1 U415 ( .A1(in[210]), .A2(in[181]), .ZN(n558) );
  AND2_X1 U415bar ( .A1(inbar[210]), .A2(inbar[181]), .ZN(n558bar);
  OR2_X1 U416 ( .A1(n556), .A2(n555), .ZN(n564) );
  AND2_X1 U416bar ( .A1(n556bar), .A2(n555bar), .ZN(n564bar);
  OR2_X1 U417 ( .A1(n554), .A2(n553), .ZN(n555) );
  AND2_X1 U417bar ( .A1(n554bar), .A2(n553bar), .ZN(n555bar);
  OR2_X1 U418 ( .A1(in_13), .A2(in[234]), .ZN(n553) );
  AND2_X1 U418bar ( .A1(in_13bar), .A2(inbar[234]), .ZN(n553bar);
  OR2_X1 U419 ( .A1(in_38), .A2(in_32), .ZN(n554) );
  AND2_X1 U419bar ( .A1(in_38bar), .A2(in_32bar), .ZN(n554bar);
  OR2_X1 U420 ( .A1(n552), .A2(n551), .ZN(n556) );
  AND2_X1 U420bar ( .A1(n552bar), .A2(n551bar), .ZN(n556bar);
  OR2_X1 U421 ( .A1(in_42), .A2(in_41), .ZN(n551) );
  AND2_X1 U421bar ( .A1(in_42bar), .A2(in_41bar), .ZN(n551bar);
  OR2_X1 U422 ( .A1(in_7), .A2(in_49), .ZN(n552) );
  AND2_X1 U422bar ( .A1(in_7bar), .A2(in_49bar), .ZN(n552bar);
  OR2_X1 U423 ( .A1(n550), .A2(n549), .ZN(n817) );
  AND2_X1 U423bar ( .A1(n550bar), .A2(n549bar), .ZN(n817bar);
  OR2_X1 U424 ( .A1(n548), .A2(n547), .ZN(n549) );
  AND2_X1 U424bar ( .A1(n548bar), .A2(n547bar), .ZN(n549bar);
  OR2_X1 U425 ( .A1(n546), .A2(n545), .ZN(n547) );
  AND2_X1 U425bar ( .A1(n546bar), .A2(n545bar), .ZN(n547bar);
  OR2_X1 U426 ( .A1(in[159]), .A2(in[105]), .ZN(n545) );
  AND2_X1 U426bar ( .A1(inbar[159]), .A2(inbar[105]), .ZN(n545bar);
  OR2_X1 U427 ( .A1(in[206]), .A2(in[183]), .ZN(n546) );
  AND2_X1 U427bar ( .A1(inbar[206]), .A2(inbar[183]), .ZN(n546bar);
  OR2_X1 U428 ( .A1(n544), .A2(n543), .ZN(n548) );
  AND2_X1 U428bar ( .A1(n544bar), .A2(n543bar), .ZN(n548bar);
  OR2_X1 U429 ( .A1(in[229]), .A2(in[219]), .ZN(n543) );
  AND2_X1 U429bar ( .A1(inbar[229]), .A2(inbar[219]), .ZN(n543bar);
  OR2_X1 U430 ( .A1(in[235]), .A2(in[232]), .ZN(n544) );
  AND2_X1 U430bar ( .A1(inbar[235]), .A2(inbar[232]), .ZN(n544bar);
  OR2_X1 U431 ( .A1(n542), .A2(n541), .ZN(n550) );
  AND2_X1 U431bar ( .A1(n542bar), .A2(n541bar), .ZN(n550bar);
  OR2_X1 U432 ( .A1(n540), .A2(n539), .ZN(n541) );
  AND2_X1 U432bar ( .A1(n540bar), .A2(n539bar), .ZN(n541bar);
  OR2_X1 U433 ( .A1(in[249]), .A2(in[242]), .ZN(n539) );
  AND2_X1 U433bar ( .A1(inbar[249]), .A2(inbar[242]), .ZN(n539bar);
  OR2_X1 U434 ( .A1(in[89]), .A2(in[254]), .ZN(n540) );
  AND2_X1 U434bar ( .A1(inbar[89]), .A2(inbar[254]), .ZN(n540bar);
  OR2_X1 U435 ( .A1(n538), .A2(n537), .ZN(n542) );
  AND2_X1 U435bar ( .A1(n538bar), .A2(n537bar), .ZN(n542bar);
  OR2_X1 U436 ( .A1(in_14), .A2(in[99]), .ZN(n537) );
  AND2_X1 U436bar ( .A1(in_14bar), .A2(inbar[99]), .ZN(n537bar);
  OR2_X1 U437 ( .A1(in_60), .A2(in_18), .ZN(n538) );
  AND2_X1 U437bar ( .A1(in_60bar), .A2(in_18bar), .ZN(n538bar);
  OR2_X1 U438 ( .A1(in[113]), .A2(n763), .ZN(n566) );
  AND2_X1 U438bar ( .A1(inbar[113]), .A2(n763bar), .ZN(n566bar);
  OR2_X1 U439 ( .A1(n536), .A2(n535), .ZN(n763) );
  AND2_X1 U439bar ( .A1(n536bar), .A2(n535bar), .ZN(n763bar);
  OR2_X1 U440 ( .A1(n534), .A2(n533), .ZN(n535) );
  AND2_X1 U440bar ( .A1(n534bar), .A2(n533bar), .ZN(n535bar);
  OR2_X1 U441 ( .A1(n532), .A2(n531), .ZN(n533) );
  AND2_X1 U441bar ( .A1(n532bar), .A2(n531bar), .ZN(n533bar);
  OR2_X1 U442 ( .A1(in[115]), .A2(in[110]), .ZN(n531) );
  AND2_X1 U442bar ( .A1(inbar[115]), .A2(inbar[110]), .ZN(n531bar);
  OR2_X1 U443 ( .A1(in[125]), .A2(in[117]), .ZN(n532) );
  AND2_X1 U443bar ( .A1(inbar[125]), .A2(inbar[117]), .ZN(n532bar);
  OR2_X1 U444 ( .A1(n530), .A2(n529), .ZN(n534) );
  AND2_X1 U444bar ( .A1(n530bar), .A2(n529bar), .ZN(n534bar);
  OR2_X1 U445 ( .A1(in[180]), .A2(in[128]), .ZN(n529) );
  AND2_X1 U445bar ( .A1(inbar[180]), .A2(inbar[128]), .ZN(n529bar);
  OR2_X1 U446 ( .A1(in[205]), .A2(in[201]), .ZN(n530) );
  AND2_X1 U446bar ( .A1(inbar[205]), .A2(inbar[201]), .ZN(n530bar);
  OR2_X1 U447 ( .A1(n528), .A2(n527), .ZN(n536) );
  AND2_X1 U447bar ( .A1(n528bar), .A2(n527bar), .ZN(n536bar);
  OR2_X1 U448 ( .A1(n526), .A2(n525), .ZN(n527) );
  AND2_X1 U448bar ( .A1(n526bar), .A2(n525bar), .ZN(n527bar);
  OR2_X1 U449 ( .A1(in[244]), .A2(in[239]), .ZN(n525) );
  AND2_X1 U449bar ( .A1(inbar[244]), .A2(inbar[239]), .ZN(n525bar);
  OR2_X1 U450 ( .A1(in[95]), .A2(in[83]), .ZN(n526) );
  AND2_X1 U450bar ( .A1(inbar[95]), .A2(inbar[83]), .ZN(n526bar);
  OR2_X1 U451 ( .A1(n524), .A2(n523), .ZN(n528) );
  AND2_X1 U451bar ( .A1(n524bar), .A2(n523bar), .ZN(n528bar);
  OR2_X1 U452 ( .A1(in_24), .A2(in[97]), .ZN(n523) );
  AND2_X1 U452bar ( .A1(in_24bar), .A2(inbar[97]), .ZN(n523bar);
  OR2_X1 U453 ( .A1(in_33), .A2(in_27), .ZN(n524) );
  AND2_X1 U453bar ( .A1(in_33bar), .A2(in_27bar), .ZN(n524bar);
  OR2_X1 U454 ( .A1(n522), .A2(n521), .ZN(n568) );
  AND2_X1 U454bar ( .A1(n522bar), .A2(n521bar), .ZN(n568bar);
  OR2_X1 U455 ( .A1(in[145]), .A2(in[126]), .ZN(n521) );
  AND2_X1 U455bar ( .A1(inbar[145]), .A2(inbar[126]), .ZN(n521bar);
  OR2_X1 U456 ( .A1(in[169]), .A2(n520), .ZN(n522) );
  AND2_X1 U456bar ( .A1(inbar[169]), .A2(n520bar), .ZN(n522bar);
  OR2_X1 U457 ( .A1(in[221]), .A2(in[172]), .ZN(n520) );
  AND2_X1 U457bar ( .A1(inbar[221]), .A2(inbar[172]), .ZN(n520bar);
  OR2_X1 U458 ( .A1(n519), .A2(n518), .ZN(n570) );
  AND2_X1 U458bar ( .A1(n519bar), .A2(n518bar), .ZN(n570bar);
  OR2_X1 U459 ( .A1(n517), .A2(n516), .ZN(n518) );
  AND2_X1 U459bar ( .A1(n517bar), .A2(n516bar), .ZN(n518bar);
  OR2_X1 U460 ( .A1(in[241]), .A2(in[224]), .ZN(n516) );
  AND2_X1 U460bar ( .A1(inbar[241]), .A2(inbar[224]), .ZN(n516bar);
  OR2_X1 U461 ( .A1(in[86]), .A2(n515), .ZN(n517) );
  AND2_X1 U461bar ( .A1(inbar[86]), .A2(n515bar), .ZN(n517bar);
  OR2_X1 U462 ( .A1(in_43), .A2(in_34), .ZN(n515) );
  AND2_X1 U462bar ( .A1(in_43bar), .A2(in_34bar), .ZN(n515bar);
  OR2_X1 U463 ( .A1(n514), .A2(n513), .ZN(n519) );
  AND2_X1 U463bar ( .A1(n514bar), .A2(n513bar), .ZN(n519bar);
  OR2_X1 U464 ( .A1(in_65), .A2(in_51), .ZN(n513) );
  AND2_X1 U464bar ( .A1(in_65bar), .A2(in_51bar), .ZN(n513bar);
  OR2_X1 U465 ( .A1(in_75), .A2(n512), .ZN(n514) );
  AND2_X1 U465bar ( .A1(in_75bar), .A2(n512bar), .ZN(n514bar);
  OR2_X1 U466 ( .A1(in_81), .A2(in_77), .ZN(n512) );
  AND2_X1 U466bar ( .A1(in_81bar), .A2(in_77bar), .ZN(n512bar);
  OR2_X1 U467 ( .A1(n511), .A2(n510), .ZN(n778) );
  AND2_X1 U467bar ( .A1(n511bar), .A2(n510bar), .ZN(n778bar);
  OR2_X1 U468 ( .A1(n509), .A2(n508), .ZN(n510) );
  AND2_X1 U468bar ( .A1(n509bar), .A2(n508bar), .ZN(n510bar);
  OR2_X1 U469 ( .A1(n507), .A2(n506), .ZN(n508) );
  AND2_X1 U469bar ( .A1(n507bar), .A2(n506bar), .ZN(n508bar);
  OR2_X1 U470 ( .A1(in[107]), .A2(in[101]), .ZN(n506) );
  AND2_X1 U470bar ( .A1(inbar[107]), .A2(inbar[101]), .ZN(n506bar);
  OR2_X1 U471 ( .A1(in[139]), .A2(in[132]), .ZN(n507) );
  AND2_X1 U471bar ( .A1(inbar[139]), .A2(inbar[132]), .ZN(n507bar);
  OR2_X1 U472 ( .A1(n505), .A2(n504), .ZN(n509) );
  AND2_X1 U472bar ( .A1(n505bar), .A2(n504bar), .ZN(n509bar);
  OR2_X1 U473 ( .A1(in[146]), .A2(in[141]), .ZN(n504) );
  AND2_X1 U473bar ( .A1(inbar[146]), .A2(inbar[141]), .ZN(n504bar);
  OR2_X1 U474 ( .A1(in[203]), .A2(in[179]), .ZN(n505) );
  AND2_X1 U474bar ( .A1(inbar[203]), .A2(inbar[179]), .ZN(n505bar);
  OR2_X1 U475 ( .A1(n503), .A2(n502), .ZN(n511) );
  AND2_X1 U475bar ( .A1(n503bar), .A2(n502bar), .ZN(n511bar);
  OR2_X1 U476 ( .A1(n501), .A2(n500), .ZN(n502) );
  AND2_X1 U476bar ( .A1(n501bar), .A2(n500bar), .ZN(n502bar);
  OR2_X1 U477 ( .A1(in[243]), .A2(in[222]), .ZN(n500) );
  AND2_X1 U477bar ( .A1(inbar[243]), .A2(inbar[222]), .ZN(n500bar);
  OR2_X1 U478 ( .A1(in[251]), .A2(in[250]), .ZN(n501) );
  AND2_X1 U478bar ( .A1(inbar[251]), .A2(inbar[250]), .ZN(n501bar);
  OR2_X1 U479 ( .A1(n499), .A2(n498), .ZN(n503) );
  AND2_X1 U479bar ( .A1(n499bar), .A2(n498bar), .ZN(n503bar);
  OR2_X1 U480 ( .A1(in_37), .A2(in_19), .ZN(n498) );
  AND2_X1 U480bar ( .A1(in_37bar), .A2(in_19bar), .ZN(n498bar);
  OR2_X1 U481 ( .A1(in_78), .A2(in_6), .ZN(n499) );
  AND2_X1 U481bar ( .A1(in_78bar), .A2(in_6bar), .ZN(n499bar);
  OR2_X1 U482 ( .A1(n497), .A2(n496), .ZN(n603) );
  AND2_X1 U482bar ( .A1(n497bar), .A2(n496bar), .ZN(n603bar);
  OR2_X1 U483 ( .A1(in[112]), .A2(in[102]), .ZN(n496) );
  AND2_X1 U483bar ( .A1(inbar[112]), .A2(inbar[102]), .ZN(n496bar);
  OR2_X1 U484 ( .A1(in[123]), .A2(n495), .ZN(n497) );
  AND2_X1 U484bar ( .A1(inbar[123]), .A2(n495bar), .ZN(n497bar);
  OR2_X1 U485 ( .A1(in[143]), .A2(in[130]), .ZN(n495) );
  AND2_X1 U485bar ( .A1(inbar[143]), .A2(inbar[130]), .ZN(n495bar);
  OR2_X1 U486 ( .A1(n494), .A2(n493), .ZN(n605) );
  AND2_X1 U486bar ( .A1(n494bar), .A2(n493bar), .ZN(n605bar);
  OR2_X1 U487 ( .A1(n492), .A2(n491), .ZN(n493) );
  AND2_X1 U487bar ( .A1(n492bar), .A2(n491bar), .ZN(n493bar);
  OR2_X1 U488 ( .A1(in[216]), .A2(in[213]), .ZN(n491) );
  AND2_X1 U488bar ( .A1(inbar[216]), .A2(inbar[213]), .ZN(n491bar);
  OR2_X1 U489 ( .A1(in[227]), .A2(n490), .ZN(n492) );
  AND2_X1 U489bar ( .A1(inbar[227]), .A2(n490bar), .ZN(n492bar);
  OR2_X1 U490 ( .A1(in_0), .A2(in[248]), .ZN(n490) );
  AND2_X1 U490bar ( .A1(in_0bar), .A2(inbar[248]), .ZN(n490bar);
  OR2_X1 U491 ( .A1(n489), .A2(n488), .ZN(n494) );
  AND2_X1 U491bar ( .A1(n489bar), .A2(n488bar), .ZN(n494bar);
  OR2_X1 U492 ( .A1(in_46), .A2(in_44), .ZN(n488) );
  AND2_X1 U492bar ( .A1(in_46bar), .A2(in_44bar), .ZN(n488bar);
  OR2_X1 U493 ( .A1(in_50), .A2(n487), .ZN(n489) );
  AND2_X1 U493bar ( .A1(in_50bar), .A2(n487bar), .ZN(n489bar);
  OR2_X1 U494 ( .A1(in_9), .A2(in_80), .ZN(n487) );
  AND2_X1 U494bar ( .A1(in_9bar), .A2(in_80bar), .ZN(n487bar);
endmodule




module sBox_8 ( in, out );
  input [7:0] in;
  //input_done

  output [7:0] out;
  //output_done

  wire   [255:0] decodeOut;
  //wire_done

  decode_8 dec ( .in(in), .out(decodeOut) );
  encode_8 enc ( .in(decodeOut), .out(out) );
endmodule


module CD2_33 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_34 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_35 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
 
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_36 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD4_17 ( a, b, y );
  input [3:0] a;
  input [3:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  //input_done

  output [15:0] y;
  reg [15:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]);
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]);
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]);
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]);
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]);
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]);
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]);
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]);
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]);
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]);
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]);
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]);
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]);
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]);
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]);
endmodule




module CD4_18 ( a, b, y );
  input [3:0] a;
  input [3:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  //input_done

  output [15:0] y;
  reg [15:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]);
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]);
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]);
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]);
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]);
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]);
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]);
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]);
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]);
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]);
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]);
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]);
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]);
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]);
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]);
endmodule




module CD16_9 ( a, b, y );
  input [15:0] a;
  input [15:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign abar[8] = ~a[8];
  assign abar[9] = ~a[9];
  assign abar[10] = ~a[10];
  assign abar[11] = ~a[11];
  assign abar[12] = ~a[12];
  assign abar[13] = ~a[13];
  assign abar[14] = ~a[14];
  assign abar[15] = ~a[15];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign bbar[8] = ~b[8];
  assign bbar[9] = ~b[9];
  assign bbar[10] = ~b[10];
  assign bbar[11] = ~b[11];
  assign bbar[12] = ~b[12];
  assign bbar[13] = ~b[13];
  assign bbar[14] = ~b[14];
  assign bbar[15] = ~b[15];
  //input_done

  output [255:0] y;
  reg [255:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[9]), .A2(a[0]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[9]), .A2(abar[0]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[3]), .A2(a[6]), .ZN(y[99]) );
  OR2_X1 U2bar ( .A1(bbar[3]), .A2(abar[6]), .ZN(ybar[99]);
  AND2_X1 U3 ( .A1(b[2]), .A2(a[6]), .ZN(y[98]) );
  OR2_X1 U3bar ( .A1(bbar[2]), .A2(abar[6]), .ZN(ybar[98]);
  AND2_X1 U4 ( .A1(b[1]), .A2(a[6]), .ZN(y[97]) );
  OR2_X1 U4bar ( .A1(bbar[1]), .A2(abar[6]), .ZN(ybar[97]);
  AND2_X1 U5 ( .A1(b[0]), .A2(a[6]), .ZN(y[96]) );
  OR2_X1 U5bar ( .A1(bbar[0]), .A2(abar[6]), .ZN(ybar[96]);
  AND2_X1 U6 ( .A1(b[15]), .A2(a[5]), .ZN(y[95]) );
  OR2_X1 U6bar ( .A1(bbar[15]), .A2(abar[5]), .ZN(ybar[95]);
  AND2_X1 U7 ( .A1(b[14]), .A2(a[5]), .ZN(y[94]) );
  OR2_X1 U7bar ( .A1(bbar[14]), .A2(abar[5]), .ZN(ybar[94]);
  AND2_X1 U8 ( .A1(b[13]), .A2(a[5]), .ZN(y[93]) );
  OR2_X1 U8bar ( .A1(bbar[13]), .A2(abar[5]), .ZN(ybar[93]);
  AND2_X1 U9 ( .A1(b[12]), .A2(a[5]), .ZN(y[92]) );
  OR2_X1 U9bar ( .A1(bbar[12]), .A2(abar[5]), .ZN(ybar[92]);
  AND2_X1 U10 ( .A1(b[11]), .A2(a[5]), .ZN(y[91]) );
  OR2_X1 U10bar ( .A1(bbar[11]), .A2(abar[5]), .ZN(ybar[91]);
  AND2_X1 U11 ( .A1(b[10]), .A2(a[5]), .ZN(y[90]) );
  OR2_X1 U11bar ( .A1(bbar[10]), .A2(abar[5]), .ZN(ybar[90]);
  AND2_X1 U12 ( .A1(b[8]), .A2(a[0]), .ZN(y[8]) );
  OR2_X1 U12bar ( .A1(bbar[8]), .A2(abar[0]), .ZN(ybar[8]);
  AND2_X1 U13 ( .A1(a[5]), .A2(b[9]), .ZN(y[89]) );
  OR2_X1 U13bar ( .A1(abar[5]), .A2(bbar[9]), .ZN(ybar[89]);
  AND2_X1 U14 ( .A1(b[8]), .A2(a[5]), .ZN(y[88]) );
  OR2_X1 U14bar ( .A1(bbar[8]), .A2(abar[5]), .ZN(ybar[88]);
  AND2_X1 U15 ( .A1(b[7]), .A2(a[5]), .ZN(y[87]) );
  OR2_X1 U15bar ( .A1(bbar[7]), .A2(abar[5]), .ZN(ybar[87]);
  AND2_X1 U16 ( .A1(b[6]), .A2(a[5]), .ZN(y[86]) );
  OR2_X1 U16bar ( .A1(bbar[6]), .A2(abar[5]), .ZN(ybar[86]);
  AND2_X1 U17 ( .A1(b[5]), .A2(a[5]), .ZN(y[85]) );
  OR2_X1 U17bar ( .A1(bbar[5]), .A2(abar[5]), .ZN(ybar[85]);
  AND2_X1 U18 ( .A1(b[4]), .A2(a[5]), .ZN(y[84]) );
  OR2_X1 U18bar ( .A1(bbar[4]), .A2(abar[5]), .ZN(ybar[84]);
  AND2_X1 U19 ( .A1(a[5]), .A2(b[3]), .ZN(y[83]) );
  OR2_X1 U19bar ( .A1(abar[5]), .A2(bbar[3]), .ZN(ybar[83]);
  AND2_X1 U20 ( .A1(a[5]), .A2(b[2]), .ZN(y[82]) );
  OR2_X1 U20bar ( .A1(abar[5]), .A2(bbar[2]), .ZN(ybar[82]);
  AND2_X1 U21 ( .A1(a[5]), .A2(b[1]), .ZN(y[81]) );
  OR2_X1 U21bar ( .A1(abar[5]), .A2(bbar[1]), .ZN(ybar[81]);
  AND2_X1 U22 ( .A1(a[5]), .A2(b[0]), .ZN(y[80]) );
  OR2_X1 U22bar ( .A1(abar[5]), .A2(bbar[0]), .ZN(ybar[80]);
  AND2_X1 U23 ( .A1(b[7]), .A2(a[0]), .ZN(y[7]) );
  OR2_X1 U23bar ( .A1(bbar[7]), .A2(abar[0]), .ZN(ybar[7]);
  AND2_X1 U24 ( .A1(a[4]), .A2(b[15]), .ZN(y[79]) );
  OR2_X1 U24bar ( .A1(abar[4]), .A2(bbar[15]), .ZN(ybar[79]);
  AND2_X1 U25 ( .A1(a[4]), .A2(b[14]), .ZN(y[78]) );
  OR2_X1 U25bar ( .A1(abar[4]), .A2(bbar[14]), .ZN(ybar[78]);
  AND2_X1 U26 ( .A1(a[4]), .A2(b[13]), .ZN(y[77]) );
  OR2_X1 U26bar ( .A1(abar[4]), .A2(bbar[13]), .ZN(ybar[77]);
  AND2_X1 U27 ( .A1(a[4]), .A2(b[12]), .ZN(y[76]) );
  OR2_X1 U27bar ( .A1(abar[4]), .A2(bbar[12]), .ZN(ybar[76]);
  AND2_X1 U28 ( .A1(a[4]), .A2(b[11]), .ZN(y[75]) );
  OR2_X1 U28bar ( .A1(abar[4]), .A2(bbar[11]), .ZN(ybar[75]);
  AND2_X1 U29 ( .A1(a[4]), .A2(b[10]), .ZN(y[74]) );
  OR2_X1 U29bar ( .A1(abar[4]), .A2(bbar[10]), .ZN(ybar[74]);
  AND2_X1 U30 ( .A1(a[4]), .A2(b[9]), .ZN(y[73]) );
  OR2_X1 U30bar ( .A1(abar[4]), .A2(bbar[9]), .ZN(ybar[73]);
  AND2_X1 U31 ( .A1(a[4]), .A2(b[8]), .ZN(y[72]) );
  OR2_X1 U31bar ( .A1(abar[4]), .A2(bbar[8]), .ZN(ybar[72]);
  AND2_X1 U32 ( .A1(a[4]), .A2(b[7]), .ZN(y[71]) );
  OR2_X1 U32bar ( .A1(abar[4]), .A2(bbar[7]), .ZN(ybar[71]);
  AND2_X1 U33 ( .A1(a[4]), .A2(b[6]), .ZN(y[70]) );
  OR2_X1 U33bar ( .A1(abar[4]), .A2(bbar[6]), .ZN(ybar[70]);
  AND2_X1 U34 ( .A1(b[6]), .A2(a[0]), .ZN(y[6]) );
  OR2_X1 U34bar ( .A1(bbar[6]), .A2(abar[0]), .ZN(ybar[6]);
  AND2_X1 U35 ( .A1(a[4]), .A2(b[5]), .ZN(y[69]) );
  OR2_X1 U35bar ( .A1(abar[4]), .A2(bbar[5]), .ZN(ybar[69]);
  AND2_X1 U36 ( .A1(a[4]), .A2(b[4]), .ZN(y[68]) );
  OR2_X1 U36bar ( .A1(abar[4]), .A2(bbar[4]), .ZN(ybar[68]);
  AND2_X1 U37 ( .A1(a[4]), .A2(b[3]), .ZN(y[67]) );
  OR2_X1 U37bar ( .A1(abar[4]), .A2(bbar[3]), .ZN(ybar[67]);
  AND2_X1 U38 ( .A1(a[4]), .A2(b[2]), .ZN(y[66]) );
  OR2_X1 U38bar ( .A1(abar[4]), .A2(bbar[2]), .ZN(ybar[66]);
  AND2_X1 U39 ( .A1(a[4]), .A2(b[1]), .ZN(y[65]) );
  OR2_X1 U39bar ( .A1(abar[4]), .A2(bbar[1]), .ZN(ybar[65]);
  AND2_X1 U40 ( .A1(a[4]), .A2(b[0]), .ZN(y[64]) );
  OR2_X1 U40bar ( .A1(abar[4]), .A2(bbar[0]), .ZN(ybar[64]);
  AND2_X1 U41 ( .A1(a[3]), .A2(b[15]), .ZN(y[63]) );
  OR2_X1 U41bar ( .A1(abar[3]), .A2(bbar[15]), .ZN(ybar[63]);
  AND2_X1 U42 ( .A1(a[3]), .A2(b[14]), .ZN(y[62]) );
  OR2_X1 U42bar ( .A1(abar[3]), .A2(bbar[14]), .ZN(ybar[62]);
  AND2_X1 U43 ( .A1(a[3]), .A2(b[13]), .ZN(y[61]) );
  OR2_X1 U43bar ( .A1(abar[3]), .A2(bbar[13]), .ZN(ybar[61]);
  AND2_X1 U44 ( .A1(a[3]), .A2(b[12]), .ZN(y[60]) );
  OR2_X1 U44bar ( .A1(abar[3]), .A2(bbar[12]), .ZN(ybar[60]);
  AND2_X1 U45 ( .A1(b[5]), .A2(a[0]), .ZN(y[5]) );
  OR2_X1 U45bar ( .A1(bbar[5]), .A2(abar[0]), .ZN(ybar[5]);
  AND2_X1 U46 ( .A1(a[3]), .A2(b[11]), .ZN(y[59]) );
  OR2_X1 U46bar ( .A1(abar[3]), .A2(bbar[11]), .ZN(ybar[59]);
  AND2_X1 U47 ( .A1(a[3]), .A2(b[10]), .ZN(y[58]) );
  OR2_X1 U47bar ( .A1(abar[3]), .A2(bbar[10]), .ZN(ybar[58]);
  AND2_X1 U48 ( .A1(a[3]), .A2(b[9]), .ZN(y[57]) );
  OR2_X1 U48bar ( .A1(abar[3]), .A2(bbar[9]), .ZN(ybar[57]);
  AND2_X1 U49 ( .A1(a[3]), .A2(b[8]), .ZN(y[56]) );
  OR2_X1 U49bar ( .A1(abar[3]), .A2(bbar[8]), .ZN(ybar[56]);
  AND2_X1 U50 ( .A1(a[3]), .A2(b[7]), .ZN(y[55]) );
  OR2_X1 U50bar ( .A1(abar[3]), .A2(bbar[7]), .ZN(ybar[55]);
  AND2_X1 U51 ( .A1(a[3]), .A2(b[6]), .ZN(y[54]) );
  OR2_X1 U51bar ( .A1(abar[3]), .A2(bbar[6]), .ZN(ybar[54]);
  AND2_X1 U52 ( .A1(a[3]), .A2(b[5]), .ZN(y[53]) );
  OR2_X1 U52bar ( .A1(abar[3]), .A2(bbar[5]), .ZN(ybar[53]);
  AND2_X1 U53 ( .A1(a[3]), .A2(b[4]), .ZN(y[52]) );
  OR2_X1 U53bar ( .A1(abar[3]), .A2(bbar[4]), .ZN(ybar[52]);
  AND2_X1 U54 ( .A1(a[3]), .A2(b[3]), .ZN(y[51]) );
  OR2_X1 U54bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[51]);
  AND2_X1 U55 ( .A1(a[3]), .A2(b[2]), .ZN(y[50]) );
  OR2_X1 U55bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[50]);
  AND2_X1 U56 ( .A1(b[4]), .A2(a[0]), .ZN(y[4]) );
  OR2_X1 U56bar ( .A1(bbar[4]), .A2(abar[0]), .ZN(ybar[4]);
  AND2_X1 U57 ( .A1(a[3]), .A2(b[1]), .ZN(y[49]) );
  OR2_X1 U57bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[49]);
  AND2_X1 U58 ( .A1(a[3]), .A2(b[0]), .ZN(y[48]) );
  OR2_X1 U58bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[48]);
  AND2_X1 U59 ( .A1(a[2]), .A2(b[15]), .ZN(y[47]) );
  OR2_X1 U59bar ( .A1(abar[2]), .A2(bbar[15]), .ZN(ybar[47]);
  AND2_X1 U60 ( .A1(a[2]), .A2(b[14]), .ZN(y[46]) );
  OR2_X1 U60bar ( .A1(abar[2]), .A2(bbar[14]), .ZN(ybar[46]);
  AND2_X1 U61 ( .A1(a[2]), .A2(b[13]), .ZN(y[45]) );
  OR2_X1 U61bar ( .A1(abar[2]), .A2(bbar[13]), .ZN(ybar[45]);
  AND2_X1 U62 ( .A1(a[2]), .A2(b[12]), .ZN(y[44]) );
  OR2_X1 U62bar ( .A1(abar[2]), .A2(bbar[12]), .ZN(ybar[44]);
  AND2_X1 U63 ( .A1(a[2]), .A2(b[11]), .ZN(y[43]) );
  OR2_X1 U63bar ( .A1(abar[2]), .A2(bbar[11]), .ZN(ybar[43]);
  AND2_X1 U64 ( .A1(a[2]), .A2(b[10]), .ZN(y[42]) );
  OR2_X1 U64bar ( .A1(abar[2]), .A2(bbar[10]), .ZN(ybar[42]);
  AND2_X1 U65 ( .A1(a[2]), .A2(b[9]), .ZN(y[41]) );
  OR2_X1 U65bar ( .A1(abar[2]), .A2(bbar[9]), .ZN(ybar[41]);
  AND2_X1 U66 ( .A1(a[2]), .A2(b[8]), .ZN(y[40]) );
  OR2_X1 U66bar ( .A1(abar[2]), .A2(bbar[8]), .ZN(ybar[40]);
  AND2_X1 U67 ( .A1(b[3]), .A2(a[0]), .ZN(y[3]) );
  OR2_X1 U67bar ( .A1(bbar[3]), .A2(abar[0]), .ZN(ybar[3]);
  AND2_X1 U68 ( .A1(a[2]), .A2(b[7]), .ZN(y[39]) );
  OR2_X1 U68bar ( .A1(abar[2]), .A2(bbar[7]), .ZN(ybar[39]);
  AND2_X1 U69 ( .A1(a[2]), .A2(b[6]), .ZN(y[38]) );
  OR2_X1 U69bar ( .A1(abar[2]), .A2(bbar[6]), .ZN(ybar[38]);
  AND2_X1 U70 ( .A1(a[2]), .A2(b[5]), .ZN(y[37]) );
  OR2_X1 U70bar ( .A1(abar[2]), .A2(bbar[5]), .ZN(ybar[37]);
  AND2_X1 U71 ( .A1(a[2]), .A2(b[4]), .ZN(y[36]) );
  OR2_X1 U71bar ( .A1(abar[2]), .A2(bbar[4]), .ZN(ybar[36]);
  AND2_X1 U72 ( .A1(a[2]), .A2(b[3]), .ZN(y[35]) );
  OR2_X1 U72bar ( .A1(abar[2]), .A2(bbar[3]), .ZN(ybar[35]);
  AND2_X1 U73 ( .A1(a[2]), .A2(b[2]), .ZN(y[34]) );
  OR2_X1 U73bar ( .A1(abar[2]), .A2(bbar[2]), .ZN(ybar[34]);
  AND2_X1 U74 ( .A1(a[2]), .A2(b[1]), .ZN(y[33]) );
  OR2_X1 U74bar ( .A1(abar[2]), .A2(bbar[1]), .ZN(ybar[33]);
  AND2_X1 U75 ( .A1(a[2]), .A2(b[0]), .ZN(y[32]) );
  OR2_X1 U75bar ( .A1(abar[2]), .A2(bbar[0]), .ZN(ybar[32]);
  AND2_X1 U76 ( .A1(a[1]), .A2(b[15]), .ZN(y[31]) );
  OR2_X1 U76bar ( .A1(abar[1]), .A2(bbar[15]), .ZN(ybar[31]);
  AND2_X1 U77 ( .A1(a[1]), .A2(b[14]), .ZN(y[30]) );
  OR2_X1 U77bar ( .A1(abar[1]), .A2(bbar[14]), .ZN(ybar[30]);
  AND2_X1 U78 ( .A1(b[2]), .A2(a[0]), .ZN(y[2]) );
  OR2_X1 U78bar ( .A1(bbar[2]), .A2(abar[0]), .ZN(ybar[2]);
  AND2_X1 U79 ( .A1(a[1]), .A2(b[13]), .ZN(y[29]) );
  OR2_X1 U79bar ( .A1(abar[1]), .A2(bbar[13]), .ZN(ybar[29]);
  AND2_X1 U80 ( .A1(a[1]), .A2(b[12]), .ZN(y[28]) );
  OR2_X1 U80bar ( .A1(abar[1]), .A2(bbar[12]), .ZN(ybar[28]);
  AND2_X1 U81 ( .A1(a[1]), .A2(b[11]), .ZN(y[27]) );
  OR2_X1 U81bar ( .A1(abar[1]), .A2(bbar[11]), .ZN(ybar[27]);
  AND2_X1 U82 ( .A1(a[1]), .A2(b[10]), .ZN(y[26]) );
  OR2_X1 U82bar ( .A1(abar[1]), .A2(bbar[10]), .ZN(ybar[26]);
  AND2_X1 U83 ( .A1(a[1]), .A2(b[9]), .ZN(y[25]) );
  OR2_X1 U83bar ( .A1(abar[1]), .A2(bbar[9]), .ZN(ybar[25]);
  AND2_X1 U84 ( .A1(a[15]), .A2(b[15]), .ZN(y[255]) );
  OR2_X1 U84bar ( .A1(abar[15]), .A2(bbar[15]), .ZN(ybar[255]);
  AND2_X1 U85 ( .A1(a[15]), .A2(b[14]), .ZN(y[254]) );
  OR2_X1 U85bar ( .A1(abar[15]), .A2(bbar[14]), .ZN(ybar[254]);
  AND2_X1 U86 ( .A1(a[15]), .A2(b[13]), .ZN(y[253]) );
  OR2_X1 U86bar ( .A1(abar[15]), .A2(bbar[13]), .ZN(ybar[253]);
  AND2_X1 U87 ( .A1(a[15]), .A2(b[12]), .ZN(y[252]) );
  OR2_X1 U87bar ( .A1(abar[15]), .A2(bbar[12]), .ZN(ybar[252]);
  AND2_X1 U88 ( .A1(a[15]), .A2(b[11]), .ZN(y[251]) );
  OR2_X1 U88bar ( .A1(abar[15]), .A2(bbar[11]), .ZN(ybar[251]);
  AND2_X1 U89 ( .A1(a[15]), .A2(b[10]), .ZN(y[250]) );
  OR2_X1 U89bar ( .A1(abar[15]), .A2(bbar[10]), .ZN(ybar[250]);
  AND2_X1 U90 ( .A1(a[1]), .A2(b[8]), .ZN(y[24]) );
  OR2_X1 U90bar ( .A1(abar[1]), .A2(bbar[8]), .ZN(ybar[24]);
  AND2_X1 U91 ( .A1(a[15]), .A2(b[9]), .ZN(y[249]) );
  OR2_X1 U91bar ( .A1(abar[15]), .A2(bbar[9]), .ZN(ybar[249]);
  AND2_X1 U92 ( .A1(a[15]), .A2(b[8]), .ZN(y[248]) );
  OR2_X1 U92bar ( .A1(abar[15]), .A2(bbar[8]), .ZN(ybar[248]);
  AND2_X1 U93 ( .A1(a[15]), .A2(b[7]), .ZN(y[247]) );
  OR2_X1 U93bar ( .A1(abar[15]), .A2(bbar[7]), .ZN(ybar[247]);
  AND2_X1 U94 ( .A1(a[15]), .A2(b[6]), .ZN(y[246]) );
  OR2_X1 U94bar ( .A1(abar[15]), .A2(bbar[6]), .ZN(ybar[246]);
  AND2_X1 U95 ( .A1(a[15]), .A2(b[5]), .ZN(y[245]) );
  OR2_X1 U95bar ( .A1(abar[15]), .A2(bbar[5]), .ZN(ybar[245]);
  AND2_X1 U96 ( .A1(a[15]), .A2(b[4]), .ZN(y[244]) );
  OR2_X1 U96bar ( .A1(abar[15]), .A2(bbar[4]), .ZN(ybar[244]);
  AND2_X1 U97 ( .A1(a[15]), .A2(b[3]), .ZN(y[243]) );
  OR2_X1 U97bar ( .A1(abar[15]), .A2(bbar[3]), .ZN(ybar[243]);
  AND2_X1 U98 ( .A1(a[15]), .A2(b[2]), .ZN(y[242]) );
  OR2_X1 U98bar ( .A1(abar[15]), .A2(bbar[2]), .ZN(ybar[242]);
  AND2_X1 U99 ( .A1(a[15]), .A2(b[1]), .ZN(y[241]) );
  OR2_X1 U99bar ( .A1(abar[15]), .A2(bbar[1]), .ZN(ybar[241]);
  AND2_X1 U100 ( .A1(a[15]), .A2(b[0]), .ZN(y[240]) );
  OR2_X1 U100bar ( .A1(abar[15]), .A2(bbar[0]), .ZN(ybar[240]);
  AND2_X1 U101 ( .A1(a[1]), .A2(b[7]), .ZN(y[23]) );
  OR2_X1 U101bar ( .A1(abar[1]), .A2(bbar[7]), .ZN(ybar[23]);
  AND2_X1 U102 ( .A1(a[14]), .A2(b[15]), .ZN(y[239]) );
  OR2_X1 U102bar ( .A1(abar[14]), .A2(bbar[15]), .ZN(ybar[239]);
  AND2_X1 U103 ( .A1(a[14]), .A2(b[14]), .ZN(y[238]) );
  OR2_X1 U103bar ( .A1(abar[14]), .A2(bbar[14]), .ZN(ybar[238]);
  AND2_X1 U104 ( .A1(a[14]), .A2(b[13]), .ZN(y[237]) );
  OR2_X1 U104bar ( .A1(abar[14]), .A2(bbar[13]), .ZN(ybar[237]);
  AND2_X1 U105 ( .A1(a[14]), .A2(b[12]), .ZN(y[236]) );
  OR2_X1 U105bar ( .A1(abar[14]), .A2(bbar[12]), .ZN(ybar[236]);
  AND2_X1 U106 ( .A1(a[14]), .A2(b[11]), .ZN(y[235]) );
  OR2_X1 U106bar ( .A1(abar[14]), .A2(bbar[11]), .ZN(ybar[235]);
  AND2_X1 U107 ( .A1(a[14]), .A2(b[10]), .ZN(y[234]) );
  OR2_X1 U107bar ( .A1(abar[14]), .A2(bbar[10]), .ZN(ybar[234]);
  AND2_X1 U108 ( .A1(a[14]), .A2(b[9]), .ZN(y[233]) );
  OR2_X1 U108bar ( .A1(abar[14]), .A2(bbar[9]), .ZN(ybar[233]);
  AND2_X1 U109 ( .A1(a[14]), .A2(b[8]), .ZN(y[232]) );
  OR2_X1 U109bar ( .A1(abar[14]), .A2(bbar[8]), .ZN(ybar[232]);
  AND2_X1 U110 ( .A1(a[14]), .A2(b[7]), .ZN(y[231]) );
  OR2_X1 U110bar ( .A1(abar[14]), .A2(bbar[7]), .ZN(ybar[231]);
  AND2_X1 U111 ( .A1(a[14]), .A2(b[6]), .ZN(y[230]) );
  OR2_X1 U111bar ( .A1(abar[14]), .A2(bbar[6]), .ZN(ybar[230]);
  AND2_X1 U112 ( .A1(a[1]), .A2(b[6]), .ZN(y[22]) );
  OR2_X1 U112bar ( .A1(abar[1]), .A2(bbar[6]), .ZN(ybar[22]);
  AND2_X1 U113 ( .A1(a[14]), .A2(b[5]), .ZN(y[229]) );
  OR2_X1 U113bar ( .A1(abar[14]), .A2(bbar[5]), .ZN(ybar[229]);
  AND2_X1 U114 ( .A1(a[14]), .A2(b[4]), .ZN(y[228]) );
  OR2_X1 U114bar ( .A1(abar[14]), .A2(bbar[4]), .ZN(ybar[228]);
  AND2_X1 U115 ( .A1(a[14]), .A2(b[3]), .ZN(y[227]) );
  OR2_X1 U115bar ( .A1(abar[14]), .A2(bbar[3]), .ZN(ybar[227]);
  AND2_X1 U116 ( .A1(a[14]), .A2(b[2]), .ZN(y[226]) );
  OR2_X1 U116bar ( .A1(abar[14]), .A2(bbar[2]), .ZN(ybar[226]);
  AND2_X1 U117 ( .A1(a[14]), .A2(b[1]), .ZN(y[225]) );
  OR2_X1 U117bar ( .A1(abar[14]), .A2(bbar[1]), .ZN(ybar[225]);
  AND2_X1 U118 ( .A1(a[14]), .A2(b[0]), .ZN(y[224]) );
  OR2_X1 U118bar ( .A1(abar[14]), .A2(bbar[0]), .ZN(ybar[224]);
  AND2_X1 U119 ( .A1(a[13]), .A2(b[15]), .ZN(y[223]) );
  OR2_X1 U119bar ( .A1(abar[13]), .A2(bbar[15]), .ZN(ybar[223]);
  AND2_X1 U120 ( .A1(a[13]), .A2(b[14]), .ZN(y[222]) );
  OR2_X1 U120bar ( .A1(abar[13]), .A2(bbar[14]), .ZN(ybar[222]);
  AND2_X1 U121 ( .A1(a[13]), .A2(b[13]), .ZN(y[221]) );
  OR2_X1 U121bar ( .A1(abar[13]), .A2(bbar[13]), .ZN(ybar[221]);
  AND2_X1 U122 ( .A1(a[13]), .A2(b[12]), .ZN(y[220]) );
  OR2_X1 U122bar ( .A1(abar[13]), .A2(bbar[12]), .ZN(ybar[220]);
  AND2_X1 U123 ( .A1(a[1]), .A2(b[5]), .ZN(y[21]) );
  OR2_X1 U123bar ( .A1(abar[1]), .A2(bbar[5]), .ZN(ybar[21]);
  AND2_X1 U124 ( .A1(a[13]), .A2(b[11]), .ZN(y[219]) );
  OR2_X1 U124bar ( .A1(abar[13]), .A2(bbar[11]), .ZN(ybar[219]);
  AND2_X1 U125 ( .A1(a[13]), .A2(b[10]), .ZN(y[218]) );
  OR2_X1 U125bar ( .A1(abar[13]), .A2(bbar[10]), .ZN(ybar[218]);
  AND2_X1 U126 ( .A1(a[13]), .A2(b[9]), .ZN(y[217]) );
  OR2_X1 U126bar ( .A1(abar[13]), .A2(bbar[9]), .ZN(ybar[217]);
  AND2_X1 U127 ( .A1(a[13]), .A2(b[8]), .ZN(y[216]) );
  OR2_X1 U127bar ( .A1(abar[13]), .A2(bbar[8]), .ZN(ybar[216]);
  AND2_X1 U128 ( .A1(a[13]), .A2(b[7]), .ZN(y[215]) );
  OR2_X1 U128bar ( .A1(abar[13]), .A2(bbar[7]), .ZN(ybar[215]);
  AND2_X1 U129 ( .A1(a[13]), .A2(b[6]), .ZN(y[214]) );
  OR2_X1 U129bar ( .A1(abar[13]), .A2(bbar[6]), .ZN(ybar[214]);
  AND2_X1 U130 ( .A1(a[13]), .A2(b[5]), .ZN(y[213]) );
  OR2_X1 U130bar ( .A1(abar[13]), .A2(bbar[5]), .ZN(ybar[213]);
  AND2_X1 U131 ( .A1(a[13]), .A2(b[4]), .ZN(y[212]) );
  OR2_X1 U131bar ( .A1(abar[13]), .A2(bbar[4]), .ZN(ybar[212]);
  AND2_X1 U132 ( .A1(a[13]), .A2(b[3]), .ZN(y[211]) );
  OR2_X1 U132bar ( .A1(abar[13]), .A2(bbar[3]), .ZN(ybar[211]);
  AND2_X1 U133 ( .A1(a[13]), .A2(b[2]), .ZN(y[210]) );
  OR2_X1 U133bar ( .A1(abar[13]), .A2(bbar[2]), .ZN(ybar[210]);
  AND2_X1 U134 ( .A1(a[1]), .A2(b[4]), .ZN(y[20]) );
  OR2_X1 U134bar ( .A1(abar[1]), .A2(bbar[4]), .ZN(ybar[20]);
  AND2_X1 U135 ( .A1(a[13]), .A2(b[1]), .ZN(y[209]) );
  OR2_X1 U135bar ( .A1(abar[13]), .A2(bbar[1]), .ZN(ybar[209]);
  AND2_X1 U136 ( .A1(a[13]), .A2(b[0]), .ZN(y[208]) );
  OR2_X1 U136bar ( .A1(abar[13]), .A2(bbar[0]), .ZN(ybar[208]);
  AND2_X1 U137 ( .A1(a[12]), .A2(b[15]), .ZN(y[207]) );
  OR2_X1 U137bar ( .A1(abar[12]), .A2(bbar[15]), .ZN(ybar[207]);
  AND2_X1 U138 ( .A1(a[12]), .A2(b[14]), .ZN(y[206]) );
  OR2_X1 U138bar ( .A1(abar[12]), .A2(bbar[14]), .ZN(ybar[206]);
  AND2_X1 U139 ( .A1(a[12]), .A2(b[13]), .ZN(y[205]) );
  OR2_X1 U139bar ( .A1(abar[12]), .A2(bbar[13]), .ZN(ybar[205]);
  AND2_X1 U140 ( .A1(a[12]), .A2(b[12]), .ZN(y[204]) );
  OR2_X1 U140bar ( .A1(abar[12]), .A2(bbar[12]), .ZN(ybar[204]);
  AND2_X1 U141 ( .A1(a[12]), .A2(b[11]), .ZN(y[203]) );
  OR2_X1 U141bar ( .A1(abar[12]), .A2(bbar[11]), .ZN(ybar[203]);
  AND2_X1 U142 ( .A1(a[12]), .A2(b[10]), .ZN(y[202]) );
  OR2_X1 U142bar ( .A1(abar[12]), .A2(bbar[10]), .ZN(ybar[202]);
  AND2_X1 U143 ( .A1(a[12]), .A2(b[9]), .ZN(y[201]) );
  OR2_X1 U143bar ( .A1(abar[12]), .A2(bbar[9]), .ZN(ybar[201]);
  AND2_X1 U144 ( .A1(a[12]), .A2(b[8]), .ZN(y[200]) );
  OR2_X1 U144bar ( .A1(abar[12]), .A2(bbar[8]), .ZN(ybar[200]);
  AND2_X1 U145 ( .A1(b[1]), .A2(a[0]), .ZN(y[1]) );
  OR2_X1 U145bar ( .A1(bbar[1]), .A2(abar[0]), .ZN(ybar[1]);
  AND2_X1 U146 ( .A1(a[1]), .A2(b[3]), .ZN(y[19]) );
  OR2_X1 U146bar ( .A1(abar[1]), .A2(bbar[3]), .ZN(ybar[19]);
  AND2_X1 U147 ( .A1(a[12]), .A2(b[7]), .ZN(y[199]) );
  OR2_X1 U147bar ( .A1(abar[12]), .A2(bbar[7]), .ZN(ybar[199]);
  AND2_X1 U148 ( .A1(a[12]), .A2(b[6]), .ZN(y[198]) );
  OR2_X1 U148bar ( .A1(abar[12]), .A2(bbar[6]), .ZN(ybar[198]);
  AND2_X1 U149 ( .A1(a[12]), .A2(b[5]), .ZN(y[197]) );
  OR2_X1 U149bar ( .A1(abar[12]), .A2(bbar[5]), .ZN(ybar[197]);
  AND2_X1 U150 ( .A1(a[12]), .A2(b[4]), .ZN(y[196]) );
  OR2_X1 U150bar ( .A1(abar[12]), .A2(bbar[4]), .ZN(ybar[196]);
  AND2_X1 U151 ( .A1(a[12]), .A2(b[3]), .ZN(y[195]) );
  OR2_X1 U151bar ( .A1(abar[12]), .A2(bbar[3]), .ZN(ybar[195]);
  AND2_X1 U152 ( .A1(a[12]), .A2(b[2]), .ZN(y[194]) );
  OR2_X1 U152bar ( .A1(abar[12]), .A2(bbar[2]), .ZN(ybar[194]);
  AND2_X1 U153 ( .A1(a[12]), .A2(b[1]), .ZN(y[193]) );
  OR2_X1 U153bar ( .A1(abar[12]), .A2(bbar[1]), .ZN(ybar[193]);
  AND2_X1 U154 ( .A1(a[12]), .A2(b[0]), .ZN(y[192]) );
  OR2_X1 U154bar ( .A1(abar[12]), .A2(bbar[0]), .ZN(ybar[192]);
  AND2_X1 U155 ( .A1(a[11]), .A2(b[15]), .ZN(y[191]) );
  OR2_X1 U155bar ( .A1(abar[11]), .A2(bbar[15]), .ZN(ybar[191]);
  AND2_X1 U156 ( .A1(a[11]), .A2(b[14]), .ZN(y[190]) );
  OR2_X1 U156bar ( .A1(abar[11]), .A2(bbar[14]), .ZN(ybar[190]);
  AND2_X1 U157 ( .A1(a[1]), .A2(b[2]), .ZN(y[18]) );
  OR2_X1 U157bar ( .A1(abar[1]), .A2(bbar[2]), .ZN(ybar[18]);
  AND2_X1 U158 ( .A1(a[11]), .A2(b[13]), .ZN(y[189]) );
  OR2_X1 U158bar ( .A1(abar[11]), .A2(bbar[13]), .ZN(ybar[189]);
  AND2_X1 U159 ( .A1(a[11]), .A2(b[12]), .ZN(y[188]) );
  OR2_X1 U159bar ( .A1(abar[11]), .A2(bbar[12]), .ZN(ybar[188]);
  AND2_X1 U160 ( .A1(a[11]), .A2(b[11]), .ZN(y[187]) );
  OR2_X1 U160bar ( .A1(abar[11]), .A2(bbar[11]), .ZN(ybar[187]);
  AND2_X1 U161 ( .A1(a[11]), .A2(b[10]), .ZN(y[186]) );
  OR2_X1 U161bar ( .A1(abar[11]), .A2(bbar[10]), .ZN(ybar[186]);
  AND2_X1 U162 ( .A1(a[11]), .A2(b[9]), .ZN(y[185]) );
  OR2_X1 U162bar ( .A1(abar[11]), .A2(bbar[9]), .ZN(ybar[185]);
  AND2_X1 U163 ( .A1(a[11]), .A2(b[8]), .ZN(y[184]) );
  OR2_X1 U163bar ( .A1(abar[11]), .A2(bbar[8]), .ZN(ybar[184]);
  AND2_X1 U164 ( .A1(a[11]), .A2(b[7]), .ZN(y[183]) );
  OR2_X1 U164bar ( .A1(abar[11]), .A2(bbar[7]), .ZN(ybar[183]);
  AND2_X1 U165 ( .A1(a[11]), .A2(b[6]), .ZN(y[182]) );
  OR2_X1 U165bar ( .A1(abar[11]), .A2(bbar[6]), .ZN(ybar[182]);
  AND2_X1 U166 ( .A1(a[11]), .A2(b[5]), .ZN(y[181]) );
  OR2_X1 U166bar ( .A1(abar[11]), .A2(bbar[5]), .ZN(ybar[181]);
  AND2_X1 U167 ( .A1(a[11]), .A2(b[4]), .ZN(y[180]) );
  OR2_X1 U167bar ( .A1(abar[11]), .A2(bbar[4]), .ZN(ybar[180]);
  AND2_X1 U168 ( .A1(a[1]), .A2(b[1]), .ZN(y[17]) );
  OR2_X1 U168bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[17]);
  AND2_X1 U169 ( .A1(a[11]), .A2(b[3]), .ZN(y[179]) );
  OR2_X1 U169bar ( .A1(abar[11]), .A2(bbar[3]), .ZN(ybar[179]);
  AND2_X1 U170 ( .A1(a[11]), .A2(b[2]), .ZN(y[178]) );
  OR2_X1 U170bar ( .A1(abar[11]), .A2(bbar[2]), .ZN(ybar[178]);
  AND2_X1 U171 ( .A1(a[11]), .A2(b[1]), .ZN(y[177]) );
  OR2_X1 U171bar ( .A1(abar[11]), .A2(bbar[1]), .ZN(ybar[177]);
  AND2_X1 U172 ( .A1(a[11]), .A2(b[0]), .ZN(y[176]) );
  OR2_X1 U172bar ( .A1(abar[11]), .A2(bbar[0]), .ZN(ybar[176]);
  AND2_X1 U173 ( .A1(a[10]), .A2(b[15]), .ZN(y[175]) );
  OR2_X1 U173bar ( .A1(abar[10]), .A2(bbar[15]), .ZN(ybar[175]);
  AND2_X1 U174 ( .A1(a[10]), .A2(b[14]), .ZN(y[174]) );
  OR2_X1 U174bar ( .A1(abar[10]), .A2(bbar[14]), .ZN(ybar[174]);
  AND2_X1 U175 ( .A1(a[10]), .A2(b[13]), .ZN(y[173]) );
  OR2_X1 U175bar ( .A1(abar[10]), .A2(bbar[13]), .ZN(ybar[173]);
  AND2_X1 U176 ( .A1(a[10]), .A2(b[12]), .ZN(y[172]) );
  OR2_X1 U176bar ( .A1(abar[10]), .A2(bbar[12]), .ZN(ybar[172]);
  AND2_X1 U177 ( .A1(a[10]), .A2(b[11]), .ZN(y[171]) );
  OR2_X1 U177bar ( .A1(abar[10]), .A2(bbar[11]), .ZN(ybar[171]);
  AND2_X1 U178 ( .A1(a[10]), .A2(b[10]), .ZN(y[170]) );
  OR2_X1 U178bar ( .A1(abar[10]), .A2(bbar[10]), .ZN(ybar[170]);
  AND2_X1 U179 ( .A1(a[1]), .A2(b[0]), .ZN(y[16]) );
  OR2_X1 U179bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[16]);
  AND2_X1 U180 ( .A1(a[10]), .A2(b[9]), .ZN(y[169]) );
  OR2_X1 U180bar ( .A1(abar[10]), .A2(bbar[9]), .ZN(ybar[169]);
  AND2_X1 U181 ( .A1(a[10]), .A2(b[8]), .ZN(y[168]) );
  OR2_X1 U181bar ( .A1(abar[10]), .A2(bbar[8]), .ZN(ybar[168]);
  AND2_X1 U182 ( .A1(a[10]), .A2(b[7]), .ZN(y[167]) );
  OR2_X1 U182bar ( .A1(abar[10]), .A2(bbar[7]), .ZN(ybar[167]);
  AND2_X1 U183 ( .A1(a[10]), .A2(b[6]), .ZN(y[166]) );
  OR2_X1 U183bar ( .A1(abar[10]), .A2(bbar[6]), .ZN(ybar[166]);
  AND2_X1 U184 ( .A1(a[10]), .A2(b[5]), .ZN(y[165]) );
  OR2_X1 U184bar ( .A1(abar[10]), .A2(bbar[5]), .ZN(ybar[165]);
  AND2_X1 U185 ( .A1(a[10]), .A2(b[4]), .ZN(y[164]) );
  OR2_X1 U185bar ( .A1(abar[10]), .A2(bbar[4]), .ZN(ybar[164]);
  AND2_X1 U186 ( .A1(a[10]), .A2(b[3]), .ZN(y[163]) );
  OR2_X1 U186bar ( .A1(abar[10]), .A2(bbar[3]), .ZN(ybar[163]);
  AND2_X1 U187 ( .A1(a[10]), .A2(b[2]), .ZN(y[162]) );
  OR2_X1 U187bar ( .A1(abar[10]), .A2(bbar[2]), .ZN(ybar[162]);
  AND2_X1 U188 ( .A1(a[10]), .A2(b[1]), .ZN(y[161]) );
  OR2_X1 U188bar ( .A1(abar[10]), .A2(bbar[1]), .ZN(ybar[161]);
  AND2_X1 U189 ( .A1(a[10]), .A2(b[0]), .ZN(y[160]) );
  OR2_X1 U189bar ( .A1(abar[10]), .A2(bbar[0]), .ZN(ybar[160]);
  AND2_X1 U190 ( .A1(b[15]), .A2(a[0]), .ZN(y[15]) );
  OR2_X1 U190bar ( .A1(bbar[15]), .A2(abar[0]), .ZN(ybar[15]);
  AND2_X1 U191 ( .A1(a[9]), .A2(b[15]), .ZN(y[159]) );
  OR2_X1 U191bar ( .A1(abar[9]), .A2(bbar[15]), .ZN(ybar[159]);
  AND2_X1 U192 ( .A1(a[9]), .A2(b[14]), .ZN(y[158]) );
  OR2_X1 U192bar ( .A1(abar[9]), .A2(bbar[14]), .ZN(ybar[158]);
  AND2_X1 U193 ( .A1(a[9]), .A2(b[13]), .ZN(y[157]) );
  OR2_X1 U193bar ( .A1(abar[9]), .A2(bbar[13]), .ZN(ybar[157]);
  AND2_X1 U194 ( .A1(a[9]), .A2(b[12]), .ZN(y[156]) );
  OR2_X1 U194bar ( .A1(abar[9]), .A2(bbar[12]), .ZN(ybar[156]);
  AND2_X1 U195 ( .A1(a[9]), .A2(b[11]), .ZN(y[155]) );
  OR2_X1 U195bar ( .A1(abar[9]), .A2(bbar[11]), .ZN(ybar[155]);
  AND2_X1 U196 ( .A1(a[9]), .A2(b[10]), .ZN(y[154]) );
  OR2_X1 U196bar ( .A1(abar[9]), .A2(bbar[10]), .ZN(ybar[154]);
  AND2_X1 U197 ( .A1(a[9]), .A2(b[9]), .ZN(y[153]) );
  OR2_X1 U197bar ( .A1(abar[9]), .A2(bbar[9]), .ZN(ybar[153]);
  AND2_X1 U198 ( .A1(a[9]), .A2(b[8]), .ZN(y[152]) );
  OR2_X1 U198bar ( .A1(abar[9]), .A2(bbar[8]), .ZN(ybar[152]);
  AND2_X1 U199 ( .A1(a[9]), .A2(b[7]), .ZN(y[151]) );
  OR2_X1 U199bar ( .A1(abar[9]), .A2(bbar[7]), .ZN(ybar[151]);
  AND2_X1 U200 ( .A1(a[9]), .A2(b[6]), .ZN(y[150]) );
  OR2_X1 U200bar ( .A1(abar[9]), .A2(bbar[6]), .ZN(ybar[150]);
  AND2_X1 U201 ( .A1(b[14]), .A2(a[0]), .ZN(y[14]) );
  OR2_X1 U201bar ( .A1(bbar[14]), .A2(abar[0]), .ZN(ybar[14]);
  AND2_X1 U202 ( .A1(a[9]), .A2(b[5]), .ZN(y[149]) );
  OR2_X1 U202bar ( .A1(abar[9]), .A2(bbar[5]), .ZN(ybar[149]);
  AND2_X1 U203 ( .A1(a[9]), .A2(b[4]), .ZN(y[148]) );
  OR2_X1 U203bar ( .A1(abar[9]), .A2(bbar[4]), .ZN(ybar[148]);
  AND2_X1 U204 ( .A1(a[9]), .A2(b[3]), .ZN(y[147]) );
  OR2_X1 U204bar ( .A1(abar[9]), .A2(bbar[3]), .ZN(ybar[147]);
  AND2_X1 U205 ( .A1(a[9]), .A2(b[2]), .ZN(y[146]) );
  OR2_X1 U205bar ( .A1(abar[9]), .A2(bbar[2]), .ZN(ybar[146]);
  AND2_X1 U206 ( .A1(a[9]), .A2(b[1]), .ZN(y[145]) );
  OR2_X1 U206bar ( .A1(abar[9]), .A2(bbar[1]), .ZN(ybar[145]);
  AND2_X1 U207 ( .A1(a[9]), .A2(b[0]), .ZN(y[144]) );
  OR2_X1 U207bar ( .A1(abar[9]), .A2(bbar[0]), .ZN(ybar[144]);
  AND2_X1 U208 ( .A1(a[8]), .A2(b[15]), .ZN(y[143]) );
  OR2_X1 U208bar ( .A1(abar[8]), .A2(bbar[15]), .ZN(ybar[143]);
  AND2_X1 U209 ( .A1(a[8]), .A2(b[14]), .ZN(y[142]) );
  OR2_X1 U209bar ( .A1(abar[8]), .A2(bbar[14]), .ZN(ybar[142]);
  AND2_X1 U210 ( .A1(a[8]), .A2(b[13]), .ZN(y[141]) );
  OR2_X1 U210bar ( .A1(abar[8]), .A2(bbar[13]), .ZN(ybar[141]);
  AND2_X1 U211 ( .A1(a[8]), .A2(b[12]), .ZN(y[140]) );
  OR2_X1 U211bar ( .A1(abar[8]), .A2(bbar[12]), .ZN(ybar[140]);
  AND2_X1 U212 ( .A1(b[13]), .A2(a[0]), .ZN(y[13]) );
  OR2_X1 U212bar ( .A1(bbar[13]), .A2(abar[0]), .ZN(ybar[13]);
  AND2_X1 U213 ( .A1(a[8]), .A2(b[11]), .ZN(y[139]) );
  OR2_X1 U213bar ( .A1(abar[8]), .A2(bbar[11]), .ZN(ybar[139]);
  AND2_X1 U214 ( .A1(a[8]), .A2(b[10]), .ZN(y[138]) );
  OR2_X1 U214bar ( .A1(abar[8]), .A2(bbar[10]), .ZN(ybar[138]);
  AND2_X1 U215 ( .A1(a[8]), .A2(b[9]), .ZN(y[137]) );
  OR2_X1 U215bar ( .A1(abar[8]), .A2(bbar[9]), .ZN(ybar[137]);
  AND2_X1 U216 ( .A1(a[8]), .A2(b[8]), .ZN(y[136]) );
  OR2_X1 U216bar ( .A1(abar[8]), .A2(bbar[8]), .ZN(ybar[136]);
  AND2_X1 U217 ( .A1(a[8]), .A2(b[7]), .ZN(y[135]) );
  OR2_X1 U217bar ( .A1(abar[8]), .A2(bbar[7]), .ZN(ybar[135]);
  AND2_X1 U218 ( .A1(a[8]), .A2(b[6]), .ZN(y[134]) );
  OR2_X1 U218bar ( .A1(abar[8]), .A2(bbar[6]), .ZN(ybar[134]);
  AND2_X1 U219 ( .A1(a[8]), .A2(b[5]), .ZN(y[133]) );
  OR2_X1 U219bar ( .A1(abar[8]), .A2(bbar[5]), .ZN(ybar[133]);
  AND2_X1 U220 ( .A1(a[8]), .A2(b[4]), .ZN(y[132]) );
  OR2_X1 U220bar ( .A1(abar[8]), .A2(bbar[4]), .ZN(ybar[132]);
  AND2_X1 U221 ( .A1(a[8]), .A2(b[3]), .ZN(y[131]) );
  OR2_X1 U221bar ( .A1(abar[8]), .A2(bbar[3]), .ZN(ybar[131]);
  AND2_X1 U222 ( .A1(a[8]), .A2(b[2]), .ZN(y[130]) );
  OR2_X1 U222bar ( .A1(abar[8]), .A2(bbar[2]), .ZN(ybar[130]);
  AND2_X1 U223 ( .A1(b[12]), .A2(a[0]), .ZN(y[12]) );
  OR2_X1 U223bar ( .A1(bbar[12]), .A2(abar[0]), .ZN(ybar[12]);
  AND2_X1 U224 ( .A1(a[8]), .A2(b[1]), .ZN(y[129]) );
  OR2_X1 U224bar ( .A1(abar[8]), .A2(bbar[1]), .ZN(ybar[129]);
  AND2_X1 U225 ( .A1(a[8]), .A2(b[0]), .ZN(y[128]) );
  OR2_X1 U225bar ( .A1(abar[8]), .A2(bbar[0]), .ZN(ybar[128]);
  AND2_X1 U226 ( .A1(a[7]), .A2(b[15]), .ZN(y[127]) );
  OR2_X1 U226bar ( .A1(abar[7]), .A2(bbar[15]), .ZN(ybar[127]);
  AND2_X1 U227 ( .A1(a[7]), .A2(b[14]), .ZN(y[126]) );
  OR2_X1 U227bar ( .A1(abar[7]), .A2(bbar[14]), .ZN(ybar[126]);
  AND2_X1 U228 ( .A1(a[7]), .A2(b[13]), .ZN(y[125]) );
  OR2_X1 U228bar ( .A1(abar[7]), .A2(bbar[13]), .ZN(ybar[125]);
  AND2_X1 U229 ( .A1(a[7]), .A2(b[12]), .ZN(y[124]) );
  OR2_X1 U229bar ( .A1(abar[7]), .A2(bbar[12]), .ZN(ybar[124]);
  AND2_X1 U230 ( .A1(a[7]), .A2(b[11]), .ZN(y[123]) );
  OR2_X1 U230bar ( .A1(abar[7]), .A2(bbar[11]), .ZN(ybar[123]);
  AND2_X1 U231 ( .A1(a[7]), .A2(b[10]), .ZN(y[122]) );
  OR2_X1 U231bar ( .A1(abar[7]), .A2(bbar[10]), .ZN(ybar[122]);
  AND2_X1 U232 ( .A1(a[7]), .A2(b[9]), .ZN(y[121]) );
  OR2_X1 U232bar ( .A1(abar[7]), .A2(bbar[9]), .ZN(ybar[121]);
  AND2_X1 U233 ( .A1(a[7]), .A2(b[8]), .ZN(y[120]) );
  OR2_X1 U233bar ( .A1(abar[7]), .A2(bbar[8]), .ZN(ybar[120]);
  AND2_X1 U234 ( .A1(b[11]), .A2(a[0]), .ZN(y[11]) );
  OR2_X1 U234bar ( .A1(bbar[11]), .A2(abar[0]), .ZN(ybar[11]);
  AND2_X1 U235 ( .A1(a[7]), .A2(b[7]), .ZN(y[119]) );
  OR2_X1 U235bar ( .A1(abar[7]), .A2(bbar[7]), .ZN(ybar[119]);
  AND2_X1 U236 ( .A1(a[7]), .A2(b[6]), .ZN(y[118]) );
  OR2_X1 U236bar ( .A1(abar[7]), .A2(bbar[6]), .ZN(ybar[118]);
  AND2_X1 U237 ( .A1(a[7]), .A2(b[5]), .ZN(y[117]) );
  OR2_X1 U237bar ( .A1(abar[7]), .A2(bbar[5]), .ZN(ybar[117]);
  AND2_X1 U238 ( .A1(a[7]), .A2(b[4]), .ZN(y[116]) );
  OR2_X1 U238bar ( .A1(abar[7]), .A2(bbar[4]), .ZN(ybar[116]);
  AND2_X1 U239 ( .A1(a[7]), .A2(b[3]), .ZN(y[115]) );
  OR2_X1 U239bar ( .A1(abar[7]), .A2(bbar[3]), .ZN(ybar[115]);
  AND2_X1 U240 ( .A1(a[7]), .A2(b[2]), .ZN(y[114]) );
  OR2_X1 U240bar ( .A1(abar[7]), .A2(bbar[2]), .ZN(ybar[114]);
  AND2_X1 U241 ( .A1(a[7]), .A2(b[1]), .ZN(y[113]) );
  OR2_X1 U241bar ( .A1(abar[7]), .A2(bbar[1]), .ZN(ybar[113]);
  AND2_X1 U242 ( .A1(a[7]), .A2(b[0]), .ZN(y[112]) );
  OR2_X1 U242bar ( .A1(abar[7]), .A2(bbar[0]), .ZN(ybar[112]);
  AND2_X1 U243 ( .A1(b[15]), .A2(a[6]), .ZN(y[111]) );
  OR2_X1 U243bar ( .A1(bbar[15]), .A2(abar[6]), .ZN(ybar[111]);
  AND2_X1 U244 ( .A1(b[14]), .A2(a[6]), .ZN(y[110]) );
  OR2_X1 U244bar ( .A1(bbar[14]), .A2(abar[6]), .ZN(ybar[110]);
  AND2_X1 U245 ( .A1(b[10]), .A2(a[0]), .ZN(y[10]) );
  OR2_X1 U245bar ( .A1(bbar[10]), .A2(abar[0]), .ZN(ybar[10]);
  AND2_X1 U246 ( .A1(b[13]), .A2(a[6]), .ZN(y[109]) );
  OR2_X1 U246bar ( .A1(bbar[13]), .A2(abar[6]), .ZN(ybar[109]);
  AND2_X1 U247 ( .A1(b[12]), .A2(a[6]), .ZN(y[108]) );
  OR2_X1 U247bar ( .A1(bbar[12]), .A2(abar[6]), .ZN(ybar[108]);
  AND2_X1 U248 ( .A1(b[11]), .A2(a[6]), .ZN(y[107]) );
  OR2_X1 U248bar ( .A1(bbar[11]), .A2(abar[6]), .ZN(ybar[107]);
  AND2_X1 U249 ( .A1(b[10]), .A2(a[6]), .ZN(y[106]) );
  OR2_X1 U249bar ( .A1(bbar[10]), .A2(abar[6]), .ZN(ybar[106]);
  AND2_X1 U250 ( .A1(a[6]), .A2(b[9]), .ZN(y[105]) );
  OR2_X1 U250bar ( .A1(abar[6]), .A2(bbar[9]), .ZN(ybar[105]);
  AND2_X1 U251 ( .A1(b[8]), .A2(a[6]), .ZN(y[104]) );
  OR2_X1 U251bar ( .A1(bbar[8]), .A2(abar[6]), .ZN(ybar[104]);
  AND2_X1 U252 ( .A1(b[7]), .A2(a[6]), .ZN(y[103]) );
  OR2_X1 U252bar ( .A1(bbar[7]), .A2(abar[6]), .ZN(ybar[103]);
  AND2_X1 U253 ( .A1(b[6]), .A2(a[6]), .ZN(y[102]) );
  OR2_X1 U253bar ( .A1(bbar[6]), .A2(abar[6]), .ZN(ybar[102]);
  AND2_X1 U254 ( .A1(b[5]), .A2(a[6]), .ZN(y[101]) );
  OR2_X1 U254bar ( .A1(bbar[5]), .A2(abar[6]), .ZN(ybar[101]);
  AND2_X1 U255 ( .A1(b[4]), .A2(a[6]), .ZN(y[100]) );
  OR2_X1 U255bar ( .A1(bbar[4]), .A2(abar[6]), .ZN(ybar[100]);
  AND2_X1 U256 ( .A1(b[0]), .A2(a[0]), .ZN(y[0]) );
  OR2_X1 U256bar ( .A1(bbar[0]), .A2(abar[0]), .ZN(ybar[0]);
endmodule




module decode_9 ( in, out );
  input [7:0] in;
  //input_done

  output [255:0] out;
  //output_done

  wire   [15:0] level1;
  wire   [31:0] level2;
  //wire_done

  CD2_36 cd_l1_1 ( .a(in[1]), .b(in[0]), .y(level1[3:0]) );
  CD2_35 cd_l1_2 ( .a(in[3]), .b(in[2]), .y(level1[7:4]) );
  CD2_34 cd_l1_3 ( .a(in[5]), .b(in[4]), .y(level1[11:8]) );
  CD2_33 cd_l1_4 ( .a(in[7]), .b(in[6]), .y(level1[15:12]) );
  CD4_18 cd_l2_1 ( .a(level1[7:4]), .b(level1[3:0]), .y(level2[15:0]) );
  CD4_17 cd_l2_2 ( .a(level1[15:12]), .b(level1[11:8]), .y(level2[31:16]) );
  CD16_9 cd_l3 ( .a(level2[31:16]), .b(level2[15:0]), .y(out) );
endmodule


module encode_9 ( in, out );
  input [255:0] in;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
  assign inbar[8] = ~in[8];
  assign inbar[9] = ~in[9];
  assign inbar[10] = ~in[10];
  assign inbar[11] = ~in[11];
  assign inbar[12] = ~in[12];
  assign inbar[13] = ~in[13];
  assign inbar[14] = ~in[14];
  assign inbar[15] = ~in[15];
  assign inbar[16] = ~in[16];
  assign inbar[17] = ~in[17];
  assign inbar[18] = ~in[18];
  assign inbar[19] = ~in[19];
  assign inbar[20] = ~in[20];
  assign inbar[21] = ~in[21];
  assign inbar[22] = ~in[22];
  assign inbar[23] = ~in[23];
  assign inbar[24] = ~in[24];
  assign inbar[25] = ~in[25];
  assign inbar[26] = ~in[26];
  assign inbar[27] = ~in[27];
  assign inbar[28] = ~in[28];
  assign inbar[29] = ~in[29];
  assign inbar[30] = ~in[30];
  assign inbar[31] = ~in[31];
  assign inbar[32] = ~in[32];
  assign inbar[33] = ~in[33];
  assign inbar[34] = ~in[34];
  assign inbar[35] = ~in[35];
  assign inbar[36] = ~in[36];
  assign inbar[37] = ~in[37];
  assign inbar[38] = ~in[38];
  assign inbar[39] = ~in[39];
  assign inbar[40] = ~in[40];
  assign inbar[41] = ~in[41];
  assign inbar[42] = ~in[42];
  assign inbar[43] = ~in[43];
  assign inbar[44] = ~in[44];
  assign inbar[45] = ~in[45];
  assign inbar[46] = ~in[46];
  assign inbar[47] = ~in[47];
  assign inbar[48] = ~in[48];
  assign inbar[49] = ~in[49];
  assign inbar[50] = ~in[50];
  assign inbar[51] = ~in[51];
  assign inbar[52] = ~in[52];
  assign inbar[53] = ~in[53];
  assign inbar[54] = ~in[54];
  assign inbar[55] = ~in[55];
  assign inbar[56] = ~in[56];
  assign inbar[57] = ~in[57];
  assign inbar[58] = ~in[58];
  assign inbar[59] = ~in[59];
  assign inbar[60] = ~in[60];
  assign inbar[61] = ~in[61];
  assign inbar[62] = ~in[62];
  assign inbar[63] = ~in[63];
  assign inbar[64] = ~in[64];
  assign inbar[65] = ~in[65];
  assign inbar[66] = ~in[66];
  assign inbar[67] = ~in[67];
  assign inbar[68] = ~in[68];
  assign inbar[69] = ~in[69];
  assign inbar[70] = ~in[70];
  assign inbar[71] = ~in[71];
  assign inbar[72] = ~in[72];
  assign inbar[73] = ~in[73];
  assign inbar[74] = ~in[74];
  assign inbar[75] = ~in[75];
  assign inbar[76] = ~in[76];
  assign inbar[77] = ~in[77];
  assign inbar[78] = ~in[78];
  assign inbar[79] = ~in[79];
  assign inbar[80] = ~in[80];
  assign inbar[81] = ~in[81];
  assign inbar[82] = ~in[82];
  assign inbar[83] = ~in[83];
  assign inbar[84] = ~in[84];
  assign inbar[85] = ~in[85];
  assign inbar[86] = ~in[86];
  assign inbar[87] = ~in[87];
  assign inbar[88] = ~in[88];
  assign inbar[89] = ~in[89];
  assign inbar[90] = ~in[90];
  assign inbar[91] = ~in[91];
  assign inbar[92] = ~in[92];
  assign inbar[93] = ~in[93];
  assign inbar[94] = ~in[94];
  assign inbar[95] = ~in[95];
  assign inbar[96] = ~in[96];
  assign inbar[97] = ~in[97];
  assign inbar[98] = ~in[98];
  assign inbar[99] = ~in[99];
  assign inbar[100] = ~in[100];
  assign inbar[101] = ~in[101];
  assign inbar[102] = ~in[102];
  assign inbar[103] = ~in[103];
  assign inbar[104] = ~in[104];
  assign inbar[105] = ~in[105];
  assign inbar[106] = ~in[106];
  assign inbar[107] = ~in[107];
  assign inbar[108] = ~in[108];
  assign inbar[109] = ~in[109];
  assign inbar[110] = ~in[110];
  assign inbar[111] = ~in[111];
  assign inbar[112] = ~in[112];
  assign inbar[113] = ~in[113];
  assign inbar[114] = ~in[114];
  assign inbar[115] = ~in[115];
  assign inbar[116] = ~in[116];
  assign inbar[117] = ~in[117];
  assign inbar[118] = ~in[118];
  assign inbar[119] = ~in[119];
  assign inbar[120] = ~in[120];
  assign inbar[121] = ~in[121];
  assign inbar[122] = ~in[122];
  assign inbar[123] = ~in[123];
  assign inbar[124] = ~in[124];
  assign inbar[125] = ~in[125];
  assign inbar[126] = ~in[126];
  assign inbar[127] = ~in[127];
  assign inbar[128] = ~in[128];
  assign inbar[129] = ~in[129];
  assign inbar[130] = ~in[130];
  assign inbar[131] = ~in[131];
  assign inbar[132] = ~in[132];
  assign inbar[133] = ~in[133];
  assign inbar[134] = ~in[134];
  assign inbar[135] = ~in[135];
  assign inbar[136] = ~in[136];
  assign inbar[137] = ~in[137];
  assign inbar[138] = ~in[138];
  assign inbar[139] = ~in[139];
  assign inbar[140] = ~in[140];
  assign inbar[141] = ~in[141];
  assign inbar[142] = ~in[142];
  assign inbar[143] = ~in[143];
  assign inbar[144] = ~in[144];
  assign inbar[145] = ~in[145];
  assign inbar[146] = ~in[146];
  assign inbar[147] = ~in[147];
  assign inbar[148] = ~in[148];
  assign inbar[149] = ~in[149];
  assign inbar[150] = ~in[150];
  assign inbar[151] = ~in[151];
  assign inbar[152] = ~in[152];
  assign inbar[153] = ~in[153];
  assign inbar[154] = ~in[154];
  assign inbar[155] = ~in[155];
  assign inbar[156] = ~in[156];
  assign inbar[157] = ~in[157];
  assign inbar[158] = ~in[158];
  assign inbar[159] = ~in[159];
  assign inbar[160] = ~in[160];
  assign inbar[161] = ~in[161];
  assign inbar[162] = ~in[162];
  assign inbar[163] = ~in[163];
  assign inbar[164] = ~in[164];
  assign inbar[165] = ~in[165];
  assign inbar[166] = ~in[166];
  assign inbar[167] = ~in[167];
  assign inbar[168] = ~in[168];
  assign inbar[169] = ~in[169];
  assign inbar[170] = ~in[170];
  assign inbar[171] = ~in[171];
  assign inbar[172] = ~in[172];
  assign inbar[173] = ~in[173];
  assign inbar[174] = ~in[174];
  assign inbar[175] = ~in[175];
  assign inbar[176] = ~in[176];
  assign inbar[177] = ~in[177];
  assign inbar[178] = ~in[178];
  assign inbar[179] = ~in[179];
  assign inbar[180] = ~in[180];
  assign inbar[181] = ~in[181];
  assign inbar[182] = ~in[182];
  assign inbar[183] = ~in[183];
  assign inbar[184] = ~in[184];
  assign inbar[185] = ~in[185];
  assign inbar[186] = ~in[186];
  assign inbar[187] = ~in[187];
  assign inbar[188] = ~in[188];
  assign inbar[189] = ~in[189];
  assign inbar[190] = ~in[190];
  assign inbar[191] = ~in[191];
  assign inbar[192] = ~in[192];
  assign inbar[193] = ~in[193];
  assign inbar[194] = ~in[194];
  assign inbar[195] = ~in[195];
  assign inbar[196] = ~in[196];
  assign inbar[197] = ~in[197];
  assign inbar[198] = ~in[198];
  assign inbar[199] = ~in[199];
  assign inbar[200] = ~in[200];
  assign inbar[201] = ~in[201];
  assign inbar[202] = ~in[202];
  assign inbar[203] = ~in[203];
  assign inbar[204] = ~in[204];
  assign inbar[205] = ~in[205];
  assign inbar[206] = ~in[206];
  assign inbar[207] = ~in[207];
  assign inbar[208] = ~in[208];
  assign inbar[209] = ~in[209];
  assign inbar[210] = ~in[210];
  assign inbar[211] = ~in[211];
  assign inbar[212] = ~in[212];
  assign inbar[213] = ~in[213];
  assign inbar[214] = ~in[214];
  assign inbar[215] = ~in[215];
  assign inbar[216] = ~in[216];
  assign inbar[217] = ~in[217];
  assign inbar[218] = ~in[218];
  assign inbar[219] = ~in[219];
  assign inbar[220] = ~in[220];
  assign inbar[221] = ~in[221];
  assign inbar[222] = ~in[222];
  assign inbar[223] = ~in[223];
  assign inbar[224] = ~in[224];
  assign inbar[225] = ~in[225];
  assign inbar[226] = ~in[226];
  assign inbar[227] = ~in[227];
  assign inbar[228] = ~in[228];
  assign inbar[229] = ~in[229];
  assign inbar[230] = ~in[230];
  assign inbar[231] = ~in[231];
  assign inbar[232] = ~in[232];
  assign inbar[233] = ~in[233];
  assign inbar[234] = ~in[234];
  assign inbar[235] = ~in[235];
  assign inbar[236] = ~in[236];
  assign inbar[237] = ~in[237];
  assign inbar[238] = ~in[238];
  assign inbar[239] = ~in[239];
  assign inbar[240] = ~in[240];
  assign inbar[241] = ~in[241];
  assign inbar[242] = ~in[242];
  assign inbar[243] = ~in[243];
  assign inbar[244] = ~in[244];
  assign inbar[245] = ~in[245];
  assign inbar[246] = ~in[246];
  assign inbar[247] = ~in[247];
  assign inbar[248] = ~in[248];
  assign inbar[249] = ~in[249];
  assign inbar[250] = ~in[250];
  assign inbar[251] = ~in[251];
  assign inbar[252] = ~in[252];
  assign inbar[253] = ~in[253];
  assign inbar[254] = ~in[254];
  assign inbar[255] = ~in[255];
  //input_done

  output [7:0] out;
  reg [7:0] outbar;
  //output_done

  wire   in_81, in_80, in_79, in_78, in_77, in_76, in_75, in_74, in_73, in_72,
         in_71, in_70, in_69, in_68, in_67, in_66, in_65, in_64, in_63, in_62,
         in_61, in_60, in_59, in_58, in_57, in_56, in_55, in_54, in_53, in_52,
         in_51, in_50, in_49, in_48, in_47, in_46, in_45, in_44, in_43, in_42,
         in_41, in_40, in_39, in_38, in_37, in_36, in_35, in_34, in_33, in_32,
         in_31, in_30, in_29, in_28, in_27, in_26, in_25, in_24, in_23, in_22,
         in_21, in_20, in_19, in_18, in_17, in_16, in_15, in_14, in_13, in_12,
         in_11, in_10, in_9, in_8, in_7, in_6, in_5, in_4, in_3, in_2, in_1,
         in_0, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972;
  wire in_81bar, in_80bar, in_79bar, in_78bar, in_77bar, in_76bar, in_75bar, in_74bar, in_73bar, in_72bar, in_71bar, in_70bar, in_69bar, in_68bar, in_67bar, in_66bar, in_65bar, in_64bar, in_63bar, in_62bar, in_61bar, in_60bar, in_59bar, in_58bar, in_57bar, in_56bar, in_55bar, in_54bar, in_53bar, in_52bar, in_51bar, in_50bar, in_49bar, in_48bar, in_47bar, in_46bar, in_45bar, in_44bar, in_43bar, in_42bar, in_41bar, in_40bar, in_39bar, in_38bar, in_37bar, in_36bar, in_35bar, in_34bar, in_33bar, in_32bar, in_31bar, in_30bar, in_29bar, in_28bar, in_27bar, in_26bar, in_25bar, in_24bar, in_23bar, in_22bar, in_21bar, in_20bar, in_19bar, in_18bar, in_17bar, in_16bar, in_15bar, in_14bar, in_13bar, in_12bar, in_11bar, in_10bar, in_9bar, in_8bar, in_7bar, in_6bar, in_5bar, in_4bar, in_3bar, in_2bar, in_1bar, in_0bar, n487bar, n488bar, n489bar, n490bar, n491bar, n492bar, n493bar, n494bar, n495bar, n496bar, n497bar, n498bar, n499bar, n500bar, n501bar, n502bar, n503bar, n504bar, n505bar, n506bar, n507bar, n508bar, n509bar, n510bar, n511bar, n512bar, n513bar, n514bar, n515bar, n516bar, n517bar, n518bar, n519bar, n520bar, n521bar, n522bar, n523bar, n524bar, n525bar, n526bar, n527bar, n528bar, n529bar, n530bar, n531bar, n532bar, n533bar, n534bar, n535bar, n536bar, n537bar, n538bar, n539bar, n540bar, n541bar, n542bar, n543bar, n544bar, n545bar, n546bar, n547bar, n548bar, n549bar, n550bar, n551bar, n552bar, n553bar, n554bar, n555bar, n556bar, n557bar, n558bar, n559bar, n560bar, n561bar, n562bar, n563bar, n564bar, n565bar, n566bar, n567bar, n568bar, n569bar, n570bar, n571bar, n572bar, n573bar, n574bar, n575bar, n576bar, n577bar, n578bar, n579bar, n580bar, n581bar, n582bar, n583bar, n584bar, n585bar, n586bar, n587bar, n588bar, n589bar, n590bar, n591bar, n592bar, n593bar, n594bar, n595bar, n596bar, n597bar, n598bar, n599bar, n600bar, n601bar, n602bar, n603bar, n604bar, n605bar, n606bar, n607bar, n608bar, n609bar, n610bar, n611bar, n612bar, n613bar, n614bar, n615bar, n616bar, n617bar, n618bar, n619bar, n620bar, n621bar, n622bar, n623bar, n624bar, n625bar, n626bar, n627bar, n628bar, n629bar, n630bar, n631bar, n632bar, n633bar, n634bar, n635bar, n636bar, n637bar, n638bar, n639bar, n640bar, n641bar, n642bar, n643bar, n644bar, n645bar, n646bar, n647bar, n648bar, n649bar, n650bar, n651bar, n652bar, n653bar, n654bar, n655bar, n656bar, n657bar, n658bar, n659bar, n660bar, n661bar, n662bar, n663bar, n664bar, n665bar, n666bar, n667bar, n668bar, n669bar, n670bar, n671bar, n672bar, n673bar, n674bar, n675bar, n676bar, n677bar, n678bar, n679bar, n680bar, n681bar, n682bar, n683bar, n684bar, n685bar, n686bar, n687bar, n688bar, n689bar, n690bar, n691bar, n692bar, n693bar, n694bar, n695bar, n696bar, n697bar, n698bar, n699bar, n700bar, n701bar, n702bar, n703bar, n704bar, n705bar, n706bar, n707bar, n708bar, n709bar, n710bar, n711bar, n712bar, n713bar, n714bar, n715bar, n716bar, n717bar, n718bar, n719bar, n720bar, n721bar, n722bar, n723bar, n724bar, n725bar, n726bar, n727bar, n728bar, n729bar, n730bar, n731bar, n732bar, n733bar, n734bar, n735bar, n736bar, n737bar, n738bar, n739bar, n740bar, n741bar, n742bar, n743bar, n744bar, n745bar, n746bar, n747bar, n748bar, n749bar, n750bar, n751bar, n752bar, n753bar, n754bar, n755bar, n756bar, n757bar, n758bar, n759bar, n760bar, n761bar, n762bar, n763bar, n764bar, n765bar, n766bar, n767bar, n768bar, n769bar, n770bar, n771bar, n772bar, n773bar, n774bar, n775bar, n776bar, n777bar, n778bar, n779bar, n780bar, n781bar, n782bar, n783bar, n784bar, n785bar, n786bar, n787bar, n788bar, n789bar, n790bar, n791bar, n792bar, n793bar, n794bar, n795bar, n796bar, n797bar, n798bar, n799bar, n800bar, n801bar, n802bar, n803bar, n804bar, n805bar, n806bar, n807bar, n808bar, n809bar, n810bar, n811bar, n812bar, n813bar, n814bar, n815bar, n816bar, n817bar, n818bar, n819bar, n820bar, n821bar, n822bar, n823bar, n824bar, n825bar, n826bar, n827bar, n828bar, n829bar, n830bar, n831bar, n832bar, n833bar, n834bar, n835bar, n836bar, n837bar, n838bar, n839bar, n840bar, n841bar, n842bar, n843bar, n844bar, n845bar, n846bar, n847bar, n848bar, n849bar, n850bar, n851bar, n852bar, n853bar, n854bar, n855bar, n856bar, n857bar, n858bar, n859bar, n860bar, n861bar, n862bar, n863bar, n864bar, n865bar, n866bar, n867bar, n868bar, n869bar, n870bar, n871bar, n872bar, n873bar, n874bar, n875bar, n876bar, n877bar, n878bar, n879bar, n880bar, n881bar, n882bar, n883bar, n884bar, n885bar, n886bar, n887bar, n888bar, n889bar, n890bar, n891bar, n892bar, n893bar, n894bar, n895bar, n896bar, n897bar, n898bar, n899bar, n900bar, n901bar, n902bar, n903bar, n904bar, n905bar, n906bar, n907bar, n908bar, n909bar, n910bar, n911bar, n912bar, n913bar, n914bar, n915bar, n916bar, n917bar, n918bar, n919bar, n920bar, n921bar, n922bar, n923bar, n924bar, n925bar, n926bar, n927bar, n928bar, n929bar, n930bar, n931bar, n932bar, n933bar, n934bar, n935bar, n936bar, n937bar, n938bar, n939bar, n940bar, n941bar, n942bar, n943bar, n944bar, n945bar, n946bar, n947bar, n948bar, n949bar, n950bar, n951bar, n952bar, n953bar, n954bar, n955bar, n956bar, n957bar, n958bar, n959bar, n960bar, n961bar, n962bar, n963bar, n964bar, n965bar, n966bar, n967bar, n968bar, n969bar, n970bar, n971bar, n972bar;
  //wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];

  OR2_X1 U1 ( .A1(n972), .A2(n971), .ZN(out[7]) );
  AND2_X1 U1bar ( .A1(n972bar), .A2(n971bar), .ZN(outbar[7]);
  OR2_X1 U2 ( .A1(n970), .A2(n969), .ZN(n971) );
  AND2_X1 U2bar ( .A1(n970bar), .A2(n969bar), .ZN(n971bar);
  OR2_X1 U3 ( .A1(n968), .A2(n967), .ZN(n969) );
  AND2_X1 U3bar ( .A1(n968bar), .A2(n967bar), .ZN(n969bar);
  OR2_X1 U4 ( .A1(n966), .A2(n965), .ZN(n967) );
  AND2_X1 U4bar ( .A1(n966bar), .A2(n965bar), .ZN(n967bar);
  OR2_X1 U5 ( .A1(n964), .A2(n963), .ZN(n968) );
  AND2_X1 U5bar ( .A1(n964bar), .A2(n963bar), .ZN(n968bar);
  OR2_X1 U6 ( .A1(in[116]), .A2(n962), .ZN(n963) );
  AND2_X1 U6bar ( .A1(inbar[116]), .A2(n962bar), .ZN(n963bar);
  OR2_X1 U7 ( .A1(n961), .A2(n960), .ZN(n970) );
  AND2_X1 U7bar ( .A1(n961bar), .A2(n960bar), .ZN(n970bar);
  OR2_X1 U8 ( .A1(in[150]), .A2(in[127]), .ZN(n960) );
  AND2_X1 U8bar ( .A1(inbar[150]), .A2(inbar[127]), .ZN(n960bar);
  OR2_X1 U9 ( .A1(in[160]), .A2(n959), .ZN(n961) );
  AND2_X1 U9bar ( .A1(inbar[160]), .A2(n959bar), .ZN(n961bar);
  OR2_X1 U10 ( .A1(in[252]), .A2(in[168]), .ZN(n959) );
  AND2_X1 U10bar ( .A1(inbar[252]), .A2(inbar[168]), .ZN(n959bar);
  OR2_X1 U11 ( .A1(n958), .A2(n957), .ZN(n972) );
  AND2_X1 U11bar ( .A1(n958bar), .A2(n957bar), .ZN(n972bar);
  OR2_X1 U12 ( .A1(n956), .A2(n955), .ZN(n957) );
  AND2_X1 U12bar ( .A1(n956bar), .A2(n955bar), .ZN(n957bar);
  OR2_X1 U13 ( .A1(in_17), .A2(in[96]), .ZN(n955) );
  AND2_X1 U13bar ( .A1(in_17bar), .A2(inbar[96]), .ZN(n955bar);
  OR2_X1 U14 ( .A1(in_23), .A2(n954), .ZN(n956) );
  AND2_X1 U14bar ( .A1(in_23bar), .A2(n954bar), .ZN(n956bar);
  OR2_X1 U15 ( .A1(in_31), .A2(in_26), .ZN(n954) );
  AND2_X1 U15bar ( .A1(in_31bar), .A2(in_26bar), .ZN(n954bar);
  OR2_X1 U16 ( .A1(n953), .A2(n952), .ZN(n958) );
  AND2_X1 U16bar ( .A1(n953bar), .A2(n952bar), .ZN(n958bar);
  OR2_X1 U17 ( .A1(in_58), .A2(in_4), .ZN(n952) );
  AND2_X1 U17bar ( .A1(in_58bar), .A2(in_4bar), .ZN(n952bar);
  OR2_X1 U18 ( .A1(in_59), .A2(n951), .ZN(n953) );
  AND2_X1 U18bar ( .A1(in_59bar), .A2(n951bar), .ZN(n953bar);
  OR2_X1 U19 ( .A1(in_71), .A2(in_62), .ZN(n951) );
  AND2_X1 U19bar ( .A1(in_71bar), .A2(in_62bar), .ZN(n951bar);
  OR2_X1 U20 ( .A1(n950), .A2(n949), .ZN(out[6]) );
  AND2_X1 U20bar ( .A1(n950bar), .A2(n949bar), .ZN(outbar[6]);
  OR2_X1 U21 ( .A1(n948), .A2(n947), .ZN(n949) );
  AND2_X1 U21bar ( .A1(n948bar), .A2(n947bar), .ZN(n949bar);
  OR2_X1 U22 ( .A1(n946), .A2(n945), .ZN(n947) );
  AND2_X1 U22bar ( .A1(n946bar), .A2(n945bar), .ZN(n947bar);
  OR2_X1 U23 ( .A1(n944), .A2(n943), .ZN(n945) );
  AND2_X1 U23bar ( .A1(n944bar), .A2(n943bar), .ZN(n945bar);
  OR2_X1 U24 ( .A1(n942), .A2(n941), .ZN(n946) );
  AND2_X1 U24bar ( .A1(n942bar), .A2(n941bar), .ZN(n946bar);
  OR2_X1 U25 ( .A1(in[101]), .A2(n940), .ZN(n941) );
  AND2_X1 U25bar ( .A1(inbar[101]), .A2(n940bar), .ZN(n941bar);
  OR2_X1 U26 ( .A1(n939), .A2(n938), .ZN(n948) );
  AND2_X1 U26bar ( .A1(n939bar), .A2(n938bar), .ZN(n948bar);
  OR2_X1 U27 ( .A1(in[114]), .A2(in[104]), .ZN(n938) );
  AND2_X1 U27bar ( .A1(inbar[114]), .A2(inbar[104]), .ZN(n938bar);
  OR2_X1 U28 ( .A1(in[128]), .A2(n937), .ZN(n939) );
  AND2_X1 U28bar ( .A1(inbar[128]), .A2(n937bar), .ZN(n939bar);
  OR2_X1 U29 ( .A1(in[136]), .A2(in[134]), .ZN(n937) );
  AND2_X1 U29bar ( .A1(inbar[136]), .A2(inbar[134]), .ZN(n937bar);
  OR2_X1 U30 ( .A1(n936), .A2(n935), .ZN(n950) );
  AND2_X1 U30bar ( .A1(n936bar), .A2(n935bar), .ZN(n950bar);
  OR2_X1 U31 ( .A1(n934), .A2(n933), .ZN(n935) );
  AND2_X1 U31bar ( .A1(n934bar), .A2(n933bar), .ZN(n935bar);
  OR2_X1 U32 ( .A1(in[177]), .A2(in[164]), .ZN(n933) );
  AND2_X1 U32bar ( .A1(inbar[177]), .A2(inbar[164]), .ZN(n933bar);
  OR2_X1 U33 ( .A1(in[212]), .A2(n932), .ZN(n934) );
  AND2_X1 U33bar ( .A1(inbar[212]), .A2(n932bar), .ZN(n934bar);
  OR2_X1 U34 ( .A1(in[248]), .A2(in[221]), .ZN(n932) );
  AND2_X1 U34bar ( .A1(inbar[248]), .A2(inbar[221]), .ZN(n932bar);
  OR2_X1 U35 ( .A1(n931), .A2(n930), .ZN(n936) );
  AND2_X1 U35bar ( .A1(n931bar), .A2(n930bar), .ZN(n936bar);
  OR2_X1 U36 ( .A1(in_18), .A2(in[93]), .ZN(n930) );
  AND2_X1 U36bar ( .A1(in_18bar), .A2(inbar[93]), .ZN(n930bar);
  OR2_X1 U37 ( .A1(in_31), .A2(n929), .ZN(n931) );
  AND2_X1 U37bar ( .A1(in_31bar), .A2(n929bar), .ZN(n931bar);
  OR2_X1 U38 ( .A1(in_7), .A2(in_39), .ZN(n929) );
  AND2_X1 U38bar ( .A1(in_7bar), .A2(in_39bar), .ZN(n929bar);
  OR2_X1 U39 ( .A1(n928), .A2(n927), .ZN(out[5]) );
  AND2_X1 U39bar ( .A1(n928bar), .A2(n927bar), .ZN(outbar[5]);
  OR2_X1 U40 ( .A1(n926), .A2(n925), .ZN(n927) );
  AND2_X1 U40bar ( .A1(n926bar), .A2(n925bar), .ZN(n927bar);
  OR2_X1 U41 ( .A1(n924), .A2(n923), .ZN(n925) );
  AND2_X1 U41bar ( .A1(n924bar), .A2(n923bar), .ZN(n925bar);
  OR2_X1 U42 ( .A1(n922), .A2(n921), .ZN(n923) );
  AND2_X1 U42bar ( .A1(n922bar), .A2(n921bar), .ZN(n923bar);
  OR2_X1 U43 ( .A1(n940), .A2(n920), .ZN(n924) );
  AND2_X1 U43bar ( .A1(n940bar), .A2(n920bar), .ZN(n924bar);
  OR2_X1 U44 ( .A1(in[111]), .A2(n919), .ZN(n920) );
  AND2_X1 U44bar ( .A1(inbar[111]), .A2(n919bar), .ZN(n920bar);
  OR2_X1 U45 ( .A1(n918), .A2(n917), .ZN(n940) );
  AND2_X1 U45bar ( .A1(n918bar), .A2(n917bar), .ZN(n940bar);
  OR2_X1 U46 ( .A1(n916), .A2(n915), .ZN(n917) );
  AND2_X1 U46bar ( .A1(n916bar), .A2(n915bar), .ZN(n917bar);
  OR2_X1 U47 ( .A1(n914), .A2(n913), .ZN(n915) );
  AND2_X1 U47bar ( .A1(n914bar), .A2(n913bar), .ZN(n915bar);
  OR2_X1 U48 ( .A1(in[140]), .A2(in[131]), .ZN(n913) );
  AND2_X1 U48bar ( .A1(inbar[140]), .A2(inbar[131]), .ZN(n913bar);
  OR2_X1 U49 ( .A1(in[160]), .A2(in[144]), .ZN(n914) );
  AND2_X1 U49bar ( .A1(inbar[160]), .A2(inbar[144]), .ZN(n914bar);
  OR2_X1 U50 ( .A1(n912), .A2(n911), .ZN(n916) );
  AND2_X1 U50bar ( .A1(n912bar), .A2(n911bar), .ZN(n916bar);
  OR2_X1 U51 ( .A1(in[179]), .A2(in[174]), .ZN(n911) );
  AND2_X1 U51bar ( .A1(inbar[179]), .A2(inbar[174]), .ZN(n911bar);
  OR2_X1 U52 ( .A1(in[188]), .A2(in[184]), .ZN(n912) );
  AND2_X1 U52bar ( .A1(inbar[188]), .A2(inbar[184]), .ZN(n912bar);
  OR2_X1 U53 ( .A1(n910), .A2(n909), .ZN(n918) );
  AND2_X1 U53bar ( .A1(n910bar), .A2(n909bar), .ZN(n918bar);
  OR2_X1 U54 ( .A1(n908), .A2(n907), .ZN(n909) );
  AND2_X1 U54bar ( .A1(n908bar), .A2(n907bar), .ZN(n909bar);
  OR2_X1 U55 ( .A1(in[216]), .A2(in[200]), .ZN(n907) );
  AND2_X1 U55bar ( .A1(inbar[216]), .A2(inbar[200]), .ZN(n907bar);
  OR2_X1 U56 ( .A1(in[228]), .A2(in[224]), .ZN(n908) );
  AND2_X1 U56bar ( .A1(inbar[228]), .A2(inbar[224]), .ZN(n908bar);
  OR2_X1 U57 ( .A1(n906), .A2(n905), .ZN(n910) );
  AND2_X1 U57bar ( .A1(n906bar), .A2(n905bar), .ZN(n910bar);
  OR2_X1 U58 ( .A1(in[247]), .A2(in[235]), .ZN(n905) );
  AND2_X1 U58bar ( .A1(inbar[247]), .A2(inbar[235]), .ZN(n905bar);
  OR2_X1 U59 ( .A1(in_42), .A2(in[83]), .ZN(n906) );
  AND2_X1 U59bar ( .A1(in_42bar), .A2(inbar[83]), .ZN(n906bar);
  OR2_X1 U60 ( .A1(n904), .A2(n903), .ZN(n926) );
  AND2_X1 U60bar ( .A1(n904bar), .A2(n903bar), .ZN(n926bar);
  OR2_X1 U61 ( .A1(in[166]), .A2(in[123]), .ZN(n903) );
  AND2_X1 U61bar ( .A1(inbar[166]), .A2(inbar[123]), .ZN(n903bar);
  OR2_X1 U62 ( .A1(in[170]), .A2(n902), .ZN(n904) );
  AND2_X1 U62bar ( .A1(inbar[170]), .A2(n902bar), .ZN(n904bar);
  OR2_X1 U63 ( .A1(in[194]), .A2(in[183]), .ZN(n902) );
  AND2_X1 U63bar ( .A1(inbar[194]), .A2(inbar[183]), .ZN(n902bar);
  OR2_X1 U64 ( .A1(n901), .A2(n900), .ZN(n928) );
  AND2_X1 U64bar ( .A1(n901bar), .A2(n900bar), .ZN(n928bar);
  OR2_X1 U65 ( .A1(n899), .A2(n898), .ZN(n900) );
  AND2_X1 U65bar ( .A1(n899bar), .A2(n898bar), .ZN(n900bar);
  OR2_X1 U66 ( .A1(in[241]), .A2(in[238]), .ZN(n898) );
  AND2_X1 U66bar ( .A1(inbar[241]), .A2(inbar[238]), .ZN(n898bar);
  OR2_X1 U67 ( .A1(in[250]), .A2(n897), .ZN(n899) );
  AND2_X1 U67bar ( .A1(inbar[250]), .A2(n897bar), .ZN(n899bar);
  OR2_X1 U68 ( .A1(in_24), .A2(in[84]), .ZN(n897) );
  AND2_X1 U68bar ( .A1(in_24bar), .A2(inbar[84]), .ZN(n897bar);
  OR2_X1 U69 ( .A1(n896), .A2(n895), .ZN(n901) );
  AND2_X1 U69bar ( .A1(n896bar), .A2(n895bar), .ZN(n901bar);
  OR2_X1 U70 ( .A1(in_41), .A2(in_29), .ZN(n895) );
  AND2_X1 U70bar ( .A1(in_41bar), .A2(in_29bar), .ZN(n895bar);
  OR2_X1 U71 ( .A1(in_66), .A2(n894), .ZN(n896) );
  AND2_X1 U71bar ( .A1(in_66bar), .A2(n894bar), .ZN(n896bar);
  OR2_X1 U72 ( .A1(in_76), .A2(in_71), .ZN(n894) );
  AND2_X1 U72bar ( .A1(in_76bar), .A2(in_71bar), .ZN(n894bar);
  OR2_X1 U73 ( .A1(n893), .A2(n892), .ZN(out[4]) );
  AND2_X1 U73bar ( .A1(n893bar), .A2(n892bar), .ZN(outbar[4]);
  OR2_X1 U74 ( .A1(n891), .A2(n890), .ZN(n892) );
  AND2_X1 U74bar ( .A1(n891bar), .A2(n890bar), .ZN(n892bar);
  OR2_X1 U75 ( .A1(n889), .A2(n888), .ZN(n890) );
  AND2_X1 U75bar ( .A1(n889bar), .A2(n888bar), .ZN(n890bar);
  OR2_X1 U76 ( .A1(n922), .A2(n887), .ZN(n888) );
  AND2_X1 U76bar ( .A1(n922bar), .A2(n887bar), .ZN(n888bar);
  OR2_X1 U77 ( .A1(n886), .A2(n885), .ZN(n922) );
  AND2_X1 U77bar ( .A1(n886bar), .A2(n885bar), .ZN(n922bar);
  OR2_X1 U78 ( .A1(n884), .A2(n883), .ZN(n885) );
  AND2_X1 U78bar ( .A1(n884bar), .A2(n883bar), .ZN(n885bar);
  OR2_X1 U79 ( .A1(n882), .A2(n881), .ZN(n883) );
  AND2_X1 U79bar ( .A1(n882bar), .A2(n881bar), .ZN(n883bar);
  OR2_X1 U80 ( .A1(in[118]), .A2(in[109]), .ZN(n881) );
  AND2_X1 U80bar ( .A1(inbar[118]), .A2(inbar[109]), .ZN(n881bar);
  OR2_X1 U81 ( .A1(in[139]), .A2(in[120]), .ZN(n882) );
  AND2_X1 U81bar ( .A1(inbar[139]), .A2(inbar[120]), .ZN(n882bar);
  OR2_X1 U82 ( .A1(n880), .A2(n879), .ZN(n884) );
  AND2_X1 U82bar ( .A1(n880bar), .A2(n879bar), .ZN(n884bar);
  OR2_X1 U83 ( .A1(in[198]), .A2(in[154]), .ZN(n879) );
  AND2_X1 U83bar ( .A1(inbar[198]), .A2(inbar[154]), .ZN(n879bar);
  OR2_X1 U84 ( .A1(in[210]), .A2(in[205]), .ZN(n880) );
  AND2_X1 U84bar ( .A1(inbar[210]), .A2(inbar[205]), .ZN(n880bar);
  OR2_X1 U85 ( .A1(n878), .A2(n877), .ZN(n886) );
  AND2_X1 U85bar ( .A1(n878bar), .A2(n877bar), .ZN(n886bar);
  OR2_X1 U86 ( .A1(n876), .A2(n875), .ZN(n877) );
  AND2_X1 U86bar ( .A1(n876bar), .A2(n875bar), .ZN(n877bar);
  OR2_X1 U87 ( .A1(in[219]), .A2(in[217]), .ZN(n875) );
  AND2_X1 U87bar ( .A1(inbar[219]), .A2(inbar[217]), .ZN(n875bar);
  OR2_X1 U88 ( .A1(in[86]), .A2(in[252]), .ZN(n876) );
  AND2_X1 U88bar ( .A1(inbar[86]), .A2(inbar[252]), .ZN(n876bar);
  OR2_X1 U89 ( .A1(n874), .A2(n873), .ZN(n878) );
  AND2_X1 U89bar ( .A1(n874bar), .A2(n873bar), .ZN(n878bar);
  OR2_X1 U90 ( .A1(in_40), .A2(in[91]), .ZN(n873) );
  AND2_X1 U90bar ( .A1(in_40bar), .A2(inbar[91]), .ZN(n873bar);
  OR2_X1 U91 ( .A1(in_8), .A2(in_46), .ZN(n874) );
  AND2_X1 U91bar ( .A1(in_8bar), .A2(in_46bar), .ZN(n874bar);
  OR2_X1 U92 ( .A1(n872), .A2(n871), .ZN(n889) );
  AND2_X1 U92bar ( .A1(n872bar), .A2(n871bar), .ZN(n889bar);
  OR2_X1 U93 ( .A1(in[117]), .A2(n943), .ZN(n871) );
  AND2_X1 U93bar ( .A1(inbar[117]), .A2(n943bar), .ZN(n871bar);
  OR2_X1 U94 ( .A1(n870), .A2(n869), .ZN(n943) );
  AND2_X1 U94bar ( .A1(n870bar), .A2(n869bar), .ZN(n943bar);
  OR2_X1 U95 ( .A1(n868), .A2(n867), .ZN(n869) );
  AND2_X1 U95bar ( .A1(n868bar), .A2(n867bar), .ZN(n869bar);
  OR2_X1 U96 ( .A1(n866), .A2(n865), .ZN(n867) );
  AND2_X1 U96bar ( .A1(n866bar), .A2(n865bar), .ZN(n867bar);
  OR2_X1 U97 ( .A1(n864), .A2(n863), .ZN(n865) );
  AND2_X1 U97bar ( .A1(n864bar), .A2(n863bar), .ZN(n865bar);
  OR2_X1 U98 ( .A1(in[108]), .A2(n919), .ZN(n866) );
  AND2_X1 U98bar ( .A1(inbar[108]), .A2(n919bar), .ZN(n866bar);
  OR2_X1 U99 ( .A1(n862), .A2(n861), .ZN(n919) );
  AND2_X1 U99bar ( .A1(n862bar), .A2(n861bar), .ZN(n919bar);
  OR2_X1 U100 ( .A1(n860), .A2(n859), .ZN(n861) );
  AND2_X1 U100bar ( .A1(n860bar), .A2(n859bar), .ZN(n861bar);
  OR2_X1 U101 ( .A1(n858), .A2(n857), .ZN(n859) );
  AND2_X1 U101bar ( .A1(n858bar), .A2(n857bar), .ZN(n859bar);
  OR2_X1 U102 ( .A1(in[119]), .A2(in[105]), .ZN(n857) );
  AND2_X1 U102bar ( .A1(inbar[119]), .A2(inbar[105]), .ZN(n857bar);
  OR2_X1 U103 ( .A1(in[186]), .A2(in[175]), .ZN(n858) );
  AND2_X1 U103bar ( .A1(inbar[186]), .A2(inbar[175]), .ZN(n858bar);
  OR2_X1 U104 ( .A1(n856), .A2(n855), .ZN(n860) );
  AND2_X1 U104bar ( .A1(n856bar), .A2(n855bar), .ZN(n860bar);
  OR2_X1 U105 ( .A1(in[202]), .A2(in[193]), .ZN(n855) );
  AND2_X1 U105bar ( .A1(inbar[202]), .A2(inbar[193]), .ZN(n855bar);
  OR2_X1 U106 ( .A1(in[225]), .A2(in[208]), .ZN(n856) );
  AND2_X1 U106bar ( .A1(inbar[225]), .A2(inbar[208]), .ZN(n856bar);
  OR2_X1 U107 ( .A1(n854), .A2(n853), .ZN(n862) );
  AND2_X1 U107bar ( .A1(n854bar), .A2(n853bar), .ZN(n862bar);
  OR2_X1 U108 ( .A1(n852), .A2(n851), .ZN(n853) );
  AND2_X1 U108bar ( .A1(n852bar), .A2(n851bar), .ZN(n853bar);
  OR2_X1 U109 ( .A1(in_1), .A2(in[85]), .ZN(n851) );
  AND2_X1 U109bar ( .A1(in_1bar), .A2(inbar[85]), .ZN(n851bar);
  OR2_X1 U110 ( .A1(in_23), .A2(in_19), .ZN(n852) );
  AND2_X1 U110bar ( .A1(in_23bar), .A2(in_19bar), .ZN(n852bar);
  OR2_X1 U111 ( .A1(n850), .A2(n849), .ZN(n854) );
  AND2_X1 U111bar ( .A1(n850bar), .A2(n849bar), .ZN(n854bar);
  OR2_X1 U112 ( .A1(in_43), .A2(in_33), .ZN(n849) );
  AND2_X1 U112bar ( .A1(in_43bar), .A2(in_33bar), .ZN(n849bar);
  OR2_X1 U113 ( .A1(in_63), .A2(in_44), .ZN(n850) );
  AND2_X1 U113bar ( .A1(in_63bar), .A2(in_44bar), .ZN(n850bar);
  OR2_X1 U114 ( .A1(n848), .A2(n847), .ZN(n868) );
  AND2_X1 U114bar ( .A1(n848bar), .A2(n847bar), .ZN(n868bar);
  OR2_X1 U115 ( .A1(in[141]), .A2(in[112]), .ZN(n847) );
  AND2_X1 U115bar ( .A1(inbar[141]), .A2(inbar[112]), .ZN(n847bar);
  OR2_X1 U116 ( .A1(in[147]), .A2(n846), .ZN(n848) );
  AND2_X1 U116bar ( .A1(inbar[147]), .A2(n846bar), .ZN(n848bar);
  OR2_X1 U117 ( .A1(in[181]), .A2(in[167]), .ZN(n846) );
  AND2_X1 U117bar ( .A1(inbar[181]), .A2(inbar[167]), .ZN(n846bar);
  OR2_X1 U118 ( .A1(n845), .A2(n844), .ZN(n870) );
  AND2_X1 U118bar ( .A1(n845bar), .A2(n844bar), .ZN(n870bar);
  OR2_X1 U119 ( .A1(n843), .A2(n842), .ZN(n844) );
  AND2_X1 U119bar ( .A1(n843bar), .A2(n842bar), .ZN(n844bar);
  OR2_X1 U120 ( .A1(in[229]), .A2(in[201]), .ZN(n842) );
  AND2_X1 U120bar ( .A1(inbar[229]), .A2(inbar[201]), .ZN(n842bar);
  OR2_X1 U121 ( .A1(in[237]), .A2(n841), .ZN(n843) );
  AND2_X1 U121bar ( .A1(inbar[237]), .A2(n841bar), .ZN(n843bar);
  OR2_X1 U122 ( .A1(in[94]), .A2(in[253]), .ZN(n841) );
  AND2_X1 U122bar ( .A1(inbar[94]), .A2(inbar[253]), .ZN(n841bar);
  OR2_X1 U123 ( .A1(n840), .A2(n839), .ZN(n845) );
  AND2_X1 U123bar ( .A1(n840bar), .A2(n839bar), .ZN(n845bar);
  OR2_X1 U124 ( .A1(in_21), .A2(in[96]), .ZN(n839) );
  AND2_X1 U124bar ( .A1(in_21bar), .A2(inbar[96]), .ZN(n839bar);
  OR2_X1 U125 ( .A1(in_25), .A2(n838), .ZN(n840) );
  AND2_X1 U125bar ( .A1(in_25bar), .A2(n838bar), .ZN(n840bar);
  OR2_X1 U126 ( .A1(in_81), .A2(in_45), .ZN(n838) );
  AND2_X1 U126bar ( .A1(in_81bar), .A2(in_45bar), .ZN(n838bar);
  OR2_X1 U127 ( .A1(n837), .A2(n836), .ZN(n891) );
  AND2_X1 U127bar ( .A1(n837bar), .A2(n836bar), .ZN(n891bar);
  OR2_X1 U128 ( .A1(in[142]), .A2(in[124]), .ZN(n836) );
  AND2_X1 U128bar ( .A1(inbar[142]), .A2(inbar[124]), .ZN(n836bar);
  OR2_X1 U129 ( .A1(in[150]), .A2(n835), .ZN(n837) );
  AND2_X1 U129bar ( .A1(inbar[150]), .A2(n835bar), .ZN(n837bar);
  OR2_X1 U130 ( .A1(in[172]), .A2(in[155]), .ZN(n835) );
  AND2_X1 U130bar ( .A1(inbar[172]), .A2(inbar[155]), .ZN(n835bar);
  OR2_X1 U131 ( .A1(n834), .A2(n833), .ZN(n893) );
  AND2_X1 U131bar ( .A1(n834bar), .A2(n833bar), .ZN(n893bar);
  OR2_X1 U132 ( .A1(n832), .A2(n831), .ZN(n833) );
  AND2_X1 U132bar ( .A1(n832bar), .A2(n831bar), .ZN(n833bar);
  OR2_X1 U133 ( .A1(in[196]), .A2(in[173]), .ZN(n831) );
  AND2_X1 U133bar ( .A1(inbar[196]), .A2(inbar[173]), .ZN(n831bar);
  OR2_X1 U134 ( .A1(in[222]), .A2(n830), .ZN(n832) );
  AND2_X1 U134bar ( .A1(inbar[222]), .A2(n830bar), .ZN(n832bar);
  OR2_X1 U135 ( .A1(in[227]), .A2(in[226]), .ZN(n830) );
  AND2_X1 U135bar ( .A1(inbar[227]), .A2(inbar[226]), .ZN(n830bar);
  OR2_X1 U136 ( .A1(n829), .A2(n828), .ZN(n834) );
  AND2_X1 U136bar ( .A1(n829bar), .A2(n828bar), .ZN(n834bar);
  OR2_X1 U137 ( .A1(in[249]), .A2(in[231]), .ZN(n828) );
  AND2_X1 U137bar ( .A1(inbar[249]), .A2(inbar[231]), .ZN(n828bar);
  OR2_X1 U138 ( .A1(in_28), .A2(n827), .ZN(n829) );
  AND2_X1 U138bar ( .A1(in_28bar), .A2(n827bar), .ZN(n829bar);
  OR2_X1 U139 ( .A1(in_52), .A2(in_47), .ZN(n827) );
  AND2_X1 U139bar ( .A1(in_52bar), .A2(in_47bar), .ZN(n827bar);
  OR2_X1 U140 ( .A1(n826), .A2(n825), .ZN(out[3]) );
  AND2_X1 U140bar ( .A1(n826bar), .A2(n825bar), .ZN(outbar[3]);
  OR2_X1 U141 ( .A1(n824), .A2(n823), .ZN(n825) );
  AND2_X1 U141bar ( .A1(n824bar), .A2(n823bar), .ZN(n825bar);
  OR2_X1 U142 ( .A1(n822), .A2(n821), .ZN(n823) );
  AND2_X1 U142bar ( .A1(n822bar), .A2(n821bar), .ZN(n823bar);
  OR2_X1 U143 ( .A1(n820), .A2(n819), .ZN(n821) );
  AND2_X1 U143bar ( .A1(n820bar), .A2(n819bar), .ZN(n821bar);
  OR2_X1 U144 ( .A1(n964), .A2(n818), .ZN(n822) );
  AND2_X1 U144bar ( .A1(n964bar), .A2(n818bar), .ZN(n822bar);
  OR2_X1 U145 ( .A1(in[118]), .A2(n817), .ZN(n818) );
  AND2_X1 U145bar ( .A1(inbar[118]), .A2(n817bar), .ZN(n818bar);
  OR2_X1 U146 ( .A1(n816), .A2(n815), .ZN(n964) );
  AND2_X1 U146bar ( .A1(n816bar), .A2(n815bar), .ZN(n964bar);
  OR2_X1 U147 ( .A1(n814), .A2(n813), .ZN(n815) );
  AND2_X1 U147bar ( .A1(n814bar), .A2(n813bar), .ZN(n815bar);
  OR2_X1 U148 ( .A1(n812), .A2(n811), .ZN(n813) );
  AND2_X1 U148bar ( .A1(n812bar), .A2(n811bar), .ZN(n813bar);
  OR2_X1 U149 ( .A1(in[122]), .A2(in[111]), .ZN(n811) );
  AND2_X1 U149bar ( .A1(inbar[122]), .A2(inbar[111]), .ZN(n811bar);
  OR2_X1 U150 ( .A1(in[154]), .A2(in[151]), .ZN(n812) );
  AND2_X1 U150bar ( .A1(inbar[154]), .A2(inbar[151]), .ZN(n812bar);
  OR2_X1 U151 ( .A1(n810), .A2(n809), .ZN(n814) );
  AND2_X1 U151bar ( .A1(n810bar), .A2(n809bar), .ZN(n814bar);
  OR2_X1 U152 ( .A1(in[187]), .A2(in[177]), .ZN(n809) );
  AND2_X1 U152bar ( .A1(inbar[187]), .A2(inbar[177]), .ZN(n809bar);
  OR2_X1 U153 ( .A1(in[200]), .A2(in[192]), .ZN(n810) );
  AND2_X1 U153bar ( .A1(inbar[200]), .A2(inbar[192]), .ZN(n810bar);
  OR2_X1 U154 ( .A1(n808), .A2(n807), .ZN(n816) );
  AND2_X1 U154bar ( .A1(n808bar), .A2(n807bar), .ZN(n816bar);
  OR2_X1 U155 ( .A1(n806), .A2(n805), .ZN(n807) );
  AND2_X1 U155bar ( .A1(n806bar), .A2(n805bar), .ZN(n807bar);
  OR2_X1 U156 ( .A1(in[225]), .A2(in[207]), .ZN(n805) );
  AND2_X1 U156bar ( .A1(inbar[225]), .A2(inbar[207]), .ZN(n805bar);
  OR2_X1 U157 ( .A1(in[98]), .A2(in[226]), .ZN(n806) );
  AND2_X1 U157bar ( .A1(inbar[98]), .A2(inbar[226]), .ZN(n806bar);
  OR2_X1 U158 ( .A1(n804), .A2(n803), .ZN(n808) );
  AND2_X1 U158bar ( .A1(n804bar), .A2(n803bar), .ZN(n808bar);
  OR2_X1 U159 ( .A1(in_20), .A2(in_16), .ZN(n803) );
  AND2_X1 U159bar ( .A1(in_20bar), .A2(in_16bar), .ZN(n803bar);
  OR2_X1 U160 ( .A1(in_55), .A2(in_45), .ZN(n804) );
  AND2_X1 U160bar ( .A1(in_55bar), .A2(in_45bar), .ZN(n804bar);
  OR2_X1 U161 ( .A1(n802), .A2(n801), .ZN(n824) );
  AND2_X1 U161bar ( .A1(n802bar), .A2(n801bar), .ZN(n824bar);
  OR2_X1 U162 ( .A1(in[162]), .A2(in[149]), .ZN(n801) );
  AND2_X1 U162bar ( .A1(inbar[162]), .A2(inbar[149]), .ZN(n801bar);
  OR2_X1 U163 ( .A1(in[163]), .A2(n800), .ZN(n802) );
  AND2_X1 U163bar ( .A1(inbar[163]), .A2(n800bar), .ZN(n802bar);
  OR2_X1 U164 ( .A1(in[191]), .A2(in[189]), .ZN(n800) );
  AND2_X1 U164bar ( .A1(inbar[191]), .A2(inbar[189]), .ZN(n800bar);
  OR2_X1 U165 ( .A1(n799), .A2(n798), .ZN(n826) );
  AND2_X1 U165bar ( .A1(n799bar), .A2(n798bar), .ZN(n826bar);
  OR2_X1 U166 ( .A1(n797), .A2(n796), .ZN(n798) );
  AND2_X1 U166bar ( .A1(n797bar), .A2(n796bar), .ZN(n798bar);
  OR2_X1 U167 ( .A1(in[212]), .A2(in[193]), .ZN(n796) );
  AND2_X1 U167bar ( .A1(inbar[212]), .A2(inbar[193]), .ZN(n796bar);
  OR2_X1 U168 ( .A1(in[238]), .A2(n795), .ZN(n797) );
  AND2_X1 U168bar ( .A1(inbar[238]), .A2(n795bar), .ZN(n797bar);
  OR2_X1 U169 ( .A1(in[88]), .A2(in[247]), .ZN(n795) );
  AND2_X1 U169bar ( .A1(inbar[88]), .A2(inbar[247]), .ZN(n795bar);
  OR2_X1 U170 ( .A1(n794), .A2(n793), .ZN(n799) );
  AND2_X1 U170bar ( .A1(n794bar), .A2(n793bar), .ZN(n799bar);
  OR2_X1 U171 ( .A1(in[94]), .A2(in[92]), .ZN(n793) );
  AND2_X1 U171bar ( .A1(inbar[94]), .A2(inbar[92]), .ZN(n793bar);
  OR2_X1 U172 ( .A1(in_52), .A2(n792), .ZN(n794) );
  AND2_X1 U172bar ( .A1(in_52bar), .A2(n792bar), .ZN(n794bar);
  OR2_X1 U173 ( .A1(in_70), .A2(in_67), .ZN(n792) );
  AND2_X1 U173bar ( .A1(in_70bar), .A2(in_67bar), .ZN(n792bar);
  OR2_X1 U174 ( .A1(n791), .A2(n790), .ZN(out[2]) );
  AND2_X1 U174bar ( .A1(n791bar), .A2(n790bar), .ZN(outbar[2]);
  OR2_X1 U175 ( .A1(n789), .A2(n788), .ZN(n790) );
  AND2_X1 U175bar ( .A1(n789bar), .A2(n788bar), .ZN(n790bar);
  OR2_X1 U176 ( .A1(n787), .A2(n786), .ZN(n788) );
  AND2_X1 U176bar ( .A1(n787bar), .A2(n786bar), .ZN(n788bar);
  OR2_X1 U177 ( .A1(n819), .A2(n785), .ZN(n786) );
  AND2_X1 U177bar ( .A1(n819bar), .A2(n785bar), .ZN(n786bar);
  OR2_X1 U178 ( .A1(n784), .A2(n783), .ZN(n819) );
  AND2_X1 U178bar ( .A1(n784bar), .A2(n783bar), .ZN(n819bar);
  OR2_X1 U179 ( .A1(n782), .A2(n781), .ZN(n783) );
  AND2_X1 U179bar ( .A1(n782bar), .A2(n781bar), .ZN(n783bar);
  OR2_X1 U180 ( .A1(n780), .A2(n779), .ZN(n781) );
  AND2_X1 U180bar ( .A1(n780bar), .A2(n779bar), .ZN(n781bar);
  OR2_X1 U181 ( .A1(n962), .A2(n778), .ZN(n779) );
  AND2_X1 U181bar ( .A1(n962bar), .A2(n778bar), .ZN(n779bar);
  OR2_X1 U182 ( .A1(n777), .A2(n776), .ZN(n962) );
  AND2_X1 U182bar ( .A1(n777bar), .A2(n776bar), .ZN(n962bar);
  OR2_X1 U183 ( .A1(n775), .A2(n774), .ZN(n776) );
  AND2_X1 U183bar ( .A1(n775bar), .A2(n774bar), .ZN(n776bar);
  OR2_X1 U184 ( .A1(n773), .A2(n772), .ZN(n774) );
  AND2_X1 U184bar ( .A1(n773bar), .A2(n772bar), .ZN(n774bar);
  OR2_X1 U185 ( .A1(in[131]), .A2(in[120]), .ZN(n772) );
  AND2_X1 U185bar ( .A1(inbar[131]), .A2(inbar[120]), .ZN(n772bar);
  OR2_X1 U186 ( .A1(in[153]), .A2(in[147]), .ZN(n773) );
  AND2_X1 U186bar ( .A1(inbar[153]), .A2(inbar[147]), .ZN(n773bar);
  OR2_X1 U187 ( .A1(n771), .A2(n770), .ZN(n775) );
  AND2_X1 U187bar ( .A1(n771bar), .A2(n770bar), .ZN(n775bar);
  OR2_X1 U188 ( .A1(in[170]), .A2(in[156]), .ZN(n770) );
  AND2_X1 U188bar ( .A1(inbar[170]), .A2(inbar[156]), .ZN(n770bar);
  OR2_X1 U189 ( .A1(in[223]), .A2(in[190]), .ZN(n771) );
  AND2_X1 U189bar ( .A1(inbar[223]), .A2(inbar[190]), .ZN(n771bar);
  OR2_X1 U190 ( .A1(n769), .A2(n768), .ZN(n777) );
  AND2_X1 U190bar ( .A1(n769bar), .A2(n768bar), .ZN(n777bar);
  OR2_X1 U191 ( .A1(n767), .A2(n766), .ZN(n768) );
  AND2_X1 U191bar ( .A1(n767bar), .A2(n766bar), .ZN(n768bar);
  OR2_X1 U192 ( .A1(in[236]), .A2(in[230]), .ZN(n766) );
  AND2_X1 U192bar ( .A1(inbar[236]), .A2(inbar[230]), .ZN(n766bar);
  OR2_X1 U193 ( .A1(in[85]), .A2(in[240]), .ZN(n767) );
  AND2_X1 U193bar ( .A1(inbar[85]), .A2(inbar[240]), .ZN(n767bar);
  OR2_X1 U194 ( .A1(n765), .A2(n764), .ZN(n769) );
  AND2_X1 U194bar ( .A1(n765bar), .A2(n764bar), .ZN(n769bar);
  OR2_X1 U195 ( .A1(in_12), .A2(in[90]), .ZN(n764) );
  AND2_X1 U195bar ( .A1(in_12bar), .A2(inbar[90]), .ZN(n764bar);
  OR2_X1 U196 ( .A1(in_39), .A2(in_28), .ZN(n765) );
  AND2_X1 U196bar ( .A1(in_39bar), .A2(in_28bar), .ZN(n765bar);
  OR2_X1 U197 ( .A1(in[109]), .A2(n763), .ZN(n780) );
  AND2_X1 U197bar ( .A1(inbar[109]), .A2(n763bar), .ZN(n780bar);
  OR2_X1 U198 ( .A1(n762), .A2(n761), .ZN(n782) );
  AND2_X1 U198bar ( .A1(n762bar), .A2(n761bar), .ZN(n782bar);
  OR2_X1 U199 ( .A1(in[138]), .A2(in[129]), .ZN(n761) );
  AND2_X1 U199bar ( .A1(inbar[138]), .A2(inbar[129]), .ZN(n761bar);
  OR2_X1 U200 ( .A1(in[157]), .A2(n760), .ZN(n762) );
  AND2_X1 U200bar ( .A1(inbar[157]), .A2(n760bar), .ZN(n762bar);
  OR2_X1 U201 ( .A1(in[182]), .A2(in[167]), .ZN(n760) );
  AND2_X1 U201bar ( .A1(inbar[182]), .A2(inbar[167]), .ZN(n760bar);
  OR2_X1 U202 ( .A1(n759), .A2(n758), .ZN(n784) );
  AND2_X1 U202bar ( .A1(n759bar), .A2(n758bar), .ZN(n784bar);
  OR2_X1 U203 ( .A1(n757), .A2(n756), .ZN(n758) );
  AND2_X1 U203bar ( .A1(n757bar), .A2(n756bar), .ZN(n758bar);
  OR2_X1 U204 ( .A1(in[195]), .A2(in[184]), .ZN(n756) );
  AND2_X1 U204bar ( .A1(inbar[195]), .A2(inbar[184]), .ZN(n756bar);
  OR2_X1 U205 ( .A1(in[196]), .A2(n755), .ZN(n757) );
  AND2_X1 U205bar ( .A1(inbar[196]), .A2(n755bar), .ZN(n757bar);
  OR2_X1 U206 ( .A1(in[215]), .A2(in[209]), .ZN(n755) );
  AND2_X1 U206bar ( .A1(inbar[215]), .A2(inbar[209]), .ZN(n755bar);
  OR2_X1 U207 ( .A1(n754), .A2(n753), .ZN(n759) );
  AND2_X1 U207bar ( .A1(n754bar), .A2(n753bar), .ZN(n759bar);
  OR2_X1 U208 ( .A1(in[93]), .A2(in[233]), .ZN(n753) );
  AND2_X1 U208bar ( .A1(inbar[93]), .A2(inbar[233]), .ZN(n753bar);
  OR2_X1 U209 ( .A1(in_1), .A2(n752), .ZN(n754) );
  AND2_X1 U209bar ( .A1(in_1bar), .A2(n752bar), .ZN(n754bar);
  OR2_X1 U210 ( .A1(in_69), .A2(in_66), .ZN(n752) );
  AND2_X1 U210bar ( .A1(in_69bar), .A2(in_66bar), .ZN(n752bar);
  OR2_X1 U211 ( .A1(n966), .A2(n751), .ZN(n787) );
  AND2_X1 U211bar ( .A1(n966bar), .A2(n751bar), .ZN(n787bar);
  OR2_X1 U212 ( .A1(in[134]), .A2(n750), .ZN(n751) );
  AND2_X1 U212bar ( .A1(inbar[134]), .A2(n750bar), .ZN(n751bar);
  OR2_X1 U213 ( .A1(n749), .A2(n748), .ZN(n966) );
  AND2_X1 U213bar ( .A1(n749bar), .A2(n748bar), .ZN(n966bar);
  OR2_X1 U214 ( .A1(n747), .A2(n746), .ZN(n748) );
  AND2_X1 U214bar ( .A1(n747bar), .A2(n746bar), .ZN(n748bar);
  OR2_X1 U215 ( .A1(n745), .A2(n744), .ZN(n746) );
  AND2_X1 U215bar ( .A1(n745bar), .A2(n744bar), .ZN(n746bar);
  OR2_X1 U216 ( .A1(in[136]), .A2(in[121]), .ZN(n744) );
  AND2_X1 U216bar ( .A1(inbar[136]), .A2(inbar[121]), .ZN(n744bar);
  OR2_X1 U217 ( .A1(in[186]), .A2(in[174]), .ZN(n745) );
  AND2_X1 U217bar ( .A1(inbar[186]), .A2(inbar[174]), .ZN(n745bar);
  OR2_X1 U218 ( .A1(n743), .A2(n742), .ZN(n747) );
  AND2_X1 U218bar ( .A1(n743bar), .A2(n742bar), .ZN(n747bar);
  OR2_X1 U219 ( .A1(in[198]), .A2(in[197]), .ZN(n742) );
  AND2_X1 U219bar ( .A1(inbar[198]), .A2(inbar[197]), .ZN(n742bar);
  OR2_X1 U220 ( .A1(in[214]), .A2(in[199]), .ZN(n743) );
  AND2_X1 U220bar ( .A1(inbar[214]), .A2(inbar[199]), .ZN(n743bar);
  OR2_X1 U221 ( .A1(n741), .A2(n740), .ZN(n749) );
  AND2_X1 U221bar ( .A1(n741bar), .A2(n740bar), .ZN(n749bar);
  OR2_X1 U222 ( .A1(n739), .A2(n738), .ZN(n740) );
  AND2_X1 U222bar ( .A1(n739bar), .A2(n738bar), .ZN(n740bar);
  OR2_X1 U223 ( .A1(in[231]), .A2(in[220]), .ZN(n738) );
  AND2_X1 U223bar ( .A1(inbar[231]), .A2(inbar[220]), .ZN(n738bar);
  OR2_X1 U224 ( .A1(in_25), .A2(in[245]), .ZN(n739) );
  AND2_X1 U224bar ( .A1(in_25bar), .A2(inbar[245]), .ZN(n739bar);
  OR2_X1 U225 ( .A1(n737), .A2(n736), .ZN(n741) );
  AND2_X1 U225bar ( .A1(n737bar), .A2(n736bar), .ZN(n741bar);
  OR2_X1 U226 ( .A1(in_53), .A2(in_29), .ZN(n736) );
  AND2_X1 U226bar ( .A1(in_53bar), .A2(in_29bar), .ZN(n736bar);
  OR2_X1 U227 ( .A1(in_79), .A2(in_74), .ZN(n737) );
  AND2_X1 U227bar ( .A1(in_79bar), .A2(in_74bar), .ZN(n737bar);
  OR2_X1 U228 ( .A1(n735), .A2(n734), .ZN(n789) );
  AND2_X1 U228bar ( .A1(n735bar), .A2(n734bar), .ZN(n789bar);
  OR2_X1 U229 ( .A1(in[152]), .A2(in[140]), .ZN(n734) );
  AND2_X1 U229bar ( .A1(inbar[152]), .A2(inbar[140]), .ZN(n734bar);
  OR2_X1 U230 ( .A1(in[155]), .A2(n733), .ZN(n735) );
  AND2_X1 U230bar ( .A1(inbar[155]), .A2(n733bar), .ZN(n735bar);
  OR2_X1 U231 ( .A1(in[166]), .A2(in[165]), .ZN(n733) );
  AND2_X1 U231bar ( .A1(inbar[166]), .A2(inbar[165]), .ZN(n733bar);
  OR2_X1 U232 ( .A1(n732), .A2(n731), .ZN(n791) );
  AND2_X1 U232bar ( .A1(n732bar), .A2(n731bar), .ZN(n791bar);
  OR2_X1 U233 ( .A1(n730), .A2(n729), .ZN(n731) );
  AND2_X1 U233bar ( .A1(n730bar), .A2(n729bar), .ZN(n731bar);
  OR2_X1 U234 ( .A1(in[202]), .A2(in[185]), .ZN(n729) );
  AND2_X1 U234bar ( .A1(inbar[202]), .A2(inbar[185]), .ZN(n729bar);
  OR2_X1 U235 ( .A1(in[211]), .A2(n728), .ZN(n730) );
  AND2_X1 U235bar ( .A1(inbar[211]), .A2(n728bar), .ZN(n730bar);
  OR2_X1 U236 ( .A1(in[255]), .A2(in[253]), .ZN(n728) );
  AND2_X1 U236bar ( .A1(inbar[255]), .A2(inbar[253]), .ZN(n728bar);
  OR2_X1 U237 ( .A1(n727), .A2(n726), .ZN(n732) );
  AND2_X1 U237bar ( .A1(n727bar), .A2(n726bar), .ZN(n732bar);
  OR2_X1 U238 ( .A1(in_35), .A2(in_15), .ZN(n726) );
  AND2_X1 U238bar ( .A1(in_35bar), .A2(in_15bar), .ZN(n726bar);
  OR2_X1 U239 ( .A1(in_36), .A2(n725), .ZN(n727) );
  AND2_X1 U239bar ( .A1(in_36bar), .A2(n725bar), .ZN(n727bar);
  OR2_X1 U240 ( .A1(in_48), .A2(in_40), .ZN(n725) );
  AND2_X1 U240bar ( .A1(in_48bar), .A2(in_40bar), .ZN(n725bar);
  OR2_X1 U241 ( .A1(n724), .A2(n723), .ZN(out[1]) );
  AND2_X1 U241bar ( .A1(n724bar), .A2(n723bar), .ZN(outbar[1]);
  OR2_X1 U242 ( .A1(n722), .A2(n721), .ZN(n723) );
  AND2_X1 U242bar ( .A1(n722bar), .A2(n721bar), .ZN(n723bar);
  OR2_X1 U243 ( .A1(n720), .A2(n719), .ZN(n721) );
  AND2_X1 U243bar ( .A1(n720bar), .A2(n719bar), .ZN(n721bar);
  OR2_X1 U244 ( .A1(n921), .A2(n887), .ZN(n719) );
  AND2_X1 U244bar ( .A1(n921bar), .A2(n887bar), .ZN(n719bar);
  OR2_X1 U245 ( .A1(n718), .A2(n717), .ZN(n887) );
  AND2_X1 U245bar ( .A1(n718bar), .A2(n717bar), .ZN(n887bar);
  OR2_X1 U246 ( .A1(n716), .A2(n715), .ZN(n717) );
  AND2_X1 U246bar ( .A1(n716bar), .A2(n715bar), .ZN(n717bar);
  OR2_X1 U247 ( .A1(n714), .A2(n713), .ZN(n715) );
  AND2_X1 U247bar ( .A1(n714bar), .A2(n713bar), .ZN(n715bar);
  OR2_X1 U248 ( .A1(in[116]), .A2(in[110]), .ZN(n713) );
  AND2_X1 U248bar ( .A1(inbar[116]), .A2(inbar[110]), .ZN(n713bar);
  OR2_X1 U249 ( .A1(in[133]), .A2(in[130]), .ZN(n714) );
  AND2_X1 U249bar ( .A1(inbar[133]), .A2(inbar[130]), .ZN(n714bar);
  OR2_X1 U250 ( .A1(n712), .A2(n711), .ZN(n716) );
  AND2_X1 U250bar ( .A1(n712bar), .A2(n711bar), .ZN(n716bar);
  OR2_X1 U251 ( .A1(in[203]), .A2(in[135]), .ZN(n711) );
  AND2_X1 U251bar ( .A1(inbar[203]), .A2(inbar[135]), .ZN(n711bar);
  OR2_X1 U252 ( .A1(in[232]), .A2(in[223]), .ZN(n712) );
  AND2_X1 U252bar ( .A1(inbar[232]), .A2(inbar[223]), .ZN(n712bar);
  OR2_X1 U253 ( .A1(n710), .A2(n709), .ZN(n718) );
  AND2_X1 U253bar ( .A1(n710bar), .A2(n709bar), .ZN(n718bar);
  OR2_X1 U254 ( .A1(n708), .A2(n707), .ZN(n709) );
  AND2_X1 U254bar ( .A1(n708bar), .A2(n707bar), .ZN(n709bar);
  OR2_X1 U255 ( .A1(in[255]), .A2(in[233]), .ZN(n707) );
  AND2_X1 U255bar ( .A1(inbar[255]), .A2(inbar[233]), .ZN(n707bar);
  OR2_X1 U256 ( .A1(in_53), .A2(in_34), .ZN(n708) );
  AND2_X1 U256bar ( .A1(in_53bar), .A2(in_34bar), .ZN(n708bar);
  OR2_X1 U257 ( .A1(n706), .A2(n705), .ZN(n710) );
  AND2_X1 U257bar ( .A1(n706bar), .A2(n705bar), .ZN(n710bar);
  OR2_X1 U258 ( .A1(in_57), .A2(in_55), .ZN(n705) );
  AND2_X1 U258bar ( .A1(in_57bar), .A2(in_55bar), .ZN(n705bar);
  OR2_X1 U259 ( .A1(in_68), .A2(in_67), .ZN(n706) );
  AND2_X1 U259bar ( .A1(in_68bar), .A2(in_67bar), .ZN(n706bar);
  OR2_X1 U260 ( .A1(n704), .A2(n703), .ZN(n921) );
  AND2_X1 U260bar ( .A1(n704bar), .A2(n703bar), .ZN(n921bar);
  OR2_X1 U261 ( .A1(n702), .A2(n701), .ZN(n703) );
  AND2_X1 U261bar ( .A1(n702bar), .A2(n701bar), .ZN(n703bar);
  OR2_X1 U262 ( .A1(n700), .A2(n699), .ZN(n701) );
  AND2_X1 U262bar ( .A1(n700bar), .A2(n699bar), .ZN(n701bar);
  OR2_X1 U263 ( .A1(n944), .A2(n872), .ZN(n699) );
  AND2_X1 U263bar ( .A1(n944bar), .A2(n872bar), .ZN(n699bar);
  OR2_X1 U264 ( .A1(n698), .A2(n697), .ZN(n872) );
  AND2_X1 U264bar ( .A1(n698bar), .A2(n697bar), .ZN(n872bar);
  OR2_X1 U265 ( .A1(n696), .A2(n695), .ZN(n697) );
  AND2_X1 U265bar ( .A1(n696bar), .A2(n695bar), .ZN(n697bar);
  OR2_X1 U266 ( .A1(n694), .A2(n693), .ZN(n695) );
  AND2_X1 U266bar ( .A1(n694bar), .A2(n693bar), .ZN(n695bar);
  OR2_X1 U267 ( .A1(in[121]), .A2(in[102]), .ZN(n693) );
  AND2_X1 U267bar ( .A1(inbar[121]), .A2(inbar[102]), .ZN(n693bar);
  OR2_X1 U268 ( .A1(in[162]), .A2(in[161]), .ZN(n694) );
  AND2_X1 U268bar ( .A1(inbar[162]), .A2(inbar[161]), .ZN(n694bar);
  OR2_X1 U269 ( .A1(n692), .A2(n691), .ZN(n696) );
  AND2_X1 U269bar ( .A1(n692bar), .A2(n691bar), .ZN(n696bar);
  OR2_X1 U270 ( .A1(in[192]), .A2(in[178]), .ZN(n691) );
  AND2_X1 U270bar ( .A1(inbar[192]), .A2(inbar[178]), .ZN(n691bar);
  OR2_X1 U271 ( .A1(in[244]), .A2(in[209]), .ZN(n692) );
  AND2_X1 U271bar ( .A1(inbar[244]), .A2(inbar[209]), .ZN(n692bar);
  OR2_X1 U272 ( .A1(n690), .A2(n689), .ZN(n698) );
  AND2_X1 U272bar ( .A1(n690bar), .A2(n689bar), .ZN(n698bar);
  OR2_X1 U273 ( .A1(n688), .A2(n687), .ZN(n689) );
  AND2_X1 U273bar ( .A1(n688bar), .A2(n687bar), .ZN(n689bar);
  OR2_X1 U274 ( .A1(in[90]), .A2(in[254]), .ZN(n687) );
  AND2_X1 U274bar ( .A1(inbar[90]), .A2(inbar[254]), .ZN(n687bar);
  OR2_X1 U275 ( .A1(in_36), .A2(in_32), .ZN(n688) );
  AND2_X1 U275bar ( .A1(in_36bar), .A2(in_32bar), .ZN(n688bar);
  OR2_X1 U276 ( .A1(n686), .A2(n685), .ZN(n690) );
  AND2_X1 U276bar ( .A1(n686bar), .A2(n685bar), .ZN(n690bar);
  OR2_X1 U277 ( .A1(in_62), .A2(in_37), .ZN(n685) );
  AND2_X1 U277bar ( .A1(in_62bar), .A2(in_37bar), .ZN(n685bar);
  OR2_X1 U278 ( .A1(in_75), .A2(in_73), .ZN(n686) );
  AND2_X1 U278bar ( .A1(in_75bar), .A2(in_73bar), .ZN(n686bar);
  OR2_X1 U279 ( .A1(n684), .A2(n683), .ZN(n944) );
  AND2_X1 U279bar ( .A1(n684bar), .A2(n683bar), .ZN(n944bar);
  OR2_X1 U280 ( .A1(n682), .A2(n681), .ZN(n683) );
  AND2_X1 U280bar ( .A1(n682bar), .A2(n681bar), .ZN(n683bar);
  OR2_X1 U281 ( .A1(n680), .A2(n679), .ZN(n681) );
  AND2_X1 U281bar ( .A1(n680bar), .A2(n679bar), .ZN(n681bar);
  OR2_X1 U282 ( .A1(in[171]), .A2(in[153]), .ZN(n679) );
  AND2_X1 U282bar ( .A1(inbar[171]), .A2(inbar[153]), .ZN(n679bar);
  OR2_X1 U283 ( .A1(in[187]), .A2(in[176]), .ZN(n680) );
  AND2_X1 U283bar ( .A1(inbar[187]), .A2(inbar[176]), .ZN(n680bar);
  OR2_X1 U284 ( .A1(n678), .A2(n677), .ZN(n682) );
  AND2_X1 U284bar ( .A1(n678bar), .A2(n677bar), .ZN(n682bar);
  OR2_X1 U285 ( .A1(in[245]), .A2(in[211]), .ZN(n677) );
  AND2_X1 U285bar ( .A1(inbar[245]), .A2(inbar[211]), .ZN(n677bar);
  OR2_X1 U286 ( .A1(in[97]), .A2(in[88]), .ZN(n678) );
  AND2_X1 U286bar ( .A1(inbar[97]), .A2(inbar[88]), .ZN(n678bar);
  OR2_X1 U287 ( .A1(n676), .A2(n675), .ZN(n684) );
  AND2_X1 U287bar ( .A1(n676bar), .A2(n675bar), .ZN(n684bar);
  OR2_X1 U288 ( .A1(n674), .A2(n673), .ZN(n675) );
  AND2_X1 U288bar ( .A1(n674bar), .A2(n673bar), .ZN(n675bar);
  OR2_X1 U289 ( .A1(in_10), .A2(in_0), .ZN(n673) );
  AND2_X1 U289bar ( .A1(in_10bar), .A2(in_0bar), .ZN(n673bar);
  OR2_X1 U290 ( .A1(in_59), .A2(in_5), .ZN(n674) );
  AND2_X1 U290bar ( .A1(in_59bar), .A2(in_5bar), .ZN(n674bar);
  OR2_X1 U291 ( .A1(n672), .A2(n671), .ZN(n676) );
  AND2_X1 U291bar ( .A1(n672bar), .A2(n671bar), .ZN(n676bar);
  OR2_X1 U292 ( .A1(in_60), .A2(in_6), .ZN(n671) );
  AND2_X1 U292bar ( .A1(in_60bar), .A2(in_6bar), .ZN(n671bar);
  OR2_X1 U293 ( .A1(in_77), .A2(in_69), .ZN(n672) );
  AND2_X1 U293bar ( .A1(in_77bar), .A2(in_69bar), .ZN(n672bar);
  OR2_X1 U294 ( .A1(in[113]), .A2(n864), .ZN(n700) );
  AND2_X1 U294bar ( .A1(inbar[113]), .A2(n864bar), .ZN(n700bar);
  OR2_X1 U295 ( .A1(n670), .A2(n669), .ZN(n864) );
  AND2_X1 U295bar ( .A1(n670bar), .A2(n669bar), .ZN(n864bar);
  OR2_X1 U296 ( .A1(n668), .A2(n667), .ZN(n669) );
  AND2_X1 U296bar ( .A1(n668bar), .A2(n667bar), .ZN(n669bar);
  OR2_X1 U297 ( .A1(n666), .A2(n665), .ZN(n667) );
  AND2_X1 U297bar ( .A1(n666bar), .A2(n665bar), .ZN(n667bar);
  OR2_X1 U298 ( .A1(in[125]), .A2(in[107]), .ZN(n665) );
  AND2_X1 U298bar ( .A1(inbar[125]), .A2(inbar[107]), .ZN(n665bar);
  OR2_X1 U299 ( .A1(in[138]), .A2(in[126]), .ZN(n666) );
  AND2_X1 U299bar ( .A1(inbar[138]), .A2(inbar[126]), .ZN(n666bar);
  OR2_X1 U300 ( .A1(n664), .A2(n663), .ZN(n668) );
  AND2_X1 U300bar ( .A1(n664bar), .A2(n663bar), .ZN(n668bar);
  OR2_X1 U301 ( .A1(in[189]), .A2(in[143]), .ZN(n663) );
  AND2_X1 U301bar ( .A1(inbar[189]), .A2(inbar[143]), .ZN(n663bar);
  OR2_X1 U302 ( .A1(in[99]), .A2(in[214]), .ZN(n664) );
  AND2_X1 U302bar ( .A1(inbar[99]), .A2(inbar[214]), .ZN(n664bar);
  OR2_X1 U303 ( .A1(n662), .A2(n661), .ZN(n670) );
  AND2_X1 U303bar ( .A1(n662bar), .A2(n661bar), .ZN(n670bar);
  OR2_X1 U304 ( .A1(n660), .A2(n659), .ZN(n661) );
  AND2_X1 U304bar ( .A1(n660bar), .A2(n659bar), .ZN(n661bar);
  OR2_X1 U305 ( .A1(in_15), .A2(in_12), .ZN(n659) );
  AND2_X1 U305bar ( .A1(in_15bar), .A2(in_12bar), .ZN(n659bar);
  OR2_X1 U306 ( .A1(in_20), .A2(in_2), .ZN(n660) );
  AND2_X1 U306bar ( .A1(in_20bar), .A2(in_2bar), .ZN(n660bar);
  OR2_X1 U307 ( .A1(n658), .A2(n657), .ZN(n662) );
  AND2_X1 U307bar ( .A1(n658bar), .A2(n657bar), .ZN(n662bar);
  OR2_X1 U308 ( .A1(in_30), .A2(in_3), .ZN(n657) );
  AND2_X1 U308bar ( .A1(in_30bar), .A2(in_3bar), .ZN(n657bar);
  OR2_X1 U309 ( .A1(in_4), .A2(in_38), .ZN(n658) );
  AND2_X1 U309bar ( .A1(in_4bar), .A2(in_38bar), .ZN(n658bar);
  OR2_X1 U310 ( .A1(n656), .A2(n655), .ZN(n702) );
  AND2_X1 U310bar ( .A1(n656bar), .A2(n655bar), .ZN(n702bar);
  OR2_X1 U311 ( .A1(in[148]), .A2(in[137]), .ZN(n655) );
  AND2_X1 U311bar ( .A1(inbar[148]), .A2(inbar[137]), .ZN(n655bar);
  OR2_X1 U312 ( .A1(in[149]), .A2(n654), .ZN(n656) );
  AND2_X1 U312bar ( .A1(inbar[149]), .A2(n654bar), .ZN(n656bar);
  OR2_X1 U313 ( .A1(in[195]), .A2(in[190]), .ZN(n654) );
  AND2_X1 U313bar ( .A1(inbar[195]), .A2(inbar[190]), .ZN(n654bar);
  OR2_X1 U314 ( .A1(n653), .A2(n652), .ZN(n704) );
  AND2_X1 U314bar ( .A1(n653bar), .A2(n652bar), .ZN(n704bar);
  OR2_X1 U315 ( .A1(n651), .A2(n650), .ZN(n652) );
  AND2_X1 U315bar ( .A1(n651bar), .A2(n650bar), .ZN(n652bar);
  OR2_X1 U316 ( .A1(in[98]), .A2(in[197]), .ZN(n650) );
  AND2_X1 U316bar ( .A1(inbar[98]), .A2(inbar[197]), .ZN(n650bar);
  OR2_X1 U317 ( .A1(in_11), .A2(n649), .ZN(n651) );
  AND2_X1 U317bar ( .A1(in_11bar), .A2(n649bar), .ZN(n651bar);
  OR2_X1 U318 ( .A1(in_26), .A2(in_14), .ZN(n649) );
  AND2_X1 U318bar ( .A1(in_26bar), .A2(in_14bar), .ZN(n649bar);
  OR2_X1 U319 ( .A1(n648), .A2(n647), .ZN(n653) );
  AND2_X1 U319bar ( .A1(n648bar), .A2(n647bar), .ZN(n653bar);
  OR2_X1 U320 ( .A1(in_35), .A2(in_27), .ZN(n647) );
  AND2_X1 U320bar ( .A1(in_35bar), .A2(in_27bar), .ZN(n647bar);
  OR2_X1 U321 ( .A1(in_50), .A2(n646), .ZN(n648) );
  AND2_X1 U321bar ( .A1(in_50bar), .A2(n646bar), .ZN(n648bar);
  OR2_X1 U322 ( .A1(in_78), .A2(in_61), .ZN(n646) );
  AND2_X1 U322bar ( .A1(in_78bar), .A2(in_61bar), .ZN(n646bar);
  OR2_X1 U323 ( .A1(n942), .A2(n645), .ZN(n720) );
  AND2_X1 U323bar ( .A1(n942bar), .A2(n645bar), .ZN(n720bar);
  OR2_X1 U324 ( .A1(in[106]), .A2(n863), .ZN(n645) );
  AND2_X1 U324bar ( .A1(inbar[106]), .A2(n863bar), .ZN(n645bar);
  OR2_X1 U325 ( .A1(n644), .A2(n643), .ZN(n863) );
  AND2_X1 U325bar ( .A1(n644bar), .A2(n643bar), .ZN(n863bar);
  OR2_X1 U326 ( .A1(n642), .A2(n641), .ZN(n643) );
  AND2_X1 U326bar ( .A1(n642bar), .A2(n641bar), .ZN(n643bar);
  OR2_X1 U327 ( .A1(n640), .A2(n639), .ZN(n641) );
  AND2_X1 U327bar ( .A1(n640bar), .A2(n639bar), .ZN(n641bar);
  OR2_X1 U328 ( .A1(in[127]), .A2(in[122]), .ZN(n639) );
  AND2_X1 U328bar ( .A1(inbar[127]), .A2(inbar[122]), .ZN(n639bar);
  OR2_X1 U329 ( .A1(in[156]), .A2(in[132]), .ZN(n640) );
  AND2_X1 U329bar ( .A1(inbar[156]), .A2(inbar[132]), .ZN(n640bar);
  OR2_X1 U330 ( .A1(n638), .A2(n637), .ZN(n642) );
  AND2_X1 U330bar ( .A1(n638bar), .A2(n637bar), .ZN(n642bar);
  OR2_X1 U331 ( .A1(in[159]), .A2(in[157]), .ZN(n637) );
  AND2_X1 U331bar ( .A1(inbar[159]), .A2(inbar[157]), .ZN(n637bar);
  OR2_X1 U332 ( .A1(in[185]), .A2(in[169]), .ZN(n638) );
  AND2_X1 U332bar ( .A1(inbar[185]), .A2(inbar[169]), .ZN(n638bar);
  OR2_X1 U333 ( .A1(n636), .A2(n635), .ZN(n644) );
  AND2_X1 U333bar ( .A1(n636bar), .A2(n635bar), .ZN(n644bar);
  OR2_X1 U334 ( .A1(n634), .A2(n633), .ZN(n635) );
  AND2_X1 U334bar ( .A1(n634bar), .A2(n633bar), .ZN(n635bar);
  OR2_X1 U335 ( .A1(in[239]), .A2(in[218]), .ZN(n633) );
  AND2_X1 U335bar ( .A1(inbar[239]), .A2(inbar[218]), .ZN(n633bar);
  OR2_X1 U336 ( .A1(in_13), .A2(in[87]), .ZN(n634) );
  AND2_X1 U336bar ( .A1(in_13bar), .A2(inbar[87]), .ZN(n634bar);
  OR2_X1 U337 ( .A1(n632), .A2(n631), .ZN(n636) );
  AND2_X1 U337bar ( .A1(n632bar), .A2(n631bar), .ZN(n636bar);
  OR2_X1 U338 ( .A1(in_72), .A2(in_70), .ZN(n631) );
  AND2_X1 U338bar ( .A1(in_72bar), .A2(in_70bar), .ZN(n631bar);
  OR2_X1 U339 ( .A1(in_80), .A2(in_74), .ZN(n632) );
  AND2_X1 U339bar ( .A1(in_80bar), .A2(in_74bar), .ZN(n632bar);
  OR2_X1 U340 ( .A1(n630), .A2(n629), .ZN(n942) );
  AND2_X1 U340bar ( .A1(n630bar), .A2(n629bar), .ZN(n942bar);
  OR2_X1 U341 ( .A1(n628), .A2(n627), .ZN(n629) );
  AND2_X1 U341bar ( .A1(n628bar), .A2(n627bar), .ZN(n629bar);
  OR2_X1 U342 ( .A1(n626), .A2(n625), .ZN(n627) );
  AND2_X1 U342bar ( .A1(n626bar), .A2(n625bar), .ZN(n627bar);
  OR2_X1 U343 ( .A1(in[146]), .A2(in[100]), .ZN(n625) );
  AND2_X1 U343bar ( .A1(inbar[146]), .A2(inbar[100]), .ZN(n625bar);
  OR2_X1 U344 ( .A1(in[168]), .A2(in[152]), .ZN(n626) );
  AND2_X1 U344bar ( .A1(inbar[168]), .A2(inbar[152]), .ZN(n626bar);
  OR2_X1 U345 ( .A1(n624), .A2(n623), .ZN(n628) );
  AND2_X1 U345bar ( .A1(n624bar), .A2(n623bar), .ZN(n628bar);
  OR2_X1 U346 ( .A1(in[199]), .A2(in[182]), .ZN(n623) );
  AND2_X1 U346bar ( .A1(inbar[199]), .A2(inbar[182]), .ZN(n623bar);
  OR2_X1 U347 ( .A1(in[236]), .A2(in[204]), .ZN(n624) );
  AND2_X1 U347bar ( .A1(inbar[236]), .A2(inbar[204]), .ZN(n624bar);
  OR2_X1 U348 ( .A1(n622), .A2(n621), .ZN(n630) );
  AND2_X1 U348bar ( .A1(n622bar), .A2(n621bar), .ZN(n630bar);
  OR2_X1 U349 ( .A1(n620), .A2(n619), .ZN(n621) );
  AND2_X1 U349bar ( .A1(n620bar), .A2(n619bar), .ZN(n621bar);
  OR2_X1 U350 ( .A1(in[89]), .A2(in[246]), .ZN(n619) );
  AND2_X1 U350bar ( .A1(inbar[89]), .A2(inbar[246]), .ZN(n619bar);
  OR2_X1 U351 ( .A1(in[95]), .A2(in[92]), .ZN(n620) );
  AND2_X1 U351bar ( .A1(inbar[95]), .A2(inbar[92]), .ZN(n620bar);
  OR2_X1 U352 ( .A1(n618), .A2(n617), .ZN(n622) );
  AND2_X1 U352bar ( .A1(n618bar), .A2(n617bar), .ZN(n622bar);
  OR2_X1 U353 ( .A1(in_22), .A2(in_16), .ZN(n617) );
  AND2_X1 U353bar ( .A1(in_22bar), .A2(in_16bar), .ZN(n617bar);
  OR2_X1 U354 ( .A1(in_51), .A2(in_49), .ZN(n618) );
  AND2_X1 U354bar ( .A1(in_51bar), .A2(in_49bar), .ZN(n618bar);
  OR2_X1 U355 ( .A1(n616), .A2(n615), .ZN(n722) );
  AND2_X1 U355bar ( .A1(n616bar), .A2(n615bar), .ZN(n722bar);
  OR2_X1 U356 ( .A1(in[158]), .A2(in[115]), .ZN(n615) );
  AND2_X1 U356bar ( .A1(inbar[158]), .A2(inbar[115]), .ZN(n615bar);
  OR2_X1 U357 ( .A1(in[163]), .A2(n614), .ZN(n616) );
  AND2_X1 U357bar ( .A1(inbar[163]), .A2(n614bar), .ZN(n616bar);
  OR2_X1 U358 ( .A1(in[206]), .A2(in[165]), .ZN(n614) );
  AND2_X1 U358bar ( .A1(inbar[206]), .A2(inbar[165]), .ZN(n614bar);
  OR2_X1 U359 ( .A1(n613), .A2(n612), .ZN(n724) );
  AND2_X1 U359bar ( .A1(n613bar), .A2(n612bar), .ZN(n724bar);
  OR2_X1 U360 ( .A1(n611), .A2(n610), .ZN(n612) );
  AND2_X1 U360bar ( .A1(n611bar), .A2(n610bar), .ZN(n612bar);
  OR2_X1 U361 ( .A1(in[213]), .A2(in[207]), .ZN(n610) );
  AND2_X1 U361bar ( .A1(inbar[213]), .A2(inbar[207]), .ZN(n610bar);
  OR2_X1 U362 ( .A1(in[215]), .A2(n609), .ZN(n611) );
  AND2_X1 U362bar ( .A1(inbar[215]), .A2(n609bar), .ZN(n611bar);
  OR2_X1 U363 ( .A1(in[230]), .A2(in[220]), .ZN(n609) );
  AND2_X1 U363bar ( .A1(inbar[230]), .A2(inbar[220]), .ZN(n609bar);
  OR2_X1 U364 ( .A1(n608), .A2(n607), .ZN(n613) );
  AND2_X1 U364bar ( .A1(n608bar), .A2(n607bar), .ZN(n613bar);
  OR2_X1 U365 ( .A1(in[251]), .A2(in[234]), .ZN(n607) );
  AND2_X1 U365bar ( .A1(inbar[251]), .A2(inbar[234]), .ZN(n607bar);
  OR2_X1 U366 ( .A1(in_17), .A2(n606), .ZN(n608) );
  AND2_X1 U366bar ( .A1(in_17bar), .A2(n606bar), .ZN(n608bar);
  OR2_X1 U367 ( .A1(in_65), .A2(in_56), .ZN(n606) );
  AND2_X1 U367bar ( .A1(in_65bar), .A2(in_56bar), .ZN(n606bar);
  OR2_X1 U368 ( .A1(n605), .A2(n604), .ZN(out[0]) );
  AND2_X1 U368bar ( .A1(n605bar), .A2(n604bar), .ZN(outbar[0]);
  OR2_X1 U369 ( .A1(n603), .A2(n602), .ZN(n604) );
  AND2_X1 U369bar ( .A1(n603bar), .A2(n602bar), .ZN(n604bar);
  OR2_X1 U370 ( .A1(n601), .A2(n600), .ZN(n602) );
  AND2_X1 U370bar ( .A1(n601bar), .A2(n600bar), .ZN(n602bar);
  OR2_X1 U371 ( .A1(n820), .A2(n785), .ZN(n600) );
  AND2_X1 U371bar ( .A1(n820bar), .A2(n785bar), .ZN(n600bar);
  OR2_X1 U372 ( .A1(n599), .A2(n598), .ZN(n785) );
  AND2_X1 U372bar ( .A1(n599bar), .A2(n598bar), .ZN(n785bar);
  OR2_X1 U373 ( .A1(n597), .A2(n596), .ZN(n598) );
  AND2_X1 U373bar ( .A1(n597bar), .A2(n596bar), .ZN(n598bar);
  OR2_X1 U374 ( .A1(n595), .A2(n594), .ZN(n596) );
  AND2_X1 U374bar ( .A1(n595bar), .A2(n594bar), .ZN(n596bar);
  OR2_X1 U375 ( .A1(in[135]), .A2(in[104]), .ZN(n594) );
  AND2_X1 U375bar ( .A1(inbar[135]), .A2(inbar[104]), .ZN(n594bar);
  OR2_X1 U376 ( .A1(in[188]), .A2(in[178]), .ZN(n595) );
  AND2_X1 U376bar ( .A1(inbar[188]), .A2(inbar[178]), .ZN(n595bar);
  OR2_X1 U377 ( .A1(n593), .A2(n592), .ZN(n597) );
  AND2_X1 U377bar ( .A1(n593bar), .A2(n592bar), .ZN(n597bar);
  OR2_X1 U378 ( .A1(in[217]), .A2(in[194]), .ZN(n592) );
  AND2_X1 U378bar ( .A1(inbar[217]), .A2(inbar[194]), .ZN(n592bar);
  OR2_X1 U379 ( .A1(in[237]), .A2(in[218]), .ZN(n593) );
  AND2_X1 U379bar ( .A1(inbar[237]), .A2(inbar[218]), .ZN(n593bar);
  OR2_X1 U380 ( .A1(n591), .A2(n590), .ZN(n599) );
  AND2_X1 U380bar ( .A1(n591bar), .A2(n590bar), .ZN(n599bar);
  OR2_X1 U381 ( .A1(n589), .A2(n588), .ZN(n590) );
  AND2_X1 U381bar ( .A1(n589bar), .A2(n588bar), .ZN(n590bar);
  OR2_X1 U382 ( .A1(in_2), .A2(in_10), .ZN(n588) );
  AND2_X1 U382bar ( .A1(in_2bar), .A2(in_10bar), .ZN(n588bar);
  OR2_X1 U383 ( .A1(in_47), .A2(in_22), .ZN(n589) );
  AND2_X1 U383bar ( .A1(in_47bar), .A2(in_22bar), .ZN(n589bar);
  OR2_X1 U384 ( .A1(n587), .A2(n586), .ZN(n591) );
  AND2_X1 U384bar ( .A1(n587bar), .A2(n586bar), .ZN(n591bar);
  OR2_X1 U385 ( .A1(in_56), .A2(in_54), .ZN(n586) );
  AND2_X1 U385bar ( .A1(in_56bar), .A2(in_54bar), .ZN(n586bar);
  OR2_X1 U386 ( .A1(in_63), .A2(in_61), .ZN(n587) );
  AND2_X1 U386bar ( .A1(in_63bar), .A2(in_61bar), .ZN(n587bar);
  OR2_X1 U387 ( .A1(n585), .A2(n584), .ZN(n820) );
  AND2_X1 U387bar ( .A1(n585bar), .A2(n584bar), .ZN(n820bar);
  OR2_X1 U388 ( .A1(n583), .A2(n582), .ZN(n584) );
  AND2_X1 U388bar ( .A1(n583bar), .A2(n582bar), .ZN(n584bar);
  OR2_X1 U389 ( .A1(n581), .A2(n580), .ZN(n582) );
  AND2_X1 U389bar ( .A1(n581bar), .A2(n580bar), .ZN(n582bar);
  OR2_X1 U390 ( .A1(in[158]), .A2(in[142]), .ZN(n580) );
  AND2_X1 U390bar ( .A1(inbar[158]), .A2(inbar[142]), .ZN(n580bar);
  OR2_X1 U391 ( .A1(in[175]), .A2(in[164]), .ZN(n581) );
  AND2_X1 U391bar ( .A1(inbar[175]), .A2(inbar[164]), .ZN(n581bar);
  OR2_X1 U392 ( .A1(n579), .A2(n578), .ZN(n583) );
  AND2_X1 U392bar ( .A1(n579bar), .A2(n578bar), .ZN(n583bar);
  OR2_X1 U393 ( .A1(in[228]), .A2(in[204]), .ZN(n578) );
  AND2_X1 U393bar ( .A1(inbar[228]), .A2(inbar[204]), .ZN(n578bar);
  OR2_X1 U394 ( .A1(in[91]), .A2(in[87]), .ZN(n579) );
  AND2_X1 U394bar ( .A1(inbar[91]), .A2(inbar[87]), .ZN(n579bar);
  OR2_X1 U395 ( .A1(n577), .A2(n576), .ZN(n585) );
  AND2_X1 U395bar ( .A1(n577bar), .A2(n576bar), .ZN(n585bar);
  OR2_X1 U396 ( .A1(n575), .A2(n574), .ZN(n576) );
  AND2_X1 U396bar ( .A1(n575bar), .A2(n574bar), .ZN(n576bar);
  OR2_X1 U397 ( .A1(in_21), .A2(in_11), .ZN(n574) );
  AND2_X1 U397bar ( .A1(in_21bar), .A2(in_11bar), .ZN(n574bar);
  OR2_X1 U398 ( .A1(in_5), .A2(in_3), .ZN(n575) );
  AND2_X1 U398bar ( .A1(in_5bar), .A2(in_3bar), .ZN(n575bar);
  OR2_X1 U399 ( .A1(n573), .A2(n572), .ZN(n577) );
  AND2_X1 U399bar ( .A1(n573bar), .A2(n572bar), .ZN(n577bar);
  OR2_X1 U400 ( .A1(in_68), .A2(in_64), .ZN(n572) );
  AND2_X1 U400bar ( .A1(in_68bar), .A2(in_64bar), .ZN(n572bar);
  OR2_X1 U401 ( .A1(in_76), .A2(in_73), .ZN(n573) );
  AND2_X1 U401bar ( .A1(in_76bar), .A2(in_73bar), .ZN(n573bar);
  OR2_X1 U402 ( .A1(n778), .A2(n571), .ZN(n601) );
  AND2_X1 U402bar ( .A1(n778bar), .A2(n571bar), .ZN(n601bar);
  OR2_X1 U403 ( .A1(in[100]), .A2(n965), .ZN(n571) );
  AND2_X1 U403bar ( .A1(inbar[100]), .A2(n965bar), .ZN(n571bar);
  OR2_X1 U404 ( .A1(n570), .A2(n569), .ZN(n965) );
  AND2_X1 U404bar ( .A1(n570bar), .A2(n569bar), .ZN(n965bar);
  OR2_X1 U405 ( .A1(n568), .A2(n567), .ZN(n569) );
  AND2_X1 U405bar ( .A1(n568bar), .A2(n567bar), .ZN(n569bar);
  OR2_X1 U406 ( .A1(n566), .A2(n565), .ZN(n567) );
  AND2_X1 U406bar ( .A1(n566bar), .A2(n565bar), .ZN(n567bar);
  OR2_X1 U407 ( .A1(n817), .A2(n750), .ZN(n565) );
  AND2_X1 U407bar ( .A1(n817bar), .A2(n750bar), .ZN(n565bar);
  OR2_X1 U408 ( .A1(n564), .A2(n563), .ZN(n750) );
  AND2_X1 U408bar ( .A1(n564bar), .A2(n563bar), .ZN(n750bar);
  OR2_X1 U409 ( .A1(n562), .A2(n561), .ZN(n563) );
  AND2_X1 U409bar ( .A1(n562bar), .A2(n561bar), .ZN(n563bar);
  OR2_X1 U410 ( .A1(n560), .A2(n559), .ZN(n561) );
  AND2_X1 U410bar ( .A1(n560bar), .A2(n559bar), .ZN(n561bar);
  OR2_X1 U411 ( .A1(in[119]), .A2(in[103]), .ZN(n559) );
  AND2_X1 U411bar ( .A1(inbar[119]), .A2(inbar[103]), .ZN(n559bar);
  OR2_X1 U412 ( .A1(in[137]), .A2(in[133]), .ZN(n560) );
  AND2_X1 U412bar ( .A1(inbar[137]), .A2(inbar[133]), .ZN(n560bar);
  OR2_X1 U413 ( .A1(n558), .A2(n557), .ZN(n562) );
  AND2_X1 U413bar ( .A1(n558bar), .A2(n557bar), .ZN(n562bar);
  OR2_X1 U414 ( .A1(in[176]), .A2(in[173]), .ZN(n557) );
  AND2_X1 U414bar ( .A1(inbar[176]), .A2(inbar[173]), .ZN(n557bar);
  OR2_X1 U415 ( .A1(in[210]), .A2(in[181]), .ZN(n558) );
  AND2_X1 U415bar ( .A1(inbar[210]), .A2(inbar[181]), .ZN(n558bar);
  OR2_X1 U416 ( .A1(n556), .A2(n555), .ZN(n564) );
  AND2_X1 U416bar ( .A1(n556bar), .A2(n555bar), .ZN(n564bar);
  OR2_X1 U417 ( .A1(n554), .A2(n553), .ZN(n555) );
  AND2_X1 U417bar ( .A1(n554bar), .A2(n553bar), .ZN(n555bar);
  OR2_X1 U418 ( .A1(in_13), .A2(in[234]), .ZN(n553) );
  AND2_X1 U418bar ( .A1(in_13bar), .A2(inbar[234]), .ZN(n553bar);
  OR2_X1 U419 ( .A1(in_38), .A2(in_32), .ZN(n554) );
  AND2_X1 U419bar ( .A1(in_38bar), .A2(in_32bar), .ZN(n554bar);
  OR2_X1 U420 ( .A1(n552), .A2(n551), .ZN(n556) );
  AND2_X1 U420bar ( .A1(n552bar), .A2(n551bar), .ZN(n556bar);
  OR2_X1 U421 ( .A1(in_42), .A2(in_41), .ZN(n551) );
  AND2_X1 U421bar ( .A1(in_42bar), .A2(in_41bar), .ZN(n551bar);
  OR2_X1 U422 ( .A1(in_7), .A2(in_49), .ZN(n552) );
  AND2_X1 U422bar ( .A1(in_7bar), .A2(in_49bar), .ZN(n552bar);
  OR2_X1 U423 ( .A1(n550), .A2(n549), .ZN(n817) );
  AND2_X1 U423bar ( .A1(n550bar), .A2(n549bar), .ZN(n817bar);
  OR2_X1 U424 ( .A1(n548), .A2(n547), .ZN(n549) );
  AND2_X1 U424bar ( .A1(n548bar), .A2(n547bar), .ZN(n549bar);
  OR2_X1 U425 ( .A1(n546), .A2(n545), .ZN(n547) );
  AND2_X1 U425bar ( .A1(n546bar), .A2(n545bar), .ZN(n547bar);
  OR2_X1 U426 ( .A1(in[159]), .A2(in[105]), .ZN(n545) );
  AND2_X1 U426bar ( .A1(inbar[159]), .A2(inbar[105]), .ZN(n545bar);
  OR2_X1 U427 ( .A1(in[206]), .A2(in[183]), .ZN(n546) );
  AND2_X1 U427bar ( .A1(inbar[206]), .A2(inbar[183]), .ZN(n546bar);
  OR2_X1 U428 ( .A1(n544), .A2(n543), .ZN(n548) );
  AND2_X1 U428bar ( .A1(n544bar), .A2(n543bar), .ZN(n548bar);
  OR2_X1 U429 ( .A1(in[229]), .A2(in[219]), .ZN(n543) );
  AND2_X1 U429bar ( .A1(inbar[229]), .A2(inbar[219]), .ZN(n543bar);
  OR2_X1 U430 ( .A1(in[235]), .A2(in[232]), .ZN(n544) );
  AND2_X1 U430bar ( .A1(inbar[235]), .A2(inbar[232]), .ZN(n544bar);
  OR2_X1 U431 ( .A1(n542), .A2(n541), .ZN(n550) );
  AND2_X1 U431bar ( .A1(n542bar), .A2(n541bar), .ZN(n550bar);
  OR2_X1 U432 ( .A1(n540), .A2(n539), .ZN(n541) );
  AND2_X1 U432bar ( .A1(n540bar), .A2(n539bar), .ZN(n541bar);
  OR2_X1 U433 ( .A1(in[249]), .A2(in[242]), .ZN(n539) );
  AND2_X1 U433bar ( .A1(inbar[249]), .A2(inbar[242]), .ZN(n539bar);
  OR2_X1 U434 ( .A1(in[89]), .A2(in[254]), .ZN(n540) );
  AND2_X1 U434bar ( .A1(inbar[89]), .A2(inbar[254]), .ZN(n540bar);
  OR2_X1 U435 ( .A1(n538), .A2(n537), .ZN(n542) );
  AND2_X1 U435bar ( .A1(n538bar), .A2(n537bar), .ZN(n542bar);
  OR2_X1 U436 ( .A1(in_14), .A2(in[99]), .ZN(n537) );
  AND2_X1 U436bar ( .A1(in_14bar), .A2(inbar[99]), .ZN(n537bar);
  OR2_X1 U437 ( .A1(in_60), .A2(in_18), .ZN(n538) );
  AND2_X1 U437bar ( .A1(in_60bar), .A2(in_18bar), .ZN(n538bar);
  OR2_X1 U438 ( .A1(in[113]), .A2(n763), .ZN(n566) );
  AND2_X1 U438bar ( .A1(inbar[113]), .A2(n763bar), .ZN(n566bar);
  OR2_X1 U439 ( .A1(n536), .A2(n535), .ZN(n763) );
  AND2_X1 U439bar ( .A1(n536bar), .A2(n535bar), .ZN(n763bar);
  OR2_X1 U440 ( .A1(n534), .A2(n533), .ZN(n535) );
  AND2_X1 U440bar ( .A1(n534bar), .A2(n533bar), .ZN(n535bar);
  OR2_X1 U441 ( .A1(n532), .A2(n531), .ZN(n533) );
  AND2_X1 U441bar ( .A1(n532bar), .A2(n531bar), .ZN(n533bar);
  OR2_X1 U442 ( .A1(in[115]), .A2(in[110]), .ZN(n531) );
  AND2_X1 U442bar ( .A1(inbar[115]), .A2(inbar[110]), .ZN(n531bar);
  OR2_X1 U443 ( .A1(in[125]), .A2(in[117]), .ZN(n532) );
  AND2_X1 U443bar ( .A1(inbar[125]), .A2(inbar[117]), .ZN(n532bar);
  OR2_X1 U444 ( .A1(n530), .A2(n529), .ZN(n534) );
  AND2_X1 U444bar ( .A1(n530bar), .A2(n529bar), .ZN(n534bar);
  OR2_X1 U445 ( .A1(in[180]), .A2(in[128]), .ZN(n529) );
  AND2_X1 U445bar ( .A1(inbar[180]), .A2(inbar[128]), .ZN(n529bar);
  OR2_X1 U446 ( .A1(in[205]), .A2(in[201]), .ZN(n530) );
  AND2_X1 U446bar ( .A1(inbar[205]), .A2(inbar[201]), .ZN(n530bar);
  OR2_X1 U447 ( .A1(n528), .A2(n527), .ZN(n536) );
  AND2_X1 U447bar ( .A1(n528bar), .A2(n527bar), .ZN(n536bar);
  OR2_X1 U448 ( .A1(n526), .A2(n525), .ZN(n527) );
  AND2_X1 U448bar ( .A1(n526bar), .A2(n525bar), .ZN(n527bar);
  OR2_X1 U449 ( .A1(in[244]), .A2(in[239]), .ZN(n525) );
  AND2_X1 U449bar ( .A1(inbar[244]), .A2(inbar[239]), .ZN(n525bar);
  OR2_X1 U450 ( .A1(in[95]), .A2(in[83]), .ZN(n526) );
  AND2_X1 U450bar ( .A1(inbar[95]), .A2(inbar[83]), .ZN(n526bar);
  OR2_X1 U451 ( .A1(n524), .A2(n523), .ZN(n528) );
  AND2_X1 U451bar ( .A1(n524bar), .A2(n523bar), .ZN(n528bar);
  OR2_X1 U452 ( .A1(in_24), .A2(in[97]), .ZN(n523) );
  AND2_X1 U452bar ( .A1(in_24bar), .A2(inbar[97]), .ZN(n523bar);
  OR2_X1 U453 ( .A1(in_33), .A2(in_27), .ZN(n524) );
  AND2_X1 U453bar ( .A1(in_33bar), .A2(in_27bar), .ZN(n524bar);
  OR2_X1 U454 ( .A1(n522), .A2(n521), .ZN(n568) );
  AND2_X1 U454bar ( .A1(n522bar), .A2(n521bar), .ZN(n568bar);
  OR2_X1 U455 ( .A1(in[145]), .A2(in[126]), .ZN(n521) );
  AND2_X1 U455bar ( .A1(inbar[145]), .A2(inbar[126]), .ZN(n521bar);
  OR2_X1 U456 ( .A1(in[169]), .A2(n520), .ZN(n522) );
  AND2_X1 U456bar ( .A1(inbar[169]), .A2(n520bar), .ZN(n522bar);
  OR2_X1 U457 ( .A1(in[221]), .A2(in[172]), .ZN(n520) );
  AND2_X1 U457bar ( .A1(inbar[221]), .A2(inbar[172]), .ZN(n520bar);
  OR2_X1 U458 ( .A1(n519), .A2(n518), .ZN(n570) );
  AND2_X1 U458bar ( .A1(n519bar), .A2(n518bar), .ZN(n570bar);
  OR2_X1 U459 ( .A1(n517), .A2(n516), .ZN(n518) );
  AND2_X1 U459bar ( .A1(n517bar), .A2(n516bar), .ZN(n518bar);
  OR2_X1 U460 ( .A1(in[241]), .A2(in[224]), .ZN(n516) );
  AND2_X1 U460bar ( .A1(inbar[241]), .A2(inbar[224]), .ZN(n516bar);
  OR2_X1 U461 ( .A1(in[86]), .A2(n515), .ZN(n517) );
  AND2_X1 U461bar ( .A1(inbar[86]), .A2(n515bar), .ZN(n517bar);
  OR2_X1 U462 ( .A1(in_43), .A2(in_34), .ZN(n515) );
  AND2_X1 U462bar ( .A1(in_43bar), .A2(in_34bar), .ZN(n515bar);
  OR2_X1 U463 ( .A1(n514), .A2(n513), .ZN(n519) );
  AND2_X1 U463bar ( .A1(n514bar), .A2(n513bar), .ZN(n519bar);
  OR2_X1 U464 ( .A1(in_65), .A2(in_51), .ZN(n513) );
  AND2_X1 U464bar ( .A1(in_65bar), .A2(in_51bar), .ZN(n513bar);
  OR2_X1 U465 ( .A1(in_75), .A2(n512), .ZN(n514) );
  AND2_X1 U465bar ( .A1(in_75bar), .A2(n512bar), .ZN(n514bar);
  OR2_X1 U466 ( .A1(in_81), .A2(in_77), .ZN(n512) );
  AND2_X1 U466bar ( .A1(in_81bar), .A2(in_77bar), .ZN(n512bar);
  OR2_X1 U467 ( .A1(n511), .A2(n510), .ZN(n778) );
  AND2_X1 U467bar ( .A1(n511bar), .A2(n510bar), .ZN(n778bar);
  OR2_X1 U468 ( .A1(n509), .A2(n508), .ZN(n510) );
  AND2_X1 U468bar ( .A1(n509bar), .A2(n508bar), .ZN(n510bar);
  OR2_X1 U469 ( .A1(n507), .A2(n506), .ZN(n508) );
  AND2_X1 U469bar ( .A1(n507bar), .A2(n506bar), .ZN(n508bar);
  OR2_X1 U470 ( .A1(in[107]), .A2(in[101]), .ZN(n506) );
  AND2_X1 U470bar ( .A1(inbar[107]), .A2(inbar[101]), .ZN(n506bar);
  OR2_X1 U471 ( .A1(in[139]), .A2(in[132]), .ZN(n507) );
  AND2_X1 U471bar ( .A1(inbar[139]), .A2(inbar[132]), .ZN(n507bar);
  OR2_X1 U472 ( .A1(n505), .A2(n504), .ZN(n509) );
  AND2_X1 U472bar ( .A1(n505bar), .A2(n504bar), .ZN(n509bar);
  OR2_X1 U473 ( .A1(in[146]), .A2(in[141]), .ZN(n504) );
  AND2_X1 U473bar ( .A1(inbar[146]), .A2(inbar[141]), .ZN(n504bar);
  OR2_X1 U474 ( .A1(in[203]), .A2(in[179]), .ZN(n505) );
  AND2_X1 U474bar ( .A1(inbar[203]), .A2(inbar[179]), .ZN(n505bar);
  OR2_X1 U475 ( .A1(n503), .A2(n502), .ZN(n511) );
  AND2_X1 U475bar ( .A1(n503bar), .A2(n502bar), .ZN(n511bar);
  OR2_X1 U476 ( .A1(n501), .A2(n500), .ZN(n502) );
  AND2_X1 U476bar ( .A1(n501bar), .A2(n500bar), .ZN(n502bar);
  OR2_X1 U477 ( .A1(in[243]), .A2(in[222]), .ZN(n500) );
  AND2_X1 U477bar ( .A1(inbar[243]), .A2(inbar[222]), .ZN(n500bar);
  OR2_X1 U478 ( .A1(in[251]), .A2(in[250]), .ZN(n501) );
  AND2_X1 U478bar ( .A1(inbar[251]), .A2(inbar[250]), .ZN(n501bar);
  OR2_X1 U479 ( .A1(n499), .A2(n498), .ZN(n503) );
  AND2_X1 U479bar ( .A1(n499bar), .A2(n498bar), .ZN(n503bar);
  OR2_X1 U480 ( .A1(in_37), .A2(in_19), .ZN(n498) );
  AND2_X1 U480bar ( .A1(in_37bar), .A2(in_19bar), .ZN(n498bar);
  OR2_X1 U481 ( .A1(in_78), .A2(in_6), .ZN(n499) );
  AND2_X1 U481bar ( .A1(in_78bar), .A2(in_6bar), .ZN(n499bar);
  OR2_X1 U482 ( .A1(n497), .A2(n496), .ZN(n603) );
  AND2_X1 U482bar ( .A1(n497bar), .A2(n496bar), .ZN(n603bar);
  OR2_X1 U483 ( .A1(in[112]), .A2(in[102]), .ZN(n496) );
  AND2_X1 U483bar ( .A1(inbar[112]), .A2(inbar[102]), .ZN(n496bar);
  OR2_X1 U484 ( .A1(in[123]), .A2(n495), .ZN(n497) );
  AND2_X1 U484bar ( .A1(inbar[123]), .A2(n495bar), .ZN(n497bar);
  OR2_X1 U485 ( .A1(in[143]), .A2(in[130]), .ZN(n495) );
  AND2_X1 U485bar ( .A1(inbar[143]), .A2(inbar[130]), .ZN(n495bar);
  OR2_X1 U486 ( .A1(n494), .A2(n493), .ZN(n605) );
  AND2_X1 U486bar ( .A1(n494bar), .A2(n493bar), .ZN(n605bar);
  OR2_X1 U487 ( .A1(n492), .A2(n491), .ZN(n493) );
  AND2_X1 U487bar ( .A1(n492bar), .A2(n491bar), .ZN(n493bar);
  OR2_X1 U488 ( .A1(in[216]), .A2(in[213]), .ZN(n491) );
  AND2_X1 U488bar ( .A1(inbar[216]), .A2(inbar[213]), .ZN(n491bar);
  OR2_X1 U489 ( .A1(in[227]), .A2(n490), .ZN(n492) );
  AND2_X1 U489bar ( .A1(inbar[227]), .A2(n490bar), .ZN(n492bar);
  OR2_X1 U490 ( .A1(in_0), .A2(in[248]), .ZN(n490) );
  AND2_X1 U490bar ( .A1(in_0bar), .A2(inbar[248]), .ZN(n490bar);
  OR2_X1 U491 ( .A1(n489), .A2(n488), .ZN(n494) );
  AND2_X1 U491bar ( .A1(n489bar), .A2(n488bar), .ZN(n494bar);
  OR2_X1 U492 ( .A1(in_46), .A2(in_44), .ZN(n488) );
  AND2_X1 U492bar ( .A1(in_46bar), .A2(in_44bar), .ZN(n488bar);
  OR2_X1 U493 ( .A1(in_50), .A2(n487), .ZN(n489) );
  AND2_X1 U493bar ( .A1(in_50bar), .A2(n487bar), .ZN(n489bar);
  OR2_X1 U494 ( .A1(in_9), .A2(in_80), .ZN(n487) );
  AND2_X1 U494bar ( .A1(in_9bar), .A2(in_80bar), .ZN(n487bar);
endmodule




module sBox_9 ( in, out );
  input [7:0] in;
  //input_done

  output [7:0] out;
  //output_done

  wire   [255:0] decodeOut;
  //wire_done

  decode_9 dec ( .in(in), .out(decodeOut) );
  encode_9 enc ( .in(decodeOut), .out(out) );
endmodule


module CD2_37 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_38 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_39 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_40 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD4_19 ( a, b, y );
  input [3:0] a;
  input [3:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  //input_done

  output [15:0] y;
  reg [15:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]);
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]);
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]);
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]);
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]);
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]);
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]);
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]);
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]);
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]);
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]);
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]);
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]);
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]);
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]);
endmodule




module CD4_20 ( a, b, y );
  input [3:0] a;
  input [3:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  //input_done

  output [15:0] y;
  reg [15:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]);
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]);
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]);
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]);
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]);
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]);
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]);
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]);
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]);
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]);
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]);
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]);
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]);
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]);
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]);
endmodule




module CD16_10 ( a, b, y );
  input [15:0] a;
  input [15:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign abar[8] = ~a[8];
  assign abar[9] = ~a[9];
  assign abar[10] = ~a[10];
  assign abar[11] = ~a[11];
  assign abar[12] = ~a[12];
  assign abar[13] = ~a[13];
  assign abar[14] = ~a[14];
  assign abar[15] = ~a[15];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign bbar[8] = ~b[8];
  assign bbar[9] = ~b[9];
  assign bbar[10] = ~b[10];
  assign bbar[11] = ~b[11];
  assign bbar[12] = ~b[12];
  assign bbar[13] = ~b[13];
  assign bbar[14] = ~b[14];
  assign bbar[15] = ~b[15];
  //input_done

  output [255:0] y;
  reg [255:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[9]), .A2(a[0]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[9]), .A2(abar[0]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[3]), .A2(a[6]), .ZN(y[99]) );
  OR2_X1 U2bar ( .A1(bbar[3]), .A2(abar[6]), .ZN(ybar[99]);
  AND2_X1 U3 ( .A1(b[2]), .A2(a[6]), .ZN(y[98]) );
  OR2_X1 U3bar ( .A1(bbar[2]), .A2(abar[6]), .ZN(ybar[98]);
  AND2_X1 U4 ( .A1(b[1]), .A2(a[6]), .ZN(y[97]) );
  OR2_X1 U4bar ( .A1(bbar[1]), .A2(abar[6]), .ZN(ybar[97]);
  AND2_X1 U5 ( .A1(b[0]), .A2(a[6]), .ZN(y[96]) );
  OR2_X1 U5bar ( .A1(bbar[0]), .A2(abar[6]), .ZN(ybar[96]);
  AND2_X1 U6 ( .A1(b[15]), .A2(a[5]), .ZN(y[95]) );
  OR2_X1 U6bar ( .A1(bbar[15]), .A2(abar[5]), .ZN(ybar[95]);
  AND2_X1 U7 ( .A1(b[14]), .A2(a[5]), .ZN(y[94]) );
  OR2_X1 U7bar ( .A1(bbar[14]), .A2(abar[5]), .ZN(ybar[94]);
  AND2_X1 U8 ( .A1(b[13]), .A2(a[5]), .ZN(y[93]) );
  OR2_X1 U8bar ( .A1(bbar[13]), .A2(abar[5]), .ZN(ybar[93]);
  AND2_X1 U9 ( .A1(b[12]), .A2(a[5]), .ZN(y[92]) );
  OR2_X1 U9bar ( .A1(bbar[12]), .A2(abar[5]), .ZN(ybar[92]);
  AND2_X1 U10 ( .A1(b[11]), .A2(a[5]), .ZN(y[91]) );
  OR2_X1 U10bar ( .A1(bbar[11]), .A2(abar[5]), .ZN(ybar[91]);
  AND2_X1 U11 ( .A1(b[10]), .A2(a[5]), .ZN(y[90]) );
  OR2_X1 U11bar ( .A1(bbar[10]), .A2(abar[5]), .ZN(ybar[90]);
  AND2_X1 U12 ( .A1(b[8]), .A2(a[0]), .ZN(y[8]) );
  OR2_X1 U12bar ( .A1(bbar[8]), .A2(abar[0]), .ZN(ybar[8]);
  AND2_X1 U13 ( .A1(a[5]), .A2(b[9]), .ZN(y[89]) );
  OR2_X1 U13bar ( .A1(abar[5]), .A2(bbar[9]), .ZN(ybar[89]);
  AND2_X1 U14 ( .A1(b[8]), .A2(a[5]), .ZN(y[88]) );
  OR2_X1 U14bar ( .A1(bbar[8]), .A2(abar[5]), .ZN(ybar[88]);
  AND2_X1 U15 ( .A1(b[7]), .A2(a[5]), .ZN(y[87]) );
  OR2_X1 U15bar ( .A1(bbar[7]), .A2(abar[5]), .ZN(ybar[87]);
  AND2_X1 U16 ( .A1(b[6]), .A2(a[5]), .ZN(y[86]) );
  OR2_X1 U16bar ( .A1(bbar[6]), .A2(abar[5]), .ZN(ybar[86]);
  AND2_X1 U17 ( .A1(b[5]), .A2(a[5]), .ZN(y[85]) );
  OR2_X1 U17bar ( .A1(bbar[5]), .A2(abar[5]), .ZN(ybar[85]);
  AND2_X1 U18 ( .A1(b[4]), .A2(a[5]), .ZN(y[84]) );
  OR2_X1 U18bar ( .A1(bbar[4]), .A2(abar[5]), .ZN(ybar[84]);
  AND2_X1 U19 ( .A1(a[5]), .A2(b[3]), .ZN(y[83]) );
  OR2_X1 U19bar ( .A1(abar[5]), .A2(bbar[3]), .ZN(ybar[83]);
  AND2_X1 U20 ( .A1(a[5]), .A2(b[2]), .ZN(y[82]) );
  OR2_X1 U20bar ( .A1(abar[5]), .A2(bbar[2]), .ZN(ybar[82]);
  AND2_X1 U21 ( .A1(a[5]), .A2(b[1]), .ZN(y[81]) );
  OR2_X1 U21bar ( .A1(abar[5]), .A2(bbar[1]), .ZN(ybar[81]);
  AND2_X1 U22 ( .A1(a[5]), .A2(b[0]), .ZN(y[80]) );
  OR2_X1 U22bar ( .A1(abar[5]), .A2(bbar[0]), .ZN(ybar[80]);
  AND2_X1 U23 ( .A1(b[7]), .A2(a[0]), .ZN(y[7]) );
  OR2_X1 U23bar ( .A1(bbar[7]), .A2(abar[0]), .ZN(ybar[7]);
  AND2_X1 U24 ( .A1(a[4]), .A2(b[15]), .ZN(y[79]) );
  OR2_X1 U24bar ( .A1(abar[4]), .A2(bbar[15]), .ZN(ybar[79]);
  AND2_X1 U25 ( .A1(a[4]), .A2(b[14]), .ZN(y[78]) );
  OR2_X1 U25bar ( .A1(abar[4]), .A2(bbar[14]), .ZN(ybar[78]);
  AND2_X1 U26 ( .A1(a[4]), .A2(b[13]), .ZN(y[77]) );
  OR2_X1 U26bar ( .A1(abar[4]), .A2(bbar[13]), .ZN(ybar[77]);
  AND2_X1 U27 ( .A1(a[4]), .A2(b[12]), .ZN(y[76]) );
  OR2_X1 U27bar ( .A1(abar[4]), .A2(bbar[12]), .ZN(ybar[76]);
  AND2_X1 U28 ( .A1(a[4]), .A2(b[11]), .ZN(y[75]) );
  OR2_X1 U28bar ( .A1(abar[4]), .A2(bbar[11]), .ZN(ybar[75]);
  AND2_X1 U29 ( .A1(a[4]), .A2(b[10]), .ZN(y[74]) );
  OR2_X1 U29bar ( .A1(abar[4]), .A2(bbar[10]), .ZN(ybar[74]);
  AND2_X1 U30 ( .A1(a[4]), .A2(b[9]), .ZN(y[73]) );
  OR2_X1 U30bar ( .A1(abar[4]), .A2(bbar[9]), .ZN(ybar[73]);
  AND2_X1 U31 ( .A1(a[4]), .A2(b[8]), .ZN(y[72]) );
  OR2_X1 U31bar ( .A1(abar[4]), .A2(bbar[8]), .ZN(ybar[72]);
  AND2_X1 U32 ( .A1(a[4]), .A2(b[7]), .ZN(y[71]) );
  OR2_X1 U32bar ( .A1(abar[4]), .A2(bbar[7]), .ZN(ybar[71]);
  AND2_X1 U33 ( .A1(a[4]), .A2(b[6]), .ZN(y[70]) );
  OR2_X1 U33bar ( .A1(abar[4]), .A2(bbar[6]), .ZN(ybar[70]);
  AND2_X1 U34 ( .A1(b[6]), .A2(a[0]), .ZN(y[6]) );
  OR2_X1 U34bar ( .A1(bbar[6]), .A2(abar[0]), .ZN(ybar[6]);
  AND2_X1 U35 ( .A1(a[4]), .A2(b[5]), .ZN(y[69]) );
  OR2_X1 U35bar ( .A1(abar[4]), .A2(bbar[5]), .ZN(ybar[69]);
  AND2_X1 U36 ( .A1(a[4]), .A2(b[4]), .ZN(y[68]) );
  OR2_X1 U36bar ( .A1(abar[4]), .A2(bbar[4]), .ZN(ybar[68]);
  AND2_X1 U37 ( .A1(a[4]), .A2(b[3]), .ZN(y[67]) );
  OR2_X1 U37bar ( .A1(abar[4]), .A2(bbar[3]), .ZN(ybar[67]);
  AND2_X1 U38 ( .A1(a[4]), .A2(b[2]), .ZN(y[66]) );
  OR2_X1 U38bar ( .A1(abar[4]), .A2(bbar[2]), .ZN(ybar[66]);
  AND2_X1 U39 ( .A1(a[4]), .A2(b[1]), .ZN(y[65]) );
  OR2_X1 U39bar ( .A1(abar[4]), .A2(bbar[1]), .ZN(ybar[65]);
  AND2_X1 U40 ( .A1(a[4]), .A2(b[0]), .ZN(y[64]) );
  OR2_X1 U40bar ( .A1(abar[4]), .A2(bbar[0]), .ZN(ybar[64]);
  AND2_X1 U41 ( .A1(a[3]), .A2(b[15]), .ZN(y[63]) );
  OR2_X1 U41bar ( .A1(abar[3]), .A2(bbar[15]), .ZN(ybar[63]);
  AND2_X1 U42 ( .A1(a[3]), .A2(b[14]), .ZN(y[62]) );
  OR2_X1 U42bar ( .A1(abar[3]), .A2(bbar[14]), .ZN(ybar[62]);
  AND2_X1 U43 ( .A1(a[3]), .A2(b[13]), .ZN(y[61]) );
  OR2_X1 U43bar ( .A1(abar[3]), .A2(bbar[13]), .ZN(ybar[61]);
  AND2_X1 U44 ( .A1(a[3]), .A2(b[12]), .ZN(y[60]) );
  OR2_X1 U44bar ( .A1(abar[3]), .A2(bbar[12]), .ZN(ybar[60]);
  AND2_X1 U45 ( .A1(b[5]), .A2(a[0]), .ZN(y[5]) );
  OR2_X1 U45bar ( .A1(bbar[5]), .A2(abar[0]), .ZN(ybar[5]);
  AND2_X1 U46 ( .A1(a[3]), .A2(b[11]), .ZN(y[59]) );
  OR2_X1 U46bar ( .A1(abar[3]), .A2(bbar[11]), .ZN(ybar[59]);
  AND2_X1 U47 ( .A1(a[3]), .A2(b[10]), .ZN(y[58]) );
  OR2_X1 U47bar ( .A1(abar[3]), .A2(bbar[10]), .ZN(ybar[58]);
  AND2_X1 U48 ( .A1(a[3]), .A2(b[9]), .ZN(y[57]) );
  OR2_X1 U48bar ( .A1(abar[3]), .A2(bbar[9]), .ZN(ybar[57]);
  AND2_X1 U49 ( .A1(a[3]), .A2(b[8]), .ZN(y[56]) );
  OR2_X1 U49bar ( .A1(abar[3]), .A2(bbar[8]), .ZN(ybar[56]);
  AND2_X1 U50 ( .A1(a[3]), .A2(b[7]), .ZN(y[55]) );
  OR2_X1 U50bar ( .A1(abar[3]), .A2(bbar[7]), .ZN(ybar[55]);
  AND2_X1 U51 ( .A1(a[3]), .A2(b[6]), .ZN(y[54]) );
  OR2_X1 U51bar ( .A1(abar[3]), .A2(bbar[6]), .ZN(ybar[54]);
  AND2_X1 U52 ( .A1(a[3]), .A2(b[5]), .ZN(y[53]) );
  OR2_X1 U52bar ( .A1(abar[3]), .A2(bbar[5]), .ZN(ybar[53]);
  AND2_X1 U53 ( .A1(a[3]), .A2(b[4]), .ZN(y[52]) );
  OR2_X1 U53bar ( .A1(abar[3]), .A2(bbar[4]), .ZN(ybar[52]);
  AND2_X1 U54 ( .A1(a[3]), .A2(b[3]), .ZN(y[51]) );
  OR2_X1 U54bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[51]);
  AND2_X1 U55 ( .A1(a[3]), .A2(b[2]), .ZN(y[50]) );
  OR2_X1 U55bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[50]);
  AND2_X1 U56 ( .A1(b[4]), .A2(a[0]), .ZN(y[4]) );
  OR2_X1 U56bar ( .A1(bbar[4]), .A2(abar[0]), .ZN(ybar[4]);
  AND2_X1 U57 ( .A1(a[3]), .A2(b[1]), .ZN(y[49]) );
  OR2_X1 U57bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[49]);
  AND2_X1 U58 ( .A1(a[3]), .A2(b[0]), .ZN(y[48]) );
  OR2_X1 U58bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[48]);
  AND2_X1 U59 ( .A1(a[2]), .A2(b[15]), .ZN(y[47]) );
  OR2_X1 U59bar ( .A1(abar[2]), .A2(bbar[15]), .ZN(ybar[47]);
  AND2_X1 U60 ( .A1(a[2]), .A2(b[14]), .ZN(y[46]) );
  OR2_X1 U60bar ( .A1(abar[2]), .A2(bbar[14]), .ZN(ybar[46]);
  AND2_X1 U61 ( .A1(a[2]), .A2(b[13]), .ZN(y[45]) );
  OR2_X1 U61bar ( .A1(abar[2]), .A2(bbar[13]), .ZN(ybar[45]);
  AND2_X1 U62 ( .A1(a[2]), .A2(b[12]), .ZN(y[44]) );
  OR2_X1 U62bar ( .A1(abar[2]), .A2(bbar[12]), .ZN(ybar[44]);
  AND2_X1 U63 ( .A1(a[2]), .A2(b[11]), .ZN(y[43]) );
  OR2_X1 U63bar ( .A1(abar[2]), .A2(bbar[11]), .ZN(ybar[43]);
  AND2_X1 U64 ( .A1(a[2]), .A2(b[10]), .ZN(y[42]) );
  OR2_X1 U64bar ( .A1(abar[2]), .A2(bbar[10]), .ZN(ybar[42]);
  AND2_X1 U65 ( .A1(a[2]), .A2(b[9]), .ZN(y[41]) );
  OR2_X1 U65bar ( .A1(abar[2]), .A2(bbar[9]), .ZN(ybar[41]);
  AND2_X1 U66 ( .A1(a[2]), .A2(b[8]), .ZN(y[40]) );
  OR2_X1 U66bar ( .A1(abar[2]), .A2(bbar[8]), .ZN(ybar[40]);
  AND2_X1 U67 ( .A1(b[3]), .A2(a[0]), .ZN(y[3]) );
  OR2_X1 U67bar ( .A1(bbar[3]), .A2(abar[0]), .ZN(ybar[3]);
  AND2_X1 U68 ( .A1(a[2]), .A2(b[7]), .ZN(y[39]) );
  OR2_X1 U68bar ( .A1(abar[2]), .A2(bbar[7]), .ZN(ybar[39]);
  AND2_X1 U69 ( .A1(a[2]), .A2(b[6]), .ZN(y[38]) );
  OR2_X1 U69bar ( .A1(abar[2]), .A2(bbar[6]), .ZN(ybar[38]);
  AND2_X1 U70 ( .A1(a[2]), .A2(b[5]), .ZN(y[37]) );
  OR2_X1 U70bar ( .A1(abar[2]), .A2(bbar[5]), .ZN(ybar[37]);
  AND2_X1 U71 ( .A1(a[2]), .A2(b[4]), .ZN(y[36]) );
  OR2_X1 U71bar ( .A1(abar[2]), .A2(bbar[4]), .ZN(ybar[36]);
  AND2_X1 U72 ( .A1(a[2]), .A2(b[3]), .ZN(y[35]) );
  OR2_X1 U72bar ( .A1(abar[2]), .A2(bbar[3]), .ZN(ybar[35]);
  AND2_X1 U73 ( .A1(a[2]), .A2(b[2]), .ZN(y[34]) );
  OR2_X1 U73bar ( .A1(abar[2]), .A2(bbar[2]), .ZN(ybar[34]);
  AND2_X1 U74 ( .A1(a[2]), .A2(b[1]), .ZN(y[33]) );
  OR2_X1 U74bar ( .A1(abar[2]), .A2(bbar[1]), .ZN(ybar[33]);
  AND2_X1 U75 ( .A1(a[2]), .A2(b[0]), .ZN(y[32]) );
  OR2_X1 U75bar ( .A1(abar[2]), .A2(bbar[0]), .ZN(ybar[32]);
  AND2_X1 U76 ( .A1(a[1]), .A2(b[15]), .ZN(y[31]) );
  OR2_X1 U76bar ( .A1(abar[1]), .A2(bbar[15]), .ZN(ybar[31]);
  AND2_X1 U77 ( .A1(a[1]), .A2(b[14]), .ZN(y[30]) );
  OR2_X1 U77bar ( .A1(abar[1]), .A2(bbar[14]), .ZN(ybar[30]);
  AND2_X1 U78 ( .A1(b[2]), .A2(a[0]), .ZN(y[2]) );
  OR2_X1 U78bar ( .A1(bbar[2]), .A2(abar[0]), .ZN(ybar[2]);
  AND2_X1 U79 ( .A1(a[1]), .A2(b[13]), .ZN(y[29]) );
  OR2_X1 U79bar ( .A1(abar[1]), .A2(bbar[13]), .ZN(ybar[29]);
  AND2_X1 U80 ( .A1(a[1]), .A2(b[12]), .ZN(y[28]) );
  OR2_X1 U80bar ( .A1(abar[1]), .A2(bbar[12]), .ZN(ybar[28]);
  AND2_X1 U81 ( .A1(a[1]), .A2(b[11]), .ZN(y[27]) );
  OR2_X1 U81bar ( .A1(abar[1]), .A2(bbar[11]), .ZN(ybar[27]);
  AND2_X1 U82 ( .A1(a[1]), .A2(b[10]), .ZN(y[26]) );
  OR2_X1 U82bar ( .A1(abar[1]), .A2(bbar[10]), .ZN(ybar[26]);
  AND2_X1 U83 ( .A1(a[1]), .A2(b[9]), .ZN(y[25]) );
  OR2_X1 U83bar ( .A1(abar[1]), .A2(bbar[9]), .ZN(ybar[25]);
  AND2_X1 U84 ( .A1(a[15]), .A2(b[15]), .ZN(y[255]) );
  OR2_X1 U84bar ( .A1(abar[15]), .A2(bbar[15]), .ZN(ybar[255]);
  AND2_X1 U85 ( .A1(a[15]), .A2(b[14]), .ZN(y[254]) );
  OR2_X1 U85bar ( .A1(abar[15]), .A2(bbar[14]), .ZN(ybar[254]);
  AND2_X1 U86 ( .A1(a[15]), .A2(b[13]), .ZN(y[253]) );
  OR2_X1 U86bar ( .A1(abar[15]), .A2(bbar[13]), .ZN(ybar[253]);
  AND2_X1 U87 ( .A1(a[15]), .A2(b[12]), .ZN(y[252]) );
  OR2_X1 U87bar ( .A1(abar[15]), .A2(bbar[12]), .ZN(ybar[252]);
  AND2_X1 U88 ( .A1(a[15]), .A2(b[11]), .ZN(y[251]) );
  OR2_X1 U88bar ( .A1(abar[15]), .A2(bbar[11]), .ZN(ybar[251]);
  AND2_X1 U89 ( .A1(a[15]), .A2(b[10]), .ZN(y[250]) );
  OR2_X1 U89bar ( .A1(abar[15]), .A2(bbar[10]), .ZN(ybar[250]);
  AND2_X1 U90 ( .A1(a[1]), .A2(b[8]), .ZN(y[24]) );
  OR2_X1 U90bar ( .A1(abar[1]), .A2(bbar[8]), .ZN(ybar[24]);
  AND2_X1 U91 ( .A1(a[15]), .A2(b[9]), .ZN(y[249]) );
  OR2_X1 U91bar ( .A1(abar[15]), .A2(bbar[9]), .ZN(ybar[249]);
  AND2_X1 U92 ( .A1(a[15]), .A2(b[8]), .ZN(y[248]) );
  OR2_X1 U92bar ( .A1(abar[15]), .A2(bbar[8]), .ZN(ybar[248]);
  AND2_X1 U93 ( .A1(a[15]), .A2(b[7]), .ZN(y[247]) );
  OR2_X1 U93bar ( .A1(abar[15]), .A2(bbar[7]), .ZN(ybar[247]);
  AND2_X1 U94 ( .A1(a[15]), .A2(b[6]), .ZN(y[246]) );
  OR2_X1 U94bar ( .A1(abar[15]), .A2(bbar[6]), .ZN(ybar[246]);
  AND2_X1 U95 ( .A1(a[15]), .A2(b[5]), .ZN(y[245]) );
  OR2_X1 U95bar ( .A1(abar[15]), .A2(bbar[5]), .ZN(ybar[245]);
  AND2_X1 U96 ( .A1(a[15]), .A2(b[4]), .ZN(y[244]) );
  OR2_X1 U96bar ( .A1(abar[15]), .A2(bbar[4]), .ZN(ybar[244]);
  AND2_X1 U97 ( .A1(a[15]), .A2(b[3]), .ZN(y[243]) );
  OR2_X1 U97bar ( .A1(abar[15]), .A2(bbar[3]), .ZN(ybar[243]);
  AND2_X1 U98 ( .A1(a[15]), .A2(b[2]), .ZN(y[242]) );
  OR2_X1 U98bar ( .A1(abar[15]), .A2(bbar[2]), .ZN(ybar[242]);
  AND2_X1 U99 ( .A1(a[15]), .A2(b[1]), .ZN(y[241]) );
  OR2_X1 U99bar ( .A1(abar[15]), .A2(bbar[1]), .ZN(ybar[241]);
  AND2_X1 U100 ( .A1(a[15]), .A2(b[0]), .ZN(y[240]) );
  OR2_X1 U100bar ( .A1(abar[15]), .A2(bbar[0]), .ZN(ybar[240]);
  AND2_X1 U101 ( .A1(a[1]), .A2(b[7]), .ZN(y[23]) );
  OR2_X1 U101bar ( .A1(abar[1]), .A2(bbar[7]), .ZN(ybar[23]);
  AND2_X1 U102 ( .A1(a[14]), .A2(b[15]), .ZN(y[239]) );
  OR2_X1 U102bar ( .A1(abar[14]), .A2(bbar[15]), .ZN(ybar[239]);
  AND2_X1 U103 ( .A1(a[14]), .A2(b[14]), .ZN(y[238]) );
  OR2_X1 U103bar ( .A1(abar[14]), .A2(bbar[14]), .ZN(ybar[238]);
  AND2_X1 U104 ( .A1(a[14]), .A2(b[13]), .ZN(y[237]) );
  OR2_X1 U104bar ( .A1(abar[14]), .A2(bbar[13]), .ZN(ybar[237]);
  AND2_X1 U105 ( .A1(a[14]), .A2(b[12]), .ZN(y[236]) );
  OR2_X1 U105bar ( .A1(abar[14]), .A2(bbar[12]), .ZN(ybar[236]);
  AND2_X1 U106 ( .A1(a[14]), .A2(b[11]), .ZN(y[235]) );
  OR2_X1 U106bar ( .A1(abar[14]), .A2(bbar[11]), .ZN(ybar[235]);
  AND2_X1 U107 ( .A1(a[14]), .A2(b[10]), .ZN(y[234]) );
  OR2_X1 U107bar ( .A1(abar[14]), .A2(bbar[10]), .ZN(ybar[234]);
  AND2_X1 U108 ( .A1(a[14]), .A2(b[9]), .ZN(y[233]) );
  OR2_X1 U108bar ( .A1(abar[14]), .A2(bbar[9]), .ZN(ybar[233]);
  AND2_X1 U109 ( .A1(a[14]), .A2(b[8]), .ZN(y[232]) );
  OR2_X1 U109bar ( .A1(abar[14]), .A2(bbar[8]), .ZN(ybar[232]);
  AND2_X1 U110 ( .A1(a[14]), .A2(b[7]), .ZN(y[231]) );
  OR2_X1 U110bar ( .A1(abar[14]), .A2(bbar[7]), .ZN(ybar[231]);
  AND2_X1 U111 ( .A1(a[14]), .A2(b[6]), .ZN(y[230]) );
  OR2_X1 U111bar ( .A1(abar[14]), .A2(bbar[6]), .ZN(ybar[230]);
  AND2_X1 U112 ( .A1(a[1]), .A2(b[6]), .ZN(y[22]) );
  OR2_X1 U112bar ( .A1(abar[1]), .A2(bbar[6]), .ZN(ybar[22]);
  AND2_X1 U113 ( .A1(a[14]), .A2(b[5]), .ZN(y[229]) );
  OR2_X1 U113bar ( .A1(abar[14]), .A2(bbar[5]), .ZN(ybar[229]);
  AND2_X1 U114 ( .A1(a[14]), .A2(b[4]), .ZN(y[228]) );
  OR2_X1 U114bar ( .A1(abar[14]), .A2(bbar[4]), .ZN(ybar[228]);
  AND2_X1 U115 ( .A1(a[14]), .A2(b[3]), .ZN(y[227]) );
  OR2_X1 U115bar ( .A1(abar[14]), .A2(bbar[3]), .ZN(ybar[227]);
  AND2_X1 U116 ( .A1(a[14]), .A2(b[2]), .ZN(y[226]) );
  OR2_X1 U116bar ( .A1(abar[14]), .A2(bbar[2]), .ZN(ybar[226]);
  AND2_X1 U117 ( .A1(a[14]), .A2(b[1]), .ZN(y[225]) );
  OR2_X1 U117bar ( .A1(abar[14]), .A2(bbar[1]), .ZN(ybar[225]);
  AND2_X1 U118 ( .A1(a[14]), .A2(b[0]), .ZN(y[224]) );
  OR2_X1 U118bar ( .A1(abar[14]), .A2(bbar[0]), .ZN(ybar[224]);
  AND2_X1 U119 ( .A1(a[13]), .A2(b[15]), .ZN(y[223]) );
  OR2_X1 U119bar ( .A1(abar[13]), .A2(bbar[15]), .ZN(ybar[223]);
  AND2_X1 U120 ( .A1(a[13]), .A2(b[14]), .ZN(y[222]) );
  OR2_X1 U120bar ( .A1(abar[13]), .A2(bbar[14]), .ZN(ybar[222]);
  AND2_X1 U121 ( .A1(a[13]), .A2(b[13]), .ZN(y[221]) );
  OR2_X1 U121bar ( .A1(abar[13]), .A2(bbar[13]), .ZN(ybar[221]);
  AND2_X1 U122 ( .A1(a[13]), .A2(b[12]), .ZN(y[220]) );
  OR2_X1 U122bar ( .A1(abar[13]), .A2(bbar[12]), .ZN(ybar[220]);
  AND2_X1 U123 ( .A1(a[1]), .A2(b[5]), .ZN(y[21]) );
  OR2_X1 U123bar ( .A1(abar[1]), .A2(bbar[5]), .ZN(ybar[21]);
  AND2_X1 U124 ( .A1(a[13]), .A2(b[11]), .ZN(y[219]) );
  OR2_X1 U124bar ( .A1(abar[13]), .A2(bbar[11]), .ZN(ybar[219]);
  AND2_X1 U125 ( .A1(a[13]), .A2(b[10]), .ZN(y[218]) );
  OR2_X1 U125bar ( .A1(abar[13]), .A2(bbar[10]), .ZN(ybar[218]);
  AND2_X1 U126 ( .A1(a[13]), .A2(b[9]), .ZN(y[217]) );
  OR2_X1 U126bar ( .A1(abar[13]), .A2(bbar[9]), .ZN(ybar[217]);
  AND2_X1 U127 ( .A1(a[13]), .A2(b[8]), .ZN(y[216]) );
  OR2_X1 U127bar ( .A1(abar[13]), .A2(bbar[8]), .ZN(ybar[216]);
  AND2_X1 U128 ( .A1(a[13]), .A2(b[7]), .ZN(y[215]) );
  OR2_X1 U128bar ( .A1(abar[13]), .A2(bbar[7]), .ZN(ybar[215]);
  AND2_X1 U129 ( .A1(a[13]), .A2(b[6]), .ZN(y[214]) );
  OR2_X1 U129bar ( .A1(abar[13]), .A2(bbar[6]), .ZN(ybar[214]);
  AND2_X1 U130 ( .A1(a[13]), .A2(b[5]), .ZN(y[213]) );
  OR2_X1 U130bar ( .A1(abar[13]), .A2(bbar[5]), .ZN(ybar[213]);
  AND2_X1 U131 ( .A1(a[13]), .A2(b[4]), .ZN(y[212]) );
  OR2_X1 U131bar ( .A1(abar[13]), .A2(bbar[4]), .ZN(ybar[212]);
  AND2_X1 U132 ( .A1(a[13]), .A2(b[3]), .ZN(y[211]) );
  OR2_X1 U132bar ( .A1(abar[13]), .A2(bbar[3]), .ZN(ybar[211]);
  AND2_X1 U133 ( .A1(a[13]), .A2(b[2]), .ZN(y[210]) );
  OR2_X1 U133bar ( .A1(abar[13]), .A2(bbar[2]), .ZN(ybar[210]);
  AND2_X1 U134 ( .A1(a[1]), .A2(b[4]), .ZN(y[20]) );
  OR2_X1 U134bar ( .A1(abar[1]), .A2(bbar[4]), .ZN(ybar[20]);
  AND2_X1 U135 ( .A1(a[13]), .A2(b[1]), .ZN(y[209]) );
  OR2_X1 U135bar ( .A1(abar[13]), .A2(bbar[1]), .ZN(ybar[209]);
  AND2_X1 U136 ( .A1(a[13]), .A2(b[0]), .ZN(y[208]) );
  OR2_X1 U136bar ( .A1(abar[13]), .A2(bbar[0]), .ZN(ybar[208]);
  AND2_X1 U137 ( .A1(a[12]), .A2(b[15]), .ZN(y[207]) );
  OR2_X1 U137bar ( .A1(abar[12]), .A2(bbar[15]), .ZN(ybar[207]);
  AND2_X1 U138 ( .A1(a[12]), .A2(b[14]), .ZN(y[206]) );
  OR2_X1 U138bar ( .A1(abar[12]), .A2(bbar[14]), .ZN(ybar[206]);
  AND2_X1 U139 ( .A1(a[12]), .A2(b[13]), .ZN(y[205]) );
  OR2_X1 U139bar ( .A1(abar[12]), .A2(bbar[13]), .ZN(ybar[205]);
  AND2_X1 U140 ( .A1(a[12]), .A2(b[12]), .ZN(y[204]) );
  OR2_X1 U140bar ( .A1(abar[12]), .A2(bbar[12]), .ZN(ybar[204]);
  AND2_X1 U141 ( .A1(a[12]), .A2(b[11]), .ZN(y[203]) );
  OR2_X1 U141bar ( .A1(abar[12]), .A2(bbar[11]), .ZN(ybar[203]);
  AND2_X1 U142 ( .A1(a[12]), .A2(b[10]), .ZN(y[202]) );
  OR2_X1 U142bar ( .A1(abar[12]), .A2(bbar[10]), .ZN(ybar[202]);
  AND2_X1 U143 ( .A1(a[12]), .A2(b[9]), .ZN(y[201]) );
  OR2_X1 U143bar ( .A1(abar[12]), .A2(bbar[9]), .ZN(ybar[201]);
  AND2_X1 U144 ( .A1(a[12]), .A2(b[8]), .ZN(y[200]) );
  OR2_X1 U144bar ( .A1(abar[12]), .A2(bbar[8]), .ZN(ybar[200]);
  AND2_X1 U145 ( .A1(b[1]), .A2(a[0]), .ZN(y[1]) );
  OR2_X1 U145bar ( .A1(bbar[1]), .A2(abar[0]), .ZN(ybar[1]);
  AND2_X1 U146 ( .A1(a[1]), .A2(b[3]), .ZN(y[19]) );
  OR2_X1 U146bar ( .A1(abar[1]), .A2(bbar[3]), .ZN(ybar[19]);
  AND2_X1 U147 ( .A1(a[12]), .A2(b[7]), .ZN(y[199]) );
  OR2_X1 U147bar ( .A1(abar[12]), .A2(bbar[7]), .ZN(ybar[199]);
  AND2_X1 U148 ( .A1(a[12]), .A2(b[6]), .ZN(y[198]) );
  OR2_X1 U148bar ( .A1(abar[12]), .A2(bbar[6]), .ZN(ybar[198]);
  AND2_X1 U149 ( .A1(a[12]), .A2(b[5]), .ZN(y[197]) );
  OR2_X1 U149bar ( .A1(abar[12]), .A2(bbar[5]), .ZN(ybar[197]);
  AND2_X1 U150 ( .A1(a[12]), .A2(b[4]), .ZN(y[196]) );
  OR2_X1 U150bar ( .A1(abar[12]), .A2(bbar[4]), .ZN(ybar[196]);
  AND2_X1 U151 ( .A1(a[12]), .A2(b[3]), .ZN(y[195]) );
  OR2_X1 U151bar ( .A1(abar[12]), .A2(bbar[3]), .ZN(ybar[195]);
  AND2_X1 U152 ( .A1(a[12]), .A2(b[2]), .ZN(y[194]) );
  OR2_X1 U152bar ( .A1(abar[12]), .A2(bbar[2]), .ZN(ybar[194]);
  AND2_X1 U153 ( .A1(a[12]), .A2(b[1]), .ZN(y[193]) );
  OR2_X1 U153bar ( .A1(abar[12]), .A2(bbar[1]), .ZN(ybar[193]);
  AND2_X1 U154 ( .A1(a[12]), .A2(b[0]), .ZN(y[192]) );
  OR2_X1 U154bar ( .A1(abar[12]), .A2(bbar[0]), .ZN(ybar[192]);
  AND2_X1 U155 ( .A1(a[11]), .A2(b[15]), .ZN(y[191]) );
  OR2_X1 U155bar ( .A1(abar[11]), .A2(bbar[15]), .ZN(ybar[191]);
  AND2_X1 U156 ( .A1(a[11]), .A2(b[14]), .ZN(y[190]) );
  OR2_X1 U156bar ( .A1(abar[11]), .A2(bbar[14]), .ZN(ybar[190]);
  AND2_X1 U157 ( .A1(a[1]), .A2(b[2]), .ZN(y[18]) );
  OR2_X1 U157bar ( .A1(abar[1]), .A2(bbar[2]), .ZN(ybar[18]);
  AND2_X1 U158 ( .A1(a[11]), .A2(b[13]), .ZN(y[189]) );
  OR2_X1 U158bar ( .A1(abar[11]), .A2(bbar[13]), .ZN(ybar[189]);
  AND2_X1 U159 ( .A1(a[11]), .A2(b[12]), .ZN(y[188]) );
  OR2_X1 U159bar ( .A1(abar[11]), .A2(bbar[12]), .ZN(ybar[188]);
  AND2_X1 U160 ( .A1(a[11]), .A2(b[11]), .ZN(y[187]) );
  OR2_X1 U160bar ( .A1(abar[11]), .A2(bbar[11]), .ZN(ybar[187]);
  AND2_X1 U161 ( .A1(a[11]), .A2(b[10]), .ZN(y[186]) );
  OR2_X1 U161bar ( .A1(abar[11]), .A2(bbar[10]), .ZN(ybar[186]);
  AND2_X1 U162 ( .A1(a[11]), .A2(b[9]), .ZN(y[185]) );
  OR2_X1 U162bar ( .A1(abar[11]), .A2(bbar[9]), .ZN(ybar[185]);
  AND2_X1 U163 ( .A1(a[11]), .A2(b[8]), .ZN(y[184]) );
  OR2_X1 U163bar ( .A1(abar[11]), .A2(bbar[8]), .ZN(ybar[184]);
  AND2_X1 U164 ( .A1(a[11]), .A2(b[7]), .ZN(y[183]) );
  OR2_X1 U164bar ( .A1(abar[11]), .A2(bbar[7]), .ZN(ybar[183]);
  AND2_X1 U165 ( .A1(a[11]), .A2(b[6]), .ZN(y[182]) );
  OR2_X1 U165bar ( .A1(abar[11]), .A2(bbar[6]), .ZN(ybar[182]);
  AND2_X1 U166 ( .A1(a[11]), .A2(b[5]), .ZN(y[181]) );
  OR2_X1 U166bar ( .A1(abar[11]), .A2(bbar[5]), .ZN(ybar[181]);
  AND2_X1 U167 ( .A1(a[11]), .A2(b[4]), .ZN(y[180]) );
  OR2_X1 U167bar ( .A1(abar[11]), .A2(bbar[4]), .ZN(ybar[180]);
  AND2_X1 U168 ( .A1(a[1]), .A2(b[1]), .ZN(y[17]) );
  OR2_X1 U168bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[17]);
  AND2_X1 U169 ( .A1(a[11]), .A2(b[3]), .ZN(y[179]) );
  OR2_X1 U169bar ( .A1(abar[11]), .A2(bbar[3]), .ZN(ybar[179]);
  AND2_X1 U170 ( .A1(a[11]), .A2(b[2]), .ZN(y[178]) );
  OR2_X1 U170bar ( .A1(abar[11]), .A2(bbar[2]), .ZN(ybar[178]);
  AND2_X1 U171 ( .A1(a[11]), .A2(b[1]), .ZN(y[177]) );
  OR2_X1 U171bar ( .A1(abar[11]), .A2(bbar[1]), .ZN(ybar[177]);
  AND2_X1 U172 ( .A1(a[11]), .A2(b[0]), .ZN(y[176]) );
  OR2_X1 U172bar ( .A1(abar[11]), .A2(bbar[0]), .ZN(ybar[176]);
  AND2_X1 U173 ( .A1(a[10]), .A2(b[15]), .ZN(y[175]) );
  OR2_X1 U173bar ( .A1(abar[10]), .A2(bbar[15]), .ZN(ybar[175]);
  AND2_X1 U174 ( .A1(a[10]), .A2(b[14]), .ZN(y[174]) );
  OR2_X1 U174bar ( .A1(abar[10]), .A2(bbar[14]), .ZN(ybar[174]);
  AND2_X1 U175 ( .A1(a[10]), .A2(b[13]), .ZN(y[173]) );
  OR2_X1 U175bar ( .A1(abar[10]), .A2(bbar[13]), .ZN(ybar[173]);
  AND2_X1 U176 ( .A1(a[10]), .A2(b[12]), .ZN(y[172]) );
  OR2_X1 U176bar ( .A1(abar[10]), .A2(bbar[12]), .ZN(ybar[172]);
  AND2_X1 U177 ( .A1(a[10]), .A2(b[11]), .ZN(y[171]) );
  OR2_X1 U177bar ( .A1(abar[10]), .A2(bbar[11]), .ZN(ybar[171]);
  AND2_X1 U178 ( .A1(a[10]), .A2(b[10]), .ZN(y[170]) );
  OR2_X1 U178bar ( .A1(abar[10]), .A2(bbar[10]), .ZN(ybar[170]);
  AND2_X1 U179 ( .A1(a[1]), .A2(b[0]), .ZN(y[16]) );
  OR2_X1 U179bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[16]);
  AND2_X1 U180 ( .A1(a[10]), .A2(b[9]), .ZN(y[169]) );
  OR2_X1 U180bar ( .A1(abar[10]), .A2(bbar[9]), .ZN(ybar[169]);
  AND2_X1 U181 ( .A1(a[10]), .A2(b[8]), .ZN(y[168]) );
  OR2_X1 U181bar ( .A1(abar[10]), .A2(bbar[8]), .ZN(ybar[168]);
  AND2_X1 U182 ( .A1(a[10]), .A2(b[7]), .ZN(y[167]) );
  OR2_X1 U182bar ( .A1(abar[10]), .A2(bbar[7]), .ZN(ybar[167]);
  AND2_X1 U183 ( .A1(a[10]), .A2(b[6]), .ZN(y[166]) );
  OR2_X1 U183bar ( .A1(abar[10]), .A2(bbar[6]), .ZN(ybar[166]);
  AND2_X1 U184 ( .A1(a[10]), .A2(b[5]), .ZN(y[165]) );
  OR2_X1 U184bar ( .A1(abar[10]), .A2(bbar[5]), .ZN(ybar[165]);
  AND2_X1 U185 ( .A1(a[10]), .A2(b[4]), .ZN(y[164]) );
  OR2_X1 U185bar ( .A1(abar[10]), .A2(bbar[4]), .ZN(ybar[164]);
  AND2_X1 U186 ( .A1(a[10]), .A2(b[3]), .ZN(y[163]) );
  OR2_X1 U186bar ( .A1(abar[10]), .A2(bbar[3]), .ZN(ybar[163]);
  AND2_X1 U187 ( .A1(a[10]), .A2(b[2]), .ZN(y[162]) );
  OR2_X1 U187bar ( .A1(abar[10]), .A2(bbar[2]), .ZN(ybar[162]);
  AND2_X1 U188 ( .A1(a[10]), .A2(b[1]), .ZN(y[161]) );
  OR2_X1 U188bar ( .A1(abar[10]), .A2(bbar[1]), .ZN(ybar[161]);
  AND2_X1 U189 ( .A1(a[10]), .A2(b[0]), .ZN(y[160]) );
  OR2_X1 U189bar ( .A1(abar[10]), .A2(bbar[0]), .ZN(ybar[160]);
  AND2_X1 U190 ( .A1(b[15]), .A2(a[0]), .ZN(y[15]) );
  OR2_X1 U190bar ( .A1(bbar[15]), .A2(abar[0]), .ZN(ybar[15]);
  AND2_X1 U191 ( .A1(a[9]), .A2(b[15]), .ZN(y[159]) );
  OR2_X1 U191bar ( .A1(abar[9]), .A2(bbar[15]), .ZN(ybar[159]);
  AND2_X1 U192 ( .A1(a[9]), .A2(b[14]), .ZN(y[158]) );
  OR2_X1 U192bar ( .A1(abar[9]), .A2(bbar[14]), .ZN(ybar[158]);
  AND2_X1 U193 ( .A1(a[9]), .A2(b[13]), .ZN(y[157]) );
  OR2_X1 U193bar ( .A1(abar[9]), .A2(bbar[13]), .ZN(ybar[157]);
  AND2_X1 U194 ( .A1(a[9]), .A2(b[12]), .ZN(y[156]) );
  OR2_X1 U194bar ( .A1(abar[9]), .A2(bbar[12]), .ZN(ybar[156]);
  AND2_X1 U195 ( .A1(a[9]), .A2(b[11]), .ZN(y[155]) );
  OR2_X1 U195bar ( .A1(abar[9]), .A2(bbar[11]), .ZN(ybar[155]);
  AND2_X1 U196 ( .A1(a[9]), .A2(b[10]), .ZN(y[154]) );
  OR2_X1 U196bar ( .A1(abar[9]), .A2(bbar[10]), .ZN(ybar[154]);
  AND2_X1 U197 ( .A1(a[9]), .A2(b[9]), .ZN(y[153]) );
  OR2_X1 U197bar ( .A1(abar[9]), .A2(bbar[9]), .ZN(ybar[153]);
  AND2_X1 U198 ( .A1(a[9]), .A2(b[8]), .ZN(y[152]) );
  OR2_X1 U198bar ( .A1(abar[9]), .A2(bbar[8]), .ZN(ybar[152]);
  AND2_X1 U199 ( .A1(a[9]), .A2(b[7]), .ZN(y[151]) );
  OR2_X1 U199bar ( .A1(abar[9]), .A2(bbar[7]), .ZN(ybar[151]);
  AND2_X1 U200 ( .A1(a[9]), .A2(b[6]), .ZN(y[150]) );
  OR2_X1 U200bar ( .A1(abar[9]), .A2(bbar[6]), .ZN(ybar[150]);
  AND2_X1 U201 ( .A1(b[14]), .A2(a[0]), .ZN(y[14]) );
  OR2_X1 U201bar ( .A1(bbar[14]), .A2(abar[0]), .ZN(ybar[14]);
  AND2_X1 U202 ( .A1(a[9]), .A2(b[5]), .ZN(y[149]) );
  OR2_X1 U202bar ( .A1(abar[9]), .A2(bbar[5]), .ZN(ybar[149]);
  AND2_X1 U203 ( .A1(a[9]), .A2(b[4]), .ZN(y[148]) );
  OR2_X1 U203bar ( .A1(abar[9]), .A2(bbar[4]), .ZN(ybar[148]);
  AND2_X1 U204 ( .A1(a[9]), .A2(b[3]), .ZN(y[147]) );
  OR2_X1 U204bar ( .A1(abar[9]), .A2(bbar[3]), .ZN(ybar[147]);
  AND2_X1 U205 ( .A1(a[9]), .A2(b[2]), .ZN(y[146]) );
  OR2_X1 U205bar ( .A1(abar[9]), .A2(bbar[2]), .ZN(ybar[146]);
  AND2_X1 U206 ( .A1(a[9]), .A2(b[1]), .ZN(y[145]) );
  OR2_X1 U206bar ( .A1(abar[9]), .A2(bbar[1]), .ZN(ybar[145]);
  AND2_X1 U207 ( .A1(a[9]), .A2(b[0]), .ZN(y[144]) );
  OR2_X1 U207bar ( .A1(abar[9]), .A2(bbar[0]), .ZN(ybar[144]);
  AND2_X1 U208 ( .A1(a[8]), .A2(b[15]), .ZN(y[143]) );
  OR2_X1 U208bar ( .A1(abar[8]), .A2(bbar[15]), .ZN(ybar[143]);
  AND2_X1 U209 ( .A1(a[8]), .A2(b[14]), .ZN(y[142]) );
  OR2_X1 U209bar ( .A1(abar[8]), .A2(bbar[14]), .ZN(ybar[142]);
  AND2_X1 U210 ( .A1(a[8]), .A2(b[13]), .ZN(y[141]) );
  OR2_X1 U210bar ( .A1(abar[8]), .A2(bbar[13]), .ZN(ybar[141]);
  AND2_X1 U211 ( .A1(a[8]), .A2(b[12]), .ZN(y[140]) );
  OR2_X1 U211bar ( .A1(abar[8]), .A2(bbar[12]), .ZN(ybar[140]);
  AND2_X1 U212 ( .A1(b[13]), .A2(a[0]), .ZN(y[13]) );
  OR2_X1 U212bar ( .A1(bbar[13]), .A2(abar[0]), .ZN(ybar[13]);
  AND2_X1 U213 ( .A1(a[8]), .A2(b[11]), .ZN(y[139]) );
  OR2_X1 U213bar ( .A1(abar[8]), .A2(bbar[11]), .ZN(ybar[139]);
  AND2_X1 U214 ( .A1(a[8]), .A2(b[10]), .ZN(y[138]) );
  OR2_X1 U214bar ( .A1(abar[8]), .A2(bbar[10]), .ZN(ybar[138]);
  AND2_X1 U215 ( .A1(a[8]), .A2(b[9]), .ZN(y[137]) );
  OR2_X1 U215bar ( .A1(abar[8]), .A2(bbar[9]), .ZN(ybar[137]);
  AND2_X1 U216 ( .A1(a[8]), .A2(b[8]), .ZN(y[136]) );
  OR2_X1 U216bar ( .A1(abar[8]), .A2(bbar[8]), .ZN(ybar[136]);
  AND2_X1 U217 ( .A1(a[8]), .A2(b[7]), .ZN(y[135]) );
  OR2_X1 U217bar ( .A1(abar[8]), .A2(bbar[7]), .ZN(ybar[135]);
  AND2_X1 U218 ( .A1(a[8]), .A2(b[6]), .ZN(y[134]) );
  OR2_X1 U218bar ( .A1(abar[8]), .A2(bbar[6]), .ZN(ybar[134]);
  AND2_X1 U219 ( .A1(a[8]), .A2(b[5]), .ZN(y[133]) );
  OR2_X1 U219bar ( .A1(abar[8]), .A2(bbar[5]), .ZN(ybar[133]);
  AND2_X1 U220 ( .A1(a[8]), .A2(b[4]), .ZN(y[132]) );
  OR2_X1 U220bar ( .A1(abar[8]), .A2(bbar[4]), .ZN(ybar[132]);
  AND2_X1 U221 ( .A1(a[8]), .A2(b[3]), .ZN(y[131]) );
  OR2_X1 U221bar ( .A1(abar[8]), .A2(bbar[3]), .ZN(ybar[131]);
  AND2_X1 U222 ( .A1(a[8]), .A2(b[2]), .ZN(y[130]) );
  OR2_X1 U222bar ( .A1(abar[8]), .A2(bbar[2]), .ZN(ybar[130]);
  AND2_X1 U223 ( .A1(b[12]), .A2(a[0]), .ZN(y[12]) );
  OR2_X1 U223bar ( .A1(bbar[12]), .A2(abar[0]), .ZN(ybar[12]);
  AND2_X1 U224 ( .A1(a[8]), .A2(b[1]), .ZN(y[129]) );
  OR2_X1 U224bar ( .A1(abar[8]), .A2(bbar[1]), .ZN(ybar[129]);
  AND2_X1 U225 ( .A1(a[8]), .A2(b[0]), .ZN(y[128]) );
  OR2_X1 U225bar ( .A1(abar[8]), .A2(bbar[0]), .ZN(ybar[128]);
  AND2_X1 U226 ( .A1(a[7]), .A2(b[15]), .ZN(y[127]) );
  OR2_X1 U226bar ( .A1(abar[7]), .A2(bbar[15]), .ZN(ybar[127]);
  AND2_X1 U227 ( .A1(a[7]), .A2(b[14]), .ZN(y[126]) );
  OR2_X1 U227bar ( .A1(abar[7]), .A2(bbar[14]), .ZN(ybar[126]);
  AND2_X1 U228 ( .A1(a[7]), .A2(b[13]), .ZN(y[125]) );
  OR2_X1 U228bar ( .A1(abar[7]), .A2(bbar[13]), .ZN(ybar[125]);
  AND2_X1 U229 ( .A1(a[7]), .A2(b[12]), .ZN(y[124]) );
  OR2_X1 U229bar ( .A1(abar[7]), .A2(bbar[12]), .ZN(ybar[124]);
  AND2_X1 U230 ( .A1(a[7]), .A2(b[11]), .ZN(y[123]) );
  OR2_X1 U230bar ( .A1(abar[7]), .A2(bbar[11]), .ZN(ybar[123]);
  AND2_X1 U231 ( .A1(a[7]), .A2(b[10]), .ZN(y[122]) );
  OR2_X1 U231bar ( .A1(abar[7]), .A2(bbar[10]), .ZN(ybar[122]);
  AND2_X1 U232 ( .A1(a[7]), .A2(b[9]), .ZN(y[121]) );
  OR2_X1 U232bar ( .A1(abar[7]), .A2(bbar[9]), .ZN(ybar[121]);
  AND2_X1 U233 ( .A1(a[7]), .A2(b[8]), .ZN(y[120]) );
  OR2_X1 U233bar ( .A1(abar[7]), .A2(bbar[8]), .ZN(ybar[120]);
  AND2_X1 U234 ( .A1(b[11]), .A2(a[0]), .ZN(y[11]) );
  OR2_X1 U234bar ( .A1(bbar[11]), .A2(abar[0]), .ZN(ybar[11]);
  AND2_X1 U235 ( .A1(a[7]), .A2(b[7]), .ZN(y[119]) );
  OR2_X1 U235bar ( .A1(abar[7]), .A2(bbar[7]), .ZN(ybar[119]);
  AND2_X1 U236 ( .A1(a[7]), .A2(b[6]), .ZN(y[118]) );
  OR2_X1 U236bar ( .A1(abar[7]), .A2(bbar[6]), .ZN(ybar[118]);
  AND2_X1 U237 ( .A1(a[7]), .A2(b[5]), .ZN(y[117]) );
  OR2_X1 U237bar ( .A1(abar[7]), .A2(bbar[5]), .ZN(ybar[117]);
  AND2_X1 U238 ( .A1(a[7]), .A2(b[4]), .ZN(y[116]) );
  OR2_X1 U238bar ( .A1(abar[7]), .A2(bbar[4]), .ZN(ybar[116]);
  AND2_X1 U239 ( .A1(a[7]), .A2(b[3]), .ZN(y[115]) );
  OR2_X1 U239bar ( .A1(abar[7]), .A2(bbar[3]), .ZN(ybar[115]);
  AND2_X1 U240 ( .A1(a[7]), .A2(b[2]), .ZN(y[114]) );
  OR2_X1 U240bar ( .A1(abar[7]), .A2(bbar[2]), .ZN(ybar[114]);
  AND2_X1 U241 ( .A1(a[7]), .A2(b[1]), .ZN(y[113]) );
  OR2_X1 U241bar ( .A1(abar[7]), .A2(bbar[1]), .ZN(ybar[113]);
  AND2_X1 U242 ( .A1(a[7]), .A2(b[0]), .ZN(y[112]) );
  OR2_X1 U242bar ( .A1(abar[7]), .A2(bbar[0]), .ZN(ybar[112]);
  AND2_X1 U243 ( .A1(b[15]), .A2(a[6]), .ZN(y[111]) );
  OR2_X1 U243bar ( .A1(bbar[15]), .A2(abar[6]), .ZN(ybar[111]);
  AND2_X1 U244 ( .A1(b[14]), .A2(a[6]), .ZN(y[110]) );
  OR2_X1 U244bar ( .A1(bbar[14]), .A2(abar[6]), .ZN(ybar[110]);
  AND2_X1 U245 ( .A1(b[10]), .A2(a[0]), .ZN(y[10]) );
  OR2_X1 U245bar ( .A1(bbar[10]), .A2(abar[0]), .ZN(ybar[10]);
  AND2_X1 U246 ( .A1(b[13]), .A2(a[6]), .ZN(y[109]) );
  OR2_X1 U246bar ( .A1(bbar[13]), .A2(abar[6]), .ZN(ybar[109]);
  AND2_X1 U247 ( .A1(b[12]), .A2(a[6]), .ZN(y[108]) );
  OR2_X1 U247bar ( .A1(bbar[12]), .A2(abar[6]), .ZN(ybar[108]);
  AND2_X1 U248 ( .A1(b[11]), .A2(a[6]), .ZN(y[107]) );
  OR2_X1 U248bar ( .A1(bbar[11]), .A2(abar[6]), .ZN(ybar[107]);
  AND2_X1 U249 ( .A1(b[10]), .A2(a[6]), .ZN(y[106]) );
  OR2_X1 U249bar ( .A1(bbar[10]), .A2(abar[6]), .ZN(ybar[106]);
  AND2_X1 U250 ( .A1(a[6]), .A2(b[9]), .ZN(y[105]) );
  OR2_X1 U250bar ( .A1(abar[6]), .A2(bbar[9]), .ZN(ybar[105]);
  AND2_X1 U251 ( .A1(b[8]), .A2(a[6]), .ZN(y[104]) );
  OR2_X1 U251bar ( .A1(bbar[8]), .A2(abar[6]), .ZN(ybar[104]);
  AND2_X1 U252 ( .A1(b[7]), .A2(a[6]), .ZN(y[103]) );
  OR2_X1 U252bar ( .A1(bbar[7]), .A2(abar[6]), .ZN(ybar[103]);
  AND2_X1 U253 ( .A1(b[6]), .A2(a[6]), .ZN(y[102]) );
  OR2_X1 U253bar ( .A1(bbar[6]), .A2(abar[6]), .ZN(ybar[102]);
  AND2_X1 U254 ( .A1(b[5]), .A2(a[6]), .ZN(y[101]) );
  OR2_X1 U254bar ( .A1(bbar[5]), .A2(abar[6]), .ZN(ybar[101]);
  AND2_X1 U255 ( .A1(b[4]), .A2(a[6]), .ZN(y[100]) );
  OR2_X1 U255bar ( .A1(bbar[4]), .A2(abar[6]), .ZN(ybar[100]);
  AND2_X1 U256 ( .A1(b[0]), .A2(a[0]), .ZN(y[0]) );
  OR2_X1 U256bar ( .A1(bbar[0]), .A2(abar[0]), .ZN(ybar[0]);
endmodule




module decode_10 ( in, out );
  input [7:0] in;
  //input_done

  output [255:0] out;
  //output_done

  wire   [15:0] level1;
  wire   [31:0] level2;
  //wire_done

  CD2_40 cd_l1_1 ( .a(in[1]), .b(in[0]), .y(level1[3:0]) );
  CD2_39 cd_l1_2 ( .a(in[3]), .b(in[2]), .y(level1[7:4]) );
  CD2_38 cd_l1_3 ( .a(in[5]), .b(in[4]), .y(level1[11:8]) );
  CD2_37 cd_l1_4 ( .a(in[7]), .b(in[6]), .y(level1[15:12]) );
  CD4_20 cd_l2_1 ( .a(level1[7:4]), .b(level1[3:0]), .y(level2[15:0]) );
  CD4_19 cd_l2_2 ( .a(level1[15:12]), .b(level1[11:8]), .y(level2[31:16]) );
  CD16_10 cd_l3 ( .a(level2[31:16]), .b(level2[15:0]), .y(out) );
endmodule


module encode_10 ( in, out );
  input [255:0] in;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
  assign inbar[8] = ~in[8];
  assign inbar[9] = ~in[9];
  assign inbar[10] = ~in[10];
  assign inbar[11] = ~in[11];
  assign inbar[12] = ~in[12];
  assign inbar[13] = ~in[13];
  assign inbar[14] = ~in[14];
  assign inbar[15] = ~in[15];
  assign inbar[16] = ~in[16];
  assign inbar[17] = ~in[17];
  assign inbar[18] = ~in[18];
  assign inbar[19] = ~in[19];
  assign inbar[20] = ~in[20];
  assign inbar[21] = ~in[21];
  assign inbar[22] = ~in[22];
  assign inbar[23] = ~in[23];
  assign inbar[24] = ~in[24];
  assign inbar[25] = ~in[25];
  assign inbar[26] = ~in[26];
  assign inbar[27] = ~in[27];
  assign inbar[28] = ~in[28];
  assign inbar[29] = ~in[29];
  assign inbar[30] = ~in[30];
  assign inbar[31] = ~in[31];
  assign inbar[32] = ~in[32];
  assign inbar[33] = ~in[33];
  assign inbar[34] = ~in[34];
  assign inbar[35] = ~in[35];
  assign inbar[36] = ~in[36];
  assign inbar[37] = ~in[37];
  assign inbar[38] = ~in[38];
  assign inbar[39] = ~in[39];
  assign inbar[40] = ~in[40];
  assign inbar[41] = ~in[41];
  assign inbar[42] = ~in[42];
  assign inbar[43] = ~in[43];
  assign inbar[44] = ~in[44];
  assign inbar[45] = ~in[45];
  assign inbar[46] = ~in[46];
  assign inbar[47] = ~in[47];
  assign inbar[48] = ~in[48];
  assign inbar[49] = ~in[49];
  assign inbar[50] = ~in[50];
  assign inbar[51] = ~in[51];
  assign inbar[52] = ~in[52];
  assign inbar[53] = ~in[53];
  assign inbar[54] = ~in[54];
  assign inbar[55] = ~in[55];
  assign inbar[56] = ~in[56];
  assign inbar[57] = ~in[57];
  assign inbar[58] = ~in[58];
  assign inbar[59] = ~in[59];
  assign inbar[60] = ~in[60];
  assign inbar[61] = ~in[61];
  assign inbar[62] = ~in[62];
  assign inbar[63] = ~in[63];
  assign inbar[64] = ~in[64];
  assign inbar[65] = ~in[65];
  assign inbar[66] = ~in[66];
  assign inbar[67] = ~in[67];
  assign inbar[68] = ~in[68];
  assign inbar[69] = ~in[69];
  assign inbar[70] = ~in[70];
  assign inbar[71] = ~in[71];
  assign inbar[72] = ~in[72];
  assign inbar[73] = ~in[73];
  assign inbar[74] = ~in[74];
  assign inbar[75] = ~in[75];
  assign inbar[76] = ~in[76];
  assign inbar[77] = ~in[77];
  assign inbar[78] = ~in[78];
  assign inbar[79] = ~in[79];
  assign inbar[80] = ~in[80];
  assign inbar[81] = ~in[81];
  assign inbar[82] = ~in[82];
  assign inbar[83] = ~in[83];
  assign inbar[84] = ~in[84];
  assign inbar[85] = ~in[85];
  assign inbar[86] = ~in[86];
  assign inbar[87] = ~in[87];
  assign inbar[88] = ~in[88];
  assign inbar[89] = ~in[89];
  assign inbar[90] = ~in[90];
  assign inbar[91] = ~in[91];
  assign inbar[92] = ~in[92];
  assign inbar[93] = ~in[93];
  assign inbar[94] = ~in[94];
  assign inbar[95] = ~in[95];
  assign inbar[96] = ~in[96];
  assign inbar[97] = ~in[97];
  assign inbar[98] = ~in[98];
  assign inbar[99] = ~in[99];
  assign inbar[100] = ~in[100];
  assign inbar[101] = ~in[101];
  assign inbar[102] = ~in[102];
  assign inbar[103] = ~in[103];
  assign inbar[104] = ~in[104];
  assign inbar[105] = ~in[105];
  assign inbar[106] = ~in[106];
  assign inbar[107] = ~in[107];
  assign inbar[108] = ~in[108];
  assign inbar[109] = ~in[109];
  assign inbar[110] = ~in[110];
  assign inbar[111] = ~in[111];
  assign inbar[112] = ~in[112];
  assign inbar[113] = ~in[113];
  assign inbar[114] = ~in[114];
  assign inbar[115] = ~in[115];
  assign inbar[116] = ~in[116];
  assign inbar[117] = ~in[117];
  assign inbar[118] = ~in[118];
  assign inbar[119] = ~in[119];
  assign inbar[120] = ~in[120];
  assign inbar[121] = ~in[121];
  assign inbar[122] = ~in[122];
  assign inbar[123] = ~in[123];
  assign inbar[124] = ~in[124];
  assign inbar[125] = ~in[125];
  assign inbar[126] = ~in[126];
  assign inbar[127] = ~in[127];
  assign inbar[128] = ~in[128];
  assign inbar[129] = ~in[129];
  assign inbar[130] = ~in[130];
  assign inbar[131] = ~in[131];
  assign inbar[132] = ~in[132];
  assign inbar[133] = ~in[133];
  assign inbar[134] = ~in[134];
  assign inbar[135] = ~in[135];
  assign inbar[136] = ~in[136];
  assign inbar[137] = ~in[137];
  assign inbar[138] = ~in[138];
  assign inbar[139] = ~in[139];
  assign inbar[140] = ~in[140];
  assign inbar[141] = ~in[141];
  assign inbar[142] = ~in[142];
  assign inbar[143] = ~in[143];
  assign inbar[144] = ~in[144];
  assign inbar[145] = ~in[145];
  assign inbar[146] = ~in[146];
  assign inbar[147] = ~in[147];
  assign inbar[148] = ~in[148];
  assign inbar[149] = ~in[149];
  assign inbar[150] = ~in[150];
  assign inbar[151] = ~in[151];
  assign inbar[152] = ~in[152];
  assign inbar[153] = ~in[153];
  assign inbar[154] = ~in[154];
  assign inbar[155] = ~in[155];
  assign inbar[156] = ~in[156];
  assign inbar[157] = ~in[157];
  assign inbar[158] = ~in[158];
  assign inbar[159] = ~in[159];
  assign inbar[160] = ~in[160];
  assign inbar[161] = ~in[161];
  assign inbar[162] = ~in[162];
  assign inbar[163] = ~in[163];
  assign inbar[164] = ~in[164];
  assign inbar[165] = ~in[165];
  assign inbar[166] = ~in[166];
  assign inbar[167] = ~in[167];
  assign inbar[168] = ~in[168];
  assign inbar[169] = ~in[169];
  assign inbar[170] = ~in[170];
  assign inbar[171] = ~in[171];
  assign inbar[172] = ~in[172];
  assign inbar[173] = ~in[173];
  assign inbar[174] = ~in[174];
  assign inbar[175] = ~in[175];
  assign inbar[176] = ~in[176];
  assign inbar[177] = ~in[177];
  assign inbar[178] = ~in[178];
  assign inbar[179] = ~in[179];
  assign inbar[180] = ~in[180];
  assign inbar[181] = ~in[181];
  assign inbar[182] = ~in[182];
  assign inbar[183] = ~in[183];
  assign inbar[184] = ~in[184];
  assign inbar[185] = ~in[185];
  assign inbar[186] = ~in[186];
  assign inbar[187] = ~in[187];
  assign inbar[188] = ~in[188];
  assign inbar[189] = ~in[189];
  assign inbar[190] = ~in[190];
  assign inbar[191] = ~in[191];
  assign inbar[192] = ~in[192];
  assign inbar[193] = ~in[193];
  assign inbar[194] = ~in[194];
  assign inbar[195] = ~in[195];
  assign inbar[196] = ~in[196];
  assign inbar[197] = ~in[197];
  assign inbar[198] = ~in[198];
  assign inbar[199] = ~in[199];
  assign inbar[200] = ~in[200];
  assign inbar[201] = ~in[201];
  assign inbar[202] = ~in[202];
  assign inbar[203] = ~in[203];
  assign inbar[204] = ~in[204];
  assign inbar[205] = ~in[205];
  assign inbar[206] = ~in[206];
  assign inbar[207] = ~in[207];
  assign inbar[208] = ~in[208];
  assign inbar[209] = ~in[209];
  assign inbar[210] = ~in[210];
  assign inbar[211] = ~in[211];
  assign inbar[212] = ~in[212];
  assign inbar[213] = ~in[213];
  assign inbar[214] = ~in[214];
  assign inbar[215] = ~in[215];
  assign inbar[216] = ~in[216];
  assign inbar[217] = ~in[217];
  assign inbar[218] = ~in[218];
  assign inbar[219] = ~in[219];
  assign inbar[220] = ~in[220];
  assign inbar[221] = ~in[221];
  assign inbar[222] = ~in[222];
  assign inbar[223] = ~in[223];
  assign inbar[224] = ~in[224];
  assign inbar[225] = ~in[225];
  assign inbar[226] = ~in[226];
  assign inbar[227] = ~in[227];
  assign inbar[228] = ~in[228];
  assign inbar[229] = ~in[229];
  assign inbar[230] = ~in[230];
  assign inbar[231] = ~in[231];
  assign inbar[232] = ~in[232];
  assign inbar[233] = ~in[233];
  assign inbar[234] = ~in[234];
  assign inbar[235] = ~in[235];
  assign inbar[236] = ~in[236];
  assign inbar[237] = ~in[237];
  assign inbar[238] = ~in[238];
  assign inbar[239] = ~in[239];
  assign inbar[240] = ~in[240];
  assign inbar[241] = ~in[241];
  assign inbar[242] = ~in[242];
  assign inbar[243] = ~in[243];
  assign inbar[244] = ~in[244];
  assign inbar[245] = ~in[245];
  assign inbar[246] = ~in[246];
  assign inbar[247] = ~in[247];
  assign inbar[248] = ~in[248];
  assign inbar[249] = ~in[249];
  assign inbar[250] = ~in[250];
  assign inbar[251] = ~in[251];
  assign inbar[252] = ~in[252];
  assign inbar[253] = ~in[253];
  assign inbar[254] = ~in[254];
  assign inbar[255] = ~in[255];
  //input_done

  output [7:0] out;
  reg [7:0] outbar;
  //output_done

  wire   in_81, in_80, in_79, in_78, in_77, in_76, in_75, in_74, in_73, in_72,
         in_71, in_70, in_69, in_68, in_67, in_66, in_65, in_64, in_63, in_62,
         in_61, in_60, in_59, in_58, in_57, in_56, in_55, in_54, in_53, in_52,
         in_51, in_50, in_49, in_48, in_47, in_46, in_45, in_44, in_43, in_42,
         in_41, in_40, in_39, in_38, in_37, in_36, in_35, in_34, in_33, in_32,
         in_31, in_30, in_29, in_28, in_27, in_26, in_25, in_24, in_23, in_22,
         in_21, in_20, in_19, in_18, in_17, in_16, in_15, in_14, in_13, in_12,
         in_11, in_10, in_9, in_8, in_7, in_6, in_5, in_4, in_3, in_2, in_1,
         in_0, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972;
  wire in_81bar, in_80bar, in_79bar, in_78bar, in_77bar, in_76bar, in_75bar, in_74bar, in_73bar, in_72bar, in_71bar, in_70bar, in_69bar, in_68bar, in_67bar, in_66bar, in_65bar, in_64bar, in_63bar, in_62bar, in_61bar, in_60bar, in_59bar, in_58bar, in_57bar, in_56bar, in_55bar, in_54bar, in_53bar, in_52bar, in_51bar, in_50bar, in_49bar, in_48bar, in_47bar, in_46bar, in_45bar, in_44bar, in_43bar, in_42bar, in_41bar, in_40bar, in_39bar, in_38bar, in_37bar, in_36bar, in_35bar, in_34bar, in_33bar, in_32bar, in_31bar, in_30bar, in_29bar, in_28bar, in_27bar, in_26bar, in_25bar, in_24bar, in_23bar, in_22bar, in_21bar, in_20bar, in_19bar, in_18bar, in_17bar, in_16bar, in_15bar, in_14bar, in_13bar, in_12bar, in_11bar, in_10bar, in_9bar, in_8bar, in_7bar, in_6bar, in_5bar, in_4bar, in_3bar, in_2bar, in_1bar, in_0bar, n487bar, n488bar, n489bar, n490bar, n491bar, n492bar, n493bar, n494bar, n495bar, n496bar, n497bar, n498bar, n499bar, n500bar, n501bar, n502bar, n503bar, n504bar, n505bar, n506bar, n507bar, n508bar, n509bar, n510bar, n511bar, n512bar, n513bar, n514bar, n515bar, n516bar, n517bar, n518bar, n519bar, n520bar, n521bar, n522bar, n523bar, n524bar, n525bar, n526bar, n527bar, n528bar, n529bar, n530bar, n531bar, n532bar, n533bar, n534bar, n535bar, n536bar, n537bar, n538bar, n539bar, n540bar, n541bar, n542bar, n543bar, n544bar, n545bar, n546bar, n547bar, n548bar, n549bar, n550bar, n551bar, n552bar, n553bar, n554bar, n555bar, n556bar, n557bar, n558bar, n559bar, n560bar, n561bar, n562bar, n563bar, n564bar, n565bar, n566bar, n567bar, n568bar, n569bar, n570bar, n571bar, n572bar, n573bar, n574bar, n575bar, n576bar, n577bar, n578bar, n579bar, n580bar, n581bar, n582bar, n583bar, n584bar, n585bar, n586bar, n587bar, n588bar, n589bar, n590bar, n591bar, n592bar, n593bar, n594bar, n595bar, n596bar, n597bar, n598bar, n599bar, n600bar, n601bar, n602bar, n603bar, n604bar, n605bar, n606bar, n607bar, n608bar, n609bar, n610bar, n611bar, n612bar, n613bar, n614bar, n615bar, n616bar, n617bar, n618bar, n619bar, n620bar, n621bar, n622bar, n623bar, n624bar, n625bar, n626bar, n627bar, n628bar, n629bar, n630bar, n631bar, n632bar, n633bar, n634bar, n635bar, n636bar, n637bar, n638bar, n639bar, n640bar, n641bar, n642bar, n643bar, n644bar, n645bar, n646bar, n647bar, n648bar, n649bar, n650bar, n651bar, n652bar, n653bar, n654bar, n655bar, n656bar, n657bar, n658bar, n659bar, n660bar, n661bar, n662bar, n663bar, n664bar, n665bar, n666bar, n667bar, n668bar, n669bar, n670bar, n671bar, n672bar, n673bar, n674bar, n675bar, n676bar, n677bar, n678bar, n679bar, n680bar, n681bar, n682bar, n683bar, n684bar, n685bar, n686bar, n687bar, n688bar, n689bar, n690bar, n691bar, n692bar, n693bar, n694bar, n695bar, n696bar, n697bar, n698bar, n699bar, n700bar, n701bar, n702bar, n703bar, n704bar, n705bar, n706bar, n707bar, n708bar, n709bar, n710bar, n711bar, n712bar, n713bar, n714bar, n715bar, n716bar, n717bar, n718bar, n719bar, n720bar, n721bar, n722bar, n723bar, n724bar, n725bar, n726bar, n727bar, n728bar, n729bar, n730bar, n731bar, n732bar, n733bar, n734bar, n735bar, n736bar, n737bar, n738bar, n739bar, n740bar, n741bar, n742bar, n743bar, n744bar, n745bar, n746bar, n747bar, n748bar, n749bar, n750bar, n751bar, n752bar, n753bar, n754bar, n755bar, n756bar, n757bar, n758bar, n759bar, n760bar, n761bar, n762bar, n763bar, n764bar, n765bar, n766bar, n767bar, n768bar, n769bar, n770bar, n771bar, n772bar, n773bar, n774bar, n775bar, n776bar, n777bar, n778bar, n779bar, n780bar, n781bar, n782bar, n783bar, n784bar, n785bar, n786bar, n787bar, n788bar, n789bar, n790bar, n791bar, n792bar, n793bar, n794bar, n795bar, n796bar, n797bar, n798bar, n799bar, n800bar, n801bar, n802bar, n803bar, n804bar, n805bar, n806bar, n807bar, n808bar, n809bar, n810bar, n811bar, n812bar, n813bar, n814bar, n815bar, n816bar, n817bar, n818bar, n819bar, n820bar, n821bar, n822bar, n823bar, n824bar, n825bar, n826bar, n827bar, n828bar, n829bar, n830bar, n831bar, n832bar, n833bar, n834bar, n835bar, n836bar, n837bar, n838bar, n839bar, n840bar, n841bar, n842bar, n843bar, n844bar, n845bar, n846bar, n847bar, n848bar, n849bar, n850bar, n851bar, n852bar, n853bar, n854bar, n855bar, n856bar, n857bar, n858bar, n859bar, n860bar, n861bar, n862bar, n863bar, n864bar, n865bar, n866bar, n867bar, n868bar, n869bar, n870bar, n871bar, n872bar, n873bar, n874bar, n875bar, n876bar, n877bar, n878bar, n879bar, n880bar, n881bar, n882bar, n883bar, n884bar, n885bar, n886bar, n887bar, n888bar, n889bar, n890bar, n891bar, n892bar, n893bar, n894bar, n895bar, n896bar, n897bar, n898bar, n899bar, n900bar, n901bar, n902bar, n903bar, n904bar, n905bar, n906bar, n907bar, n908bar, n909bar, n910bar, n911bar, n912bar, n913bar, n914bar, n915bar, n916bar, n917bar, n918bar, n919bar, n920bar, n921bar, n922bar, n923bar, n924bar, n925bar, n926bar, n927bar, n928bar, n929bar, n930bar, n931bar, n932bar, n933bar, n934bar, n935bar, n936bar, n937bar, n938bar, n939bar, n940bar, n941bar, n942bar, n943bar, n944bar, n945bar, n946bar, n947bar, n948bar, n949bar, n950bar, n951bar, n952bar, n953bar, n954bar, n955bar, n956bar, n957bar, n958bar, n959bar, n960bar, n961bar, n962bar, n963bar, n964bar, n965bar, n966bar, n967bar, n968bar, n969bar, n970bar, n971bar, n972bar;
  //wire_done
  
  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];

  OR2_X1 U1 ( .A1(n972), .A2(n971), .ZN(out[7]) );
  AND2_X1 U1bar ( .A1(n972bar), .A2(n971bar), .ZN(outbar[7]);
  OR2_X1 U2 ( .A1(n970), .A2(n969), .ZN(n971) );
  AND2_X1 U2bar ( .A1(n970bar), .A2(n969bar), .ZN(n971bar);
  OR2_X1 U3 ( .A1(n968), .A2(n967), .ZN(n969) );
  AND2_X1 U3bar ( .A1(n968bar), .A2(n967bar), .ZN(n969bar);
  OR2_X1 U4 ( .A1(n966), .A2(n965), .ZN(n967) );
  AND2_X1 U4bar ( .A1(n966bar), .A2(n965bar), .ZN(n967bar);
  OR2_X1 U5 ( .A1(n964), .A2(n963), .ZN(n968) );
  AND2_X1 U5bar ( .A1(n964bar), .A2(n963bar), .ZN(n968bar);
  OR2_X1 U6 ( .A1(in[116]), .A2(n962), .ZN(n963) );
  AND2_X1 U6bar ( .A1(inbar[116]), .A2(n962bar), .ZN(n963bar);
  OR2_X1 U7 ( .A1(n961), .A2(n960), .ZN(n970) );
  AND2_X1 U7bar ( .A1(n961bar), .A2(n960bar), .ZN(n970bar);
  OR2_X1 U8 ( .A1(in[150]), .A2(in[127]), .ZN(n960) );
  AND2_X1 U8bar ( .A1(inbar[150]), .A2(inbar[127]), .ZN(n960bar);
  OR2_X1 U9 ( .A1(in[160]), .A2(n959), .ZN(n961) );
  AND2_X1 U9bar ( .A1(inbar[160]), .A2(n959bar), .ZN(n961bar);
  OR2_X1 U10 ( .A1(in[252]), .A2(in[168]), .ZN(n959) );
  AND2_X1 U10bar ( .A1(inbar[252]), .A2(inbar[168]), .ZN(n959bar);
  OR2_X1 U11 ( .A1(n958), .A2(n957), .ZN(n972) );
  AND2_X1 U11bar ( .A1(n958bar), .A2(n957bar), .ZN(n972bar);
  OR2_X1 U12 ( .A1(n956), .A2(n955), .ZN(n957) );
  AND2_X1 U12bar ( .A1(n956bar), .A2(n955bar), .ZN(n957bar);
  OR2_X1 U13 ( .A1(in_17), .A2(in[96]), .ZN(n955) );
  AND2_X1 U13bar ( .A1(in_17bar), .A2(inbar[96]), .ZN(n955bar);
  OR2_X1 U14 ( .A1(in_23), .A2(n954), .ZN(n956) );
  AND2_X1 U14bar ( .A1(in_23bar), .A2(n954bar), .ZN(n956bar);
  OR2_X1 U15 ( .A1(in_31), .A2(in_26), .ZN(n954) );
  AND2_X1 U15bar ( .A1(in_31bar), .A2(in_26bar), .ZN(n954bar);
  OR2_X1 U16 ( .A1(n953), .A2(n952), .ZN(n958) );
  AND2_X1 U16bar ( .A1(n953bar), .A2(n952bar), .ZN(n958bar);
  OR2_X1 U17 ( .A1(in_58), .A2(in_4), .ZN(n952) );
  AND2_X1 U17bar ( .A1(in_58bar), .A2(in_4bar), .ZN(n952bar);
  OR2_X1 U18 ( .A1(in_59), .A2(n951), .ZN(n953) );
  AND2_X1 U18bar ( .A1(in_59bar), .A2(n951bar), .ZN(n953bar);
  OR2_X1 U19 ( .A1(in_71), .A2(in_62), .ZN(n951) );
  AND2_X1 U19bar ( .A1(in_71bar), .A2(in_62bar), .ZN(n951bar);
  OR2_X1 U20 ( .A1(n950), .A2(n949), .ZN(out[6]) );
  AND2_X1 U20bar ( .A1(n950bar), .A2(n949bar), .ZN(outbar[6]);
  OR2_X1 U21 ( .A1(n948), .A2(n947), .ZN(n949) );
  AND2_X1 U21bar ( .A1(n948bar), .A2(n947bar), .ZN(n949bar);
  OR2_X1 U22 ( .A1(n946), .A2(n945), .ZN(n947) );
  AND2_X1 U22bar ( .A1(n946bar), .A2(n945bar), .ZN(n947bar);
  OR2_X1 U23 ( .A1(n944), .A2(n943), .ZN(n945) );
  AND2_X1 U23bar ( .A1(n944bar), .A2(n943bar), .ZN(n945bar);
  OR2_X1 U24 ( .A1(n942), .A2(n941), .ZN(n946) );
  AND2_X1 U24bar ( .A1(n942bar), .A2(n941bar), .ZN(n946bar);
  OR2_X1 U25 ( .A1(in[101]), .A2(n940), .ZN(n941) );
  AND2_X1 U25bar ( .A1(inbar[101]), .A2(n940bar), .ZN(n941bar);
  OR2_X1 U26 ( .A1(n939), .A2(n938), .ZN(n948) );
  AND2_X1 U26bar ( .A1(n939bar), .A2(n938bar), .ZN(n948bar);
  OR2_X1 U27 ( .A1(in[114]), .A2(in[104]), .ZN(n938) );
  AND2_X1 U27bar ( .A1(inbar[114]), .A2(inbar[104]), .ZN(n938bar);
  OR2_X1 U28 ( .A1(in[128]), .A2(n937), .ZN(n939) );
  AND2_X1 U28bar ( .A1(inbar[128]), .A2(n937bar), .ZN(n939bar);
  OR2_X1 U29 ( .A1(in[136]), .A2(in[134]), .ZN(n937) );
  AND2_X1 U29bar ( .A1(inbar[136]), .A2(inbar[134]), .ZN(n937bar);
  OR2_X1 U30 ( .A1(n936), .A2(n935), .ZN(n950) );
  AND2_X1 U30bar ( .A1(n936bar), .A2(n935bar), .ZN(n950bar);
  OR2_X1 U31 ( .A1(n934), .A2(n933), .ZN(n935) );
  AND2_X1 U31bar ( .A1(n934bar), .A2(n933bar), .ZN(n935bar);
  OR2_X1 U32 ( .A1(in[177]), .A2(in[164]), .ZN(n933) );
  AND2_X1 U32bar ( .A1(inbar[177]), .A2(inbar[164]), .ZN(n933bar);
  OR2_X1 U33 ( .A1(in[212]), .A2(n932), .ZN(n934) );
  AND2_X1 U33bar ( .A1(inbar[212]), .A2(n932bar), .ZN(n934bar);
  OR2_X1 U34 ( .A1(in[248]), .A2(in[221]), .ZN(n932) );
  AND2_X1 U34bar ( .A1(inbar[248]), .A2(inbar[221]), .ZN(n932bar);
  OR2_X1 U35 ( .A1(n931), .A2(n930), .ZN(n936) );
  AND2_X1 U35bar ( .A1(n931bar), .A2(n930bar), .ZN(n936bar);
  OR2_X1 U36 ( .A1(in_18), .A2(in[93]), .ZN(n930) );
  AND2_X1 U36bar ( .A1(in_18bar), .A2(inbar[93]), .ZN(n930bar);
  OR2_X1 U37 ( .A1(in_31), .A2(n929), .ZN(n931) );
  AND2_X1 U37bar ( .A1(in_31bar), .A2(n929bar), .ZN(n931bar);
  OR2_X1 U38 ( .A1(in_7), .A2(in_39), .ZN(n929) );
  AND2_X1 U38bar ( .A1(in_7bar), .A2(in_39bar), .ZN(n929bar);
  OR2_X1 U39 ( .A1(n928), .A2(n927), .ZN(out[5]) );
  AND2_X1 U39bar ( .A1(n928bar), .A2(n927bar), .ZN(outbar[5]);
  OR2_X1 U40 ( .A1(n926), .A2(n925), .ZN(n927) );
  AND2_X1 U40bar ( .A1(n926bar), .A2(n925bar), .ZN(n927bar);
  OR2_X1 U41 ( .A1(n924), .A2(n923), .ZN(n925) );
  AND2_X1 U41bar ( .A1(n924bar), .A2(n923bar), .ZN(n925bar);
  OR2_X1 U42 ( .A1(n922), .A2(n921), .ZN(n923) );
  AND2_X1 U42bar ( .A1(n922bar), .A2(n921bar), .ZN(n923bar);
  OR2_X1 U43 ( .A1(n940), .A2(n920), .ZN(n924) );
  AND2_X1 U43bar ( .A1(n940bar), .A2(n920bar), .ZN(n924bar);
  OR2_X1 U44 ( .A1(in[111]), .A2(n919), .ZN(n920) );
  AND2_X1 U44bar ( .A1(inbar[111]), .A2(n919bar), .ZN(n920bar);
  OR2_X1 U45 ( .A1(n918), .A2(n917), .ZN(n940) );
  AND2_X1 U45bar ( .A1(n918bar), .A2(n917bar), .ZN(n940bar);
  OR2_X1 U46 ( .A1(n916), .A2(n915), .ZN(n917) );
  AND2_X1 U46bar ( .A1(n916bar), .A2(n915bar), .ZN(n917bar);
  OR2_X1 U47 ( .A1(n914), .A2(n913), .ZN(n915) );
  AND2_X1 U47bar ( .A1(n914bar), .A2(n913bar), .ZN(n915bar);
  OR2_X1 U48 ( .A1(in[140]), .A2(in[131]), .ZN(n913) );
  AND2_X1 U48bar ( .A1(inbar[140]), .A2(inbar[131]), .ZN(n913bar);
  OR2_X1 U49 ( .A1(in[160]), .A2(in[144]), .ZN(n914) );
  AND2_X1 U49bar ( .A1(inbar[160]), .A2(inbar[144]), .ZN(n914bar);
  OR2_X1 U50 ( .A1(n912), .A2(n911), .ZN(n916) );
  AND2_X1 U50bar ( .A1(n912bar), .A2(n911bar), .ZN(n916bar);
  OR2_X1 U51 ( .A1(in[179]), .A2(in[174]), .ZN(n911) );
  AND2_X1 U51bar ( .A1(inbar[179]), .A2(inbar[174]), .ZN(n911bar);
  OR2_X1 U52 ( .A1(in[188]), .A2(in[184]), .ZN(n912) );
  AND2_X1 U52bar ( .A1(inbar[188]), .A2(inbar[184]), .ZN(n912bar);
  OR2_X1 U53 ( .A1(n910), .A2(n909), .ZN(n918) );
  AND2_X1 U53bar ( .A1(n910bar), .A2(n909bar), .ZN(n918bar);
  OR2_X1 U54 ( .A1(n908), .A2(n907), .ZN(n909) );
  AND2_X1 U54bar ( .A1(n908bar), .A2(n907bar), .ZN(n909bar);
  OR2_X1 U55 ( .A1(in[216]), .A2(in[200]), .ZN(n907) );
  AND2_X1 U55bar ( .A1(inbar[216]), .A2(inbar[200]), .ZN(n907bar);
  OR2_X1 U56 ( .A1(in[228]), .A2(in[224]), .ZN(n908) );
  AND2_X1 U56bar ( .A1(inbar[228]), .A2(inbar[224]), .ZN(n908bar);
  OR2_X1 U57 ( .A1(n906), .A2(n905), .ZN(n910) );
  AND2_X1 U57bar ( .A1(n906bar), .A2(n905bar), .ZN(n910bar);
  OR2_X1 U58 ( .A1(in[247]), .A2(in[235]), .ZN(n905) );
  AND2_X1 U58bar ( .A1(inbar[247]), .A2(inbar[235]), .ZN(n905bar);
  OR2_X1 U59 ( .A1(in_42), .A2(in[83]), .ZN(n906) );
  AND2_X1 U59bar ( .A1(in_42bar), .A2(inbar[83]), .ZN(n906bar);
  OR2_X1 U60 ( .A1(n904), .A2(n903), .ZN(n926) );
  AND2_X1 U60bar ( .A1(n904bar), .A2(n903bar), .ZN(n926bar);
  OR2_X1 U61 ( .A1(in[166]), .A2(in[123]), .ZN(n903) );
  AND2_X1 U61bar ( .A1(inbar[166]), .A2(inbar[123]), .ZN(n903bar);
  OR2_X1 U62 ( .A1(in[170]), .A2(n902), .ZN(n904) );
  AND2_X1 U62bar ( .A1(inbar[170]), .A2(n902bar), .ZN(n904bar);
  OR2_X1 U63 ( .A1(in[194]), .A2(in[183]), .ZN(n902) );
  AND2_X1 U63bar ( .A1(inbar[194]), .A2(inbar[183]), .ZN(n902bar);
  OR2_X1 U64 ( .A1(n901), .A2(n900), .ZN(n928) );
  AND2_X1 U64bar ( .A1(n901bar), .A2(n900bar), .ZN(n928bar);
  OR2_X1 U65 ( .A1(n899), .A2(n898), .ZN(n900) );
  AND2_X1 U65bar ( .A1(n899bar), .A2(n898bar), .ZN(n900bar);
  OR2_X1 U66 ( .A1(in[241]), .A2(in[238]), .ZN(n898) );
  AND2_X1 U66bar ( .A1(inbar[241]), .A2(inbar[238]), .ZN(n898bar);
  OR2_X1 U67 ( .A1(in[250]), .A2(n897), .ZN(n899) );
  AND2_X1 U67bar ( .A1(inbar[250]), .A2(n897bar), .ZN(n899bar);
  OR2_X1 U68 ( .A1(in_24), .A2(in[84]), .ZN(n897) );
  AND2_X1 U68bar ( .A1(in_24bar), .A2(inbar[84]), .ZN(n897bar);
  OR2_X1 U69 ( .A1(n896), .A2(n895), .ZN(n901) );
  AND2_X1 U69bar ( .A1(n896bar), .A2(n895bar), .ZN(n901bar);
  OR2_X1 U70 ( .A1(in_41), .A2(in_29), .ZN(n895) );
  AND2_X1 U70bar ( .A1(in_41bar), .A2(in_29bar), .ZN(n895bar);
  OR2_X1 U71 ( .A1(in_66), .A2(n894), .ZN(n896) );
  AND2_X1 U71bar ( .A1(in_66bar), .A2(n894bar), .ZN(n896bar);
  OR2_X1 U72 ( .A1(in_76), .A2(in_71), .ZN(n894) );
  AND2_X1 U72bar ( .A1(in_76bar), .A2(in_71bar), .ZN(n894bar);
  OR2_X1 U73 ( .A1(n893), .A2(n892), .ZN(out[4]) );
  AND2_X1 U73bar ( .A1(n893bar), .A2(n892bar), .ZN(outbar[4]);
  OR2_X1 U74 ( .A1(n891), .A2(n890), .ZN(n892) );
  AND2_X1 U74bar ( .A1(n891bar), .A2(n890bar), .ZN(n892bar);
  OR2_X1 U75 ( .A1(n889), .A2(n888), .ZN(n890) );
  AND2_X1 U75bar ( .A1(n889bar), .A2(n888bar), .ZN(n890bar);
  OR2_X1 U76 ( .A1(n922), .A2(n887), .ZN(n888) );
  AND2_X1 U76bar ( .A1(n922bar), .A2(n887bar), .ZN(n888bar);
  OR2_X1 U77 ( .A1(n886), .A2(n885), .ZN(n922) );
  AND2_X1 U77bar ( .A1(n886bar), .A2(n885bar), .ZN(n922bar);
  OR2_X1 U78 ( .A1(n884), .A2(n883), .ZN(n885) );
  AND2_X1 U78bar ( .A1(n884bar), .A2(n883bar), .ZN(n885bar);
  OR2_X1 U79 ( .A1(n882), .A2(n881), .ZN(n883) );
  AND2_X1 U79bar ( .A1(n882bar), .A2(n881bar), .ZN(n883bar);
  OR2_X1 U80 ( .A1(in[118]), .A2(in[109]), .ZN(n881) );
  AND2_X1 U80bar ( .A1(inbar[118]), .A2(inbar[109]), .ZN(n881bar);
  OR2_X1 U81 ( .A1(in[139]), .A2(in[120]), .ZN(n882) );
  AND2_X1 U81bar ( .A1(inbar[139]), .A2(inbar[120]), .ZN(n882bar);
  OR2_X1 U82 ( .A1(n880), .A2(n879), .ZN(n884) );
  AND2_X1 U82bar ( .A1(n880bar), .A2(n879bar), .ZN(n884bar);
  OR2_X1 U83 ( .A1(in[198]), .A2(in[154]), .ZN(n879) );
  AND2_X1 U83bar ( .A1(inbar[198]), .A2(inbar[154]), .ZN(n879bar);
  OR2_X1 U84 ( .A1(in[210]), .A2(in[205]), .ZN(n880) );
  AND2_X1 U84bar ( .A1(inbar[210]), .A2(inbar[205]), .ZN(n880bar);
  OR2_X1 U85 ( .A1(n878), .A2(n877), .ZN(n886) );
  AND2_X1 U85bar ( .A1(n878bar), .A2(n877bar), .ZN(n886bar);
  OR2_X1 U86 ( .A1(n876), .A2(n875), .ZN(n877) );
  AND2_X1 U86bar ( .A1(n876bar), .A2(n875bar), .ZN(n877bar);
  OR2_X1 U87 ( .A1(in[219]), .A2(in[217]), .ZN(n875) );
  AND2_X1 U87bar ( .A1(inbar[219]), .A2(inbar[217]), .ZN(n875bar);
  OR2_X1 U88 ( .A1(in[86]), .A2(in[252]), .ZN(n876) );
  AND2_X1 U88bar ( .A1(inbar[86]), .A2(inbar[252]), .ZN(n876bar);
  OR2_X1 U89 ( .A1(n874), .A2(n873), .ZN(n878) );
  AND2_X1 U89bar ( .A1(n874bar), .A2(n873bar), .ZN(n878bar);
  OR2_X1 U90 ( .A1(in_40), .A2(in[91]), .ZN(n873) );
  AND2_X1 U90bar ( .A1(in_40bar), .A2(inbar[91]), .ZN(n873bar);
  OR2_X1 U91 ( .A1(in_8), .A2(in_46), .ZN(n874) );
  AND2_X1 U91bar ( .A1(in_8bar), .A2(in_46bar), .ZN(n874bar);
  OR2_X1 U92 ( .A1(n872), .A2(n871), .ZN(n889) );
  AND2_X1 U92bar ( .A1(n872bar), .A2(n871bar), .ZN(n889bar);
  OR2_X1 U93 ( .A1(in[117]), .A2(n943), .ZN(n871) );
  AND2_X1 U93bar ( .A1(inbar[117]), .A2(n943bar), .ZN(n871bar);
  OR2_X1 U94 ( .A1(n870), .A2(n869), .ZN(n943) );
  AND2_X1 U94bar ( .A1(n870bar), .A2(n869bar), .ZN(n943bar);
  OR2_X1 U95 ( .A1(n868), .A2(n867), .ZN(n869) );
  AND2_X1 U95bar ( .A1(n868bar), .A2(n867bar), .ZN(n869bar);
  OR2_X1 U96 ( .A1(n866), .A2(n865), .ZN(n867) );
  AND2_X1 U96bar ( .A1(n866bar), .A2(n865bar), .ZN(n867bar);
  OR2_X1 U97 ( .A1(n864), .A2(n863), .ZN(n865) );
  AND2_X1 U97bar ( .A1(n864bar), .A2(n863bar), .ZN(n865bar);
  OR2_X1 U98 ( .A1(in[108]), .A2(n919), .ZN(n866) );
  AND2_X1 U98bar ( .A1(inbar[108]), .A2(n919bar), .ZN(n866bar);
  OR2_X1 U99 ( .A1(n862), .A2(n861), .ZN(n919) );
  AND2_X1 U99bar ( .A1(n862bar), .A2(n861bar), .ZN(n919bar);
  OR2_X1 U100 ( .A1(n860), .A2(n859), .ZN(n861) );
  AND2_X1 U100bar ( .A1(n860bar), .A2(n859bar), .ZN(n861bar);
  OR2_X1 U101 ( .A1(n858), .A2(n857), .ZN(n859) );
  AND2_X1 U101bar ( .A1(n858bar), .A2(n857bar), .ZN(n859bar);
  OR2_X1 U102 ( .A1(in[119]), .A2(in[105]), .ZN(n857) );
  AND2_X1 U102bar ( .A1(inbar[119]), .A2(inbar[105]), .ZN(n857bar);
  OR2_X1 U103 ( .A1(in[186]), .A2(in[175]), .ZN(n858) );
  AND2_X1 U103bar ( .A1(inbar[186]), .A2(inbar[175]), .ZN(n858bar);
  OR2_X1 U104 ( .A1(n856), .A2(n855), .ZN(n860) );
  AND2_X1 U104bar ( .A1(n856bar), .A2(n855bar), .ZN(n860bar);
  OR2_X1 U105 ( .A1(in[202]), .A2(in[193]), .ZN(n855) );
  AND2_X1 U105bar ( .A1(inbar[202]), .A2(inbar[193]), .ZN(n855bar);
  OR2_X1 U106 ( .A1(in[225]), .A2(in[208]), .ZN(n856) );
  AND2_X1 U106bar ( .A1(inbar[225]), .A2(inbar[208]), .ZN(n856bar);
  OR2_X1 U107 ( .A1(n854), .A2(n853), .ZN(n862) );
  AND2_X1 U107bar ( .A1(n854bar), .A2(n853bar), .ZN(n862bar);
  OR2_X1 U108 ( .A1(n852), .A2(n851), .ZN(n853) );
  AND2_X1 U108bar ( .A1(n852bar), .A2(n851bar), .ZN(n853bar);
  OR2_X1 U109 ( .A1(in_1), .A2(in[85]), .ZN(n851) );
  AND2_X1 U109bar ( .A1(in_1bar), .A2(inbar[85]), .ZN(n851bar);
  OR2_X1 U110 ( .A1(in_23), .A2(in_19), .ZN(n852) );
  AND2_X1 U110bar ( .A1(in_23bar), .A2(in_19bar), .ZN(n852bar);
  OR2_X1 U111 ( .A1(n850), .A2(n849), .ZN(n854) );
  AND2_X1 U111bar ( .A1(n850bar), .A2(n849bar), .ZN(n854bar);
  OR2_X1 U112 ( .A1(in_43), .A2(in_33), .ZN(n849) );
  AND2_X1 U112bar ( .A1(in_43bar), .A2(in_33bar), .ZN(n849bar);
  OR2_X1 U113 ( .A1(in_63), .A2(in_44), .ZN(n850) );
  AND2_X1 U113bar ( .A1(in_63bar), .A2(in_44bar), .ZN(n850bar);
  OR2_X1 U114 ( .A1(n848), .A2(n847), .ZN(n868) );
  AND2_X1 U114bar ( .A1(n848bar), .A2(n847bar), .ZN(n868bar);
  OR2_X1 U115 ( .A1(in[141]), .A2(in[112]), .ZN(n847) );
  AND2_X1 U115bar ( .A1(inbar[141]), .A2(inbar[112]), .ZN(n847bar);
  OR2_X1 U116 ( .A1(in[147]), .A2(n846), .ZN(n848) );
  AND2_X1 U116bar ( .A1(inbar[147]), .A2(n846bar), .ZN(n848bar);
  OR2_X1 U117 ( .A1(in[181]), .A2(in[167]), .ZN(n846) );
  AND2_X1 U117bar ( .A1(inbar[181]), .A2(inbar[167]), .ZN(n846bar);
  OR2_X1 U118 ( .A1(n845), .A2(n844), .ZN(n870) );
  AND2_X1 U118bar ( .A1(n845bar), .A2(n844bar), .ZN(n870bar);
  OR2_X1 U119 ( .A1(n843), .A2(n842), .ZN(n844) );
  AND2_X1 U119bar ( .A1(n843bar), .A2(n842bar), .ZN(n844bar);
  OR2_X1 U120 ( .A1(in[229]), .A2(in[201]), .ZN(n842) );
  AND2_X1 U120bar ( .A1(inbar[229]), .A2(inbar[201]), .ZN(n842bar);
  OR2_X1 U121 ( .A1(in[237]), .A2(n841), .ZN(n843) );
  AND2_X1 U121bar ( .A1(inbar[237]), .A2(n841bar), .ZN(n843bar);
  OR2_X1 U122 ( .A1(in[94]), .A2(in[253]), .ZN(n841) );
  AND2_X1 U122bar ( .A1(inbar[94]), .A2(inbar[253]), .ZN(n841bar);
  OR2_X1 U123 ( .A1(n840), .A2(n839), .ZN(n845) );
  AND2_X1 U123bar ( .A1(n840bar), .A2(n839bar), .ZN(n845bar);
  OR2_X1 U124 ( .A1(in_21), .A2(in[96]), .ZN(n839) );
  AND2_X1 U124bar ( .A1(in_21bar), .A2(inbar[96]), .ZN(n839bar);
  OR2_X1 U125 ( .A1(in_25), .A2(n838), .ZN(n840) );
  AND2_X1 U125bar ( .A1(in_25bar), .A2(n838bar), .ZN(n840bar);
  OR2_X1 U126 ( .A1(in_81), .A2(in_45), .ZN(n838) );
  AND2_X1 U126bar ( .A1(in_81bar), .A2(in_45bar), .ZN(n838bar);
  OR2_X1 U127 ( .A1(n837), .A2(n836), .ZN(n891) );
  AND2_X1 U127bar ( .A1(n837bar), .A2(n836bar), .ZN(n891bar);
  OR2_X1 U128 ( .A1(in[142]), .A2(in[124]), .ZN(n836) );
  AND2_X1 U128bar ( .A1(inbar[142]), .A2(inbar[124]), .ZN(n836bar);
  OR2_X1 U129 ( .A1(in[150]), .A2(n835), .ZN(n837) );
  AND2_X1 U129bar ( .A1(inbar[150]), .A2(n835bar), .ZN(n837bar);
  OR2_X1 U130 ( .A1(in[172]), .A2(in[155]), .ZN(n835) );
  AND2_X1 U130bar ( .A1(inbar[172]), .A2(inbar[155]), .ZN(n835bar);
  OR2_X1 U131 ( .A1(n834), .A2(n833), .ZN(n893) );
  AND2_X1 U131bar ( .A1(n834bar), .A2(n833bar), .ZN(n893bar);
  OR2_X1 U132 ( .A1(n832), .A2(n831), .ZN(n833) );
  AND2_X1 U132bar ( .A1(n832bar), .A2(n831bar), .ZN(n833bar);
  OR2_X1 U133 ( .A1(in[196]), .A2(in[173]), .ZN(n831) );
  AND2_X1 U133bar ( .A1(inbar[196]), .A2(inbar[173]), .ZN(n831bar);
  OR2_X1 U134 ( .A1(in[222]), .A2(n830), .ZN(n832) );
  AND2_X1 U134bar ( .A1(inbar[222]), .A2(n830bar), .ZN(n832bar);
  OR2_X1 U135 ( .A1(in[227]), .A2(in[226]), .ZN(n830) );
  AND2_X1 U135bar ( .A1(inbar[227]), .A2(inbar[226]), .ZN(n830bar);
  OR2_X1 U136 ( .A1(n829), .A2(n828), .ZN(n834) );
  AND2_X1 U136bar ( .A1(n829bar), .A2(n828bar), .ZN(n834bar);
  OR2_X1 U137 ( .A1(in[249]), .A2(in[231]), .ZN(n828) );
  AND2_X1 U137bar ( .A1(inbar[249]), .A2(inbar[231]), .ZN(n828bar);
  OR2_X1 U138 ( .A1(in_28), .A2(n827), .ZN(n829) );
  AND2_X1 U138bar ( .A1(in_28bar), .A2(n827bar), .ZN(n829bar);
  OR2_X1 U139 ( .A1(in_52), .A2(in_47), .ZN(n827) );
  AND2_X1 U139bar ( .A1(in_52bar), .A2(in_47bar), .ZN(n827bar);
  OR2_X1 U140 ( .A1(n826), .A2(n825), .ZN(out[3]) );
  AND2_X1 U140bar ( .A1(n826bar), .A2(n825bar), .ZN(outbar[3]);
  OR2_X1 U141 ( .A1(n824), .A2(n823), .ZN(n825) );
  AND2_X1 U141bar ( .A1(n824bar), .A2(n823bar), .ZN(n825bar);
  OR2_X1 U142 ( .A1(n822), .A2(n821), .ZN(n823) );
  AND2_X1 U142bar ( .A1(n822bar), .A2(n821bar), .ZN(n823bar);
  OR2_X1 U143 ( .A1(n820), .A2(n819), .ZN(n821) );
  AND2_X1 U143bar ( .A1(n820bar), .A2(n819bar), .ZN(n821bar);
  OR2_X1 U144 ( .A1(n964), .A2(n818), .ZN(n822) );
  AND2_X1 U144bar ( .A1(n964bar), .A2(n818bar), .ZN(n822bar);
  OR2_X1 U145 ( .A1(in[118]), .A2(n817), .ZN(n818) );
  AND2_X1 U145bar ( .A1(inbar[118]), .A2(n817bar), .ZN(n818bar);
  OR2_X1 U146 ( .A1(n816), .A2(n815), .ZN(n964) );
  AND2_X1 U146bar ( .A1(n816bar), .A2(n815bar), .ZN(n964bar);
  OR2_X1 U147 ( .A1(n814), .A2(n813), .ZN(n815) );
  AND2_X1 U147bar ( .A1(n814bar), .A2(n813bar), .ZN(n815bar);
  OR2_X1 U148 ( .A1(n812), .A2(n811), .ZN(n813) );
  AND2_X1 U148bar ( .A1(n812bar), .A2(n811bar), .ZN(n813bar);
  OR2_X1 U149 ( .A1(in[122]), .A2(in[111]), .ZN(n811) );
  AND2_X1 U149bar ( .A1(inbar[122]), .A2(inbar[111]), .ZN(n811bar);
  OR2_X1 U150 ( .A1(in[154]), .A2(in[151]), .ZN(n812) );
  AND2_X1 U150bar ( .A1(inbar[154]), .A2(inbar[151]), .ZN(n812bar);
  OR2_X1 U151 ( .A1(n810), .A2(n809), .ZN(n814) );
  AND2_X1 U151bar ( .A1(n810bar), .A2(n809bar), .ZN(n814bar);
  OR2_X1 U152 ( .A1(in[187]), .A2(in[177]), .ZN(n809) );
  AND2_X1 U152bar ( .A1(inbar[187]), .A2(inbar[177]), .ZN(n809bar);
  OR2_X1 U153 ( .A1(in[200]), .A2(in[192]), .ZN(n810) );
  AND2_X1 U153bar ( .A1(inbar[200]), .A2(inbar[192]), .ZN(n810bar);
  OR2_X1 U154 ( .A1(n808), .A2(n807), .ZN(n816) );
  AND2_X1 U154bar ( .A1(n808bar), .A2(n807bar), .ZN(n816bar);
  OR2_X1 U155 ( .A1(n806), .A2(n805), .ZN(n807) );
  AND2_X1 U155bar ( .A1(n806bar), .A2(n805bar), .ZN(n807bar);
  OR2_X1 U156 ( .A1(in[225]), .A2(in[207]), .ZN(n805) );
  AND2_X1 U156bar ( .A1(inbar[225]), .A2(inbar[207]), .ZN(n805bar);
  OR2_X1 U157 ( .A1(in[98]), .A2(in[226]), .ZN(n806) );
  AND2_X1 U157bar ( .A1(inbar[98]), .A2(inbar[226]), .ZN(n806bar);
  OR2_X1 U158 ( .A1(n804), .A2(n803), .ZN(n808) );
  AND2_X1 U158bar ( .A1(n804bar), .A2(n803bar), .ZN(n808bar);
  OR2_X1 U159 ( .A1(in_20), .A2(in_16), .ZN(n803) );
  AND2_X1 U159bar ( .A1(in_20bar), .A2(in_16bar), .ZN(n803bar);
  OR2_X1 U160 ( .A1(in_55), .A2(in_45), .ZN(n804) );
  AND2_X1 U160bar ( .A1(in_55bar), .A2(in_45bar), .ZN(n804bar);
  OR2_X1 U161 ( .A1(n802), .A2(n801), .ZN(n824) );
  AND2_X1 U161bar ( .A1(n802bar), .A2(n801bar), .ZN(n824bar);
  OR2_X1 U162 ( .A1(in[162]), .A2(in[149]), .ZN(n801) );
  AND2_X1 U162bar ( .A1(inbar[162]), .A2(inbar[149]), .ZN(n801bar);
  OR2_X1 U163 ( .A1(in[163]), .A2(n800), .ZN(n802) );
  AND2_X1 U163bar ( .A1(inbar[163]), .A2(n800bar), .ZN(n802bar);
  OR2_X1 U164 ( .A1(in[191]), .A2(in[189]), .ZN(n800) );
  AND2_X1 U164bar ( .A1(inbar[191]), .A2(inbar[189]), .ZN(n800bar);
  OR2_X1 U165 ( .A1(n799), .A2(n798), .ZN(n826) );
  AND2_X1 U165bar ( .A1(n799bar), .A2(n798bar), .ZN(n826bar);
  OR2_X1 U166 ( .A1(n797), .A2(n796), .ZN(n798) );
  AND2_X1 U166bar ( .A1(n797bar), .A2(n796bar), .ZN(n798bar);
  OR2_X1 U167 ( .A1(in[212]), .A2(in[193]), .ZN(n796) );
  AND2_X1 U167bar ( .A1(inbar[212]), .A2(inbar[193]), .ZN(n796bar);
  OR2_X1 U168 ( .A1(in[238]), .A2(n795), .ZN(n797) );
  AND2_X1 U168bar ( .A1(inbar[238]), .A2(n795bar), .ZN(n797bar);
  OR2_X1 U169 ( .A1(in[88]), .A2(in[247]), .ZN(n795) );
  AND2_X1 U169bar ( .A1(inbar[88]), .A2(inbar[247]), .ZN(n795bar);
  OR2_X1 U170 ( .A1(n794), .A2(n793), .ZN(n799) );
  AND2_X1 U170bar ( .A1(n794bar), .A2(n793bar), .ZN(n799bar);
  OR2_X1 U171 ( .A1(in[94]), .A2(in[92]), .ZN(n793) );
  AND2_X1 U171bar ( .A1(inbar[94]), .A2(inbar[92]), .ZN(n793bar);
  OR2_X1 U172 ( .A1(in_52), .A2(n792), .ZN(n794) );
  AND2_X1 U172bar ( .A1(in_52bar), .A2(n792bar), .ZN(n794bar);
  OR2_X1 U173 ( .A1(in_70), .A2(in_67), .ZN(n792) );
  AND2_X1 U173bar ( .A1(in_70bar), .A2(in_67bar), .ZN(n792bar);
  OR2_X1 U174 ( .A1(n791), .A2(n790), .ZN(out[2]) );
  AND2_X1 U174bar ( .A1(n791bar), .A2(n790bar), .ZN(outbar[2]);
  OR2_X1 U175 ( .A1(n789), .A2(n788), .ZN(n790) );
  AND2_X1 U175bar ( .A1(n789bar), .A2(n788bar), .ZN(n790bar);
  OR2_X1 U176 ( .A1(n787), .A2(n786), .ZN(n788) );
  AND2_X1 U176bar ( .A1(n787bar), .A2(n786bar), .ZN(n788bar);
  OR2_X1 U177 ( .A1(n819), .A2(n785), .ZN(n786) );
  AND2_X1 U177bar ( .A1(n819bar), .A2(n785bar), .ZN(n786bar);
  OR2_X1 U178 ( .A1(n784), .A2(n783), .ZN(n819) );
  AND2_X1 U178bar ( .A1(n784bar), .A2(n783bar), .ZN(n819bar);
  OR2_X1 U179 ( .A1(n782), .A2(n781), .ZN(n783) );
  AND2_X1 U179bar ( .A1(n782bar), .A2(n781bar), .ZN(n783bar);
  OR2_X1 U180 ( .A1(n780), .A2(n779), .ZN(n781) );
  AND2_X1 U180bar ( .A1(n780bar), .A2(n779bar), .ZN(n781bar);
  OR2_X1 U181 ( .A1(n962), .A2(n778), .ZN(n779) );
  AND2_X1 U181bar ( .A1(n962bar), .A2(n778bar), .ZN(n779bar);
  OR2_X1 U182 ( .A1(n777), .A2(n776), .ZN(n962) );
  AND2_X1 U182bar ( .A1(n777bar), .A2(n776bar), .ZN(n962bar);
  OR2_X1 U183 ( .A1(n775), .A2(n774), .ZN(n776) );
  AND2_X1 U183bar ( .A1(n775bar), .A2(n774bar), .ZN(n776bar);
  OR2_X1 U184 ( .A1(n773), .A2(n772), .ZN(n774) );
  AND2_X1 U184bar ( .A1(n773bar), .A2(n772bar), .ZN(n774bar);
  OR2_X1 U185 ( .A1(in[131]), .A2(in[120]), .ZN(n772) );
  AND2_X1 U185bar ( .A1(inbar[131]), .A2(inbar[120]), .ZN(n772bar);
  OR2_X1 U186 ( .A1(in[153]), .A2(in[147]), .ZN(n773) );
  AND2_X1 U186bar ( .A1(inbar[153]), .A2(inbar[147]), .ZN(n773bar);
  OR2_X1 U187 ( .A1(n771), .A2(n770), .ZN(n775) );
  AND2_X1 U187bar ( .A1(n771bar), .A2(n770bar), .ZN(n775bar);
  OR2_X1 U188 ( .A1(in[170]), .A2(in[156]), .ZN(n770) );
  AND2_X1 U188bar ( .A1(inbar[170]), .A2(inbar[156]), .ZN(n770bar);
  OR2_X1 U189 ( .A1(in[223]), .A2(in[190]), .ZN(n771) );
  AND2_X1 U189bar ( .A1(inbar[223]), .A2(inbar[190]), .ZN(n771bar);
  OR2_X1 U190 ( .A1(n769), .A2(n768), .ZN(n777) );
  AND2_X1 U190bar ( .A1(n769bar), .A2(n768bar), .ZN(n777bar);
  OR2_X1 U191 ( .A1(n767), .A2(n766), .ZN(n768) );
  AND2_X1 U191bar ( .A1(n767bar), .A2(n766bar), .ZN(n768bar);
  OR2_X1 U192 ( .A1(in[236]), .A2(in[230]), .ZN(n766) );
  AND2_X1 U192bar ( .A1(inbar[236]), .A2(inbar[230]), .ZN(n766bar);
  OR2_X1 U193 ( .A1(in[85]), .A2(in[240]), .ZN(n767) );
  AND2_X1 U193bar ( .A1(inbar[85]), .A2(inbar[240]), .ZN(n767bar);
  OR2_X1 U194 ( .A1(n765), .A2(n764), .ZN(n769) );
  AND2_X1 U194bar ( .A1(n765bar), .A2(n764bar), .ZN(n769bar);
  OR2_X1 U195 ( .A1(in_12), .A2(in[90]), .ZN(n764) );
  AND2_X1 U195bar ( .A1(in_12bar), .A2(inbar[90]), .ZN(n764bar);
  OR2_X1 U196 ( .A1(in_39), .A2(in_28), .ZN(n765) );
  AND2_X1 U196bar ( .A1(in_39bar), .A2(in_28bar), .ZN(n765bar);
  OR2_X1 U197 ( .A1(in[109]), .A2(n763), .ZN(n780) );
  AND2_X1 U197bar ( .A1(inbar[109]), .A2(n763bar), .ZN(n780bar);
  OR2_X1 U198 ( .A1(n762), .A2(n761), .ZN(n782) );
  AND2_X1 U198bar ( .A1(n762bar), .A2(n761bar), .ZN(n782bar);
  OR2_X1 U199 ( .A1(in[138]), .A2(in[129]), .ZN(n761) );
  AND2_X1 U199bar ( .A1(inbar[138]), .A2(inbar[129]), .ZN(n761bar);
  OR2_X1 U200 ( .A1(in[157]), .A2(n760), .ZN(n762) );
  AND2_X1 U200bar ( .A1(inbar[157]), .A2(n760bar), .ZN(n762bar);
  OR2_X1 U201 ( .A1(in[182]), .A2(in[167]), .ZN(n760) );
  AND2_X1 U201bar ( .A1(inbar[182]), .A2(inbar[167]), .ZN(n760bar);
  OR2_X1 U202 ( .A1(n759), .A2(n758), .ZN(n784) );
  AND2_X1 U202bar ( .A1(n759bar), .A2(n758bar), .ZN(n784bar);
  OR2_X1 U203 ( .A1(n757), .A2(n756), .ZN(n758) );
  AND2_X1 U203bar ( .A1(n757bar), .A2(n756bar), .ZN(n758bar);
  OR2_X1 U204 ( .A1(in[195]), .A2(in[184]), .ZN(n756) );
  AND2_X1 U204bar ( .A1(inbar[195]), .A2(inbar[184]), .ZN(n756bar);
  OR2_X1 U205 ( .A1(in[196]), .A2(n755), .ZN(n757) );
  AND2_X1 U205bar ( .A1(inbar[196]), .A2(n755bar), .ZN(n757bar);
  OR2_X1 U206 ( .A1(in[215]), .A2(in[209]), .ZN(n755) );
  AND2_X1 U206bar ( .A1(inbar[215]), .A2(inbar[209]), .ZN(n755bar);
  OR2_X1 U207 ( .A1(n754), .A2(n753), .ZN(n759) );
  AND2_X1 U207bar ( .A1(n754bar), .A2(n753bar), .ZN(n759bar);
  OR2_X1 U208 ( .A1(in[93]), .A2(in[233]), .ZN(n753) );
  AND2_X1 U208bar ( .A1(inbar[93]), .A2(inbar[233]), .ZN(n753bar);
  OR2_X1 U209 ( .A1(in_1), .A2(n752), .ZN(n754) );
  AND2_X1 U209bar ( .A1(in_1bar), .A2(n752bar), .ZN(n754bar);
  OR2_X1 U210 ( .A1(in_69), .A2(in_66), .ZN(n752) );
  AND2_X1 U210bar ( .A1(in_69bar), .A2(in_66bar), .ZN(n752bar);
  OR2_X1 U211 ( .A1(n966), .A2(n751), .ZN(n787) );
  AND2_X1 U211bar ( .A1(n966bar), .A2(n751bar), .ZN(n787bar);
  OR2_X1 U212 ( .A1(in[134]), .A2(n750), .ZN(n751) );
  AND2_X1 U212bar ( .A1(inbar[134]), .A2(n750bar), .ZN(n751bar);
  OR2_X1 U213 ( .A1(n749), .A2(n748), .ZN(n966) );
  AND2_X1 U213bar ( .A1(n749bar), .A2(n748bar), .ZN(n966bar);
  OR2_X1 U214 ( .A1(n747), .A2(n746), .ZN(n748) );
  AND2_X1 U214bar ( .A1(n747bar), .A2(n746bar), .ZN(n748bar);
  OR2_X1 U215 ( .A1(n745), .A2(n744), .ZN(n746) );
  AND2_X1 U215bar ( .A1(n745bar), .A2(n744bar), .ZN(n746bar);
  OR2_X1 U216 ( .A1(in[136]), .A2(in[121]), .ZN(n744) );
  AND2_X1 U216bar ( .A1(inbar[136]), .A2(inbar[121]), .ZN(n744bar);
  OR2_X1 U217 ( .A1(in[186]), .A2(in[174]), .ZN(n745) );
  AND2_X1 U217bar ( .A1(inbar[186]), .A2(inbar[174]), .ZN(n745bar);
  OR2_X1 U218 ( .A1(n743), .A2(n742), .ZN(n747) );
  AND2_X1 U218bar ( .A1(n743bar), .A2(n742bar), .ZN(n747bar);
  OR2_X1 U219 ( .A1(in[198]), .A2(in[197]), .ZN(n742) );
  AND2_X1 U219bar ( .A1(inbar[198]), .A2(inbar[197]), .ZN(n742bar);
  OR2_X1 U220 ( .A1(in[214]), .A2(in[199]), .ZN(n743) );
  AND2_X1 U220bar ( .A1(inbar[214]), .A2(inbar[199]), .ZN(n743bar);
  OR2_X1 U221 ( .A1(n741), .A2(n740), .ZN(n749) );
  AND2_X1 U221bar ( .A1(n741bar), .A2(n740bar), .ZN(n749bar);
  OR2_X1 U222 ( .A1(n739), .A2(n738), .ZN(n740) );
  AND2_X1 U222bar ( .A1(n739bar), .A2(n738bar), .ZN(n740bar);
  OR2_X1 U223 ( .A1(in[231]), .A2(in[220]), .ZN(n738) );
  AND2_X1 U223bar ( .A1(inbar[231]), .A2(inbar[220]), .ZN(n738bar);
  OR2_X1 U224 ( .A1(in_25), .A2(in[245]), .ZN(n739) );
  AND2_X1 U224bar ( .A1(in_25bar), .A2(inbar[245]), .ZN(n739bar);
  OR2_X1 U225 ( .A1(n737), .A2(n736), .ZN(n741) );
  AND2_X1 U225bar ( .A1(n737bar), .A2(n736bar), .ZN(n741bar);
  OR2_X1 U226 ( .A1(in_53), .A2(in_29), .ZN(n736) );
  AND2_X1 U226bar ( .A1(in_53bar), .A2(in_29bar), .ZN(n736bar);
  OR2_X1 U227 ( .A1(in_79), .A2(in_74), .ZN(n737) );
  AND2_X1 U227bar ( .A1(in_79bar), .A2(in_74bar), .ZN(n737bar);
  OR2_X1 U228 ( .A1(n735), .A2(n734), .ZN(n789) );
  AND2_X1 U228bar ( .A1(n735bar), .A2(n734bar), .ZN(n789bar);
  OR2_X1 U229 ( .A1(in[152]), .A2(in[140]), .ZN(n734) );
  AND2_X1 U229bar ( .A1(inbar[152]), .A2(inbar[140]), .ZN(n734bar);
  OR2_X1 U230 ( .A1(in[155]), .A2(n733), .ZN(n735) );
  AND2_X1 U230bar ( .A1(inbar[155]), .A2(n733bar), .ZN(n735bar);
  OR2_X1 U231 ( .A1(in[166]), .A2(in[165]), .ZN(n733) );
  AND2_X1 U231bar ( .A1(inbar[166]), .A2(inbar[165]), .ZN(n733bar);
  OR2_X1 U232 ( .A1(n732), .A2(n731), .ZN(n791) );
  AND2_X1 U232bar ( .A1(n732bar), .A2(n731bar), .ZN(n791bar);
  OR2_X1 U233 ( .A1(n730), .A2(n729), .ZN(n731) );
  AND2_X1 U233bar ( .A1(n730bar), .A2(n729bar), .ZN(n731bar);
  OR2_X1 U234 ( .A1(in[202]), .A2(in[185]), .ZN(n729) );
  AND2_X1 U234bar ( .A1(inbar[202]), .A2(inbar[185]), .ZN(n729bar);
  OR2_X1 U235 ( .A1(in[211]), .A2(n728), .ZN(n730) );
  AND2_X1 U235bar ( .A1(inbar[211]), .A2(n728bar), .ZN(n730bar);
  OR2_X1 U236 ( .A1(in[255]), .A2(in[253]), .ZN(n728) );
  AND2_X1 U236bar ( .A1(inbar[255]), .A2(inbar[253]), .ZN(n728bar);
  OR2_X1 U237 ( .A1(n727), .A2(n726), .ZN(n732) );
  AND2_X1 U237bar ( .A1(n727bar), .A2(n726bar), .ZN(n732bar);
  OR2_X1 U238 ( .A1(in_35), .A2(in_15), .ZN(n726) );
  AND2_X1 U238bar ( .A1(in_35bar), .A2(in_15bar), .ZN(n726bar);
  OR2_X1 U239 ( .A1(in_36), .A2(n725), .ZN(n727) );
  AND2_X1 U239bar ( .A1(in_36bar), .A2(n725bar), .ZN(n727bar);
  OR2_X1 U240 ( .A1(in_48), .A2(in_40), .ZN(n725) );
  AND2_X1 U240bar ( .A1(in_48bar), .A2(in_40bar), .ZN(n725bar);
  OR2_X1 U241 ( .A1(n724), .A2(n723), .ZN(out[1]) );
  AND2_X1 U241bar ( .A1(n724bar), .A2(n723bar), .ZN(outbar[1]);
  OR2_X1 U242 ( .A1(n722), .A2(n721), .ZN(n723) );
  AND2_X1 U242bar ( .A1(n722bar), .A2(n721bar), .ZN(n723bar);
  OR2_X1 U243 ( .A1(n720), .A2(n719), .ZN(n721) );
  AND2_X1 U243bar ( .A1(n720bar), .A2(n719bar), .ZN(n721bar);
  OR2_X1 U244 ( .A1(n921), .A2(n887), .ZN(n719) );
  AND2_X1 U244bar ( .A1(n921bar), .A2(n887bar), .ZN(n719bar);
  OR2_X1 U245 ( .A1(n718), .A2(n717), .ZN(n887) );
  AND2_X1 U245bar ( .A1(n718bar), .A2(n717bar), .ZN(n887bar);
  OR2_X1 U246 ( .A1(n716), .A2(n715), .ZN(n717) );
  AND2_X1 U246bar ( .A1(n716bar), .A2(n715bar), .ZN(n717bar);
  OR2_X1 U247 ( .A1(n714), .A2(n713), .ZN(n715) );
  AND2_X1 U247bar ( .A1(n714bar), .A2(n713bar), .ZN(n715bar);
  OR2_X1 U248 ( .A1(in[116]), .A2(in[110]), .ZN(n713) );
  AND2_X1 U248bar ( .A1(inbar[116]), .A2(inbar[110]), .ZN(n713bar);
  OR2_X1 U249 ( .A1(in[133]), .A2(in[130]), .ZN(n714) );
  AND2_X1 U249bar ( .A1(inbar[133]), .A2(inbar[130]), .ZN(n714bar);
  OR2_X1 U250 ( .A1(n712), .A2(n711), .ZN(n716) );
  AND2_X1 U250bar ( .A1(n712bar), .A2(n711bar), .ZN(n716bar);
  OR2_X1 U251 ( .A1(in[203]), .A2(in[135]), .ZN(n711) );
  AND2_X1 U251bar ( .A1(inbar[203]), .A2(inbar[135]), .ZN(n711bar);
  OR2_X1 U252 ( .A1(in[232]), .A2(in[223]), .ZN(n712) );
  AND2_X1 U252bar ( .A1(inbar[232]), .A2(inbar[223]), .ZN(n712bar);
  OR2_X1 U253 ( .A1(n710), .A2(n709), .ZN(n718) );
  AND2_X1 U253bar ( .A1(n710bar), .A2(n709bar), .ZN(n718bar);
  OR2_X1 U254 ( .A1(n708), .A2(n707), .ZN(n709) );
  AND2_X1 U254bar ( .A1(n708bar), .A2(n707bar), .ZN(n709bar);
  OR2_X1 U255 ( .A1(in[255]), .A2(in[233]), .ZN(n707) );
  AND2_X1 U255bar ( .A1(inbar[255]), .A2(inbar[233]), .ZN(n707bar);
  OR2_X1 U256 ( .A1(in_53), .A2(in_34), .ZN(n708) );
  AND2_X1 U256bar ( .A1(in_53bar), .A2(in_34bar), .ZN(n708bar);
  OR2_X1 U257 ( .A1(n706), .A2(n705), .ZN(n710) );
  AND2_X1 U257bar ( .A1(n706bar), .A2(n705bar), .ZN(n710bar);
  OR2_X1 U258 ( .A1(in_57), .A2(in_55), .ZN(n705) );
  AND2_X1 U258bar ( .A1(in_57bar), .A2(in_55bar), .ZN(n705bar);
  OR2_X1 U259 ( .A1(in_68), .A2(in_67), .ZN(n706) );
  AND2_X1 U259bar ( .A1(in_68bar), .A2(in_67bar), .ZN(n706bar);
  OR2_X1 U260 ( .A1(n704), .A2(n703), .ZN(n921) );
  AND2_X1 U260bar ( .A1(n704bar), .A2(n703bar), .ZN(n921bar);
  OR2_X1 U261 ( .A1(n702), .A2(n701), .ZN(n703) );
  AND2_X1 U261bar ( .A1(n702bar), .A2(n701bar), .ZN(n703bar);
  OR2_X1 U262 ( .A1(n700), .A2(n699), .ZN(n701) );
  AND2_X1 U262bar ( .A1(n700bar), .A2(n699bar), .ZN(n701bar);
  OR2_X1 U263 ( .A1(n944), .A2(n872), .ZN(n699) );
  AND2_X1 U263bar ( .A1(n944bar), .A2(n872bar), .ZN(n699bar);
  OR2_X1 U264 ( .A1(n698), .A2(n697), .ZN(n872) );
  AND2_X1 U264bar ( .A1(n698bar), .A2(n697bar), .ZN(n872bar);
  OR2_X1 U265 ( .A1(n696), .A2(n695), .ZN(n697) );
  AND2_X1 U265bar ( .A1(n696bar), .A2(n695bar), .ZN(n697bar);
  OR2_X1 U266 ( .A1(n694), .A2(n693), .ZN(n695) );
  AND2_X1 U266bar ( .A1(n694bar), .A2(n693bar), .ZN(n695bar);
  OR2_X1 U267 ( .A1(in[121]), .A2(in[102]), .ZN(n693) );
  AND2_X1 U267bar ( .A1(inbar[121]), .A2(inbar[102]), .ZN(n693bar);
  OR2_X1 U268 ( .A1(in[162]), .A2(in[161]), .ZN(n694) );
  AND2_X1 U268bar ( .A1(inbar[162]), .A2(inbar[161]), .ZN(n694bar);
  OR2_X1 U269 ( .A1(n692), .A2(n691), .ZN(n696) );
  AND2_X1 U269bar ( .A1(n692bar), .A2(n691bar), .ZN(n696bar);
  OR2_X1 U270 ( .A1(in[192]), .A2(in[178]), .ZN(n691) );
  AND2_X1 U270bar ( .A1(inbar[192]), .A2(inbar[178]), .ZN(n691bar);
  OR2_X1 U271 ( .A1(in[244]), .A2(in[209]), .ZN(n692) );
  AND2_X1 U271bar ( .A1(inbar[244]), .A2(inbar[209]), .ZN(n692bar);
  OR2_X1 U272 ( .A1(n690), .A2(n689), .ZN(n698) );
  AND2_X1 U272bar ( .A1(n690bar), .A2(n689bar), .ZN(n698bar);
  OR2_X1 U273 ( .A1(n688), .A2(n687), .ZN(n689) );
  AND2_X1 U273bar ( .A1(n688bar), .A2(n687bar), .ZN(n689bar);
  OR2_X1 U274 ( .A1(in[90]), .A2(in[254]), .ZN(n687) );
  AND2_X1 U274bar ( .A1(inbar[90]), .A2(inbar[254]), .ZN(n687bar);
  OR2_X1 U275 ( .A1(in_36), .A2(in_32), .ZN(n688) );
  AND2_X1 U275bar ( .A1(in_36bar), .A2(in_32bar), .ZN(n688bar);
  OR2_X1 U276 ( .A1(n686), .A2(n685), .ZN(n690) );
  AND2_X1 U276bar ( .A1(n686bar), .A2(n685bar), .ZN(n690bar);
  OR2_X1 U277 ( .A1(in_62), .A2(in_37), .ZN(n685) );
  AND2_X1 U277bar ( .A1(in_62bar), .A2(in_37bar), .ZN(n685bar);
  OR2_X1 U278 ( .A1(in_75), .A2(in_73), .ZN(n686) );
  AND2_X1 U278bar ( .A1(in_75bar), .A2(in_73bar), .ZN(n686bar);
  OR2_X1 U279 ( .A1(n684), .A2(n683), .ZN(n944) );
  AND2_X1 U279bar ( .A1(n684bar), .A2(n683bar), .ZN(n944bar);
  OR2_X1 U280 ( .A1(n682), .A2(n681), .ZN(n683) );
  AND2_X1 U280bar ( .A1(n682bar), .A2(n681bar), .ZN(n683bar);
  OR2_X1 U281 ( .A1(n680), .A2(n679), .ZN(n681) );
  AND2_X1 U281bar ( .A1(n680bar), .A2(n679bar), .ZN(n681bar);
  OR2_X1 U282 ( .A1(in[171]), .A2(in[153]), .ZN(n679) );
  AND2_X1 U282bar ( .A1(inbar[171]), .A2(inbar[153]), .ZN(n679bar);
  OR2_X1 U283 ( .A1(in[187]), .A2(in[176]), .ZN(n680) );
  AND2_X1 U283bar ( .A1(inbar[187]), .A2(inbar[176]), .ZN(n680bar);
  OR2_X1 U284 ( .A1(n678), .A2(n677), .ZN(n682) );
  AND2_X1 U284bar ( .A1(n678bar), .A2(n677bar), .ZN(n682bar);
  OR2_X1 U285 ( .A1(in[245]), .A2(in[211]), .ZN(n677) );
  AND2_X1 U285bar ( .A1(inbar[245]), .A2(inbar[211]), .ZN(n677bar);
  OR2_X1 U286 ( .A1(in[97]), .A2(in[88]), .ZN(n678) );
  AND2_X1 U286bar ( .A1(inbar[97]), .A2(inbar[88]), .ZN(n678bar);
  OR2_X1 U287 ( .A1(n676), .A2(n675), .ZN(n684) );
  AND2_X1 U287bar ( .A1(n676bar), .A2(n675bar), .ZN(n684bar);
  OR2_X1 U288 ( .A1(n674), .A2(n673), .ZN(n675) );
  AND2_X1 U288bar ( .A1(n674bar), .A2(n673bar), .ZN(n675bar);
  OR2_X1 U289 ( .A1(in_10), .A2(in_0), .ZN(n673) );
  AND2_X1 U289bar ( .A1(in_10bar), .A2(in_0bar), .ZN(n673bar);
  OR2_X1 U290 ( .A1(in_59), .A2(in_5), .ZN(n674) );
  AND2_X1 U290bar ( .A1(in_59bar), .A2(in_5bar), .ZN(n674bar);
  OR2_X1 U291 ( .A1(n672), .A2(n671), .ZN(n676) );
  AND2_X1 U291bar ( .A1(n672bar), .A2(n671bar), .ZN(n676bar);
  OR2_X1 U292 ( .A1(in_60), .A2(in_6), .ZN(n671) );
  AND2_X1 U292bar ( .A1(in_60bar), .A2(in_6bar), .ZN(n671bar);
  OR2_X1 U293 ( .A1(in_77), .A2(in_69), .ZN(n672) );
  AND2_X1 U293bar ( .A1(in_77bar), .A2(in_69bar), .ZN(n672bar);
  OR2_X1 U294 ( .A1(in[113]), .A2(n864), .ZN(n700) );
  AND2_X1 U294bar ( .A1(inbar[113]), .A2(n864bar), .ZN(n700bar);
  OR2_X1 U295 ( .A1(n670), .A2(n669), .ZN(n864) );
  AND2_X1 U295bar ( .A1(n670bar), .A2(n669bar), .ZN(n864bar);
  OR2_X1 U296 ( .A1(n668), .A2(n667), .ZN(n669) );
  AND2_X1 U296bar ( .A1(n668bar), .A2(n667bar), .ZN(n669bar);
  OR2_X1 U297 ( .A1(n666), .A2(n665), .ZN(n667) );
  AND2_X1 U297bar ( .A1(n666bar), .A2(n665bar), .ZN(n667bar);
  OR2_X1 U298 ( .A1(in[125]), .A2(in[107]), .ZN(n665) );
  AND2_X1 U298bar ( .A1(inbar[125]), .A2(inbar[107]), .ZN(n665bar);
  OR2_X1 U299 ( .A1(in[138]), .A2(in[126]), .ZN(n666) );
  AND2_X1 U299bar ( .A1(inbar[138]), .A2(inbar[126]), .ZN(n666bar);
  OR2_X1 U300 ( .A1(n664), .A2(n663), .ZN(n668) );
  AND2_X1 U300bar ( .A1(n664bar), .A2(n663bar), .ZN(n668bar);
  OR2_X1 U301 ( .A1(in[189]), .A2(in[143]), .ZN(n663) );
  AND2_X1 U301bar ( .A1(inbar[189]), .A2(inbar[143]), .ZN(n663bar);
  OR2_X1 U302 ( .A1(in[99]), .A2(in[214]), .ZN(n664) );
  AND2_X1 U302bar ( .A1(inbar[99]), .A2(inbar[214]), .ZN(n664bar);
  OR2_X1 U303 ( .A1(n662), .A2(n661), .ZN(n670) );
  AND2_X1 U303bar ( .A1(n662bar), .A2(n661bar), .ZN(n670bar);
  OR2_X1 U304 ( .A1(n660), .A2(n659), .ZN(n661) );
  AND2_X1 U304bar ( .A1(n660bar), .A2(n659bar), .ZN(n661bar);
  OR2_X1 U305 ( .A1(in_15), .A2(in_12), .ZN(n659) );
  AND2_X1 U305bar ( .A1(in_15bar), .A2(in_12bar), .ZN(n659bar);
  OR2_X1 U306 ( .A1(in_20), .A2(in_2), .ZN(n660) );
  AND2_X1 U306bar ( .A1(in_20bar), .A2(in_2bar), .ZN(n660bar);
  OR2_X1 U307 ( .A1(n658), .A2(n657), .ZN(n662) );
  AND2_X1 U307bar ( .A1(n658bar), .A2(n657bar), .ZN(n662bar);
  OR2_X1 U308 ( .A1(in_30), .A2(in_3), .ZN(n657) );
  AND2_X1 U308bar ( .A1(in_30bar), .A2(in_3bar), .ZN(n657bar);
  OR2_X1 U309 ( .A1(in_4), .A2(in_38), .ZN(n658) );
  AND2_X1 U309bar ( .A1(in_4bar), .A2(in_38bar), .ZN(n658bar);
  OR2_X1 U310 ( .A1(n656), .A2(n655), .ZN(n702) );
  AND2_X1 U310bar ( .A1(n656bar), .A2(n655bar), .ZN(n702bar);
  OR2_X1 U311 ( .A1(in[148]), .A2(in[137]), .ZN(n655) );
  AND2_X1 U311bar ( .A1(inbar[148]), .A2(inbar[137]), .ZN(n655bar);
  OR2_X1 U312 ( .A1(in[149]), .A2(n654), .ZN(n656) );
  AND2_X1 U312bar ( .A1(inbar[149]), .A2(n654bar), .ZN(n656bar);
  OR2_X1 U313 ( .A1(in[195]), .A2(in[190]), .ZN(n654) );
  AND2_X1 U313bar ( .A1(inbar[195]), .A2(inbar[190]), .ZN(n654bar);
  OR2_X1 U314 ( .A1(n653), .A2(n652), .ZN(n704) );
  AND2_X1 U314bar ( .A1(n653bar), .A2(n652bar), .ZN(n704bar);
  OR2_X1 U315 ( .A1(n651), .A2(n650), .ZN(n652) );
  AND2_X1 U315bar ( .A1(n651bar), .A2(n650bar), .ZN(n652bar);
  OR2_X1 U316 ( .A1(in[98]), .A2(in[197]), .ZN(n650) );
  AND2_X1 U316bar ( .A1(inbar[98]), .A2(inbar[197]), .ZN(n650bar);
  OR2_X1 U317 ( .A1(in_11), .A2(n649), .ZN(n651) );
  AND2_X1 U317bar ( .A1(in_11bar), .A2(n649bar), .ZN(n651bar);
  OR2_X1 U318 ( .A1(in_26), .A2(in_14), .ZN(n649) );
  AND2_X1 U318bar ( .A1(in_26bar), .A2(in_14bar), .ZN(n649bar);
  OR2_X1 U319 ( .A1(n648), .A2(n647), .ZN(n653) );
  AND2_X1 U319bar ( .A1(n648bar), .A2(n647bar), .ZN(n653bar);
  OR2_X1 U320 ( .A1(in_35), .A2(in_27), .ZN(n647) );
  AND2_X1 U320bar ( .A1(in_35bar), .A2(in_27bar), .ZN(n647bar);
  OR2_X1 U321 ( .A1(in_50), .A2(n646), .ZN(n648) );
  AND2_X1 U321bar ( .A1(in_50bar), .A2(n646bar), .ZN(n648bar);
  OR2_X1 U322 ( .A1(in_78), .A2(in_61), .ZN(n646) );
  AND2_X1 U322bar ( .A1(in_78bar), .A2(in_61bar), .ZN(n646bar);
  OR2_X1 U323 ( .A1(n942), .A2(n645), .ZN(n720) );
  AND2_X1 U323bar ( .A1(n942bar), .A2(n645bar), .ZN(n720bar);
  OR2_X1 U324 ( .A1(in[106]), .A2(n863), .ZN(n645) );
  AND2_X1 U324bar ( .A1(inbar[106]), .A2(n863bar), .ZN(n645bar);
  OR2_X1 U325 ( .A1(n644), .A2(n643), .ZN(n863) );
  AND2_X1 U325bar ( .A1(n644bar), .A2(n643bar), .ZN(n863bar);
  OR2_X1 U326 ( .A1(n642), .A2(n641), .ZN(n643) );
  AND2_X1 U326bar ( .A1(n642bar), .A2(n641bar), .ZN(n643bar);
  OR2_X1 U327 ( .A1(n640), .A2(n639), .ZN(n641) );
  AND2_X1 U327bar ( .A1(n640bar), .A2(n639bar), .ZN(n641bar);
  OR2_X1 U328 ( .A1(in[127]), .A2(in[122]), .ZN(n639) );
  AND2_X1 U328bar ( .A1(inbar[127]), .A2(inbar[122]), .ZN(n639bar);
  OR2_X1 U329 ( .A1(in[156]), .A2(in[132]), .ZN(n640) );
  AND2_X1 U329bar ( .A1(inbar[156]), .A2(inbar[132]), .ZN(n640bar);
  OR2_X1 U330 ( .A1(n638), .A2(n637), .ZN(n642) );
  AND2_X1 U330bar ( .A1(n638bar), .A2(n637bar), .ZN(n642bar);
  OR2_X1 U331 ( .A1(in[159]), .A2(in[157]), .ZN(n637) );
  AND2_X1 U331bar ( .A1(inbar[159]), .A2(inbar[157]), .ZN(n637bar);
  OR2_X1 U332 ( .A1(in[185]), .A2(in[169]), .ZN(n638) );
  AND2_X1 U332bar ( .A1(inbar[185]), .A2(inbar[169]), .ZN(n638bar);
  OR2_X1 U333 ( .A1(n636), .A2(n635), .ZN(n644) );
  AND2_X1 U333bar ( .A1(n636bar), .A2(n635bar), .ZN(n644bar);
  OR2_X1 U334 ( .A1(n634), .A2(n633), .ZN(n635) );
  AND2_X1 U334bar ( .A1(n634bar), .A2(n633bar), .ZN(n635bar);
  OR2_X1 U335 ( .A1(in[239]), .A2(in[218]), .ZN(n633) );
  AND2_X1 U335bar ( .A1(inbar[239]), .A2(inbar[218]), .ZN(n633bar);
  OR2_X1 U336 ( .A1(in_13), .A2(in[87]), .ZN(n634) );
  AND2_X1 U336bar ( .A1(in_13bar), .A2(inbar[87]), .ZN(n634bar);
  OR2_X1 U337 ( .A1(n632), .A2(n631), .ZN(n636) );
  AND2_X1 U337bar ( .A1(n632bar), .A2(n631bar), .ZN(n636bar);
  OR2_X1 U338 ( .A1(in_72), .A2(in_70), .ZN(n631) );
  AND2_X1 U338bar ( .A1(in_72bar), .A2(in_70bar), .ZN(n631bar);
  OR2_X1 U339 ( .A1(in_80), .A2(in_74), .ZN(n632) );
  AND2_X1 U339bar ( .A1(in_80bar), .A2(in_74bar), .ZN(n632bar);
  OR2_X1 U340 ( .A1(n630), .A2(n629), .ZN(n942) );
  AND2_X1 U340bar ( .A1(n630bar), .A2(n629bar), .ZN(n942bar);
  OR2_X1 U341 ( .A1(n628), .A2(n627), .ZN(n629) );
  AND2_X1 U341bar ( .A1(n628bar), .A2(n627bar), .ZN(n629bar);
  OR2_X1 U342 ( .A1(n626), .A2(n625), .ZN(n627) );
  AND2_X1 U342bar ( .A1(n626bar), .A2(n625bar), .ZN(n627bar);
  OR2_X1 U343 ( .A1(in[146]), .A2(in[100]), .ZN(n625) );
  AND2_X1 U343bar ( .A1(inbar[146]), .A2(inbar[100]), .ZN(n625bar);
  OR2_X1 U344 ( .A1(in[168]), .A2(in[152]), .ZN(n626) );
  AND2_X1 U344bar ( .A1(inbar[168]), .A2(inbar[152]), .ZN(n626bar);
  OR2_X1 U345 ( .A1(n624), .A2(n623), .ZN(n628) );
  AND2_X1 U345bar ( .A1(n624bar), .A2(n623bar), .ZN(n628bar);
  OR2_X1 U346 ( .A1(in[199]), .A2(in[182]), .ZN(n623) );
  AND2_X1 U346bar ( .A1(inbar[199]), .A2(inbar[182]), .ZN(n623bar);
  OR2_X1 U347 ( .A1(in[236]), .A2(in[204]), .ZN(n624) );
  AND2_X1 U347bar ( .A1(inbar[236]), .A2(inbar[204]), .ZN(n624bar);
  OR2_X1 U348 ( .A1(n622), .A2(n621), .ZN(n630) );
  AND2_X1 U348bar ( .A1(n622bar), .A2(n621bar), .ZN(n630bar);
  OR2_X1 U349 ( .A1(n620), .A2(n619), .ZN(n621) );
  AND2_X1 U349bar ( .A1(n620bar), .A2(n619bar), .ZN(n621bar);
  OR2_X1 U350 ( .A1(in[89]), .A2(in[246]), .ZN(n619) );
  AND2_X1 U350bar ( .A1(inbar[89]), .A2(inbar[246]), .ZN(n619bar);
  OR2_X1 U351 ( .A1(in[95]), .A2(in[92]), .ZN(n620) );
  AND2_X1 U351bar ( .A1(inbar[95]), .A2(inbar[92]), .ZN(n620bar);
  OR2_X1 U352 ( .A1(n618), .A2(n617), .ZN(n622) );
  AND2_X1 U352bar ( .A1(n618bar), .A2(n617bar), .ZN(n622bar);
  OR2_X1 U353 ( .A1(in_22), .A2(in_16), .ZN(n617) );
  AND2_X1 U353bar ( .A1(in_22bar), .A2(in_16bar), .ZN(n617bar);
  OR2_X1 U354 ( .A1(in_51), .A2(in_49), .ZN(n618) );
  AND2_X1 U354bar ( .A1(in_51bar), .A2(in_49bar), .ZN(n618bar);
  OR2_X1 U355 ( .A1(n616), .A2(n615), .ZN(n722) );
  AND2_X1 U355bar ( .A1(n616bar), .A2(n615bar), .ZN(n722bar);
  OR2_X1 U356 ( .A1(in[158]), .A2(in[115]), .ZN(n615) );
  AND2_X1 U356bar ( .A1(inbar[158]), .A2(inbar[115]), .ZN(n615bar);
  OR2_X1 U357 ( .A1(in[163]), .A2(n614), .ZN(n616) );
  AND2_X1 U357bar ( .A1(inbar[163]), .A2(n614bar), .ZN(n616bar);
  OR2_X1 U358 ( .A1(in[206]), .A2(in[165]), .ZN(n614) );
  AND2_X1 U358bar ( .A1(inbar[206]), .A2(inbar[165]), .ZN(n614bar);
  OR2_X1 U359 ( .A1(n613), .A2(n612), .ZN(n724) );
  AND2_X1 U359bar ( .A1(n613bar), .A2(n612bar), .ZN(n724bar);
  OR2_X1 U360 ( .A1(n611), .A2(n610), .ZN(n612) );
  AND2_X1 U360bar ( .A1(n611bar), .A2(n610bar), .ZN(n612bar);
  OR2_X1 U361 ( .A1(in[213]), .A2(in[207]), .ZN(n610) );
  AND2_X1 U361bar ( .A1(inbar[213]), .A2(inbar[207]), .ZN(n610bar);
  OR2_X1 U362 ( .A1(in[215]), .A2(n609), .ZN(n611) );
  AND2_X1 U362bar ( .A1(inbar[215]), .A2(n609bar), .ZN(n611bar);
  OR2_X1 U363 ( .A1(in[230]), .A2(in[220]), .ZN(n609) );
  AND2_X1 U363bar ( .A1(inbar[230]), .A2(inbar[220]), .ZN(n609bar);
  OR2_X1 U364 ( .A1(n608), .A2(n607), .ZN(n613) );
  AND2_X1 U364bar ( .A1(n608bar), .A2(n607bar), .ZN(n613bar);
  OR2_X1 U365 ( .A1(in[251]), .A2(in[234]), .ZN(n607) );
  AND2_X1 U365bar ( .A1(inbar[251]), .A2(inbar[234]), .ZN(n607bar);
  OR2_X1 U366 ( .A1(in_17), .A2(n606), .ZN(n608) );
  AND2_X1 U366bar ( .A1(in_17bar), .A2(n606bar), .ZN(n608bar);
  OR2_X1 U367 ( .A1(in_65), .A2(in_56), .ZN(n606) );
  AND2_X1 U367bar ( .A1(in_65bar), .A2(in_56bar), .ZN(n606bar);
  OR2_X1 U368 ( .A1(n605), .A2(n604), .ZN(out[0]) );
  AND2_X1 U368bar ( .A1(n605bar), .A2(n604bar), .ZN(outbar[0]);
  OR2_X1 U369 ( .A1(n603), .A2(n602), .ZN(n604) );
  AND2_X1 U369bar ( .A1(n603bar), .A2(n602bar), .ZN(n604bar);
  OR2_X1 U370 ( .A1(n601), .A2(n600), .ZN(n602) );
  AND2_X1 U370bar ( .A1(n601bar), .A2(n600bar), .ZN(n602bar);
  OR2_X1 U371 ( .A1(n820), .A2(n785), .ZN(n600) );
  AND2_X1 U371bar ( .A1(n820bar), .A2(n785bar), .ZN(n600bar);
  OR2_X1 U372 ( .A1(n599), .A2(n598), .ZN(n785) );
  AND2_X1 U372bar ( .A1(n599bar), .A2(n598bar), .ZN(n785bar);
  OR2_X1 U373 ( .A1(n597), .A2(n596), .ZN(n598) );
  AND2_X1 U373bar ( .A1(n597bar), .A2(n596bar), .ZN(n598bar);
  OR2_X1 U374 ( .A1(n595), .A2(n594), .ZN(n596) );
  AND2_X1 U374bar ( .A1(n595bar), .A2(n594bar), .ZN(n596bar);
  OR2_X1 U375 ( .A1(in[135]), .A2(in[104]), .ZN(n594) );
  AND2_X1 U375bar ( .A1(inbar[135]), .A2(inbar[104]), .ZN(n594bar);
  OR2_X1 U376 ( .A1(in[188]), .A2(in[178]), .ZN(n595) );
  AND2_X1 U376bar ( .A1(inbar[188]), .A2(inbar[178]), .ZN(n595bar);
  OR2_X1 U377 ( .A1(n593), .A2(n592), .ZN(n597) );
  AND2_X1 U377bar ( .A1(n593bar), .A2(n592bar), .ZN(n597bar);
  OR2_X1 U378 ( .A1(in[217]), .A2(in[194]), .ZN(n592) );
  AND2_X1 U378bar ( .A1(inbar[217]), .A2(inbar[194]), .ZN(n592bar);
  OR2_X1 U379 ( .A1(in[237]), .A2(in[218]), .ZN(n593) );
  AND2_X1 U379bar ( .A1(inbar[237]), .A2(inbar[218]), .ZN(n593bar);
  OR2_X1 U380 ( .A1(n591), .A2(n590), .ZN(n599) );
  AND2_X1 U380bar ( .A1(n591bar), .A2(n590bar), .ZN(n599bar);
  OR2_X1 U381 ( .A1(n589), .A2(n588), .ZN(n590) );
  AND2_X1 U381bar ( .A1(n589bar), .A2(n588bar), .ZN(n590bar);
  OR2_X1 U382 ( .A1(in_2), .A2(in_10), .ZN(n588) );
  AND2_X1 U382bar ( .A1(in_2bar), .A2(in_10bar), .ZN(n588bar);
  OR2_X1 U383 ( .A1(in_47), .A2(in_22), .ZN(n589) );
  AND2_X1 U383bar ( .A1(in_47bar), .A2(in_22bar), .ZN(n589bar);
  OR2_X1 U384 ( .A1(n587), .A2(n586), .ZN(n591) );
  AND2_X1 U384bar ( .A1(n587bar), .A2(n586bar), .ZN(n591bar);
  OR2_X1 U385 ( .A1(in_56), .A2(in_54), .ZN(n586) );
  AND2_X1 U385bar ( .A1(in_56bar), .A2(in_54bar), .ZN(n586bar);
  OR2_X1 U386 ( .A1(in_63), .A2(in_61), .ZN(n587) );
  AND2_X1 U386bar ( .A1(in_63bar), .A2(in_61bar), .ZN(n587bar);
  OR2_X1 U387 ( .A1(n585), .A2(n584), .ZN(n820) );
  AND2_X1 U387bar ( .A1(n585bar), .A2(n584bar), .ZN(n820bar);
  OR2_X1 U388 ( .A1(n583), .A2(n582), .ZN(n584) );
  AND2_X1 U388bar ( .A1(n583bar), .A2(n582bar), .ZN(n584bar);
  OR2_X1 U389 ( .A1(n581), .A2(n580), .ZN(n582) );
  AND2_X1 U389bar ( .A1(n581bar), .A2(n580bar), .ZN(n582bar);
  OR2_X1 U390 ( .A1(in[158]), .A2(in[142]), .ZN(n580) );
  AND2_X1 U390bar ( .A1(inbar[158]), .A2(inbar[142]), .ZN(n580bar);
  OR2_X1 U391 ( .A1(in[175]), .A2(in[164]), .ZN(n581) );
  AND2_X1 U391bar ( .A1(inbar[175]), .A2(inbar[164]), .ZN(n581bar);
  OR2_X1 U392 ( .A1(n579), .A2(n578), .ZN(n583) );
  AND2_X1 U392bar ( .A1(n579bar), .A2(n578bar), .ZN(n583bar);
  OR2_X1 U393 ( .A1(in[228]), .A2(in[204]), .ZN(n578) );
  AND2_X1 U393bar ( .A1(inbar[228]), .A2(inbar[204]), .ZN(n578bar);
  OR2_X1 U394 ( .A1(in[91]), .A2(in[87]), .ZN(n579) );
  AND2_X1 U394bar ( .A1(inbar[91]), .A2(inbar[87]), .ZN(n579bar);
  OR2_X1 U395 ( .A1(n577), .A2(n576), .ZN(n585) );
  AND2_X1 U395bar ( .A1(n577bar), .A2(n576bar), .ZN(n585bar);
  OR2_X1 U396 ( .A1(n575), .A2(n574), .ZN(n576) );
  AND2_X1 U396bar ( .A1(n575bar), .A2(n574bar), .ZN(n576bar);
  OR2_X1 U397 ( .A1(in_21), .A2(in_11), .ZN(n574) );
  AND2_X1 U397bar ( .A1(in_21bar), .A2(in_11bar), .ZN(n574bar);
  OR2_X1 U398 ( .A1(in_5), .A2(in_3), .ZN(n575) );
  AND2_X1 U398bar ( .A1(in_5bar), .A2(in_3bar), .ZN(n575bar);
  OR2_X1 U399 ( .A1(n573), .A2(n572), .ZN(n577) );
  AND2_X1 U399bar ( .A1(n573bar), .A2(n572bar), .ZN(n577bar);
  OR2_X1 U400 ( .A1(in_68), .A2(in_64), .ZN(n572) );
  AND2_X1 U400bar ( .A1(in_68bar), .A2(in_64bar), .ZN(n572bar);
  OR2_X1 U401 ( .A1(in_76), .A2(in_73), .ZN(n573) );
  AND2_X1 U401bar ( .A1(in_76bar), .A2(in_73bar), .ZN(n573bar);
  OR2_X1 U402 ( .A1(n778), .A2(n571), .ZN(n601) );
  AND2_X1 U402bar ( .A1(n778bar), .A2(n571bar), .ZN(n601bar);
  OR2_X1 U403 ( .A1(in[100]), .A2(n965), .ZN(n571) );
  AND2_X1 U403bar ( .A1(inbar[100]), .A2(n965bar), .ZN(n571bar);
  OR2_X1 U404 ( .A1(n570), .A2(n569), .ZN(n965) );
  AND2_X1 U404bar ( .A1(n570bar), .A2(n569bar), .ZN(n965bar);
  OR2_X1 U405 ( .A1(n568), .A2(n567), .ZN(n569) );
  AND2_X1 U405bar ( .A1(n568bar), .A2(n567bar), .ZN(n569bar);
  OR2_X1 U406 ( .A1(n566), .A2(n565), .ZN(n567) );
  AND2_X1 U406bar ( .A1(n566bar), .A2(n565bar), .ZN(n567bar);
  OR2_X1 U407 ( .A1(n817), .A2(n750), .ZN(n565) );
  AND2_X1 U407bar ( .A1(n817bar), .A2(n750bar), .ZN(n565bar);
  OR2_X1 U408 ( .A1(n564), .A2(n563), .ZN(n750) );
  AND2_X1 U408bar ( .A1(n564bar), .A2(n563bar), .ZN(n750bar);
  OR2_X1 U409 ( .A1(n562), .A2(n561), .ZN(n563) );
  AND2_X1 U409bar ( .A1(n562bar), .A2(n561bar), .ZN(n563bar);
  OR2_X1 U410 ( .A1(n560), .A2(n559), .ZN(n561) );
  AND2_X1 U410bar ( .A1(n560bar), .A2(n559bar), .ZN(n561bar);
  OR2_X1 U411 ( .A1(in[119]), .A2(in[103]), .ZN(n559) );
  AND2_X1 U411bar ( .A1(inbar[119]), .A2(inbar[103]), .ZN(n559bar);
  OR2_X1 U412 ( .A1(in[137]), .A2(in[133]), .ZN(n560) );
  AND2_X1 U412bar ( .A1(inbar[137]), .A2(inbar[133]), .ZN(n560bar);
  OR2_X1 U413 ( .A1(n558), .A2(n557), .ZN(n562) );
  AND2_X1 U413bar ( .A1(n558bar), .A2(n557bar), .ZN(n562bar);
  OR2_X1 U414 ( .A1(in[176]), .A2(in[173]), .ZN(n557) );
  AND2_X1 U414bar ( .A1(inbar[176]), .A2(inbar[173]), .ZN(n557bar);
  OR2_X1 U415 ( .A1(in[210]), .A2(in[181]), .ZN(n558) );
  AND2_X1 U415bar ( .A1(inbar[210]), .A2(inbar[181]), .ZN(n558bar);
  OR2_X1 U416 ( .A1(n556), .A2(n555), .ZN(n564) );
  AND2_X1 U416bar ( .A1(n556bar), .A2(n555bar), .ZN(n564bar);
  OR2_X1 U417 ( .A1(n554), .A2(n553), .ZN(n555) );
  AND2_X1 U417bar ( .A1(n554bar), .A2(n553bar), .ZN(n555bar);
  OR2_X1 U418 ( .A1(in_13), .A2(in[234]), .ZN(n553) );
  AND2_X1 U418bar ( .A1(in_13bar), .A2(inbar[234]), .ZN(n553bar);
  OR2_X1 U419 ( .A1(in_38), .A2(in_32), .ZN(n554) );
  AND2_X1 U419bar ( .A1(in_38bar), .A2(in_32bar), .ZN(n554bar);
  OR2_X1 U420 ( .A1(n552), .A2(n551), .ZN(n556) );
  AND2_X1 U420bar ( .A1(n552bar), .A2(n551bar), .ZN(n556bar);
  OR2_X1 U421 ( .A1(in_42), .A2(in_41), .ZN(n551) );
  AND2_X1 U421bar ( .A1(in_42bar), .A2(in_41bar), .ZN(n551bar);
  OR2_X1 U422 ( .A1(in_7), .A2(in_49), .ZN(n552) );
  AND2_X1 U422bar ( .A1(in_7bar), .A2(in_49bar), .ZN(n552bar);
  OR2_X1 U423 ( .A1(n550), .A2(n549), .ZN(n817) );
  AND2_X1 U423bar ( .A1(n550bar), .A2(n549bar), .ZN(n817bar);
  OR2_X1 U424 ( .A1(n548), .A2(n547), .ZN(n549) );
  AND2_X1 U424bar ( .A1(n548bar), .A2(n547bar), .ZN(n549bar);
  OR2_X1 U425 ( .A1(n546), .A2(n545), .ZN(n547) );
  AND2_X1 U425bar ( .A1(n546bar), .A2(n545bar), .ZN(n547bar);
  OR2_X1 U426 ( .A1(in[159]), .A2(in[105]), .ZN(n545) );
  AND2_X1 U426bar ( .A1(inbar[159]), .A2(inbar[105]), .ZN(n545bar);
  OR2_X1 U427 ( .A1(in[206]), .A2(in[183]), .ZN(n546) );
  AND2_X1 U427bar ( .A1(inbar[206]), .A2(inbar[183]), .ZN(n546bar);
  OR2_X1 U428 ( .A1(n544), .A2(n543), .ZN(n548) );
  AND2_X1 U428bar ( .A1(n544bar), .A2(n543bar), .ZN(n548bar);
  OR2_X1 U429 ( .A1(in[229]), .A2(in[219]), .ZN(n543) );
  AND2_X1 U429bar ( .A1(inbar[229]), .A2(inbar[219]), .ZN(n543bar);
  OR2_X1 U430 ( .A1(in[235]), .A2(in[232]), .ZN(n544) );
  AND2_X1 U430bar ( .A1(inbar[235]), .A2(inbar[232]), .ZN(n544bar);
  OR2_X1 U431 ( .A1(n542), .A2(n541), .ZN(n550) );
  AND2_X1 U431bar ( .A1(n542bar), .A2(n541bar), .ZN(n550bar);
  OR2_X1 U432 ( .A1(n540), .A2(n539), .ZN(n541) );
  AND2_X1 U432bar ( .A1(n540bar), .A2(n539bar), .ZN(n541bar);
  OR2_X1 U433 ( .A1(in[249]), .A2(in[242]), .ZN(n539) );
  AND2_X1 U433bar ( .A1(inbar[249]), .A2(inbar[242]), .ZN(n539bar);
  OR2_X1 U434 ( .A1(in[89]), .A2(in[254]), .ZN(n540) );
  AND2_X1 U434bar ( .A1(inbar[89]), .A2(inbar[254]), .ZN(n540bar);
  OR2_X1 U435 ( .A1(n538), .A2(n537), .ZN(n542) );
  AND2_X1 U435bar ( .A1(n538bar), .A2(n537bar), .ZN(n542bar);
  OR2_X1 U436 ( .A1(in_14), .A2(in[99]), .ZN(n537) );
  AND2_X1 U436bar ( .A1(in_14bar), .A2(inbar[99]), .ZN(n537bar);
  OR2_X1 U437 ( .A1(in_60), .A2(in_18), .ZN(n538) );
  AND2_X1 U437bar ( .A1(in_60bar), .A2(in_18bar), .ZN(n538bar);
  OR2_X1 U438 ( .A1(in[113]), .A2(n763), .ZN(n566) );
  AND2_X1 U438bar ( .A1(inbar[113]), .A2(n763bar), .ZN(n566bar);
  OR2_X1 U439 ( .A1(n536), .A2(n535), .ZN(n763) );
  AND2_X1 U439bar ( .A1(n536bar), .A2(n535bar), .ZN(n763bar);
  OR2_X1 U440 ( .A1(n534), .A2(n533), .ZN(n535) );
  AND2_X1 U440bar ( .A1(n534bar), .A2(n533bar), .ZN(n535bar);
  OR2_X1 U441 ( .A1(n532), .A2(n531), .ZN(n533) );
  AND2_X1 U441bar ( .A1(n532bar), .A2(n531bar), .ZN(n533bar);
  OR2_X1 U442 ( .A1(in[115]), .A2(in[110]), .ZN(n531) );
  AND2_X1 U442bar ( .A1(inbar[115]), .A2(inbar[110]), .ZN(n531bar);
  OR2_X1 U443 ( .A1(in[125]), .A2(in[117]), .ZN(n532) );
  AND2_X1 U443bar ( .A1(inbar[125]), .A2(inbar[117]), .ZN(n532bar);
  OR2_X1 U444 ( .A1(n530), .A2(n529), .ZN(n534) );
  AND2_X1 U444bar ( .A1(n530bar), .A2(n529bar), .ZN(n534bar);
  OR2_X1 U445 ( .A1(in[180]), .A2(in[128]), .ZN(n529) );
  AND2_X1 U445bar ( .A1(inbar[180]), .A2(inbar[128]), .ZN(n529bar);
  OR2_X1 U446 ( .A1(in[205]), .A2(in[201]), .ZN(n530) );
  AND2_X1 U446bar ( .A1(inbar[205]), .A2(inbar[201]), .ZN(n530bar);
  OR2_X1 U447 ( .A1(n528), .A2(n527), .ZN(n536) );
  AND2_X1 U447bar ( .A1(n528bar), .A2(n527bar), .ZN(n536bar);
  OR2_X1 U448 ( .A1(n526), .A2(n525), .ZN(n527) );
  AND2_X1 U448bar ( .A1(n526bar), .A2(n525bar), .ZN(n527bar);
  OR2_X1 U449 ( .A1(in[244]), .A2(in[239]), .ZN(n525) );
  AND2_X1 U449bar ( .A1(inbar[244]), .A2(inbar[239]), .ZN(n525bar);
  OR2_X1 U450 ( .A1(in[95]), .A2(in[83]), .ZN(n526) );
  AND2_X1 U450bar ( .A1(inbar[95]), .A2(inbar[83]), .ZN(n526bar);
  OR2_X1 U451 ( .A1(n524), .A2(n523), .ZN(n528) );
  AND2_X1 U451bar ( .A1(n524bar), .A2(n523bar), .ZN(n528bar);
  OR2_X1 U452 ( .A1(in_24), .A2(in[97]), .ZN(n523) );
  AND2_X1 U452bar ( .A1(in_24bar), .A2(inbar[97]), .ZN(n523bar);
  OR2_X1 U453 ( .A1(in_33), .A2(in_27), .ZN(n524) );
  AND2_X1 U453bar ( .A1(in_33bar), .A2(in_27bar), .ZN(n524bar);
  OR2_X1 U454 ( .A1(n522), .A2(n521), .ZN(n568) );
  AND2_X1 U454bar ( .A1(n522bar), .A2(n521bar), .ZN(n568bar);
  OR2_X1 U455 ( .A1(in[145]), .A2(in[126]), .ZN(n521) );
  AND2_X1 U455bar ( .A1(inbar[145]), .A2(inbar[126]), .ZN(n521bar);
  OR2_X1 U456 ( .A1(in[169]), .A2(n520), .ZN(n522) );
  AND2_X1 U456bar ( .A1(inbar[169]), .A2(n520bar), .ZN(n522bar);
  OR2_X1 U457 ( .A1(in[221]), .A2(in[172]), .ZN(n520) );
  AND2_X1 U457bar ( .A1(inbar[221]), .A2(inbar[172]), .ZN(n520bar);
  OR2_X1 U458 ( .A1(n519), .A2(n518), .ZN(n570) );
  AND2_X1 U458bar ( .A1(n519bar), .A2(n518bar), .ZN(n570bar);
  OR2_X1 U459 ( .A1(n517), .A2(n516), .ZN(n518) );
  AND2_X1 U459bar ( .A1(n517bar), .A2(n516bar), .ZN(n518bar);
  OR2_X1 U460 ( .A1(in[241]), .A2(in[224]), .ZN(n516) );
  AND2_X1 U460bar ( .A1(inbar[241]), .A2(inbar[224]), .ZN(n516bar);
  OR2_X1 U461 ( .A1(in[86]), .A2(n515), .ZN(n517) );
  AND2_X1 U461bar ( .A1(inbar[86]), .A2(n515bar), .ZN(n517bar);
  OR2_X1 U462 ( .A1(in_43), .A2(in_34), .ZN(n515) );
  AND2_X1 U462bar ( .A1(in_43bar), .A2(in_34bar), .ZN(n515bar);
  OR2_X1 U463 ( .A1(n514), .A2(n513), .ZN(n519) );
  AND2_X1 U463bar ( .A1(n514bar), .A2(n513bar), .ZN(n519bar);
  OR2_X1 U464 ( .A1(in_65), .A2(in_51), .ZN(n513) );
  AND2_X1 U464bar ( .A1(in_65bar), .A2(in_51bar), .ZN(n513bar);
  OR2_X1 U465 ( .A1(in_75), .A2(n512), .ZN(n514) );
  AND2_X1 U465bar ( .A1(in_75bar), .A2(n512bar), .ZN(n514bar);
  OR2_X1 U466 ( .A1(in_81), .A2(in_77), .ZN(n512) );
  AND2_X1 U466bar ( .A1(in_81bar), .A2(in_77bar), .ZN(n512bar);
  OR2_X1 U467 ( .A1(n511), .A2(n510), .ZN(n778) );
  AND2_X1 U467bar ( .A1(n511bar), .A2(n510bar), .ZN(n778bar);
  OR2_X1 U468 ( .A1(n509), .A2(n508), .ZN(n510) );
  AND2_X1 U468bar ( .A1(n509bar), .A2(n508bar), .ZN(n510bar);
  OR2_X1 U469 ( .A1(n507), .A2(n506), .ZN(n508) );
  AND2_X1 U469bar ( .A1(n507bar), .A2(n506bar), .ZN(n508bar);
  OR2_X1 U470 ( .A1(in[107]), .A2(in[101]), .ZN(n506) );
  AND2_X1 U470bar ( .A1(inbar[107]), .A2(inbar[101]), .ZN(n506bar);
  OR2_X1 U471 ( .A1(in[139]), .A2(in[132]), .ZN(n507) );
  AND2_X1 U471bar ( .A1(inbar[139]), .A2(inbar[132]), .ZN(n507bar);
  OR2_X1 U472 ( .A1(n505), .A2(n504), .ZN(n509) );
  AND2_X1 U472bar ( .A1(n505bar), .A2(n504bar), .ZN(n509bar);
  OR2_X1 U473 ( .A1(in[146]), .A2(in[141]), .ZN(n504) );
  AND2_X1 U473bar ( .A1(inbar[146]), .A2(inbar[141]), .ZN(n504bar);
  OR2_X1 U474 ( .A1(in[203]), .A2(in[179]), .ZN(n505) );
  AND2_X1 U474bar ( .A1(inbar[203]), .A2(inbar[179]), .ZN(n505bar);
  OR2_X1 U475 ( .A1(n503), .A2(n502), .ZN(n511) );
  AND2_X1 U475bar ( .A1(n503bar), .A2(n502bar), .ZN(n511bar);
  OR2_X1 U476 ( .A1(n501), .A2(n500), .ZN(n502) );
  AND2_X1 U476bar ( .A1(n501bar), .A2(n500bar), .ZN(n502bar);
  OR2_X1 U477 ( .A1(in[243]), .A2(in[222]), .ZN(n500) );
  AND2_X1 U477bar ( .A1(inbar[243]), .A2(inbar[222]), .ZN(n500bar);
  OR2_X1 U478 ( .A1(in[251]), .A2(in[250]), .ZN(n501) );
  AND2_X1 U478bar ( .A1(inbar[251]), .A2(inbar[250]), .ZN(n501bar);
  OR2_X1 U479 ( .A1(n499), .A2(n498), .ZN(n503) );
  AND2_X1 U479bar ( .A1(n499bar), .A2(n498bar), .ZN(n503bar);
  OR2_X1 U480 ( .A1(in_37), .A2(in_19), .ZN(n498) );
  AND2_X1 U480bar ( .A1(in_37bar), .A2(in_19bar), .ZN(n498bar);
  OR2_X1 U481 ( .A1(in_78), .A2(in_6), .ZN(n499) );
  AND2_X1 U481bar ( .A1(in_78bar), .A2(in_6bar), .ZN(n499bar);
  OR2_X1 U482 ( .A1(n497), .A2(n496), .ZN(n603) );
  AND2_X1 U482bar ( .A1(n497bar), .A2(n496bar), .ZN(n603bar);
  OR2_X1 U483 ( .A1(in[112]), .A2(in[102]), .ZN(n496) );
  AND2_X1 U483bar ( .A1(inbar[112]), .A2(inbar[102]), .ZN(n496bar);
  OR2_X1 U484 ( .A1(in[123]), .A2(n495), .ZN(n497) );
  AND2_X1 U484bar ( .A1(inbar[123]), .A2(n495bar), .ZN(n497bar);
  OR2_X1 U485 ( .A1(in[143]), .A2(in[130]), .ZN(n495) );
  AND2_X1 U485bar ( .A1(inbar[143]), .A2(inbar[130]), .ZN(n495bar);
  OR2_X1 U486 ( .A1(n494), .A2(n493), .ZN(n605) );
  AND2_X1 U486bar ( .A1(n494bar), .A2(n493bar), .ZN(n605bar);
  OR2_X1 U487 ( .A1(n492), .A2(n491), .ZN(n493) );
  AND2_X1 U487bar ( .A1(n492bar), .A2(n491bar), .ZN(n493bar);
  OR2_X1 U488 ( .A1(in[216]), .A2(in[213]), .ZN(n491) );
  AND2_X1 U488bar ( .A1(inbar[216]), .A2(inbar[213]), .ZN(n491bar);
  OR2_X1 U489 ( .A1(in[227]), .A2(n490), .ZN(n492) );
  AND2_X1 U489bar ( .A1(inbar[227]), .A2(n490bar), .ZN(n492bar);
  OR2_X1 U490 ( .A1(in_0), .A2(in[248]), .ZN(n490) );
  AND2_X1 U490bar ( .A1(in_0bar), .A2(inbar[248]), .ZN(n490bar);
  OR2_X1 U491 ( .A1(n489), .A2(n488), .ZN(n494) );
  AND2_X1 U491bar ( .A1(n489bar), .A2(n488bar), .ZN(n494bar);
  OR2_X1 U492 ( .A1(in_46), .A2(in_44), .ZN(n488) );
  AND2_X1 U492bar ( .A1(in_46bar), .A2(in_44bar), .ZN(n488bar);
  OR2_X1 U493 ( .A1(in_50), .A2(n487), .ZN(n489) );
  AND2_X1 U493bar ( .A1(in_50bar), .A2(n487bar), .ZN(n489bar);
  OR2_X1 U494 ( .A1(in_9), .A2(in_80), .ZN(n487) );
  AND2_X1 U494bar ( .A1(in_9bar), .A2(in_80bar), .ZN(n487bar);
endmodule




module sBox_10 ( in, out );
  input [7:0] in;
  //input_done

  output [7:0] out;
  //output_done

  wire   [255:0] decodeOut;
  //wire_done

  decode_10 dec ( .in(in), .out(decodeOut) );
  encode_10 enc ( .in(decodeOut), .out(out) );
endmodule


module CD2_41 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_42 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_43 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_44 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD4_21 ( a, b, y );
  input [3:0] a;
  input [3:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  //input_done

  output [15:0] y;
  reg [15:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]);
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]);
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]);
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]);
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]);
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]);
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]);
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]);
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]);
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]);
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]);
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]);
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]);
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]);
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]);
endmodule




module CD4_22 ( a, b, y );
  input [3:0] a;
  input [3:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  //input_done

  output [15:0] y;
  reg [15:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]);
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]);
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]);
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]);
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]);
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]);
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]);
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]);
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]);
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]);
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]);
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]);
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]);
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]);
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]);
endmodule




module CD16_11 ( a, b, y );
  input [15:0] a;
  input [15:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign abar[8] = ~a[8];
  assign abar[9] = ~a[9];
  assign abar[10] = ~a[10];
  assign abar[11] = ~a[11];
  assign abar[12] = ~a[12];
  assign abar[13] = ~a[13];
  assign abar[14] = ~a[14];
  assign abar[15] = ~a[15];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign bbar[8] = ~b[8];
  assign bbar[9] = ~b[9];
  assign bbar[10] = ~b[10];
  assign bbar[11] = ~b[11];
  assign bbar[12] = ~b[12];
  assign bbar[13] = ~b[13];
  assign bbar[14] = ~b[14];
  assign bbar[15] = ~b[15];
  //input_done

  output [255:0] y;
  reg [255:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[9]), .A2(a[0]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[9]), .A2(abar[0]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[3]), .A2(a[6]), .ZN(y[99]) );
  OR2_X1 U2bar ( .A1(bbar[3]), .A2(abar[6]), .ZN(ybar[99]);
  AND2_X1 U3 ( .A1(b[2]), .A2(a[6]), .ZN(y[98]) );
  OR2_X1 U3bar ( .A1(bbar[2]), .A2(abar[6]), .ZN(ybar[98]);
  AND2_X1 U4 ( .A1(b[1]), .A2(a[6]), .ZN(y[97]) );
  OR2_X1 U4bar ( .A1(bbar[1]), .A2(abar[6]), .ZN(ybar[97]);
  AND2_X1 U5 ( .A1(b[0]), .A2(a[6]), .ZN(y[96]) );
  OR2_X1 U5bar ( .A1(bbar[0]), .A2(abar[6]), .ZN(ybar[96]);
  AND2_X1 U6 ( .A1(b[15]), .A2(a[5]), .ZN(y[95]) );
  OR2_X1 U6bar ( .A1(bbar[15]), .A2(abar[5]), .ZN(ybar[95]);
  AND2_X1 U7 ( .A1(b[14]), .A2(a[5]), .ZN(y[94]) );
  OR2_X1 U7bar ( .A1(bbar[14]), .A2(abar[5]), .ZN(ybar[94]);
  AND2_X1 U8 ( .A1(b[13]), .A2(a[5]), .ZN(y[93]) );
  OR2_X1 U8bar ( .A1(bbar[13]), .A2(abar[5]), .ZN(ybar[93]);
  AND2_X1 U9 ( .A1(b[12]), .A2(a[5]), .ZN(y[92]) );
  OR2_X1 U9bar ( .A1(bbar[12]), .A2(abar[5]), .ZN(ybar[92]);
  AND2_X1 U10 ( .A1(b[11]), .A2(a[5]), .ZN(y[91]) );
  OR2_X1 U10bar ( .A1(bbar[11]), .A2(abar[5]), .ZN(ybar[91]);
  AND2_X1 U11 ( .A1(b[10]), .A2(a[5]), .ZN(y[90]) );
  OR2_X1 U11bar ( .A1(bbar[10]), .A2(abar[5]), .ZN(ybar[90]);
  AND2_X1 U12 ( .A1(b[8]), .A2(a[0]), .ZN(y[8]) );
  OR2_X1 U12bar ( .A1(bbar[8]), .A2(abar[0]), .ZN(ybar[8]);
  AND2_X1 U13 ( .A1(a[5]), .A2(b[9]), .ZN(y[89]) );
  OR2_X1 U13bar ( .A1(abar[5]), .A2(bbar[9]), .ZN(ybar[89]);
  AND2_X1 U14 ( .A1(b[8]), .A2(a[5]), .ZN(y[88]) );
  OR2_X1 U14bar ( .A1(bbar[8]), .A2(abar[5]), .ZN(ybar[88]);
  AND2_X1 U15 ( .A1(b[7]), .A2(a[5]), .ZN(y[87]) );
  OR2_X1 U15bar ( .A1(bbar[7]), .A2(abar[5]), .ZN(ybar[87]);
  AND2_X1 U16 ( .A1(b[6]), .A2(a[5]), .ZN(y[86]) );
  OR2_X1 U16bar ( .A1(bbar[6]), .A2(abar[5]), .ZN(ybar[86]);
  AND2_X1 U17 ( .A1(b[5]), .A2(a[5]), .ZN(y[85]) );
  OR2_X1 U17bar ( .A1(bbar[5]), .A2(abar[5]), .ZN(ybar[85]);
  AND2_X1 U18 ( .A1(b[4]), .A2(a[5]), .ZN(y[84]) );
  OR2_X1 U18bar ( .A1(bbar[4]), .A2(abar[5]), .ZN(ybar[84]);
  AND2_X1 U19 ( .A1(a[5]), .A2(b[3]), .ZN(y[83]) );
  OR2_X1 U19bar ( .A1(abar[5]), .A2(bbar[3]), .ZN(ybar[83]);
  AND2_X1 U20 ( .A1(a[5]), .A2(b[2]), .ZN(y[82]) );
  OR2_X1 U20bar ( .A1(abar[5]), .A2(bbar[2]), .ZN(ybar[82]);
  AND2_X1 U21 ( .A1(a[5]), .A2(b[1]), .ZN(y[81]) );
  OR2_X1 U21bar ( .A1(abar[5]), .A2(bbar[1]), .ZN(ybar[81]);
  AND2_X1 U22 ( .A1(a[5]), .A2(b[0]), .ZN(y[80]) );
  OR2_X1 U22bar ( .A1(abar[5]), .A2(bbar[0]), .ZN(ybar[80]);
  AND2_X1 U23 ( .A1(b[7]), .A2(a[0]), .ZN(y[7]) );
  OR2_X1 U23bar ( .A1(bbar[7]), .A2(abar[0]), .ZN(ybar[7]);
  AND2_X1 U24 ( .A1(a[4]), .A2(b[15]), .ZN(y[79]) );
  OR2_X1 U24bar ( .A1(abar[4]), .A2(bbar[15]), .ZN(ybar[79]);
  AND2_X1 U25 ( .A1(a[4]), .A2(b[14]), .ZN(y[78]) );
  OR2_X1 U25bar ( .A1(abar[4]), .A2(bbar[14]), .ZN(ybar[78]);
  AND2_X1 U26 ( .A1(a[4]), .A2(b[13]), .ZN(y[77]) );
  OR2_X1 U26bar ( .A1(abar[4]), .A2(bbar[13]), .ZN(ybar[77]);
  AND2_X1 U27 ( .A1(a[4]), .A2(b[12]), .ZN(y[76]) );
  OR2_X1 U27bar ( .A1(abar[4]), .A2(bbar[12]), .ZN(ybar[76]);
  AND2_X1 U28 ( .A1(a[4]), .A2(b[11]), .ZN(y[75]) );
  OR2_X1 U28bar ( .A1(abar[4]), .A2(bbar[11]), .ZN(ybar[75]);
  AND2_X1 U29 ( .A1(a[4]), .A2(b[10]), .ZN(y[74]) );
  OR2_X1 U29bar ( .A1(abar[4]), .A2(bbar[10]), .ZN(ybar[74]);
  AND2_X1 U30 ( .A1(a[4]), .A2(b[9]), .ZN(y[73]) );
  OR2_X1 U30bar ( .A1(abar[4]), .A2(bbar[9]), .ZN(ybar[73]);
  AND2_X1 U31 ( .A1(a[4]), .A2(b[8]), .ZN(y[72]) );
  OR2_X1 U31bar ( .A1(abar[4]), .A2(bbar[8]), .ZN(ybar[72]);
  AND2_X1 U32 ( .A1(a[4]), .A2(b[7]), .ZN(y[71]) );
  OR2_X1 U32bar ( .A1(abar[4]), .A2(bbar[7]), .ZN(ybar[71]);
  AND2_X1 U33 ( .A1(a[4]), .A2(b[6]), .ZN(y[70]) );
  OR2_X1 U33bar ( .A1(abar[4]), .A2(bbar[6]), .ZN(ybar[70]);
  AND2_X1 U34 ( .A1(b[6]), .A2(a[0]), .ZN(y[6]) );
  OR2_X1 U34bar ( .A1(bbar[6]), .A2(abar[0]), .ZN(ybar[6]);
  AND2_X1 U35 ( .A1(a[4]), .A2(b[5]), .ZN(y[69]) );
  OR2_X1 U35bar ( .A1(abar[4]), .A2(bbar[5]), .ZN(ybar[69]);
  AND2_X1 U36 ( .A1(a[4]), .A2(b[4]), .ZN(y[68]) );
  OR2_X1 U36bar ( .A1(abar[4]), .A2(bbar[4]), .ZN(ybar[68]);
  AND2_X1 U37 ( .A1(a[4]), .A2(b[3]), .ZN(y[67]) );
  OR2_X1 U37bar ( .A1(abar[4]), .A2(bbar[3]), .ZN(ybar[67]);
  AND2_X1 U38 ( .A1(a[4]), .A2(b[2]), .ZN(y[66]) );
  OR2_X1 U38bar ( .A1(abar[4]), .A2(bbar[2]), .ZN(ybar[66]);
  AND2_X1 U39 ( .A1(a[4]), .A2(b[1]), .ZN(y[65]) );
  OR2_X1 U39bar ( .A1(abar[4]), .A2(bbar[1]), .ZN(ybar[65]);
  AND2_X1 U40 ( .A1(a[4]), .A2(b[0]), .ZN(y[64]) );
  OR2_X1 U40bar ( .A1(abar[4]), .A2(bbar[0]), .ZN(ybar[64]);
  AND2_X1 U41 ( .A1(a[3]), .A2(b[15]), .ZN(y[63]) );
  OR2_X1 U41bar ( .A1(abar[3]), .A2(bbar[15]), .ZN(ybar[63]);
  AND2_X1 U42 ( .A1(a[3]), .A2(b[14]), .ZN(y[62]) );
  OR2_X1 U42bar ( .A1(abar[3]), .A2(bbar[14]), .ZN(ybar[62]);
  AND2_X1 U43 ( .A1(a[3]), .A2(b[13]), .ZN(y[61]) );
  OR2_X1 U43bar ( .A1(abar[3]), .A2(bbar[13]), .ZN(ybar[61]);
  AND2_X1 U44 ( .A1(a[3]), .A2(b[12]), .ZN(y[60]) );
  OR2_X1 U44bar ( .A1(abar[3]), .A2(bbar[12]), .ZN(ybar[60]);
  AND2_X1 U45 ( .A1(b[5]), .A2(a[0]), .ZN(y[5]) );
  OR2_X1 U45bar ( .A1(bbar[5]), .A2(abar[0]), .ZN(ybar[5]);
  AND2_X1 U46 ( .A1(a[3]), .A2(b[11]), .ZN(y[59]) );
  OR2_X1 U46bar ( .A1(abar[3]), .A2(bbar[11]), .ZN(ybar[59]);
  AND2_X1 U47 ( .A1(a[3]), .A2(b[10]), .ZN(y[58]) );
  OR2_X1 U47bar ( .A1(abar[3]), .A2(bbar[10]), .ZN(ybar[58]);
  AND2_X1 U48 ( .A1(a[3]), .A2(b[9]), .ZN(y[57]) );
  OR2_X1 U48bar ( .A1(abar[3]), .A2(bbar[9]), .ZN(ybar[57]);
  AND2_X1 U49 ( .A1(a[3]), .A2(b[8]), .ZN(y[56]) );
  OR2_X1 U49bar ( .A1(abar[3]), .A2(bbar[8]), .ZN(ybar[56]);
  AND2_X1 U50 ( .A1(a[3]), .A2(b[7]), .ZN(y[55]) );
  OR2_X1 U50bar ( .A1(abar[3]), .A2(bbar[7]), .ZN(ybar[55]);
  AND2_X1 U51 ( .A1(a[3]), .A2(b[6]), .ZN(y[54]) );
  OR2_X1 U51bar ( .A1(abar[3]), .A2(bbar[6]), .ZN(ybar[54]);
  AND2_X1 U52 ( .A1(a[3]), .A2(b[5]), .ZN(y[53]) );
  OR2_X1 U52bar ( .A1(abar[3]), .A2(bbar[5]), .ZN(ybar[53]);
  AND2_X1 U53 ( .A1(a[3]), .A2(b[4]), .ZN(y[52]) );
  OR2_X1 U53bar ( .A1(abar[3]), .A2(bbar[4]), .ZN(ybar[52]);
  AND2_X1 U54 ( .A1(a[3]), .A2(b[3]), .ZN(y[51]) );
  OR2_X1 U54bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[51]);
  AND2_X1 U55 ( .A1(a[3]), .A2(b[2]), .ZN(y[50]) );
  OR2_X1 U55bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[50]);
  AND2_X1 U56 ( .A1(b[4]), .A2(a[0]), .ZN(y[4]) );
  OR2_X1 U56bar ( .A1(bbar[4]), .A2(abar[0]), .ZN(ybar[4]);
  AND2_X1 U57 ( .A1(a[3]), .A2(b[1]), .ZN(y[49]) );
  OR2_X1 U57bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[49]);
  AND2_X1 U58 ( .A1(a[3]), .A2(b[0]), .ZN(y[48]) );
  OR2_X1 U58bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[48]);
  AND2_X1 U59 ( .A1(a[2]), .A2(b[15]), .ZN(y[47]) );
  OR2_X1 U59bar ( .A1(abar[2]), .A2(bbar[15]), .ZN(ybar[47]);
  AND2_X1 U60 ( .A1(a[2]), .A2(b[14]), .ZN(y[46]) );
  OR2_X1 U60bar ( .A1(abar[2]), .A2(bbar[14]), .ZN(ybar[46]);
  AND2_X1 U61 ( .A1(a[2]), .A2(b[13]), .ZN(y[45]) );
  OR2_X1 U61bar ( .A1(abar[2]), .A2(bbar[13]), .ZN(ybar[45]);
  AND2_X1 U62 ( .A1(a[2]), .A2(b[12]), .ZN(y[44]) );
  OR2_X1 U62bar ( .A1(abar[2]), .A2(bbar[12]), .ZN(ybar[44]);
  AND2_X1 U63 ( .A1(a[2]), .A2(b[11]), .ZN(y[43]) );
  OR2_X1 U63bar ( .A1(abar[2]), .A2(bbar[11]), .ZN(ybar[43]);
  AND2_X1 U64 ( .A1(a[2]), .A2(b[10]), .ZN(y[42]) );
  OR2_X1 U64bar ( .A1(abar[2]), .A2(bbar[10]), .ZN(ybar[42]);
  AND2_X1 U65 ( .A1(a[2]), .A2(b[9]), .ZN(y[41]) );
  OR2_X1 U65bar ( .A1(abar[2]), .A2(bbar[9]), .ZN(ybar[41]);
  AND2_X1 U66 ( .A1(a[2]), .A2(b[8]), .ZN(y[40]) );
  OR2_X1 U66bar ( .A1(abar[2]), .A2(bbar[8]), .ZN(ybar[40]);
  AND2_X1 U67 ( .A1(b[3]), .A2(a[0]), .ZN(y[3]) );
  OR2_X1 U67bar ( .A1(bbar[3]), .A2(abar[0]), .ZN(ybar[3]);
  AND2_X1 U68 ( .A1(a[2]), .A2(b[7]), .ZN(y[39]) );
  OR2_X1 U68bar ( .A1(abar[2]), .A2(bbar[7]), .ZN(ybar[39]);
  AND2_X1 U69 ( .A1(a[2]), .A2(b[6]), .ZN(y[38]) );
  OR2_X1 U69bar ( .A1(abar[2]), .A2(bbar[6]), .ZN(ybar[38]);
  AND2_X1 U70 ( .A1(a[2]), .A2(b[5]), .ZN(y[37]) );
  OR2_X1 U70bar ( .A1(abar[2]), .A2(bbar[5]), .ZN(ybar[37]);
  AND2_X1 U71 ( .A1(a[2]), .A2(b[4]), .ZN(y[36]) );
  OR2_X1 U71bar ( .A1(abar[2]), .A2(bbar[4]), .ZN(ybar[36]);
  AND2_X1 U72 ( .A1(a[2]), .A2(b[3]), .ZN(y[35]) );
  OR2_X1 U72bar ( .A1(abar[2]), .A2(bbar[3]), .ZN(ybar[35]);
  AND2_X1 U73 ( .A1(a[2]), .A2(b[2]), .ZN(y[34]) );
  OR2_X1 U73bar ( .A1(abar[2]), .A2(bbar[2]), .ZN(ybar[34]);
  AND2_X1 U74 ( .A1(a[2]), .A2(b[1]), .ZN(y[33]) );
  OR2_X1 U74bar ( .A1(abar[2]), .A2(bbar[1]), .ZN(ybar[33]);
  AND2_X1 U75 ( .A1(a[2]), .A2(b[0]), .ZN(y[32]) );
  OR2_X1 U75bar ( .A1(abar[2]), .A2(bbar[0]), .ZN(ybar[32]);
  AND2_X1 U76 ( .A1(a[1]), .A2(b[15]), .ZN(y[31]) );
  OR2_X1 U76bar ( .A1(abar[1]), .A2(bbar[15]), .ZN(ybar[31]);
  AND2_X1 U77 ( .A1(a[1]), .A2(b[14]), .ZN(y[30]) );
  OR2_X1 U77bar ( .A1(abar[1]), .A2(bbar[14]), .ZN(ybar[30]);
  AND2_X1 U78 ( .A1(b[2]), .A2(a[0]), .ZN(y[2]) );
  OR2_X1 U78bar ( .A1(bbar[2]), .A2(abar[0]), .ZN(ybar[2]);
  AND2_X1 U79 ( .A1(a[1]), .A2(b[13]), .ZN(y[29]) );
  OR2_X1 U79bar ( .A1(abar[1]), .A2(bbar[13]), .ZN(ybar[29]);
  AND2_X1 U80 ( .A1(a[1]), .A2(b[12]), .ZN(y[28]) );
  OR2_X1 U80bar ( .A1(abar[1]), .A2(bbar[12]), .ZN(ybar[28]);
  AND2_X1 U81 ( .A1(a[1]), .A2(b[11]), .ZN(y[27]) );
  OR2_X1 U81bar ( .A1(abar[1]), .A2(bbar[11]), .ZN(ybar[27]);
  AND2_X1 U82 ( .A1(a[1]), .A2(b[10]), .ZN(y[26]) );
  OR2_X1 U82bar ( .A1(abar[1]), .A2(bbar[10]), .ZN(ybar[26]);
  AND2_X1 U83 ( .A1(a[1]), .A2(b[9]), .ZN(y[25]) );
  OR2_X1 U83bar ( .A1(abar[1]), .A2(bbar[9]), .ZN(ybar[25]);
  AND2_X1 U84 ( .A1(a[15]), .A2(b[15]), .ZN(y[255]) );
  OR2_X1 U84bar ( .A1(abar[15]), .A2(bbar[15]), .ZN(ybar[255]);
  AND2_X1 U85 ( .A1(a[15]), .A2(b[14]), .ZN(y[254]) );
  OR2_X1 U85bar ( .A1(abar[15]), .A2(bbar[14]), .ZN(ybar[254]);
  AND2_X1 U86 ( .A1(a[15]), .A2(b[13]), .ZN(y[253]) );
  OR2_X1 U86bar ( .A1(abar[15]), .A2(bbar[13]), .ZN(ybar[253]);
  AND2_X1 U87 ( .A1(a[15]), .A2(b[12]), .ZN(y[252]) );
  OR2_X1 U87bar ( .A1(abar[15]), .A2(bbar[12]), .ZN(ybar[252]);
  AND2_X1 U88 ( .A1(a[15]), .A2(b[11]), .ZN(y[251]) );
  OR2_X1 U88bar ( .A1(abar[15]), .A2(bbar[11]), .ZN(ybar[251]);
  AND2_X1 U89 ( .A1(a[15]), .A2(b[10]), .ZN(y[250]) );
  OR2_X1 U89bar ( .A1(abar[15]), .A2(bbar[10]), .ZN(ybar[250]);
  AND2_X1 U90 ( .A1(a[1]), .A2(b[8]), .ZN(y[24]) );
  OR2_X1 U90bar ( .A1(abar[1]), .A2(bbar[8]), .ZN(ybar[24]);
  AND2_X1 U91 ( .A1(a[15]), .A2(b[9]), .ZN(y[249]) );
  OR2_X1 U91bar ( .A1(abar[15]), .A2(bbar[9]), .ZN(ybar[249]);
  AND2_X1 U92 ( .A1(a[15]), .A2(b[8]), .ZN(y[248]) );
  OR2_X1 U92bar ( .A1(abar[15]), .A2(bbar[8]), .ZN(ybar[248]);
  AND2_X1 U93 ( .A1(a[15]), .A2(b[7]), .ZN(y[247]) );
  OR2_X1 U93bar ( .A1(abar[15]), .A2(bbar[7]), .ZN(ybar[247]);
  AND2_X1 U94 ( .A1(a[15]), .A2(b[6]), .ZN(y[246]) );
  OR2_X1 U94bar ( .A1(abar[15]), .A2(bbar[6]), .ZN(ybar[246]);
  AND2_X1 U95 ( .A1(a[15]), .A2(b[5]), .ZN(y[245]) );
  OR2_X1 U95bar ( .A1(abar[15]), .A2(bbar[5]), .ZN(ybar[245]);
  AND2_X1 U96 ( .A1(a[15]), .A2(b[4]), .ZN(y[244]) );
  OR2_X1 U96bar ( .A1(abar[15]), .A2(bbar[4]), .ZN(ybar[244]);
  AND2_X1 U97 ( .A1(a[15]), .A2(b[3]), .ZN(y[243]) );
  OR2_X1 U97bar ( .A1(abar[15]), .A2(bbar[3]), .ZN(ybar[243]);
  AND2_X1 U98 ( .A1(a[15]), .A2(b[2]), .ZN(y[242]) );
  OR2_X1 U98bar ( .A1(abar[15]), .A2(bbar[2]), .ZN(ybar[242]);
  AND2_X1 U99 ( .A1(a[15]), .A2(b[1]), .ZN(y[241]) );
  OR2_X1 U99bar ( .A1(abar[15]), .A2(bbar[1]), .ZN(ybar[241]);
  AND2_X1 U100 ( .A1(a[15]), .A2(b[0]), .ZN(y[240]) );
  OR2_X1 U100bar ( .A1(abar[15]), .A2(bbar[0]), .ZN(ybar[240]);
  AND2_X1 U101 ( .A1(a[1]), .A2(b[7]), .ZN(y[23]) );
  OR2_X1 U101bar ( .A1(abar[1]), .A2(bbar[7]), .ZN(ybar[23]);
  AND2_X1 U102 ( .A1(a[14]), .A2(b[15]), .ZN(y[239]) );
  OR2_X1 U102bar ( .A1(abar[14]), .A2(bbar[15]), .ZN(ybar[239]);
  AND2_X1 U103 ( .A1(a[14]), .A2(b[14]), .ZN(y[238]) );
  OR2_X1 U103bar ( .A1(abar[14]), .A2(bbar[14]), .ZN(ybar[238]);
  AND2_X1 U104 ( .A1(a[14]), .A2(b[13]), .ZN(y[237]) );
  OR2_X1 U104bar ( .A1(abar[14]), .A2(bbar[13]), .ZN(ybar[237]);
  AND2_X1 U105 ( .A1(a[14]), .A2(b[12]), .ZN(y[236]) );
  OR2_X1 U105bar ( .A1(abar[14]), .A2(bbar[12]), .ZN(ybar[236]);
  AND2_X1 U106 ( .A1(a[14]), .A2(b[11]), .ZN(y[235]) );
  OR2_X1 U106bar ( .A1(abar[14]), .A2(bbar[11]), .ZN(ybar[235]);
  AND2_X1 U107 ( .A1(a[14]), .A2(b[10]), .ZN(y[234]) );
  OR2_X1 U107bar ( .A1(abar[14]), .A2(bbar[10]), .ZN(ybar[234]);
  AND2_X1 U108 ( .A1(a[14]), .A2(b[9]), .ZN(y[233]) );
  OR2_X1 U108bar ( .A1(abar[14]), .A2(bbar[9]), .ZN(ybar[233]);
  AND2_X1 U109 ( .A1(a[14]), .A2(b[8]), .ZN(y[232]) );
  OR2_X1 U109bar ( .A1(abar[14]), .A2(bbar[8]), .ZN(ybar[232]);
  AND2_X1 U110 ( .A1(a[14]), .A2(b[7]), .ZN(y[231]) );
  OR2_X1 U110bar ( .A1(abar[14]), .A2(bbar[7]), .ZN(ybar[231]);
  AND2_X1 U111 ( .A1(a[14]), .A2(b[6]), .ZN(y[230]) );
  OR2_X1 U111bar ( .A1(abar[14]), .A2(bbar[6]), .ZN(ybar[230]);
  AND2_X1 U112 ( .A1(a[1]), .A2(b[6]), .ZN(y[22]) );
  OR2_X1 U112bar ( .A1(abar[1]), .A2(bbar[6]), .ZN(ybar[22]);
  AND2_X1 U113 ( .A1(a[14]), .A2(b[5]), .ZN(y[229]) );
  OR2_X1 U113bar ( .A1(abar[14]), .A2(bbar[5]), .ZN(ybar[229]);
  AND2_X1 U114 ( .A1(a[14]), .A2(b[4]), .ZN(y[228]) );
  OR2_X1 U114bar ( .A1(abar[14]), .A2(bbar[4]), .ZN(ybar[228]);
  AND2_X1 U115 ( .A1(a[14]), .A2(b[3]), .ZN(y[227]) );
  OR2_X1 U115bar ( .A1(abar[14]), .A2(bbar[3]), .ZN(ybar[227]);
  AND2_X1 U116 ( .A1(a[14]), .A2(b[2]), .ZN(y[226]) );
  OR2_X1 U116bar ( .A1(abar[14]), .A2(bbar[2]), .ZN(ybar[226]);
  AND2_X1 U117 ( .A1(a[14]), .A2(b[1]), .ZN(y[225]) );
  OR2_X1 U117bar ( .A1(abar[14]), .A2(bbar[1]), .ZN(ybar[225]);
  AND2_X1 U118 ( .A1(a[14]), .A2(b[0]), .ZN(y[224]) );
  OR2_X1 U118bar ( .A1(abar[14]), .A2(bbar[0]), .ZN(ybar[224]);
  AND2_X1 U119 ( .A1(a[13]), .A2(b[15]), .ZN(y[223]) );
  OR2_X1 U119bar ( .A1(abar[13]), .A2(bbar[15]), .ZN(ybar[223]);
  AND2_X1 U120 ( .A1(a[13]), .A2(b[14]), .ZN(y[222]) );
  OR2_X1 U120bar ( .A1(abar[13]), .A2(bbar[14]), .ZN(ybar[222]);
  AND2_X1 U121 ( .A1(a[13]), .A2(b[13]), .ZN(y[221]) );
  OR2_X1 U121bar ( .A1(abar[13]), .A2(bbar[13]), .ZN(ybar[221]);
  AND2_X1 U122 ( .A1(a[13]), .A2(b[12]), .ZN(y[220]) );
  OR2_X1 U122bar ( .A1(abar[13]), .A2(bbar[12]), .ZN(ybar[220]);
  AND2_X1 U123 ( .A1(a[1]), .A2(b[5]), .ZN(y[21]) );
  OR2_X1 U123bar ( .A1(abar[1]), .A2(bbar[5]), .ZN(ybar[21]);
  AND2_X1 U124 ( .A1(a[13]), .A2(b[11]), .ZN(y[219]) );
  OR2_X1 U124bar ( .A1(abar[13]), .A2(bbar[11]), .ZN(ybar[219]);
  AND2_X1 U125 ( .A1(a[13]), .A2(b[10]), .ZN(y[218]) );
  OR2_X1 U125bar ( .A1(abar[13]), .A2(bbar[10]), .ZN(ybar[218]);
  AND2_X1 U126 ( .A1(a[13]), .A2(b[9]), .ZN(y[217]) );
  OR2_X1 U126bar ( .A1(abar[13]), .A2(bbar[9]), .ZN(ybar[217]);
  AND2_X1 U127 ( .A1(a[13]), .A2(b[8]), .ZN(y[216]) );
  OR2_X1 U127bar ( .A1(abar[13]), .A2(bbar[8]), .ZN(ybar[216]);
  AND2_X1 U128 ( .A1(a[13]), .A2(b[7]), .ZN(y[215]) );
  OR2_X1 U128bar ( .A1(abar[13]), .A2(bbar[7]), .ZN(ybar[215]);
  AND2_X1 U129 ( .A1(a[13]), .A2(b[6]), .ZN(y[214]) );
  OR2_X1 U129bar ( .A1(abar[13]), .A2(bbar[6]), .ZN(ybar[214]);
  AND2_X1 U130 ( .A1(a[13]), .A2(b[5]), .ZN(y[213]) );
  OR2_X1 U130bar ( .A1(abar[13]), .A2(bbar[5]), .ZN(ybar[213]);
  AND2_X1 U131 ( .A1(a[13]), .A2(b[4]), .ZN(y[212]) );
  OR2_X1 U131bar ( .A1(abar[13]), .A2(bbar[4]), .ZN(ybar[212]);
  AND2_X1 U132 ( .A1(a[13]), .A2(b[3]), .ZN(y[211]) );
  OR2_X1 U132bar ( .A1(abar[13]), .A2(bbar[3]), .ZN(ybar[211]);
  AND2_X1 U133 ( .A1(a[13]), .A2(b[2]), .ZN(y[210]) );
  OR2_X1 U133bar ( .A1(abar[13]), .A2(bbar[2]), .ZN(ybar[210]);
  AND2_X1 U134 ( .A1(a[1]), .A2(b[4]), .ZN(y[20]) );
  OR2_X1 U134bar ( .A1(abar[1]), .A2(bbar[4]), .ZN(ybar[20]);
  AND2_X1 U135 ( .A1(a[13]), .A2(b[1]), .ZN(y[209]) );
  OR2_X1 U135bar ( .A1(abar[13]), .A2(bbar[1]), .ZN(ybar[209]);
  AND2_X1 U136 ( .A1(a[13]), .A2(b[0]), .ZN(y[208]) );
  OR2_X1 U136bar ( .A1(abar[13]), .A2(bbar[0]), .ZN(ybar[208]);
  AND2_X1 U137 ( .A1(a[12]), .A2(b[15]), .ZN(y[207]) );
  OR2_X1 U137bar ( .A1(abar[12]), .A2(bbar[15]), .ZN(ybar[207]);
  AND2_X1 U138 ( .A1(a[12]), .A2(b[14]), .ZN(y[206]) );
  OR2_X1 U138bar ( .A1(abar[12]), .A2(bbar[14]), .ZN(ybar[206]);
  AND2_X1 U139 ( .A1(a[12]), .A2(b[13]), .ZN(y[205]) );
  OR2_X1 U139bar ( .A1(abar[12]), .A2(bbar[13]), .ZN(ybar[205]);
  AND2_X1 U140 ( .A1(a[12]), .A2(b[12]), .ZN(y[204]) );
  OR2_X1 U140bar ( .A1(abar[12]), .A2(bbar[12]), .ZN(ybar[204]);
  AND2_X1 U141 ( .A1(a[12]), .A2(b[11]), .ZN(y[203]) );
  OR2_X1 U141bar ( .A1(abar[12]), .A2(bbar[11]), .ZN(ybar[203]);
  AND2_X1 U142 ( .A1(a[12]), .A2(b[10]), .ZN(y[202]) );
  OR2_X1 U142bar ( .A1(abar[12]), .A2(bbar[10]), .ZN(ybar[202]);
  AND2_X1 U143 ( .A1(a[12]), .A2(b[9]), .ZN(y[201]) );
  OR2_X1 U143bar ( .A1(abar[12]), .A2(bbar[9]), .ZN(ybar[201]);
  AND2_X1 U144 ( .A1(a[12]), .A2(b[8]), .ZN(y[200]) );
  OR2_X1 U144bar ( .A1(abar[12]), .A2(bbar[8]), .ZN(ybar[200]);
  AND2_X1 U145 ( .A1(b[1]), .A2(a[0]), .ZN(y[1]) );
  OR2_X1 U145bar ( .A1(bbar[1]), .A2(abar[0]), .ZN(ybar[1]);
  AND2_X1 U146 ( .A1(a[1]), .A2(b[3]), .ZN(y[19]) );
  OR2_X1 U146bar ( .A1(abar[1]), .A2(bbar[3]), .ZN(ybar[19]);
  AND2_X1 U147 ( .A1(a[12]), .A2(b[7]), .ZN(y[199]) );
  OR2_X1 U147bar ( .A1(abar[12]), .A2(bbar[7]), .ZN(ybar[199]);
  AND2_X1 U148 ( .A1(a[12]), .A2(b[6]), .ZN(y[198]) );
  OR2_X1 U148bar ( .A1(abar[12]), .A2(bbar[6]), .ZN(ybar[198]);
  AND2_X1 U149 ( .A1(a[12]), .A2(b[5]), .ZN(y[197]) );
  OR2_X1 U149bar ( .A1(abar[12]), .A2(bbar[5]), .ZN(ybar[197]);
  AND2_X1 U150 ( .A1(a[12]), .A2(b[4]), .ZN(y[196]) );
  OR2_X1 U150bar ( .A1(abar[12]), .A2(bbar[4]), .ZN(ybar[196]);
  AND2_X1 U151 ( .A1(a[12]), .A2(b[3]), .ZN(y[195]) );
  OR2_X1 U151bar ( .A1(abar[12]), .A2(bbar[3]), .ZN(ybar[195]);
  AND2_X1 U152 ( .A1(a[12]), .A2(b[2]), .ZN(y[194]) );
  OR2_X1 U152bar ( .A1(abar[12]), .A2(bbar[2]), .ZN(ybar[194]);
  AND2_X1 U153 ( .A1(a[12]), .A2(b[1]), .ZN(y[193]) );
  OR2_X1 U153bar ( .A1(abar[12]), .A2(bbar[1]), .ZN(ybar[193]);
  AND2_X1 U154 ( .A1(a[12]), .A2(b[0]), .ZN(y[192]) );
  OR2_X1 U154bar ( .A1(abar[12]), .A2(bbar[0]), .ZN(ybar[192]);
  AND2_X1 U155 ( .A1(a[11]), .A2(b[15]), .ZN(y[191]) );
  OR2_X1 U155bar ( .A1(abar[11]), .A2(bbar[15]), .ZN(ybar[191]);
  AND2_X1 U156 ( .A1(a[11]), .A2(b[14]), .ZN(y[190]) );
  OR2_X1 U156bar ( .A1(abar[11]), .A2(bbar[14]), .ZN(ybar[190]);
  AND2_X1 U157 ( .A1(a[1]), .A2(b[2]), .ZN(y[18]) );
  OR2_X1 U157bar ( .A1(abar[1]), .A2(bbar[2]), .ZN(ybar[18]);
  AND2_X1 U158 ( .A1(a[11]), .A2(b[13]), .ZN(y[189]) );
  OR2_X1 U158bar ( .A1(abar[11]), .A2(bbar[13]), .ZN(ybar[189]);
  AND2_X1 U159 ( .A1(a[11]), .A2(b[12]), .ZN(y[188]) );
  OR2_X1 U159bar ( .A1(abar[11]), .A2(bbar[12]), .ZN(ybar[188]);
  AND2_X1 U160 ( .A1(a[11]), .A2(b[11]), .ZN(y[187]) );
  OR2_X1 U160bar ( .A1(abar[11]), .A2(bbar[11]), .ZN(ybar[187]);
  AND2_X1 U161 ( .A1(a[11]), .A2(b[10]), .ZN(y[186]) );
  OR2_X1 U161bar ( .A1(abar[11]), .A2(bbar[10]), .ZN(ybar[186]);
  AND2_X1 U162 ( .A1(a[11]), .A2(b[9]), .ZN(y[185]) );
  OR2_X1 U162bar ( .A1(abar[11]), .A2(bbar[9]), .ZN(ybar[185]);
  AND2_X1 U163 ( .A1(a[11]), .A2(b[8]), .ZN(y[184]) );
  OR2_X1 U163bar ( .A1(abar[11]), .A2(bbar[8]), .ZN(ybar[184]);
  AND2_X1 U164 ( .A1(a[11]), .A2(b[7]), .ZN(y[183]) );
  OR2_X1 U164bar ( .A1(abar[11]), .A2(bbar[7]), .ZN(ybar[183]);
  AND2_X1 U165 ( .A1(a[11]), .A2(b[6]), .ZN(y[182]) );
  OR2_X1 U165bar ( .A1(abar[11]), .A2(bbar[6]), .ZN(ybar[182]);
  AND2_X1 U166 ( .A1(a[11]), .A2(b[5]), .ZN(y[181]) );
  OR2_X1 U166bar ( .A1(abar[11]), .A2(bbar[5]), .ZN(ybar[181]);
  AND2_X1 U167 ( .A1(a[11]), .A2(b[4]), .ZN(y[180]) );
  OR2_X1 U167bar ( .A1(abar[11]), .A2(bbar[4]), .ZN(ybar[180]);
  AND2_X1 U168 ( .A1(a[1]), .A2(b[1]), .ZN(y[17]) );
  OR2_X1 U168bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[17]);
  AND2_X1 U169 ( .A1(a[11]), .A2(b[3]), .ZN(y[179]) );
  OR2_X1 U169bar ( .A1(abar[11]), .A2(bbar[3]), .ZN(ybar[179]);
  AND2_X1 U170 ( .A1(a[11]), .A2(b[2]), .ZN(y[178]) );
  OR2_X1 U170bar ( .A1(abar[11]), .A2(bbar[2]), .ZN(ybar[178]);
  AND2_X1 U171 ( .A1(a[11]), .A2(b[1]), .ZN(y[177]) );
  OR2_X1 U171bar ( .A1(abar[11]), .A2(bbar[1]), .ZN(ybar[177]);
  AND2_X1 U172 ( .A1(a[11]), .A2(b[0]), .ZN(y[176]) );
  OR2_X1 U172bar ( .A1(abar[11]), .A2(bbar[0]), .ZN(ybar[176]);
  AND2_X1 U173 ( .A1(a[10]), .A2(b[15]), .ZN(y[175]) );
  OR2_X1 U173bar ( .A1(abar[10]), .A2(bbar[15]), .ZN(ybar[175]);
  AND2_X1 U174 ( .A1(a[10]), .A2(b[14]), .ZN(y[174]) );
  OR2_X1 U174bar ( .A1(abar[10]), .A2(bbar[14]), .ZN(ybar[174]);
  AND2_X1 U175 ( .A1(a[10]), .A2(b[13]), .ZN(y[173]) );
  OR2_X1 U175bar ( .A1(abar[10]), .A2(bbar[13]), .ZN(ybar[173]);
  AND2_X1 U176 ( .A1(a[10]), .A2(b[12]), .ZN(y[172]) );
  OR2_X1 U176bar ( .A1(abar[10]), .A2(bbar[12]), .ZN(ybar[172]);
  AND2_X1 U177 ( .A1(a[10]), .A2(b[11]), .ZN(y[171]) );
  OR2_X1 U177bar ( .A1(abar[10]), .A2(bbar[11]), .ZN(ybar[171]);
  AND2_X1 U178 ( .A1(a[10]), .A2(b[10]), .ZN(y[170]) );
  OR2_X1 U178bar ( .A1(abar[10]), .A2(bbar[10]), .ZN(ybar[170]);
  AND2_X1 U179 ( .A1(a[1]), .A2(b[0]), .ZN(y[16]) );
  OR2_X1 U179bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[16]);
  AND2_X1 U180 ( .A1(a[10]), .A2(b[9]), .ZN(y[169]) );
  OR2_X1 U180bar ( .A1(abar[10]), .A2(bbar[9]), .ZN(ybar[169]);
  AND2_X1 U181 ( .A1(a[10]), .A2(b[8]), .ZN(y[168]) );
  OR2_X1 U181bar ( .A1(abar[10]), .A2(bbar[8]), .ZN(ybar[168]);
  AND2_X1 U182 ( .A1(a[10]), .A2(b[7]), .ZN(y[167]) );
  OR2_X1 U182bar ( .A1(abar[10]), .A2(bbar[7]), .ZN(ybar[167]);
  AND2_X1 U183 ( .A1(a[10]), .A2(b[6]), .ZN(y[166]) );
  OR2_X1 U183bar ( .A1(abar[10]), .A2(bbar[6]), .ZN(ybar[166]);
  AND2_X1 U184 ( .A1(a[10]), .A2(b[5]), .ZN(y[165]) );
  OR2_X1 U184bar ( .A1(abar[10]), .A2(bbar[5]), .ZN(ybar[165]);
  AND2_X1 U185 ( .A1(a[10]), .A2(b[4]), .ZN(y[164]) );
  OR2_X1 U185bar ( .A1(abar[10]), .A2(bbar[4]), .ZN(ybar[164]);
  AND2_X1 U186 ( .A1(a[10]), .A2(b[3]), .ZN(y[163]) );
  OR2_X1 U186bar ( .A1(abar[10]), .A2(bbar[3]), .ZN(ybar[163]);
  AND2_X1 U187 ( .A1(a[10]), .A2(b[2]), .ZN(y[162]) );
  OR2_X1 U187bar ( .A1(abar[10]), .A2(bbar[2]), .ZN(ybar[162]);
  AND2_X1 U188 ( .A1(a[10]), .A2(b[1]), .ZN(y[161]) );
  OR2_X1 U188bar ( .A1(abar[10]), .A2(bbar[1]), .ZN(ybar[161]);
  AND2_X1 U189 ( .A1(a[10]), .A2(b[0]), .ZN(y[160]) );
  OR2_X1 U189bar ( .A1(abar[10]), .A2(bbar[0]), .ZN(ybar[160]);
  AND2_X1 U190 ( .A1(b[15]), .A2(a[0]), .ZN(y[15]) );
  OR2_X1 U190bar ( .A1(bbar[15]), .A2(abar[0]), .ZN(ybar[15]);
  AND2_X1 U191 ( .A1(a[9]), .A2(b[15]), .ZN(y[159]) );
  OR2_X1 U191bar ( .A1(abar[9]), .A2(bbar[15]), .ZN(ybar[159]);
  AND2_X1 U192 ( .A1(a[9]), .A2(b[14]), .ZN(y[158]) );
  OR2_X1 U192bar ( .A1(abar[9]), .A2(bbar[14]), .ZN(ybar[158]);
  AND2_X1 U193 ( .A1(a[9]), .A2(b[13]), .ZN(y[157]) );
  OR2_X1 U193bar ( .A1(abar[9]), .A2(bbar[13]), .ZN(ybar[157]);
  AND2_X1 U194 ( .A1(a[9]), .A2(b[12]), .ZN(y[156]) );
  OR2_X1 U194bar ( .A1(abar[9]), .A2(bbar[12]), .ZN(ybar[156]);
  AND2_X1 U195 ( .A1(a[9]), .A2(b[11]), .ZN(y[155]) );
  OR2_X1 U195bar ( .A1(abar[9]), .A2(bbar[11]), .ZN(ybar[155]);
  AND2_X1 U196 ( .A1(a[9]), .A2(b[10]), .ZN(y[154]) );
  OR2_X1 U196bar ( .A1(abar[9]), .A2(bbar[10]), .ZN(ybar[154]);
  AND2_X1 U197 ( .A1(a[9]), .A2(b[9]), .ZN(y[153]) );
  OR2_X1 U197bar ( .A1(abar[9]), .A2(bbar[9]), .ZN(ybar[153]);
  AND2_X1 U198 ( .A1(a[9]), .A2(b[8]), .ZN(y[152]) );
  OR2_X1 U198bar ( .A1(abar[9]), .A2(bbar[8]), .ZN(ybar[152]);
  AND2_X1 U199 ( .A1(a[9]), .A2(b[7]), .ZN(y[151]) );
  OR2_X1 U199bar ( .A1(abar[9]), .A2(bbar[7]), .ZN(ybar[151]);
  AND2_X1 U200 ( .A1(a[9]), .A2(b[6]), .ZN(y[150]) );
  OR2_X1 U200bar ( .A1(abar[9]), .A2(bbar[6]), .ZN(ybar[150]);
  AND2_X1 U201 ( .A1(b[14]), .A2(a[0]), .ZN(y[14]) );
  OR2_X1 U201bar ( .A1(bbar[14]), .A2(abar[0]), .ZN(ybar[14]);
  AND2_X1 U202 ( .A1(a[9]), .A2(b[5]), .ZN(y[149]) );
  OR2_X1 U202bar ( .A1(abar[9]), .A2(bbar[5]), .ZN(ybar[149]);
  AND2_X1 U203 ( .A1(a[9]), .A2(b[4]), .ZN(y[148]) );
  OR2_X1 U203bar ( .A1(abar[9]), .A2(bbar[4]), .ZN(ybar[148]);
  AND2_X1 U204 ( .A1(a[9]), .A2(b[3]), .ZN(y[147]) );
  OR2_X1 U204bar ( .A1(abar[9]), .A2(bbar[3]), .ZN(ybar[147]);
  AND2_X1 U205 ( .A1(a[9]), .A2(b[2]), .ZN(y[146]) );
  OR2_X1 U205bar ( .A1(abar[9]), .A2(bbar[2]), .ZN(ybar[146]);
  AND2_X1 U206 ( .A1(a[9]), .A2(b[1]), .ZN(y[145]) );
  OR2_X1 U206bar ( .A1(abar[9]), .A2(bbar[1]), .ZN(ybar[145]);
  AND2_X1 U207 ( .A1(a[9]), .A2(b[0]), .ZN(y[144]) );
  OR2_X1 U207bar ( .A1(abar[9]), .A2(bbar[0]), .ZN(ybar[144]);
  AND2_X1 U208 ( .A1(a[8]), .A2(b[15]), .ZN(y[143]) );
  OR2_X1 U208bar ( .A1(abar[8]), .A2(bbar[15]), .ZN(ybar[143]);
  AND2_X1 U209 ( .A1(a[8]), .A2(b[14]), .ZN(y[142]) );
  OR2_X1 U209bar ( .A1(abar[8]), .A2(bbar[14]), .ZN(ybar[142]);
  AND2_X1 U210 ( .A1(a[8]), .A2(b[13]), .ZN(y[141]) );
  OR2_X1 U210bar ( .A1(abar[8]), .A2(bbar[13]), .ZN(ybar[141]);
  AND2_X1 U211 ( .A1(a[8]), .A2(b[12]), .ZN(y[140]) );
  OR2_X1 U211bar ( .A1(abar[8]), .A2(bbar[12]), .ZN(ybar[140]);
  AND2_X1 U212 ( .A1(b[13]), .A2(a[0]), .ZN(y[13]) );
  OR2_X1 U212bar ( .A1(bbar[13]), .A2(abar[0]), .ZN(ybar[13]);
  AND2_X1 U213 ( .A1(a[8]), .A2(b[11]), .ZN(y[139]) );
  OR2_X1 U213bar ( .A1(abar[8]), .A2(bbar[11]), .ZN(ybar[139]);
  AND2_X1 U214 ( .A1(a[8]), .A2(b[10]), .ZN(y[138]) );
  OR2_X1 U214bar ( .A1(abar[8]), .A2(bbar[10]), .ZN(ybar[138]);
  AND2_X1 U215 ( .A1(a[8]), .A2(b[9]), .ZN(y[137]) );
  OR2_X1 U215bar ( .A1(abar[8]), .A2(bbar[9]), .ZN(ybar[137]);
  AND2_X1 U216 ( .A1(a[8]), .A2(b[8]), .ZN(y[136]) );
  OR2_X1 U216bar ( .A1(abar[8]), .A2(bbar[8]), .ZN(ybar[136]);
  AND2_X1 U217 ( .A1(a[8]), .A2(b[7]), .ZN(y[135]) );
  OR2_X1 U217bar ( .A1(abar[8]), .A2(bbar[7]), .ZN(ybar[135]);
  AND2_X1 U218 ( .A1(a[8]), .A2(b[6]), .ZN(y[134]) );
  OR2_X1 U218bar ( .A1(abar[8]), .A2(bbar[6]), .ZN(ybar[134]);
  AND2_X1 U219 ( .A1(a[8]), .A2(b[5]), .ZN(y[133]) );
  OR2_X1 U219bar ( .A1(abar[8]), .A2(bbar[5]), .ZN(ybar[133]);
  AND2_X1 U220 ( .A1(a[8]), .A2(b[4]), .ZN(y[132]) );
  OR2_X1 U220bar ( .A1(abar[8]), .A2(bbar[4]), .ZN(ybar[132]);
  AND2_X1 U221 ( .A1(a[8]), .A2(b[3]), .ZN(y[131]) );
  OR2_X1 U221bar ( .A1(abar[8]), .A2(bbar[3]), .ZN(ybar[131]);
  AND2_X1 U222 ( .A1(a[8]), .A2(b[2]), .ZN(y[130]) );
  OR2_X1 U222bar ( .A1(abar[8]), .A2(bbar[2]), .ZN(ybar[130]);
  AND2_X1 U223 ( .A1(b[12]), .A2(a[0]), .ZN(y[12]) );
  OR2_X1 U223bar ( .A1(bbar[12]), .A2(abar[0]), .ZN(ybar[12]);
  AND2_X1 U224 ( .A1(a[8]), .A2(b[1]), .ZN(y[129]) );
  OR2_X1 U224bar ( .A1(abar[8]), .A2(bbar[1]), .ZN(ybar[129]);
  AND2_X1 U225 ( .A1(a[8]), .A2(b[0]), .ZN(y[128]) );
  OR2_X1 U225bar ( .A1(abar[8]), .A2(bbar[0]), .ZN(ybar[128]);
  AND2_X1 U226 ( .A1(a[7]), .A2(b[15]), .ZN(y[127]) );
  OR2_X1 U226bar ( .A1(abar[7]), .A2(bbar[15]), .ZN(ybar[127]);
  AND2_X1 U227 ( .A1(a[7]), .A2(b[14]), .ZN(y[126]) );
  OR2_X1 U227bar ( .A1(abar[7]), .A2(bbar[14]), .ZN(ybar[126]);
  AND2_X1 U228 ( .A1(a[7]), .A2(b[13]), .ZN(y[125]) );
  OR2_X1 U228bar ( .A1(abar[7]), .A2(bbar[13]), .ZN(ybar[125]);
  AND2_X1 U229 ( .A1(a[7]), .A2(b[12]), .ZN(y[124]) );
  OR2_X1 U229bar ( .A1(abar[7]), .A2(bbar[12]), .ZN(ybar[124]);
  AND2_X1 U230 ( .A1(a[7]), .A2(b[11]), .ZN(y[123]) );
  OR2_X1 U230bar ( .A1(abar[7]), .A2(bbar[11]), .ZN(ybar[123]);
  AND2_X1 U231 ( .A1(a[7]), .A2(b[10]), .ZN(y[122]) );
  OR2_X1 U231bar ( .A1(abar[7]), .A2(bbar[10]), .ZN(ybar[122]);
  AND2_X1 U232 ( .A1(a[7]), .A2(b[9]), .ZN(y[121]) );
  OR2_X1 U232bar ( .A1(abar[7]), .A2(bbar[9]), .ZN(ybar[121]);
  AND2_X1 U233 ( .A1(a[7]), .A2(b[8]), .ZN(y[120]) );
  OR2_X1 U233bar ( .A1(abar[7]), .A2(bbar[8]), .ZN(ybar[120]);
  AND2_X1 U234 ( .A1(b[11]), .A2(a[0]), .ZN(y[11]) );
  OR2_X1 U234bar ( .A1(bbar[11]), .A2(abar[0]), .ZN(ybar[11]);
  AND2_X1 U235 ( .A1(a[7]), .A2(b[7]), .ZN(y[119]) );
  OR2_X1 U235bar ( .A1(abar[7]), .A2(bbar[7]), .ZN(ybar[119]);
  AND2_X1 U236 ( .A1(a[7]), .A2(b[6]), .ZN(y[118]) );
  OR2_X1 U236bar ( .A1(abar[7]), .A2(bbar[6]), .ZN(ybar[118]);
  AND2_X1 U237 ( .A1(a[7]), .A2(b[5]), .ZN(y[117]) );
  OR2_X1 U237bar ( .A1(abar[7]), .A2(bbar[5]), .ZN(ybar[117]);
  AND2_X1 U238 ( .A1(a[7]), .A2(b[4]), .ZN(y[116]) );
  OR2_X1 U238bar ( .A1(abar[7]), .A2(bbar[4]), .ZN(ybar[116]);
  AND2_X1 U239 ( .A1(a[7]), .A2(b[3]), .ZN(y[115]) );
  OR2_X1 U239bar ( .A1(abar[7]), .A2(bbar[3]), .ZN(ybar[115]);
  AND2_X1 U240 ( .A1(a[7]), .A2(b[2]), .ZN(y[114]) );
  OR2_X1 U240bar ( .A1(abar[7]), .A2(bbar[2]), .ZN(ybar[114]);
  AND2_X1 U241 ( .A1(a[7]), .A2(b[1]), .ZN(y[113]) );
  OR2_X1 U241bar ( .A1(abar[7]), .A2(bbar[1]), .ZN(ybar[113]);
  AND2_X1 U242 ( .A1(a[7]), .A2(b[0]), .ZN(y[112]) );
  OR2_X1 U242bar ( .A1(abar[7]), .A2(bbar[0]), .ZN(ybar[112]);
  AND2_X1 U243 ( .A1(b[15]), .A2(a[6]), .ZN(y[111]) );
  OR2_X1 U243bar ( .A1(bbar[15]), .A2(abar[6]), .ZN(ybar[111]);
  AND2_X1 U244 ( .A1(b[14]), .A2(a[6]), .ZN(y[110]) );
  OR2_X1 U244bar ( .A1(bbar[14]), .A2(abar[6]), .ZN(ybar[110]);
  AND2_X1 U245 ( .A1(b[10]), .A2(a[0]), .ZN(y[10]) );
  OR2_X1 U245bar ( .A1(bbar[10]), .A2(abar[0]), .ZN(ybar[10]);
  AND2_X1 U246 ( .A1(b[13]), .A2(a[6]), .ZN(y[109]) );
  OR2_X1 U246bar ( .A1(bbar[13]), .A2(abar[6]), .ZN(ybar[109]);
  AND2_X1 U247 ( .A1(b[12]), .A2(a[6]), .ZN(y[108]) );
  OR2_X1 U247bar ( .A1(bbar[12]), .A2(abar[6]), .ZN(ybar[108]);
  AND2_X1 U248 ( .A1(b[11]), .A2(a[6]), .ZN(y[107]) );
  OR2_X1 U248bar ( .A1(bbar[11]), .A2(abar[6]), .ZN(ybar[107]);
  AND2_X1 U249 ( .A1(b[10]), .A2(a[6]), .ZN(y[106]) );
  OR2_X1 U249bar ( .A1(bbar[10]), .A2(abar[6]), .ZN(ybar[106]);
  AND2_X1 U250 ( .A1(a[6]), .A2(b[9]), .ZN(y[105]) );
  OR2_X1 U250bar ( .A1(abar[6]), .A2(bbar[9]), .ZN(ybar[105]);
  AND2_X1 U251 ( .A1(b[8]), .A2(a[6]), .ZN(y[104]) );
  OR2_X1 U251bar ( .A1(bbar[8]), .A2(abar[6]), .ZN(ybar[104]);
  AND2_X1 U252 ( .A1(b[7]), .A2(a[6]), .ZN(y[103]) );
  OR2_X1 U252bar ( .A1(bbar[7]), .A2(abar[6]), .ZN(ybar[103]);
  AND2_X1 U253 ( .A1(b[6]), .A2(a[6]), .ZN(y[102]) );
  OR2_X1 U253bar ( .A1(bbar[6]), .A2(abar[6]), .ZN(ybar[102]);
  AND2_X1 U254 ( .A1(b[5]), .A2(a[6]), .ZN(y[101]) );
  OR2_X1 U254bar ( .A1(bbar[5]), .A2(abar[6]), .ZN(ybar[101]);
  AND2_X1 U255 ( .A1(b[4]), .A2(a[6]), .ZN(y[100]) );
  OR2_X1 U255bar ( .A1(bbar[4]), .A2(abar[6]), .ZN(ybar[100]);
  AND2_X1 U256 ( .A1(b[0]), .A2(a[0]), .ZN(y[0]) );
  OR2_X1 U256bar ( .A1(bbar[0]), .A2(abar[0]), .ZN(ybar[0]);
endmodule




module decode_11 ( in, out );
  input [7:0] in;
  //input_done

  output [255:0] out;
  //output_done

  wire   [15:0] level1;
  wire   [31:0] level2;
  //wire_done

  CD2_44 cd_l1_1 ( .a(in[1]), .b(in[0]), .y(level1[3:0]) );
  CD2_43 cd_l1_2 ( .a(in[3]), .b(in[2]), .y(level1[7:4]) );
  CD2_42 cd_l1_3 ( .a(in[5]), .b(in[4]), .y(level1[11:8]) );
  CD2_41 cd_l1_4 ( .a(in[7]), .b(in[6]), .y(level1[15:12]) );
  CD4_22 cd_l2_1 ( .a(level1[7:4]), .b(level1[3:0]), .y(level2[15:0]) );
  CD4_21 cd_l2_2 ( .a(level1[15:12]), .b(level1[11:8]), .y(level2[31:16]) );
  CD16_11 cd_l3 ( .a(level2[31:16]), .b(level2[15:0]), .y(out) );
endmodule


module encode_11 ( in, out );
  input [255:0] in;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
  assign inbar[8] = ~in[8];
  assign inbar[9] = ~in[9];
  assign inbar[10] = ~in[10];
  assign inbar[11] = ~in[11];
  assign inbar[12] = ~in[12];
  assign inbar[13] = ~in[13];
  assign inbar[14] = ~in[14];
  assign inbar[15] = ~in[15];
  assign inbar[16] = ~in[16];
  assign inbar[17] = ~in[17];
  assign inbar[18] = ~in[18];
  assign inbar[19] = ~in[19];
  assign inbar[20] = ~in[20];
  assign inbar[21] = ~in[21];
  assign inbar[22] = ~in[22];
  assign inbar[23] = ~in[23];
  assign inbar[24] = ~in[24];
  assign inbar[25] = ~in[25];
  assign inbar[26] = ~in[26];
  assign inbar[27] = ~in[27];
  assign inbar[28] = ~in[28];
  assign inbar[29] = ~in[29];
  assign inbar[30] = ~in[30];
  assign inbar[31] = ~in[31];
  assign inbar[32] = ~in[32];
  assign inbar[33] = ~in[33];
  assign inbar[34] = ~in[34];
  assign inbar[35] = ~in[35];
  assign inbar[36] = ~in[36];
  assign inbar[37] = ~in[37];
  assign inbar[38] = ~in[38];
  assign inbar[39] = ~in[39];
  assign inbar[40] = ~in[40];
  assign inbar[41] = ~in[41];
  assign inbar[42] = ~in[42];
  assign inbar[43] = ~in[43];
  assign inbar[44] = ~in[44];
  assign inbar[45] = ~in[45];
  assign inbar[46] = ~in[46];
  assign inbar[47] = ~in[47];
  assign inbar[48] = ~in[48];
  assign inbar[49] = ~in[49];
  assign inbar[50] = ~in[50];
  assign inbar[51] = ~in[51];
  assign inbar[52] = ~in[52];
  assign inbar[53] = ~in[53];
  assign inbar[54] = ~in[54];
  assign inbar[55] = ~in[55];
  assign inbar[56] = ~in[56];
  assign inbar[57] = ~in[57];
  assign inbar[58] = ~in[58];
  assign inbar[59] = ~in[59];
  assign inbar[60] = ~in[60];
  assign inbar[61] = ~in[61];
  assign inbar[62] = ~in[62];
  assign inbar[63] = ~in[63];
  assign inbar[64] = ~in[64];
  assign inbar[65] = ~in[65];
  assign inbar[66] = ~in[66];
  assign inbar[67] = ~in[67];
  assign inbar[68] = ~in[68];
  assign inbar[69] = ~in[69];
  assign inbar[70] = ~in[70];
  assign inbar[71] = ~in[71];
  assign inbar[72] = ~in[72];
  assign inbar[73] = ~in[73];
  assign inbar[74] = ~in[74];
  assign inbar[75] = ~in[75];
  assign inbar[76] = ~in[76];
  assign inbar[77] = ~in[77];
  assign inbar[78] = ~in[78];
  assign inbar[79] = ~in[79];
  assign inbar[80] = ~in[80];
  assign inbar[81] = ~in[81];
  assign inbar[82] = ~in[82];
  assign inbar[83] = ~in[83];
  assign inbar[84] = ~in[84];
  assign inbar[85] = ~in[85];
  assign inbar[86] = ~in[86];
  assign inbar[87] = ~in[87];
  assign inbar[88] = ~in[88];
  assign inbar[89] = ~in[89];
  assign inbar[90] = ~in[90];
  assign inbar[91] = ~in[91];
  assign inbar[92] = ~in[92];
  assign inbar[93] = ~in[93];
  assign inbar[94] = ~in[94];
  assign inbar[95] = ~in[95];
  assign inbar[96] = ~in[96];
  assign inbar[97] = ~in[97];
  assign inbar[98] = ~in[98];
  assign inbar[99] = ~in[99];
  assign inbar[100] = ~in[100];
  assign inbar[101] = ~in[101];
  assign inbar[102] = ~in[102];
  assign inbar[103] = ~in[103];
  assign inbar[104] = ~in[104];
  assign inbar[105] = ~in[105];
  assign inbar[106] = ~in[106];
  assign inbar[107] = ~in[107];
  assign inbar[108] = ~in[108];
  assign inbar[109] = ~in[109];
  assign inbar[110] = ~in[110];
  assign inbar[111] = ~in[111];
  assign inbar[112] = ~in[112];
  assign inbar[113] = ~in[113];
  assign inbar[114] = ~in[114];
  assign inbar[115] = ~in[115];
  assign inbar[116] = ~in[116];
  assign inbar[117] = ~in[117];
  assign inbar[118] = ~in[118];
  assign inbar[119] = ~in[119];
  assign inbar[120] = ~in[120];
  assign inbar[121] = ~in[121];
  assign inbar[122] = ~in[122];
  assign inbar[123] = ~in[123];
  assign inbar[124] = ~in[124];
  assign inbar[125] = ~in[125];
  assign inbar[126] = ~in[126];
  assign inbar[127] = ~in[127];
  assign inbar[128] = ~in[128];
  assign inbar[129] = ~in[129];
  assign inbar[130] = ~in[130];
  assign inbar[131] = ~in[131];
  assign inbar[132] = ~in[132];
  assign inbar[133] = ~in[133];
  assign inbar[134] = ~in[134];
  assign inbar[135] = ~in[135];
  assign inbar[136] = ~in[136];
  assign inbar[137] = ~in[137];
  assign inbar[138] = ~in[138];
  assign inbar[139] = ~in[139];
  assign inbar[140] = ~in[140];
  assign inbar[141] = ~in[141];
  assign inbar[142] = ~in[142];
  assign inbar[143] = ~in[143];
  assign inbar[144] = ~in[144];
  assign inbar[145] = ~in[145];
  assign inbar[146] = ~in[146];
  assign inbar[147] = ~in[147];
  assign inbar[148] = ~in[148];
  assign inbar[149] = ~in[149];
  assign inbar[150] = ~in[150];
  assign inbar[151] = ~in[151];
  assign inbar[152] = ~in[152];
  assign inbar[153] = ~in[153];
  assign inbar[154] = ~in[154];
  assign inbar[155] = ~in[155];
  assign inbar[156] = ~in[156];
  assign inbar[157] = ~in[157];
  assign inbar[158] = ~in[158];
  assign inbar[159] = ~in[159];
  assign inbar[160] = ~in[160];
  assign inbar[161] = ~in[161];
  assign inbar[162] = ~in[162];
  assign inbar[163] = ~in[163];
  assign inbar[164] = ~in[164];
  assign inbar[165] = ~in[165];
  assign inbar[166] = ~in[166];
  assign inbar[167] = ~in[167];
  assign inbar[168] = ~in[168];
  assign inbar[169] = ~in[169];
  assign inbar[170] = ~in[170];
  assign inbar[171] = ~in[171];
  assign inbar[172] = ~in[172];
  assign inbar[173] = ~in[173];
  assign inbar[174] = ~in[174];
  assign inbar[175] = ~in[175];
  assign inbar[176] = ~in[176];
  assign inbar[177] = ~in[177];
  assign inbar[178] = ~in[178];
  assign inbar[179] = ~in[179];
  assign inbar[180] = ~in[180];
  assign inbar[181] = ~in[181];
  assign inbar[182] = ~in[182];
  assign inbar[183] = ~in[183];
  assign inbar[184] = ~in[184];
  assign inbar[185] = ~in[185];
  assign inbar[186] = ~in[186];
  assign inbar[187] = ~in[187];
  assign inbar[188] = ~in[188];
  assign inbar[189] = ~in[189];
  assign inbar[190] = ~in[190];
  assign inbar[191] = ~in[191];
  assign inbar[192] = ~in[192];
  assign inbar[193] = ~in[193];
  assign inbar[194] = ~in[194];
  assign inbar[195] = ~in[195];
  assign inbar[196] = ~in[196];
  assign inbar[197] = ~in[197];
  assign inbar[198] = ~in[198];
  assign inbar[199] = ~in[199];
  assign inbar[200] = ~in[200];
  assign inbar[201] = ~in[201];
  assign inbar[202] = ~in[202];
  assign inbar[203] = ~in[203];
  assign inbar[204] = ~in[204];
  assign inbar[205] = ~in[205];
  assign inbar[206] = ~in[206];
  assign inbar[207] = ~in[207];
  assign inbar[208] = ~in[208];
  assign inbar[209] = ~in[209];
  assign inbar[210] = ~in[210];
  assign inbar[211] = ~in[211];
  assign inbar[212] = ~in[212];
  assign inbar[213] = ~in[213];
  assign inbar[214] = ~in[214];
  assign inbar[215] = ~in[215];
  assign inbar[216] = ~in[216];
  assign inbar[217] = ~in[217];
  assign inbar[218] = ~in[218];
  assign inbar[219] = ~in[219];
  assign inbar[220] = ~in[220];
  assign inbar[221] = ~in[221];
  assign inbar[222] = ~in[222];
  assign inbar[223] = ~in[223];
  assign inbar[224] = ~in[224];
  assign inbar[225] = ~in[225];
  assign inbar[226] = ~in[226];
  assign inbar[227] = ~in[227];
  assign inbar[228] = ~in[228];
  assign inbar[229] = ~in[229];
  assign inbar[230] = ~in[230];
  assign inbar[231] = ~in[231];
  assign inbar[232] = ~in[232];
  assign inbar[233] = ~in[233];
  assign inbar[234] = ~in[234];
  assign inbar[235] = ~in[235];
  assign inbar[236] = ~in[236];
  assign inbar[237] = ~in[237];
  assign inbar[238] = ~in[238];
  assign inbar[239] = ~in[239];
  assign inbar[240] = ~in[240];
  assign inbar[241] = ~in[241];
  assign inbar[242] = ~in[242];
  assign inbar[243] = ~in[243];
  assign inbar[244] = ~in[244];
  assign inbar[245] = ~in[245];
  assign inbar[246] = ~in[246];
  assign inbar[247] = ~in[247];
  assign inbar[248] = ~in[248];
  assign inbar[249] = ~in[249];
  assign inbar[250] = ~in[250];
  assign inbar[251] = ~in[251];
  assign inbar[252] = ~in[252];
  assign inbar[253] = ~in[253];
  assign inbar[254] = ~in[254];
  assign inbar[255] = ~in[255];
  //input_done

  output [7:0] out;
  reg [7:0] outbar;
  //output_done

  wire   in_81, in_80, in_79, in_78, in_77, in_76, in_75, in_74, in_73, in_72,
         in_71, in_70, in_69, in_68, in_67, in_66, in_65, in_64, in_63, in_62,
         in_61, in_60, in_59, in_58, in_57, in_56, in_55, in_54, in_53, in_52,
         in_51, in_50, in_49, in_48, in_47, in_46, in_45, in_44, in_43, in_42,
         in_41, in_40, in_39, in_38, in_37, in_36, in_35, in_34, in_33, in_32,
         in_31, in_30, in_29, in_28, in_27, in_26, in_25, in_24, in_23, in_22,
         in_21, in_20, in_19, in_18, in_17, in_16, in_15, in_14, in_13, in_12,
         in_11, in_10, in_9, in_8, in_7, in_6, in_5, in_4, in_3, in_2, in_1,
         in_0, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972;
  wire in_81bar, in_80bar, in_79bar, in_78bar, in_77bar, in_76bar, in_75bar, in_74bar, in_73bar, in_72bar, in_71bar, in_70bar, in_69bar, in_68bar, in_67bar, in_66bar, in_65bar, in_64bar, in_63bar, in_62bar, in_61bar, in_60bar, in_59bar, in_58bar, in_57bar, in_56bar, in_55bar, in_54bar, in_53bar, in_52bar, in_51bar, in_50bar, in_49bar, in_48bar, in_47bar, in_46bar, in_45bar, in_44bar, in_43bar, in_42bar, in_41bar, in_40bar, in_39bar, in_38bar, in_37bar, in_36bar, in_35bar, in_34bar, in_33bar, in_32bar, in_31bar, in_30bar, in_29bar, in_28bar, in_27bar, in_26bar, in_25bar, in_24bar, in_23bar, in_22bar, in_21bar, in_20bar, in_19bar, in_18bar, in_17bar, in_16bar, in_15bar, in_14bar, in_13bar, in_12bar, in_11bar, in_10bar, in_9bar, in_8bar, in_7bar, in_6bar, in_5bar, in_4bar, in_3bar, in_2bar, in_1bar, in_0bar, n487bar, n488bar, n489bar, n490bar, n491bar, n492bar, n493bar, n494bar, n495bar, n496bar, n497bar, n498bar, n499bar, n500bar, n501bar, n502bar, n503bar, n504bar, n505bar, n506bar, n507bar, n508bar, n509bar, n510bar, n511bar, n512bar, n513bar, n514bar, n515bar, n516bar, n517bar, n518bar, n519bar, n520bar, n521bar, n522bar, n523bar, n524bar, n525bar, n526bar, n527bar, n528bar, n529bar, n530bar, n531bar, n532bar, n533bar, n534bar, n535bar, n536bar, n537bar, n538bar, n539bar, n540bar, n541bar, n542bar, n543bar, n544bar, n545bar, n546bar, n547bar, n548bar, n549bar, n550bar, n551bar, n552bar, n553bar, n554bar, n555bar, n556bar, n557bar, n558bar, n559bar, n560bar, n561bar, n562bar, n563bar, n564bar, n565bar, n566bar, n567bar, n568bar, n569bar, n570bar, n571bar, n572bar, n573bar, n574bar, n575bar, n576bar, n577bar, n578bar, n579bar, n580bar, n581bar, n582bar, n583bar, n584bar, n585bar, n586bar, n587bar, n588bar, n589bar, n590bar, n591bar, n592bar, n593bar, n594bar, n595bar, n596bar, n597bar, n598bar, n599bar, n600bar, n601bar, n602bar, n603bar, n604bar, n605bar, n606bar, n607bar, n608bar, n609bar, n610bar, n611bar, n612bar, n613bar, n614bar, n615bar, n616bar, n617bar, n618bar, n619bar, n620bar, n621bar, n622bar, n623bar, n624bar, n625bar, n626bar, n627bar, n628bar, n629bar, n630bar, n631bar, n632bar, n633bar, n634bar, n635bar, n636bar, n637bar, n638bar, n639bar, n640bar, n641bar, n642bar, n643bar, n644bar, n645bar, n646bar, n647bar, n648bar, n649bar, n650bar, n651bar, n652bar, n653bar, n654bar, n655bar, n656bar, n657bar, n658bar, n659bar, n660bar, n661bar, n662bar, n663bar, n664bar, n665bar, n666bar, n667bar, n668bar, n669bar, n670bar, n671bar, n672bar, n673bar, n674bar, n675bar, n676bar, n677bar, n678bar, n679bar, n680bar, n681bar, n682bar, n683bar, n684bar, n685bar, n686bar, n687bar, n688bar, n689bar, n690bar, n691bar, n692bar, n693bar, n694bar, n695bar, n696bar, n697bar, n698bar, n699bar, n700bar, n701bar, n702bar, n703bar, n704bar, n705bar, n706bar, n707bar, n708bar, n709bar, n710bar, n711bar, n712bar, n713bar, n714bar, n715bar, n716bar, n717bar, n718bar, n719bar, n720bar, n721bar, n722bar, n723bar, n724bar, n725bar, n726bar, n727bar, n728bar, n729bar, n730bar, n731bar, n732bar, n733bar, n734bar, n735bar, n736bar, n737bar, n738bar, n739bar, n740bar, n741bar, n742bar, n743bar, n744bar, n745bar, n746bar, n747bar, n748bar, n749bar, n750bar, n751bar, n752bar, n753bar, n754bar, n755bar, n756bar, n757bar, n758bar, n759bar, n760bar, n761bar, n762bar, n763bar, n764bar, n765bar, n766bar, n767bar, n768bar, n769bar, n770bar, n771bar, n772bar, n773bar, n774bar, n775bar, n776bar, n777bar, n778bar, n779bar, n780bar, n781bar, n782bar, n783bar, n784bar, n785bar, n786bar, n787bar, n788bar, n789bar, n790bar, n791bar, n792bar, n793bar, n794bar, n795bar, n796bar, n797bar, n798bar, n799bar, n800bar, n801bar, n802bar, n803bar, n804bar, n805bar, n806bar, n807bar, n808bar, n809bar, n810bar, n811bar, n812bar, n813bar, n814bar, n815bar, n816bar, n817bar, n818bar, n819bar, n820bar, n821bar, n822bar, n823bar, n824bar, n825bar, n826bar, n827bar, n828bar, n829bar, n830bar, n831bar, n832bar, n833bar, n834bar, n835bar, n836bar, n837bar, n838bar, n839bar, n840bar, n841bar, n842bar, n843bar, n844bar, n845bar, n846bar, n847bar, n848bar, n849bar, n850bar, n851bar, n852bar, n853bar, n854bar, n855bar, n856bar, n857bar, n858bar, n859bar, n860bar, n861bar, n862bar, n863bar, n864bar, n865bar, n866bar, n867bar, n868bar, n869bar, n870bar, n871bar, n872bar, n873bar, n874bar, n875bar, n876bar, n877bar, n878bar, n879bar, n880bar, n881bar, n882bar, n883bar, n884bar, n885bar, n886bar, n887bar, n888bar, n889bar, n890bar, n891bar, n892bar, n893bar, n894bar, n895bar, n896bar, n897bar, n898bar, n899bar, n900bar, n901bar, n902bar, n903bar, n904bar, n905bar, n906bar, n907bar, n908bar, n909bar, n910bar, n911bar, n912bar, n913bar, n914bar, n915bar, n916bar, n917bar, n918bar, n919bar, n920bar, n921bar, n922bar, n923bar, n924bar, n925bar, n926bar, n927bar, n928bar, n929bar, n930bar, n931bar, n932bar, n933bar, n934bar, n935bar, n936bar, n937bar, n938bar, n939bar, n940bar, n941bar, n942bar, n943bar, n944bar, n945bar, n946bar, n947bar, n948bar, n949bar, n950bar, n951bar, n952bar, n953bar, n954bar, n955bar, n956bar, n957bar, n958bar, n959bar, n960bar, n961bar, n962bar, n963bar, n964bar, n965bar, n966bar, n967bar, n968bar, n969bar, n970bar, n971bar, n972bar;
  //wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];

  OR2_X1 U1 ( .A1(n972), .A2(n971), .ZN(out[7]) );
  AND2_X1 U1bar ( .A1(n972bar), .A2(n971bar), .ZN(outbar[7]);
  OR2_X1 U2 ( .A1(n970), .A2(n969), .ZN(n971) );
  AND2_X1 U2bar ( .A1(n970bar), .A2(n969bar), .ZN(n971bar);
  OR2_X1 U3 ( .A1(n968), .A2(n967), .ZN(n969) );
  AND2_X1 U3bar ( .A1(n968bar), .A2(n967bar), .ZN(n969bar);
  OR2_X1 U4 ( .A1(n966), .A2(n965), .ZN(n967) );
  AND2_X1 U4bar ( .A1(n966bar), .A2(n965bar), .ZN(n967bar);
  OR2_X1 U5 ( .A1(n964), .A2(n963), .ZN(n968) );
  AND2_X1 U5bar ( .A1(n964bar), .A2(n963bar), .ZN(n968bar);
  OR2_X1 U6 ( .A1(in[116]), .A2(n962), .ZN(n963) );
  AND2_X1 U6bar ( .A1(inbar[116]), .A2(n962bar), .ZN(n963bar);
  OR2_X1 U7 ( .A1(n961), .A2(n960), .ZN(n970) );
  AND2_X1 U7bar ( .A1(n961bar), .A2(n960bar), .ZN(n970bar);
  OR2_X1 U8 ( .A1(in[150]), .A2(in[127]), .ZN(n960) );
  AND2_X1 U8bar ( .A1(inbar[150]), .A2(inbar[127]), .ZN(n960bar);
  OR2_X1 U9 ( .A1(in[160]), .A2(n959), .ZN(n961) );
  AND2_X1 U9bar ( .A1(inbar[160]), .A2(n959bar), .ZN(n961bar);
  OR2_X1 U10 ( .A1(in[252]), .A2(in[168]), .ZN(n959) );
  AND2_X1 U10bar ( .A1(inbar[252]), .A2(inbar[168]), .ZN(n959bar);
  OR2_X1 U11 ( .A1(n958), .A2(n957), .ZN(n972) );
  AND2_X1 U11bar ( .A1(n958bar), .A2(n957bar), .ZN(n972bar);
  OR2_X1 U12 ( .A1(n956), .A2(n955), .ZN(n957) );
  AND2_X1 U12bar ( .A1(n956bar), .A2(n955bar), .ZN(n957bar);
  OR2_X1 U13 ( .A1(in_17), .A2(in[96]), .ZN(n955) );
  AND2_X1 U13bar ( .A1(in_17bar), .A2(inbar[96]), .ZN(n955bar);
  OR2_X1 U14 ( .A1(in_23), .A2(n954), .ZN(n956) );
  AND2_X1 U14bar ( .A1(in_23bar), .A2(n954bar), .ZN(n956bar);
  OR2_X1 U15 ( .A1(in_31), .A2(in_26), .ZN(n954) );
  AND2_X1 U15bar ( .A1(in_31bar), .A2(in_26bar), .ZN(n954bar);
  OR2_X1 U16 ( .A1(n953), .A2(n952), .ZN(n958) );
  AND2_X1 U16bar ( .A1(n953bar), .A2(n952bar), .ZN(n958bar);
  OR2_X1 U17 ( .A1(in_58), .A2(in_4), .ZN(n952) );
  AND2_X1 U17bar ( .A1(in_58bar), .A2(in_4bar), .ZN(n952bar);
  OR2_X1 U18 ( .A1(in_59), .A2(n951), .ZN(n953) );
  AND2_X1 U18bar ( .A1(in_59bar), .A2(n951bar), .ZN(n953bar);
  OR2_X1 U19 ( .A1(in_71), .A2(in_62), .ZN(n951) );
  AND2_X1 U19bar ( .A1(in_71bar), .A2(in_62bar), .ZN(n951bar);
  OR2_X1 U20 ( .A1(n950), .A2(n949), .ZN(out[6]) );
  AND2_X1 U20bar ( .A1(n950bar), .A2(n949bar), .ZN(outbar[6]);
  OR2_X1 U21 ( .A1(n948), .A2(n947), .ZN(n949) );
  AND2_X1 U21bar ( .A1(n948bar), .A2(n947bar), .ZN(n949bar);
  OR2_X1 U22 ( .A1(n946), .A2(n945), .ZN(n947) );
  AND2_X1 U22bar ( .A1(n946bar), .A2(n945bar), .ZN(n947bar);
  OR2_X1 U23 ( .A1(n944), .A2(n943), .ZN(n945) );
  AND2_X1 U23bar ( .A1(n944bar), .A2(n943bar), .ZN(n945bar);
  OR2_X1 U24 ( .A1(n942), .A2(n941), .ZN(n946) );
  AND2_X1 U24bar ( .A1(n942bar), .A2(n941bar), .ZN(n946bar);
  OR2_X1 U25 ( .A1(in[101]), .A2(n940), .ZN(n941) );
  AND2_X1 U25bar ( .A1(inbar[101]), .A2(n940bar), .ZN(n941bar);
  OR2_X1 U26 ( .A1(n939), .A2(n938), .ZN(n948) );
  AND2_X1 U26bar ( .A1(n939bar), .A2(n938bar), .ZN(n948bar);
  OR2_X1 U27 ( .A1(in[114]), .A2(in[104]), .ZN(n938) );
  AND2_X1 U27bar ( .A1(inbar[114]), .A2(inbar[104]), .ZN(n938bar);
  OR2_X1 U28 ( .A1(in[128]), .A2(n937), .ZN(n939) );
  AND2_X1 U28bar ( .A1(inbar[128]), .A2(n937bar), .ZN(n939bar);
  OR2_X1 U29 ( .A1(in[136]), .A2(in[134]), .ZN(n937) );
  AND2_X1 U29bar ( .A1(inbar[136]), .A2(inbar[134]), .ZN(n937bar);
  OR2_X1 U30 ( .A1(n936), .A2(n935), .ZN(n950) );
  AND2_X1 U30bar ( .A1(n936bar), .A2(n935bar), .ZN(n950bar);
  OR2_X1 U31 ( .A1(n934), .A2(n933), .ZN(n935) );
  AND2_X1 U31bar ( .A1(n934bar), .A2(n933bar), .ZN(n935bar);
  OR2_X1 U32 ( .A1(in[177]), .A2(in[164]), .ZN(n933) );
  AND2_X1 U32bar ( .A1(inbar[177]), .A2(inbar[164]), .ZN(n933bar);
  OR2_X1 U33 ( .A1(in[212]), .A2(n932), .ZN(n934) );
  AND2_X1 U33bar ( .A1(inbar[212]), .A2(n932bar), .ZN(n934bar);
  OR2_X1 U34 ( .A1(in[248]), .A2(in[221]), .ZN(n932) );
  AND2_X1 U34bar ( .A1(inbar[248]), .A2(inbar[221]), .ZN(n932bar);
  OR2_X1 U35 ( .A1(n931), .A2(n930), .ZN(n936) );
  AND2_X1 U35bar ( .A1(n931bar), .A2(n930bar), .ZN(n936bar);
  OR2_X1 U36 ( .A1(in_18), .A2(in[93]), .ZN(n930) );
  AND2_X1 U36bar ( .A1(in_18bar), .A2(inbar[93]), .ZN(n930bar);
  OR2_X1 U37 ( .A1(in_31), .A2(n929), .ZN(n931) );
  AND2_X1 U37bar ( .A1(in_31bar), .A2(n929bar), .ZN(n931bar);
  OR2_X1 U38 ( .A1(in_7), .A2(in_39), .ZN(n929) );
  AND2_X1 U38bar ( .A1(in_7bar), .A2(in_39bar), .ZN(n929bar);
  OR2_X1 U39 ( .A1(n928), .A2(n927), .ZN(out[5]) );
  AND2_X1 U39bar ( .A1(n928bar), .A2(n927bar), .ZN(outbar[5]);
  OR2_X1 U40 ( .A1(n926), .A2(n925), .ZN(n927) );
  AND2_X1 U40bar ( .A1(n926bar), .A2(n925bar), .ZN(n927bar);
  OR2_X1 U41 ( .A1(n924), .A2(n923), .ZN(n925) );
  AND2_X1 U41bar ( .A1(n924bar), .A2(n923bar), .ZN(n925bar);
  OR2_X1 U42 ( .A1(n922), .A2(n921), .ZN(n923) );
  AND2_X1 U42bar ( .A1(n922bar), .A2(n921bar), .ZN(n923bar);
  OR2_X1 U43 ( .A1(n940), .A2(n920), .ZN(n924) );
  AND2_X1 U43bar ( .A1(n940bar), .A2(n920bar), .ZN(n924bar);
  OR2_X1 U44 ( .A1(in[111]), .A2(n919), .ZN(n920) );
  AND2_X1 U44bar ( .A1(inbar[111]), .A2(n919bar), .ZN(n920bar);
  OR2_X1 U45 ( .A1(n918), .A2(n917), .ZN(n940) );
  AND2_X1 U45bar ( .A1(n918bar), .A2(n917bar), .ZN(n940bar);
  OR2_X1 U46 ( .A1(n916), .A2(n915), .ZN(n917) );
  AND2_X1 U46bar ( .A1(n916bar), .A2(n915bar), .ZN(n917bar);
  OR2_X1 U47 ( .A1(n914), .A2(n913), .ZN(n915) );
  AND2_X1 U47bar ( .A1(n914bar), .A2(n913bar), .ZN(n915bar);
  OR2_X1 U48 ( .A1(in[140]), .A2(in[131]), .ZN(n913) );
  AND2_X1 U48bar ( .A1(inbar[140]), .A2(inbar[131]), .ZN(n913bar);
  OR2_X1 U49 ( .A1(in[160]), .A2(in[144]), .ZN(n914) );
  AND2_X1 U49bar ( .A1(inbar[160]), .A2(inbar[144]), .ZN(n914bar);
  OR2_X1 U50 ( .A1(n912), .A2(n911), .ZN(n916) );
  AND2_X1 U50bar ( .A1(n912bar), .A2(n911bar), .ZN(n916bar);
  OR2_X1 U51 ( .A1(in[179]), .A2(in[174]), .ZN(n911) );
  AND2_X1 U51bar ( .A1(inbar[179]), .A2(inbar[174]), .ZN(n911bar);
  OR2_X1 U52 ( .A1(in[188]), .A2(in[184]), .ZN(n912) );
  AND2_X1 U52bar ( .A1(inbar[188]), .A2(inbar[184]), .ZN(n912bar);
  OR2_X1 U53 ( .A1(n910), .A2(n909), .ZN(n918) );
  AND2_X1 U53bar ( .A1(n910bar), .A2(n909bar), .ZN(n918bar);
  OR2_X1 U54 ( .A1(n908), .A2(n907), .ZN(n909) );
  AND2_X1 U54bar ( .A1(n908bar), .A2(n907bar), .ZN(n909bar);
  OR2_X1 U55 ( .A1(in[216]), .A2(in[200]), .ZN(n907) );
  AND2_X1 U55bar ( .A1(inbar[216]), .A2(inbar[200]), .ZN(n907bar);
  OR2_X1 U56 ( .A1(in[228]), .A2(in[224]), .ZN(n908) );
  AND2_X1 U56bar ( .A1(inbar[228]), .A2(inbar[224]), .ZN(n908bar);
  OR2_X1 U57 ( .A1(n906), .A2(n905), .ZN(n910) );
  AND2_X1 U57bar ( .A1(n906bar), .A2(n905bar), .ZN(n910bar);
  OR2_X1 U58 ( .A1(in[247]), .A2(in[235]), .ZN(n905) );
  AND2_X1 U58bar ( .A1(inbar[247]), .A2(inbar[235]), .ZN(n905bar);
  OR2_X1 U59 ( .A1(in_42), .A2(in[83]), .ZN(n906) );
  AND2_X1 U59bar ( .A1(in_42bar), .A2(inbar[83]), .ZN(n906bar);
  OR2_X1 U60 ( .A1(n904), .A2(n903), .ZN(n926) );
  AND2_X1 U60bar ( .A1(n904bar), .A2(n903bar), .ZN(n926bar);
  OR2_X1 U61 ( .A1(in[166]), .A2(in[123]), .ZN(n903) );
  AND2_X1 U61bar ( .A1(inbar[166]), .A2(inbar[123]), .ZN(n903bar);
  OR2_X1 U62 ( .A1(in[170]), .A2(n902), .ZN(n904) );
  AND2_X1 U62bar ( .A1(inbar[170]), .A2(n902bar), .ZN(n904bar);
  OR2_X1 U63 ( .A1(in[194]), .A2(in[183]), .ZN(n902) );
  AND2_X1 U63bar ( .A1(inbar[194]), .A2(inbar[183]), .ZN(n902bar);
  OR2_X1 U64 ( .A1(n901), .A2(n900), .ZN(n928) );
  AND2_X1 U64bar ( .A1(n901bar), .A2(n900bar), .ZN(n928bar);
  OR2_X1 U65 ( .A1(n899), .A2(n898), .ZN(n900) );
  AND2_X1 U65bar ( .A1(n899bar), .A2(n898bar), .ZN(n900bar);
  OR2_X1 U66 ( .A1(in[241]), .A2(in[238]), .ZN(n898) );
  AND2_X1 U66bar ( .A1(inbar[241]), .A2(inbar[238]), .ZN(n898bar);
  OR2_X1 U67 ( .A1(in[250]), .A2(n897), .ZN(n899) );
  AND2_X1 U67bar ( .A1(inbar[250]), .A2(n897bar), .ZN(n899bar);
  OR2_X1 U68 ( .A1(in_24), .A2(in[84]), .ZN(n897) );
  AND2_X1 U68bar ( .A1(in_24bar), .A2(inbar[84]), .ZN(n897bar);
  OR2_X1 U69 ( .A1(n896), .A2(n895), .ZN(n901) );
  AND2_X1 U69bar ( .A1(n896bar), .A2(n895bar), .ZN(n901bar);
  OR2_X1 U70 ( .A1(in_41), .A2(in_29), .ZN(n895) );
  AND2_X1 U70bar ( .A1(in_41bar), .A2(in_29bar), .ZN(n895bar);
  OR2_X1 U71 ( .A1(in_66), .A2(n894), .ZN(n896) );
  AND2_X1 U71bar ( .A1(in_66bar), .A2(n894bar), .ZN(n896bar);
  OR2_X1 U72 ( .A1(in_76), .A2(in_71), .ZN(n894) );
  AND2_X1 U72bar ( .A1(in_76bar), .A2(in_71bar), .ZN(n894bar);
  OR2_X1 U73 ( .A1(n893), .A2(n892), .ZN(out[4]) );
  AND2_X1 U73bar ( .A1(n893bar), .A2(n892bar), .ZN(outbar[4]);
  OR2_X1 U74 ( .A1(n891), .A2(n890), .ZN(n892) );
  AND2_X1 U74bar ( .A1(n891bar), .A2(n890bar), .ZN(n892bar);
  OR2_X1 U75 ( .A1(n889), .A2(n888), .ZN(n890) );
  AND2_X1 U75bar ( .A1(n889bar), .A2(n888bar), .ZN(n890bar);
  OR2_X1 U76 ( .A1(n922), .A2(n887), .ZN(n888) );
  AND2_X1 U76bar ( .A1(n922bar), .A2(n887bar), .ZN(n888bar);
  OR2_X1 U77 ( .A1(n886), .A2(n885), .ZN(n922) );
  AND2_X1 U77bar ( .A1(n886bar), .A2(n885bar), .ZN(n922bar);
  OR2_X1 U78 ( .A1(n884), .A2(n883), .ZN(n885) );
  AND2_X1 U78bar ( .A1(n884bar), .A2(n883bar), .ZN(n885bar);
  OR2_X1 U79 ( .A1(n882), .A2(n881), .ZN(n883) );
  AND2_X1 U79bar ( .A1(n882bar), .A2(n881bar), .ZN(n883bar);
  OR2_X1 U80 ( .A1(in[118]), .A2(in[109]), .ZN(n881) );
  AND2_X1 U80bar ( .A1(inbar[118]), .A2(inbar[109]), .ZN(n881bar);
  OR2_X1 U81 ( .A1(in[139]), .A2(in[120]), .ZN(n882) );
  AND2_X1 U81bar ( .A1(inbar[139]), .A2(inbar[120]), .ZN(n882bar);
  OR2_X1 U82 ( .A1(n880), .A2(n879), .ZN(n884) );
  AND2_X1 U82bar ( .A1(n880bar), .A2(n879bar), .ZN(n884bar);
  OR2_X1 U83 ( .A1(in[198]), .A2(in[154]), .ZN(n879) );
  AND2_X1 U83bar ( .A1(inbar[198]), .A2(inbar[154]), .ZN(n879bar);
  OR2_X1 U84 ( .A1(in[210]), .A2(in[205]), .ZN(n880) );
  AND2_X1 U84bar ( .A1(inbar[210]), .A2(inbar[205]), .ZN(n880bar);
  OR2_X1 U85 ( .A1(n878), .A2(n877), .ZN(n886) );
  AND2_X1 U85bar ( .A1(n878bar), .A2(n877bar), .ZN(n886bar);
  OR2_X1 U86 ( .A1(n876), .A2(n875), .ZN(n877) );
  AND2_X1 U86bar ( .A1(n876bar), .A2(n875bar), .ZN(n877bar);
  OR2_X1 U87 ( .A1(in[219]), .A2(in[217]), .ZN(n875) );
  AND2_X1 U87bar ( .A1(inbar[219]), .A2(inbar[217]), .ZN(n875bar);
  OR2_X1 U88 ( .A1(in[86]), .A2(in[252]), .ZN(n876) );
  AND2_X1 U88bar ( .A1(inbar[86]), .A2(inbar[252]), .ZN(n876bar);
  OR2_X1 U89 ( .A1(n874), .A2(n873), .ZN(n878) );
  AND2_X1 U89bar ( .A1(n874bar), .A2(n873bar), .ZN(n878bar);
  OR2_X1 U90 ( .A1(in_40), .A2(in[91]), .ZN(n873) );
  AND2_X1 U90bar ( .A1(in_40bar), .A2(inbar[91]), .ZN(n873bar);
  OR2_X1 U91 ( .A1(in_8), .A2(in_46), .ZN(n874) );
  AND2_X1 U91bar ( .A1(in_8bar), .A2(in_46bar), .ZN(n874bar);
  OR2_X1 U92 ( .A1(n872), .A2(n871), .ZN(n889) );
  AND2_X1 U92bar ( .A1(n872bar), .A2(n871bar), .ZN(n889bar);
  OR2_X1 U93 ( .A1(in[117]), .A2(n943), .ZN(n871) );
  AND2_X1 U93bar ( .A1(inbar[117]), .A2(n943bar), .ZN(n871bar);
  OR2_X1 U94 ( .A1(n870), .A2(n869), .ZN(n943) );
  AND2_X1 U94bar ( .A1(n870bar), .A2(n869bar), .ZN(n943bar);
  OR2_X1 U95 ( .A1(n868), .A2(n867), .ZN(n869) );
  AND2_X1 U95bar ( .A1(n868bar), .A2(n867bar), .ZN(n869bar);
  OR2_X1 U96 ( .A1(n866), .A2(n865), .ZN(n867) );
  AND2_X1 U96bar ( .A1(n866bar), .A2(n865bar), .ZN(n867bar);
  OR2_X1 U97 ( .A1(n864), .A2(n863), .ZN(n865) );
  AND2_X1 U97bar ( .A1(n864bar), .A2(n863bar), .ZN(n865bar);
  OR2_X1 U98 ( .A1(in[108]), .A2(n919), .ZN(n866) );
  AND2_X1 U98bar ( .A1(inbar[108]), .A2(n919bar), .ZN(n866bar);
  OR2_X1 U99 ( .A1(n862), .A2(n861), .ZN(n919) );
  AND2_X1 U99bar ( .A1(n862bar), .A2(n861bar), .ZN(n919bar);
  OR2_X1 U100 ( .A1(n860), .A2(n859), .ZN(n861) );
  AND2_X1 U100bar ( .A1(n860bar), .A2(n859bar), .ZN(n861bar);
  OR2_X1 U101 ( .A1(n858), .A2(n857), .ZN(n859) );
  AND2_X1 U101bar ( .A1(n858bar), .A2(n857bar), .ZN(n859bar);
  OR2_X1 U102 ( .A1(in[119]), .A2(in[105]), .ZN(n857) );
  AND2_X1 U102bar ( .A1(inbar[119]), .A2(inbar[105]), .ZN(n857bar);
  OR2_X1 U103 ( .A1(in[186]), .A2(in[175]), .ZN(n858) );
  AND2_X1 U103bar ( .A1(inbar[186]), .A2(inbar[175]), .ZN(n858bar);
  OR2_X1 U104 ( .A1(n856), .A2(n855), .ZN(n860) );
  AND2_X1 U104bar ( .A1(n856bar), .A2(n855bar), .ZN(n860bar);
  OR2_X1 U105 ( .A1(in[202]), .A2(in[193]), .ZN(n855) );
  AND2_X1 U105bar ( .A1(inbar[202]), .A2(inbar[193]), .ZN(n855bar);
  OR2_X1 U106 ( .A1(in[225]), .A2(in[208]), .ZN(n856) );
  AND2_X1 U106bar ( .A1(inbar[225]), .A2(inbar[208]), .ZN(n856bar);
  OR2_X1 U107 ( .A1(n854), .A2(n853), .ZN(n862) );
  AND2_X1 U107bar ( .A1(n854bar), .A2(n853bar), .ZN(n862bar);
  OR2_X1 U108 ( .A1(n852), .A2(n851), .ZN(n853) );
  AND2_X1 U108bar ( .A1(n852bar), .A2(n851bar), .ZN(n853bar);
  OR2_X1 U109 ( .A1(in_1), .A2(in[85]), .ZN(n851) );
  AND2_X1 U109bar ( .A1(in_1bar), .A2(inbar[85]), .ZN(n851bar);
  OR2_X1 U110 ( .A1(in_23), .A2(in_19), .ZN(n852) );
  AND2_X1 U110bar ( .A1(in_23bar), .A2(in_19bar), .ZN(n852bar);
  OR2_X1 U111 ( .A1(n850), .A2(n849), .ZN(n854) );
  AND2_X1 U111bar ( .A1(n850bar), .A2(n849bar), .ZN(n854bar);
  OR2_X1 U112 ( .A1(in_43), .A2(in_33), .ZN(n849) );
  AND2_X1 U112bar ( .A1(in_43bar), .A2(in_33bar), .ZN(n849bar);
  OR2_X1 U113 ( .A1(in_63), .A2(in_44), .ZN(n850) );
  AND2_X1 U113bar ( .A1(in_63bar), .A2(in_44bar), .ZN(n850bar);
  OR2_X1 U114 ( .A1(n848), .A2(n847), .ZN(n868) );
  AND2_X1 U114bar ( .A1(n848bar), .A2(n847bar), .ZN(n868bar);
  OR2_X1 U115 ( .A1(in[141]), .A2(in[112]), .ZN(n847) );
  AND2_X1 U115bar ( .A1(inbar[141]), .A2(inbar[112]), .ZN(n847bar);
  OR2_X1 U116 ( .A1(in[147]), .A2(n846), .ZN(n848) );
  AND2_X1 U116bar ( .A1(inbar[147]), .A2(n846bar), .ZN(n848bar);
  OR2_X1 U117 ( .A1(in[181]), .A2(in[167]), .ZN(n846) );
  AND2_X1 U117bar ( .A1(inbar[181]), .A2(inbar[167]), .ZN(n846bar);
  OR2_X1 U118 ( .A1(n845), .A2(n844), .ZN(n870) );
  AND2_X1 U118bar ( .A1(n845bar), .A2(n844bar), .ZN(n870bar);
  OR2_X1 U119 ( .A1(n843), .A2(n842), .ZN(n844) );
  AND2_X1 U119bar ( .A1(n843bar), .A2(n842bar), .ZN(n844bar);
  OR2_X1 U120 ( .A1(in[229]), .A2(in[201]), .ZN(n842) );
  AND2_X1 U120bar ( .A1(inbar[229]), .A2(inbar[201]), .ZN(n842bar);
  OR2_X1 U121 ( .A1(in[237]), .A2(n841), .ZN(n843) );
  AND2_X1 U121bar ( .A1(inbar[237]), .A2(n841bar), .ZN(n843bar);
  OR2_X1 U122 ( .A1(in[94]), .A2(in[253]), .ZN(n841) );
  AND2_X1 U122bar ( .A1(inbar[94]), .A2(inbar[253]), .ZN(n841bar);
  OR2_X1 U123 ( .A1(n840), .A2(n839), .ZN(n845) );
  AND2_X1 U123bar ( .A1(n840bar), .A2(n839bar), .ZN(n845bar);
  OR2_X1 U124 ( .A1(in_21), .A2(in[96]), .ZN(n839) );
  AND2_X1 U124bar ( .A1(in_21bar), .A2(inbar[96]), .ZN(n839bar);
  OR2_X1 U125 ( .A1(in_25), .A2(n838), .ZN(n840) );
  AND2_X1 U125bar ( .A1(in_25bar), .A2(n838bar), .ZN(n840bar);
  OR2_X1 U126 ( .A1(in_81), .A2(in_45), .ZN(n838) );
  AND2_X1 U126bar ( .A1(in_81bar), .A2(in_45bar), .ZN(n838bar);
  OR2_X1 U127 ( .A1(n837), .A2(n836), .ZN(n891) );
  AND2_X1 U127bar ( .A1(n837bar), .A2(n836bar), .ZN(n891bar);
  OR2_X1 U128 ( .A1(in[142]), .A2(in[124]), .ZN(n836) );
  AND2_X1 U128bar ( .A1(inbar[142]), .A2(inbar[124]), .ZN(n836bar);
  OR2_X1 U129 ( .A1(in[150]), .A2(n835), .ZN(n837) );
  AND2_X1 U129bar ( .A1(inbar[150]), .A2(n835bar), .ZN(n837bar);
  OR2_X1 U130 ( .A1(in[172]), .A2(in[155]), .ZN(n835) );
  AND2_X1 U130bar ( .A1(inbar[172]), .A2(inbar[155]), .ZN(n835bar);
  OR2_X1 U131 ( .A1(n834), .A2(n833), .ZN(n893) );
  AND2_X1 U131bar ( .A1(n834bar), .A2(n833bar), .ZN(n893bar);
  OR2_X1 U132 ( .A1(n832), .A2(n831), .ZN(n833) );
  AND2_X1 U132bar ( .A1(n832bar), .A2(n831bar), .ZN(n833bar);
  OR2_X1 U133 ( .A1(in[196]), .A2(in[173]), .ZN(n831) );
  AND2_X1 U133bar ( .A1(inbar[196]), .A2(inbar[173]), .ZN(n831bar);
  OR2_X1 U134 ( .A1(in[222]), .A2(n830), .ZN(n832) );
  AND2_X1 U134bar ( .A1(inbar[222]), .A2(n830bar), .ZN(n832bar);
  OR2_X1 U135 ( .A1(in[227]), .A2(in[226]), .ZN(n830) );
  AND2_X1 U135bar ( .A1(inbar[227]), .A2(inbar[226]), .ZN(n830bar);
  OR2_X1 U136 ( .A1(n829), .A2(n828), .ZN(n834) );
  AND2_X1 U136bar ( .A1(n829bar), .A2(n828bar), .ZN(n834bar);
  OR2_X1 U137 ( .A1(in[249]), .A2(in[231]), .ZN(n828) );
  AND2_X1 U137bar ( .A1(inbar[249]), .A2(inbar[231]), .ZN(n828bar);
  OR2_X1 U138 ( .A1(in_28), .A2(n827), .ZN(n829) );
  AND2_X1 U138bar ( .A1(in_28bar), .A2(n827bar), .ZN(n829bar);
  OR2_X1 U139 ( .A1(in_52), .A2(in_47), .ZN(n827) );
  AND2_X1 U139bar ( .A1(in_52bar), .A2(in_47bar), .ZN(n827bar);
  OR2_X1 U140 ( .A1(n826), .A2(n825), .ZN(out[3]) );
  AND2_X1 U140bar ( .A1(n826bar), .A2(n825bar), .ZN(outbar[3]);
  OR2_X1 U141 ( .A1(n824), .A2(n823), .ZN(n825) );
  AND2_X1 U141bar ( .A1(n824bar), .A2(n823bar), .ZN(n825bar);
  OR2_X1 U142 ( .A1(n822), .A2(n821), .ZN(n823) );
  AND2_X1 U142bar ( .A1(n822bar), .A2(n821bar), .ZN(n823bar);
  OR2_X1 U143 ( .A1(n820), .A2(n819), .ZN(n821) );
  AND2_X1 U143bar ( .A1(n820bar), .A2(n819bar), .ZN(n821bar);
  OR2_X1 U144 ( .A1(n964), .A2(n818), .ZN(n822) );
  AND2_X1 U144bar ( .A1(n964bar), .A2(n818bar), .ZN(n822bar);
  OR2_X1 U145 ( .A1(in[118]), .A2(n817), .ZN(n818) );
  AND2_X1 U145bar ( .A1(inbar[118]), .A2(n817bar), .ZN(n818bar);
  OR2_X1 U146 ( .A1(n816), .A2(n815), .ZN(n964) );
  AND2_X1 U146bar ( .A1(n816bar), .A2(n815bar), .ZN(n964bar);
  OR2_X1 U147 ( .A1(n814), .A2(n813), .ZN(n815) );
  AND2_X1 U147bar ( .A1(n814bar), .A2(n813bar), .ZN(n815bar);
  OR2_X1 U148 ( .A1(n812), .A2(n811), .ZN(n813) );
  AND2_X1 U148bar ( .A1(n812bar), .A2(n811bar), .ZN(n813bar);
  OR2_X1 U149 ( .A1(in[122]), .A2(in[111]), .ZN(n811) );
  AND2_X1 U149bar ( .A1(inbar[122]), .A2(inbar[111]), .ZN(n811bar);
  OR2_X1 U150 ( .A1(in[154]), .A2(in[151]), .ZN(n812) );
  AND2_X1 U150bar ( .A1(inbar[154]), .A2(inbar[151]), .ZN(n812bar);
  OR2_X1 U151 ( .A1(n810), .A2(n809), .ZN(n814) );
  AND2_X1 U151bar ( .A1(n810bar), .A2(n809bar), .ZN(n814bar);
  OR2_X1 U152 ( .A1(in[187]), .A2(in[177]), .ZN(n809) );
  AND2_X1 U152bar ( .A1(inbar[187]), .A2(inbar[177]), .ZN(n809bar);
  OR2_X1 U153 ( .A1(in[200]), .A2(in[192]), .ZN(n810) );
  AND2_X1 U153bar ( .A1(inbar[200]), .A2(inbar[192]), .ZN(n810bar);
  OR2_X1 U154 ( .A1(n808), .A2(n807), .ZN(n816) );
  AND2_X1 U154bar ( .A1(n808bar), .A2(n807bar), .ZN(n816bar);
  OR2_X1 U155 ( .A1(n806), .A2(n805), .ZN(n807) );
  AND2_X1 U155bar ( .A1(n806bar), .A2(n805bar), .ZN(n807bar);
  OR2_X1 U156 ( .A1(in[225]), .A2(in[207]), .ZN(n805) );
  AND2_X1 U156bar ( .A1(inbar[225]), .A2(inbar[207]), .ZN(n805bar);
  OR2_X1 U157 ( .A1(in[98]), .A2(in[226]), .ZN(n806) );
  AND2_X1 U157bar ( .A1(inbar[98]), .A2(inbar[226]), .ZN(n806bar);
  OR2_X1 U158 ( .A1(n804), .A2(n803), .ZN(n808) );
  AND2_X1 U158bar ( .A1(n804bar), .A2(n803bar), .ZN(n808bar);
  OR2_X1 U159 ( .A1(in_20), .A2(in_16), .ZN(n803) );
  AND2_X1 U159bar ( .A1(in_20bar), .A2(in_16bar), .ZN(n803bar);
  OR2_X1 U160 ( .A1(in_55), .A2(in_45), .ZN(n804) );
  AND2_X1 U160bar ( .A1(in_55bar), .A2(in_45bar), .ZN(n804bar);
  OR2_X1 U161 ( .A1(n802), .A2(n801), .ZN(n824) );
  AND2_X1 U161bar ( .A1(n802bar), .A2(n801bar), .ZN(n824bar);
  OR2_X1 U162 ( .A1(in[162]), .A2(in[149]), .ZN(n801) );
  AND2_X1 U162bar ( .A1(inbar[162]), .A2(inbar[149]), .ZN(n801bar);
  OR2_X1 U163 ( .A1(in[163]), .A2(n800), .ZN(n802) );
  AND2_X1 U163bar ( .A1(inbar[163]), .A2(n800bar), .ZN(n802bar);
  OR2_X1 U164 ( .A1(in[191]), .A2(in[189]), .ZN(n800) );
  AND2_X1 U164bar ( .A1(inbar[191]), .A2(inbar[189]), .ZN(n800bar);
  OR2_X1 U165 ( .A1(n799), .A2(n798), .ZN(n826) );
  AND2_X1 U165bar ( .A1(n799bar), .A2(n798bar), .ZN(n826bar);
  OR2_X1 U166 ( .A1(n797), .A2(n796), .ZN(n798) );
  AND2_X1 U166bar ( .A1(n797bar), .A2(n796bar), .ZN(n798bar);
  OR2_X1 U167 ( .A1(in[212]), .A2(in[193]), .ZN(n796) );
  AND2_X1 U167bar ( .A1(inbar[212]), .A2(inbar[193]), .ZN(n796bar);
  OR2_X1 U168 ( .A1(in[238]), .A2(n795), .ZN(n797) );
  AND2_X1 U168bar ( .A1(inbar[238]), .A2(n795bar), .ZN(n797bar);
  OR2_X1 U169 ( .A1(in[88]), .A2(in[247]), .ZN(n795) );
  AND2_X1 U169bar ( .A1(inbar[88]), .A2(inbar[247]), .ZN(n795bar);
  OR2_X1 U170 ( .A1(n794), .A2(n793), .ZN(n799) );
  AND2_X1 U170bar ( .A1(n794bar), .A2(n793bar), .ZN(n799bar);
  OR2_X1 U171 ( .A1(in[94]), .A2(in[92]), .ZN(n793) );
  AND2_X1 U171bar ( .A1(inbar[94]), .A2(inbar[92]), .ZN(n793bar);
  OR2_X1 U172 ( .A1(in_52), .A2(n792), .ZN(n794) );
  AND2_X1 U172bar ( .A1(in_52bar), .A2(n792bar), .ZN(n794bar);
  OR2_X1 U173 ( .A1(in_70), .A2(in_67), .ZN(n792) );
  AND2_X1 U173bar ( .A1(in_70bar), .A2(in_67bar), .ZN(n792bar);
  OR2_X1 U174 ( .A1(n791), .A2(n790), .ZN(out[2]) );
  AND2_X1 U174bar ( .A1(n791bar), .A2(n790bar), .ZN(outbar[2]);
  OR2_X1 U175 ( .A1(n789), .A2(n788), .ZN(n790) );
  AND2_X1 U175bar ( .A1(n789bar), .A2(n788bar), .ZN(n790bar);
  OR2_X1 U176 ( .A1(n787), .A2(n786), .ZN(n788) );
  AND2_X1 U176bar ( .A1(n787bar), .A2(n786bar), .ZN(n788bar);
  OR2_X1 U177 ( .A1(n819), .A2(n785), .ZN(n786) );
  AND2_X1 U177bar ( .A1(n819bar), .A2(n785bar), .ZN(n786bar);
  OR2_X1 U178 ( .A1(n784), .A2(n783), .ZN(n819) );
  AND2_X1 U178bar ( .A1(n784bar), .A2(n783bar), .ZN(n819bar);
  OR2_X1 U179 ( .A1(n782), .A2(n781), .ZN(n783) );
  AND2_X1 U179bar ( .A1(n782bar), .A2(n781bar), .ZN(n783bar);
  OR2_X1 U180 ( .A1(n780), .A2(n779), .ZN(n781) );
  AND2_X1 U180bar ( .A1(n780bar), .A2(n779bar), .ZN(n781bar);
  OR2_X1 U181 ( .A1(n962), .A2(n778), .ZN(n779) );
  AND2_X1 U181bar ( .A1(n962bar), .A2(n778bar), .ZN(n779bar);
  OR2_X1 U182 ( .A1(n777), .A2(n776), .ZN(n962) );
  AND2_X1 U182bar ( .A1(n777bar), .A2(n776bar), .ZN(n962bar);
  OR2_X1 U183 ( .A1(n775), .A2(n774), .ZN(n776) );
  AND2_X1 U183bar ( .A1(n775bar), .A2(n774bar), .ZN(n776bar);
  OR2_X1 U184 ( .A1(n773), .A2(n772), .ZN(n774) );
  AND2_X1 U184bar ( .A1(n773bar), .A2(n772bar), .ZN(n774bar);
  OR2_X1 U185 ( .A1(in[131]), .A2(in[120]), .ZN(n772) );
  AND2_X1 U185bar ( .A1(inbar[131]), .A2(inbar[120]), .ZN(n772bar);
  OR2_X1 U186 ( .A1(in[153]), .A2(in[147]), .ZN(n773) );
  AND2_X1 U186bar ( .A1(inbar[153]), .A2(inbar[147]), .ZN(n773bar);
  OR2_X1 U187 ( .A1(n771), .A2(n770), .ZN(n775) );
  AND2_X1 U187bar ( .A1(n771bar), .A2(n770bar), .ZN(n775bar);
  OR2_X1 U188 ( .A1(in[170]), .A2(in[156]), .ZN(n770) );
  AND2_X1 U188bar ( .A1(inbar[170]), .A2(inbar[156]), .ZN(n770bar);
  OR2_X1 U189 ( .A1(in[223]), .A2(in[190]), .ZN(n771) );
  AND2_X1 U189bar ( .A1(inbar[223]), .A2(inbar[190]), .ZN(n771bar);
  OR2_X1 U190 ( .A1(n769), .A2(n768), .ZN(n777) );
  AND2_X1 U190bar ( .A1(n769bar), .A2(n768bar), .ZN(n777bar);
  OR2_X1 U191 ( .A1(n767), .A2(n766), .ZN(n768) );
  AND2_X1 U191bar ( .A1(n767bar), .A2(n766bar), .ZN(n768bar);
  OR2_X1 U192 ( .A1(in[236]), .A2(in[230]), .ZN(n766) );
  AND2_X1 U192bar ( .A1(inbar[236]), .A2(inbar[230]), .ZN(n766bar);
  OR2_X1 U193 ( .A1(in[85]), .A2(in[240]), .ZN(n767) );
  AND2_X1 U193bar ( .A1(inbar[85]), .A2(inbar[240]), .ZN(n767bar);
  OR2_X1 U194 ( .A1(n765), .A2(n764), .ZN(n769) );
  AND2_X1 U194bar ( .A1(n765bar), .A2(n764bar), .ZN(n769bar);
  OR2_X1 U195 ( .A1(in_12), .A2(in[90]), .ZN(n764) );
  AND2_X1 U195bar ( .A1(in_12bar), .A2(inbar[90]), .ZN(n764bar);
  OR2_X1 U196 ( .A1(in_39), .A2(in_28), .ZN(n765) );
  AND2_X1 U196bar ( .A1(in_39bar), .A2(in_28bar), .ZN(n765bar);
  OR2_X1 U197 ( .A1(in[109]), .A2(n763), .ZN(n780) );
  AND2_X1 U197bar ( .A1(inbar[109]), .A2(n763bar), .ZN(n780bar);
  OR2_X1 U198 ( .A1(n762), .A2(n761), .ZN(n782) );
  AND2_X1 U198bar ( .A1(n762bar), .A2(n761bar), .ZN(n782bar);
  OR2_X1 U199 ( .A1(in[138]), .A2(in[129]), .ZN(n761) );
  AND2_X1 U199bar ( .A1(inbar[138]), .A2(inbar[129]), .ZN(n761bar);
  OR2_X1 U200 ( .A1(in[157]), .A2(n760), .ZN(n762) );
  AND2_X1 U200bar ( .A1(inbar[157]), .A2(n760bar), .ZN(n762bar);
  OR2_X1 U201 ( .A1(in[182]), .A2(in[167]), .ZN(n760) );
  AND2_X1 U201bar ( .A1(inbar[182]), .A2(inbar[167]), .ZN(n760bar);
  OR2_X1 U202 ( .A1(n759), .A2(n758), .ZN(n784) );
  AND2_X1 U202bar ( .A1(n759bar), .A2(n758bar), .ZN(n784bar);
  OR2_X1 U203 ( .A1(n757), .A2(n756), .ZN(n758) );
  AND2_X1 U203bar ( .A1(n757bar), .A2(n756bar), .ZN(n758bar);
  OR2_X1 U204 ( .A1(in[195]), .A2(in[184]), .ZN(n756) );
  AND2_X1 U204bar ( .A1(inbar[195]), .A2(inbar[184]), .ZN(n756bar);
  OR2_X1 U205 ( .A1(in[196]), .A2(n755), .ZN(n757) );
  AND2_X1 U205bar ( .A1(inbar[196]), .A2(n755bar), .ZN(n757bar);
  OR2_X1 U206 ( .A1(in[215]), .A2(in[209]), .ZN(n755) );
  AND2_X1 U206bar ( .A1(inbar[215]), .A2(inbar[209]), .ZN(n755bar);
  OR2_X1 U207 ( .A1(n754), .A2(n753), .ZN(n759) );
  AND2_X1 U207bar ( .A1(n754bar), .A2(n753bar), .ZN(n759bar);
  OR2_X1 U208 ( .A1(in[93]), .A2(in[233]), .ZN(n753) );
  AND2_X1 U208bar ( .A1(inbar[93]), .A2(inbar[233]), .ZN(n753bar);
  OR2_X1 U209 ( .A1(in_1), .A2(n752), .ZN(n754) );
  AND2_X1 U209bar ( .A1(in_1bar), .A2(n752bar), .ZN(n754bar);
  OR2_X1 U210 ( .A1(in_69), .A2(in_66), .ZN(n752) );
  AND2_X1 U210bar ( .A1(in_69bar), .A2(in_66bar), .ZN(n752bar);
  OR2_X1 U211 ( .A1(n966), .A2(n751), .ZN(n787) );
  AND2_X1 U211bar ( .A1(n966bar), .A2(n751bar), .ZN(n787bar);
  OR2_X1 U212 ( .A1(in[134]), .A2(n750), .ZN(n751) );
  AND2_X1 U212bar ( .A1(inbar[134]), .A2(n750bar), .ZN(n751bar);
  OR2_X1 U213 ( .A1(n749), .A2(n748), .ZN(n966) );
  AND2_X1 U213bar ( .A1(n749bar), .A2(n748bar), .ZN(n966bar);
  OR2_X1 U214 ( .A1(n747), .A2(n746), .ZN(n748) );
  AND2_X1 U214bar ( .A1(n747bar), .A2(n746bar), .ZN(n748bar);
  OR2_X1 U215 ( .A1(n745), .A2(n744), .ZN(n746) );
  AND2_X1 U215bar ( .A1(n745bar), .A2(n744bar), .ZN(n746bar);
  OR2_X1 U216 ( .A1(in[136]), .A2(in[121]), .ZN(n744) );
  AND2_X1 U216bar ( .A1(inbar[136]), .A2(inbar[121]), .ZN(n744bar);
  OR2_X1 U217 ( .A1(in[186]), .A2(in[174]), .ZN(n745) );
  AND2_X1 U217bar ( .A1(inbar[186]), .A2(inbar[174]), .ZN(n745bar);
  OR2_X1 U218 ( .A1(n743), .A2(n742), .ZN(n747) );
  AND2_X1 U218bar ( .A1(n743bar), .A2(n742bar), .ZN(n747bar);
  OR2_X1 U219 ( .A1(in[198]), .A2(in[197]), .ZN(n742) );
  AND2_X1 U219bar ( .A1(inbar[198]), .A2(inbar[197]), .ZN(n742bar);
  OR2_X1 U220 ( .A1(in[214]), .A2(in[199]), .ZN(n743) );
  AND2_X1 U220bar ( .A1(inbar[214]), .A2(inbar[199]), .ZN(n743bar);
  OR2_X1 U221 ( .A1(n741), .A2(n740), .ZN(n749) );
  AND2_X1 U221bar ( .A1(n741bar), .A2(n740bar), .ZN(n749bar);
  OR2_X1 U222 ( .A1(n739), .A2(n738), .ZN(n740) );
  AND2_X1 U222bar ( .A1(n739bar), .A2(n738bar), .ZN(n740bar);
  OR2_X1 U223 ( .A1(in[231]), .A2(in[220]), .ZN(n738) );
  AND2_X1 U223bar ( .A1(inbar[231]), .A2(inbar[220]), .ZN(n738bar);
  OR2_X1 U224 ( .A1(in_25), .A2(in[245]), .ZN(n739) );
  AND2_X1 U224bar ( .A1(in_25bar), .A2(inbar[245]), .ZN(n739bar);
  OR2_X1 U225 ( .A1(n737), .A2(n736), .ZN(n741) );
  AND2_X1 U225bar ( .A1(n737bar), .A2(n736bar), .ZN(n741bar);
  OR2_X1 U226 ( .A1(in_53), .A2(in_29), .ZN(n736) );
  AND2_X1 U226bar ( .A1(in_53bar), .A2(in_29bar), .ZN(n736bar);
  OR2_X1 U227 ( .A1(in_79), .A2(in_74), .ZN(n737) );
  AND2_X1 U227bar ( .A1(in_79bar), .A2(in_74bar), .ZN(n737bar);
  OR2_X1 U228 ( .A1(n735), .A2(n734), .ZN(n789) );
  AND2_X1 U228bar ( .A1(n735bar), .A2(n734bar), .ZN(n789bar);
  OR2_X1 U229 ( .A1(in[152]), .A2(in[140]), .ZN(n734) );
  AND2_X1 U229bar ( .A1(inbar[152]), .A2(inbar[140]), .ZN(n734bar);
  OR2_X1 U230 ( .A1(in[155]), .A2(n733), .ZN(n735) );
  AND2_X1 U230bar ( .A1(inbar[155]), .A2(n733bar), .ZN(n735bar);
  OR2_X1 U231 ( .A1(in[166]), .A2(in[165]), .ZN(n733) );
  AND2_X1 U231bar ( .A1(inbar[166]), .A2(inbar[165]), .ZN(n733bar);
  OR2_X1 U232 ( .A1(n732), .A2(n731), .ZN(n791) );
  AND2_X1 U232bar ( .A1(n732bar), .A2(n731bar), .ZN(n791bar);
  OR2_X1 U233 ( .A1(n730), .A2(n729), .ZN(n731) );
  AND2_X1 U233bar ( .A1(n730bar), .A2(n729bar), .ZN(n731bar);
  OR2_X1 U234 ( .A1(in[202]), .A2(in[185]), .ZN(n729) );
  AND2_X1 U234bar ( .A1(inbar[202]), .A2(inbar[185]), .ZN(n729bar);
  OR2_X1 U235 ( .A1(in[211]), .A2(n728), .ZN(n730) );
  AND2_X1 U235bar ( .A1(inbar[211]), .A2(n728bar), .ZN(n730bar);
  OR2_X1 U236 ( .A1(in[255]), .A2(in[253]), .ZN(n728) );
  AND2_X1 U236bar ( .A1(inbar[255]), .A2(inbar[253]), .ZN(n728bar);
  OR2_X1 U237 ( .A1(n727), .A2(n726), .ZN(n732) );
  AND2_X1 U237bar ( .A1(n727bar), .A2(n726bar), .ZN(n732bar);
  OR2_X1 U238 ( .A1(in_35), .A2(in_15), .ZN(n726) );
  AND2_X1 U238bar ( .A1(in_35bar), .A2(in_15bar), .ZN(n726bar);
  OR2_X1 U239 ( .A1(in_36), .A2(n725), .ZN(n727) );
  AND2_X1 U239bar ( .A1(in_36bar), .A2(n725bar), .ZN(n727bar);
  OR2_X1 U240 ( .A1(in_48), .A2(in_40), .ZN(n725) );
  AND2_X1 U240bar ( .A1(in_48bar), .A2(in_40bar), .ZN(n725bar);
  OR2_X1 U241 ( .A1(n724), .A2(n723), .ZN(out[1]) );
  AND2_X1 U241bar ( .A1(n724bar), .A2(n723bar), .ZN(outbar[1]);
  OR2_X1 U242 ( .A1(n722), .A2(n721), .ZN(n723) );
  AND2_X1 U242bar ( .A1(n722bar), .A2(n721bar), .ZN(n723bar);
  OR2_X1 U243 ( .A1(n720), .A2(n719), .ZN(n721) );
  AND2_X1 U243bar ( .A1(n720bar), .A2(n719bar), .ZN(n721bar);
  OR2_X1 U244 ( .A1(n921), .A2(n887), .ZN(n719) );
  AND2_X1 U244bar ( .A1(n921bar), .A2(n887bar), .ZN(n719bar);
  OR2_X1 U245 ( .A1(n718), .A2(n717), .ZN(n887) );
  AND2_X1 U245bar ( .A1(n718bar), .A2(n717bar), .ZN(n887bar);
  OR2_X1 U246 ( .A1(n716), .A2(n715), .ZN(n717) );
  AND2_X1 U246bar ( .A1(n716bar), .A2(n715bar), .ZN(n717bar);
  OR2_X1 U247 ( .A1(n714), .A2(n713), .ZN(n715) );
  AND2_X1 U247bar ( .A1(n714bar), .A2(n713bar), .ZN(n715bar);
  OR2_X1 U248 ( .A1(in[116]), .A2(in[110]), .ZN(n713) );
  AND2_X1 U248bar ( .A1(inbar[116]), .A2(inbar[110]), .ZN(n713bar);
  OR2_X1 U249 ( .A1(in[133]), .A2(in[130]), .ZN(n714) );
  AND2_X1 U249bar ( .A1(inbar[133]), .A2(inbar[130]), .ZN(n714bar);
  OR2_X1 U250 ( .A1(n712), .A2(n711), .ZN(n716) );
  AND2_X1 U250bar ( .A1(n712bar), .A2(n711bar), .ZN(n716bar);
  OR2_X1 U251 ( .A1(in[203]), .A2(in[135]), .ZN(n711) );
  AND2_X1 U251bar ( .A1(inbar[203]), .A2(inbar[135]), .ZN(n711bar);
  OR2_X1 U252 ( .A1(in[232]), .A2(in[223]), .ZN(n712) );
  AND2_X1 U252bar ( .A1(inbar[232]), .A2(inbar[223]), .ZN(n712bar);
  OR2_X1 U253 ( .A1(n710), .A2(n709), .ZN(n718) );
  AND2_X1 U253bar ( .A1(n710bar), .A2(n709bar), .ZN(n718bar);
  OR2_X1 U254 ( .A1(n708), .A2(n707), .ZN(n709) );
  AND2_X1 U254bar ( .A1(n708bar), .A2(n707bar), .ZN(n709bar);
  OR2_X1 U255 ( .A1(in[255]), .A2(in[233]), .ZN(n707) );
  AND2_X1 U255bar ( .A1(inbar[255]), .A2(inbar[233]), .ZN(n707bar);
  OR2_X1 U256 ( .A1(in_53), .A2(in_34), .ZN(n708) );
  AND2_X1 U256bar ( .A1(in_53bar), .A2(in_34bar), .ZN(n708bar);
  OR2_X1 U257 ( .A1(n706), .A2(n705), .ZN(n710) );
  AND2_X1 U257bar ( .A1(n706bar), .A2(n705bar), .ZN(n710bar);
  OR2_X1 U258 ( .A1(in_57), .A2(in_55), .ZN(n705) );
  AND2_X1 U258bar ( .A1(in_57bar), .A2(in_55bar), .ZN(n705bar);
  OR2_X1 U259 ( .A1(in_68), .A2(in_67), .ZN(n706) );
  AND2_X1 U259bar ( .A1(in_68bar), .A2(in_67bar), .ZN(n706bar);
  OR2_X1 U260 ( .A1(n704), .A2(n703), .ZN(n921) );
  AND2_X1 U260bar ( .A1(n704bar), .A2(n703bar), .ZN(n921bar);
  OR2_X1 U261 ( .A1(n702), .A2(n701), .ZN(n703) );
  AND2_X1 U261bar ( .A1(n702bar), .A2(n701bar), .ZN(n703bar);
  OR2_X1 U262 ( .A1(n700), .A2(n699), .ZN(n701) );
  AND2_X1 U262bar ( .A1(n700bar), .A2(n699bar), .ZN(n701bar);
  OR2_X1 U263 ( .A1(n944), .A2(n872), .ZN(n699) );
  AND2_X1 U263bar ( .A1(n944bar), .A2(n872bar), .ZN(n699bar);
  OR2_X1 U264 ( .A1(n698), .A2(n697), .ZN(n872) );
  AND2_X1 U264bar ( .A1(n698bar), .A2(n697bar), .ZN(n872bar);
  OR2_X1 U265 ( .A1(n696), .A2(n695), .ZN(n697) );
  AND2_X1 U265bar ( .A1(n696bar), .A2(n695bar), .ZN(n697bar);
  OR2_X1 U266 ( .A1(n694), .A2(n693), .ZN(n695) );
  AND2_X1 U266bar ( .A1(n694bar), .A2(n693bar), .ZN(n695bar);
  OR2_X1 U267 ( .A1(in[121]), .A2(in[102]), .ZN(n693) );
  AND2_X1 U267bar ( .A1(inbar[121]), .A2(inbar[102]), .ZN(n693bar);
  OR2_X1 U268 ( .A1(in[162]), .A2(in[161]), .ZN(n694) );
  AND2_X1 U268bar ( .A1(inbar[162]), .A2(inbar[161]), .ZN(n694bar);
  OR2_X1 U269 ( .A1(n692), .A2(n691), .ZN(n696) );
  AND2_X1 U269bar ( .A1(n692bar), .A2(n691bar), .ZN(n696bar);
  OR2_X1 U270 ( .A1(in[192]), .A2(in[178]), .ZN(n691) );
  AND2_X1 U270bar ( .A1(inbar[192]), .A2(inbar[178]), .ZN(n691bar);
  OR2_X1 U271 ( .A1(in[244]), .A2(in[209]), .ZN(n692) );
  AND2_X1 U271bar ( .A1(inbar[244]), .A2(inbar[209]), .ZN(n692bar);
  OR2_X1 U272 ( .A1(n690), .A2(n689), .ZN(n698) );
  AND2_X1 U272bar ( .A1(n690bar), .A2(n689bar), .ZN(n698bar);
  OR2_X1 U273 ( .A1(n688), .A2(n687), .ZN(n689) );
  AND2_X1 U273bar ( .A1(n688bar), .A2(n687bar), .ZN(n689bar);
  OR2_X1 U274 ( .A1(in[90]), .A2(in[254]), .ZN(n687) );
  AND2_X1 U274bar ( .A1(inbar[90]), .A2(inbar[254]), .ZN(n687bar);
  OR2_X1 U275 ( .A1(in_36), .A2(in_32), .ZN(n688) );
  AND2_X1 U275bar ( .A1(in_36bar), .A2(in_32bar), .ZN(n688bar);
  OR2_X1 U276 ( .A1(n686), .A2(n685), .ZN(n690) );
  AND2_X1 U276bar ( .A1(n686bar), .A2(n685bar), .ZN(n690bar);
  OR2_X1 U277 ( .A1(in_62), .A2(in_37), .ZN(n685) );
  AND2_X1 U277bar ( .A1(in_62bar), .A2(in_37bar), .ZN(n685bar);
  OR2_X1 U278 ( .A1(in_75), .A2(in_73), .ZN(n686) );
  AND2_X1 U278bar ( .A1(in_75bar), .A2(in_73bar), .ZN(n686bar);
  OR2_X1 U279 ( .A1(n684), .A2(n683), .ZN(n944) );
  AND2_X1 U279bar ( .A1(n684bar), .A2(n683bar), .ZN(n944bar);
  OR2_X1 U280 ( .A1(n682), .A2(n681), .ZN(n683) );
  AND2_X1 U280bar ( .A1(n682bar), .A2(n681bar), .ZN(n683bar);
  OR2_X1 U281 ( .A1(n680), .A2(n679), .ZN(n681) );
  AND2_X1 U281bar ( .A1(n680bar), .A2(n679bar), .ZN(n681bar);
  OR2_X1 U282 ( .A1(in[171]), .A2(in[153]), .ZN(n679) );
  AND2_X1 U282bar ( .A1(inbar[171]), .A2(inbar[153]), .ZN(n679bar);
  OR2_X1 U283 ( .A1(in[187]), .A2(in[176]), .ZN(n680) );
  AND2_X1 U283bar ( .A1(inbar[187]), .A2(inbar[176]), .ZN(n680bar);
  OR2_X1 U284 ( .A1(n678), .A2(n677), .ZN(n682) );
  AND2_X1 U284bar ( .A1(n678bar), .A2(n677bar), .ZN(n682bar);
  OR2_X1 U285 ( .A1(in[245]), .A2(in[211]), .ZN(n677) );
  AND2_X1 U285bar ( .A1(inbar[245]), .A2(inbar[211]), .ZN(n677bar);
  OR2_X1 U286 ( .A1(in[97]), .A2(in[88]), .ZN(n678) );
  AND2_X1 U286bar ( .A1(inbar[97]), .A2(inbar[88]), .ZN(n678bar);
  OR2_X1 U287 ( .A1(n676), .A2(n675), .ZN(n684) );
  AND2_X1 U287bar ( .A1(n676bar), .A2(n675bar), .ZN(n684bar);
  OR2_X1 U288 ( .A1(n674), .A2(n673), .ZN(n675) );
  AND2_X1 U288bar ( .A1(n674bar), .A2(n673bar), .ZN(n675bar);
  OR2_X1 U289 ( .A1(in_10), .A2(in_0), .ZN(n673) );
  AND2_X1 U289bar ( .A1(in_10bar), .A2(in_0bar), .ZN(n673bar);
  OR2_X1 U290 ( .A1(in_59), .A2(in_5), .ZN(n674) );
  AND2_X1 U290bar ( .A1(in_59bar), .A2(in_5bar), .ZN(n674bar);
  OR2_X1 U291 ( .A1(n672), .A2(n671), .ZN(n676) );
  AND2_X1 U291bar ( .A1(n672bar), .A2(n671bar), .ZN(n676bar);
  OR2_X1 U292 ( .A1(in_60), .A2(in_6), .ZN(n671) );
  AND2_X1 U292bar ( .A1(in_60bar), .A2(in_6bar), .ZN(n671bar);
  OR2_X1 U293 ( .A1(in_77), .A2(in_69), .ZN(n672) );
  AND2_X1 U293bar ( .A1(in_77bar), .A2(in_69bar), .ZN(n672bar);
  OR2_X1 U294 ( .A1(in[113]), .A2(n864), .ZN(n700) );
  AND2_X1 U294bar ( .A1(inbar[113]), .A2(n864bar), .ZN(n700bar);
  OR2_X1 U295 ( .A1(n670), .A2(n669), .ZN(n864) );
  AND2_X1 U295bar ( .A1(n670bar), .A2(n669bar), .ZN(n864bar);
  OR2_X1 U296 ( .A1(n668), .A2(n667), .ZN(n669) );
  AND2_X1 U296bar ( .A1(n668bar), .A2(n667bar), .ZN(n669bar);
  OR2_X1 U297 ( .A1(n666), .A2(n665), .ZN(n667) );
  AND2_X1 U297bar ( .A1(n666bar), .A2(n665bar), .ZN(n667bar);
  OR2_X1 U298 ( .A1(in[125]), .A2(in[107]), .ZN(n665) );
  AND2_X1 U298bar ( .A1(inbar[125]), .A2(inbar[107]), .ZN(n665bar);
  OR2_X1 U299 ( .A1(in[138]), .A2(in[126]), .ZN(n666) );
  AND2_X1 U299bar ( .A1(inbar[138]), .A2(inbar[126]), .ZN(n666bar);
  OR2_X1 U300 ( .A1(n664), .A2(n663), .ZN(n668) );
  AND2_X1 U300bar ( .A1(n664bar), .A2(n663bar), .ZN(n668bar);
  OR2_X1 U301 ( .A1(in[189]), .A2(in[143]), .ZN(n663) );
  AND2_X1 U301bar ( .A1(inbar[189]), .A2(inbar[143]), .ZN(n663bar);
  OR2_X1 U302 ( .A1(in[99]), .A2(in[214]), .ZN(n664) );
  AND2_X1 U302bar ( .A1(inbar[99]), .A2(inbar[214]), .ZN(n664bar);
  OR2_X1 U303 ( .A1(n662), .A2(n661), .ZN(n670) );
  AND2_X1 U303bar ( .A1(n662bar), .A2(n661bar), .ZN(n670bar);
  OR2_X1 U304 ( .A1(n660), .A2(n659), .ZN(n661) );
  AND2_X1 U304bar ( .A1(n660bar), .A2(n659bar), .ZN(n661bar);
  OR2_X1 U305 ( .A1(in_15), .A2(in_12), .ZN(n659) );
  AND2_X1 U305bar ( .A1(in_15bar), .A2(in_12bar), .ZN(n659bar);
  OR2_X1 U306 ( .A1(in_20), .A2(in_2), .ZN(n660) );
  AND2_X1 U306bar ( .A1(in_20bar), .A2(in_2bar), .ZN(n660bar);
  OR2_X1 U307 ( .A1(n658), .A2(n657), .ZN(n662) );
  AND2_X1 U307bar ( .A1(n658bar), .A2(n657bar), .ZN(n662bar);
  OR2_X1 U308 ( .A1(in_30), .A2(in_3), .ZN(n657) );
  AND2_X1 U308bar ( .A1(in_30bar), .A2(in_3bar), .ZN(n657bar);
  OR2_X1 U309 ( .A1(in_4), .A2(in_38), .ZN(n658) );
  AND2_X1 U309bar ( .A1(in_4bar), .A2(in_38bar), .ZN(n658bar);
  OR2_X1 U310 ( .A1(n656), .A2(n655), .ZN(n702) );
  AND2_X1 U310bar ( .A1(n656bar), .A2(n655bar), .ZN(n702bar);
  OR2_X1 U311 ( .A1(in[148]), .A2(in[137]), .ZN(n655) );
  AND2_X1 U311bar ( .A1(inbar[148]), .A2(inbar[137]), .ZN(n655bar);
  OR2_X1 U312 ( .A1(in[149]), .A2(n654), .ZN(n656) );
  AND2_X1 U312bar ( .A1(inbar[149]), .A2(n654bar), .ZN(n656bar);
  OR2_X1 U313 ( .A1(in[195]), .A2(in[190]), .ZN(n654) );
  AND2_X1 U313bar ( .A1(inbar[195]), .A2(inbar[190]), .ZN(n654bar);
  OR2_X1 U314 ( .A1(n653), .A2(n652), .ZN(n704) );
  AND2_X1 U314bar ( .A1(n653bar), .A2(n652bar), .ZN(n704bar);
  OR2_X1 U315 ( .A1(n651), .A2(n650), .ZN(n652) );
  AND2_X1 U315bar ( .A1(n651bar), .A2(n650bar), .ZN(n652bar);
  OR2_X1 U316 ( .A1(in[98]), .A2(in[197]), .ZN(n650) );
  AND2_X1 U316bar ( .A1(inbar[98]), .A2(inbar[197]), .ZN(n650bar);
  OR2_X1 U317 ( .A1(in_11), .A2(n649), .ZN(n651) );
  AND2_X1 U317bar ( .A1(in_11bar), .A2(n649bar), .ZN(n651bar);
  OR2_X1 U318 ( .A1(in_26), .A2(in_14), .ZN(n649) );
  AND2_X1 U318bar ( .A1(in_26bar), .A2(in_14bar), .ZN(n649bar);
  OR2_X1 U319 ( .A1(n648), .A2(n647), .ZN(n653) );
  AND2_X1 U319bar ( .A1(n648bar), .A2(n647bar), .ZN(n653bar);
  OR2_X1 U320 ( .A1(in_35), .A2(in_27), .ZN(n647) );
  AND2_X1 U320bar ( .A1(in_35bar), .A2(in_27bar), .ZN(n647bar);
  OR2_X1 U321 ( .A1(in_50), .A2(n646), .ZN(n648) );
  AND2_X1 U321bar ( .A1(in_50bar), .A2(n646bar), .ZN(n648bar);
  OR2_X1 U322 ( .A1(in_78), .A2(in_61), .ZN(n646) );
  AND2_X1 U322bar ( .A1(in_78bar), .A2(in_61bar), .ZN(n646bar);
  OR2_X1 U323 ( .A1(n942), .A2(n645), .ZN(n720) );
  AND2_X1 U323bar ( .A1(n942bar), .A2(n645bar), .ZN(n720bar);
  OR2_X1 U324 ( .A1(in[106]), .A2(n863), .ZN(n645) );
  AND2_X1 U324bar ( .A1(inbar[106]), .A2(n863bar), .ZN(n645bar);
  OR2_X1 U325 ( .A1(n644), .A2(n643), .ZN(n863) );
  AND2_X1 U325bar ( .A1(n644bar), .A2(n643bar), .ZN(n863bar);
  OR2_X1 U326 ( .A1(n642), .A2(n641), .ZN(n643) );
  AND2_X1 U326bar ( .A1(n642bar), .A2(n641bar), .ZN(n643bar);
  OR2_X1 U327 ( .A1(n640), .A2(n639), .ZN(n641) );
  AND2_X1 U327bar ( .A1(n640bar), .A2(n639bar), .ZN(n641bar);
  OR2_X1 U328 ( .A1(in[127]), .A2(in[122]), .ZN(n639) );
  AND2_X1 U328bar ( .A1(inbar[127]), .A2(inbar[122]), .ZN(n639bar);
  OR2_X1 U329 ( .A1(in[156]), .A2(in[132]), .ZN(n640) );
  AND2_X1 U329bar ( .A1(inbar[156]), .A2(inbar[132]), .ZN(n640bar);
  OR2_X1 U330 ( .A1(n638), .A2(n637), .ZN(n642) );
  AND2_X1 U330bar ( .A1(n638bar), .A2(n637bar), .ZN(n642bar);
  OR2_X1 U331 ( .A1(in[159]), .A2(in[157]), .ZN(n637) );
  AND2_X1 U331bar ( .A1(inbar[159]), .A2(inbar[157]), .ZN(n637bar);
  OR2_X1 U332 ( .A1(in[185]), .A2(in[169]), .ZN(n638) );
  AND2_X1 U332bar ( .A1(inbar[185]), .A2(inbar[169]), .ZN(n638bar);
  OR2_X1 U333 ( .A1(n636), .A2(n635), .ZN(n644) );
  AND2_X1 U333bar ( .A1(n636bar), .A2(n635bar), .ZN(n644bar);
  OR2_X1 U334 ( .A1(n634), .A2(n633), .ZN(n635) );
  AND2_X1 U334bar ( .A1(n634bar), .A2(n633bar), .ZN(n635bar);
  OR2_X1 U335 ( .A1(in[239]), .A2(in[218]), .ZN(n633) );
  AND2_X1 U335bar ( .A1(inbar[239]), .A2(inbar[218]), .ZN(n633bar);
  OR2_X1 U336 ( .A1(in_13), .A2(in[87]), .ZN(n634) );
  AND2_X1 U336bar ( .A1(in_13bar), .A2(inbar[87]), .ZN(n634bar);
  OR2_X1 U337 ( .A1(n632), .A2(n631), .ZN(n636) );
  AND2_X1 U337bar ( .A1(n632bar), .A2(n631bar), .ZN(n636bar);
  OR2_X1 U338 ( .A1(in_72), .A2(in_70), .ZN(n631) );
  AND2_X1 U338bar ( .A1(in_72bar), .A2(in_70bar), .ZN(n631bar);
  OR2_X1 U339 ( .A1(in_80), .A2(in_74), .ZN(n632) );
  AND2_X1 U339bar ( .A1(in_80bar), .A2(in_74bar), .ZN(n632bar);
  OR2_X1 U340 ( .A1(n630), .A2(n629), .ZN(n942) );
  AND2_X1 U340bar ( .A1(n630bar), .A2(n629bar), .ZN(n942bar);
  OR2_X1 U341 ( .A1(n628), .A2(n627), .ZN(n629) );
  AND2_X1 U341bar ( .A1(n628bar), .A2(n627bar), .ZN(n629bar);
  OR2_X1 U342 ( .A1(n626), .A2(n625), .ZN(n627) );
  AND2_X1 U342bar ( .A1(n626bar), .A2(n625bar), .ZN(n627bar);
  OR2_X1 U343 ( .A1(in[146]), .A2(in[100]), .ZN(n625) );
  AND2_X1 U343bar ( .A1(inbar[146]), .A2(inbar[100]), .ZN(n625bar);
  OR2_X1 U344 ( .A1(in[168]), .A2(in[152]), .ZN(n626) );
  AND2_X1 U344bar ( .A1(inbar[168]), .A2(inbar[152]), .ZN(n626bar);
  OR2_X1 U345 ( .A1(n624), .A2(n623), .ZN(n628) );
  AND2_X1 U345bar ( .A1(n624bar), .A2(n623bar), .ZN(n628bar);
  OR2_X1 U346 ( .A1(in[199]), .A2(in[182]), .ZN(n623) );
  AND2_X1 U346bar ( .A1(inbar[199]), .A2(inbar[182]), .ZN(n623bar);
  OR2_X1 U347 ( .A1(in[236]), .A2(in[204]), .ZN(n624) );
  AND2_X1 U347bar ( .A1(inbar[236]), .A2(inbar[204]), .ZN(n624bar);
  OR2_X1 U348 ( .A1(n622), .A2(n621), .ZN(n630) );
  AND2_X1 U348bar ( .A1(n622bar), .A2(n621bar), .ZN(n630bar);
  OR2_X1 U349 ( .A1(n620), .A2(n619), .ZN(n621) );
  AND2_X1 U349bar ( .A1(n620bar), .A2(n619bar), .ZN(n621bar);
  OR2_X1 U350 ( .A1(in[89]), .A2(in[246]), .ZN(n619) );
  AND2_X1 U350bar ( .A1(inbar[89]), .A2(inbar[246]), .ZN(n619bar);
  OR2_X1 U351 ( .A1(in[95]), .A2(in[92]), .ZN(n620) );
  AND2_X1 U351bar ( .A1(inbar[95]), .A2(inbar[92]), .ZN(n620bar);
  OR2_X1 U352 ( .A1(n618), .A2(n617), .ZN(n622) );
  AND2_X1 U352bar ( .A1(n618bar), .A2(n617bar), .ZN(n622bar);
  OR2_X1 U353 ( .A1(in_22), .A2(in_16), .ZN(n617) );
  AND2_X1 U353bar ( .A1(in_22bar), .A2(in_16bar), .ZN(n617bar);
  OR2_X1 U354 ( .A1(in_51), .A2(in_49), .ZN(n618) );
  AND2_X1 U354bar ( .A1(in_51bar), .A2(in_49bar), .ZN(n618bar);
  OR2_X1 U355 ( .A1(n616), .A2(n615), .ZN(n722) );
  AND2_X1 U355bar ( .A1(n616bar), .A2(n615bar), .ZN(n722bar);
  OR2_X1 U356 ( .A1(in[158]), .A2(in[115]), .ZN(n615) );
  AND2_X1 U356bar ( .A1(inbar[158]), .A2(inbar[115]), .ZN(n615bar);
  OR2_X1 U357 ( .A1(in[163]), .A2(n614), .ZN(n616) );
  AND2_X1 U357bar ( .A1(inbar[163]), .A2(n614bar), .ZN(n616bar);
  OR2_X1 U358 ( .A1(in[206]), .A2(in[165]), .ZN(n614) );
  AND2_X1 U358bar ( .A1(inbar[206]), .A2(inbar[165]), .ZN(n614bar);
  OR2_X1 U359 ( .A1(n613), .A2(n612), .ZN(n724) );
  AND2_X1 U359bar ( .A1(n613bar), .A2(n612bar), .ZN(n724bar);
  OR2_X1 U360 ( .A1(n611), .A2(n610), .ZN(n612) );
  AND2_X1 U360bar ( .A1(n611bar), .A2(n610bar), .ZN(n612bar);
  OR2_X1 U361 ( .A1(in[213]), .A2(in[207]), .ZN(n610) );
  AND2_X1 U361bar ( .A1(inbar[213]), .A2(inbar[207]), .ZN(n610bar);
  OR2_X1 U362 ( .A1(in[215]), .A2(n609), .ZN(n611) );
  AND2_X1 U362bar ( .A1(inbar[215]), .A2(n609bar), .ZN(n611bar);
  OR2_X1 U363 ( .A1(in[230]), .A2(in[220]), .ZN(n609) );
  AND2_X1 U363bar ( .A1(inbar[230]), .A2(inbar[220]), .ZN(n609bar);
  OR2_X1 U364 ( .A1(n608), .A2(n607), .ZN(n613) );
  AND2_X1 U364bar ( .A1(n608bar), .A2(n607bar), .ZN(n613bar);
  OR2_X1 U365 ( .A1(in[251]), .A2(in[234]), .ZN(n607) );
  AND2_X1 U365bar ( .A1(inbar[251]), .A2(inbar[234]), .ZN(n607bar);
  OR2_X1 U366 ( .A1(in_17), .A2(n606), .ZN(n608) );
  AND2_X1 U366bar ( .A1(in_17bar), .A2(n606bar), .ZN(n608bar);
  OR2_X1 U367 ( .A1(in_65), .A2(in_56), .ZN(n606) );
  AND2_X1 U367bar ( .A1(in_65bar), .A2(in_56bar), .ZN(n606bar);
  OR2_X1 U368 ( .A1(n605), .A2(n604), .ZN(out[0]) );
  AND2_X1 U368bar ( .A1(n605bar), .A2(n604bar), .ZN(outbar[0]);
  OR2_X1 U369 ( .A1(n603), .A2(n602), .ZN(n604) );
  AND2_X1 U369bar ( .A1(n603bar), .A2(n602bar), .ZN(n604bar);
  OR2_X1 U370 ( .A1(n601), .A2(n600), .ZN(n602) );
  AND2_X1 U370bar ( .A1(n601bar), .A2(n600bar), .ZN(n602bar);
  OR2_X1 U371 ( .A1(n820), .A2(n785), .ZN(n600) );
  AND2_X1 U371bar ( .A1(n820bar), .A2(n785bar), .ZN(n600bar);
  OR2_X1 U372 ( .A1(n599), .A2(n598), .ZN(n785) );
  AND2_X1 U372bar ( .A1(n599bar), .A2(n598bar), .ZN(n785bar);
  OR2_X1 U373 ( .A1(n597), .A2(n596), .ZN(n598) );
  AND2_X1 U373bar ( .A1(n597bar), .A2(n596bar), .ZN(n598bar);
  OR2_X1 U374 ( .A1(n595), .A2(n594), .ZN(n596) );
  AND2_X1 U374bar ( .A1(n595bar), .A2(n594bar), .ZN(n596bar);
  OR2_X1 U375 ( .A1(in[135]), .A2(in[104]), .ZN(n594) );
  AND2_X1 U375bar ( .A1(inbar[135]), .A2(inbar[104]), .ZN(n594bar);
  OR2_X1 U376 ( .A1(in[188]), .A2(in[178]), .ZN(n595) );
  AND2_X1 U376bar ( .A1(inbar[188]), .A2(inbar[178]), .ZN(n595bar);
  OR2_X1 U377 ( .A1(n593), .A2(n592), .ZN(n597) );
  AND2_X1 U377bar ( .A1(n593bar), .A2(n592bar), .ZN(n597bar);
  OR2_X1 U378 ( .A1(in[217]), .A2(in[194]), .ZN(n592) );
  AND2_X1 U378bar ( .A1(inbar[217]), .A2(inbar[194]), .ZN(n592bar);
  OR2_X1 U379 ( .A1(in[237]), .A2(in[218]), .ZN(n593) );
  AND2_X1 U379bar ( .A1(inbar[237]), .A2(inbar[218]), .ZN(n593bar);
  OR2_X1 U380 ( .A1(n591), .A2(n590), .ZN(n599) );
  AND2_X1 U380bar ( .A1(n591bar), .A2(n590bar), .ZN(n599bar);
  OR2_X1 U381 ( .A1(n589), .A2(n588), .ZN(n590) );
  AND2_X1 U381bar ( .A1(n589bar), .A2(n588bar), .ZN(n590bar);
  OR2_X1 U382 ( .A1(in_2), .A2(in_10), .ZN(n588) );
  AND2_X1 U382bar ( .A1(in_2bar), .A2(in_10bar), .ZN(n588bar);
  OR2_X1 U383 ( .A1(in_47), .A2(in_22), .ZN(n589) );
  AND2_X1 U383bar ( .A1(in_47bar), .A2(in_22bar), .ZN(n589bar);
  OR2_X1 U384 ( .A1(n587), .A2(n586), .ZN(n591) );
  AND2_X1 U384bar ( .A1(n587bar), .A2(n586bar), .ZN(n591bar);
  OR2_X1 U385 ( .A1(in_56), .A2(in_54), .ZN(n586) );
  AND2_X1 U385bar ( .A1(in_56bar), .A2(in_54bar), .ZN(n586bar);
  OR2_X1 U386 ( .A1(in_63), .A2(in_61), .ZN(n587) );
  AND2_X1 U386bar ( .A1(in_63bar), .A2(in_61bar), .ZN(n587bar);
  OR2_X1 U387 ( .A1(n585), .A2(n584), .ZN(n820) );
  AND2_X1 U387bar ( .A1(n585bar), .A2(n584bar), .ZN(n820bar);
  OR2_X1 U388 ( .A1(n583), .A2(n582), .ZN(n584) );
  AND2_X1 U388bar ( .A1(n583bar), .A2(n582bar), .ZN(n584bar);
  OR2_X1 U389 ( .A1(n581), .A2(n580), .ZN(n582) );
  AND2_X1 U389bar ( .A1(n581bar), .A2(n580bar), .ZN(n582bar);
  OR2_X1 U390 ( .A1(in[158]), .A2(in[142]), .ZN(n580) );
  AND2_X1 U390bar ( .A1(inbar[158]), .A2(inbar[142]), .ZN(n580bar);
  OR2_X1 U391 ( .A1(in[175]), .A2(in[164]), .ZN(n581) );
  AND2_X1 U391bar ( .A1(inbar[175]), .A2(inbar[164]), .ZN(n581bar);
  OR2_X1 U392 ( .A1(n579), .A2(n578), .ZN(n583) );
  AND2_X1 U392bar ( .A1(n579bar), .A2(n578bar), .ZN(n583bar);
  OR2_X1 U393 ( .A1(in[228]), .A2(in[204]), .ZN(n578) );
  AND2_X1 U393bar ( .A1(inbar[228]), .A2(inbar[204]), .ZN(n578bar);
  OR2_X1 U394 ( .A1(in[91]), .A2(in[87]), .ZN(n579) );
  AND2_X1 U394bar ( .A1(inbar[91]), .A2(inbar[87]), .ZN(n579bar);
  OR2_X1 U395 ( .A1(n577), .A2(n576), .ZN(n585) );
  AND2_X1 U395bar ( .A1(n577bar), .A2(n576bar), .ZN(n585bar);
  OR2_X1 U396 ( .A1(n575), .A2(n574), .ZN(n576) );
  AND2_X1 U396bar ( .A1(n575bar), .A2(n574bar), .ZN(n576bar);
  OR2_X1 U397 ( .A1(in_21), .A2(in_11), .ZN(n574) );
  AND2_X1 U397bar ( .A1(in_21bar), .A2(in_11bar), .ZN(n574bar);
  OR2_X1 U398 ( .A1(in_5), .A2(in_3), .ZN(n575) );
  AND2_X1 U398bar ( .A1(in_5bar), .A2(in_3bar), .ZN(n575bar);
  OR2_X1 U399 ( .A1(n573), .A2(n572), .ZN(n577) );
  AND2_X1 U399bar ( .A1(n573bar), .A2(n572bar), .ZN(n577bar);
  OR2_X1 U400 ( .A1(in_68), .A2(in_64), .ZN(n572) );
  AND2_X1 U400bar ( .A1(in_68bar), .A2(in_64bar), .ZN(n572bar);
  OR2_X1 U401 ( .A1(in_76), .A2(in_73), .ZN(n573) );
  AND2_X1 U401bar ( .A1(in_76bar), .A2(in_73bar), .ZN(n573bar);
  OR2_X1 U402 ( .A1(n778), .A2(n571), .ZN(n601) );
  AND2_X1 U402bar ( .A1(n778bar), .A2(n571bar), .ZN(n601bar);
  OR2_X1 U403 ( .A1(in[100]), .A2(n965), .ZN(n571) );
  AND2_X1 U403bar ( .A1(inbar[100]), .A2(n965bar), .ZN(n571bar);
  OR2_X1 U404 ( .A1(n570), .A2(n569), .ZN(n965) );
  AND2_X1 U404bar ( .A1(n570bar), .A2(n569bar), .ZN(n965bar);
  OR2_X1 U405 ( .A1(n568), .A2(n567), .ZN(n569) );
  AND2_X1 U405bar ( .A1(n568bar), .A2(n567bar), .ZN(n569bar);
  OR2_X1 U406 ( .A1(n566), .A2(n565), .ZN(n567) );
  AND2_X1 U406bar ( .A1(n566bar), .A2(n565bar), .ZN(n567bar);
  OR2_X1 U407 ( .A1(n817), .A2(n750), .ZN(n565) );
  AND2_X1 U407bar ( .A1(n817bar), .A2(n750bar), .ZN(n565bar);
  OR2_X1 U408 ( .A1(n564), .A2(n563), .ZN(n750) );
  AND2_X1 U408bar ( .A1(n564bar), .A2(n563bar), .ZN(n750bar);
  OR2_X1 U409 ( .A1(n562), .A2(n561), .ZN(n563) );
  AND2_X1 U409bar ( .A1(n562bar), .A2(n561bar), .ZN(n563bar);
  OR2_X1 U410 ( .A1(n560), .A2(n559), .ZN(n561) );
  AND2_X1 U410bar ( .A1(n560bar), .A2(n559bar), .ZN(n561bar);
  OR2_X1 U411 ( .A1(in[119]), .A2(in[103]), .ZN(n559) );
  AND2_X1 U411bar ( .A1(inbar[119]), .A2(inbar[103]), .ZN(n559bar);
  OR2_X1 U412 ( .A1(in[137]), .A2(in[133]), .ZN(n560) );
  AND2_X1 U412bar ( .A1(inbar[137]), .A2(inbar[133]), .ZN(n560bar);
  OR2_X1 U413 ( .A1(n558), .A2(n557), .ZN(n562) );
  AND2_X1 U413bar ( .A1(n558bar), .A2(n557bar), .ZN(n562bar);
  OR2_X1 U414 ( .A1(in[176]), .A2(in[173]), .ZN(n557) );
  AND2_X1 U414bar ( .A1(inbar[176]), .A2(inbar[173]), .ZN(n557bar);
  OR2_X1 U415 ( .A1(in[210]), .A2(in[181]), .ZN(n558) );
  AND2_X1 U415bar ( .A1(inbar[210]), .A2(inbar[181]), .ZN(n558bar);
  OR2_X1 U416 ( .A1(n556), .A2(n555), .ZN(n564) );
  AND2_X1 U416bar ( .A1(n556bar), .A2(n555bar), .ZN(n564bar);
  OR2_X1 U417 ( .A1(n554), .A2(n553), .ZN(n555) );
  AND2_X1 U417bar ( .A1(n554bar), .A2(n553bar), .ZN(n555bar);
  OR2_X1 U418 ( .A1(in_13), .A2(in[234]), .ZN(n553) );
  AND2_X1 U418bar ( .A1(in_13bar), .A2(inbar[234]), .ZN(n553bar);
  OR2_X1 U419 ( .A1(in_38), .A2(in_32), .ZN(n554) );
  AND2_X1 U419bar ( .A1(in_38bar), .A2(in_32bar), .ZN(n554bar);
  OR2_X1 U420 ( .A1(n552), .A2(n551), .ZN(n556) );
  AND2_X1 U420bar ( .A1(n552bar), .A2(n551bar), .ZN(n556bar);
  OR2_X1 U421 ( .A1(in_42), .A2(in_41), .ZN(n551) );
  AND2_X1 U421bar ( .A1(in_42bar), .A2(in_41bar), .ZN(n551bar);
  OR2_X1 U422 ( .A1(in_7), .A2(in_49), .ZN(n552) );
  AND2_X1 U422bar ( .A1(in_7bar), .A2(in_49bar), .ZN(n552bar);
  OR2_X1 U423 ( .A1(n550), .A2(n549), .ZN(n817) );
  AND2_X1 U423bar ( .A1(n550bar), .A2(n549bar), .ZN(n817bar);
  OR2_X1 U424 ( .A1(n548), .A2(n547), .ZN(n549) );
  AND2_X1 U424bar ( .A1(n548bar), .A2(n547bar), .ZN(n549bar);
  OR2_X1 U425 ( .A1(n546), .A2(n545), .ZN(n547) );
  AND2_X1 U425bar ( .A1(n546bar), .A2(n545bar), .ZN(n547bar);
  OR2_X1 U426 ( .A1(in[159]), .A2(in[105]), .ZN(n545) );
  AND2_X1 U426bar ( .A1(inbar[159]), .A2(inbar[105]), .ZN(n545bar);
  OR2_X1 U427 ( .A1(in[206]), .A2(in[183]), .ZN(n546) );
  AND2_X1 U427bar ( .A1(inbar[206]), .A2(inbar[183]), .ZN(n546bar);
  OR2_X1 U428 ( .A1(n544), .A2(n543), .ZN(n548) );
  AND2_X1 U428bar ( .A1(n544bar), .A2(n543bar), .ZN(n548bar);
  OR2_X1 U429 ( .A1(in[229]), .A2(in[219]), .ZN(n543) );
  AND2_X1 U429bar ( .A1(inbar[229]), .A2(inbar[219]), .ZN(n543bar);
  OR2_X1 U430 ( .A1(in[235]), .A2(in[232]), .ZN(n544) );
  AND2_X1 U430bar ( .A1(inbar[235]), .A2(inbar[232]), .ZN(n544bar);
  OR2_X1 U431 ( .A1(n542), .A2(n541), .ZN(n550) );
  AND2_X1 U431bar ( .A1(n542bar), .A2(n541bar), .ZN(n550bar);
  OR2_X1 U432 ( .A1(n540), .A2(n539), .ZN(n541) );
  AND2_X1 U432bar ( .A1(n540bar), .A2(n539bar), .ZN(n541bar);
  OR2_X1 U433 ( .A1(in[249]), .A2(in[242]), .ZN(n539) );
  AND2_X1 U433bar ( .A1(inbar[249]), .A2(inbar[242]), .ZN(n539bar);
  OR2_X1 U434 ( .A1(in[89]), .A2(in[254]), .ZN(n540) );
  AND2_X1 U434bar ( .A1(inbar[89]), .A2(inbar[254]), .ZN(n540bar);
  OR2_X1 U435 ( .A1(n538), .A2(n537), .ZN(n542) );
  AND2_X1 U435bar ( .A1(n538bar), .A2(n537bar), .ZN(n542bar);
  OR2_X1 U436 ( .A1(in_14), .A2(in[99]), .ZN(n537) );
  AND2_X1 U436bar ( .A1(in_14bar), .A2(inbar[99]), .ZN(n537bar);
  OR2_X1 U437 ( .A1(in_60), .A2(in_18), .ZN(n538) );
  AND2_X1 U437bar ( .A1(in_60bar), .A2(in_18bar), .ZN(n538bar);
  OR2_X1 U438 ( .A1(in[113]), .A2(n763), .ZN(n566) );
  AND2_X1 U438bar ( .A1(inbar[113]), .A2(n763bar), .ZN(n566bar);
  OR2_X1 U439 ( .A1(n536), .A2(n535), .ZN(n763) );
  AND2_X1 U439bar ( .A1(n536bar), .A2(n535bar), .ZN(n763bar);
  OR2_X1 U440 ( .A1(n534), .A2(n533), .ZN(n535) );
  AND2_X1 U440bar ( .A1(n534bar), .A2(n533bar), .ZN(n535bar);
  OR2_X1 U441 ( .A1(n532), .A2(n531), .ZN(n533) );
  AND2_X1 U441bar ( .A1(n532bar), .A2(n531bar), .ZN(n533bar);
  OR2_X1 U442 ( .A1(in[115]), .A2(in[110]), .ZN(n531) );
  AND2_X1 U442bar ( .A1(inbar[115]), .A2(inbar[110]), .ZN(n531bar);
  OR2_X1 U443 ( .A1(in[125]), .A2(in[117]), .ZN(n532) );
  AND2_X1 U443bar ( .A1(inbar[125]), .A2(inbar[117]), .ZN(n532bar);
  OR2_X1 U444 ( .A1(n530), .A2(n529), .ZN(n534) );
  AND2_X1 U444bar ( .A1(n530bar), .A2(n529bar), .ZN(n534bar);
  OR2_X1 U445 ( .A1(in[180]), .A2(in[128]), .ZN(n529) );
  AND2_X1 U445bar ( .A1(inbar[180]), .A2(inbar[128]), .ZN(n529bar);
  OR2_X1 U446 ( .A1(in[205]), .A2(in[201]), .ZN(n530) );
  AND2_X1 U446bar ( .A1(inbar[205]), .A2(inbar[201]), .ZN(n530bar);
  OR2_X1 U447 ( .A1(n528), .A2(n527), .ZN(n536) );
  AND2_X1 U447bar ( .A1(n528bar), .A2(n527bar), .ZN(n536bar);
  OR2_X1 U448 ( .A1(n526), .A2(n525), .ZN(n527) );
  AND2_X1 U448bar ( .A1(n526bar), .A2(n525bar), .ZN(n527bar);
  OR2_X1 U449 ( .A1(in[244]), .A2(in[239]), .ZN(n525) );
  AND2_X1 U449bar ( .A1(inbar[244]), .A2(inbar[239]), .ZN(n525bar);
  OR2_X1 U450 ( .A1(in[95]), .A2(in[83]), .ZN(n526) );
  AND2_X1 U450bar ( .A1(inbar[95]), .A2(inbar[83]), .ZN(n526bar);
  OR2_X1 U451 ( .A1(n524), .A2(n523), .ZN(n528) );
  AND2_X1 U451bar ( .A1(n524bar), .A2(n523bar), .ZN(n528bar);
  OR2_X1 U452 ( .A1(in_24), .A2(in[97]), .ZN(n523) );
  AND2_X1 U452bar ( .A1(in_24bar), .A2(inbar[97]), .ZN(n523bar);
  OR2_X1 U453 ( .A1(in_33), .A2(in_27), .ZN(n524) );
  AND2_X1 U453bar ( .A1(in_33bar), .A2(in_27bar), .ZN(n524bar);
  OR2_X1 U454 ( .A1(n522), .A2(n521), .ZN(n568) );
  AND2_X1 U454bar ( .A1(n522bar), .A2(n521bar), .ZN(n568bar);
  OR2_X1 U455 ( .A1(in[145]), .A2(in[126]), .ZN(n521) );
  AND2_X1 U455bar ( .A1(inbar[145]), .A2(inbar[126]), .ZN(n521bar);
  OR2_X1 U456 ( .A1(in[169]), .A2(n520), .ZN(n522) );
  AND2_X1 U456bar ( .A1(inbar[169]), .A2(n520bar), .ZN(n522bar);
  OR2_X1 U457 ( .A1(in[221]), .A2(in[172]), .ZN(n520) );
  AND2_X1 U457bar ( .A1(inbar[221]), .A2(inbar[172]), .ZN(n520bar);
  OR2_X1 U458 ( .A1(n519), .A2(n518), .ZN(n570) );
  AND2_X1 U458bar ( .A1(n519bar), .A2(n518bar), .ZN(n570bar);
  OR2_X1 U459 ( .A1(n517), .A2(n516), .ZN(n518) );
  AND2_X1 U459bar ( .A1(n517bar), .A2(n516bar), .ZN(n518bar);
  OR2_X1 U460 ( .A1(in[241]), .A2(in[224]), .ZN(n516) );
  AND2_X1 U460bar ( .A1(inbar[241]), .A2(inbar[224]), .ZN(n516bar);
  OR2_X1 U461 ( .A1(in[86]), .A2(n515), .ZN(n517) );
  AND2_X1 U461bar ( .A1(inbar[86]), .A2(n515bar), .ZN(n517bar);
  OR2_X1 U462 ( .A1(in_43), .A2(in_34), .ZN(n515) );
  AND2_X1 U462bar ( .A1(in_43bar), .A2(in_34bar), .ZN(n515bar);
  OR2_X1 U463 ( .A1(n514), .A2(n513), .ZN(n519) );
  AND2_X1 U463bar ( .A1(n514bar), .A2(n513bar), .ZN(n519bar);
  OR2_X1 U464 ( .A1(in_65), .A2(in_51), .ZN(n513) );
  AND2_X1 U464bar ( .A1(in_65bar), .A2(in_51bar), .ZN(n513bar);
  OR2_X1 U465 ( .A1(in_75), .A2(n512), .ZN(n514) );
  AND2_X1 U465bar ( .A1(in_75bar), .A2(n512bar), .ZN(n514bar);
  OR2_X1 U466 ( .A1(in_81), .A2(in_77), .ZN(n512) );
  AND2_X1 U466bar ( .A1(in_81bar), .A2(in_77bar), .ZN(n512bar);
  OR2_X1 U467 ( .A1(n511), .A2(n510), .ZN(n778) );
  AND2_X1 U467bar ( .A1(n511bar), .A2(n510bar), .ZN(n778bar);
  OR2_X1 U468 ( .A1(n509), .A2(n508), .ZN(n510) );
  AND2_X1 U468bar ( .A1(n509bar), .A2(n508bar), .ZN(n510bar);
  OR2_X1 U469 ( .A1(n507), .A2(n506), .ZN(n508) );
  AND2_X1 U469bar ( .A1(n507bar), .A2(n506bar), .ZN(n508bar);
  OR2_X1 U470 ( .A1(in[107]), .A2(in[101]), .ZN(n506) );
  AND2_X1 U470bar ( .A1(inbar[107]), .A2(inbar[101]), .ZN(n506bar);
  OR2_X1 U471 ( .A1(in[139]), .A2(in[132]), .ZN(n507) );
  AND2_X1 U471bar ( .A1(inbar[139]), .A2(inbar[132]), .ZN(n507bar);
  OR2_X1 U472 ( .A1(n505), .A2(n504), .ZN(n509) );
  AND2_X1 U472bar ( .A1(n505bar), .A2(n504bar), .ZN(n509bar);
  OR2_X1 U473 ( .A1(in[146]), .A2(in[141]), .ZN(n504) );
  AND2_X1 U473bar ( .A1(inbar[146]), .A2(inbar[141]), .ZN(n504bar);
  OR2_X1 U474 ( .A1(in[203]), .A2(in[179]), .ZN(n505) );
  AND2_X1 U474bar ( .A1(inbar[203]), .A2(inbar[179]), .ZN(n505bar);
  OR2_X1 U475 ( .A1(n503), .A2(n502), .ZN(n511) );
  AND2_X1 U475bar ( .A1(n503bar), .A2(n502bar), .ZN(n511bar);
  OR2_X1 U476 ( .A1(n501), .A2(n500), .ZN(n502) );
  AND2_X1 U476bar ( .A1(n501bar), .A2(n500bar), .ZN(n502bar);
  OR2_X1 U477 ( .A1(in[243]), .A2(in[222]), .ZN(n500) );
  AND2_X1 U477bar ( .A1(inbar[243]), .A2(inbar[222]), .ZN(n500bar);
  OR2_X1 U478 ( .A1(in[251]), .A2(in[250]), .ZN(n501) );
  AND2_X1 U478bar ( .A1(inbar[251]), .A2(inbar[250]), .ZN(n501bar);
  OR2_X1 U479 ( .A1(n499), .A2(n498), .ZN(n503) );
  AND2_X1 U479bar ( .A1(n499bar), .A2(n498bar), .ZN(n503bar);
  OR2_X1 U480 ( .A1(in_37), .A2(in_19), .ZN(n498) );
  AND2_X1 U480bar ( .A1(in_37bar), .A2(in_19bar), .ZN(n498bar);
  OR2_X1 U481 ( .A1(in_78), .A2(in_6), .ZN(n499) );
  AND2_X1 U481bar ( .A1(in_78bar), .A2(in_6bar), .ZN(n499bar);
  OR2_X1 U482 ( .A1(n497), .A2(n496), .ZN(n603) );
  AND2_X1 U482bar ( .A1(n497bar), .A2(n496bar), .ZN(n603bar);
  OR2_X1 U483 ( .A1(in[112]), .A2(in[102]), .ZN(n496) );
  AND2_X1 U483bar ( .A1(inbar[112]), .A2(inbar[102]), .ZN(n496bar);
  OR2_X1 U484 ( .A1(in[123]), .A2(n495), .ZN(n497) );
  AND2_X1 U484bar ( .A1(inbar[123]), .A2(n495bar), .ZN(n497bar);
  OR2_X1 U485 ( .A1(in[143]), .A2(in[130]), .ZN(n495) );
  AND2_X1 U485bar ( .A1(inbar[143]), .A2(inbar[130]), .ZN(n495bar);
  OR2_X1 U486 ( .A1(n494), .A2(n493), .ZN(n605) );
  AND2_X1 U486bar ( .A1(n494bar), .A2(n493bar), .ZN(n605bar);
  OR2_X1 U487 ( .A1(n492), .A2(n491), .ZN(n493) );
  AND2_X1 U487bar ( .A1(n492bar), .A2(n491bar), .ZN(n493bar);
  OR2_X1 U488 ( .A1(in[216]), .A2(in[213]), .ZN(n491) );
  AND2_X1 U488bar ( .A1(inbar[216]), .A2(inbar[213]), .ZN(n491bar);
  OR2_X1 U489 ( .A1(in[227]), .A2(n490), .ZN(n492) );
  AND2_X1 U489bar ( .A1(inbar[227]), .A2(n490bar), .ZN(n492bar);
  OR2_X1 U490 ( .A1(in_0), .A2(in[248]), .ZN(n490) );
  AND2_X1 U490bar ( .A1(in_0bar), .A2(inbar[248]), .ZN(n490bar);
  OR2_X1 U491 ( .A1(n489), .A2(n488), .ZN(n494) );
  AND2_X1 U491bar ( .A1(n489bar), .A2(n488bar), .ZN(n494bar);
  OR2_X1 U492 ( .A1(in_46), .A2(in_44), .ZN(n488) );
  AND2_X1 U492bar ( .A1(in_46bar), .A2(in_44bar), .ZN(n488bar);
  OR2_X1 U493 ( .A1(in_50), .A2(n487), .ZN(n489) );
  AND2_X1 U493bar ( .A1(in_50bar), .A2(n487bar), .ZN(n489bar);
  OR2_X1 U494 ( .A1(in_9), .A2(in_80), .ZN(n487) );
  AND2_X1 U494bar ( .A1(in_9bar), .A2(in_80bar), .ZN(n487bar);
endmodule




module sBox_11 ( in, out );
  input [7:0] in;
  //input_done

  output [7:0] out;
  //output_done

  wire   [255:0] decodeOut;
  //wire_done

  decode_11 dec ( .in(in), .out(decodeOut) );
  encode_11 enc ( .in(decodeOut), .out(out) );
endmodule


module CD2_45 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_46 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_47 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_48 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD4_23 ( a, b, y );
  input [3:0] a;
  input [3:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  //input_done

  output [15:0] y;
  reg [15:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]);
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]);
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]);
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]);
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]);
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]);
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]);
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]);
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]);
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]);
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]);
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]);
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]);
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]);
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]);
endmodule




module CD4_24 ( a, b, y );
  input [3:0] a;
  input [3:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  //input_done

  output [15:0] y;
  reg [15:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]);
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]);
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]);
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]);
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]);
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]);
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]);
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]);
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]);
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]);
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]);
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]);
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]);
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]);
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]);
endmodule




module CD16_12 ( a, b, y );
  input [15:0] a;
  input [15:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign abar[8] = ~a[8];
  assign abar[9] = ~a[9];
  assign abar[10] = ~a[10];
  assign abar[11] = ~a[11];
  assign abar[12] = ~a[12];
  assign abar[13] = ~a[13];
  assign abar[14] = ~a[14];
  assign abar[15] = ~a[15];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign bbar[8] = ~b[8];
  assign bbar[9] = ~b[9];
  assign bbar[10] = ~b[10];
  assign bbar[11] = ~b[11];
  assign bbar[12] = ~b[12];
  assign bbar[13] = ~b[13];
  assign bbar[14] = ~b[14];
  assign bbar[15] = ~b[15];
  //input_done

  output [255:0] y;
  reg [255:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[9]), .A2(a[0]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[9]), .A2(abar[0]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[3]), .A2(a[6]), .ZN(y[99]) );
  OR2_X1 U2bar ( .A1(bbar[3]), .A2(abar[6]), .ZN(ybar[99]);
  AND2_X1 U3 ( .A1(b[2]), .A2(a[6]), .ZN(y[98]) );
  OR2_X1 U3bar ( .A1(bbar[2]), .A2(abar[6]), .ZN(ybar[98]);
  AND2_X1 U4 ( .A1(b[1]), .A2(a[6]), .ZN(y[97]) );
  OR2_X1 U4bar ( .A1(bbar[1]), .A2(abar[6]), .ZN(ybar[97]);
  AND2_X1 U5 ( .A1(b[0]), .A2(a[6]), .ZN(y[96]) );
  OR2_X1 U5bar ( .A1(bbar[0]), .A2(abar[6]), .ZN(ybar[96]);
  AND2_X1 U6 ( .A1(b[15]), .A2(a[5]), .ZN(y[95]) );
  OR2_X1 U6bar ( .A1(bbar[15]), .A2(abar[5]), .ZN(ybar[95]);
  AND2_X1 U7 ( .A1(b[14]), .A2(a[5]), .ZN(y[94]) );
  OR2_X1 U7bar ( .A1(bbar[14]), .A2(abar[5]), .ZN(ybar[94]);
  AND2_X1 U8 ( .A1(b[13]), .A2(a[5]), .ZN(y[93]) );
  OR2_X1 U8bar ( .A1(bbar[13]), .A2(abar[5]), .ZN(ybar[93]);
  AND2_X1 U9 ( .A1(b[12]), .A2(a[5]), .ZN(y[92]) );
  OR2_X1 U9bar ( .A1(bbar[12]), .A2(abar[5]), .ZN(ybar[92]);
  AND2_X1 U10 ( .A1(b[11]), .A2(a[5]), .ZN(y[91]) );
  OR2_X1 U10bar ( .A1(bbar[11]), .A2(abar[5]), .ZN(ybar[91]);
  AND2_X1 U11 ( .A1(b[10]), .A2(a[5]), .ZN(y[90]) );
  OR2_X1 U11bar ( .A1(bbar[10]), .A2(abar[5]), .ZN(ybar[90]);
  AND2_X1 U12 ( .A1(b[8]), .A2(a[0]), .ZN(y[8]) );
  OR2_X1 U12bar ( .A1(bbar[8]), .A2(abar[0]), .ZN(ybar[8]);
  AND2_X1 U13 ( .A1(a[5]), .A2(b[9]), .ZN(y[89]) );
  OR2_X1 U13bar ( .A1(abar[5]), .A2(bbar[9]), .ZN(ybar[89]);
  AND2_X1 U14 ( .A1(b[8]), .A2(a[5]), .ZN(y[88]) );
  OR2_X1 U14bar ( .A1(bbar[8]), .A2(abar[5]), .ZN(ybar[88]);
  AND2_X1 U15 ( .A1(b[7]), .A2(a[5]), .ZN(y[87]) );
  OR2_X1 U15bar ( .A1(bbar[7]), .A2(abar[5]), .ZN(ybar[87]);
  AND2_X1 U16 ( .A1(b[6]), .A2(a[5]), .ZN(y[86]) );
  OR2_X1 U16bar ( .A1(bbar[6]), .A2(abar[5]), .ZN(ybar[86]);
  AND2_X1 U17 ( .A1(b[5]), .A2(a[5]), .ZN(y[85]) );
  OR2_X1 U17bar ( .A1(bbar[5]), .A2(abar[5]), .ZN(ybar[85]);
  AND2_X1 U18 ( .A1(b[4]), .A2(a[5]), .ZN(y[84]) );
  OR2_X1 U18bar ( .A1(bbar[4]), .A2(abar[5]), .ZN(ybar[84]);
  AND2_X1 U19 ( .A1(a[5]), .A2(b[3]), .ZN(y[83]) );
  OR2_X1 U19bar ( .A1(abar[5]), .A2(bbar[3]), .ZN(ybar[83]);
  AND2_X1 U20 ( .A1(a[5]), .A2(b[2]), .ZN(y[82]) );
  OR2_X1 U20bar ( .A1(abar[5]), .A2(bbar[2]), .ZN(ybar[82]);
  AND2_X1 U21 ( .A1(a[5]), .A2(b[1]), .ZN(y[81]) );
  OR2_X1 U21bar ( .A1(abar[5]), .A2(bbar[1]), .ZN(ybar[81]);
  AND2_X1 U22 ( .A1(a[5]), .A2(b[0]), .ZN(y[80]) );
  OR2_X1 U22bar ( .A1(abar[5]), .A2(bbar[0]), .ZN(ybar[80]);
  AND2_X1 U23 ( .A1(b[7]), .A2(a[0]), .ZN(y[7]) );
  OR2_X1 U23bar ( .A1(bbar[7]), .A2(abar[0]), .ZN(ybar[7]);
  AND2_X1 U24 ( .A1(a[4]), .A2(b[15]), .ZN(y[79]) );
  OR2_X1 U24bar ( .A1(abar[4]), .A2(bbar[15]), .ZN(ybar[79]);
  AND2_X1 U25 ( .A1(a[4]), .A2(b[14]), .ZN(y[78]) );
  OR2_X1 U25bar ( .A1(abar[4]), .A2(bbar[14]), .ZN(ybar[78]);
  AND2_X1 U26 ( .A1(a[4]), .A2(b[13]), .ZN(y[77]) );
  OR2_X1 U26bar ( .A1(abar[4]), .A2(bbar[13]), .ZN(ybar[77]);
  AND2_X1 U27 ( .A1(a[4]), .A2(b[12]), .ZN(y[76]) );
  OR2_X1 U27bar ( .A1(abar[4]), .A2(bbar[12]), .ZN(ybar[76]);
  AND2_X1 U28 ( .A1(a[4]), .A2(b[11]), .ZN(y[75]) );
  OR2_X1 U28bar ( .A1(abar[4]), .A2(bbar[11]), .ZN(ybar[75]);
  AND2_X1 U29 ( .A1(a[4]), .A2(b[10]), .ZN(y[74]) );
  OR2_X1 U29bar ( .A1(abar[4]), .A2(bbar[10]), .ZN(ybar[74]);
  AND2_X1 U30 ( .A1(a[4]), .A2(b[9]), .ZN(y[73]) );
  OR2_X1 U30bar ( .A1(abar[4]), .A2(bbar[9]), .ZN(ybar[73]);
  AND2_X1 U31 ( .A1(a[4]), .A2(b[8]), .ZN(y[72]) );
  OR2_X1 U31bar ( .A1(abar[4]), .A2(bbar[8]), .ZN(ybar[72]);
  AND2_X1 U32 ( .A1(a[4]), .A2(b[7]), .ZN(y[71]) );
  OR2_X1 U32bar ( .A1(abar[4]), .A2(bbar[7]), .ZN(ybar[71]);
  AND2_X1 U33 ( .A1(a[4]), .A2(b[6]), .ZN(y[70]) );
  OR2_X1 U33bar ( .A1(abar[4]), .A2(bbar[6]), .ZN(ybar[70]);
  AND2_X1 U34 ( .A1(b[6]), .A2(a[0]), .ZN(y[6]) );
  OR2_X1 U34bar ( .A1(bbar[6]), .A2(abar[0]), .ZN(ybar[6]);
  AND2_X1 U35 ( .A1(a[4]), .A2(b[5]), .ZN(y[69]) );
  OR2_X1 U35bar ( .A1(abar[4]), .A2(bbar[5]), .ZN(ybar[69]);
  AND2_X1 U36 ( .A1(a[4]), .A2(b[4]), .ZN(y[68]) );
  OR2_X1 U36bar ( .A1(abar[4]), .A2(bbar[4]), .ZN(ybar[68]);
  AND2_X1 U37 ( .A1(a[4]), .A2(b[3]), .ZN(y[67]) );
  OR2_X1 U37bar ( .A1(abar[4]), .A2(bbar[3]), .ZN(ybar[67]);
  AND2_X1 U38 ( .A1(a[4]), .A2(b[2]), .ZN(y[66]) );
  OR2_X1 U38bar ( .A1(abar[4]), .A2(bbar[2]), .ZN(ybar[66]);
  AND2_X1 U39 ( .A1(a[4]), .A2(b[1]), .ZN(y[65]) );
  OR2_X1 U39bar ( .A1(abar[4]), .A2(bbar[1]), .ZN(ybar[65]);
  AND2_X1 U40 ( .A1(a[4]), .A2(b[0]), .ZN(y[64]) );
  OR2_X1 U40bar ( .A1(abar[4]), .A2(bbar[0]), .ZN(ybar[64]);
  AND2_X1 U41 ( .A1(a[3]), .A2(b[15]), .ZN(y[63]) );
  OR2_X1 U41bar ( .A1(abar[3]), .A2(bbar[15]), .ZN(ybar[63]);
  AND2_X1 U42 ( .A1(a[3]), .A2(b[14]), .ZN(y[62]) );
  OR2_X1 U42bar ( .A1(abar[3]), .A2(bbar[14]), .ZN(ybar[62]);
  AND2_X1 U43 ( .A1(a[3]), .A2(b[13]), .ZN(y[61]) );
  OR2_X1 U43bar ( .A1(abar[3]), .A2(bbar[13]), .ZN(ybar[61]);
  AND2_X1 U44 ( .A1(a[3]), .A2(b[12]), .ZN(y[60]) );
  OR2_X1 U44bar ( .A1(abar[3]), .A2(bbar[12]), .ZN(ybar[60]);
  AND2_X1 U45 ( .A1(b[5]), .A2(a[0]), .ZN(y[5]) );
  OR2_X1 U45bar ( .A1(bbar[5]), .A2(abar[0]), .ZN(ybar[5]);
  AND2_X1 U46 ( .A1(a[3]), .A2(b[11]), .ZN(y[59]) );
  OR2_X1 U46bar ( .A1(abar[3]), .A2(bbar[11]), .ZN(ybar[59]);
  AND2_X1 U47 ( .A1(a[3]), .A2(b[10]), .ZN(y[58]) );
  OR2_X1 U47bar ( .A1(abar[3]), .A2(bbar[10]), .ZN(ybar[58]);
  AND2_X1 U48 ( .A1(a[3]), .A2(b[9]), .ZN(y[57]) );
  OR2_X1 U48bar ( .A1(abar[3]), .A2(bbar[9]), .ZN(ybar[57]);
  AND2_X1 U49 ( .A1(a[3]), .A2(b[8]), .ZN(y[56]) );
  OR2_X1 U49bar ( .A1(abar[3]), .A2(bbar[8]), .ZN(ybar[56]);
  AND2_X1 U50 ( .A1(a[3]), .A2(b[7]), .ZN(y[55]) );
  OR2_X1 U50bar ( .A1(abar[3]), .A2(bbar[7]), .ZN(ybar[55]);
  AND2_X1 U51 ( .A1(a[3]), .A2(b[6]), .ZN(y[54]) );
  OR2_X1 U51bar ( .A1(abar[3]), .A2(bbar[6]), .ZN(ybar[54]);
  AND2_X1 U52 ( .A1(a[3]), .A2(b[5]), .ZN(y[53]) );
  OR2_X1 U52bar ( .A1(abar[3]), .A2(bbar[5]), .ZN(ybar[53]);
  AND2_X1 U53 ( .A1(a[3]), .A2(b[4]), .ZN(y[52]) );
  OR2_X1 U53bar ( .A1(abar[3]), .A2(bbar[4]), .ZN(ybar[52]);
  AND2_X1 U54 ( .A1(a[3]), .A2(b[3]), .ZN(y[51]) );
  OR2_X1 U54bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[51]);
  AND2_X1 U55 ( .A1(a[3]), .A2(b[2]), .ZN(y[50]) );
  OR2_X1 U55bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[50]);
  AND2_X1 U56 ( .A1(b[4]), .A2(a[0]), .ZN(y[4]) );
  OR2_X1 U56bar ( .A1(bbar[4]), .A2(abar[0]), .ZN(ybar[4]);
  AND2_X1 U57 ( .A1(a[3]), .A2(b[1]), .ZN(y[49]) );
  OR2_X1 U57bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[49]);
  AND2_X1 U58 ( .A1(a[3]), .A2(b[0]), .ZN(y[48]) );
  OR2_X1 U58bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[48]);
  AND2_X1 U59 ( .A1(a[2]), .A2(b[15]), .ZN(y[47]) );
  OR2_X1 U59bar ( .A1(abar[2]), .A2(bbar[15]), .ZN(ybar[47]);
  AND2_X1 U60 ( .A1(a[2]), .A2(b[14]), .ZN(y[46]) );
  OR2_X1 U60bar ( .A1(abar[2]), .A2(bbar[14]), .ZN(ybar[46]);
  AND2_X1 U61 ( .A1(a[2]), .A2(b[13]), .ZN(y[45]) );
  OR2_X1 U61bar ( .A1(abar[2]), .A2(bbar[13]), .ZN(ybar[45]);
  AND2_X1 U62 ( .A1(a[2]), .A2(b[12]), .ZN(y[44]) );
  OR2_X1 U62bar ( .A1(abar[2]), .A2(bbar[12]), .ZN(ybar[44]);
  AND2_X1 U63 ( .A1(a[2]), .A2(b[11]), .ZN(y[43]) );
  OR2_X1 U63bar ( .A1(abar[2]), .A2(bbar[11]), .ZN(ybar[43]);
  AND2_X1 U64 ( .A1(a[2]), .A2(b[10]), .ZN(y[42]) );
  OR2_X1 U64bar ( .A1(abar[2]), .A2(bbar[10]), .ZN(ybar[42]);
  AND2_X1 U65 ( .A1(a[2]), .A2(b[9]), .ZN(y[41]) );
  OR2_X1 U65bar ( .A1(abar[2]), .A2(bbar[9]), .ZN(ybar[41]);
  AND2_X1 U66 ( .A1(a[2]), .A2(b[8]), .ZN(y[40]) );
  OR2_X1 U66bar ( .A1(abar[2]), .A2(bbar[8]), .ZN(ybar[40]);
  AND2_X1 U67 ( .A1(b[3]), .A2(a[0]), .ZN(y[3]) );
  OR2_X1 U67bar ( .A1(bbar[3]), .A2(abar[0]), .ZN(ybar[3]);
  AND2_X1 U68 ( .A1(a[2]), .A2(b[7]), .ZN(y[39]) );
  OR2_X1 U68bar ( .A1(abar[2]), .A2(bbar[7]), .ZN(ybar[39]);
  AND2_X1 U69 ( .A1(a[2]), .A2(b[6]), .ZN(y[38]) );
  OR2_X1 U69bar ( .A1(abar[2]), .A2(bbar[6]), .ZN(ybar[38]);
  AND2_X1 U70 ( .A1(a[2]), .A2(b[5]), .ZN(y[37]) );
  OR2_X1 U70bar ( .A1(abar[2]), .A2(bbar[5]), .ZN(ybar[37]);
  AND2_X1 U71 ( .A1(a[2]), .A2(b[4]), .ZN(y[36]) );
  OR2_X1 U71bar ( .A1(abar[2]), .A2(bbar[4]), .ZN(ybar[36]);
  AND2_X1 U72 ( .A1(a[2]), .A2(b[3]), .ZN(y[35]) );
  OR2_X1 U72bar ( .A1(abar[2]), .A2(bbar[3]), .ZN(ybar[35]);
  AND2_X1 U73 ( .A1(a[2]), .A2(b[2]), .ZN(y[34]) );
  OR2_X1 U73bar ( .A1(abar[2]), .A2(bbar[2]), .ZN(ybar[34]);
  AND2_X1 U74 ( .A1(a[2]), .A2(b[1]), .ZN(y[33]) );
  OR2_X1 U74bar ( .A1(abar[2]), .A2(bbar[1]), .ZN(ybar[33]);
  AND2_X1 U75 ( .A1(a[2]), .A2(b[0]), .ZN(y[32]) );
  OR2_X1 U75bar ( .A1(abar[2]), .A2(bbar[0]), .ZN(ybar[32]);
  AND2_X1 U76 ( .A1(a[1]), .A2(b[15]), .ZN(y[31]) );
  OR2_X1 U76bar ( .A1(abar[1]), .A2(bbar[15]), .ZN(ybar[31]);
  AND2_X1 U77 ( .A1(a[1]), .A2(b[14]), .ZN(y[30]) );
  OR2_X1 U77bar ( .A1(abar[1]), .A2(bbar[14]), .ZN(ybar[30]);
  AND2_X1 U78 ( .A1(b[2]), .A2(a[0]), .ZN(y[2]) );
  OR2_X1 U78bar ( .A1(bbar[2]), .A2(abar[0]), .ZN(ybar[2]);
  AND2_X1 U79 ( .A1(a[1]), .A2(b[13]), .ZN(y[29]) );
  OR2_X1 U79bar ( .A1(abar[1]), .A2(bbar[13]), .ZN(ybar[29]);
  AND2_X1 U80 ( .A1(a[1]), .A2(b[12]), .ZN(y[28]) );
  OR2_X1 U80bar ( .A1(abar[1]), .A2(bbar[12]), .ZN(ybar[28]);
  AND2_X1 U81 ( .A1(a[1]), .A2(b[11]), .ZN(y[27]) );
  OR2_X1 U81bar ( .A1(abar[1]), .A2(bbar[11]), .ZN(ybar[27]);
  AND2_X1 U82 ( .A1(a[1]), .A2(b[10]), .ZN(y[26]) );
  OR2_X1 U82bar ( .A1(abar[1]), .A2(bbar[10]), .ZN(ybar[26]);
  AND2_X1 U83 ( .A1(a[1]), .A2(b[9]), .ZN(y[25]) );
  OR2_X1 U83bar ( .A1(abar[1]), .A2(bbar[9]), .ZN(ybar[25]);
  AND2_X1 U84 ( .A1(a[15]), .A2(b[15]), .ZN(y[255]) );
  OR2_X1 U84bar ( .A1(abar[15]), .A2(bbar[15]), .ZN(ybar[255]);
  AND2_X1 U85 ( .A1(a[15]), .A2(b[14]), .ZN(y[254]) );
  OR2_X1 U85bar ( .A1(abar[15]), .A2(bbar[14]), .ZN(ybar[254]);
  AND2_X1 U86 ( .A1(a[15]), .A2(b[13]), .ZN(y[253]) );
  OR2_X1 U86bar ( .A1(abar[15]), .A2(bbar[13]), .ZN(ybar[253]);
  AND2_X1 U87 ( .A1(a[15]), .A2(b[12]), .ZN(y[252]) );
  OR2_X1 U87bar ( .A1(abar[15]), .A2(bbar[12]), .ZN(ybar[252]);
  AND2_X1 U88 ( .A1(a[15]), .A2(b[11]), .ZN(y[251]) );
  OR2_X1 U88bar ( .A1(abar[15]), .A2(bbar[11]), .ZN(ybar[251]);
  AND2_X1 U89 ( .A1(a[15]), .A2(b[10]), .ZN(y[250]) );
  OR2_X1 U89bar ( .A1(abar[15]), .A2(bbar[10]), .ZN(ybar[250]);
  AND2_X1 U90 ( .A1(a[1]), .A2(b[8]), .ZN(y[24]) );
  OR2_X1 U90bar ( .A1(abar[1]), .A2(bbar[8]), .ZN(ybar[24]);
  AND2_X1 U91 ( .A1(a[15]), .A2(b[9]), .ZN(y[249]) );
  OR2_X1 U91bar ( .A1(abar[15]), .A2(bbar[9]), .ZN(ybar[249]);
  AND2_X1 U92 ( .A1(a[15]), .A2(b[8]), .ZN(y[248]) );
  OR2_X1 U92bar ( .A1(abar[15]), .A2(bbar[8]), .ZN(ybar[248]);
  AND2_X1 U93 ( .A1(a[15]), .A2(b[7]), .ZN(y[247]) );
  OR2_X1 U93bar ( .A1(abar[15]), .A2(bbar[7]), .ZN(ybar[247]);
  AND2_X1 U94 ( .A1(a[15]), .A2(b[6]), .ZN(y[246]) );
  OR2_X1 U94bar ( .A1(abar[15]), .A2(bbar[6]), .ZN(ybar[246]);
  AND2_X1 U95 ( .A1(a[15]), .A2(b[5]), .ZN(y[245]) );
  OR2_X1 U95bar ( .A1(abar[15]), .A2(bbar[5]), .ZN(ybar[245]);
  AND2_X1 U96 ( .A1(a[15]), .A2(b[4]), .ZN(y[244]) );
  OR2_X1 U96bar ( .A1(abar[15]), .A2(bbar[4]), .ZN(ybar[244]);
  AND2_X1 U97 ( .A1(a[15]), .A2(b[3]), .ZN(y[243]) );
  OR2_X1 U97bar ( .A1(abar[15]), .A2(bbar[3]), .ZN(ybar[243]);
  AND2_X1 U98 ( .A1(a[15]), .A2(b[2]), .ZN(y[242]) );
  OR2_X1 U98bar ( .A1(abar[15]), .A2(bbar[2]), .ZN(ybar[242]);
  AND2_X1 U99 ( .A1(a[15]), .A2(b[1]), .ZN(y[241]) );
  OR2_X1 U99bar ( .A1(abar[15]), .A2(bbar[1]), .ZN(ybar[241]);
  AND2_X1 U100 ( .A1(a[15]), .A2(b[0]), .ZN(y[240]) );
  OR2_X1 U100bar ( .A1(abar[15]), .A2(bbar[0]), .ZN(ybar[240]);
  AND2_X1 U101 ( .A1(a[1]), .A2(b[7]), .ZN(y[23]) );
  OR2_X1 U101bar ( .A1(abar[1]), .A2(bbar[7]), .ZN(ybar[23]);
  AND2_X1 U102 ( .A1(a[14]), .A2(b[15]), .ZN(y[239]) );
  OR2_X1 U102bar ( .A1(abar[14]), .A2(bbar[15]), .ZN(ybar[239]);
  AND2_X1 U103 ( .A1(a[14]), .A2(b[14]), .ZN(y[238]) );
  OR2_X1 U103bar ( .A1(abar[14]), .A2(bbar[14]), .ZN(ybar[238]);
  AND2_X1 U104 ( .A1(a[14]), .A2(b[13]), .ZN(y[237]) );
  OR2_X1 U104bar ( .A1(abar[14]), .A2(bbar[13]), .ZN(ybar[237]);
  AND2_X1 U105 ( .A1(a[14]), .A2(b[12]), .ZN(y[236]) );
  OR2_X1 U105bar ( .A1(abar[14]), .A2(bbar[12]), .ZN(ybar[236]);
  AND2_X1 U106 ( .A1(a[14]), .A2(b[11]), .ZN(y[235]) );
  OR2_X1 U106bar ( .A1(abar[14]), .A2(bbar[11]), .ZN(ybar[235]);
  AND2_X1 U107 ( .A1(a[14]), .A2(b[10]), .ZN(y[234]) );
  OR2_X1 U107bar ( .A1(abar[14]), .A2(bbar[10]), .ZN(ybar[234]);
  AND2_X1 U108 ( .A1(a[14]), .A2(b[9]), .ZN(y[233]) );
  OR2_X1 U108bar ( .A1(abar[14]), .A2(bbar[9]), .ZN(ybar[233]);
  AND2_X1 U109 ( .A1(a[14]), .A2(b[8]), .ZN(y[232]) );
  OR2_X1 U109bar ( .A1(abar[14]), .A2(bbar[8]), .ZN(ybar[232]);
  AND2_X1 U110 ( .A1(a[14]), .A2(b[7]), .ZN(y[231]) );
  OR2_X1 U110bar ( .A1(abar[14]), .A2(bbar[7]), .ZN(ybar[231]);
  AND2_X1 U111 ( .A1(a[14]), .A2(b[6]), .ZN(y[230]) );
  OR2_X1 U111bar ( .A1(abar[14]), .A2(bbar[6]), .ZN(ybar[230]);
  AND2_X1 U112 ( .A1(a[1]), .A2(b[6]), .ZN(y[22]) );
  OR2_X1 U112bar ( .A1(abar[1]), .A2(bbar[6]), .ZN(ybar[22]);
  AND2_X1 U113 ( .A1(a[14]), .A2(b[5]), .ZN(y[229]) );
  OR2_X1 U113bar ( .A1(abar[14]), .A2(bbar[5]), .ZN(ybar[229]);
  AND2_X1 U114 ( .A1(a[14]), .A2(b[4]), .ZN(y[228]) );
  OR2_X1 U114bar ( .A1(abar[14]), .A2(bbar[4]), .ZN(ybar[228]);
  AND2_X1 U115 ( .A1(a[14]), .A2(b[3]), .ZN(y[227]) );
  OR2_X1 U115bar ( .A1(abar[14]), .A2(bbar[3]), .ZN(ybar[227]);
  AND2_X1 U116 ( .A1(a[14]), .A2(b[2]), .ZN(y[226]) );
  OR2_X1 U116bar ( .A1(abar[14]), .A2(bbar[2]), .ZN(ybar[226]);
  AND2_X1 U117 ( .A1(a[14]), .A2(b[1]), .ZN(y[225]) );
  OR2_X1 U117bar ( .A1(abar[14]), .A2(bbar[1]), .ZN(ybar[225]);
  AND2_X1 U118 ( .A1(a[14]), .A2(b[0]), .ZN(y[224]) );
  OR2_X1 U118bar ( .A1(abar[14]), .A2(bbar[0]), .ZN(ybar[224]);
  AND2_X1 U119 ( .A1(a[13]), .A2(b[15]), .ZN(y[223]) );
  OR2_X1 U119bar ( .A1(abar[13]), .A2(bbar[15]), .ZN(ybar[223]);
  AND2_X1 U120 ( .A1(a[13]), .A2(b[14]), .ZN(y[222]) );
  OR2_X1 U120bar ( .A1(abar[13]), .A2(bbar[14]), .ZN(ybar[222]);
  AND2_X1 U121 ( .A1(a[13]), .A2(b[13]), .ZN(y[221]) );
  OR2_X1 U121bar ( .A1(abar[13]), .A2(bbar[13]), .ZN(ybar[221]);
  AND2_X1 U122 ( .A1(a[13]), .A2(b[12]), .ZN(y[220]) );
  OR2_X1 U122bar ( .A1(abar[13]), .A2(bbar[12]), .ZN(ybar[220]);
  AND2_X1 U123 ( .A1(a[1]), .A2(b[5]), .ZN(y[21]) );
  OR2_X1 U123bar ( .A1(abar[1]), .A2(bbar[5]), .ZN(ybar[21]);
  AND2_X1 U124 ( .A1(a[13]), .A2(b[11]), .ZN(y[219]) );
  OR2_X1 U124bar ( .A1(abar[13]), .A2(bbar[11]), .ZN(ybar[219]);
  AND2_X1 U125 ( .A1(a[13]), .A2(b[10]), .ZN(y[218]) );
  OR2_X1 U125bar ( .A1(abar[13]), .A2(bbar[10]), .ZN(ybar[218]);
  AND2_X1 U126 ( .A1(a[13]), .A2(b[9]), .ZN(y[217]) );
  OR2_X1 U126bar ( .A1(abar[13]), .A2(bbar[9]), .ZN(ybar[217]);
  AND2_X1 U127 ( .A1(a[13]), .A2(b[8]), .ZN(y[216]) );
  OR2_X1 U127bar ( .A1(abar[13]), .A2(bbar[8]), .ZN(ybar[216]);
  AND2_X1 U128 ( .A1(a[13]), .A2(b[7]), .ZN(y[215]) );
  OR2_X1 U128bar ( .A1(abar[13]), .A2(bbar[7]), .ZN(ybar[215]);
  AND2_X1 U129 ( .A1(a[13]), .A2(b[6]), .ZN(y[214]) );
  OR2_X1 U129bar ( .A1(abar[13]), .A2(bbar[6]), .ZN(ybar[214]);
  AND2_X1 U130 ( .A1(a[13]), .A2(b[5]), .ZN(y[213]) );
  OR2_X1 U130bar ( .A1(abar[13]), .A2(bbar[5]), .ZN(ybar[213]);
  AND2_X1 U131 ( .A1(a[13]), .A2(b[4]), .ZN(y[212]) );
  OR2_X1 U131bar ( .A1(abar[13]), .A2(bbar[4]), .ZN(ybar[212]);
  AND2_X1 U132 ( .A1(a[13]), .A2(b[3]), .ZN(y[211]) );
  OR2_X1 U132bar ( .A1(abar[13]), .A2(bbar[3]), .ZN(ybar[211]);
  AND2_X1 U133 ( .A1(a[13]), .A2(b[2]), .ZN(y[210]) );
  OR2_X1 U133bar ( .A1(abar[13]), .A2(bbar[2]), .ZN(ybar[210]);
  AND2_X1 U134 ( .A1(a[1]), .A2(b[4]), .ZN(y[20]) );
  OR2_X1 U134bar ( .A1(abar[1]), .A2(bbar[4]), .ZN(ybar[20]);
  AND2_X1 U135 ( .A1(a[13]), .A2(b[1]), .ZN(y[209]) );
  OR2_X1 U135bar ( .A1(abar[13]), .A2(bbar[1]), .ZN(ybar[209]);
  AND2_X1 U136 ( .A1(a[13]), .A2(b[0]), .ZN(y[208]) );
  OR2_X1 U136bar ( .A1(abar[13]), .A2(bbar[0]), .ZN(ybar[208]);
  AND2_X1 U137 ( .A1(a[12]), .A2(b[15]), .ZN(y[207]) );
  OR2_X1 U137bar ( .A1(abar[12]), .A2(bbar[15]), .ZN(ybar[207]);
  AND2_X1 U138 ( .A1(a[12]), .A2(b[14]), .ZN(y[206]) );
  OR2_X1 U138bar ( .A1(abar[12]), .A2(bbar[14]), .ZN(ybar[206]);
  AND2_X1 U139 ( .A1(a[12]), .A2(b[13]), .ZN(y[205]) );
  OR2_X1 U139bar ( .A1(abar[12]), .A2(bbar[13]), .ZN(ybar[205]);
  AND2_X1 U140 ( .A1(a[12]), .A2(b[12]), .ZN(y[204]) );
  OR2_X1 U140bar ( .A1(abar[12]), .A2(bbar[12]), .ZN(ybar[204]);
  AND2_X1 U141 ( .A1(a[12]), .A2(b[11]), .ZN(y[203]) );
  OR2_X1 U141bar ( .A1(abar[12]), .A2(bbar[11]), .ZN(ybar[203]);
  AND2_X1 U142 ( .A1(a[12]), .A2(b[10]), .ZN(y[202]) );
  OR2_X1 U142bar ( .A1(abar[12]), .A2(bbar[10]), .ZN(ybar[202]);
  AND2_X1 U143 ( .A1(a[12]), .A2(b[9]), .ZN(y[201]) );
  OR2_X1 U143bar ( .A1(abar[12]), .A2(bbar[9]), .ZN(ybar[201]);
  AND2_X1 U144 ( .A1(a[12]), .A2(b[8]), .ZN(y[200]) );
  OR2_X1 U144bar ( .A1(abar[12]), .A2(bbar[8]), .ZN(ybar[200]);
  AND2_X1 U145 ( .A1(b[1]), .A2(a[0]), .ZN(y[1]) );
  OR2_X1 U145bar ( .A1(bbar[1]), .A2(abar[0]), .ZN(ybar[1]);
  AND2_X1 U146 ( .A1(a[1]), .A2(b[3]), .ZN(y[19]) );
  OR2_X1 U146bar ( .A1(abar[1]), .A2(bbar[3]), .ZN(ybar[19]);
  AND2_X1 U147 ( .A1(a[12]), .A2(b[7]), .ZN(y[199]) );
  OR2_X1 U147bar ( .A1(abar[12]), .A2(bbar[7]), .ZN(ybar[199]);
  AND2_X1 U148 ( .A1(a[12]), .A2(b[6]), .ZN(y[198]) );
  OR2_X1 U148bar ( .A1(abar[12]), .A2(bbar[6]), .ZN(ybar[198]);
  AND2_X1 U149 ( .A1(a[12]), .A2(b[5]), .ZN(y[197]) );
  OR2_X1 U149bar ( .A1(abar[12]), .A2(bbar[5]), .ZN(ybar[197]);
  AND2_X1 U150 ( .A1(a[12]), .A2(b[4]), .ZN(y[196]) );
  OR2_X1 U150bar ( .A1(abar[12]), .A2(bbar[4]), .ZN(ybar[196]);
  AND2_X1 U151 ( .A1(a[12]), .A2(b[3]), .ZN(y[195]) );
  OR2_X1 U151bar ( .A1(abar[12]), .A2(bbar[3]), .ZN(ybar[195]);
  AND2_X1 U152 ( .A1(a[12]), .A2(b[2]), .ZN(y[194]) );
  OR2_X1 U152bar ( .A1(abar[12]), .A2(bbar[2]), .ZN(ybar[194]);
  AND2_X1 U153 ( .A1(a[12]), .A2(b[1]), .ZN(y[193]) );
  OR2_X1 U153bar ( .A1(abar[12]), .A2(bbar[1]), .ZN(ybar[193]);
  AND2_X1 U154 ( .A1(a[12]), .A2(b[0]), .ZN(y[192]) );
  OR2_X1 U154bar ( .A1(abar[12]), .A2(bbar[0]), .ZN(ybar[192]);
  AND2_X1 U155 ( .A1(a[11]), .A2(b[15]), .ZN(y[191]) );
  OR2_X1 U155bar ( .A1(abar[11]), .A2(bbar[15]), .ZN(ybar[191]);
  AND2_X1 U156 ( .A1(a[11]), .A2(b[14]), .ZN(y[190]) );
  OR2_X1 U156bar ( .A1(abar[11]), .A2(bbar[14]), .ZN(ybar[190]);
  AND2_X1 U157 ( .A1(a[1]), .A2(b[2]), .ZN(y[18]) );
  OR2_X1 U157bar ( .A1(abar[1]), .A2(bbar[2]), .ZN(ybar[18]);
  AND2_X1 U158 ( .A1(a[11]), .A2(b[13]), .ZN(y[189]) );
  OR2_X1 U158bar ( .A1(abar[11]), .A2(bbar[13]), .ZN(ybar[189]);
  AND2_X1 U159 ( .A1(a[11]), .A2(b[12]), .ZN(y[188]) );
  OR2_X1 U159bar ( .A1(abar[11]), .A2(bbar[12]), .ZN(ybar[188]);
  AND2_X1 U160 ( .A1(a[11]), .A2(b[11]), .ZN(y[187]) );
  OR2_X1 U160bar ( .A1(abar[11]), .A2(bbar[11]), .ZN(ybar[187]);
  AND2_X1 U161 ( .A1(a[11]), .A2(b[10]), .ZN(y[186]) );
  OR2_X1 U161bar ( .A1(abar[11]), .A2(bbar[10]), .ZN(ybar[186]);
  AND2_X1 U162 ( .A1(a[11]), .A2(b[9]), .ZN(y[185]) );
  OR2_X1 U162bar ( .A1(abar[11]), .A2(bbar[9]), .ZN(ybar[185]);
  AND2_X1 U163 ( .A1(a[11]), .A2(b[8]), .ZN(y[184]) );
  OR2_X1 U163bar ( .A1(abar[11]), .A2(bbar[8]), .ZN(ybar[184]);
  AND2_X1 U164 ( .A1(a[11]), .A2(b[7]), .ZN(y[183]) );
  OR2_X1 U164bar ( .A1(abar[11]), .A2(bbar[7]), .ZN(ybar[183]);
  AND2_X1 U165 ( .A1(a[11]), .A2(b[6]), .ZN(y[182]) );
  OR2_X1 U165bar ( .A1(abar[11]), .A2(bbar[6]), .ZN(ybar[182]);
  AND2_X1 U166 ( .A1(a[11]), .A2(b[5]), .ZN(y[181]) );
  OR2_X1 U166bar ( .A1(abar[11]), .A2(bbar[5]), .ZN(ybar[181]);
  AND2_X1 U167 ( .A1(a[11]), .A2(b[4]), .ZN(y[180]) );
  OR2_X1 U167bar ( .A1(abar[11]), .A2(bbar[4]), .ZN(ybar[180]);
  AND2_X1 U168 ( .A1(a[1]), .A2(b[1]), .ZN(y[17]) );
  OR2_X1 U168bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[17]);
  AND2_X1 U169 ( .A1(a[11]), .A2(b[3]), .ZN(y[179]) );
  OR2_X1 U169bar ( .A1(abar[11]), .A2(bbar[3]), .ZN(ybar[179]);
  AND2_X1 U170 ( .A1(a[11]), .A2(b[2]), .ZN(y[178]) );
  OR2_X1 U170bar ( .A1(abar[11]), .A2(bbar[2]), .ZN(ybar[178]);
  AND2_X1 U171 ( .A1(a[11]), .A2(b[1]), .ZN(y[177]) );
  OR2_X1 U171bar ( .A1(abar[11]), .A2(bbar[1]), .ZN(ybar[177]);
  AND2_X1 U172 ( .A1(a[11]), .A2(b[0]), .ZN(y[176]) );
  OR2_X1 U172bar ( .A1(abar[11]), .A2(bbar[0]), .ZN(ybar[176]);
  AND2_X1 U173 ( .A1(a[10]), .A2(b[15]), .ZN(y[175]) );
  OR2_X1 U173bar ( .A1(abar[10]), .A2(bbar[15]), .ZN(ybar[175]);
  AND2_X1 U174 ( .A1(a[10]), .A2(b[14]), .ZN(y[174]) );
  OR2_X1 U174bar ( .A1(abar[10]), .A2(bbar[14]), .ZN(ybar[174]);
  AND2_X1 U175 ( .A1(a[10]), .A2(b[13]), .ZN(y[173]) );
  OR2_X1 U175bar ( .A1(abar[10]), .A2(bbar[13]), .ZN(ybar[173]);
  AND2_X1 U176 ( .A1(a[10]), .A2(b[12]), .ZN(y[172]) );
  OR2_X1 U176bar ( .A1(abar[10]), .A2(bbar[12]), .ZN(ybar[172]);
  AND2_X1 U177 ( .A1(a[10]), .A2(b[11]), .ZN(y[171]) );
  OR2_X1 U177bar ( .A1(abar[10]), .A2(bbar[11]), .ZN(ybar[171]);
  AND2_X1 U178 ( .A1(a[10]), .A2(b[10]), .ZN(y[170]) );
  OR2_X1 U178bar ( .A1(abar[10]), .A2(bbar[10]), .ZN(ybar[170]);
  AND2_X1 U179 ( .A1(a[1]), .A2(b[0]), .ZN(y[16]) );
  OR2_X1 U179bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[16]);
  AND2_X1 U180 ( .A1(a[10]), .A2(b[9]), .ZN(y[169]) );
  OR2_X1 U180bar ( .A1(abar[10]), .A2(bbar[9]), .ZN(ybar[169]);
  AND2_X1 U181 ( .A1(a[10]), .A2(b[8]), .ZN(y[168]) );
  OR2_X1 U181bar ( .A1(abar[10]), .A2(bbar[8]), .ZN(ybar[168]);
  AND2_X1 U182 ( .A1(a[10]), .A2(b[7]), .ZN(y[167]) );
  OR2_X1 U182bar ( .A1(abar[10]), .A2(bbar[7]), .ZN(ybar[167]);
  AND2_X1 U183 ( .A1(a[10]), .A2(b[6]), .ZN(y[166]) );
  OR2_X1 U183bar ( .A1(abar[10]), .A2(bbar[6]), .ZN(ybar[166]);
  AND2_X1 U184 ( .A1(a[10]), .A2(b[5]), .ZN(y[165]) );
  OR2_X1 U184bar ( .A1(abar[10]), .A2(bbar[5]), .ZN(ybar[165]);
  AND2_X1 U185 ( .A1(a[10]), .A2(b[4]), .ZN(y[164]) );
  OR2_X1 U185bar ( .A1(abar[10]), .A2(bbar[4]), .ZN(ybar[164]);
  AND2_X1 U186 ( .A1(a[10]), .A2(b[3]), .ZN(y[163]) );
  OR2_X1 U186bar ( .A1(abar[10]), .A2(bbar[3]), .ZN(ybar[163]);
  AND2_X1 U187 ( .A1(a[10]), .A2(b[2]), .ZN(y[162]) );
  OR2_X1 U187bar ( .A1(abar[10]), .A2(bbar[2]), .ZN(ybar[162]);
  AND2_X1 U188 ( .A1(a[10]), .A2(b[1]), .ZN(y[161]) );
  OR2_X1 U188bar ( .A1(abar[10]), .A2(bbar[1]), .ZN(ybar[161]);
  AND2_X1 U189 ( .A1(a[10]), .A2(b[0]), .ZN(y[160]) );
  OR2_X1 U189bar ( .A1(abar[10]), .A2(bbar[0]), .ZN(ybar[160]);
  AND2_X1 U190 ( .A1(b[15]), .A2(a[0]), .ZN(y[15]) );
  OR2_X1 U190bar ( .A1(bbar[15]), .A2(abar[0]), .ZN(ybar[15]);
  AND2_X1 U191 ( .A1(a[9]), .A2(b[15]), .ZN(y[159]) );
  OR2_X1 U191bar ( .A1(abar[9]), .A2(bbar[15]), .ZN(ybar[159]);
  AND2_X1 U192 ( .A1(a[9]), .A2(b[14]), .ZN(y[158]) );
  OR2_X1 U192bar ( .A1(abar[9]), .A2(bbar[14]), .ZN(ybar[158]);
  AND2_X1 U193 ( .A1(a[9]), .A2(b[13]), .ZN(y[157]) );
  OR2_X1 U193bar ( .A1(abar[9]), .A2(bbar[13]), .ZN(ybar[157]);
  AND2_X1 U194 ( .A1(a[9]), .A2(b[12]), .ZN(y[156]) );
  OR2_X1 U194bar ( .A1(abar[9]), .A2(bbar[12]), .ZN(ybar[156]);
  AND2_X1 U195 ( .A1(a[9]), .A2(b[11]), .ZN(y[155]) );
  OR2_X1 U195bar ( .A1(abar[9]), .A2(bbar[11]), .ZN(ybar[155]);
  AND2_X1 U196 ( .A1(a[9]), .A2(b[10]), .ZN(y[154]) );
  OR2_X1 U196bar ( .A1(abar[9]), .A2(bbar[10]), .ZN(ybar[154]);
  AND2_X1 U197 ( .A1(a[9]), .A2(b[9]), .ZN(y[153]) );
  OR2_X1 U197bar ( .A1(abar[9]), .A2(bbar[9]), .ZN(ybar[153]);
  AND2_X1 U198 ( .A1(a[9]), .A2(b[8]), .ZN(y[152]) );
  OR2_X1 U198bar ( .A1(abar[9]), .A2(bbar[8]), .ZN(ybar[152]);
  AND2_X1 U199 ( .A1(a[9]), .A2(b[7]), .ZN(y[151]) );
  OR2_X1 U199bar ( .A1(abar[9]), .A2(bbar[7]), .ZN(ybar[151]);
  AND2_X1 U200 ( .A1(a[9]), .A2(b[6]), .ZN(y[150]) );
  OR2_X1 U200bar ( .A1(abar[9]), .A2(bbar[6]), .ZN(ybar[150]);
  AND2_X1 U201 ( .A1(b[14]), .A2(a[0]), .ZN(y[14]) );
  OR2_X1 U201bar ( .A1(bbar[14]), .A2(abar[0]), .ZN(ybar[14]);
  AND2_X1 U202 ( .A1(a[9]), .A2(b[5]), .ZN(y[149]) );
  OR2_X1 U202bar ( .A1(abar[9]), .A2(bbar[5]), .ZN(ybar[149]);
  AND2_X1 U203 ( .A1(a[9]), .A2(b[4]), .ZN(y[148]) );
  OR2_X1 U203bar ( .A1(abar[9]), .A2(bbar[4]), .ZN(ybar[148]);
  AND2_X1 U204 ( .A1(a[9]), .A2(b[3]), .ZN(y[147]) );
  OR2_X1 U204bar ( .A1(abar[9]), .A2(bbar[3]), .ZN(ybar[147]);
  AND2_X1 U205 ( .A1(a[9]), .A2(b[2]), .ZN(y[146]) );
  OR2_X1 U205bar ( .A1(abar[9]), .A2(bbar[2]), .ZN(ybar[146]);
  AND2_X1 U206 ( .A1(a[9]), .A2(b[1]), .ZN(y[145]) );
  OR2_X1 U206bar ( .A1(abar[9]), .A2(bbar[1]), .ZN(ybar[145]);
  AND2_X1 U207 ( .A1(a[9]), .A2(b[0]), .ZN(y[144]) );
  OR2_X1 U207bar ( .A1(abar[9]), .A2(bbar[0]), .ZN(ybar[144]);
  AND2_X1 U208 ( .A1(a[8]), .A2(b[15]), .ZN(y[143]) );
  OR2_X1 U208bar ( .A1(abar[8]), .A2(bbar[15]), .ZN(ybar[143]);
  AND2_X1 U209 ( .A1(a[8]), .A2(b[14]), .ZN(y[142]) );
  OR2_X1 U209bar ( .A1(abar[8]), .A2(bbar[14]), .ZN(ybar[142]);
  AND2_X1 U210 ( .A1(a[8]), .A2(b[13]), .ZN(y[141]) );
  OR2_X1 U210bar ( .A1(abar[8]), .A2(bbar[13]), .ZN(ybar[141]);
  AND2_X1 U211 ( .A1(a[8]), .A2(b[12]), .ZN(y[140]) );
  OR2_X1 U211bar ( .A1(abar[8]), .A2(bbar[12]), .ZN(ybar[140]);
  AND2_X1 U212 ( .A1(b[13]), .A2(a[0]), .ZN(y[13]) );
  OR2_X1 U212bar ( .A1(bbar[13]), .A2(abar[0]), .ZN(ybar[13]);
  AND2_X1 U213 ( .A1(a[8]), .A2(b[11]), .ZN(y[139]) );
  OR2_X1 U213bar ( .A1(abar[8]), .A2(bbar[11]), .ZN(ybar[139]);
  AND2_X1 U214 ( .A1(a[8]), .A2(b[10]), .ZN(y[138]) );
  OR2_X1 U214bar ( .A1(abar[8]), .A2(bbar[10]), .ZN(ybar[138]);
  AND2_X1 U215 ( .A1(a[8]), .A2(b[9]), .ZN(y[137]) );
  OR2_X1 U215bar ( .A1(abar[8]), .A2(bbar[9]), .ZN(ybar[137]);
  AND2_X1 U216 ( .A1(a[8]), .A2(b[8]), .ZN(y[136]) );
  OR2_X1 U216bar ( .A1(abar[8]), .A2(bbar[8]), .ZN(ybar[136]);
  AND2_X1 U217 ( .A1(a[8]), .A2(b[7]), .ZN(y[135]) );
  OR2_X1 U217bar ( .A1(abar[8]), .A2(bbar[7]), .ZN(ybar[135]);
  AND2_X1 U218 ( .A1(a[8]), .A2(b[6]), .ZN(y[134]) );
  OR2_X1 U218bar ( .A1(abar[8]), .A2(bbar[6]), .ZN(ybar[134]);
  AND2_X1 U219 ( .A1(a[8]), .A2(b[5]), .ZN(y[133]) );
  OR2_X1 U219bar ( .A1(abar[8]), .A2(bbar[5]), .ZN(ybar[133]);
  AND2_X1 U220 ( .A1(a[8]), .A2(b[4]), .ZN(y[132]) );
  OR2_X1 U220bar ( .A1(abar[8]), .A2(bbar[4]), .ZN(ybar[132]);
  AND2_X1 U221 ( .A1(a[8]), .A2(b[3]), .ZN(y[131]) );
  OR2_X1 U221bar ( .A1(abar[8]), .A2(bbar[3]), .ZN(ybar[131]);
  AND2_X1 U222 ( .A1(a[8]), .A2(b[2]), .ZN(y[130]) );
  OR2_X1 U222bar ( .A1(abar[8]), .A2(bbar[2]), .ZN(ybar[130]);
  AND2_X1 U223 ( .A1(b[12]), .A2(a[0]), .ZN(y[12]) );
  OR2_X1 U223bar ( .A1(bbar[12]), .A2(abar[0]), .ZN(ybar[12]);
  AND2_X1 U224 ( .A1(a[8]), .A2(b[1]), .ZN(y[129]) );
  OR2_X1 U224bar ( .A1(abar[8]), .A2(bbar[1]), .ZN(ybar[129]);
  AND2_X1 U225 ( .A1(a[8]), .A2(b[0]), .ZN(y[128]) );
  OR2_X1 U225bar ( .A1(abar[8]), .A2(bbar[0]), .ZN(ybar[128]);
  AND2_X1 U226 ( .A1(a[7]), .A2(b[15]), .ZN(y[127]) );
  OR2_X1 U226bar ( .A1(abar[7]), .A2(bbar[15]), .ZN(ybar[127]);
  AND2_X1 U227 ( .A1(a[7]), .A2(b[14]), .ZN(y[126]) );
  OR2_X1 U227bar ( .A1(abar[7]), .A2(bbar[14]), .ZN(ybar[126]);
  AND2_X1 U228 ( .A1(a[7]), .A2(b[13]), .ZN(y[125]) );
  OR2_X1 U228bar ( .A1(abar[7]), .A2(bbar[13]), .ZN(ybar[125]);
  AND2_X1 U229 ( .A1(a[7]), .A2(b[12]), .ZN(y[124]) );
  OR2_X1 U229bar ( .A1(abar[7]), .A2(bbar[12]), .ZN(ybar[124]);
  AND2_X1 U230 ( .A1(a[7]), .A2(b[11]), .ZN(y[123]) );
  OR2_X1 U230bar ( .A1(abar[7]), .A2(bbar[11]), .ZN(ybar[123]);
  AND2_X1 U231 ( .A1(a[7]), .A2(b[10]), .ZN(y[122]) );
  OR2_X1 U231bar ( .A1(abar[7]), .A2(bbar[10]), .ZN(ybar[122]);
  AND2_X1 U232 ( .A1(a[7]), .A2(b[9]), .ZN(y[121]) );
  OR2_X1 U232bar ( .A1(abar[7]), .A2(bbar[9]), .ZN(ybar[121]);
  AND2_X1 U233 ( .A1(a[7]), .A2(b[8]), .ZN(y[120]) );
  OR2_X1 U233bar ( .A1(abar[7]), .A2(bbar[8]), .ZN(ybar[120]);
  AND2_X1 U234 ( .A1(b[11]), .A2(a[0]), .ZN(y[11]) );
  OR2_X1 U234bar ( .A1(bbar[11]), .A2(abar[0]), .ZN(ybar[11]);
  AND2_X1 U235 ( .A1(a[7]), .A2(b[7]), .ZN(y[119]) );
  OR2_X1 U235bar ( .A1(abar[7]), .A2(bbar[7]), .ZN(ybar[119]);
  AND2_X1 U236 ( .A1(a[7]), .A2(b[6]), .ZN(y[118]) );
  OR2_X1 U236bar ( .A1(abar[7]), .A2(bbar[6]), .ZN(ybar[118]);
  AND2_X1 U237 ( .A1(a[7]), .A2(b[5]), .ZN(y[117]) );
  OR2_X1 U237bar ( .A1(abar[7]), .A2(bbar[5]), .ZN(ybar[117]);
  AND2_X1 U238 ( .A1(a[7]), .A2(b[4]), .ZN(y[116]) );
  OR2_X1 U238bar ( .A1(abar[7]), .A2(bbar[4]), .ZN(ybar[116]);
  AND2_X1 U239 ( .A1(a[7]), .A2(b[3]), .ZN(y[115]) );
  OR2_X1 U239bar ( .A1(abar[7]), .A2(bbar[3]), .ZN(ybar[115]);
  AND2_X1 U240 ( .A1(a[7]), .A2(b[2]), .ZN(y[114]) );
  OR2_X1 U240bar ( .A1(abar[7]), .A2(bbar[2]), .ZN(ybar[114]);
  AND2_X1 U241 ( .A1(a[7]), .A2(b[1]), .ZN(y[113]) );
  OR2_X1 U241bar ( .A1(abar[7]), .A2(bbar[1]), .ZN(ybar[113]);
  AND2_X1 U242 ( .A1(a[7]), .A2(b[0]), .ZN(y[112]) );
  OR2_X1 U242bar ( .A1(abar[7]), .A2(bbar[0]), .ZN(ybar[112]);
  AND2_X1 U243 ( .A1(b[15]), .A2(a[6]), .ZN(y[111]) );
  OR2_X1 U243bar ( .A1(bbar[15]), .A2(abar[6]), .ZN(ybar[111]);
  AND2_X1 U244 ( .A1(b[14]), .A2(a[6]), .ZN(y[110]) );
  OR2_X1 U244bar ( .A1(bbar[14]), .A2(abar[6]), .ZN(ybar[110]);
  AND2_X1 U245 ( .A1(b[10]), .A2(a[0]), .ZN(y[10]) );
  OR2_X1 U245bar ( .A1(bbar[10]), .A2(abar[0]), .ZN(ybar[10]);
  AND2_X1 U246 ( .A1(b[13]), .A2(a[6]), .ZN(y[109]) );
  OR2_X1 U246bar ( .A1(bbar[13]), .A2(abar[6]), .ZN(ybar[109]);
  AND2_X1 U247 ( .A1(b[12]), .A2(a[6]), .ZN(y[108]) );
  OR2_X1 U247bar ( .A1(bbar[12]), .A2(abar[6]), .ZN(ybar[108]);
  AND2_X1 U248 ( .A1(b[11]), .A2(a[6]), .ZN(y[107]) );
  OR2_X1 U248bar ( .A1(bbar[11]), .A2(abar[6]), .ZN(ybar[107]);
  AND2_X1 U249 ( .A1(b[10]), .A2(a[6]), .ZN(y[106]) );
  OR2_X1 U249bar ( .A1(bbar[10]), .A2(abar[6]), .ZN(ybar[106]);
  AND2_X1 U250 ( .A1(a[6]), .A2(b[9]), .ZN(y[105]) );
  OR2_X1 U250bar ( .A1(abar[6]), .A2(bbar[9]), .ZN(ybar[105]);
  AND2_X1 U251 ( .A1(b[8]), .A2(a[6]), .ZN(y[104]) );
  OR2_X1 U251bar ( .A1(bbar[8]), .A2(abar[6]), .ZN(ybar[104]);
  AND2_X1 U252 ( .A1(b[7]), .A2(a[6]), .ZN(y[103]) );
  OR2_X1 U252bar ( .A1(bbar[7]), .A2(abar[6]), .ZN(ybar[103]);
  AND2_X1 U253 ( .A1(b[6]), .A2(a[6]), .ZN(y[102]) );
  OR2_X1 U253bar ( .A1(bbar[6]), .A2(abar[6]), .ZN(ybar[102]);
  AND2_X1 U254 ( .A1(b[5]), .A2(a[6]), .ZN(y[101]) );
  OR2_X1 U254bar ( .A1(bbar[5]), .A2(abar[6]), .ZN(ybar[101]);
  AND2_X1 U255 ( .A1(b[4]), .A2(a[6]), .ZN(y[100]) );
  OR2_X1 U255bar ( .A1(bbar[4]), .A2(abar[6]), .ZN(ybar[100]);
  AND2_X1 U256 ( .A1(b[0]), .A2(a[0]), .ZN(y[0]) );
  OR2_X1 U256bar ( .A1(bbar[0]), .A2(abar[0]), .ZN(ybar[0]);
endmodule




module decode_12 ( in, out );
  input [7:0] in;
  //input_done

  output [255:0] out;
  //output_done

  wire   [15:0] level1;
  wire   [31:0] level2;
  //wire_done

  CD2_48 cd_l1_1 ( .a(in[1]), .b(in[0]), .y(level1[3:0]) );
  CD2_47 cd_l1_2 ( .a(in[3]), .b(in[2]), .y(level1[7:4]) );
  CD2_46 cd_l1_3 ( .a(in[5]), .b(in[4]), .y(level1[11:8]) );
  CD2_45 cd_l1_4 ( .a(in[7]), .b(in[6]), .y(level1[15:12]) );
  CD4_24 cd_l2_1 ( .a(level1[7:4]), .b(level1[3:0]), .y(level2[15:0]) );
  CD4_23 cd_l2_2 ( .a(level1[15:12]), .b(level1[11:8]), .y(level2[31:16]) );
  CD16_12 cd_l3 ( .a(level2[31:16]), .b(level2[15:0]), .y(out) );
endmodule


module encode_12 ( in, out );
  input [255:0] in;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
  assign inbar[8] = ~in[8];
  assign inbar[9] = ~in[9];
  assign inbar[10] = ~in[10];
  assign inbar[11] = ~in[11];
  assign inbar[12] = ~in[12];
  assign inbar[13] = ~in[13];
  assign inbar[14] = ~in[14];
  assign inbar[15] = ~in[15];
  assign inbar[16] = ~in[16];
  assign inbar[17] = ~in[17];
  assign inbar[18] = ~in[18];
  assign inbar[19] = ~in[19];
  assign inbar[20] = ~in[20];
  assign inbar[21] = ~in[21];
  assign inbar[22] = ~in[22];
  assign inbar[23] = ~in[23];
  assign inbar[24] = ~in[24];
  assign inbar[25] = ~in[25];
  assign inbar[26] = ~in[26];
  assign inbar[27] = ~in[27];
  assign inbar[28] = ~in[28];
  assign inbar[29] = ~in[29];
  assign inbar[30] = ~in[30];
  assign inbar[31] = ~in[31];
  assign inbar[32] = ~in[32];
  assign inbar[33] = ~in[33];
  assign inbar[34] = ~in[34];
  assign inbar[35] = ~in[35];
  assign inbar[36] = ~in[36];
  assign inbar[37] = ~in[37];
  assign inbar[38] = ~in[38];
  assign inbar[39] = ~in[39];
  assign inbar[40] = ~in[40];
  assign inbar[41] = ~in[41];
  assign inbar[42] = ~in[42];
  assign inbar[43] = ~in[43];
  assign inbar[44] = ~in[44];
  assign inbar[45] = ~in[45];
  assign inbar[46] = ~in[46];
  assign inbar[47] = ~in[47];
  assign inbar[48] = ~in[48];
  assign inbar[49] = ~in[49];
  assign inbar[50] = ~in[50];
  assign inbar[51] = ~in[51];
  assign inbar[52] = ~in[52];
  assign inbar[53] = ~in[53];
  assign inbar[54] = ~in[54];
  assign inbar[55] = ~in[55];
  assign inbar[56] = ~in[56];
  assign inbar[57] = ~in[57];
  assign inbar[58] = ~in[58];
  assign inbar[59] = ~in[59];
  assign inbar[60] = ~in[60];
  assign inbar[61] = ~in[61];
  assign inbar[62] = ~in[62];
  assign inbar[63] = ~in[63];
  assign inbar[64] = ~in[64];
  assign inbar[65] = ~in[65];
  assign inbar[66] = ~in[66];
  assign inbar[67] = ~in[67];
  assign inbar[68] = ~in[68];
  assign inbar[69] = ~in[69];
  assign inbar[70] = ~in[70];
  assign inbar[71] = ~in[71];
  assign inbar[72] = ~in[72];
  assign inbar[73] = ~in[73];
  assign inbar[74] = ~in[74];
  assign inbar[75] = ~in[75];
  assign inbar[76] = ~in[76];
  assign inbar[77] = ~in[77];
  assign inbar[78] = ~in[78];
  assign inbar[79] = ~in[79];
  assign inbar[80] = ~in[80];
  assign inbar[81] = ~in[81];
  assign inbar[82] = ~in[82];
  assign inbar[83] = ~in[83];
  assign inbar[84] = ~in[84];
  assign inbar[85] = ~in[85];
  assign inbar[86] = ~in[86];
  assign inbar[87] = ~in[87];
  assign inbar[88] = ~in[88];
  assign inbar[89] = ~in[89];
  assign inbar[90] = ~in[90];
  assign inbar[91] = ~in[91];
  assign inbar[92] = ~in[92];
  assign inbar[93] = ~in[93];
  assign inbar[94] = ~in[94];
  assign inbar[95] = ~in[95];
  assign inbar[96] = ~in[96];
  assign inbar[97] = ~in[97];
  assign inbar[98] = ~in[98];
  assign inbar[99] = ~in[99];
  assign inbar[100] = ~in[100];
  assign inbar[101] = ~in[101];
  assign inbar[102] = ~in[102];
  assign inbar[103] = ~in[103];
  assign inbar[104] = ~in[104];
  assign inbar[105] = ~in[105];
  assign inbar[106] = ~in[106];
  assign inbar[107] = ~in[107];
  assign inbar[108] = ~in[108];
  assign inbar[109] = ~in[109];
  assign inbar[110] = ~in[110];
  assign inbar[111] = ~in[111];
  assign inbar[112] = ~in[112];
  assign inbar[113] = ~in[113];
  assign inbar[114] = ~in[114];
  assign inbar[115] = ~in[115];
  assign inbar[116] = ~in[116];
  assign inbar[117] = ~in[117];
  assign inbar[118] = ~in[118];
  assign inbar[119] = ~in[119];
  assign inbar[120] = ~in[120];
  assign inbar[121] = ~in[121];
  assign inbar[122] = ~in[122];
  assign inbar[123] = ~in[123];
  assign inbar[124] = ~in[124];
  assign inbar[125] = ~in[125];
  assign inbar[126] = ~in[126];
  assign inbar[127] = ~in[127];
  assign inbar[128] = ~in[128];
  assign inbar[129] = ~in[129];
  assign inbar[130] = ~in[130];
  assign inbar[131] = ~in[131];
  assign inbar[132] = ~in[132];
  assign inbar[133] = ~in[133];
  assign inbar[134] = ~in[134];
  assign inbar[135] = ~in[135];
  assign inbar[136] = ~in[136];
  assign inbar[137] = ~in[137];
  assign inbar[138] = ~in[138];
  assign inbar[139] = ~in[139];
  assign inbar[140] = ~in[140];
  assign inbar[141] = ~in[141];
  assign inbar[142] = ~in[142];
  assign inbar[143] = ~in[143];
  assign inbar[144] = ~in[144];
  assign inbar[145] = ~in[145];
  assign inbar[146] = ~in[146];
  assign inbar[147] = ~in[147];
  assign inbar[148] = ~in[148];
  assign inbar[149] = ~in[149];
  assign inbar[150] = ~in[150];
  assign inbar[151] = ~in[151];
  assign inbar[152] = ~in[152];
  assign inbar[153] = ~in[153];
  assign inbar[154] = ~in[154];
  assign inbar[155] = ~in[155];
  assign inbar[156] = ~in[156];
  assign inbar[157] = ~in[157];
  assign inbar[158] = ~in[158];
  assign inbar[159] = ~in[159];
  assign inbar[160] = ~in[160];
  assign inbar[161] = ~in[161];
  assign inbar[162] = ~in[162];
  assign inbar[163] = ~in[163];
  assign inbar[164] = ~in[164];
  assign inbar[165] = ~in[165];
  assign inbar[166] = ~in[166];
  assign inbar[167] = ~in[167];
  assign inbar[168] = ~in[168];
  assign inbar[169] = ~in[169];
  assign inbar[170] = ~in[170];
  assign inbar[171] = ~in[171];
  assign inbar[172] = ~in[172];
  assign inbar[173] = ~in[173];
  assign inbar[174] = ~in[174];
  assign inbar[175] = ~in[175];
  assign inbar[176] = ~in[176];
  assign inbar[177] = ~in[177];
  assign inbar[178] = ~in[178];
  assign inbar[179] = ~in[179];
  assign inbar[180] = ~in[180];
  assign inbar[181] = ~in[181];
  assign inbar[182] = ~in[182];
  assign inbar[183] = ~in[183];
  assign inbar[184] = ~in[184];
  assign inbar[185] = ~in[185];
  assign inbar[186] = ~in[186];
  assign inbar[187] = ~in[187];
  assign inbar[188] = ~in[188];
  assign inbar[189] = ~in[189];
  assign inbar[190] = ~in[190];
  assign inbar[191] = ~in[191];
  assign inbar[192] = ~in[192];
  assign inbar[193] = ~in[193];
  assign inbar[194] = ~in[194];
  assign inbar[195] = ~in[195];
  assign inbar[196] = ~in[196];
  assign inbar[197] = ~in[197];
  assign inbar[198] = ~in[198];
  assign inbar[199] = ~in[199];
  assign inbar[200] = ~in[200];
  assign inbar[201] = ~in[201];
  assign inbar[202] = ~in[202];
  assign inbar[203] = ~in[203];
  assign inbar[204] = ~in[204];
  assign inbar[205] = ~in[205];
  assign inbar[206] = ~in[206];
  assign inbar[207] = ~in[207];
  assign inbar[208] = ~in[208];
  assign inbar[209] = ~in[209];
  assign inbar[210] = ~in[210];
  assign inbar[211] = ~in[211];
  assign inbar[212] = ~in[212];
  assign inbar[213] = ~in[213];
  assign inbar[214] = ~in[214];
  assign inbar[215] = ~in[215];
  assign inbar[216] = ~in[216];
  assign inbar[217] = ~in[217];
  assign inbar[218] = ~in[218];
  assign inbar[219] = ~in[219];
  assign inbar[220] = ~in[220];
  assign inbar[221] = ~in[221];
  assign inbar[222] = ~in[222];
  assign inbar[223] = ~in[223];
  assign inbar[224] = ~in[224];
  assign inbar[225] = ~in[225];
  assign inbar[226] = ~in[226];
  assign inbar[227] = ~in[227];
  assign inbar[228] = ~in[228];
  assign inbar[229] = ~in[229];
  assign inbar[230] = ~in[230];
  assign inbar[231] = ~in[231];
  assign inbar[232] = ~in[232];
  assign inbar[233] = ~in[233];
  assign inbar[234] = ~in[234];
  assign inbar[235] = ~in[235];
  assign inbar[236] = ~in[236];
  assign inbar[237] = ~in[237];
  assign inbar[238] = ~in[238];
  assign inbar[239] = ~in[239];
  assign inbar[240] = ~in[240];
  assign inbar[241] = ~in[241];
  assign inbar[242] = ~in[242];
  assign inbar[243] = ~in[243];
  assign inbar[244] = ~in[244];
  assign inbar[245] = ~in[245];
  assign inbar[246] = ~in[246];
  assign inbar[247] = ~in[247];
  assign inbar[248] = ~in[248];
  assign inbar[249] = ~in[249];
  assign inbar[250] = ~in[250];
  assign inbar[251] = ~in[251];
  assign inbar[252] = ~in[252];
  assign inbar[253] = ~in[253];
  assign inbar[254] = ~in[254];
  assign inbar[255] = ~in[255];
  //input_done

  output [7:0] out;
  reg [7:0] outbar;
  //output_done

  wire   in_81, in_80, in_79, in_78, in_77, in_76, in_75, in_74, in_73, in_72,
         in_71, in_70, in_69, in_68, in_67, in_66, in_65, in_64, in_63, in_62,
         in_61, in_60, in_59, in_58, in_57, in_56, in_55, in_54, in_53, in_52,
         in_51, in_50, in_49, in_48, in_47, in_46, in_45, in_44, in_43, in_42,
         in_41, in_40, in_39, in_38, in_37, in_36, in_35, in_34, in_33, in_32,
         in_31, in_30, in_29, in_28, in_27, in_26, in_25, in_24, in_23, in_22,
         in_21, in_20, in_19, in_18, in_17, in_16, in_15, in_14, in_13, in_12,
         in_11, in_10, in_9, in_8, in_7, in_6, in_5, in_4, in_3, in_2, in_1,
         in_0, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972;
  wire in_81bar, in_80bar, in_79bar, in_78bar, in_77bar, in_76bar, in_75bar, in_74bar, in_73bar, in_72bar, in_71bar, in_70bar, in_69bar, in_68bar, in_67bar, in_66bar, in_65bar, in_64bar, in_63bar, in_62bar, in_61bar, in_60bar, in_59bar, in_58bar, in_57bar, in_56bar, in_55bar, in_54bar, in_53bar, in_52bar, in_51bar, in_50bar, in_49bar, in_48bar, in_47bar, in_46bar, in_45bar, in_44bar, in_43bar, in_42bar, in_41bar, in_40bar, in_39bar, in_38bar, in_37bar, in_36bar, in_35bar, in_34bar, in_33bar, in_32bar, in_31bar, in_30bar, in_29bar, in_28bar, in_27bar, in_26bar, in_25bar, in_24bar, in_23bar, in_22bar, in_21bar, in_20bar, in_19bar, in_18bar, in_17bar, in_16bar, in_15bar, in_14bar, in_13bar, in_12bar, in_11bar, in_10bar, in_9bar, in_8bar, in_7bar, in_6bar, in_5bar, in_4bar, in_3bar, in_2bar, in_1bar, in_0bar, n487bar, n488bar, n489bar, n490bar, n491bar, n492bar, n493bar, n494bar, n495bar, n496bar, n497bar, n498bar, n499bar, n500bar, n501bar, n502bar, n503bar, n504bar, n505bar, n506bar, n507bar, n508bar, n509bar, n510bar, n511bar, n512bar, n513bar, n514bar, n515bar, n516bar, n517bar, n518bar, n519bar, n520bar, n521bar, n522bar, n523bar, n524bar, n525bar, n526bar, n527bar, n528bar, n529bar, n530bar, n531bar, n532bar, n533bar, n534bar, n535bar, n536bar, n537bar, n538bar, n539bar, n540bar, n541bar, n542bar, n543bar, n544bar, n545bar, n546bar, n547bar, n548bar, n549bar, n550bar, n551bar, n552bar, n553bar, n554bar, n555bar, n556bar, n557bar, n558bar, n559bar, n560bar, n561bar, n562bar, n563bar, n564bar, n565bar, n566bar, n567bar, n568bar, n569bar, n570bar, n571bar, n572bar, n573bar, n574bar, n575bar, n576bar, n577bar, n578bar, n579bar, n580bar, n581bar, n582bar, n583bar, n584bar, n585bar, n586bar, n587bar, n588bar, n589bar, n590bar, n591bar, n592bar, n593bar, n594bar, n595bar, n596bar, n597bar, n598bar, n599bar, n600bar, n601bar, n602bar, n603bar, n604bar, n605bar, n606bar, n607bar, n608bar, n609bar, n610bar, n611bar, n612bar, n613bar, n614bar, n615bar, n616bar, n617bar, n618bar, n619bar, n620bar, n621bar, n622bar, n623bar, n624bar, n625bar, n626bar, n627bar, n628bar, n629bar, n630bar, n631bar, n632bar, n633bar, n634bar, n635bar, n636bar, n637bar, n638bar, n639bar, n640bar, n641bar, n642bar, n643bar, n644bar, n645bar, n646bar, n647bar, n648bar, n649bar, n650bar, n651bar, n652bar, n653bar, n654bar, n655bar, n656bar, n657bar, n658bar, n659bar, n660bar, n661bar, n662bar, n663bar, n664bar, n665bar, n666bar, n667bar, n668bar, n669bar, n670bar, n671bar, n672bar, n673bar, n674bar, n675bar, n676bar, n677bar, n678bar, n679bar, n680bar, n681bar, n682bar, n683bar, n684bar, n685bar, n686bar, n687bar, n688bar, n689bar, n690bar, n691bar, n692bar, n693bar, n694bar, n695bar, n696bar, n697bar, n698bar, n699bar, n700bar, n701bar, n702bar, n703bar, n704bar, n705bar, n706bar, n707bar, n708bar, n709bar, n710bar, n711bar, n712bar, n713bar, n714bar, n715bar, n716bar, n717bar, n718bar, n719bar, n720bar, n721bar, n722bar, n723bar, n724bar, n725bar, n726bar, n727bar, n728bar, n729bar, n730bar, n731bar, n732bar, n733bar, n734bar, n735bar, n736bar, n737bar, n738bar, n739bar, n740bar, n741bar, n742bar, n743bar, n744bar, n745bar, n746bar, n747bar, n748bar, n749bar, n750bar, n751bar, n752bar, n753bar, n754bar, n755bar, n756bar, n757bar, n758bar, n759bar, n760bar, n761bar, n762bar, n763bar, n764bar, n765bar, n766bar, n767bar, n768bar, n769bar, n770bar, n771bar, n772bar, n773bar, n774bar, n775bar, n776bar, n777bar, n778bar, n779bar, n780bar, n781bar, n782bar, n783bar, n784bar, n785bar, n786bar, n787bar, n788bar, n789bar, n790bar, n791bar, n792bar, n793bar, n794bar, n795bar, n796bar, n797bar, n798bar, n799bar, n800bar, n801bar, n802bar, n803bar, n804bar, n805bar, n806bar, n807bar, n808bar, n809bar, n810bar, n811bar, n812bar, n813bar, n814bar, n815bar, n816bar, n817bar, n818bar, n819bar, n820bar, n821bar, n822bar, n823bar, n824bar, n825bar, n826bar, n827bar, n828bar, n829bar, n830bar, n831bar, n832bar, n833bar, n834bar, n835bar, n836bar, n837bar, n838bar, n839bar, n840bar, n841bar, n842bar, n843bar, n844bar, n845bar, n846bar, n847bar, n848bar, n849bar, n850bar, n851bar, n852bar, n853bar, n854bar, n855bar, n856bar, n857bar, n858bar, n859bar, n860bar, n861bar, n862bar, n863bar, n864bar, n865bar, n866bar, n867bar, n868bar, n869bar, n870bar, n871bar, n872bar, n873bar, n874bar, n875bar, n876bar, n877bar, n878bar, n879bar, n880bar, n881bar, n882bar, n883bar, n884bar, n885bar, n886bar, n887bar, n888bar, n889bar, n890bar, n891bar, n892bar, n893bar, n894bar, n895bar, n896bar, n897bar, n898bar, n899bar, n900bar, n901bar, n902bar, n903bar, n904bar, n905bar, n906bar, n907bar, n908bar, n909bar, n910bar, n911bar, n912bar, n913bar, n914bar, n915bar, n916bar, n917bar, n918bar, n919bar, n920bar, n921bar, n922bar, n923bar, n924bar, n925bar, n926bar, n927bar, n928bar, n929bar, n930bar, n931bar, n932bar, n933bar, n934bar, n935bar, n936bar, n937bar, n938bar, n939bar, n940bar, n941bar, n942bar, n943bar, n944bar, n945bar, n946bar, n947bar, n948bar, n949bar, n950bar, n951bar, n952bar, n953bar, n954bar, n955bar, n956bar, n957bar, n958bar, n959bar, n960bar, n961bar, n962bar, n963bar, n964bar, n965bar, n966bar, n967bar, n968bar, n969bar, n970bar, n971bar, n972bar;
  //wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];

  OR2_X1 U1 ( .A1(n972), .A2(n971), .ZN(out[7]) );
  AND2_X1 U1bar ( .A1(n972bar), .A2(n971bar), .ZN(outbar[7]);
  OR2_X1 U2 ( .A1(n970), .A2(n969), .ZN(n971) );
  AND2_X1 U2bar ( .A1(n970bar), .A2(n969bar), .ZN(n971bar);
  OR2_X1 U3 ( .A1(n968), .A2(n967), .ZN(n969) );
  AND2_X1 U3bar ( .A1(n968bar), .A2(n967bar), .ZN(n969bar);
  OR2_X1 U4 ( .A1(n966), .A2(n965), .ZN(n967) );
  AND2_X1 U4bar ( .A1(n966bar), .A2(n965bar), .ZN(n967bar);
  OR2_X1 U5 ( .A1(n964), .A2(n963), .ZN(n968) );
  AND2_X1 U5bar ( .A1(n964bar), .A2(n963bar), .ZN(n968bar);
  OR2_X1 U6 ( .A1(in[116]), .A2(n962), .ZN(n963) );
  AND2_X1 U6bar ( .A1(inbar[116]), .A2(n962bar), .ZN(n963bar);
  OR2_X1 U7 ( .A1(n961), .A2(n960), .ZN(n970) );
  AND2_X1 U7bar ( .A1(n961bar), .A2(n960bar), .ZN(n970bar);
  OR2_X1 U8 ( .A1(in[150]), .A2(in[127]), .ZN(n960) );
  AND2_X1 U8bar ( .A1(inbar[150]), .A2(inbar[127]), .ZN(n960bar);
  OR2_X1 U9 ( .A1(in[160]), .A2(n959), .ZN(n961) );
  AND2_X1 U9bar ( .A1(inbar[160]), .A2(n959bar), .ZN(n961bar);
  OR2_X1 U10 ( .A1(in[252]), .A2(in[168]), .ZN(n959) );
  AND2_X1 U10bar ( .A1(inbar[252]), .A2(inbar[168]), .ZN(n959bar);
  OR2_X1 U11 ( .A1(n958), .A2(n957), .ZN(n972) );
  AND2_X1 U11bar ( .A1(n958bar), .A2(n957bar), .ZN(n972bar);
  OR2_X1 U12 ( .A1(n956), .A2(n955), .ZN(n957) );
  AND2_X1 U12bar ( .A1(n956bar), .A2(n955bar), .ZN(n957bar);
  OR2_X1 U13 ( .A1(in_17), .A2(in[96]), .ZN(n955) );
  AND2_X1 U13bar ( .A1(in_17bar), .A2(inbar[96]), .ZN(n955bar);
  OR2_X1 U14 ( .A1(in_23), .A2(n954), .ZN(n956) );
  AND2_X1 U14bar ( .A1(in_23bar), .A2(n954bar), .ZN(n956bar);
  OR2_X1 U15 ( .A1(in_31), .A2(in_26), .ZN(n954) );
  AND2_X1 U15bar ( .A1(in_31bar), .A2(in_26bar), .ZN(n954bar);
  OR2_X1 U16 ( .A1(n953), .A2(n952), .ZN(n958) );
  AND2_X1 U16bar ( .A1(n953bar), .A2(n952bar), .ZN(n958bar);
  OR2_X1 U17 ( .A1(in_58), .A2(in_4), .ZN(n952) );
  AND2_X1 U17bar ( .A1(in_58bar), .A2(in_4bar), .ZN(n952bar);
  OR2_X1 U18 ( .A1(in_59), .A2(n951), .ZN(n953) );
  AND2_X1 U18bar ( .A1(in_59bar), .A2(n951bar), .ZN(n953bar);
  OR2_X1 U19 ( .A1(in_71), .A2(in_62), .ZN(n951) );
  AND2_X1 U19bar ( .A1(in_71bar), .A2(in_62bar), .ZN(n951bar);
  OR2_X1 U20 ( .A1(n950), .A2(n949), .ZN(out[6]) );
  AND2_X1 U20bar ( .A1(n950bar), .A2(n949bar), .ZN(outbar[6]);
  OR2_X1 U21 ( .A1(n948), .A2(n947), .ZN(n949) );
  AND2_X1 U21bar ( .A1(n948bar), .A2(n947bar), .ZN(n949bar);
  OR2_X1 U22 ( .A1(n946), .A2(n945), .ZN(n947) );
  AND2_X1 U22bar ( .A1(n946bar), .A2(n945bar), .ZN(n947bar);
  OR2_X1 U23 ( .A1(n944), .A2(n943), .ZN(n945) );
  AND2_X1 U23bar ( .A1(n944bar), .A2(n943bar), .ZN(n945bar);
  OR2_X1 U24 ( .A1(n942), .A2(n941), .ZN(n946) );
  AND2_X1 U24bar ( .A1(n942bar), .A2(n941bar), .ZN(n946bar);
  OR2_X1 U25 ( .A1(in[101]), .A2(n940), .ZN(n941) );
  AND2_X1 U25bar ( .A1(inbar[101]), .A2(n940bar), .ZN(n941bar);
  OR2_X1 U26 ( .A1(n939), .A2(n938), .ZN(n948) );
  AND2_X1 U26bar ( .A1(n939bar), .A2(n938bar), .ZN(n948bar);
  OR2_X1 U27 ( .A1(in[114]), .A2(in[104]), .ZN(n938) );
  AND2_X1 U27bar ( .A1(inbar[114]), .A2(inbar[104]), .ZN(n938bar);
  OR2_X1 U28 ( .A1(in[128]), .A2(n937), .ZN(n939) );
  AND2_X1 U28bar ( .A1(inbar[128]), .A2(n937bar), .ZN(n939bar);
  OR2_X1 U29 ( .A1(in[136]), .A2(in[134]), .ZN(n937) );
  AND2_X1 U29bar ( .A1(inbar[136]), .A2(inbar[134]), .ZN(n937bar);
  OR2_X1 U30 ( .A1(n936), .A2(n935), .ZN(n950) );
  AND2_X1 U30bar ( .A1(n936bar), .A2(n935bar), .ZN(n950bar);
  OR2_X1 U31 ( .A1(n934), .A2(n933), .ZN(n935) );
  AND2_X1 U31bar ( .A1(n934bar), .A2(n933bar), .ZN(n935bar);
  OR2_X1 U32 ( .A1(in[177]), .A2(in[164]), .ZN(n933) );
  AND2_X1 U32bar ( .A1(inbar[177]), .A2(inbar[164]), .ZN(n933bar);
  OR2_X1 U33 ( .A1(in[212]), .A2(n932), .ZN(n934) );
  AND2_X1 U33bar ( .A1(inbar[212]), .A2(n932bar), .ZN(n934bar);
  OR2_X1 U34 ( .A1(in[248]), .A2(in[221]), .ZN(n932) );
  AND2_X1 U34bar ( .A1(inbar[248]), .A2(inbar[221]), .ZN(n932bar);
  OR2_X1 U35 ( .A1(n931), .A2(n930), .ZN(n936) );
  AND2_X1 U35bar ( .A1(n931bar), .A2(n930bar), .ZN(n936bar);
  OR2_X1 U36 ( .A1(in_18), .A2(in[93]), .ZN(n930) );
  AND2_X1 U36bar ( .A1(in_18bar), .A2(inbar[93]), .ZN(n930bar);
  OR2_X1 U37 ( .A1(in_31), .A2(n929), .ZN(n931) );
  AND2_X1 U37bar ( .A1(in_31bar), .A2(n929bar), .ZN(n931bar);
  OR2_X1 U38 ( .A1(in_7), .A2(in_39), .ZN(n929) );
  AND2_X1 U38bar ( .A1(in_7bar), .A2(in_39bar), .ZN(n929bar);
  OR2_X1 U39 ( .A1(n928), .A2(n927), .ZN(out[5]) );
  AND2_X1 U39bar ( .A1(n928bar), .A2(n927bar), .ZN(outbar[5]);
  OR2_X1 U40 ( .A1(n926), .A2(n925), .ZN(n927) );
  AND2_X1 U40bar ( .A1(n926bar), .A2(n925bar), .ZN(n927bar);
  OR2_X1 U41 ( .A1(n924), .A2(n923), .ZN(n925) );
  AND2_X1 U41bar ( .A1(n924bar), .A2(n923bar), .ZN(n925bar);
  OR2_X1 U42 ( .A1(n922), .A2(n921), .ZN(n923) );
  AND2_X1 U42bar ( .A1(n922bar), .A2(n921bar), .ZN(n923bar);
  OR2_X1 U43 ( .A1(n940), .A2(n920), .ZN(n924) );
  AND2_X1 U43bar ( .A1(n940bar), .A2(n920bar), .ZN(n924bar);
  OR2_X1 U44 ( .A1(in[111]), .A2(n919), .ZN(n920) );
  AND2_X1 U44bar ( .A1(inbar[111]), .A2(n919bar), .ZN(n920bar);
  OR2_X1 U45 ( .A1(n918), .A2(n917), .ZN(n940) );
  AND2_X1 U45bar ( .A1(n918bar), .A2(n917bar), .ZN(n940bar);
  OR2_X1 U46 ( .A1(n916), .A2(n915), .ZN(n917) );
  AND2_X1 U46bar ( .A1(n916bar), .A2(n915bar), .ZN(n917bar);
  OR2_X1 U47 ( .A1(n914), .A2(n913), .ZN(n915) );
  AND2_X1 U47bar ( .A1(n914bar), .A2(n913bar), .ZN(n915bar);
  OR2_X1 U48 ( .A1(in[140]), .A2(in[131]), .ZN(n913) );
  AND2_X1 U48bar ( .A1(inbar[140]), .A2(inbar[131]), .ZN(n913bar);
  OR2_X1 U49 ( .A1(in[160]), .A2(in[144]), .ZN(n914) );
  AND2_X1 U49bar ( .A1(inbar[160]), .A2(inbar[144]), .ZN(n914bar);
  OR2_X1 U50 ( .A1(n912), .A2(n911), .ZN(n916) );
  AND2_X1 U50bar ( .A1(n912bar), .A2(n911bar), .ZN(n916bar);
  OR2_X1 U51 ( .A1(in[179]), .A2(in[174]), .ZN(n911) );
  AND2_X1 U51bar ( .A1(inbar[179]), .A2(inbar[174]), .ZN(n911bar);
  OR2_X1 U52 ( .A1(in[188]), .A2(in[184]), .ZN(n912) );
  AND2_X1 U52bar ( .A1(inbar[188]), .A2(inbar[184]), .ZN(n912bar);
  OR2_X1 U53 ( .A1(n910), .A2(n909), .ZN(n918) );
  AND2_X1 U53bar ( .A1(n910bar), .A2(n909bar), .ZN(n918bar);
  OR2_X1 U54 ( .A1(n908), .A2(n907), .ZN(n909) );
  AND2_X1 U54bar ( .A1(n908bar), .A2(n907bar), .ZN(n909bar);
  OR2_X1 U55 ( .A1(in[216]), .A2(in[200]), .ZN(n907) );
  AND2_X1 U55bar ( .A1(inbar[216]), .A2(inbar[200]), .ZN(n907bar);
  OR2_X1 U56 ( .A1(in[228]), .A2(in[224]), .ZN(n908) );
  AND2_X1 U56bar ( .A1(inbar[228]), .A2(inbar[224]), .ZN(n908bar);
  OR2_X1 U57 ( .A1(n906), .A2(n905), .ZN(n910) );
  AND2_X1 U57bar ( .A1(n906bar), .A2(n905bar), .ZN(n910bar);
  OR2_X1 U58 ( .A1(in[247]), .A2(in[235]), .ZN(n905) );
  AND2_X1 U58bar ( .A1(inbar[247]), .A2(inbar[235]), .ZN(n905bar);
  OR2_X1 U59 ( .A1(in_42), .A2(in[83]), .ZN(n906) );
  AND2_X1 U59bar ( .A1(in_42bar), .A2(inbar[83]), .ZN(n906bar);
  OR2_X1 U60 ( .A1(n904), .A2(n903), .ZN(n926) );
  AND2_X1 U60bar ( .A1(n904bar), .A2(n903bar), .ZN(n926bar);
  OR2_X1 U61 ( .A1(in[166]), .A2(in[123]), .ZN(n903) );
  AND2_X1 U61bar ( .A1(inbar[166]), .A2(inbar[123]), .ZN(n903bar);
  OR2_X1 U62 ( .A1(in[170]), .A2(n902), .ZN(n904) );
  AND2_X1 U62bar ( .A1(inbar[170]), .A2(n902bar), .ZN(n904bar);
  OR2_X1 U63 ( .A1(in[194]), .A2(in[183]), .ZN(n902) );
  AND2_X1 U63bar ( .A1(inbar[194]), .A2(inbar[183]), .ZN(n902bar);
  OR2_X1 U64 ( .A1(n901), .A2(n900), .ZN(n928) );
  AND2_X1 U64bar ( .A1(n901bar), .A2(n900bar), .ZN(n928bar);
  OR2_X1 U65 ( .A1(n899), .A2(n898), .ZN(n900) );
  AND2_X1 U65bar ( .A1(n899bar), .A2(n898bar), .ZN(n900bar);
  OR2_X1 U66 ( .A1(in[241]), .A2(in[238]), .ZN(n898) );
  AND2_X1 U66bar ( .A1(inbar[241]), .A2(inbar[238]), .ZN(n898bar);
  OR2_X1 U67 ( .A1(in[250]), .A2(n897), .ZN(n899) );
  AND2_X1 U67bar ( .A1(inbar[250]), .A2(n897bar), .ZN(n899bar);
  OR2_X1 U68 ( .A1(in_24), .A2(in[84]), .ZN(n897) );
  AND2_X1 U68bar ( .A1(in_24bar), .A2(inbar[84]), .ZN(n897bar);
  OR2_X1 U69 ( .A1(n896), .A2(n895), .ZN(n901) );
  AND2_X1 U69bar ( .A1(n896bar), .A2(n895bar), .ZN(n901bar);
  OR2_X1 U70 ( .A1(in_41), .A2(in_29), .ZN(n895) );
  AND2_X1 U70bar ( .A1(in_41bar), .A2(in_29bar), .ZN(n895bar);
  OR2_X1 U71 ( .A1(in_66), .A2(n894), .ZN(n896) );
  AND2_X1 U71bar ( .A1(in_66bar), .A2(n894bar), .ZN(n896bar);
  OR2_X1 U72 ( .A1(in_76), .A2(in_71), .ZN(n894) );
  AND2_X1 U72bar ( .A1(in_76bar), .A2(in_71bar), .ZN(n894bar);
  OR2_X1 U73 ( .A1(n893), .A2(n892), .ZN(out[4]) );
  AND2_X1 U73bar ( .A1(n893bar), .A2(n892bar), .ZN(outbar[4]);
  OR2_X1 U74 ( .A1(n891), .A2(n890), .ZN(n892) );
  AND2_X1 U74bar ( .A1(n891bar), .A2(n890bar), .ZN(n892bar);
  OR2_X1 U75 ( .A1(n889), .A2(n888), .ZN(n890) );
  AND2_X1 U75bar ( .A1(n889bar), .A2(n888bar), .ZN(n890bar);
  OR2_X1 U76 ( .A1(n922), .A2(n887), .ZN(n888) );
  AND2_X1 U76bar ( .A1(n922bar), .A2(n887bar), .ZN(n888bar);
  OR2_X1 U77 ( .A1(n886), .A2(n885), .ZN(n922) );
  AND2_X1 U77bar ( .A1(n886bar), .A2(n885bar), .ZN(n922bar);
  OR2_X1 U78 ( .A1(n884), .A2(n883), .ZN(n885) );
  AND2_X1 U78bar ( .A1(n884bar), .A2(n883bar), .ZN(n885bar);
  OR2_X1 U79 ( .A1(n882), .A2(n881), .ZN(n883) );
  AND2_X1 U79bar ( .A1(n882bar), .A2(n881bar), .ZN(n883bar);
  OR2_X1 U80 ( .A1(in[118]), .A2(in[109]), .ZN(n881) );
  AND2_X1 U80bar ( .A1(inbar[118]), .A2(inbar[109]), .ZN(n881bar);
  OR2_X1 U81 ( .A1(in[139]), .A2(in[120]), .ZN(n882) );
  AND2_X1 U81bar ( .A1(inbar[139]), .A2(inbar[120]), .ZN(n882bar);
  OR2_X1 U82 ( .A1(n880), .A2(n879), .ZN(n884) );
  AND2_X1 U82bar ( .A1(n880bar), .A2(n879bar), .ZN(n884bar);
  OR2_X1 U83 ( .A1(in[198]), .A2(in[154]), .ZN(n879) );
  AND2_X1 U83bar ( .A1(inbar[198]), .A2(inbar[154]), .ZN(n879bar);
  OR2_X1 U84 ( .A1(in[210]), .A2(in[205]), .ZN(n880) );
  AND2_X1 U84bar ( .A1(inbar[210]), .A2(inbar[205]), .ZN(n880bar);
  OR2_X1 U85 ( .A1(n878), .A2(n877), .ZN(n886) );
  AND2_X1 U85bar ( .A1(n878bar), .A2(n877bar), .ZN(n886bar);
  OR2_X1 U86 ( .A1(n876), .A2(n875), .ZN(n877) );
  AND2_X1 U86bar ( .A1(n876bar), .A2(n875bar), .ZN(n877bar);
  OR2_X1 U87 ( .A1(in[219]), .A2(in[217]), .ZN(n875) );
  AND2_X1 U87bar ( .A1(inbar[219]), .A2(inbar[217]), .ZN(n875bar);
  OR2_X1 U88 ( .A1(in[86]), .A2(in[252]), .ZN(n876) );
  AND2_X1 U88bar ( .A1(inbar[86]), .A2(inbar[252]), .ZN(n876bar);
  OR2_X1 U89 ( .A1(n874), .A2(n873), .ZN(n878) );
  AND2_X1 U89bar ( .A1(n874bar), .A2(n873bar), .ZN(n878bar);
  OR2_X1 U90 ( .A1(in_40), .A2(in[91]), .ZN(n873) );
  AND2_X1 U90bar ( .A1(in_40bar), .A2(inbar[91]), .ZN(n873bar);
  OR2_X1 U91 ( .A1(in_8), .A2(in_46), .ZN(n874) );
  AND2_X1 U91bar ( .A1(in_8bar), .A2(in_46bar), .ZN(n874bar);
  OR2_X1 U92 ( .A1(n872), .A2(n871), .ZN(n889) );
  AND2_X1 U92bar ( .A1(n872bar), .A2(n871bar), .ZN(n889bar);
  OR2_X1 U93 ( .A1(in[117]), .A2(n943), .ZN(n871) );
  AND2_X1 U93bar ( .A1(inbar[117]), .A2(n943bar), .ZN(n871bar);
  OR2_X1 U94 ( .A1(n870), .A2(n869), .ZN(n943) );
  AND2_X1 U94bar ( .A1(n870bar), .A2(n869bar), .ZN(n943bar);
  OR2_X1 U95 ( .A1(n868), .A2(n867), .ZN(n869) );
  AND2_X1 U95bar ( .A1(n868bar), .A2(n867bar), .ZN(n869bar);
  OR2_X1 U96 ( .A1(n866), .A2(n865), .ZN(n867) );
  AND2_X1 U96bar ( .A1(n866bar), .A2(n865bar), .ZN(n867bar);
  OR2_X1 U97 ( .A1(n864), .A2(n863), .ZN(n865) );
  AND2_X1 U97bar ( .A1(n864bar), .A2(n863bar), .ZN(n865bar);
  OR2_X1 U98 ( .A1(in[108]), .A2(n919), .ZN(n866) );
  AND2_X1 U98bar ( .A1(inbar[108]), .A2(n919bar), .ZN(n866bar);
  OR2_X1 U99 ( .A1(n862), .A2(n861), .ZN(n919) );
  AND2_X1 U99bar ( .A1(n862bar), .A2(n861bar), .ZN(n919bar);
  OR2_X1 U100 ( .A1(n860), .A2(n859), .ZN(n861) );
  AND2_X1 U100bar ( .A1(n860bar), .A2(n859bar), .ZN(n861bar);
  OR2_X1 U101 ( .A1(n858), .A2(n857), .ZN(n859) );
  AND2_X1 U101bar ( .A1(n858bar), .A2(n857bar), .ZN(n859bar);
  OR2_X1 U102 ( .A1(in[119]), .A2(in[105]), .ZN(n857) );
  AND2_X1 U102bar ( .A1(inbar[119]), .A2(inbar[105]), .ZN(n857bar);
  OR2_X1 U103 ( .A1(in[186]), .A2(in[175]), .ZN(n858) );
  AND2_X1 U103bar ( .A1(inbar[186]), .A2(inbar[175]), .ZN(n858bar);
  OR2_X1 U104 ( .A1(n856), .A2(n855), .ZN(n860) );
  AND2_X1 U104bar ( .A1(n856bar), .A2(n855bar), .ZN(n860bar);
  OR2_X1 U105 ( .A1(in[202]), .A2(in[193]), .ZN(n855) );
  AND2_X1 U105bar ( .A1(inbar[202]), .A2(inbar[193]), .ZN(n855bar);
  OR2_X1 U106 ( .A1(in[225]), .A2(in[208]), .ZN(n856) );
  AND2_X1 U106bar ( .A1(inbar[225]), .A2(inbar[208]), .ZN(n856bar);
  OR2_X1 U107 ( .A1(n854), .A2(n853), .ZN(n862) );
  AND2_X1 U107bar ( .A1(n854bar), .A2(n853bar), .ZN(n862bar);
  OR2_X1 U108 ( .A1(n852), .A2(n851), .ZN(n853) );
  AND2_X1 U108bar ( .A1(n852bar), .A2(n851bar), .ZN(n853bar);
  OR2_X1 U109 ( .A1(in_1), .A2(in[85]), .ZN(n851) );
  AND2_X1 U109bar ( .A1(in_1bar), .A2(inbar[85]), .ZN(n851bar);
  OR2_X1 U110 ( .A1(in_23), .A2(in_19), .ZN(n852) );
  AND2_X1 U110bar ( .A1(in_23bar), .A2(in_19bar), .ZN(n852bar);
  OR2_X1 U111 ( .A1(n850), .A2(n849), .ZN(n854) );
  AND2_X1 U111bar ( .A1(n850bar), .A2(n849bar), .ZN(n854bar);
  OR2_X1 U112 ( .A1(in_43), .A2(in_33), .ZN(n849) );
  AND2_X1 U112bar ( .A1(in_43bar), .A2(in_33bar), .ZN(n849bar);
  OR2_X1 U113 ( .A1(in_63), .A2(in_44), .ZN(n850) );
  AND2_X1 U113bar ( .A1(in_63bar), .A2(in_44bar), .ZN(n850bar);
  OR2_X1 U114 ( .A1(n848), .A2(n847), .ZN(n868) );
  AND2_X1 U114bar ( .A1(n848bar), .A2(n847bar), .ZN(n868bar);
  OR2_X1 U115 ( .A1(in[141]), .A2(in[112]), .ZN(n847) );
  AND2_X1 U115bar ( .A1(inbar[141]), .A2(inbar[112]), .ZN(n847bar);
  OR2_X1 U116 ( .A1(in[147]), .A2(n846), .ZN(n848) );
  AND2_X1 U116bar ( .A1(inbar[147]), .A2(n846bar), .ZN(n848bar);
  OR2_X1 U117 ( .A1(in[181]), .A2(in[167]), .ZN(n846) );
  AND2_X1 U117bar ( .A1(inbar[181]), .A2(inbar[167]), .ZN(n846bar);
  OR2_X1 U118 ( .A1(n845), .A2(n844), .ZN(n870) );
  AND2_X1 U118bar ( .A1(n845bar), .A2(n844bar), .ZN(n870bar);
  OR2_X1 U119 ( .A1(n843), .A2(n842), .ZN(n844) );
  AND2_X1 U119bar ( .A1(n843bar), .A2(n842bar), .ZN(n844bar);
  OR2_X1 U120 ( .A1(in[229]), .A2(in[201]), .ZN(n842) );
  AND2_X1 U120bar ( .A1(inbar[229]), .A2(inbar[201]), .ZN(n842bar);
  OR2_X1 U121 ( .A1(in[237]), .A2(n841), .ZN(n843) );
  AND2_X1 U121bar ( .A1(inbar[237]), .A2(n841bar), .ZN(n843bar);
  OR2_X1 U122 ( .A1(in[94]), .A2(in[253]), .ZN(n841) );
  AND2_X1 U122bar ( .A1(inbar[94]), .A2(inbar[253]), .ZN(n841bar);
  OR2_X1 U123 ( .A1(n840), .A2(n839), .ZN(n845) );
  AND2_X1 U123bar ( .A1(n840bar), .A2(n839bar), .ZN(n845bar);
  OR2_X1 U124 ( .A1(in_21), .A2(in[96]), .ZN(n839) );
  AND2_X1 U124bar ( .A1(in_21bar), .A2(inbar[96]), .ZN(n839bar);
  OR2_X1 U125 ( .A1(in_25), .A2(n838), .ZN(n840) );
  AND2_X1 U125bar ( .A1(in_25bar), .A2(n838bar), .ZN(n840bar);
  OR2_X1 U126 ( .A1(in_81), .A2(in_45), .ZN(n838) );
  AND2_X1 U126bar ( .A1(in_81bar), .A2(in_45bar), .ZN(n838bar);
  OR2_X1 U127 ( .A1(n837), .A2(n836), .ZN(n891) );
  AND2_X1 U127bar ( .A1(n837bar), .A2(n836bar), .ZN(n891bar);
  OR2_X1 U128 ( .A1(in[142]), .A2(in[124]), .ZN(n836) );
  AND2_X1 U128bar ( .A1(inbar[142]), .A2(inbar[124]), .ZN(n836bar);
  OR2_X1 U129 ( .A1(in[150]), .A2(n835), .ZN(n837) );
  AND2_X1 U129bar ( .A1(inbar[150]), .A2(n835bar), .ZN(n837bar);
  OR2_X1 U130 ( .A1(in[172]), .A2(in[155]), .ZN(n835) );
  AND2_X1 U130bar ( .A1(inbar[172]), .A2(inbar[155]), .ZN(n835bar);
  OR2_X1 U131 ( .A1(n834), .A2(n833), .ZN(n893) );
  AND2_X1 U131bar ( .A1(n834bar), .A2(n833bar), .ZN(n893bar);
  OR2_X1 U132 ( .A1(n832), .A2(n831), .ZN(n833) );
  AND2_X1 U132bar ( .A1(n832bar), .A2(n831bar), .ZN(n833bar);
  OR2_X1 U133 ( .A1(in[196]), .A2(in[173]), .ZN(n831) );
  AND2_X1 U133bar ( .A1(inbar[196]), .A2(inbar[173]), .ZN(n831bar);
  OR2_X1 U134 ( .A1(in[222]), .A2(n830), .ZN(n832) );
  AND2_X1 U134bar ( .A1(inbar[222]), .A2(n830bar), .ZN(n832bar);
  OR2_X1 U135 ( .A1(in[227]), .A2(in[226]), .ZN(n830) );
  AND2_X1 U135bar ( .A1(inbar[227]), .A2(inbar[226]), .ZN(n830bar);
  OR2_X1 U136 ( .A1(n829), .A2(n828), .ZN(n834) );
  AND2_X1 U136bar ( .A1(n829bar), .A2(n828bar), .ZN(n834bar);
  OR2_X1 U137 ( .A1(in[249]), .A2(in[231]), .ZN(n828) );
  AND2_X1 U137bar ( .A1(inbar[249]), .A2(inbar[231]), .ZN(n828bar);
  OR2_X1 U138 ( .A1(in_28), .A2(n827), .ZN(n829) );
  AND2_X1 U138bar ( .A1(in_28bar), .A2(n827bar), .ZN(n829bar);
  OR2_X1 U139 ( .A1(in_52), .A2(in_47), .ZN(n827) );
  AND2_X1 U139bar ( .A1(in_52bar), .A2(in_47bar), .ZN(n827bar);
  OR2_X1 U140 ( .A1(n826), .A2(n825), .ZN(out[3]) );
  AND2_X1 U140bar ( .A1(n826bar), .A2(n825bar), .ZN(outbar[3]);
  OR2_X1 U141 ( .A1(n824), .A2(n823), .ZN(n825) );
  AND2_X1 U141bar ( .A1(n824bar), .A2(n823bar), .ZN(n825bar);
  OR2_X1 U142 ( .A1(n822), .A2(n821), .ZN(n823) );
  AND2_X1 U142bar ( .A1(n822bar), .A2(n821bar), .ZN(n823bar);
  OR2_X1 U143 ( .A1(n820), .A2(n819), .ZN(n821) );
  AND2_X1 U143bar ( .A1(n820bar), .A2(n819bar), .ZN(n821bar);
  OR2_X1 U144 ( .A1(n964), .A2(n818), .ZN(n822) );
  AND2_X1 U144bar ( .A1(n964bar), .A2(n818bar), .ZN(n822bar);
  OR2_X1 U145 ( .A1(in[118]), .A2(n817), .ZN(n818) );
  AND2_X1 U145bar ( .A1(inbar[118]), .A2(n817bar), .ZN(n818bar);
  OR2_X1 U146 ( .A1(n816), .A2(n815), .ZN(n964) );
  AND2_X1 U146bar ( .A1(n816bar), .A2(n815bar), .ZN(n964bar);
  OR2_X1 U147 ( .A1(n814), .A2(n813), .ZN(n815) );
  AND2_X1 U147bar ( .A1(n814bar), .A2(n813bar), .ZN(n815bar);
  OR2_X1 U148 ( .A1(n812), .A2(n811), .ZN(n813) );
  AND2_X1 U148bar ( .A1(n812bar), .A2(n811bar), .ZN(n813bar);
  OR2_X1 U149 ( .A1(in[122]), .A2(in[111]), .ZN(n811) );
  AND2_X1 U149bar ( .A1(inbar[122]), .A2(inbar[111]), .ZN(n811bar);
  OR2_X1 U150 ( .A1(in[154]), .A2(in[151]), .ZN(n812) );
  AND2_X1 U150bar ( .A1(inbar[154]), .A2(inbar[151]), .ZN(n812bar);
  OR2_X1 U151 ( .A1(n810), .A2(n809), .ZN(n814) );
  AND2_X1 U151bar ( .A1(n810bar), .A2(n809bar), .ZN(n814bar);
  OR2_X1 U152 ( .A1(in[187]), .A2(in[177]), .ZN(n809) );
  AND2_X1 U152bar ( .A1(inbar[187]), .A2(inbar[177]), .ZN(n809bar);
  OR2_X1 U153 ( .A1(in[200]), .A2(in[192]), .ZN(n810) );
  AND2_X1 U153bar ( .A1(inbar[200]), .A2(inbar[192]), .ZN(n810bar);
  OR2_X1 U154 ( .A1(n808), .A2(n807), .ZN(n816) );
  AND2_X1 U154bar ( .A1(n808bar), .A2(n807bar), .ZN(n816bar);
  OR2_X1 U155 ( .A1(n806), .A2(n805), .ZN(n807) );
  AND2_X1 U155bar ( .A1(n806bar), .A2(n805bar), .ZN(n807bar);
  OR2_X1 U156 ( .A1(in[225]), .A2(in[207]), .ZN(n805) );
  AND2_X1 U156bar ( .A1(inbar[225]), .A2(inbar[207]), .ZN(n805bar);
  OR2_X1 U157 ( .A1(in[98]), .A2(in[226]), .ZN(n806) );
  AND2_X1 U157bar ( .A1(inbar[98]), .A2(inbar[226]), .ZN(n806bar);
  OR2_X1 U158 ( .A1(n804), .A2(n803), .ZN(n808) );
  AND2_X1 U158bar ( .A1(n804bar), .A2(n803bar), .ZN(n808bar);
  OR2_X1 U159 ( .A1(in_20), .A2(in_16), .ZN(n803) );
  AND2_X1 U159bar ( .A1(in_20bar), .A2(in_16bar), .ZN(n803bar);
  OR2_X1 U160 ( .A1(in_55), .A2(in_45), .ZN(n804) );
  AND2_X1 U160bar ( .A1(in_55bar), .A2(in_45bar), .ZN(n804bar);
  OR2_X1 U161 ( .A1(n802), .A2(n801), .ZN(n824) );
  AND2_X1 U161bar ( .A1(n802bar), .A2(n801bar), .ZN(n824bar);
  OR2_X1 U162 ( .A1(in[162]), .A2(in[149]), .ZN(n801) );
  AND2_X1 U162bar ( .A1(inbar[162]), .A2(inbar[149]), .ZN(n801bar);
  OR2_X1 U163 ( .A1(in[163]), .A2(n800), .ZN(n802) );
  AND2_X1 U163bar ( .A1(inbar[163]), .A2(n800bar), .ZN(n802bar);
  OR2_X1 U164 ( .A1(in[191]), .A2(in[189]), .ZN(n800) );
  AND2_X1 U164bar ( .A1(inbar[191]), .A2(inbar[189]), .ZN(n800bar);
  OR2_X1 U165 ( .A1(n799), .A2(n798), .ZN(n826) );
  AND2_X1 U165bar ( .A1(n799bar), .A2(n798bar), .ZN(n826bar);
  OR2_X1 U166 ( .A1(n797), .A2(n796), .ZN(n798) );
  AND2_X1 U166bar ( .A1(n797bar), .A2(n796bar), .ZN(n798bar);
  OR2_X1 U167 ( .A1(in[212]), .A2(in[193]), .ZN(n796) );
  AND2_X1 U167bar ( .A1(inbar[212]), .A2(inbar[193]), .ZN(n796bar);
  OR2_X1 U168 ( .A1(in[238]), .A2(n795), .ZN(n797) );
  AND2_X1 U168bar ( .A1(inbar[238]), .A2(n795bar), .ZN(n797bar);
  OR2_X1 U169 ( .A1(in[88]), .A2(in[247]), .ZN(n795) );
  AND2_X1 U169bar ( .A1(inbar[88]), .A2(inbar[247]), .ZN(n795bar);
  OR2_X1 U170 ( .A1(n794), .A2(n793), .ZN(n799) );
  AND2_X1 U170bar ( .A1(n794bar), .A2(n793bar), .ZN(n799bar);
  OR2_X1 U171 ( .A1(in[94]), .A2(in[92]), .ZN(n793) );
  AND2_X1 U171bar ( .A1(inbar[94]), .A2(inbar[92]), .ZN(n793bar);
  OR2_X1 U172 ( .A1(in_52), .A2(n792), .ZN(n794) );
  AND2_X1 U172bar ( .A1(in_52bar), .A2(n792bar), .ZN(n794bar);
  OR2_X1 U173 ( .A1(in_70), .A2(in_67), .ZN(n792) );
  AND2_X1 U173bar ( .A1(in_70bar), .A2(in_67bar), .ZN(n792bar);
  OR2_X1 U174 ( .A1(n791), .A2(n790), .ZN(out[2]) );
  AND2_X1 U174bar ( .A1(n791bar), .A2(n790bar), .ZN(outbar[2]);
  OR2_X1 U175 ( .A1(n789), .A2(n788), .ZN(n790) );
  AND2_X1 U175bar ( .A1(n789bar), .A2(n788bar), .ZN(n790bar);
  OR2_X1 U176 ( .A1(n787), .A2(n786), .ZN(n788) );
  AND2_X1 U176bar ( .A1(n787bar), .A2(n786bar), .ZN(n788bar);
  OR2_X1 U177 ( .A1(n819), .A2(n785), .ZN(n786) );
  AND2_X1 U177bar ( .A1(n819bar), .A2(n785bar), .ZN(n786bar);
  OR2_X1 U178 ( .A1(n784), .A2(n783), .ZN(n819) );
  AND2_X1 U178bar ( .A1(n784bar), .A2(n783bar), .ZN(n819bar);
  OR2_X1 U179 ( .A1(n782), .A2(n781), .ZN(n783) );
  AND2_X1 U179bar ( .A1(n782bar), .A2(n781bar), .ZN(n783bar);
  OR2_X1 U180 ( .A1(n780), .A2(n779), .ZN(n781) );
  AND2_X1 U180bar ( .A1(n780bar), .A2(n779bar), .ZN(n781bar);
  OR2_X1 U181 ( .A1(n962), .A2(n778), .ZN(n779) );
  AND2_X1 U181bar ( .A1(n962bar), .A2(n778bar), .ZN(n779bar);
  OR2_X1 U182 ( .A1(n777), .A2(n776), .ZN(n962) );
  AND2_X1 U182bar ( .A1(n777bar), .A2(n776bar), .ZN(n962bar);
  OR2_X1 U183 ( .A1(n775), .A2(n774), .ZN(n776) );
  AND2_X1 U183bar ( .A1(n775bar), .A2(n774bar), .ZN(n776bar);
  OR2_X1 U184 ( .A1(n773), .A2(n772), .ZN(n774) );
  AND2_X1 U184bar ( .A1(n773bar), .A2(n772bar), .ZN(n774bar);
  OR2_X1 U185 ( .A1(in[131]), .A2(in[120]), .ZN(n772) );
  AND2_X1 U185bar ( .A1(inbar[131]), .A2(inbar[120]), .ZN(n772bar);
  OR2_X1 U186 ( .A1(in[153]), .A2(in[147]), .ZN(n773) );
  AND2_X1 U186bar ( .A1(inbar[153]), .A2(inbar[147]), .ZN(n773bar);
  OR2_X1 U187 ( .A1(n771), .A2(n770), .ZN(n775) );
  AND2_X1 U187bar ( .A1(n771bar), .A2(n770bar), .ZN(n775bar);
  OR2_X1 U188 ( .A1(in[170]), .A2(in[156]), .ZN(n770) );
  AND2_X1 U188bar ( .A1(inbar[170]), .A2(inbar[156]), .ZN(n770bar);
  OR2_X1 U189 ( .A1(in[223]), .A2(in[190]), .ZN(n771) );
  AND2_X1 U189bar ( .A1(inbar[223]), .A2(inbar[190]), .ZN(n771bar);
  OR2_X1 U190 ( .A1(n769), .A2(n768), .ZN(n777) );
  AND2_X1 U190bar ( .A1(n769bar), .A2(n768bar), .ZN(n777bar);
  OR2_X1 U191 ( .A1(n767), .A2(n766), .ZN(n768) );
  AND2_X1 U191bar ( .A1(n767bar), .A2(n766bar), .ZN(n768bar);
  OR2_X1 U192 ( .A1(in[236]), .A2(in[230]), .ZN(n766) );
  AND2_X1 U192bar ( .A1(inbar[236]), .A2(inbar[230]), .ZN(n766bar);
  OR2_X1 U193 ( .A1(in[85]), .A2(in[240]), .ZN(n767) );
  AND2_X1 U193bar ( .A1(inbar[85]), .A2(inbar[240]), .ZN(n767bar);
  OR2_X1 U194 ( .A1(n765), .A2(n764), .ZN(n769) );
  AND2_X1 U194bar ( .A1(n765bar), .A2(n764bar), .ZN(n769bar);
  OR2_X1 U195 ( .A1(in_12), .A2(in[90]), .ZN(n764) );
  AND2_X1 U195bar ( .A1(in_12bar), .A2(inbar[90]), .ZN(n764bar);
  OR2_X1 U196 ( .A1(in_39), .A2(in_28), .ZN(n765) );
  AND2_X1 U196bar ( .A1(in_39bar), .A2(in_28bar), .ZN(n765bar);
  OR2_X1 U197 ( .A1(in[109]), .A2(n763), .ZN(n780) );
  AND2_X1 U197bar ( .A1(inbar[109]), .A2(n763bar), .ZN(n780bar);
  OR2_X1 U198 ( .A1(n762), .A2(n761), .ZN(n782) );
  AND2_X1 U198bar ( .A1(n762bar), .A2(n761bar), .ZN(n782bar);
  OR2_X1 U199 ( .A1(in[138]), .A2(in[129]), .ZN(n761) );
  AND2_X1 U199bar ( .A1(inbar[138]), .A2(inbar[129]), .ZN(n761bar);
  OR2_X1 U200 ( .A1(in[157]), .A2(n760), .ZN(n762) );
  AND2_X1 U200bar ( .A1(inbar[157]), .A2(n760bar), .ZN(n762bar);
  OR2_X1 U201 ( .A1(in[182]), .A2(in[167]), .ZN(n760) );
  AND2_X1 U201bar ( .A1(inbar[182]), .A2(inbar[167]), .ZN(n760bar);
  OR2_X1 U202 ( .A1(n759), .A2(n758), .ZN(n784) );
  AND2_X1 U202bar ( .A1(n759bar), .A2(n758bar), .ZN(n784bar);
  OR2_X1 U203 ( .A1(n757), .A2(n756), .ZN(n758) );
  AND2_X1 U203bar ( .A1(n757bar), .A2(n756bar), .ZN(n758bar);
  OR2_X1 U204 ( .A1(in[195]), .A2(in[184]), .ZN(n756) );
  AND2_X1 U204bar ( .A1(inbar[195]), .A2(inbar[184]), .ZN(n756bar);
  OR2_X1 U205 ( .A1(in[196]), .A2(n755), .ZN(n757) );
  AND2_X1 U205bar ( .A1(inbar[196]), .A2(n755bar), .ZN(n757bar);
  OR2_X1 U206 ( .A1(in[215]), .A2(in[209]), .ZN(n755) );
  AND2_X1 U206bar ( .A1(inbar[215]), .A2(inbar[209]), .ZN(n755bar);
  OR2_X1 U207 ( .A1(n754), .A2(n753), .ZN(n759) );
  AND2_X1 U207bar ( .A1(n754bar), .A2(n753bar), .ZN(n759bar);
  OR2_X1 U208 ( .A1(in[93]), .A2(in[233]), .ZN(n753) );
  AND2_X1 U208bar ( .A1(inbar[93]), .A2(inbar[233]), .ZN(n753bar);
  OR2_X1 U209 ( .A1(in_1), .A2(n752), .ZN(n754) );
  AND2_X1 U209bar ( .A1(in_1bar), .A2(n752bar), .ZN(n754bar);
  OR2_X1 U210 ( .A1(in_69), .A2(in_66), .ZN(n752) );
  AND2_X1 U210bar ( .A1(in_69bar), .A2(in_66bar), .ZN(n752bar);
  OR2_X1 U211 ( .A1(n966), .A2(n751), .ZN(n787) );
  AND2_X1 U211bar ( .A1(n966bar), .A2(n751bar), .ZN(n787bar);
  OR2_X1 U212 ( .A1(in[134]), .A2(n750), .ZN(n751) );
  AND2_X1 U212bar ( .A1(inbar[134]), .A2(n750bar), .ZN(n751bar);
  OR2_X1 U213 ( .A1(n749), .A2(n748), .ZN(n966) );
  AND2_X1 U213bar ( .A1(n749bar), .A2(n748bar), .ZN(n966bar);
  OR2_X1 U214 ( .A1(n747), .A2(n746), .ZN(n748) );
  AND2_X1 U214bar ( .A1(n747bar), .A2(n746bar), .ZN(n748bar);
  OR2_X1 U215 ( .A1(n745), .A2(n744), .ZN(n746) );
  AND2_X1 U215bar ( .A1(n745bar), .A2(n744bar), .ZN(n746bar);
  OR2_X1 U216 ( .A1(in[136]), .A2(in[121]), .ZN(n744) );
  AND2_X1 U216bar ( .A1(inbar[136]), .A2(inbar[121]), .ZN(n744bar);
  OR2_X1 U217 ( .A1(in[186]), .A2(in[174]), .ZN(n745) );
  AND2_X1 U217bar ( .A1(inbar[186]), .A2(inbar[174]), .ZN(n745bar);
  OR2_X1 U218 ( .A1(n743), .A2(n742), .ZN(n747) );
  AND2_X1 U218bar ( .A1(n743bar), .A2(n742bar), .ZN(n747bar);
  OR2_X1 U219 ( .A1(in[198]), .A2(in[197]), .ZN(n742) );
  AND2_X1 U219bar ( .A1(inbar[198]), .A2(inbar[197]), .ZN(n742bar);
  OR2_X1 U220 ( .A1(in[214]), .A2(in[199]), .ZN(n743) );
  AND2_X1 U220bar ( .A1(inbar[214]), .A2(inbar[199]), .ZN(n743bar);
  OR2_X1 U221 ( .A1(n741), .A2(n740), .ZN(n749) );
  AND2_X1 U221bar ( .A1(n741bar), .A2(n740bar), .ZN(n749bar);
  OR2_X1 U222 ( .A1(n739), .A2(n738), .ZN(n740) );
  AND2_X1 U222bar ( .A1(n739bar), .A2(n738bar), .ZN(n740bar);
  OR2_X1 U223 ( .A1(in[231]), .A2(in[220]), .ZN(n738) );
  AND2_X1 U223bar ( .A1(inbar[231]), .A2(inbar[220]), .ZN(n738bar);
  OR2_X1 U224 ( .A1(in_25), .A2(in[245]), .ZN(n739) );
  AND2_X1 U224bar ( .A1(in_25bar), .A2(inbar[245]), .ZN(n739bar);
  OR2_X1 U225 ( .A1(n737), .A2(n736), .ZN(n741) );
  AND2_X1 U225bar ( .A1(n737bar), .A2(n736bar), .ZN(n741bar);
  OR2_X1 U226 ( .A1(in_53), .A2(in_29), .ZN(n736) );
  AND2_X1 U226bar ( .A1(in_53bar), .A2(in_29bar), .ZN(n736bar);
  OR2_X1 U227 ( .A1(in_79), .A2(in_74), .ZN(n737) );
  AND2_X1 U227bar ( .A1(in_79bar), .A2(in_74bar), .ZN(n737bar);
  OR2_X1 U228 ( .A1(n735), .A2(n734), .ZN(n789) );
  AND2_X1 U228bar ( .A1(n735bar), .A2(n734bar), .ZN(n789bar);
  OR2_X1 U229 ( .A1(in[152]), .A2(in[140]), .ZN(n734) );
  AND2_X1 U229bar ( .A1(inbar[152]), .A2(inbar[140]), .ZN(n734bar);
  OR2_X1 U230 ( .A1(in[155]), .A2(n733), .ZN(n735) );
  AND2_X1 U230bar ( .A1(inbar[155]), .A2(n733bar), .ZN(n735bar);
  OR2_X1 U231 ( .A1(in[166]), .A2(in[165]), .ZN(n733) );
  AND2_X1 U231bar ( .A1(inbar[166]), .A2(inbar[165]), .ZN(n733bar);
  OR2_X1 U232 ( .A1(n732), .A2(n731), .ZN(n791) );
  AND2_X1 U232bar ( .A1(n732bar), .A2(n731bar), .ZN(n791bar);
  OR2_X1 U233 ( .A1(n730), .A2(n729), .ZN(n731) );
  AND2_X1 U233bar ( .A1(n730bar), .A2(n729bar), .ZN(n731bar);
  OR2_X1 U234 ( .A1(in[202]), .A2(in[185]), .ZN(n729) );
  AND2_X1 U234bar ( .A1(inbar[202]), .A2(inbar[185]), .ZN(n729bar);
  OR2_X1 U235 ( .A1(in[211]), .A2(n728), .ZN(n730) );
  AND2_X1 U235bar ( .A1(inbar[211]), .A2(n728bar), .ZN(n730bar);
  OR2_X1 U236 ( .A1(in[255]), .A2(in[253]), .ZN(n728) );
  AND2_X1 U236bar ( .A1(inbar[255]), .A2(inbar[253]), .ZN(n728bar);
  OR2_X1 U237 ( .A1(n727), .A2(n726), .ZN(n732) );
  AND2_X1 U237bar ( .A1(n727bar), .A2(n726bar), .ZN(n732bar);
  OR2_X1 U238 ( .A1(in_35), .A2(in_15), .ZN(n726) );
  AND2_X1 U238bar ( .A1(in_35bar), .A2(in_15bar), .ZN(n726bar);
  OR2_X1 U239 ( .A1(in_36), .A2(n725), .ZN(n727) );
  AND2_X1 U239bar ( .A1(in_36bar), .A2(n725bar), .ZN(n727bar);
  OR2_X1 U240 ( .A1(in_48), .A2(in_40), .ZN(n725) );
  AND2_X1 U240bar ( .A1(in_48bar), .A2(in_40bar), .ZN(n725bar);
  OR2_X1 U241 ( .A1(n724), .A2(n723), .ZN(out[1]) );
  AND2_X1 U241bar ( .A1(n724bar), .A2(n723bar), .ZN(outbar[1]);
  OR2_X1 U242 ( .A1(n722), .A2(n721), .ZN(n723) );
  AND2_X1 U242bar ( .A1(n722bar), .A2(n721bar), .ZN(n723bar);
  OR2_X1 U243 ( .A1(n720), .A2(n719), .ZN(n721) );
  AND2_X1 U243bar ( .A1(n720bar), .A2(n719bar), .ZN(n721bar);
  OR2_X1 U244 ( .A1(n921), .A2(n887), .ZN(n719) );
  AND2_X1 U244bar ( .A1(n921bar), .A2(n887bar), .ZN(n719bar);
  OR2_X1 U245 ( .A1(n718), .A2(n717), .ZN(n887) );
  AND2_X1 U245bar ( .A1(n718bar), .A2(n717bar), .ZN(n887bar);
  OR2_X1 U246 ( .A1(n716), .A2(n715), .ZN(n717) );
  AND2_X1 U246bar ( .A1(n716bar), .A2(n715bar), .ZN(n717bar);
  OR2_X1 U247 ( .A1(n714), .A2(n713), .ZN(n715) );
  AND2_X1 U247bar ( .A1(n714bar), .A2(n713bar), .ZN(n715bar);
  OR2_X1 U248 ( .A1(in[116]), .A2(in[110]), .ZN(n713) );
  AND2_X1 U248bar ( .A1(inbar[116]), .A2(inbar[110]), .ZN(n713bar);
  OR2_X1 U249 ( .A1(in[133]), .A2(in[130]), .ZN(n714) );
  AND2_X1 U249bar ( .A1(inbar[133]), .A2(inbar[130]), .ZN(n714bar);
  OR2_X1 U250 ( .A1(n712), .A2(n711), .ZN(n716) );
  AND2_X1 U250bar ( .A1(n712bar), .A2(n711bar), .ZN(n716bar);
  OR2_X1 U251 ( .A1(in[203]), .A2(in[135]), .ZN(n711) );
  AND2_X1 U251bar ( .A1(inbar[203]), .A2(inbar[135]), .ZN(n711bar);
  OR2_X1 U252 ( .A1(in[232]), .A2(in[223]), .ZN(n712) );
  AND2_X1 U252bar ( .A1(inbar[232]), .A2(inbar[223]), .ZN(n712bar);
  OR2_X1 U253 ( .A1(n710), .A2(n709), .ZN(n718) );
  AND2_X1 U253bar ( .A1(n710bar), .A2(n709bar), .ZN(n718bar);
  OR2_X1 U254 ( .A1(n708), .A2(n707), .ZN(n709) );
  AND2_X1 U254bar ( .A1(n708bar), .A2(n707bar), .ZN(n709bar);
  OR2_X1 U255 ( .A1(in[255]), .A2(in[233]), .ZN(n707) );
  AND2_X1 U255bar ( .A1(inbar[255]), .A2(inbar[233]), .ZN(n707bar);
  OR2_X1 U256 ( .A1(in_53), .A2(in_34), .ZN(n708) );
  AND2_X1 U256bar ( .A1(in_53bar), .A2(in_34bar), .ZN(n708bar);
  OR2_X1 U257 ( .A1(n706), .A2(n705), .ZN(n710) );
  AND2_X1 U257bar ( .A1(n706bar), .A2(n705bar), .ZN(n710bar);
  OR2_X1 U258 ( .A1(in_57), .A2(in_55), .ZN(n705) );
  AND2_X1 U258bar ( .A1(in_57bar), .A2(in_55bar), .ZN(n705bar);
  OR2_X1 U259 ( .A1(in_68), .A2(in_67), .ZN(n706) );
  AND2_X1 U259bar ( .A1(in_68bar), .A2(in_67bar), .ZN(n706bar);
  OR2_X1 U260 ( .A1(n704), .A2(n703), .ZN(n921) );
  AND2_X1 U260bar ( .A1(n704bar), .A2(n703bar), .ZN(n921bar);
  OR2_X1 U261 ( .A1(n702), .A2(n701), .ZN(n703) );
  AND2_X1 U261bar ( .A1(n702bar), .A2(n701bar), .ZN(n703bar);
  OR2_X1 U262 ( .A1(n700), .A2(n699), .ZN(n701) );
  AND2_X1 U262bar ( .A1(n700bar), .A2(n699bar), .ZN(n701bar);
  OR2_X1 U263 ( .A1(n944), .A2(n872), .ZN(n699) );
  AND2_X1 U263bar ( .A1(n944bar), .A2(n872bar), .ZN(n699bar);
  OR2_X1 U264 ( .A1(n698), .A2(n697), .ZN(n872) );
  AND2_X1 U264bar ( .A1(n698bar), .A2(n697bar), .ZN(n872bar);
  OR2_X1 U265 ( .A1(n696), .A2(n695), .ZN(n697) );
  AND2_X1 U265bar ( .A1(n696bar), .A2(n695bar), .ZN(n697bar);
  OR2_X1 U266 ( .A1(n694), .A2(n693), .ZN(n695) );
  AND2_X1 U266bar ( .A1(n694bar), .A2(n693bar), .ZN(n695bar);
  OR2_X1 U267 ( .A1(in[121]), .A2(in[102]), .ZN(n693) );
  AND2_X1 U267bar ( .A1(inbar[121]), .A2(inbar[102]), .ZN(n693bar);
  OR2_X1 U268 ( .A1(in[162]), .A2(in[161]), .ZN(n694) );
  AND2_X1 U268bar ( .A1(inbar[162]), .A2(inbar[161]), .ZN(n694bar);
  OR2_X1 U269 ( .A1(n692), .A2(n691), .ZN(n696) );
  AND2_X1 U269bar ( .A1(n692bar), .A2(n691bar), .ZN(n696bar);
  OR2_X1 U270 ( .A1(in[192]), .A2(in[178]), .ZN(n691) );
  AND2_X1 U270bar ( .A1(inbar[192]), .A2(inbar[178]), .ZN(n691bar);
  OR2_X1 U271 ( .A1(in[244]), .A2(in[209]), .ZN(n692) );
  AND2_X1 U271bar ( .A1(inbar[244]), .A2(inbar[209]), .ZN(n692bar);
  OR2_X1 U272 ( .A1(n690), .A2(n689), .ZN(n698) );
  AND2_X1 U272bar ( .A1(n690bar), .A2(n689bar), .ZN(n698bar);
  OR2_X1 U273 ( .A1(n688), .A2(n687), .ZN(n689) );
  AND2_X1 U273bar ( .A1(n688bar), .A2(n687bar), .ZN(n689bar);
  OR2_X1 U274 ( .A1(in[90]), .A2(in[254]), .ZN(n687) );
  AND2_X1 U274bar ( .A1(inbar[90]), .A2(inbar[254]), .ZN(n687bar);
  OR2_X1 U275 ( .A1(in_36), .A2(in_32), .ZN(n688) );
  AND2_X1 U275bar ( .A1(in_36bar), .A2(in_32bar), .ZN(n688bar);
  OR2_X1 U276 ( .A1(n686), .A2(n685), .ZN(n690) );
  AND2_X1 U276bar ( .A1(n686bar), .A2(n685bar), .ZN(n690bar);
  OR2_X1 U277 ( .A1(in_62), .A2(in_37), .ZN(n685) );
  AND2_X1 U277bar ( .A1(in_62bar), .A2(in_37bar), .ZN(n685bar);
  OR2_X1 U278 ( .A1(in_75), .A2(in_73), .ZN(n686) );
  AND2_X1 U278bar ( .A1(in_75bar), .A2(in_73bar), .ZN(n686bar);
  OR2_X1 U279 ( .A1(n684), .A2(n683), .ZN(n944) );
  AND2_X1 U279bar ( .A1(n684bar), .A2(n683bar), .ZN(n944bar);
  OR2_X1 U280 ( .A1(n682), .A2(n681), .ZN(n683) );
  AND2_X1 U280bar ( .A1(n682bar), .A2(n681bar), .ZN(n683bar);
  OR2_X1 U281 ( .A1(n680), .A2(n679), .ZN(n681) );
  AND2_X1 U281bar ( .A1(n680bar), .A2(n679bar), .ZN(n681bar);
  OR2_X1 U282 ( .A1(in[171]), .A2(in[153]), .ZN(n679) );
  AND2_X1 U282bar ( .A1(inbar[171]), .A2(inbar[153]), .ZN(n679bar);
  OR2_X1 U283 ( .A1(in[187]), .A2(in[176]), .ZN(n680) );
  AND2_X1 U283bar ( .A1(inbar[187]), .A2(inbar[176]), .ZN(n680bar);
  OR2_X1 U284 ( .A1(n678), .A2(n677), .ZN(n682) );
  AND2_X1 U284bar ( .A1(n678bar), .A2(n677bar), .ZN(n682bar);
  OR2_X1 U285 ( .A1(in[245]), .A2(in[211]), .ZN(n677) );
  AND2_X1 U285bar ( .A1(inbar[245]), .A2(inbar[211]), .ZN(n677bar);
  OR2_X1 U286 ( .A1(in[97]), .A2(in[88]), .ZN(n678) );
  AND2_X1 U286bar ( .A1(inbar[97]), .A2(inbar[88]), .ZN(n678bar);
  OR2_X1 U287 ( .A1(n676), .A2(n675), .ZN(n684) );
  AND2_X1 U287bar ( .A1(n676bar), .A2(n675bar), .ZN(n684bar);
  OR2_X1 U288 ( .A1(n674), .A2(n673), .ZN(n675) );
  AND2_X1 U288bar ( .A1(n674bar), .A2(n673bar), .ZN(n675bar);
  OR2_X1 U289 ( .A1(in_10), .A2(in_0), .ZN(n673) );
  AND2_X1 U289bar ( .A1(in_10bar), .A2(in_0bar), .ZN(n673bar);
  OR2_X1 U290 ( .A1(in_59), .A2(in_5), .ZN(n674) );
  AND2_X1 U290bar ( .A1(in_59bar), .A2(in_5bar), .ZN(n674bar);
  OR2_X1 U291 ( .A1(n672), .A2(n671), .ZN(n676) );
  AND2_X1 U291bar ( .A1(n672bar), .A2(n671bar), .ZN(n676bar);
  OR2_X1 U292 ( .A1(in_60), .A2(in_6), .ZN(n671) );
  AND2_X1 U292bar ( .A1(in_60bar), .A2(in_6bar), .ZN(n671bar);
  OR2_X1 U293 ( .A1(in_77), .A2(in_69), .ZN(n672) );
  AND2_X1 U293bar ( .A1(in_77bar), .A2(in_69bar), .ZN(n672bar);
  OR2_X1 U294 ( .A1(in[113]), .A2(n864), .ZN(n700) );
  AND2_X1 U294bar ( .A1(inbar[113]), .A2(n864bar), .ZN(n700bar);
  OR2_X1 U295 ( .A1(n670), .A2(n669), .ZN(n864) );
  AND2_X1 U295bar ( .A1(n670bar), .A2(n669bar), .ZN(n864bar);
  OR2_X1 U296 ( .A1(n668), .A2(n667), .ZN(n669) );
  AND2_X1 U296bar ( .A1(n668bar), .A2(n667bar), .ZN(n669bar);
  OR2_X1 U297 ( .A1(n666), .A2(n665), .ZN(n667) );
  AND2_X1 U297bar ( .A1(n666bar), .A2(n665bar), .ZN(n667bar);
  OR2_X1 U298 ( .A1(in[125]), .A2(in[107]), .ZN(n665) );
  AND2_X1 U298bar ( .A1(inbar[125]), .A2(inbar[107]), .ZN(n665bar);
  OR2_X1 U299 ( .A1(in[138]), .A2(in[126]), .ZN(n666) );
  AND2_X1 U299bar ( .A1(inbar[138]), .A2(inbar[126]), .ZN(n666bar);
  OR2_X1 U300 ( .A1(n664), .A2(n663), .ZN(n668) );
  AND2_X1 U300bar ( .A1(n664bar), .A2(n663bar), .ZN(n668bar);
  OR2_X1 U301 ( .A1(in[189]), .A2(in[143]), .ZN(n663) );
  AND2_X1 U301bar ( .A1(inbar[189]), .A2(inbar[143]), .ZN(n663bar);
  OR2_X1 U302 ( .A1(in[99]), .A2(in[214]), .ZN(n664) );
  AND2_X1 U302bar ( .A1(inbar[99]), .A2(inbar[214]), .ZN(n664bar);
  OR2_X1 U303 ( .A1(n662), .A2(n661), .ZN(n670) );
  AND2_X1 U303bar ( .A1(n662bar), .A2(n661bar), .ZN(n670bar);
  OR2_X1 U304 ( .A1(n660), .A2(n659), .ZN(n661) );
  AND2_X1 U304bar ( .A1(n660bar), .A2(n659bar), .ZN(n661bar);
  OR2_X1 U305 ( .A1(in_15), .A2(in_12), .ZN(n659) );
  AND2_X1 U305bar ( .A1(in_15bar), .A2(in_12bar), .ZN(n659bar);
  OR2_X1 U306 ( .A1(in_20), .A2(in_2), .ZN(n660) );
  AND2_X1 U306bar ( .A1(in_20bar), .A2(in_2bar), .ZN(n660bar);
  OR2_X1 U307 ( .A1(n658), .A2(n657), .ZN(n662) );
  AND2_X1 U307bar ( .A1(n658bar), .A2(n657bar), .ZN(n662bar);
  OR2_X1 U308 ( .A1(in_30), .A2(in_3), .ZN(n657) );
  AND2_X1 U308bar ( .A1(in_30bar), .A2(in_3bar), .ZN(n657bar);
  OR2_X1 U309 ( .A1(in_4), .A2(in_38), .ZN(n658) );
  AND2_X1 U309bar ( .A1(in_4bar), .A2(in_38bar), .ZN(n658bar);
  OR2_X1 U310 ( .A1(n656), .A2(n655), .ZN(n702) );
  AND2_X1 U310bar ( .A1(n656bar), .A2(n655bar), .ZN(n702bar);
  OR2_X1 U311 ( .A1(in[148]), .A2(in[137]), .ZN(n655) );
  AND2_X1 U311bar ( .A1(inbar[148]), .A2(inbar[137]), .ZN(n655bar);
  OR2_X1 U312 ( .A1(in[149]), .A2(n654), .ZN(n656) );
  AND2_X1 U312bar ( .A1(inbar[149]), .A2(n654bar), .ZN(n656bar);
  OR2_X1 U313 ( .A1(in[195]), .A2(in[190]), .ZN(n654) );
  AND2_X1 U313bar ( .A1(inbar[195]), .A2(inbar[190]), .ZN(n654bar);
  OR2_X1 U314 ( .A1(n653), .A2(n652), .ZN(n704) );
  AND2_X1 U314bar ( .A1(n653bar), .A2(n652bar), .ZN(n704bar);
  OR2_X1 U315 ( .A1(n651), .A2(n650), .ZN(n652) );
  AND2_X1 U315bar ( .A1(n651bar), .A2(n650bar), .ZN(n652bar);
  OR2_X1 U316 ( .A1(in[98]), .A2(in[197]), .ZN(n650) );
  AND2_X1 U316bar ( .A1(inbar[98]), .A2(inbar[197]), .ZN(n650bar);
  OR2_X1 U317 ( .A1(in_11), .A2(n649), .ZN(n651) );
  AND2_X1 U317bar ( .A1(in_11bar), .A2(n649bar), .ZN(n651bar);
  OR2_X1 U318 ( .A1(in_26), .A2(in_14), .ZN(n649) );
  AND2_X1 U318bar ( .A1(in_26bar), .A2(in_14bar), .ZN(n649bar);
  OR2_X1 U319 ( .A1(n648), .A2(n647), .ZN(n653) );
  AND2_X1 U319bar ( .A1(n648bar), .A2(n647bar), .ZN(n653bar);
  OR2_X1 U320 ( .A1(in_35), .A2(in_27), .ZN(n647) );
  AND2_X1 U320bar ( .A1(in_35bar), .A2(in_27bar), .ZN(n647bar);
  OR2_X1 U321 ( .A1(in_50), .A2(n646), .ZN(n648) );
  AND2_X1 U321bar ( .A1(in_50bar), .A2(n646bar), .ZN(n648bar);
  OR2_X1 U322 ( .A1(in_78), .A2(in_61), .ZN(n646) );
  AND2_X1 U322bar ( .A1(in_78bar), .A2(in_61bar), .ZN(n646bar);
  OR2_X1 U323 ( .A1(n942), .A2(n645), .ZN(n720) );
  AND2_X1 U323bar ( .A1(n942bar), .A2(n645bar), .ZN(n720bar);
  OR2_X1 U324 ( .A1(in[106]), .A2(n863), .ZN(n645) );
  AND2_X1 U324bar ( .A1(inbar[106]), .A2(n863bar), .ZN(n645bar);
  OR2_X1 U325 ( .A1(n644), .A2(n643), .ZN(n863) );
  AND2_X1 U325bar ( .A1(n644bar), .A2(n643bar), .ZN(n863bar);
  OR2_X1 U326 ( .A1(n642), .A2(n641), .ZN(n643) );
  AND2_X1 U326bar ( .A1(n642bar), .A2(n641bar), .ZN(n643bar);
  OR2_X1 U327 ( .A1(n640), .A2(n639), .ZN(n641) );
  AND2_X1 U327bar ( .A1(n640bar), .A2(n639bar), .ZN(n641bar);
  OR2_X1 U328 ( .A1(in[127]), .A2(in[122]), .ZN(n639) );
  AND2_X1 U328bar ( .A1(inbar[127]), .A2(inbar[122]), .ZN(n639bar);
  OR2_X1 U329 ( .A1(in[156]), .A2(in[132]), .ZN(n640) );
  AND2_X1 U329bar ( .A1(inbar[156]), .A2(inbar[132]), .ZN(n640bar);
  OR2_X1 U330 ( .A1(n638), .A2(n637), .ZN(n642) );
  AND2_X1 U330bar ( .A1(n638bar), .A2(n637bar), .ZN(n642bar);
  OR2_X1 U331 ( .A1(in[159]), .A2(in[157]), .ZN(n637) );
  AND2_X1 U331bar ( .A1(inbar[159]), .A2(inbar[157]), .ZN(n637bar);
  OR2_X1 U332 ( .A1(in[185]), .A2(in[169]), .ZN(n638) );
  AND2_X1 U332bar ( .A1(inbar[185]), .A2(inbar[169]), .ZN(n638bar);
  OR2_X1 U333 ( .A1(n636), .A2(n635), .ZN(n644) );
  AND2_X1 U333bar ( .A1(n636bar), .A2(n635bar), .ZN(n644bar);
  OR2_X1 U334 ( .A1(n634), .A2(n633), .ZN(n635) );
  AND2_X1 U334bar ( .A1(n634bar), .A2(n633bar), .ZN(n635bar);
  OR2_X1 U335 ( .A1(in[239]), .A2(in[218]), .ZN(n633) );
  AND2_X1 U335bar ( .A1(inbar[239]), .A2(inbar[218]), .ZN(n633bar);
  OR2_X1 U336 ( .A1(in_13), .A2(in[87]), .ZN(n634) );
  AND2_X1 U336bar ( .A1(in_13bar), .A2(inbar[87]), .ZN(n634bar);
  OR2_X1 U337 ( .A1(n632), .A2(n631), .ZN(n636) );
  AND2_X1 U337bar ( .A1(n632bar), .A2(n631bar), .ZN(n636bar);
  OR2_X1 U338 ( .A1(in_72), .A2(in_70), .ZN(n631) );
  AND2_X1 U338bar ( .A1(in_72bar), .A2(in_70bar), .ZN(n631bar);
  OR2_X1 U339 ( .A1(in_80), .A2(in_74), .ZN(n632) );
  AND2_X1 U339bar ( .A1(in_80bar), .A2(in_74bar), .ZN(n632bar);
  OR2_X1 U340 ( .A1(n630), .A2(n629), .ZN(n942) );
  AND2_X1 U340bar ( .A1(n630bar), .A2(n629bar), .ZN(n942bar);
  OR2_X1 U341 ( .A1(n628), .A2(n627), .ZN(n629) );
  AND2_X1 U341bar ( .A1(n628bar), .A2(n627bar), .ZN(n629bar);
  OR2_X1 U342 ( .A1(n626), .A2(n625), .ZN(n627) );
  AND2_X1 U342bar ( .A1(n626bar), .A2(n625bar), .ZN(n627bar);
  OR2_X1 U343 ( .A1(in[146]), .A2(in[100]), .ZN(n625) );
  AND2_X1 U343bar ( .A1(inbar[146]), .A2(inbar[100]), .ZN(n625bar);
  OR2_X1 U344 ( .A1(in[168]), .A2(in[152]), .ZN(n626) );
  AND2_X1 U344bar ( .A1(inbar[168]), .A2(inbar[152]), .ZN(n626bar);
  OR2_X1 U345 ( .A1(n624), .A2(n623), .ZN(n628) );
  AND2_X1 U345bar ( .A1(n624bar), .A2(n623bar), .ZN(n628bar);
  OR2_X1 U346 ( .A1(in[199]), .A2(in[182]), .ZN(n623) );
  AND2_X1 U346bar ( .A1(inbar[199]), .A2(inbar[182]), .ZN(n623bar);
  OR2_X1 U347 ( .A1(in[236]), .A2(in[204]), .ZN(n624) );
  AND2_X1 U347bar ( .A1(inbar[236]), .A2(inbar[204]), .ZN(n624bar);
  OR2_X1 U348 ( .A1(n622), .A2(n621), .ZN(n630) );
  AND2_X1 U348bar ( .A1(n622bar), .A2(n621bar), .ZN(n630bar);
  OR2_X1 U349 ( .A1(n620), .A2(n619), .ZN(n621) );
  AND2_X1 U349bar ( .A1(n620bar), .A2(n619bar), .ZN(n621bar);
  OR2_X1 U350 ( .A1(in[89]), .A2(in[246]), .ZN(n619) );
  AND2_X1 U350bar ( .A1(inbar[89]), .A2(inbar[246]), .ZN(n619bar);
  OR2_X1 U351 ( .A1(in[95]), .A2(in[92]), .ZN(n620) );
  AND2_X1 U351bar ( .A1(inbar[95]), .A2(inbar[92]), .ZN(n620bar);
  OR2_X1 U352 ( .A1(n618), .A2(n617), .ZN(n622) );
  AND2_X1 U352bar ( .A1(n618bar), .A2(n617bar), .ZN(n622bar);
  OR2_X1 U353 ( .A1(in_22), .A2(in_16), .ZN(n617) );
  AND2_X1 U353bar ( .A1(in_22bar), .A2(in_16bar), .ZN(n617bar);
  OR2_X1 U354 ( .A1(in_51), .A2(in_49), .ZN(n618) );
  AND2_X1 U354bar ( .A1(in_51bar), .A2(in_49bar), .ZN(n618bar);
  OR2_X1 U355 ( .A1(n616), .A2(n615), .ZN(n722) );
  AND2_X1 U355bar ( .A1(n616bar), .A2(n615bar), .ZN(n722bar);
  OR2_X1 U356 ( .A1(in[158]), .A2(in[115]), .ZN(n615) );
  AND2_X1 U356bar ( .A1(inbar[158]), .A2(inbar[115]), .ZN(n615bar);
  OR2_X1 U357 ( .A1(in[163]), .A2(n614), .ZN(n616) );
  AND2_X1 U357bar ( .A1(inbar[163]), .A2(n614bar), .ZN(n616bar);
  OR2_X1 U358 ( .A1(in[206]), .A2(in[165]), .ZN(n614) );
  AND2_X1 U358bar ( .A1(inbar[206]), .A2(inbar[165]), .ZN(n614bar);
  OR2_X1 U359 ( .A1(n613), .A2(n612), .ZN(n724) );
  AND2_X1 U359bar ( .A1(n613bar), .A2(n612bar), .ZN(n724bar);
  OR2_X1 U360 ( .A1(n611), .A2(n610), .ZN(n612) );
  AND2_X1 U360bar ( .A1(n611bar), .A2(n610bar), .ZN(n612bar);
  OR2_X1 U361 ( .A1(in[213]), .A2(in[207]), .ZN(n610) );
  AND2_X1 U361bar ( .A1(inbar[213]), .A2(inbar[207]), .ZN(n610bar);
  OR2_X1 U362 ( .A1(in[215]), .A2(n609), .ZN(n611) );
  AND2_X1 U362bar ( .A1(inbar[215]), .A2(n609bar), .ZN(n611bar);
  OR2_X1 U363 ( .A1(in[230]), .A2(in[220]), .ZN(n609) );
  AND2_X1 U363bar ( .A1(inbar[230]), .A2(inbar[220]), .ZN(n609bar);
  OR2_X1 U364 ( .A1(n608), .A2(n607), .ZN(n613) );
  AND2_X1 U364bar ( .A1(n608bar), .A2(n607bar), .ZN(n613bar);
  OR2_X1 U365 ( .A1(in[251]), .A2(in[234]), .ZN(n607) );
  AND2_X1 U365bar ( .A1(inbar[251]), .A2(inbar[234]), .ZN(n607bar);
  OR2_X1 U366 ( .A1(in_17), .A2(n606), .ZN(n608) );
  AND2_X1 U366bar ( .A1(in_17bar), .A2(n606bar), .ZN(n608bar);
  OR2_X1 U367 ( .A1(in_65), .A2(in_56), .ZN(n606) );
  AND2_X1 U367bar ( .A1(in_65bar), .A2(in_56bar), .ZN(n606bar);
  OR2_X1 U368 ( .A1(n605), .A2(n604), .ZN(out[0]) );
  AND2_X1 U368bar ( .A1(n605bar), .A2(n604bar), .ZN(outbar[0]);
  OR2_X1 U369 ( .A1(n603), .A2(n602), .ZN(n604) );
  AND2_X1 U369bar ( .A1(n603bar), .A2(n602bar), .ZN(n604bar);
  OR2_X1 U370 ( .A1(n601), .A2(n600), .ZN(n602) );
  AND2_X1 U370bar ( .A1(n601bar), .A2(n600bar), .ZN(n602bar);
  OR2_X1 U371 ( .A1(n820), .A2(n785), .ZN(n600) );
  AND2_X1 U371bar ( .A1(n820bar), .A2(n785bar), .ZN(n600bar);
  OR2_X1 U372 ( .A1(n599), .A2(n598), .ZN(n785) );
  AND2_X1 U372bar ( .A1(n599bar), .A2(n598bar), .ZN(n785bar);
  OR2_X1 U373 ( .A1(n597), .A2(n596), .ZN(n598) );
  AND2_X1 U373bar ( .A1(n597bar), .A2(n596bar), .ZN(n598bar);
  OR2_X1 U374 ( .A1(n595), .A2(n594), .ZN(n596) );
  AND2_X1 U374bar ( .A1(n595bar), .A2(n594bar), .ZN(n596bar);
  OR2_X1 U375 ( .A1(in[135]), .A2(in[104]), .ZN(n594) );
  AND2_X1 U375bar ( .A1(inbar[135]), .A2(inbar[104]), .ZN(n594bar);
  OR2_X1 U376 ( .A1(in[188]), .A2(in[178]), .ZN(n595) );
  AND2_X1 U376bar ( .A1(inbar[188]), .A2(inbar[178]), .ZN(n595bar);
  OR2_X1 U377 ( .A1(n593), .A2(n592), .ZN(n597) );
  AND2_X1 U377bar ( .A1(n593bar), .A2(n592bar), .ZN(n597bar);
  OR2_X1 U378 ( .A1(in[217]), .A2(in[194]), .ZN(n592) );
  AND2_X1 U378bar ( .A1(inbar[217]), .A2(inbar[194]), .ZN(n592bar);
  OR2_X1 U379 ( .A1(in[237]), .A2(in[218]), .ZN(n593) );
  AND2_X1 U379bar ( .A1(inbar[237]), .A2(inbar[218]), .ZN(n593bar);
  OR2_X1 U380 ( .A1(n591), .A2(n590), .ZN(n599) );
  AND2_X1 U380bar ( .A1(n591bar), .A2(n590bar), .ZN(n599bar);
  OR2_X1 U381 ( .A1(n589), .A2(n588), .ZN(n590) );
  AND2_X1 U381bar ( .A1(n589bar), .A2(n588bar), .ZN(n590bar);
  OR2_X1 U382 ( .A1(in_2), .A2(in_10), .ZN(n588) );
  AND2_X1 U382bar ( .A1(in_2bar), .A2(in_10bar), .ZN(n588bar);
  OR2_X1 U383 ( .A1(in_47), .A2(in_22), .ZN(n589) );
  AND2_X1 U383bar ( .A1(in_47bar), .A2(in_22bar), .ZN(n589bar);
  OR2_X1 U384 ( .A1(n587), .A2(n586), .ZN(n591) );
  AND2_X1 U384bar ( .A1(n587bar), .A2(n586bar), .ZN(n591bar);
  OR2_X1 U385 ( .A1(in_56), .A2(in_54), .ZN(n586) );
  AND2_X1 U385bar ( .A1(in_56bar), .A2(in_54bar), .ZN(n586bar);
  OR2_X1 U386 ( .A1(in_63), .A2(in_61), .ZN(n587) );
  AND2_X1 U386bar ( .A1(in_63bar), .A2(in_61bar), .ZN(n587bar);
  OR2_X1 U387 ( .A1(n585), .A2(n584), .ZN(n820) );
  AND2_X1 U387bar ( .A1(n585bar), .A2(n584bar), .ZN(n820bar);
  OR2_X1 U388 ( .A1(n583), .A2(n582), .ZN(n584) );
  AND2_X1 U388bar ( .A1(n583bar), .A2(n582bar), .ZN(n584bar);
  OR2_X1 U389 ( .A1(n581), .A2(n580), .ZN(n582) );
  AND2_X1 U389bar ( .A1(n581bar), .A2(n580bar), .ZN(n582bar);
  OR2_X1 U390 ( .A1(in[158]), .A2(in[142]), .ZN(n580) );
  AND2_X1 U390bar ( .A1(inbar[158]), .A2(inbar[142]), .ZN(n580bar);
  OR2_X1 U391 ( .A1(in[175]), .A2(in[164]), .ZN(n581) );
  AND2_X1 U391bar ( .A1(inbar[175]), .A2(inbar[164]), .ZN(n581bar);
  OR2_X1 U392 ( .A1(n579), .A2(n578), .ZN(n583) );
  AND2_X1 U392bar ( .A1(n579bar), .A2(n578bar), .ZN(n583bar);
  OR2_X1 U393 ( .A1(in[228]), .A2(in[204]), .ZN(n578) );
  AND2_X1 U393bar ( .A1(inbar[228]), .A2(inbar[204]), .ZN(n578bar);
  OR2_X1 U394 ( .A1(in[91]), .A2(in[87]), .ZN(n579) );
  AND2_X1 U394bar ( .A1(inbar[91]), .A2(inbar[87]), .ZN(n579bar);
  OR2_X1 U395 ( .A1(n577), .A2(n576), .ZN(n585) );
  AND2_X1 U395bar ( .A1(n577bar), .A2(n576bar), .ZN(n585bar);
  OR2_X1 U396 ( .A1(n575), .A2(n574), .ZN(n576) );
  AND2_X1 U396bar ( .A1(n575bar), .A2(n574bar), .ZN(n576bar);
  OR2_X1 U397 ( .A1(in_21), .A2(in_11), .ZN(n574) );
  AND2_X1 U397bar ( .A1(in_21bar), .A2(in_11bar), .ZN(n574bar);
  OR2_X1 U398 ( .A1(in_5), .A2(in_3), .ZN(n575) );
  AND2_X1 U398bar ( .A1(in_5bar), .A2(in_3bar), .ZN(n575bar);
  OR2_X1 U399 ( .A1(n573), .A2(n572), .ZN(n577) );
  AND2_X1 U399bar ( .A1(n573bar), .A2(n572bar), .ZN(n577bar);
  OR2_X1 U400 ( .A1(in_68), .A2(in_64), .ZN(n572) );
  AND2_X1 U400bar ( .A1(in_68bar), .A2(in_64bar), .ZN(n572bar);
  OR2_X1 U401 ( .A1(in_76), .A2(in_73), .ZN(n573) );
  AND2_X1 U401bar ( .A1(in_76bar), .A2(in_73bar), .ZN(n573bar);
  OR2_X1 U402 ( .A1(n778), .A2(n571), .ZN(n601) );
  AND2_X1 U402bar ( .A1(n778bar), .A2(n571bar), .ZN(n601bar);
  OR2_X1 U403 ( .A1(in[100]), .A2(n965), .ZN(n571) );
  AND2_X1 U403bar ( .A1(inbar[100]), .A2(n965bar), .ZN(n571bar);
  OR2_X1 U404 ( .A1(n570), .A2(n569), .ZN(n965) );
  AND2_X1 U404bar ( .A1(n570bar), .A2(n569bar), .ZN(n965bar);
  OR2_X1 U405 ( .A1(n568), .A2(n567), .ZN(n569) );
  AND2_X1 U405bar ( .A1(n568bar), .A2(n567bar), .ZN(n569bar);
  OR2_X1 U406 ( .A1(n566), .A2(n565), .ZN(n567) );
  AND2_X1 U406bar ( .A1(n566bar), .A2(n565bar), .ZN(n567bar);
  OR2_X1 U407 ( .A1(n817), .A2(n750), .ZN(n565) );
  AND2_X1 U407bar ( .A1(n817bar), .A2(n750bar), .ZN(n565bar);
  OR2_X1 U408 ( .A1(n564), .A2(n563), .ZN(n750) );
  AND2_X1 U408bar ( .A1(n564bar), .A2(n563bar), .ZN(n750bar);
  OR2_X1 U409 ( .A1(n562), .A2(n561), .ZN(n563) );
  AND2_X1 U409bar ( .A1(n562bar), .A2(n561bar), .ZN(n563bar);
  OR2_X1 U410 ( .A1(n560), .A2(n559), .ZN(n561) );
  AND2_X1 U410bar ( .A1(n560bar), .A2(n559bar), .ZN(n561bar);
  OR2_X1 U411 ( .A1(in[119]), .A2(in[103]), .ZN(n559) );
  AND2_X1 U411bar ( .A1(inbar[119]), .A2(inbar[103]), .ZN(n559bar);
  OR2_X1 U412 ( .A1(in[137]), .A2(in[133]), .ZN(n560) );
  AND2_X1 U412bar ( .A1(inbar[137]), .A2(inbar[133]), .ZN(n560bar);
  OR2_X1 U413 ( .A1(n558), .A2(n557), .ZN(n562) );
  AND2_X1 U413bar ( .A1(n558bar), .A2(n557bar), .ZN(n562bar);
  OR2_X1 U414 ( .A1(in[176]), .A2(in[173]), .ZN(n557) );
  AND2_X1 U414bar ( .A1(inbar[176]), .A2(inbar[173]), .ZN(n557bar);
  OR2_X1 U415 ( .A1(in[210]), .A2(in[181]), .ZN(n558) );
  AND2_X1 U415bar ( .A1(inbar[210]), .A2(inbar[181]), .ZN(n558bar);
  OR2_X1 U416 ( .A1(n556), .A2(n555), .ZN(n564) );
  AND2_X1 U416bar ( .A1(n556bar), .A2(n555bar), .ZN(n564bar);
  OR2_X1 U417 ( .A1(n554), .A2(n553), .ZN(n555) );
  AND2_X1 U417bar ( .A1(n554bar), .A2(n553bar), .ZN(n555bar);
  OR2_X1 U418 ( .A1(in_13), .A2(in[234]), .ZN(n553) );
  AND2_X1 U418bar ( .A1(in_13bar), .A2(inbar[234]), .ZN(n553bar);
  OR2_X1 U419 ( .A1(in_38), .A2(in_32), .ZN(n554) );
  AND2_X1 U419bar ( .A1(in_38bar), .A2(in_32bar), .ZN(n554bar);
  OR2_X1 U420 ( .A1(n552), .A2(n551), .ZN(n556) );
  AND2_X1 U420bar ( .A1(n552bar), .A2(n551bar), .ZN(n556bar);
  OR2_X1 U421 ( .A1(in_42), .A2(in_41), .ZN(n551) );
  AND2_X1 U421bar ( .A1(in_42bar), .A2(in_41bar), .ZN(n551bar);
  OR2_X1 U422 ( .A1(in_7), .A2(in_49), .ZN(n552) );
  AND2_X1 U422bar ( .A1(in_7bar), .A2(in_49bar), .ZN(n552bar);
  OR2_X1 U423 ( .A1(n550), .A2(n549), .ZN(n817) );
  AND2_X1 U423bar ( .A1(n550bar), .A2(n549bar), .ZN(n817bar);
  OR2_X1 U424 ( .A1(n548), .A2(n547), .ZN(n549) );
  AND2_X1 U424bar ( .A1(n548bar), .A2(n547bar), .ZN(n549bar);
  OR2_X1 U425 ( .A1(n546), .A2(n545), .ZN(n547) );
  AND2_X1 U425bar ( .A1(n546bar), .A2(n545bar), .ZN(n547bar);
  OR2_X1 U426 ( .A1(in[159]), .A2(in[105]), .ZN(n545) );
  AND2_X1 U426bar ( .A1(inbar[159]), .A2(inbar[105]), .ZN(n545bar);
  OR2_X1 U427 ( .A1(in[206]), .A2(in[183]), .ZN(n546) );
  AND2_X1 U427bar ( .A1(inbar[206]), .A2(inbar[183]), .ZN(n546bar);
  OR2_X1 U428 ( .A1(n544), .A2(n543), .ZN(n548) );
  AND2_X1 U428bar ( .A1(n544bar), .A2(n543bar), .ZN(n548bar);
  OR2_X1 U429 ( .A1(in[229]), .A2(in[219]), .ZN(n543) );
  AND2_X1 U429bar ( .A1(inbar[229]), .A2(inbar[219]), .ZN(n543bar);
  OR2_X1 U430 ( .A1(in[235]), .A2(in[232]), .ZN(n544) );
  AND2_X1 U430bar ( .A1(inbar[235]), .A2(inbar[232]), .ZN(n544bar);
  OR2_X1 U431 ( .A1(n542), .A2(n541), .ZN(n550) );
  AND2_X1 U431bar ( .A1(n542bar), .A2(n541bar), .ZN(n550bar);
  OR2_X1 U432 ( .A1(n540), .A2(n539), .ZN(n541) );
  AND2_X1 U432bar ( .A1(n540bar), .A2(n539bar), .ZN(n541bar);
  OR2_X1 U433 ( .A1(in[249]), .A2(in[242]), .ZN(n539) );
  AND2_X1 U433bar ( .A1(inbar[249]), .A2(inbar[242]), .ZN(n539bar);
  OR2_X1 U434 ( .A1(in[89]), .A2(in[254]), .ZN(n540) );
  AND2_X1 U434bar ( .A1(inbar[89]), .A2(inbar[254]), .ZN(n540bar);
  OR2_X1 U435 ( .A1(n538), .A2(n537), .ZN(n542) );
  AND2_X1 U435bar ( .A1(n538bar), .A2(n537bar), .ZN(n542bar);
  OR2_X1 U436 ( .A1(in_14), .A2(in[99]), .ZN(n537) );
  AND2_X1 U436bar ( .A1(in_14bar), .A2(inbar[99]), .ZN(n537bar);
  OR2_X1 U437 ( .A1(in_60), .A2(in_18), .ZN(n538) );
  AND2_X1 U437bar ( .A1(in_60bar), .A2(in_18bar), .ZN(n538bar);
  OR2_X1 U438 ( .A1(in[113]), .A2(n763), .ZN(n566) );
  AND2_X1 U438bar ( .A1(inbar[113]), .A2(n763bar), .ZN(n566bar);
  OR2_X1 U439 ( .A1(n536), .A2(n535), .ZN(n763) );
  AND2_X1 U439bar ( .A1(n536bar), .A2(n535bar), .ZN(n763bar);
  OR2_X1 U440 ( .A1(n534), .A2(n533), .ZN(n535) );
  AND2_X1 U440bar ( .A1(n534bar), .A2(n533bar), .ZN(n535bar);
  OR2_X1 U441 ( .A1(n532), .A2(n531), .ZN(n533) );
  AND2_X1 U441bar ( .A1(n532bar), .A2(n531bar), .ZN(n533bar);
  OR2_X1 U442 ( .A1(in[115]), .A2(in[110]), .ZN(n531) );
  AND2_X1 U442bar ( .A1(inbar[115]), .A2(inbar[110]), .ZN(n531bar);
  OR2_X1 U443 ( .A1(in[125]), .A2(in[117]), .ZN(n532) );
  AND2_X1 U443bar ( .A1(inbar[125]), .A2(inbar[117]), .ZN(n532bar);
  OR2_X1 U444 ( .A1(n530), .A2(n529), .ZN(n534) );
  AND2_X1 U444bar ( .A1(n530bar), .A2(n529bar), .ZN(n534bar);
  OR2_X1 U445 ( .A1(in[180]), .A2(in[128]), .ZN(n529) );
  AND2_X1 U445bar ( .A1(inbar[180]), .A2(inbar[128]), .ZN(n529bar);
  OR2_X1 U446 ( .A1(in[205]), .A2(in[201]), .ZN(n530) );
  AND2_X1 U446bar ( .A1(inbar[205]), .A2(inbar[201]), .ZN(n530bar);
  OR2_X1 U447 ( .A1(n528), .A2(n527), .ZN(n536) );
  AND2_X1 U447bar ( .A1(n528bar), .A2(n527bar), .ZN(n536bar);
  OR2_X1 U448 ( .A1(n526), .A2(n525), .ZN(n527) );
  AND2_X1 U448bar ( .A1(n526bar), .A2(n525bar), .ZN(n527bar);
  OR2_X1 U449 ( .A1(in[244]), .A2(in[239]), .ZN(n525) );
  AND2_X1 U449bar ( .A1(inbar[244]), .A2(inbar[239]), .ZN(n525bar);
  OR2_X1 U450 ( .A1(in[95]), .A2(in[83]), .ZN(n526) );
  AND2_X1 U450bar ( .A1(inbar[95]), .A2(inbar[83]), .ZN(n526bar);
  OR2_X1 U451 ( .A1(n524), .A2(n523), .ZN(n528) );
  AND2_X1 U451bar ( .A1(n524bar), .A2(n523bar), .ZN(n528bar);
  OR2_X1 U452 ( .A1(in_24), .A2(in[97]), .ZN(n523) );
  AND2_X1 U452bar ( .A1(in_24bar), .A2(inbar[97]), .ZN(n523bar);
  OR2_X1 U453 ( .A1(in_33), .A2(in_27), .ZN(n524) );
  AND2_X1 U453bar ( .A1(in_33bar), .A2(in_27bar), .ZN(n524bar);
  OR2_X1 U454 ( .A1(n522), .A2(n521), .ZN(n568) );
  AND2_X1 U454bar ( .A1(n522bar), .A2(n521bar), .ZN(n568bar);
  OR2_X1 U455 ( .A1(in[145]), .A2(in[126]), .ZN(n521) );
  AND2_X1 U455bar ( .A1(inbar[145]), .A2(inbar[126]), .ZN(n521bar);
  OR2_X1 U456 ( .A1(in[169]), .A2(n520), .ZN(n522) );
  AND2_X1 U456bar ( .A1(inbar[169]), .A2(n520bar), .ZN(n522bar);
  OR2_X1 U457 ( .A1(in[221]), .A2(in[172]), .ZN(n520) );
  AND2_X1 U457bar ( .A1(inbar[221]), .A2(inbar[172]), .ZN(n520bar);
  OR2_X1 U458 ( .A1(n519), .A2(n518), .ZN(n570) );
  AND2_X1 U458bar ( .A1(n519bar), .A2(n518bar), .ZN(n570bar);
  OR2_X1 U459 ( .A1(n517), .A2(n516), .ZN(n518) );
  AND2_X1 U459bar ( .A1(n517bar), .A2(n516bar), .ZN(n518bar);
  OR2_X1 U460 ( .A1(in[241]), .A2(in[224]), .ZN(n516) );
  AND2_X1 U460bar ( .A1(inbar[241]), .A2(inbar[224]), .ZN(n516bar);
  OR2_X1 U461 ( .A1(in[86]), .A2(n515), .ZN(n517) );
  AND2_X1 U461bar ( .A1(inbar[86]), .A2(n515bar), .ZN(n517bar);
  OR2_X1 U462 ( .A1(in_43), .A2(in_34), .ZN(n515) );
  AND2_X1 U462bar ( .A1(in_43bar), .A2(in_34bar), .ZN(n515bar);
  OR2_X1 U463 ( .A1(n514), .A2(n513), .ZN(n519) );
  AND2_X1 U463bar ( .A1(n514bar), .A2(n513bar), .ZN(n519bar);
  OR2_X1 U464 ( .A1(in_65), .A2(in_51), .ZN(n513) );
  AND2_X1 U464bar ( .A1(in_65bar), .A2(in_51bar), .ZN(n513bar);
  OR2_X1 U465 ( .A1(in_75), .A2(n512), .ZN(n514) );
  AND2_X1 U465bar ( .A1(in_75bar), .A2(n512bar), .ZN(n514bar);
  OR2_X1 U466 ( .A1(in_81), .A2(in_77), .ZN(n512) );
  AND2_X1 U466bar ( .A1(in_81bar), .A2(in_77bar), .ZN(n512bar);
  OR2_X1 U467 ( .A1(n511), .A2(n510), .ZN(n778) );
  AND2_X1 U467bar ( .A1(n511bar), .A2(n510bar), .ZN(n778bar);
  OR2_X1 U468 ( .A1(n509), .A2(n508), .ZN(n510) );
  AND2_X1 U468bar ( .A1(n509bar), .A2(n508bar), .ZN(n510bar);
  OR2_X1 U469 ( .A1(n507), .A2(n506), .ZN(n508) );
  AND2_X1 U469bar ( .A1(n507bar), .A2(n506bar), .ZN(n508bar);
  OR2_X1 U470 ( .A1(in[107]), .A2(in[101]), .ZN(n506) );
  AND2_X1 U470bar ( .A1(inbar[107]), .A2(inbar[101]), .ZN(n506bar);
  OR2_X1 U471 ( .A1(in[139]), .A2(in[132]), .ZN(n507) );
  AND2_X1 U471bar ( .A1(inbar[139]), .A2(inbar[132]), .ZN(n507bar);
  OR2_X1 U472 ( .A1(n505), .A2(n504), .ZN(n509) );
  AND2_X1 U472bar ( .A1(n505bar), .A2(n504bar), .ZN(n509bar);
  OR2_X1 U473 ( .A1(in[146]), .A2(in[141]), .ZN(n504) );
  AND2_X1 U473bar ( .A1(inbar[146]), .A2(inbar[141]), .ZN(n504bar);
  OR2_X1 U474 ( .A1(in[203]), .A2(in[179]), .ZN(n505) );
  AND2_X1 U474bar ( .A1(inbar[203]), .A2(inbar[179]), .ZN(n505bar);
  OR2_X1 U475 ( .A1(n503), .A2(n502), .ZN(n511) );
  AND2_X1 U475bar ( .A1(n503bar), .A2(n502bar), .ZN(n511bar);
  OR2_X1 U476 ( .A1(n501), .A2(n500), .ZN(n502) );
  AND2_X1 U476bar ( .A1(n501bar), .A2(n500bar), .ZN(n502bar);
  OR2_X1 U477 ( .A1(in[243]), .A2(in[222]), .ZN(n500) );
  AND2_X1 U477bar ( .A1(inbar[243]), .A2(inbar[222]), .ZN(n500bar);
  OR2_X1 U478 ( .A1(in[251]), .A2(in[250]), .ZN(n501) );
  AND2_X1 U478bar ( .A1(inbar[251]), .A2(inbar[250]), .ZN(n501bar);
  OR2_X1 U479 ( .A1(n499), .A2(n498), .ZN(n503) );
  AND2_X1 U479bar ( .A1(n499bar), .A2(n498bar), .ZN(n503bar);
  OR2_X1 U480 ( .A1(in_37), .A2(in_19), .ZN(n498) );
  AND2_X1 U480bar ( .A1(in_37bar), .A2(in_19bar), .ZN(n498bar);
  OR2_X1 U481 ( .A1(in_78), .A2(in_6), .ZN(n499) );
  AND2_X1 U481bar ( .A1(in_78bar), .A2(in_6bar), .ZN(n499bar);
  OR2_X1 U482 ( .A1(n497), .A2(n496), .ZN(n603) );
  AND2_X1 U482bar ( .A1(n497bar), .A2(n496bar), .ZN(n603bar);
  OR2_X1 U483 ( .A1(in[112]), .A2(in[102]), .ZN(n496) );
  AND2_X1 U483bar ( .A1(inbar[112]), .A2(inbar[102]), .ZN(n496bar);
  OR2_X1 U484 ( .A1(in[123]), .A2(n495), .ZN(n497) );
  AND2_X1 U484bar ( .A1(inbar[123]), .A2(n495bar), .ZN(n497bar);
  OR2_X1 U485 ( .A1(in[143]), .A2(in[130]), .ZN(n495) );
  AND2_X1 U485bar ( .A1(inbar[143]), .A2(inbar[130]), .ZN(n495bar);
  OR2_X1 U486 ( .A1(n494), .A2(n493), .ZN(n605) );
  AND2_X1 U486bar ( .A1(n494bar), .A2(n493bar), .ZN(n605bar);
  OR2_X1 U487 ( .A1(n492), .A2(n491), .ZN(n493) );
  AND2_X1 U487bar ( .A1(n492bar), .A2(n491bar), .ZN(n493bar);
  OR2_X1 U488 ( .A1(in[216]), .A2(in[213]), .ZN(n491) );
  AND2_X1 U488bar ( .A1(inbar[216]), .A2(inbar[213]), .ZN(n491bar);
  OR2_X1 U489 ( .A1(in[227]), .A2(n490), .ZN(n492) );
  AND2_X1 U489bar ( .A1(inbar[227]), .A2(n490bar), .ZN(n492bar);
  OR2_X1 U490 ( .A1(in_0), .A2(in[248]), .ZN(n490) );
  AND2_X1 U490bar ( .A1(in_0bar), .A2(inbar[248]), .ZN(n490bar);
  OR2_X1 U491 ( .A1(n489), .A2(n488), .ZN(n494) );
  AND2_X1 U491bar ( .A1(n489bar), .A2(n488bar), .ZN(n494bar);
  OR2_X1 U492 ( .A1(in_46), .A2(in_44), .ZN(n488) );
  AND2_X1 U492bar ( .A1(in_46bar), .A2(in_44bar), .ZN(n488bar);
  OR2_X1 U493 ( .A1(in_50), .A2(n487), .ZN(n489) );
  AND2_X1 U493bar ( .A1(in_50bar), .A2(n487bar), .ZN(n489bar);
  OR2_X1 U494 ( .A1(in_9), .A2(in_80), .ZN(n487) );
  AND2_X1 U494bar ( .A1(in_9bar), .A2(in_80bar), .ZN(n487bar);
endmodule




module sBox_12 ( in, out );
  input [7:0] in;
  //input_done

  output [7:0] out;
  //output_done

  wire   [255:0] decodeOut;
  //wire_done

  decode_12 dec ( .in(in), .out(decodeOut) );
  encode_12 enc ( .in(decodeOut), .out(out) );
endmodule


module CD2_49 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_50 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_51 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_52 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD4_25 ( a, b, y );
  input [3:0] a;
  input [3:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  //input_done

  output [15:0] y;
  reg [15:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]);
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]);
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]);
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]);
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]);
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]);
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]);
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]);
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]);
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]);
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]);
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]);
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]);
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]);
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]);
endmodule




module CD4_26 ( a, b, y );
  input [3:0] a;
  input [3:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  //input_done

  output [15:0] y;
  reg [15:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]);
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]);
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]);
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]);
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]);
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]);
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]);
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]);
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]);
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]);
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]);
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]);
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]);
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]);
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]);
endmodule




module CD16_13 ( a, b, y );
  input [15:0] a;
  input [15:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign abar[8] = ~a[8];
  assign abar[9] = ~a[9];
  assign abar[10] = ~a[10];
  assign abar[11] = ~a[11];
  assign abar[12] = ~a[12];
  assign abar[13] = ~a[13];
  assign abar[14] = ~a[14];
  assign abar[15] = ~a[15];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign bbar[8] = ~b[8];
  assign bbar[9] = ~b[9];
  assign bbar[10] = ~b[10];
  assign bbar[11] = ~b[11];
  assign bbar[12] = ~b[12];
  assign bbar[13] = ~b[13];
  assign bbar[14] = ~b[14];
  assign bbar[15] = ~b[15];
  //input_done

  output [255:0] y;
  reg [255:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[9]), .A2(a[0]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[9]), .A2(abar[0]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[3]), .A2(a[6]), .ZN(y[99]) );
  OR2_X1 U2bar ( .A1(bbar[3]), .A2(abar[6]), .ZN(ybar[99]);
  AND2_X1 U3 ( .A1(b[2]), .A2(a[6]), .ZN(y[98]) );
  OR2_X1 U3bar ( .A1(bbar[2]), .A2(abar[6]), .ZN(ybar[98]);
  AND2_X1 U4 ( .A1(b[1]), .A2(a[6]), .ZN(y[97]) );
  OR2_X1 U4bar ( .A1(bbar[1]), .A2(abar[6]), .ZN(ybar[97]);
  AND2_X1 U5 ( .A1(b[0]), .A2(a[6]), .ZN(y[96]) );
  OR2_X1 U5bar ( .A1(bbar[0]), .A2(abar[6]), .ZN(ybar[96]);
  AND2_X1 U6 ( .A1(b[15]), .A2(a[5]), .ZN(y[95]) );
  OR2_X1 U6bar ( .A1(bbar[15]), .A2(abar[5]), .ZN(ybar[95]);
  AND2_X1 U7 ( .A1(b[14]), .A2(a[5]), .ZN(y[94]) );
  OR2_X1 U7bar ( .A1(bbar[14]), .A2(abar[5]), .ZN(ybar[94]);
  AND2_X1 U8 ( .A1(b[13]), .A2(a[5]), .ZN(y[93]) );
  OR2_X1 U8bar ( .A1(bbar[13]), .A2(abar[5]), .ZN(ybar[93]);
  AND2_X1 U9 ( .A1(b[12]), .A2(a[5]), .ZN(y[92]) );
  OR2_X1 U9bar ( .A1(bbar[12]), .A2(abar[5]), .ZN(ybar[92]);
  AND2_X1 U10 ( .A1(b[11]), .A2(a[5]), .ZN(y[91]) );
  OR2_X1 U10bar ( .A1(bbar[11]), .A2(abar[5]), .ZN(ybar[91]);
  AND2_X1 U11 ( .A1(b[10]), .A2(a[5]), .ZN(y[90]) );
  OR2_X1 U11bar ( .A1(bbar[10]), .A2(abar[5]), .ZN(ybar[90]);
  AND2_X1 U12 ( .A1(b[8]), .A2(a[0]), .ZN(y[8]) );
  OR2_X1 U12bar ( .A1(bbar[8]), .A2(abar[0]), .ZN(ybar[8]);
  AND2_X1 U13 ( .A1(a[5]), .A2(b[9]), .ZN(y[89]) );
  OR2_X1 U13bar ( .A1(abar[5]), .A2(bbar[9]), .ZN(ybar[89]);
  AND2_X1 U14 ( .A1(b[8]), .A2(a[5]), .ZN(y[88]) );
  OR2_X1 U14bar ( .A1(bbar[8]), .A2(abar[5]), .ZN(ybar[88]);
  AND2_X1 U15 ( .A1(b[7]), .A2(a[5]), .ZN(y[87]) );
  OR2_X1 U15bar ( .A1(bbar[7]), .A2(abar[5]), .ZN(ybar[87]);
  AND2_X1 U16 ( .A1(b[6]), .A2(a[5]), .ZN(y[86]) );
  OR2_X1 U16bar ( .A1(bbar[6]), .A2(abar[5]), .ZN(ybar[86]);
  AND2_X1 U17 ( .A1(b[5]), .A2(a[5]), .ZN(y[85]) );
  OR2_X1 U17bar ( .A1(bbar[5]), .A2(abar[5]), .ZN(ybar[85]);
  AND2_X1 U18 ( .A1(b[4]), .A2(a[5]), .ZN(y[84]) );
  OR2_X1 U18bar ( .A1(bbar[4]), .A2(abar[5]), .ZN(ybar[84]);
  AND2_X1 U19 ( .A1(a[5]), .A2(b[3]), .ZN(y[83]) );
  OR2_X1 U19bar ( .A1(abar[5]), .A2(bbar[3]), .ZN(ybar[83]);
  AND2_X1 U20 ( .A1(a[5]), .A2(b[2]), .ZN(y[82]) );
  OR2_X1 U20bar ( .A1(abar[5]), .A2(bbar[2]), .ZN(ybar[82]);
  AND2_X1 U21 ( .A1(a[5]), .A2(b[1]), .ZN(y[81]) );
  OR2_X1 U21bar ( .A1(abar[5]), .A2(bbar[1]), .ZN(ybar[81]);
  AND2_X1 U22 ( .A1(a[5]), .A2(b[0]), .ZN(y[80]) );
  OR2_X1 U22bar ( .A1(abar[5]), .A2(bbar[0]), .ZN(ybar[80]);
  AND2_X1 U23 ( .A1(b[7]), .A2(a[0]), .ZN(y[7]) );
  OR2_X1 U23bar ( .A1(bbar[7]), .A2(abar[0]), .ZN(ybar[7]);
  AND2_X1 U24 ( .A1(a[4]), .A2(b[15]), .ZN(y[79]) );
  OR2_X1 U24bar ( .A1(abar[4]), .A2(bbar[15]), .ZN(ybar[79]);
  AND2_X1 U25 ( .A1(a[4]), .A2(b[14]), .ZN(y[78]) );
  OR2_X1 U25bar ( .A1(abar[4]), .A2(bbar[14]), .ZN(ybar[78]);
  AND2_X1 U26 ( .A1(a[4]), .A2(b[13]), .ZN(y[77]) );
  OR2_X1 U26bar ( .A1(abar[4]), .A2(bbar[13]), .ZN(ybar[77]);
  AND2_X1 U27 ( .A1(a[4]), .A2(b[12]), .ZN(y[76]) );
  OR2_X1 U27bar ( .A1(abar[4]), .A2(bbar[12]), .ZN(ybar[76]);
  AND2_X1 U28 ( .A1(a[4]), .A2(b[11]), .ZN(y[75]) );
  OR2_X1 U28bar ( .A1(abar[4]), .A2(bbar[11]), .ZN(ybar[75]);
  AND2_X1 U29 ( .A1(a[4]), .A2(b[10]), .ZN(y[74]) );
  OR2_X1 U29bar ( .A1(abar[4]), .A2(bbar[10]), .ZN(ybar[74]);
  AND2_X1 U30 ( .A1(a[4]), .A2(b[9]), .ZN(y[73]) );
  OR2_X1 U30bar ( .A1(abar[4]), .A2(bbar[9]), .ZN(ybar[73]);
  AND2_X1 U31 ( .A1(a[4]), .A2(b[8]), .ZN(y[72]) );
  OR2_X1 U31bar ( .A1(abar[4]), .A2(bbar[8]), .ZN(ybar[72]);
  AND2_X1 U32 ( .A1(a[4]), .A2(b[7]), .ZN(y[71]) );
  OR2_X1 U32bar ( .A1(abar[4]), .A2(bbar[7]), .ZN(ybar[71]);
  AND2_X1 U33 ( .A1(a[4]), .A2(b[6]), .ZN(y[70]) );
  OR2_X1 U33bar ( .A1(abar[4]), .A2(bbar[6]), .ZN(ybar[70]);
  AND2_X1 U34 ( .A1(b[6]), .A2(a[0]), .ZN(y[6]) );
  OR2_X1 U34bar ( .A1(bbar[6]), .A2(abar[0]), .ZN(ybar[6]);
  AND2_X1 U35 ( .A1(a[4]), .A2(b[5]), .ZN(y[69]) );
  OR2_X1 U35bar ( .A1(abar[4]), .A2(bbar[5]), .ZN(ybar[69]);
  AND2_X1 U36 ( .A1(a[4]), .A2(b[4]), .ZN(y[68]) );
  OR2_X1 U36bar ( .A1(abar[4]), .A2(bbar[4]), .ZN(ybar[68]);
  AND2_X1 U37 ( .A1(a[4]), .A2(b[3]), .ZN(y[67]) );
  OR2_X1 U37bar ( .A1(abar[4]), .A2(bbar[3]), .ZN(ybar[67]);
  AND2_X1 U38 ( .A1(a[4]), .A2(b[2]), .ZN(y[66]) );
  OR2_X1 U38bar ( .A1(abar[4]), .A2(bbar[2]), .ZN(ybar[66]);
  AND2_X1 U39 ( .A1(a[4]), .A2(b[1]), .ZN(y[65]) );
  OR2_X1 U39bar ( .A1(abar[4]), .A2(bbar[1]), .ZN(ybar[65]);
  AND2_X1 U40 ( .A1(a[4]), .A2(b[0]), .ZN(y[64]) );
  OR2_X1 U40bar ( .A1(abar[4]), .A2(bbar[0]), .ZN(ybar[64]);
  AND2_X1 U41 ( .A1(a[3]), .A2(b[15]), .ZN(y[63]) );
  OR2_X1 U41bar ( .A1(abar[3]), .A2(bbar[15]), .ZN(ybar[63]);
  AND2_X1 U42 ( .A1(a[3]), .A2(b[14]), .ZN(y[62]) );
  OR2_X1 U42bar ( .A1(abar[3]), .A2(bbar[14]), .ZN(ybar[62]);
  AND2_X1 U43 ( .A1(a[3]), .A2(b[13]), .ZN(y[61]) );
  OR2_X1 U43bar ( .A1(abar[3]), .A2(bbar[13]), .ZN(ybar[61]);
  AND2_X1 U44 ( .A1(a[3]), .A2(b[12]), .ZN(y[60]) );
  OR2_X1 U44bar ( .A1(abar[3]), .A2(bbar[12]), .ZN(ybar[60]);
  AND2_X1 U45 ( .A1(b[5]), .A2(a[0]), .ZN(y[5]) );
  OR2_X1 U45bar ( .A1(bbar[5]), .A2(abar[0]), .ZN(ybar[5]);
  AND2_X1 U46 ( .A1(a[3]), .A2(b[11]), .ZN(y[59]) );
  OR2_X1 U46bar ( .A1(abar[3]), .A2(bbar[11]), .ZN(ybar[59]);
  AND2_X1 U47 ( .A1(a[3]), .A2(b[10]), .ZN(y[58]) );
  OR2_X1 U47bar ( .A1(abar[3]), .A2(bbar[10]), .ZN(ybar[58]);
  AND2_X1 U48 ( .A1(a[3]), .A2(b[9]), .ZN(y[57]) );
  OR2_X1 U48bar ( .A1(abar[3]), .A2(bbar[9]), .ZN(ybar[57]);
  AND2_X1 U49 ( .A1(a[3]), .A2(b[8]), .ZN(y[56]) );
  OR2_X1 U49bar ( .A1(abar[3]), .A2(bbar[8]), .ZN(ybar[56]);
  AND2_X1 U50 ( .A1(a[3]), .A2(b[7]), .ZN(y[55]) );
  OR2_X1 U50bar ( .A1(abar[3]), .A2(bbar[7]), .ZN(ybar[55]);
  AND2_X1 U51 ( .A1(a[3]), .A2(b[6]), .ZN(y[54]) );
  OR2_X1 U51bar ( .A1(abar[3]), .A2(bbar[6]), .ZN(ybar[54]);
  AND2_X1 U52 ( .A1(a[3]), .A2(b[5]), .ZN(y[53]) );
  OR2_X1 U52bar ( .A1(abar[3]), .A2(bbar[5]), .ZN(ybar[53]);
  AND2_X1 U53 ( .A1(a[3]), .A2(b[4]), .ZN(y[52]) );
  OR2_X1 U53bar ( .A1(abar[3]), .A2(bbar[4]), .ZN(ybar[52]);
  AND2_X1 U54 ( .A1(a[3]), .A2(b[3]), .ZN(y[51]) );
  OR2_X1 U54bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[51]);
  AND2_X1 U55 ( .A1(a[3]), .A2(b[2]), .ZN(y[50]) );
  OR2_X1 U55bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[50]);
  AND2_X1 U56 ( .A1(b[4]), .A2(a[0]), .ZN(y[4]) );
  OR2_X1 U56bar ( .A1(bbar[4]), .A2(abar[0]), .ZN(ybar[4]);
  AND2_X1 U57 ( .A1(a[3]), .A2(b[1]), .ZN(y[49]) );
  OR2_X1 U57bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[49]);
  AND2_X1 U58 ( .A1(a[3]), .A2(b[0]), .ZN(y[48]) );
  OR2_X1 U58bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[48]);
  AND2_X1 U59 ( .A1(a[2]), .A2(b[15]), .ZN(y[47]) );
  OR2_X1 U59bar ( .A1(abar[2]), .A2(bbar[15]), .ZN(ybar[47]);
  AND2_X1 U60 ( .A1(a[2]), .A2(b[14]), .ZN(y[46]) );
  OR2_X1 U60bar ( .A1(abar[2]), .A2(bbar[14]), .ZN(ybar[46]);
  AND2_X1 U61 ( .A1(a[2]), .A2(b[13]), .ZN(y[45]) );
  OR2_X1 U61bar ( .A1(abar[2]), .A2(bbar[13]), .ZN(ybar[45]);
  AND2_X1 U62 ( .A1(a[2]), .A2(b[12]), .ZN(y[44]) );
  OR2_X1 U62bar ( .A1(abar[2]), .A2(bbar[12]), .ZN(ybar[44]);
  AND2_X1 U63 ( .A1(a[2]), .A2(b[11]), .ZN(y[43]) );
  OR2_X1 U63bar ( .A1(abar[2]), .A2(bbar[11]), .ZN(ybar[43]);
  AND2_X1 U64 ( .A1(a[2]), .A2(b[10]), .ZN(y[42]) );
  OR2_X1 U64bar ( .A1(abar[2]), .A2(bbar[10]), .ZN(ybar[42]);
  AND2_X1 U65 ( .A1(a[2]), .A2(b[9]), .ZN(y[41]) );
  OR2_X1 U65bar ( .A1(abar[2]), .A2(bbar[9]), .ZN(ybar[41]);
  AND2_X1 U66 ( .A1(a[2]), .A2(b[8]), .ZN(y[40]) );
  OR2_X1 U66bar ( .A1(abar[2]), .A2(bbar[8]), .ZN(ybar[40]);
  AND2_X1 U67 ( .A1(b[3]), .A2(a[0]), .ZN(y[3]) );
  OR2_X1 U67bar ( .A1(bbar[3]), .A2(abar[0]), .ZN(ybar[3]);
  AND2_X1 U68 ( .A1(a[2]), .A2(b[7]), .ZN(y[39]) );
  OR2_X1 U68bar ( .A1(abar[2]), .A2(bbar[7]), .ZN(ybar[39]);
  AND2_X1 U69 ( .A1(a[2]), .A2(b[6]), .ZN(y[38]) );
  OR2_X1 U69bar ( .A1(abar[2]), .A2(bbar[6]), .ZN(ybar[38]);
  AND2_X1 U70 ( .A1(a[2]), .A2(b[5]), .ZN(y[37]) );
  OR2_X1 U70bar ( .A1(abar[2]), .A2(bbar[5]), .ZN(ybar[37]);
  AND2_X1 U71 ( .A1(a[2]), .A2(b[4]), .ZN(y[36]) );
  OR2_X1 U71bar ( .A1(abar[2]), .A2(bbar[4]), .ZN(ybar[36]);
  AND2_X1 U72 ( .A1(a[2]), .A2(b[3]), .ZN(y[35]) );
  OR2_X1 U72bar ( .A1(abar[2]), .A2(bbar[3]), .ZN(ybar[35]);
  AND2_X1 U73 ( .A1(a[2]), .A2(b[2]), .ZN(y[34]) );
  OR2_X1 U73bar ( .A1(abar[2]), .A2(bbar[2]), .ZN(ybar[34]);
  AND2_X1 U74 ( .A1(a[2]), .A2(b[1]), .ZN(y[33]) );
  OR2_X1 U74bar ( .A1(abar[2]), .A2(bbar[1]), .ZN(ybar[33]);
  AND2_X1 U75 ( .A1(a[2]), .A2(b[0]), .ZN(y[32]) );
  OR2_X1 U75bar ( .A1(abar[2]), .A2(bbar[0]), .ZN(ybar[32]);
  AND2_X1 U76 ( .A1(a[1]), .A2(b[15]), .ZN(y[31]) );
  OR2_X1 U76bar ( .A1(abar[1]), .A2(bbar[15]), .ZN(ybar[31]);
  AND2_X1 U77 ( .A1(a[1]), .A2(b[14]), .ZN(y[30]) );
  OR2_X1 U77bar ( .A1(abar[1]), .A2(bbar[14]), .ZN(ybar[30]);
  AND2_X1 U78 ( .A1(b[2]), .A2(a[0]), .ZN(y[2]) );
  OR2_X1 U78bar ( .A1(bbar[2]), .A2(abar[0]), .ZN(ybar[2]);
  AND2_X1 U79 ( .A1(a[1]), .A2(b[13]), .ZN(y[29]) );
  OR2_X1 U79bar ( .A1(abar[1]), .A2(bbar[13]), .ZN(ybar[29]);
  AND2_X1 U80 ( .A1(a[1]), .A2(b[12]), .ZN(y[28]) );
  OR2_X1 U80bar ( .A1(abar[1]), .A2(bbar[12]), .ZN(ybar[28]);
  AND2_X1 U81 ( .A1(a[1]), .A2(b[11]), .ZN(y[27]) );
  OR2_X1 U81bar ( .A1(abar[1]), .A2(bbar[11]), .ZN(ybar[27]);
  AND2_X1 U82 ( .A1(a[1]), .A2(b[10]), .ZN(y[26]) );
  OR2_X1 U82bar ( .A1(abar[1]), .A2(bbar[10]), .ZN(ybar[26]);
  AND2_X1 U83 ( .A1(a[1]), .A2(b[9]), .ZN(y[25]) );
  OR2_X1 U83bar ( .A1(abar[1]), .A2(bbar[9]), .ZN(ybar[25]);
  AND2_X1 U84 ( .A1(a[15]), .A2(b[15]), .ZN(y[255]) );
  OR2_X1 U84bar ( .A1(abar[15]), .A2(bbar[15]), .ZN(ybar[255]);
  AND2_X1 U85 ( .A1(a[15]), .A2(b[14]), .ZN(y[254]) );
  OR2_X1 U85bar ( .A1(abar[15]), .A2(bbar[14]), .ZN(ybar[254]);
  AND2_X1 U86 ( .A1(a[15]), .A2(b[13]), .ZN(y[253]) );
  OR2_X1 U86bar ( .A1(abar[15]), .A2(bbar[13]), .ZN(ybar[253]);
  AND2_X1 U87 ( .A1(a[15]), .A2(b[12]), .ZN(y[252]) );
  OR2_X1 U87bar ( .A1(abar[15]), .A2(bbar[12]), .ZN(ybar[252]);
  AND2_X1 U88 ( .A1(a[15]), .A2(b[11]), .ZN(y[251]) );
  OR2_X1 U88bar ( .A1(abar[15]), .A2(bbar[11]), .ZN(ybar[251]);
  AND2_X1 U89 ( .A1(a[15]), .A2(b[10]), .ZN(y[250]) );
  OR2_X1 U89bar ( .A1(abar[15]), .A2(bbar[10]), .ZN(ybar[250]);
  AND2_X1 U90 ( .A1(a[1]), .A2(b[8]), .ZN(y[24]) );
  OR2_X1 U90bar ( .A1(abar[1]), .A2(bbar[8]), .ZN(ybar[24]);
  AND2_X1 U91 ( .A1(a[15]), .A2(b[9]), .ZN(y[249]) );
  OR2_X1 U91bar ( .A1(abar[15]), .A2(bbar[9]), .ZN(ybar[249]);
  AND2_X1 U92 ( .A1(a[15]), .A2(b[8]), .ZN(y[248]) );
  OR2_X1 U92bar ( .A1(abar[15]), .A2(bbar[8]), .ZN(ybar[248]);
  AND2_X1 U93 ( .A1(a[15]), .A2(b[7]), .ZN(y[247]) );
  OR2_X1 U93bar ( .A1(abar[15]), .A2(bbar[7]), .ZN(ybar[247]);
  AND2_X1 U94 ( .A1(a[15]), .A2(b[6]), .ZN(y[246]) );
  OR2_X1 U94bar ( .A1(abar[15]), .A2(bbar[6]), .ZN(ybar[246]);
  AND2_X1 U95 ( .A1(a[15]), .A2(b[5]), .ZN(y[245]) );
  OR2_X1 U95bar ( .A1(abar[15]), .A2(bbar[5]), .ZN(ybar[245]);
  AND2_X1 U96 ( .A1(a[15]), .A2(b[4]), .ZN(y[244]) );
  OR2_X1 U96bar ( .A1(abar[15]), .A2(bbar[4]), .ZN(ybar[244]);
  AND2_X1 U97 ( .A1(a[15]), .A2(b[3]), .ZN(y[243]) );
  OR2_X1 U97bar ( .A1(abar[15]), .A2(bbar[3]), .ZN(ybar[243]);
  AND2_X1 U98 ( .A1(a[15]), .A2(b[2]), .ZN(y[242]) );
  OR2_X1 U98bar ( .A1(abar[15]), .A2(bbar[2]), .ZN(ybar[242]);
  AND2_X1 U99 ( .A1(a[15]), .A2(b[1]), .ZN(y[241]) );
  OR2_X1 U99bar ( .A1(abar[15]), .A2(bbar[1]), .ZN(ybar[241]);
  AND2_X1 U100 ( .A1(a[15]), .A2(b[0]), .ZN(y[240]) );
  OR2_X1 U100bar ( .A1(abar[15]), .A2(bbar[0]), .ZN(ybar[240]);
  AND2_X1 U101 ( .A1(a[1]), .A2(b[7]), .ZN(y[23]) );
  OR2_X1 U101bar ( .A1(abar[1]), .A2(bbar[7]), .ZN(ybar[23]);
  AND2_X1 U102 ( .A1(a[14]), .A2(b[15]), .ZN(y[239]) );
  OR2_X1 U102bar ( .A1(abar[14]), .A2(bbar[15]), .ZN(ybar[239]);
  AND2_X1 U103 ( .A1(a[14]), .A2(b[14]), .ZN(y[238]) );
  OR2_X1 U103bar ( .A1(abar[14]), .A2(bbar[14]), .ZN(ybar[238]);
  AND2_X1 U104 ( .A1(a[14]), .A2(b[13]), .ZN(y[237]) );
  OR2_X1 U104bar ( .A1(abar[14]), .A2(bbar[13]), .ZN(ybar[237]);
  AND2_X1 U105 ( .A1(a[14]), .A2(b[12]), .ZN(y[236]) );
  OR2_X1 U105bar ( .A1(abar[14]), .A2(bbar[12]), .ZN(ybar[236]);
  AND2_X1 U106 ( .A1(a[14]), .A2(b[11]), .ZN(y[235]) );
  OR2_X1 U106bar ( .A1(abar[14]), .A2(bbar[11]), .ZN(ybar[235]);
  AND2_X1 U107 ( .A1(a[14]), .A2(b[10]), .ZN(y[234]) );
  OR2_X1 U107bar ( .A1(abar[14]), .A2(bbar[10]), .ZN(ybar[234]);
  AND2_X1 U108 ( .A1(a[14]), .A2(b[9]), .ZN(y[233]) );
  OR2_X1 U108bar ( .A1(abar[14]), .A2(bbar[9]), .ZN(ybar[233]);
  AND2_X1 U109 ( .A1(a[14]), .A2(b[8]), .ZN(y[232]) );
  OR2_X1 U109bar ( .A1(abar[14]), .A2(bbar[8]), .ZN(ybar[232]);
  AND2_X1 U110 ( .A1(a[14]), .A2(b[7]), .ZN(y[231]) );
  OR2_X1 U110bar ( .A1(abar[14]), .A2(bbar[7]), .ZN(ybar[231]);
  AND2_X1 U111 ( .A1(a[14]), .A2(b[6]), .ZN(y[230]) );
  OR2_X1 U111bar ( .A1(abar[14]), .A2(bbar[6]), .ZN(ybar[230]);
  AND2_X1 U112 ( .A1(a[1]), .A2(b[6]), .ZN(y[22]) );
  OR2_X1 U112bar ( .A1(abar[1]), .A2(bbar[6]), .ZN(ybar[22]);
  AND2_X1 U113 ( .A1(a[14]), .A2(b[5]), .ZN(y[229]) );
  OR2_X1 U113bar ( .A1(abar[14]), .A2(bbar[5]), .ZN(ybar[229]);
  AND2_X1 U114 ( .A1(a[14]), .A2(b[4]), .ZN(y[228]) );
  OR2_X1 U114bar ( .A1(abar[14]), .A2(bbar[4]), .ZN(ybar[228]);
  AND2_X1 U115 ( .A1(a[14]), .A2(b[3]), .ZN(y[227]) );
  OR2_X1 U115bar ( .A1(abar[14]), .A2(bbar[3]), .ZN(ybar[227]);
  AND2_X1 U116 ( .A1(a[14]), .A2(b[2]), .ZN(y[226]) );
  OR2_X1 U116bar ( .A1(abar[14]), .A2(bbar[2]), .ZN(ybar[226]);
  AND2_X1 U117 ( .A1(a[14]), .A2(b[1]), .ZN(y[225]) );
  OR2_X1 U117bar ( .A1(abar[14]), .A2(bbar[1]), .ZN(ybar[225]);
  AND2_X1 U118 ( .A1(a[14]), .A2(b[0]), .ZN(y[224]) );
  OR2_X1 U118bar ( .A1(abar[14]), .A2(bbar[0]), .ZN(ybar[224]);
  AND2_X1 U119 ( .A1(a[13]), .A2(b[15]), .ZN(y[223]) );
  OR2_X1 U119bar ( .A1(abar[13]), .A2(bbar[15]), .ZN(ybar[223]);
  AND2_X1 U120 ( .A1(a[13]), .A2(b[14]), .ZN(y[222]) );
  OR2_X1 U120bar ( .A1(abar[13]), .A2(bbar[14]), .ZN(ybar[222]);
  AND2_X1 U121 ( .A1(a[13]), .A2(b[13]), .ZN(y[221]) );
  OR2_X1 U121bar ( .A1(abar[13]), .A2(bbar[13]), .ZN(ybar[221]);
  AND2_X1 U122 ( .A1(a[13]), .A2(b[12]), .ZN(y[220]) );
  OR2_X1 U122bar ( .A1(abar[13]), .A2(bbar[12]), .ZN(ybar[220]);
  AND2_X1 U123 ( .A1(a[1]), .A2(b[5]), .ZN(y[21]) );
  OR2_X1 U123bar ( .A1(abar[1]), .A2(bbar[5]), .ZN(ybar[21]);
  AND2_X1 U124 ( .A1(a[13]), .A2(b[11]), .ZN(y[219]) );
  OR2_X1 U124bar ( .A1(abar[13]), .A2(bbar[11]), .ZN(ybar[219]);
  AND2_X1 U125 ( .A1(a[13]), .A2(b[10]), .ZN(y[218]) );
  OR2_X1 U125bar ( .A1(abar[13]), .A2(bbar[10]), .ZN(ybar[218]);
  AND2_X1 U126 ( .A1(a[13]), .A2(b[9]), .ZN(y[217]) );
  OR2_X1 U126bar ( .A1(abar[13]), .A2(bbar[9]), .ZN(ybar[217]);
  AND2_X1 U127 ( .A1(a[13]), .A2(b[8]), .ZN(y[216]) );
  OR2_X1 U127bar ( .A1(abar[13]), .A2(bbar[8]), .ZN(ybar[216]);
  AND2_X1 U128 ( .A1(a[13]), .A2(b[7]), .ZN(y[215]) );
  OR2_X1 U128bar ( .A1(abar[13]), .A2(bbar[7]), .ZN(ybar[215]);
  AND2_X1 U129 ( .A1(a[13]), .A2(b[6]), .ZN(y[214]) );
  OR2_X1 U129bar ( .A1(abar[13]), .A2(bbar[6]), .ZN(ybar[214]);
  AND2_X1 U130 ( .A1(a[13]), .A2(b[5]), .ZN(y[213]) );
  OR2_X1 U130bar ( .A1(abar[13]), .A2(bbar[5]), .ZN(ybar[213]);
  AND2_X1 U131 ( .A1(a[13]), .A2(b[4]), .ZN(y[212]) );
  OR2_X1 U131bar ( .A1(abar[13]), .A2(bbar[4]), .ZN(ybar[212]);
  AND2_X1 U132 ( .A1(a[13]), .A2(b[3]), .ZN(y[211]) );
  OR2_X1 U132bar ( .A1(abar[13]), .A2(bbar[3]), .ZN(ybar[211]);
  AND2_X1 U133 ( .A1(a[13]), .A2(b[2]), .ZN(y[210]) );
  OR2_X1 U133bar ( .A1(abar[13]), .A2(bbar[2]), .ZN(ybar[210]);
  AND2_X1 U134 ( .A1(a[1]), .A2(b[4]), .ZN(y[20]) );
  OR2_X1 U134bar ( .A1(abar[1]), .A2(bbar[4]), .ZN(ybar[20]);
  AND2_X1 U135 ( .A1(a[13]), .A2(b[1]), .ZN(y[209]) );
  OR2_X1 U135bar ( .A1(abar[13]), .A2(bbar[1]), .ZN(ybar[209]);
  AND2_X1 U136 ( .A1(a[13]), .A2(b[0]), .ZN(y[208]) );
  OR2_X1 U136bar ( .A1(abar[13]), .A2(bbar[0]), .ZN(ybar[208]);
  AND2_X1 U137 ( .A1(a[12]), .A2(b[15]), .ZN(y[207]) );
  OR2_X1 U137bar ( .A1(abar[12]), .A2(bbar[15]), .ZN(ybar[207]);
  AND2_X1 U138 ( .A1(a[12]), .A2(b[14]), .ZN(y[206]) );
  OR2_X1 U138bar ( .A1(abar[12]), .A2(bbar[14]), .ZN(ybar[206]);
  AND2_X1 U139 ( .A1(a[12]), .A2(b[13]), .ZN(y[205]) );
  OR2_X1 U139bar ( .A1(abar[12]), .A2(bbar[13]), .ZN(ybar[205]);
  AND2_X1 U140 ( .A1(a[12]), .A2(b[12]), .ZN(y[204]) );
  OR2_X1 U140bar ( .A1(abar[12]), .A2(bbar[12]), .ZN(ybar[204]);
  AND2_X1 U141 ( .A1(a[12]), .A2(b[11]), .ZN(y[203]) );
  OR2_X1 U141bar ( .A1(abar[12]), .A2(bbar[11]), .ZN(ybar[203]);
  AND2_X1 U142 ( .A1(a[12]), .A2(b[10]), .ZN(y[202]) );
  OR2_X1 U142bar ( .A1(abar[12]), .A2(bbar[10]), .ZN(ybar[202]);
  AND2_X1 U143 ( .A1(a[12]), .A2(b[9]), .ZN(y[201]) );
  OR2_X1 U143bar ( .A1(abar[12]), .A2(bbar[9]), .ZN(ybar[201]);
  AND2_X1 U144 ( .A1(a[12]), .A2(b[8]), .ZN(y[200]) );
  OR2_X1 U144bar ( .A1(abar[12]), .A2(bbar[8]), .ZN(ybar[200]);
  AND2_X1 U145 ( .A1(b[1]), .A2(a[0]), .ZN(y[1]) );
  OR2_X1 U145bar ( .A1(bbar[1]), .A2(abar[0]), .ZN(ybar[1]);
  AND2_X1 U146 ( .A1(a[1]), .A2(b[3]), .ZN(y[19]) );
  OR2_X1 U146bar ( .A1(abar[1]), .A2(bbar[3]), .ZN(ybar[19]);
  AND2_X1 U147 ( .A1(a[12]), .A2(b[7]), .ZN(y[199]) );
  OR2_X1 U147bar ( .A1(abar[12]), .A2(bbar[7]), .ZN(ybar[199]);
  AND2_X1 U148 ( .A1(a[12]), .A2(b[6]), .ZN(y[198]) );
  OR2_X1 U148bar ( .A1(abar[12]), .A2(bbar[6]), .ZN(ybar[198]);
  AND2_X1 U149 ( .A1(a[12]), .A2(b[5]), .ZN(y[197]) );
  OR2_X1 U149bar ( .A1(abar[12]), .A2(bbar[5]), .ZN(ybar[197]);
  AND2_X1 U150 ( .A1(a[12]), .A2(b[4]), .ZN(y[196]) );
  OR2_X1 U150bar ( .A1(abar[12]), .A2(bbar[4]), .ZN(ybar[196]);
  AND2_X1 U151 ( .A1(a[12]), .A2(b[3]), .ZN(y[195]) );
  OR2_X1 U151bar ( .A1(abar[12]), .A2(bbar[3]), .ZN(ybar[195]);
  AND2_X1 U152 ( .A1(a[12]), .A2(b[2]), .ZN(y[194]) );
  OR2_X1 U152bar ( .A1(abar[12]), .A2(bbar[2]), .ZN(ybar[194]);
  AND2_X1 U153 ( .A1(a[12]), .A2(b[1]), .ZN(y[193]) );
  OR2_X1 U153bar ( .A1(abar[12]), .A2(bbar[1]), .ZN(ybar[193]);
  AND2_X1 U154 ( .A1(a[12]), .A2(b[0]), .ZN(y[192]) );
  OR2_X1 U154bar ( .A1(abar[12]), .A2(bbar[0]), .ZN(ybar[192]);
  AND2_X1 U155 ( .A1(a[11]), .A2(b[15]), .ZN(y[191]) );
  OR2_X1 U155bar ( .A1(abar[11]), .A2(bbar[15]), .ZN(ybar[191]);
  AND2_X1 U156 ( .A1(a[11]), .A2(b[14]), .ZN(y[190]) );
  OR2_X1 U156bar ( .A1(abar[11]), .A2(bbar[14]), .ZN(ybar[190]);
  AND2_X1 U157 ( .A1(a[1]), .A2(b[2]), .ZN(y[18]) );
  OR2_X1 U157bar ( .A1(abar[1]), .A2(bbar[2]), .ZN(ybar[18]);
  AND2_X1 U158 ( .A1(a[11]), .A2(b[13]), .ZN(y[189]) );
  OR2_X1 U158bar ( .A1(abar[11]), .A2(bbar[13]), .ZN(ybar[189]);
  AND2_X1 U159 ( .A1(a[11]), .A2(b[12]), .ZN(y[188]) );
  OR2_X1 U159bar ( .A1(abar[11]), .A2(bbar[12]), .ZN(ybar[188]);
  AND2_X1 U160 ( .A1(a[11]), .A2(b[11]), .ZN(y[187]) );
  OR2_X1 U160bar ( .A1(abar[11]), .A2(bbar[11]), .ZN(ybar[187]);
  AND2_X1 U161 ( .A1(a[11]), .A2(b[10]), .ZN(y[186]) );
  OR2_X1 U161bar ( .A1(abar[11]), .A2(bbar[10]), .ZN(ybar[186]);
  AND2_X1 U162 ( .A1(a[11]), .A2(b[9]), .ZN(y[185]) );
  OR2_X1 U162bar ( .A1(abar[11]), .A2(bbar[9]), .ZN(ybar[185]);
  AND2_X1 U163 ( .A1(a[11]), .A2(b[8]), .ZN(y[184]) );
  OR2_X1 U163bar ( .A1(abar[11]), .A2(bbar[8]), .ZN(ybar[184]);
  AND2_X1 U164 ( .A1(a[11]), .A2(b[7]), .ZN(y[183]) );
  OR2_X1 U164bar ( .A1(abar[11]), .A2(bbar[7]), .ZN(ybar[183]);
  AND2_X1 U165 ( .A1(a[11]), .A2(b[6]), .ZN(y[182]) );
  OR2_X1 U165bar ( .A1(abar[11]), .A2(bbar[6]), .ZN(ybar[182]);
  AND2_X1 U166 ( .A1(a[11]), .A2(b[5]), .ZN(y[181]) );
  OR2_X1 U166bar ( .A1(abar[11]), .A2(bbar[5]), .ZN(ybar[181]);
  AND2_X1 U167 ( .A1(a[11]), .A2(b[4]), .ZN(y[180]) );
  OR2_X1 U167bar ( .A1(abar[11]), .A2(bbar[4]), .ZN(ybar[180]);
  AND2_X1 U168 ( .A1(a[1]), .A2(b[1]), .ZN(y[17]) );
  OR2_X1 U168bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[17]);
  AND2_X1 U169 ( .A1(a[11]), .A2(b[3]), .ZN(y[179]) );
  OR2_X1 U169bar ( .A1(abar[11]), .A2(bbar[3]), .ZN(ybar[179]);
  AND2_X1 U170 ( .A1(a[11]), .A2(b[2]), .ZN(y[178]) );
  OR2_X1 U170bar ( .A1(abar[11]), .A2(bbar[2]), .ZN(ybar[178]);
  AND2_X1 U171 ( .A1(a[11]), .A2(b[1]), .ZN(y[177]) );
  OR2_X1 U171bar ( .A1(abar[11]), .A2(bbar[1]), .ZN(ybar[177]);
  AND2_X1 U172 ( .A1(a[11]), .A2(b[0]), .ZN(y[176]) );
  OR2_X1 U172bar ( .A1(abar[11]), .A2(bbar[0]), .ZN(ybar[176]);
  AND2_X1 U173 ( .A1(a[10]), .A2(b[15]), .ZN(y[175]) );
  OR2_X1 U173bar ( .A1(abar[10]), .A2(bbar[15]), .ZN(ybar[175]);
  AND2_X1 U174 ( .A1(a[10]), .A2(b[14]), .ZN(y[174]) );
  OR2_X1 U174bar ( .A1(abar[10]), .A2(bbar[14]), .ZN(ybar[174]);
  AND2_X1 U175 ( .A1(a[10]), .A2(b[13]), .ZN(y[173]) );
  OR2_X1 U175bar ( .A1(abar[10]), .A2(bbar[13]), .ZN(ybar[173]);
  AND2_X1 U176 ( .A1(a[10]), .A2(b[12]), .ZN(y[172]) );
  OR2_X1 U176bar ( .A1(abar[10]), .A2(bbar[12]), .ZN(ybar[172]);
  AND2_X1 U177 ( .A1(a[10]), .A2(b[11]), .ZN(y[171]) );
  OR2_X1 U177bar ( .A1(abar[10]), .A2(bbar[11]), .ZN(ybar[171]);
  AND2_X1 U178 ( .A1(a[10]), .A2(b[10]), .ZN(y[170]) );
  OR2_X1 U178bar ( .A1(abar[10]), .A2(bbar[10]), .ZN(ybar[170]);
  AND2_X1 U179 ( .A1(a[1]), .A2(b[0]), .ZN(y[16]) );
  OR2_X1 U179bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[16]);
  AND2_X1 U180 ( .A1(a[10]), .A2(b[9]), .ZN(y[169]) );
  OR2_X1 U180bar ( .A1(abar[10]), .A2(bbar[9]), .ZN(ybar[169]);
  AND2_X1 U181 ( .A1(a[10]), .A2(b[8]), .ZN(y[168]) );
  OR2_X1 U181bar ( .A1(abar[10]), .A2(bbar[8]), .ZN(ybar[168]);
  AND2_X1 U182 ( .A1(a[10]), .A2(b[7]), .ZN(y[167]) );
  OR2_X1 U182bar ( .A1(abar[10]), .A2(bbar[7]), .ZN(ybar[167]);
  AND2_X1 U183 ( .A1(a[10]), .A2(b[6]), .ZN(y[166]) );
  OR2_X1 U183bar ( .A1(abar[10]), .A2(bbar[6]), .ZN(ybar[166]);
  AND2_X1 U184 ( .A1(a[10]), .A2(b[5]), .ZN(y[165]) );
  OR2_X1 U184bar ( .A1(abar[10]), .A2(bbar[5]), .ZN(ybar[165]);
  AND2_X1 U185 ( .A1(a[10]), .A2(b[4]), .ZN(y[164]) );
  OR2_X1 U185bar ( .A1(abar[10]), .A2(bbar[4]), .ZN(ybar[164]);
  AND2_X1 U186 ( .A1(a[10]), .A2(b[3]), .ZN(y[163]) );
  OR2_X1 U186bar ( .A1(abar[10]), .A2(bbar[3]), .ZN(ybar[163]);
  AND2_X1 U187 ( .A1(a[10]), .A2(b[2]), .ZN(y[162]) );
  OR2_X1 U187bar ( .A1(abar[10]), .A2(bbar[2]), .ZN(ybar[162]);
  AND2_X1 U188 ( .A1(a[10]), .A2(b[1]), .ZN(y[161]) );
  OR2_X1 U188bar ( .A1(abar[10]), .A2(bbar[1]), .ZN(ybar[161]);
  AND2_X1 U189 ( .A1(a[10]), .A2(b[0]), .ZN(y[160]) );
  OR2_X1 U189bar ( .A1(abar[10]), .A2(bbar[0]), .ZN(ybar[160]);
  AND2_X1 U190 ( .A1(b[15]), .A2(a[0]), .ZN(y[15]) );
  OR2_X1 U190bar ( .A1(bbar[15]), .A2(abar[0]), .ZN(ybar[15]);
  AND2_X1 U191 ( .A1(a[9]), .A2(b[15]), .ZN(y[159]) );
  OR2_X1 U191bar ( .A1(abar[9]), .A2(bbar[15]), .ZN(ybar[159]);
  AND2_X1 U192 ( .A1(a[9]), .A2(b[14]), .ZN(y[158]) );
  OR2_X1 U192bar ( .A1(abar[9]), .A2(bbar[14]), .ZN(ybar[158]);
  AND2_X1 U193 ( .A1(a[9]), .A2(b[13]), .ZN(y[157]) );
  OR2_X1 U193bar ( .A1(abar[9]), .A2(bbar[13]), .ZN(ybar[157]);
  AND2_X1 U194 ( .A1(a[9]), .A2(b[12]), .ZN(y[156]) );
  OR2_X1 U194bar ( .A1(abar[9]), .A2(bbar[12]), .ZN(ybar[156]);
  AND2_X1 U195 ( .A1(a[9]), .A2(b[11]), .ZN(y[155]) );
  OR2_X1 U195bar ( .A1(abar[9]), .A2(bbar[11]), .ZN(ybar[155]);
  AND2_X1 U196 ( .A1(a[9]), .A2(b[10]), .ZN(y[154]) );
  OR2_X1 U196bar ( .A1(abar[9]), .A2(bbar[10]), .ZN(ybar[154]);
  AND2_X1 U197 ( .A1(a[9]), .A2(b[9]), .ZN(y[153]) );
  OR2_X1 U197bar ( .A1(abar[9]), .A2(bbar[9]), .ZN(ybar[153]);
  AND2_X1 U198 ( .A1(a[9]), .A2(b[8]), .ZN(y[152]) );
  OR2_X1 U198bar ( .A1(abar[9]), .A2(bbar[8]), .ZN(ybar[152]);
  AND2_X1 U199 ( .A1(a[9]), .A2(b[7]), .ZN(y[151]) );
  OR2_X1 U199bar ( .A1(abar[9]), .A2(bbar[7]), .ZN(ybar[151]);
  AND2_X1 U200 ( .A1(a[9]), .A2(b[6]), .ZN(y[150]) );
  OR2_X1 U200bar ( .A1(abar[9]), .A2(bbar[6]), .ZN(ybar[150]);
  AND2_X1 U201 ( .A1(b[14]), .A2(a[0]), .ZN(y[14]) );
  OR2_X1 U201bar ( .A1(bbar[14]), .A2(abar[0]), .ZN(ybar[14]);
  AND2_X1 U202 ( .A1(a[9]), .A2(b[5]), .ZN(y[149]) );
  OR2_X1 U202bar ( .A1(abar[9]), .A2(bbar[5]), .ZN(ybar[149]);
  AND2_X1 U203 ( .A1(a[9]), .A2(b[4]), .ZN(y[148]) );
  OR2_X1 U203bar ( .A1(abar[9]), .A2(bbar[4]), .ZN(ybar[148]);
  AND2_X1 U204 ( .A1(a[9]), .A2(b[3]), .ZN(y[147]) );
  OR2_X1 U204bar ( .A1(abar[9]), .A2(bbar[3]), .ZN(ybar[147]);
  AND2_X1 U205 ( .A1(a[9]), .A2(b[2]), .ZN(y[146]) );
  OR2_X1 U205bar ( .A1(abar[9]), .A2(bbar[2]), .ZN(ybar[146]);
  AND2_X1 U206 ( .A1(a[9]), .A2(b[1]), .ZN(y[145]) );
  OR2_X1 U206bar ( .A1(abar[9]), .A2(bbar[1]), .ZN(ybar[145]);
  AND2_X1 U207 ( .A1(a[9]), .A2(b[0]), .ZN(y[144]) );
  OR2_X1 U207bar ( .A1(abar[9]), .A2(bbar[0]), .ZN(ybar[144]);
  AND2_X1 U208 ( .A1(a[8]), .A2(b[15]), .ZN(y[143]) );
  OR2_X1 U208bar ( .A1(abar[8]), .A2(bbar[15]), .ZN(ybar[143]);
  AND2_X1 U209 ( .A1(a[8]), .A2(b[14]), .ZN(y[142]) );
  OR2_X1 U209bar ( .A1(abar[8]), .A2(bbar[14]), .ZN(ybar[142]);
  AND2_X1 U210 ( .A1(a[8]), .A2(b[13]), .ZN(y[141]) );
  OR2_X1 U210bar ( .A1(abar[8]), .A2(bbar[13]), .ZN(ybar[141]);
  AND2_X1 U211 ( .A1(a[8]), .A2(b[12]), .ZN(y[140]) );
  OR2_X1 U211bar ( .A1(abar[8]), .A2(bbar[12]), .ZN(ybar[140]);
  AND2_X1 U212 ( .A1(b[13]), .A2(a[0]), .ZN(y[13]) );
  OR2_X1 U212bar ( .A1(bbar[13]), .A2(abar[0]), .ZN(ybar[13]);
  AND2_X1 U213 ( .A1(a[8]), .A2(b[11]), .ZN(y[139]) );
  OR2_X1 U213bar ( .A1(abar[8]), .A2(bbar[11]), .ZN(ybar[139]);
  AND2_X1 U214 ( .A1(a[8]), .A2(b[10]), .ZN(y[138]) );
  OR2_X1 U214bar ( .A1(abar[8]), .A2(bbar[10]), .ZN(ybar[138]);
  AND2_X1 U215 ( .A1(a[8]), .A2(b[9]), .ZN(y[137]) );
  OR2_X1 U215bar ( .A1(abar[8]), .A2(bbar[9]), .ZN(ybar[137]);
  AND2_X1 U216 ( .A1(a[8]), .A2(b[8]), .ZN(y[136]) );
  OR2_X1 U216bar ( .A1(abar[8]), .A2(bbar[8]), .ZN(ybar[136]);
  AND2_X1 U217 ( .A1(a[8]), .A2(b[7]), .ZN(y[135]) );
  OR2_X1 U217bar ( .A1(abar[8]), .A2(bbar[7]), .ZN(ybar[135]);
  AND2_X1 U218 ( .A1(a[8]), .A2(b[6]), .ZN(y[134]) );
  OR2_X1 U218bar ( .A1(abar[8]), .A2(bbar[6]), .ZN(ybar[134]);
  AND2_X1 U219 ( .A1(a[8]), .A2(b[5]), .ZN(y[133]) );
  OR2_X1 U219bar ( .A1(abar[8]), .A2(bbar[5]), .ZN(ybar[133]);
  AND2_X1 U220 ( .A1(a[8]), .A2(b[4]), .ZN(y[132]) );
  OR2_X1 U220bar ( .A1(abar[8]), .A2(bbar[4]), .ZN(ybar[132]);
  AND2_X1 U221 ( .A1(a[8]), .A2(b[3]), .ZN(y[131]) );
  OR2_X1 U221bar ( .A1(abar[8]), .A2(bbar[3]), .ZN(ybar[131]);
  AND2_X1 U222 ( .A1(a[8]), .A2(b[2]), .ZN(y[130]) );
  OR2_X1 U222bar ( .A1(abar[8]), .A2(bbar[2]), .ZN(ybar[130]);
  AND2_X1 U223 ( .A1(b[12]), .A2(a[0]), .ZN(y[12]) );
  OR2_X1 U223bar ( .A1(bbar[12]), .A2(abar[0]), .ZN(ybar[12]);
  AND2_X1 U224 ( .A1(a[8]), .A2(b[1]), .ZN(y[129]) );
  OR2_X1 U224bar ( .A1(abar[8]), .A2(bbar[1]), .ZN(ybar[129]);
  AND2_X1 U225 ( .A1(a[8]), .A2(b[0]), .ZN(y[128]) );
  OR2_X1 U225bar ( .A1(abar[8]), .A2(bbar[0]), .ZN(ybar[128]);
  AND2_X1 U226 ( .A1(a[7]), .A2(b[15]), .ZN(y[127]) );
  OR2_X1 U226bar ( .A1(abar[7]), .A2(bbar[15]), .ZN(ybar[127]);
  AND2_X1 U227 ( .A1(a[7]), .A2(b[14]), .ZN(y[126]) );
  OR2_X1 U227bar ( .A1(abar[7]), .A2(bbar[14]), .ZN(ybar[126]);
  AND2_X1 U228 ( .A1(a[7]), .A2(b[13]), .ZN(y[125]) );
  OR2_X1 U228bar ( .A1(abar[7]), .A2(bbar[13]), .ZN(ybar[125]);
  AND2_X1 U229 ( .A1(a[7]), .A2(b[12]), .ZN(y[124]) );
  OR2_X1 U229bar ( .A1(abar[7]), .A2(bbar[12]), .ZN(ybar[124]);
  AND2_X1 U230 ( .A1(a[7]), .A2(b[11]), .ZN(y[123]) );
  OR2_X1 U230bar ( .A1(abar[7]), .A2(bbar[11]), .ZN(ybar[123]);
  AND2_X1 U231 ( .A1(a[7]), .A2(b[10]), .ZN(y[122]) );
  OR2_X1 U231bar ( .A1(abar[7]), .A2(bbar[10]), .ZN(ybar[122]);
  AND2_X1 U232 ( .A1(a[7]), .A2(b[9]), .ZN(y[121]) );
  OR2_X1 U232bar ( .A1(abar[7]), .A2(bbar[9]), .ZN(ybar[121]);
  AND2_X1 U233 ( .A1(a[7]), .A2(b[8]), .ZN(y[120]) );
  OR2_X1 U233bar ( .A1(abar[7]), .A2(bbar[8]), .ZN(ybar[120]);
  AND2_X1 U234 ( .A1(b[11]), .A2(a[0]), .ZN(y[11]) );
  OR2_X1 U234bar ( .A1(bbar[11]), .A2(abar[0]), .ZN(ybar[11]);
  AND2_X1 U235 ( .A1(a[7]), .A2(b[7]), .ZN(y[119]) );
  OR2_X1 U235bar ( .A1(abar[7]), .A2(bbar[7]), .ZN(ybar[119]);
  AND2_X1 U236 ( .A1(a[7]), .A2(b[6]), .ZN(y[118]) );
  OR2_X1 U236bar ( .A1(abar[7]), .A2(bbar[6]), .ZN(ybar[118]);
  AND2_X1 U237 ( .A1(a[7]), .A2(b[5]), .ZN(y[117]) );
  OR2_X1 U237bar ( .A1(abar[7]), .A2(bbar[5]), .ZN(ybar[117]);
  AND2_X1 U238 ( .A1(a[7]), .A2(b[4]), .ZN(y[116]) );
  OR2_X1 U238bar ( .A1(abar[7]), .A2(bbar[4]), .ZN(ybar[116]);
  AND2_X1 U239 ( .A1(a[7]), .A2(b[3]), .ZN(y[115]) );
  OR2_X1 U239bar ( .A1(abar[7]), .A2(bbar[3]), .ZN(ybar[115]);
  AND2_X1 U240 ( .A1(a[7]), .A2(b[2]), .ZN(y[114]) );
  OR2_X1 U240bar ( .A1(abar[7]), .A2(bbar[2]), .ZN(ybar[114]);
  AND2_X1 U241 ( .A1(a[7]), .A2(b[1]), .ZN(y[113]) );
  OR2_X1 U241bar ( .A1(abar[7]), .A2(bbar[1]), .ZN(ybar[113]);
  AND2_X1 U242 ( .A1(a[7]), .A2(b[0]), .ZN(y[112]) );
  OR2_X1 U242bar ( .A1(abar[7]), .A2(bbar[0]), .ZN(ybar[112]);
  AND2_X1 U243 ( .A1(b[15]), .A2(a[6]), .ZN(y[111]) );
  OR2_X1 U243bar ( .A1(bbar[15]), .A2(abar[6]), .ZN(ybar[111]);
  AND2_X1 U244 ( .A1(b[14]), .A2(a[6]), .ZN(y[110]) );
  OR2_X1 U244bar ( .A1(bbar[14]), .A2(abar[6]), .ZN(ybar[110]);
  AND2_X1 U245 ( .A1(b[10]), .A2(a[0]), .ZN(y[10]) );
  OR2_X1 U245bar ( .A1(bbar[10]), .A2(abar[0]), .ZN(ybar[10]);
  AND2_X1 U246 ( .A1(b[13]), .A2(a[6]), .ZN(y[109]) );
  OR2_X1 U246bar ( .A1(bbar[13]), .A2(abar[6]), .ZN(ybar[109]);
  AND2_X1 U247 ( .A1(b[12]), .A2(a[6]), .ZN(y[108]) );
  OR2_X1 U247bar ( .A1(bbar[12]), .A2(abar[6]), .ZN(ybar[108]);
  AND2_X1 U248 ( .A1(b[11]), .A2(a[6]), .ZN(y[107]) );
  OR2_X1 U248bar ( .A1(bbar[11]), .A2(abar[6]), .ZN(ybar[107]);
  AND2_X1 U249 ( .A1(b[10]), .A2(a[6]), .ZN(y[106]) );
  OR2_X1 U249bar ( .A1(bbar[10]), .A2(abar[6]), .ZN(ybar[106]);
  AND2_X1 U250 ( .A1(a[6]), .A2(b[9]), .ZN(y[105]) );
  OR2_X1 U250bar ( .A1(abar[6]), .A2(bbar[9]), .ZN(ybar[105]);
  AND2_X1 U251 ( .A1(b[8]), .A2(a[6]), .ZN(y[104]) );
  OR2_X1 U251bar ( .A1(bbar[8]), .A2(abar[6]), .ZN(ybar[104]);
  AND2_X1 U252 ( .A1(b[7]), .A2(a[6]), .ZN(y[103]) );
  OR2_X1 U252bar ( .A1(bbar[7]), .A2(abar[6]), .ZN(ybar[103]);
  AND2_X1 U253 ( .A1(b[6]), .A2(a[6]), .ZN(y[102]) );
  OR2_X1 U253bar ( .A1(bbar[6]), .A2(abar[6]), .ZN(ybar[102]);
  AND2_X1 U254 ( .A1(b[5]), .A2(a[6]), .ZN(y[101]) );
  OR2_X1 U254bar ( .A1(bbar[5]), .A2(abar[6]), .ZN(ybar[101]);
  AND2_X1 U255 ( .A1(b[4]), .A2(a[6]), .ZN(y[100]) );
  OR2_X1 U255bar ( .A1(bbar[4]), .A2(abar[6]), .ZN(ybar[100]);
  AND2_X1 U256 ( .A1(b[0]), .A2(a[0]), .ZN(y[0]) );
  OR2_X1 U256bar ( .A1(bbar[0]), .A2(abar[0]), .ZN(ybar[0]);
endmodule




module decode_13 ( in, out );
  input [7:0] in;
  //input_done

  output [255:0] out;
  //output_done

  wire   [15:0] level1;
  wire   [31:0] level2;
  //wire_done

  CD2_52 cd_l1_1 ( .a(in[1]), .b(in[0]), .y(level1[3:0]) );
  CD2_51 cd_l1_2 ( .a(in[3]), .b(in[2]), .y(level1[7:4]) );
  CD2_50 cd_l1_3 ( .a(in[5]), .b(in[4]), .y(level1[11:8]) );
  CD2_49 cd_l1_4 ( .a(in[7]), .b(in[6]), .y(level1[15:12]) );
  CD4_26 cd_l2_1 ( .a(level1[7:4]), .b(level1[3:0]), .y(level2[15:0]) );
  CD4_25 cd_l2_2 ( .a(level1[15:12]), .b(level1[11:8]), .y(level2[31:16]) );
  CD16_13 cd_l3 ( .a(level2[31:16]), .b(level2[15:0]), .y(out) );
endmodule


module encode_13 ( in, out );
  input [255:0] in;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
  assign inbar[8] = ~in[8];
  assign inbar[9] = ~in[9];
  assign inbar[10] = ~in[10];
  assign inbar[11] = ~in[11];
  assign inbar[12] = ~in[12];
  assign inbar[13] = ~in[13];
  assign inbar[14] = ~in[14];
  assign inbar[15] = ~in[15];
  assign inbar[16] = ~in[16];
  assign inbar[17] = ~in[17];
  assign inbar[18] = ~in[18];
  assign inbar[19] = ~in[19];
  assign inbar[20] = ~in[20];
  assign inbar[21] = ~in[21];
  assign inbar[22] = ~in[22];
  assign inbar[23] = ~in[23];
  assign inbar[24] = ~in[24];
  assign inbar[25] = ~in[25];
  assign inbar[26] = ~in[26];
  assign inbar[27] = ~in[27];
  assign inbar[28] = ~in[28];
  assign inbar[29] = ~in[29];
  assign inbar[30] = ~in[30];
  assign inbar[31] = ~in[31];
  assign inbar[32] = ~in[32];
  assign inbar[33] = ~in[33];
  assign inbar[34] = ~in[34];
  assign inbar[35] = ~in[35];
  assign inbar[36] = ~in[36];
  assign inbar[37] = ~in[37];
  assign inbar[38] = ~in[38];
  assign inbar[39] = ~in[39];
  assign inbar[40] = ~in[40];
  assign inbar[41] = ~in[41];
  assign inbar[42] = ~in[42];
  assign inbar[43] = ~in[43];
  assign inbar[44] = ~in[44];
  assign inbar[45] = ~in[45];
  assign inbar[46] = ~in[46];
  assign inbar[47] = ~in[47];
  assign inbar[48] = ~in[48];
  assign inbar[49] = ~in[49];
  assign inbar[50] = ~in[50];
  assign inbar[51] = ~in[51];
  assign inbar[52] = ~in[52];
  assign inbar[53] = ~in[53];
  assign inbar[54] = ~in[54];
  assign inbar[55] = ~in[55];
  assign inbar[56] = ~in[56];
  assign inbar[57] = ~in[57];
  assign inbar[58] = ~in[58];
  assign inbar[59] = ~in[59];
  assign inbar[60] = ~in[60];
  assign inbar[61] = ~in[61];
  assign inbar[62] = ~in[62];
  assign inbar[63] = ~in[63];
  assign inbar[64] = ~in[64];
  assign inbar[65] = ~in[65];
  assign inbar[66] = ~in[66];
  assign inbar[67] = ~in[67];
  assign inbar[68] = ~in[68];
  assign inbar[69] = ~in[69];
  assign inbar[70] = ~in[70];
  assign inbar[71] = ~in[71];
  assign inbar[72] = ~in[72];
  assign inbar[73] = ~in[73];
  assign inbar[74] = ~in[74];
  assign inbar[75] = ~in[75];
  assign inbar[76] = ~in[76];
  assign inbar[77] = ~in[77];
  assign inbar[78] = ~in[78];
  assign inbar[79] = ~in[79];
  assign inbar[80] = ~in[80];
  assign inbar[81] = ~in[81];
  assign inbar[82] = ~in[82];
  assign inbar[83] = ~in[83];
  assign inbar[84] = ~in[84];
  assign inbar[85] = ~in[85];
  assign inbar[86] = ~in[86];
  assign inbar[87] = ~in[87];
  assign inbar[88] = ~in[88];
  assign inbar[89] = ~in[89];
  assign inbar[90] = ~in[90];
  assign inbar[91] = ~in[91];
  assign inbar[92] = ~in[92];
  assign inbar[93] = ~in[93];
  assign inbar[94] = ~in[94];
  assign inbar[95] = ~in[95];
  assign inbar[96] = ~in[96];
  assign inbar[97] = ~in[97];
  assign inbar[98] = ~in[98];
  assign inbar[99] = ~in[99];
  assign inbar[100] = ~in[100];
  assign inbar[101] = ~in[101];
  assign inbar[102] = ~in[102];
  assign inbar[103] = ~in[103];
  assign inbar[104] = ~in[104];
  assign inbar[105] = ~in[105];
  assign inbar[106] = ~in[106];
  assign inbar[107] = ~in[107];
  assign inbar[108] = ~in[108];
  assign inbar[109] = ~in[109];
  assign inbar[110] = ~in[110];
  assign inbar[111] = ~in[111];
  assign inbar[112] = ~in[112];
  assign inbar[113] = ~in[113];
  assign inbar[114] = ~in[114];
  assign inbar[115] = ~in[115];
  assign inbar[116] = ~in[116];
  assign inbar[117] = ~in[117];
  assign inbar[118] = ~in[118];
  assign inbar[119] = ~in[119];
  assign inbar[120] = ~in[120];
  assign inbar[121] = ~in[121];
  assign inbar[122] = ~in[122];
  assign inbar[123] = ~in[123];
  assign inbar[124] = ~in[124];
  assign inbar[125] = ~in[125];
  assign inbar[126] = ~in[126];
  assign inbar[127] = ~in[127];
  assign inbar[128] = ~in[128];
  assign inbar[129] = ~in[129];
  assign inbar[130] = ~in[130];
  assign inbar[131] = ~in[131];
  assign inbar[132] = ~in[132];
  assign inbar[133] = ~in[133];
  assign inbar[134] = ~in[134];
  assign inbar[135] = ~in[135];
  assign inbar[136] = ~in[136];
  assign inbar[137] = ~in[137];
  assign inbar[138] = ~in[138];
  assign inbar[139] = ~in[139];
  assign inbar[140] = ~in[140];
  assign inbar[141] = ~in[141];
  assign inbar[142] = ~in[142];
  assign inbar[143] = ~in[143];
  assign inbar[144] = ~in[144];
  assign inbar[145] = ~in[145];
  assign inbar[146] = ~in[146];
  assign inbar[147] = ~in[147];
  assign inbar[148] = ~in[148];
  assign inbar[149] = ~in[149];
  assign inbar[150] = ~in[150];
  assign inbar[151] = ~in[151];
  assign inbar[152] = ~in[152];
  assign inbar[153] = ~in[153];
  assign inbar[154] = ~in[154];
  assign inbar[155] = ~in[155];
  assign inbar[156] = ~in[156];
  assign inbar[157] = ~in[157];
  assign inbar[158] = ~in[158];
  assign inbar[159] = ~in[159];
  assign inbar[160] = ~in[160];
  assign inbar[161] = ~in[161];
  assign inbar[162] = ~in[162];
  assign inbar[163] = ~in[163];
  assign inbar[164] = ~in[164];
  assign inbar[165] = ~in[165];
  assign inbar[166] = ~in[166];
  assign inbar[167] = ~in[167];
  assign inbar[168] = ~in[168];
  assign inbar[169] = ~in[169];
  assign inbar[170] = ~in[170];
  assign inbar[171] = ~in[171];
  assign inbar[172] = ~in[172];
  assign inbar[173] = ~in[173];
  assign inbar[174] = ~in[174];
  assign inbar[175] = ~in[175];
  assign inbar[176] = ~in[176];
  assign inbar[177] = ~in[177];
  assign inbar[178] = ~in[178];
  assign inbar[179] = ~in[179];
  assign inbar[180] = ~in[180];
  assign inbar[181] = ~in[181];
  assign inbar[182] = ~in[182];
  assign inbar[183] = ~in[183];
  assign inbar[184] = ~in[184];
  assign inbar[185] = ~in[185];
  assign inbar[186] = ~in[186];
  assign inbar[187] = ~in[187];
  assign inbar[188] = ~in[188];
  assign inbar[189] = ~in[189];
  assign inbar[190] = ~in[190];
  assign inbar[191] = ~in[191];
  assign inbar[192] = ~in[192];
  assign inbar[193] = ~in[193];
  assign inbar[194] = ~in[194];
  assign inbar[195] = ~in[195];
  assign inbar[196] = ~in[196];
  assign inbar[197] = ~in[197];
  assign inbar[198] = ~in[198];
  assign inbar[199] = ~in[199];
  assign inbar[200] = ~in[200];
  assign inbar[201] = ~in[201];
  assign inbar[202] = ~in[202];
  assign inbar[203] = ~in[203];
  assign inbar[204] = ~in[204];
  assign inbar[205] = ~in[205];
  assign inbar[206] = ~in[206];
  assign inbar[207] = ~in[207];
  assign inbar[208] = ~in[208];
  assign inbar[209] = ~in[209];
  assign inbar[210] = ~in[210];
  assign inbar[211] = ~in[211];
  assign inbar[212] = ~in[212];
  assign inbar[213] = ~in[213];
  assign inbar[214] = ~in[214];
  assign inbar[215] = ~in[215];
  assign inbar[216] = ~in[216];
  assign inbar[217] = ~in[217];
  assign inbar[218] = ~in[218];
  assign inbar[219] = ~in[219];
  assign inbar[220] = ~in[220];
  assign inbar[221] = ~in[221];
  assign inbar[222] = ~in[222];
  assign inbar[223] = ~in[223];
  assign inbar[224] = ~in[224];
  assign inbar[225] = ~in[225];
  assign inbar[226] = ~in[226];
  assign inbar[227] = ~in[227];
  assign inbar[228] = ~in[228];
  assign inbar[229] = ~in[229];
  assign inbar[230] = ~in[230];
  assign inbar[231] = ~in[231];
  assign inbar[232] = ~in[232];
  assign inbar[233] = ~in[233];
  assign inbar[234] = ~in[234];
  assign inbar[235] = ~in[235];
  assign inbar[236] = ~in[236];
  assign inbar[237] = ~in[237];
  assign inbar[238] = ~in[238];
  assign inbar[239] = ~in[239];
  assign inbar[240] = ~in[240];
  assign inbar[241] = ~in[241];
  assign inbar[242] = ~in[242];
  assign inbar[243] = ~in[243];
  assign inbar[244] = ~in[244];
  assign inbar[245] = ~in[245];
  assign inbar[246] = ~in[246];
  assign inbar[247] = ~in[247];
  assign inbar[248] = ~in[248];
  assign inbar[249] = ~in[249];
  assign inbar[250] = ~in[250];
  assign inbar[251] = ~in[251];
  assign inbar[252] = ~in[252];
  assign inbar[253] = ~in[253];
  assign inbar[254] = ~in[254];
  assign inbar[255] = ~in[255];
  //input_done

  output [7:0] out;
  reg [7:0] outbar;
  //output_done

  wire   in_81, in_80, in_79, in_78, in_77, in_76, in_75, in_74, in_73, in_72,
         in_71, in_70, in_69, in_68, in_67, in_66, in_65, in_64, in_63, in_62,
         in_61, in_60, in_59, in_58, in_57, in_56, in_55, in_54, in_53, in_52,
         in_51, in_50, in_49, in_48, in_47, in_46, in_45, in_44, in_43, in_42,
         in_41, in_40, in_39, in_38, in_37, in_36, in_35, in_34, in_33, in_32,
         in_31, in_30, in_29, in_28, in_27, in_26, in_25, in_24, in_23, in_22,
         in_21, in_20, in_19, in_18, in_17, in_16, in_15, in_14, in_13, in_12,
         in_11, in_10, in_9, in_8, in_7, in_6, in_5, in_4, in_3, in_2, in_1,
         in_0, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972;
  wire in_81bar, in_80bar, in_79bar, in_78bar, in_77bar, in_76bar, in_75bar, in_74bar, in_73bar, in_72bar, in_71bar, in_70bar, in_69bar, in_68bar, in_67bar, in_66bar, in_65bar, in_64bar, in_63bar, in_62bar, in_61bar, in_60bar, in_59bar, in_58bar, in_57bar, in_56bar, in_55bar, in_54bar, in_53bar, in_52bar, in_51bar, in_50bar, in_49bar, in_48bar, in_47bar, in_46bar, in_45bar, in_44bar, in_43bar, in_42bar, in_41bar, in_40bar, in_39bar, in_38bar, in_37bar, in_36bar, in_35bar, in_34bar, in_33bar, in_32bar, in_31bar, in_30bar, in_29bar, in_28bar, in_27bar, in_26bar, in_25bar, in_24bar, in_23bar, in_22bar, in_21bar, in_20bar, in_19bar, in_18bar, in_17bar, in_16bar, in_15bar, in_14bar, in_13bar, in_12bar, in_11bar, in_10bar, in_9bar, in_8bar, in_7bar, in_6bar, in_5bar, in_4bar, in_3bar, in_2bar, in_1bar, in_0bar, n487bar, n488bar, n489bar, n490bar, n491bar, n492bar, n493bar, n494bar, n495bar, n496bar, n497bar, n498bar, n499bar, n500bar, n501bar, n502bar, n503bar, n504bar, n505bar, n506bar, n507bar, n508bar, n509bar, n510bar, n511bar, n512bar, n513bar, n514bar, n515bar, n516bar, n517bar, n518bar, n519bar, n520bar, n521bar, n522bar, n523bar, n524bar, n525bar, n526bar, n527bar, n528bar, n529bar, n530bar, n531bar, n532bar, n533bar, n534bar, n535bar, n536bar, n537bar, n538bar, n539bar, n540bar, n541bar, n542bar, n543bar, n544bar, n545bar, n546bar, n547bar, n548bar, n549bar, n550bar, n551bar, n552bar, n553bar, n554bar, n555bar, n556bar, n557bar, n558bar, n559bar, n560bar, n561bar, n562bar, n563bar, n564bar, n565bar, n566bar, n567bar, n568bar, n569bar, n570bar, n571bar, n572bar, n573bar, n574bar, n575bar, n576bar, n577bar, n578bar, n579bar, n580bar, n581bar, n582bar, n583bar, n584bar, n585bar, n586bar, n587bar, n588bar, n589bar, n590bar, n591bar, n592bar, n593bar, n594bar, n595bar, n596bar, n597bar, n598bar, n599bar, n600bar, n601bar, n602bar, n603bar, n604bar, n605bar, n606bar, n607bar, n608bar, n609bar, n610bar, n611bar, n612bar, n613bar, n614bar, n615bar, n616bar, n617bar, n618bar, n619bar, n620bar, n621bar, n622bar, n623bar, n624bar, n625bar, n626bar, n627bar, n628bar, n629bar, n630bar, n631bar, n632bar, n633bar, n634bar, n635bar, n636bar, n637bar, n638bar, n639bar, n640bar, n641bar, n642bar, n643bar, n644bar, n645bar, n646bar, n647bar, n648bar, n649bar, n650bar, n651bar, n652bar, n653bar, n654bar, n655bar, n656bar, n657bar, n658bar, n659bar, n660bar, n661bar, n662bar, n663bar, n664bar, n665bar, n666bar, n667bar, n668bar, n669bar, n670bar, n671bar, n672bar, n673bar, n674bar, n675bar, n676bar, n677bar, n678bar, n679bar, n680bar, n681bar, n682bar, n683bar, n684bar, n685bar, n686bar, n687bar, n688bar, n689bar, n690bar, n691bar, n692bar, n693bar, n694bar, n695bar, n696bar, n697bar, n698bar, n699bar, n700bar, n701bar, n702bar, n703bar, n704bar, n705bar, n706bar, n707bar, n708bar, n709bar, n710bar, n711bar, n712bar, n713bar, n714bar, n715bar, n716bar, n717bar, n718bar, n719bar, n720bar, n721bar, n722bar, n723bar, n724bar, n725bar, n726bar, n727bar, n728bar, n729bar, n730bar, n731bar, n732bar, n733bar, n734bar, n735bar, n736bar, n737bar, n738bar, n739bar, n740bar, n741bar, n742bar, n743bar, n744bar, n745bar, n746bar, n747bar, n748bar, n749bar, n750bar, n751bar, n752bar, n753bar, n754bar, n755bar, n756bar, n757bar, n758bar, n759bar, n760bar, n761bar, n762bar, n763bar, n764bar, n765bar, n766bar, n767bar, n768bar, n769bar, n770bar, n771bar, n772bar, n773bar, n774bar, n775bar, n776bar, n777bar, n778bar, n779bar, n780bar, n781bar, n782bar, n783bar, n784bar, n785bar, n786bar, n787bar, n788bar, n789bar, n790bar, n791bar, n792bar, n793bar, n794bar, n795bar, n796bar, n797bar, n798bar, n799bar, n800bar, n801bar, n802bar, n803bar, n804bar, n805bar, n806bar, n807bar, n808bar, n809bar, n810bar, n811bar, n812bar, n813bar, n814bar, n815bar, n816bar, n817bar, n818bar, n819bar, n820bar, n821bar, n822bar, n823bar, n824bar, n825bar, n826bar, n827bar, n828bar, n829bar, n830bar, n831bar, n832bar, n833bar, n834bar, n835bar, n836bar, n837bar, n838bar, n839bar, n840bar, n841bar, n842bar, n843bar, n844bar, n845bar, n846bar, n847bar, n848bar, n849bar, n850bar, n851bar, n852bar, n853bar, n854bar, n855bar, n856bar, n857bar, n858bar, n859bar, n860bar, n861bar, n862bar, n863bar, n864bar, n865bar, n866bar, n867bar, n868bar, n869bar, n870bar, n871bar, n872bar, n873bar, n874bar, n875bar, n876bar, n877bar, n878bar, n879bar, n880bar, n881bar, n882bar, n883bar, n884bar, n885bar, n886bar, n887bar, n888bar, n889bar, n890bar, n891bar, n892bar, n893bar, n894bar, n895bar, n896bar, n897bar, n898bar, n899bar, n900bar, n901bar, n902bar, n903bar, n904bar, n905bar, n906bar, n907bar, n908bar, n909bar, n910bar, n911bar, n912bar, n913bar, n914bar, n915bar, n916bar, n917bar, n918bar, n919bar, n920bar, n921bar, n922bar, n923bar, n924bar, n925bar, n926bar, n927bar, n928bar, n929bar, n930bar, n931bar, n932bar, n933bar, n934bar, n935bar, n936bar, n937bar, n938bar, n939bar, n940bar, n941bar, n942bar, n943bar, n944bar, n945bar, n946bar, n947bar, n948bar, n949bar, n950bar, n951bar, n952bar, n953bar, n954bar, n955bar, n956bar, n957bar, n958bar, n959bar, n960bar, n961bar, n962bar, n963bar, n964bar, n965bar, n966bar, n967bar, n968bar, n969bar, n970bar, n971bar, n972bar;
  //wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];

  OR2_X1 U1 ( .A1(n972), .A2(n971), .ZN(out[7]) );
  AND2_X1 U1bar ( .A1(n972bar), .A2(n971bar), .ZN(outbar[7]);
  OR2_X1 U2 ( .A1(n970), .A2(n969), .ZN(n971) );
  AND2_X1 U2bar ( .A1(n970bar), .A2(n969bar), .ZN(n971bar);
  OR2_X1 U3 ( .A1(n968), .A2(n967), .ZN(n969) );
  AND2_X1 U3bar ( .A1(n968bar), .A2(n967bar), .ZN(n969bar);
  OR2_X1 U4 ( .A1(n966), .A2(n965), .ZN(n967) );
  AND2_X1 U4bar ( .A1(n966bar), .A2(n965bar), .ZN(n967bar);
  OR2_X1 U5 ( .A1(n964), .A2(n963), .ZN(n968) );
  AND2_X1 U5bar ( .A1(n964bar), .A2(n963bar), .ZN(n968bar);
  OR2_X1 U6 ( .A1(in[116]), .A2(n962), .ZN(n963) );
  AND2_X1 U6bar ( .A1(inbar[116]), .A2(n962bar), .ZN(n963bar);
  OR2_X1 U7 ( .A1(n961), .A2(n960), .ZN(n970) );
  AND2_X1 U7bar ( .A1(n961bar), .A2(n960bar), .ZN(n970bar);
  OR2_X1 U8 ( .A1(in[150]), .A2(in[127]), .ZN(n960) );
  AND2_X1 U8bar ( .A1(inbar[150]), .A2(inbar[127]), .ZN(n960bar);
  OR2_X1 U9 ( .A1(in[160]), .A2(n959), .ZN(n961) );
  AND2_X1 U9bar ( .A1(inbar[160]), .A2(n959bar), .ZN(n961bar);
  OR2_X1 U10 ( .A1(in[252]), .A2(in[168]), .ZN(n959) );
  AND2_X1 U10bar ( .A1(inbar[252]), .A2(inbar[168]), .ZN(n959bar);
  OR2_X1 U11 ( .A1(n958), .A2(n957), .ZN(n972) );
  AND2_X1 U11bar ( .A1(n958bar), .A2(n957bar), .ZN(n972bar);
  OR2_X1 U12 ( .A1(n956), .A2(n955), .ZN(n957) );
  AND2_X1 U12bar ( .A1(n956bar), .A2(n955bar), .ZN(n957bar);
  OR2_X1 U13 ( .A1(in_17), .A2(in[96]), .ZN(n955) );
  AND2_X1 U13bar ( .A1(in_17bar), .A2(inbar[96]), .ZN(n955bar);
  OR2_X1 U14 ( .A1(in_23), .A2(n954), .ZN(n956) );
  AND2_X1 U14bar ( .A1(in_23bar), .A2(n954bar), .ZN(n956bar);
  OR2_X1 U15 ( .A1(in_31), .A2(in_26), .ZN(n954) );
  AND2_X1 U15bar ( .A1(in_31bar), .A2(in_26bar), .ZN(n954bar);
  OR2_X1 U16 ( .A1(n953), .A2(n952), .ZN(n958) );
  AND2_X1 U16bar ( .A1(n953bar), .A2(n952bar), .ZN(n958bar);
  OR2_X1 U17 ( .A1(in_58), .A2(in_4), .ZN(n952) );
  AND2_X1 U17bar ( .A1(in_58bar), .A2(in_4bar), .ZN(n952bar);
  OR2_X1 U18 ( .A1(in_59), .A2(n951), .ZN(n953) );
  AND2_X1 U18bar ( .A1(in_59bar), .A2(n951bar), .ZN(n953bar);
  OR2_X1 U19 ( .A1(in_71), .A2(in_62), .ZN(n951) );
  AND2_X1 U19bar ( .A1(in_71bar), .A2(in_62bar), .ZN(n951bar);
  OR2_X1 U20 ( .A1(n950), .A2(n949), .ZN(out[6]) );
  AND2_X1 U20bar ( .A1(n950bar), .A2(n949bar), .ZN(outbar[6]);
  OR2_X1 U21 ( .A1(n948), .A2(n947), .ZN(n949) );
  AND2_X1 U21bar ( .A1(n948bar), .A2(n947bar), .ZN(n949bar);
  OR2_X1 U22 ( .A1(n946), .A2(n945), .ZN(n947) );
  AND2_X1 U22bar ( .A1(n946bar), .A2(n945bar), .ZN(n947bar);
  OR2_X1 U23 ( .A1(n944), .A2(n943), .ZN(n945) );
  AND2_X1 U23bar ( .A1(n944bar), .A2(n943bar), .ZN(n945bar);
  OR2_X1 U24 ( .A1(n942), .A2(n941), .ZN(n946) );
  AND2_X1 U24bar ( .A1(n942bar), .A2(n941bar), .ZN(n946bar);
  OR2_X1 U25 ( .A1(in[101]), .A2(n940), .ZN(n941) );
  AND2_X1 U25bar ( .A1(inbar[101]), .A2(n940bar), .ZN(n941bar);
  OR2_X1 U26 ( .A1(n939), .A2(n938), .ZN(n948) );
  AND2_X1 U26bar ( .A1(n939bar), .A2(n938bar), .ZN(n948bar);
  OR2_X1 U27 ( .A1(in[114]), .A2(in[104]), .ZN(n938) );
  AND2_X1 U27bar ( .A1(inbar[114]), .A2(inbar[104]), .ZN(n938bar);
  OR2_X1 U28 ( .A1(in[128]), .A2(n937), .ZN(n939) );
  AND2_X1 U28bar ( .A1(inbar[128]), .A2(n937bar), .ZN(n939bar);
  OR2_X1 U29 ( .A1(in[136]), .A2(in[134]), .ZN(n937) );
  AND2_X1 U29bar ( .A1(inbar[136]), .A2(inbar[134]), .ZN(n937bar);
  OR2_X1 U30 ( .A1(n936), .A2(n935), .ZN(n950) );
  AND2_X1 U30bar ( .A1(n936bar), .A2(n935bar), .ZN(n950bar);
  OR2_X1 U31 ( .A1(n934), .A2(n933), .ZN(n935) );
  AND2_X1 U31bar ( .A1(n934bar), .A2(n933bar), .ZN(n935bar);
  OR2_X1 U32 ( .A1(in[177]), .A2(in[164]), .ZN(n933) );
  AND2_X1 U32bar ( .A1(inbar[177]), .A2(inbar[164]), .ZN(n933bar);
  OR2_X1 U33 ( .A1(in[212]), .A2(n932), .ZN(n934) );
  AND2_X1 U33bar ( .A1(inbar[212]), .A2(n932bar), .ZN(n934bar);
  OR2_X1 U34 ( .A1(in[248]), .A2(in[221]), .ZN(n932) );
  AND2_X1 U34bar ( .A1(inbar[248]), .A2(inbar[221]), .ZN(n932bar);
  OR2_X1 U35 ( .A1(n931), .A2(n930), .ZN(n936) );
  AND2_X1 U35bar ( .A1(n931bar), .A2(n930bar), .ZN(n936bar);
  OR2_X1 U36 ( .A1(in_18), .A2(in[93]), .ZN(n930) );
  AND2_X1 U36bar ( .A1(in_18bar), .A2(inbar[93]), .ZN(n930bar);
  OR2_X1 U37 ( .A1(in_31), .A2(n929), .ZN(n931) );
  AND2_X1 U37bar ( .A1(in_31bar), .A2(n929bar), .ZN(n931bar);
  OR2_X1 U38 ( .A1(in_7), .A2(in_39), .ZN(n929) );
  AND2_X1 U38bar ( .A1(in_7bar), .A2(in_39bar), .ZN(n929bar);
  OR2_X1 U39 ( .A1(n928), .A2(n927), .ZN(out[5]) );
  AND2_X1 U39bar ( .A1(n928bar), .A2(n927bar), .ZN(outbar[5]);
  OR2_X1 U40 ( .A1(n926), .A2(n925), .ZN(n927) );
  AND2_X1 U40bar ( .A1(n926bar), .A2(n925bar), .ZN(n927bar);
  OR2_X1 U41 ( .A1(n924), .A2(n923), .ZN(n925) );
  AND2_X1 U41bar ( .A1(n924bar), .A2(n923bar), .ZN(n925bar);
  OR2_X1 U42 ( .A1(n922), .A2(n921), .ZN(n923) );
  AND2_X1 U42bar ( .A1(n922bar), .A2(n921bar), .ZN(n923bar);
  OR2_X1 U43 ( .A1(n940), .A2(n920), .ZN(n924) );
  AND2_X1 U43bar ( .A1(n940bar), .A2(n920bar), .ZN(n924bar);
  OR2_X1 U44 ( .A1(in[111]), .A2(n919), .ZN(n920) );
  AND2_X1 U44bar ( .A1(inbar[111]), .A2(n919bar), .ZN(n920bar);
  OR2_X1 U45 ( .A1(n918), .A2(n917), .ZN(n940) );
  AND2_X1 U45bar ( .A1(n918bar), .A2(n917bar), .ZN(n940bar);
  OR2_X1 U46 ( .A1(n916), .A2(n915), .ZN(n917) );
  AND2_X1 U46bar ( .A1(n916bar), .A2(n915bar), .ZN(n917bar);
  OR2_X1 U47 ( .A1(n914), .A2(n913), .ZN(n915) );
  AND2_X1 U47bar ( .A1(n914bar), .A2(n913bar), .ZN(n915bar);
  OR2_X1 U48 ( .A1(in[140]), .A2(in[131]), .ZN(n913) );
  AND2_X1 U48bar ( .A1(inbar[140]), .A2(inbar[131]), .ZN(n913bar);
  OR2_X1 U49 ( .A1(in[160]), .A2(in[144]), .ZN(n914) );
  AND2_X1 U49bar ( .A1(inbar[160]), .A2(inbar[144]), .ZN(n914bar);
  OR2_X1 U50 ( .A1(n912), .A2(n911), .ZN(n916) );
  AND2_X1 U50bar ( .A1(n912bar), .A2(n911bar), .ZN(n916bar);
  OR2_X1 U51 ( .A1(in[179]), .A2(in[174]), .ZN(n911) );
  AND2_X1 U51bar ( .A1(inbar[179]), .A2(inbar[174]), .ZN(n911bar);
  OR2_X1 U52 ( .A1(in[188]), .A2(in[184]), .ZN(n912) );
  AND2_X1 U52bar ( .A1(inbar[188]), .A2(inbar[184]), .ZN(n912bar);
  OR2_X1 U53 ( .A1(n910), .A2(n909), .ZN(n918) );
  AND2_X1 U53bar ( .A1(n910bar), .A2(n909bar), .ZN(n918bar);
  OR2_X1 U54 ( .A1(n908), .A2(n907), .ZN(n909) );
  AND2_X1 U54bar ( .A1(n908bar), .A2(n907bar), .ZN(n909bar);
  OR2_X1 U55 ( .A1(in[216]), .A2(in[200]), .ZN(n907) );
  AND2_X1 U55bar ( .A1(inbar[216]), .A2(inbar[200]), .ZN(n907bar);
  OR2_X1 U56 ( .A1(in[228]), .A2(in[224]), .ZN(n908) );
  AND2_X1 U56bar ( .A1(inbar[228]), .A2(inbar[224]), .ZN(n908bar);
  OR2_X1 U57 ( .A1(n906), .A2(n905), .ZN(n910) );
  AND2_X1 U57bar ( .A1(n906bar), .A2(n905bar), .ZN(n910bar);
  OR2_X1 U58 ( .A1(in[247]), .A2(in[235]), .ZN(n905) );
  AND2_X1 U58bar ( .A1(inbar[247]), .A2(inbar[235]), .ZN(n905bar);
  OR2_X1 U59 ( .A1(in_42), .A2(in[83]), .ZN(n906) );
  AND2_X1 U59bar ( .A1(in_42bar), .A2(inbar[83]), .ZN(n906bar);
  OR2_X1 U60 ( .A1(n904), .A2(n903), .ZN(n926) );
  AND2_X1 U60bar ( .A1(n904bar), .A2(n903bar), .ZN(n926bar);
  OR2_X1 U61 ( .A1(in[166]), .A2(in[123]), .ZN(n903) );
  AND2_X1 U61bar ( .A1(inbar[166]), .A2(inbar[123]), .ZN(n903bar);
  OR2_X1 U62 ( .A1(in[170]), .A2(n902), .ZN(n904) );
  AND2_X1 U62bar ( .A1(inbar[170]), .A2(n902bar), .ZN(n904bar);
  OR2_X1 U63 ( .A1(in[194]), .A2(in[183]), .ZN(n902) );
  AND2_X1 U63bar ( .A1(inbar[194]), .A2(inbar[183]), .ZN(n902bar);
  OR2_X1 U64 ( .A1(n901), .A2(n900), .ZN(n928) );
  AND2_X1 U64bar ( .A1(n901bar), .A2(n900bar), .ZN(n928bar);
  OR2_X1 U65 ( .A1(n899), .A2(n898), .ZN(n900) );
  AND2_X1 U65bar ( .A1(n899bar), .A2(n898bar), .ZN(n900bar);
  OR2_X1 U66 ( .A1(in[241]), .A2(in[238]), .ZN(n898) );
  AND2_X1 U66bar ( .A1(inbar[241]), .A2(inbar[238]), .ZN(n898bar);
  OR2_X1 U67 ( .A1(in[250]), .A2(n897), .ZN(n899) );
  AND2_X1 U67bar ( .A1(inbar[250]), .A2(n897bar), .ZN(n899bar);
  OR2_X1 U68 ( .A1(in_24), .A2(in[84]), .ZN(n897) );
  AND2_X1 U68bar ( .A1(in_24bar), .A2(inbar[84]), .ZN(n897bar);
  OR2_X1 U69 ( .A1(n896), .A2(n895), .ZN(n901) );
  AND2_X1 U69bar ( .A1(n896bar), .A2(n895bar), .ZN(n901bar);
  OR2_X1 U70 ( .A1(in_41), .A2(in_29), .ZN(n895) );
  AND2_X1 U70bar ( .A1(in_41bar), .A2(in_29bar), .ZN(n895bar);
  OR2_X1 U71 ( .A1(in_66), .A2(n894), .ZN(n896) );
  AND2_X1 U71bar ( .A1(in_66bar), .A2(n894bar), .ZN(n896bar);
  OR2_X1 U72 ( .A1(in_76), .A2(in_71), .ZN(n894) );
  AND2_X1 U72bar ( .A1(in_76bar), .A2(in_71bar), .ZN(n894bar);
  OR2_X1 U73 ( .A1(n893), .A2(n892), .ZN(out[4]) );
  AND2_X1 U73bar ( .A1(n893bar), .A2(n892bar), .ZN(outbar[4]);
  OR2_X1 U74 ( .A1(n891), .A2(n890), .ZN(n892) );
  AND2_X1 U74bar ( .A1(n891bar), .A2(n890bar), .ZN(n892bar);
  OR2_X1 U75 ( .A1(n889), .A2(n888), .ZN(n890) );
  AND2_X1 U75bar ( .A1(n889bar), .A2(n888bar), .ZN(n890bar);
  OR2_X1 U76 ( .A1(n922), .A2(n887), .ZN(n888) );
  AND2_X1 U76bar ( .A1(n922bar), .A2(n887bar), .ZN(n888bar);
  OR2_X1 U77 ( .A1(n886), .A2(n885), .ZN(n922) );
  AND2_X1 U77bar ( .A1(n886bar), .A2(n885bar), .ZN(n922bar);
  OR2_X1 U78 ( .A1(n884), .A2(n883), .ZN(n885) );
  AND2_X1 U78bar ( .A1(n884bar), .A2(n883bar), .ZN(n885bar);
  OR2_X1 U79 ( .A1(n882), .A2(n881), .ZN(n883) );
  AND2_X1 U79bar ( .A1(n882bar), .A2(n881bar), .ZN(n883bar);
  OR2_X1 U80 ( .A1(in[118]), .A2(in[109]), .ZN(n881) );
  AND2_X1 U80bar ( .A1(inbar[118]), .A2(inbar[109]), .ZN(n881bar);
  OR2_X1 U81 ( .A1(in[139]), .A2(in[120]), .ZN(n882) );
  AND2_X1 U81bar ( .A1(inbar[139]), .A2(inbar[120]), .ZN(n882bar);
  OR2_X1 U82 ( .A1(n880), .A2(n879), .ZN(n884) );
  AND2_X1 U82bar ( .A1(n880bar), .A2(n879bar), .ZN(n884bar);
  OR2_X1 U83 ( .A1(in[198]), .A2(in[154]), .ZN(n879) );
  AND2_X1 U83bar ( .A1(inbar[198]), .A2(inbar[154]), .ZN(n879bar);
  OR2_X1 U84 ( .A1(in[210]), .A2(in[205]), .ZN(n880) );
  AND2_X1 U84bar ( .A1(inbar[210]), .A2(inbar[205]), .ZN(n880bar);
  OR2_X1 U85 ( .A1(n878), .A2(n877), .ZN(n886) );
  AND2_X1 U85bar ( .A1(n878bar), .A2(n877bar), .ZN(n886bar);
  OR2_X1 U86 ( .A1(n876), .A2(n875), .ZN(n877) );
  AND2_X1 U86bar ( .A1(n876bar), .A2(n875bar), .ZN(n877bar);
  OR2_X1 U87 ( .A1(in[219]), .A2(in[217]), .ZN(n875) );
  AND2_X1 U87bar ( .A1(inbar[219]), .A2(inbar[217]), .ZN(n875bar);
  OR2_X1 U88 ( .A1(in[86]), .A2(in[252]), .ZN(n876) );
  AND2_X1 U88bar ( .A1(inbar[86]), .A2(inbar[252]), .ZN(n876bar);
  OR2_X1 U89 ( .A1(n874), .A2(n873), .ZN(n878) );
  AND2_X1 U89bar ( .A1(n874bar), .A2(n873bar), .ZN(n878bar);
  OR2_X1 U90 ( .A1(in_40), .A2(in[91]), .ZN(n873) );
  AND2_X1 U90bar ( .A1(in_40bar), .A2(inbar[91]), .ZN(n873bar);
  OR2_X1 U91 ( .A1(in_8), .A2(in_46), .ZN(n874) );
  AND2_X1 U91bar ( .A1(in_8bar), .A2(in_46bar), .ZN(n874bar);
  OR2_X1 U92 ( .A1(n872), .A2(n871), .ZN(n889) );
  AND2_X1 U92bar ( .A1(n872bar), .A2(n871bar), .ZN(n889bar);
  OR2_X1 U93 ( .A1(in[117]), .A2(n943), .ZN(n871) );
  AND2_X1 U93bar ( .A1(inbar[117]), .A2(n943bar), .ZN(n871bar);
  OR2_X1 U94 ( .A1(n870), .A2(n869), .ZN(n943) );
  AND2_X1 U94bar ( .A1(n870bar), .A2(n869bar), .ZN(n943bar);
  OR2_X1 U95 ( .A1(n868), .A2(n867), .ZN(n869) );
  AND2_X1 U95bar ( .A1(n868bar), .A2(n867bar), .ZN(n869bar);
  OR2_X1 U96 ( .A1(n866), .A2(n865), .ZN(n867) );
  AND2_X1 U96bar ( .A1(n866bar), .A2(n865bar), .ZN(n867bar);
  OR2_X1 U97 ( .A1(n864), .A2(n863), .ZN(n865) );
  AND2_X1 U97bar ( .A1(n864bar), .A2(n863bar), .ZN(n865bar);
  OR2_X1 U98 ( .A1(in[108]), .A2(n919), .ZN(n866) );
  AND2_X1 U98bar ( .A1(inbar[108]), .A2(n919bar), .ZN(n866bar);
  OR2_X1 U99 ( .A1(n862), .A2(n861), .ZN(n919) );
  AND2_X1 U99bar ( .A1(n862bar), .A2(n861bar), .ZN(n919bar);
  OR2_X1 U100 ( .A1(n860), .A2(n859), .ZN(n861) );
  AND2_X1 U100bar ( .A1(n860bar), .A2(n859bar), .ZN(n861bar);
  OR2_X1 U101 ( .A1(n858), .A2(n857), .ZN(n859) );
  AND2_X1 U101bar ( .A1(n858bar), .A2(n857bar), .ZN(n859bar);
  OR2_X1 U102 ( .A1(in[119]), .A2(in[105]), .ZN(n857) );
  AND2_X1 U102bar ( .A1(inbar[119]), .A2(inbar[105]), .ZN(n857bar);
  OR2_X1 U103 ( .A1(in[186]), .A2(in[175]), .ZN(n858) );
  AND2_X1 U103bar ( .A1(inbar[186]), .A2(inbar[175]), .ZN(n858bar);
  OR2_X1 U104 ( .A1(n856), .A2(n855), .ZN(n860) );
  AND2_X1 U104bar ( .A1(n856bar), .A2(n855bar), .ZN(n860bar);
  OR2_X1 U105 ( .A1(in[202]), .A2(in[193]), .ZN(n855) );
  AND2_X1 U105bar ( .A1(inbar[202]), .A2(inbar[193]), .ZN(n855bar);
  OR2_X1 U106 ( .A1(in[225]), .A2(in[208]), .ZN(n856) );
  AND2_X1 U106bar ( .A1(inbar[225]), .A2(inbar[208]), .ZN(n856bar);
  OR2_X1 U107 ( .A1(n854), .A2(n853), .ZN(n862) );
  AND2_X1 U107bar ( .A1(n854bar), .A2(n853bar), .ZN(n862bar);
  OR2_X1 U108 ( .A1(n852), .A2(n851), .ZN(n853) );
  AND2_X1 U108bar ( .A1(n852bar), .A2(n851bar), .ZN(n853bar);
  OR2_X1 U109 ( .A1(in_1), .A2(in[85]), .ZN(n851) );
  AND2_X1 U109bar ( .A1(in_1bar), .A2(inbar[85]), .ZN(n851bar);
  OR2_X1 U110 ( .A1(in_23), .A2(in_19), .ZN(n852) );
  AND2_X1 U110bar ( .A1(in_23bar), .A2(in_19bar), .ZN(n852bar);
  OR2_X1 U111 ( .A1(n850), .A2(n849), .ZN(n854) );
  AND2_X1 U111bar ( .A1(n850bar), .A2(n849bar), .ZN(n854bar);
  OR2_X1 U112 ( .A1(in_43), .A2(in_33), .ZN(n849) );
  AND2_X1 U112bar ( .A1(in_43bar), .A2(in_33bar), .ZN(n849bar);
  OR2_X1 U113 ( .A1(in_63), .A2(in_44), .ZN(n850) );
  AND2_X1 U113bar ( .A1(in_63bar), .A2(in_44bar), .ZN(n850bar);
  OR2_X1 U114 ( .A1(n848), .A2(n847), .ZN(n868) );
  AND2_X1 U114bar ( .A1(n848bar), .A2(n847bar), .ZN(n868bar);
  OR2_X1 U115 ( .A1(in[141]), .A2(in[112]), .ZN(n847) );
  AND2_X1 U115bar ( .A1(inbar[141]), .A2(inbar[112]), .ZN(n847bar);
  OR2_X1 U116 ( .A1(in[147]), .A2(n846), .ZN(n848) );
  AND2_X1 U116bar ( .A1(inbar[147]), .A2(n846bar), .ZN(n848bar);
  OR2_X1 U117 ( .A1(in[181]), .A2(in[167]), .ZN(n846) );
  AND2_X1 U117bar ( .A1(inbar[181]), .A2(inbar[167]), .ZN(n846bar);
  OR2_X1 U118 ( .A1(n845), .A2(n844), .ZN(n870) );
  AND2_X1 U118bar ( .A1(n845bar), .A2(n844bar), .ZN(n870bar);
  OR2_X1 U119 ( .A1(n843), .A2(n842), .ZN(n844) );
  AND2_X1 U119bar ( .A1(n843bar), .A2(n842bar), .ZN(n844bar);
  OR2_X1 U120 ( .A1(in[229]), .A2(in[201]), .ZN(n842) );
  AND2_X1 U120bar ( .A1(inbar[229]), .A2(inbar[201]), .ZN(n842bar);
  OR2_X1 U121 ( .A1(in[237]), .A2(n841), .ZN(n843) );
  AND2_X1 U121bar ( .A1(inbar[237]), .A2(n841bar), .ZN(n843bar);
  OR2_X1 U122 ( .A1(in[94]), .A2(in[253]), .ZN(n841) );
  AND2_X1 U122bar ( .A1(inbar[94]), .A2(inbar[253]), .ZN(n841bar);
  OR2_X1 U123 ( .A1(n840), .A2(n839), .ZN(n845) );
  AND2_X1 U123bar ( .A1(n840bar), .A2(n839bar), .ZN(n845bar);
  OR2_X1 U124 ( .A1(in_21), .A2(in[96]), .ZN(n839) );
  AND2_X1 U124bar ( .A1(in_21bar), .A2(inbar[96]), .ZN(n839bar);
  OR2_X1 U125 ( .A1(in_25), .A2(n838), .ZN(n840) );
  AND2_X1 U125bar ( .A1(in_25bar), .A2(n838bar), .ZN(n840bar);
  OR2_X1 U126 ( .A1(in_81), .A2(in_45), .ZN(n838) );
  AND2_X1 U126bar ( .A1(in_81bar), .A2(in_45bar), .ZN(n838bar);
  OR2_X1 U127 ( .A1(n837), .A2(n836), .ZN(n891) );
  AND2_X1 U127bar ( .A1(n837bar), .A2(n836bar), .ZN(n891bar);
  OR2_X1 U128 ( .A1(in[142]), .A2(in[124]), .ZN(n836) );
  AND2_X1 U128bar ( .A1(inbar[142]), .A2(inbar[124]), .ZN(n836bar);
  OR2_X1 U129 ( .A1(in[150]), .A2(n835), .ZN(n837) );
  AND2_X1 U129bar ( .A1(inbar[150]), .A2(n835bar), .ZN(n837bar);
  OR2_X1 U130 ( .A1(in[172]), .A2(in[155]), .ZN(n835) );
  AND2_X1 U130bar ( .A1(inbar[172]), .A2(inbar[155]), .ZN(n835bar);
  OR2_X1 U131 ( .A1(n834), .A2(n833), .ZN(n893) );
  AND2_X1 U131bar ( .A1(n834bar), .A2(n833bar), .ZN(n893bar);
  OR2_X1 U132 ( .A1(n832), .A2(n831), .ZN(n833) );
  AND2_X1 U132bar ( .A1(n832bar), .A2(n831bar), .ZN(n833bar);
  OR2_X1 U133 ( .A1(in[196]), .A2(in[173]), .ZN(n831) );
  AND2_X1 U133bar ( .A1(inbar[196]), .A2(inbar[173]), .ZN(n831bar);
  OR2_X1 U134 ( .A1(in[222]), .A2(n830), .ZN(n832) );
  AND2_X1 U134bar ( .A1(inbar[222]), .A2(n830bar), .ZN(n832bar);
  OR2_X1 U135 ( .A1(in[227]), .A2(in[226]), .ZN(n830) );
  AND2_X1 U135bar ( .A1(inbar[227]), .A2(inbar[226]), .ZN(n830bar);
  OR2_X1 U136 ( .A1(n829), .A2(n828), .ZN(n834) );
  AND2_X1 U136bar ( .A1(n829bar), .A2(n828bar), .ZN(n834bar);
  OR2_X1 U137 ( .A1(in[249]), .A2(in[231]), .ZN(n828) );
  AND2_X1 U137bar ( .A1(inbar[249]), .A2(inbar[231]), .ZN(n828bar);
  OR2_X1 U138 ( .A1(in_28), .A2(n827), .ZN(n829) );
  AND2_X1 U138bar ( .A1(in_28bar), .A2(n827bar), .ZN(n829bar);
  OR2_X1 U139 ( .A1(in_52), .A2(in_47), .ZN(n827) );
  AND2_X1 U139bar ( .A1(in_52bar), .A2(in_47bar), .ZN(n827bar);
  OR2_X1 U140 ( .A1(n826), .A2(n825), .ZN(out[3]) );
  AND2_X1 U140bar ( .A1(n826bar), .A2(n825bar), .ZN(outbar[3]);
  OR2_X1 U141 ( .A1(n824), .A2(n823), .ZN(n825) );
  AND2_X1 U141bar ( .A1(n824bar), .A2(n823bar), .ZN(n825bar);
  OR2_X1 U142 ( .A1(n822), .A2(n821), .ZN(n823) );
  AND2_X1 U142bar ( .A1(n822bar), .A2(n821bar), .ZN(n823bar);
  OR2_X1 U143 ( .A1(n820), .A2(n819), .ZN(n821) );
  AND2_X1 U143bar ( .A1(n820bar), .A2(n819bar), .ZN(n821bar);
  OR2_X1 U144 ( .A1(n964), .A2(n818), .ZN(n822) );
  AND2_X1 U144bar ( .A1(n964bar), .A2(n818bar), .ZN(n822bar);
  OR2_X1 U145 ( .A1(in[118]), .A2(n817), .ZN(n818) );
  AND2_X1 U145bar ( .A1(inbar[118]), .A2(n817bar), .ZN(n818bar);
  OR2_X1 U146 ( .A1(n816), .A2(n815), .ZN(n964) );
  AND2_X1 U146bar ( .A1(n816bar), .A2(n815bar), .ZN(n964bar);
  OR2_X1 U147 ( .A1(n814), .A2(n813), .ZN(n815) );
  AND2_X1 U147bar ( .A1(n814bar), .A2(n813bar), .ZN(n815bar);
  OR2_X1 U148 ( .A1(n812), .A2(n811), .ZN(n813) );
  AND2_X1 U148bar ( .A1(n812bar), .A2(n811bar), .ZN(n813bar);
  OR2_X1 U149 ( .A1(in[122]), .A2(in[111]), .ZN(n811) );
  AND2_X1 U149bar ( .A1(inbar[122]), .A2(inbar[111]), .ZN(n811bar);
  OR2_X1 U150 ( .A1(in[154]), .A2(in[151]), .ZN(n812) );
  AND2_X1 U150bar ( .A1(inbar[154]), .A2(inbar[151]), .ZN(n812bar);
  OR2_X1 U151 ( .A1(n810), .A2(n809), .ZN(n814) );
  AND2_X1 U151bar ( .A1(n810bar), .A2(n809bar), .ZN(n814bar);
  OR2_X1 U152 ( .A1(in[187]), .A2(in[177]), .ZN(n809) );
  AND2_X1 U152bar ( .A1(inbar[187]), .A2(inbar[177]), .ZN(n809bar);
  OR2_X1 U153 ( .A1(in[200]), .A2(in[192]), .ZN(n810) );
  AND2_X1 U153bar ( .A1(inbar[200]), .A2(inbar[192]), .ZN(n810bar);
  OR2_X1 U154 ( .A1(n808), .A2(n807), .ZN(n816) );
  AND2_X1 U154bar ( .A1(n808bar), .A2(n807bar), .ZN(n816bar);
  OR2_X1 U155 ( .A1(n806), .A2(n805), .ZN(n807) );
  AND2_X1 U155bar ( .A1(n806bar), .A2(n805bar), .ZN(n807bar);
  OR2_X1 U156 ( .A1(in[225]), .A2(in[207]), .ZN(n805) );
  AND2_X1 U156bar ( .A1(inbar[225]), .A2(inbar[207]), .ZN(n805bar);
  OR2_X1 U157 ( .A1(in[98]), .A2(in[226]), .ZN(n806) );
  AND2_X1 U157bar ( .A1(inbar[98]), .A2(inbar[226]), .ZN(n806bar);
  OR2_X1 U158 ( .A1(n804), .A2(n803), .ZN(n808) );
  AND2_X1 U158bar ( .A1(n804bar), .A2(n803bar), .ZN(n808bar);
  OR2_X1 U159 ( .A1(in_20), .A2(in_16), .ZN(n803) );
  AND2_X1 U159bar ( .A1(in_20bar), .A2(in_16bar), .ZN(n803bar);
  OR2_X1 U160 ( .A1(in_55), .A2(in_45), .ZN(n804) );
  AND2_X1 U160bar ( .A1(in_55bar), .A2(in_45bar), .ZN(n804bar);
  OR2_X1 U161 ( .A1(n802), .A2(n801), .ZN(n824) );
  AND2_X1 U161bar ( .A1(n802bar), .A2(n801bar), .ZN(n824bar);
  OR2_X1 U162 ( .A1(in[162]), .A2(in[149]), .ZN(n801) );
  AND2_X1 U162bar ( .A1(inbar[162]), .A2(inbar[149]), .ZN(n801bar);
  OR2_X1 U163 ( .A1(in[163]), .A2(n800), .ZN(n802) );
  AND2_X1 U163bar ( .A1(inbar[163]), .A2(n800bar), .ZN(n802bar);
  OR2_X1 U164 ( .A1(in[191]), .A2(in[189]), .ZN(n800) );
  AND2_X1 U164bar ( .A1(inbar[191]), .A2(inbar[189]), .ZN(n800bar);
  OR2_X1 U165 ( .A1(n799), .A2(n798), .ZN(n826) );
  AND2_X1 U165bar ( .A1(n799bar), .A2(n798bar), .ZN(n826bar);
  OR2_X1 U166 ( .A1(n797), .A2(n796), .ZN(n798) );
  AND2_X1 U166bar ( .A1(n797bar), .A2(n796bar), .ZN(n798bar);
  OR2_X1 U167 ( .A1(in[212]), .A2(in[193]), .ZN(n796) );
  AND2_X1 U167bar ( .A1(inbar[212]), .A2(inbar[193]), .ZN(n796bar);
  OR2_X1 U168 ( .A1(in[238]), .A2(n795), .ZN(n797) );
  AND2_X1 U168bar ( .A1(inbar[238]), .A2(n795bar), .ZN(n797bar);
  OR2_X1 U169 ( .A1(in[88]), .A2(in[247]), .ZN(n795) );
  AND2_X1 U169bar ( .A1(inbar[88]), .A2(inbar[247]), .ZN(n795bar);
  OR2_X1 U170 ( .A1(n794), .A2(n793), .ZN(n799) );
  AND2_X1 U170bar ( .A1(n794bar), .A2(n793bar), .ZN(n799bar);
  OR2_X1 U171 ( .A1(in[94]), .A2(in[92]), .ZN(n793) );
  AND2_X1 U171bar ( .A1(inbar[94]), .A2(inbar[92]), .ZN(n793bar);
  OR2_X1 U172 ( .A1(in_52), .A2(n792), .ZN(n794) );
  AND2_X1 U172bar ( .A1(in_52bar), .A2(n792bar), .ZN(n794bar);
  OR2_X1 U173 ( .A1(in_70), .A2(in_67), .ZN(n792) );
  AND2_X1 U173bar ( .A1(in_70bar), .A2(in_67bar), .ZN(n792bar);
  OR2_X1 U174 ( .A1(n791), .A2(n790), .ZN(out[2]) );
  AND2_X1 U174bar ( .A1(n791bar), .A2(n790bar), .ZN(outbar[2]);
  OR2_X1 U175 ( .A1(n789), .A2(n788), .ZN(n790) );
  AND2_X1 U175bar ( .A1(n789bar), .A2(n788bar), .ZN(n790bar);
  OR2_X1 U176 ( .A1(n787), .A2(n786), .ZN(n788) );
  AND2_X1 U176bar ( .A1(n787bar), .A2(n786bar), .ZN(n788bar);
  OR2_X1 U177 ( .A1(n819), .A2(n785), .ZN(n786) );
  AND2_X1 U177bar ( .A1(n819bar), .A2(n785bar), .ZN(n786bar);
  OR2_X1 U178 ( .A1(n784), .A2(n783), .ZN(n819) );
  AND2_X1 U178bar ( .A1(n784bar), .A2(n783bar), .ZN(n819bar);
  OR2_X1 U179 ( .A1(n782), .A2(n781), .ZN(n783) );
  AND2_X1 U179bar ( .A1(n782bar), .A2(n781bar), .ZN(n783bar);
  OR2_X1 U180 ( .A1(n780), .A2(n779), .ZN(n781) );
  AND2_X1 U180bar ( .A1(n780bar), .A2(n779bar), .ZN(n781bar);
  OR2_X1 U181 ( .A1(n962), .A2(n778), .ZN(n779) );
  AND2_X1 U181bar ( .A1(n962bar), .A2(n778bar), .ZN(n779bar);
  OR2_X1 U182 ( .A1(n777), .A2(n776), .ZN(n962) );
  AND2_X1 U182bar ( .A1(n777bar), .A2(n776bar), .ZN(n962bar);
  OR2_X1 U183 ( .A1(n775), .A2(n774), .ZN(n776) );
  AND2_X1 U183bar ( .A1(n775bar), .A2(n774bar), .ZN(n776bar);
  OR2_X1 U184 ( .A1(n773), .A2(n772), .ZN(n774) );
  AND2_X1 U184bar ( .A1(n773bar), .A2(n772bar), .ZN(n774bar);
  OR2_X1 U185 ( .A1(in[131]), .A2(in[120]), .ZN(n772) );
  AND2_X1 U185bar ( .A1(inbar[131]), .A2(inbar[120]), .ZN(n772bar);
  OR2_X1 U186 ( .A1(in[153]), .A2(in[147]), .ZN(n773) );
  AND2_X1 U186bar ( .A1(inbar[153]), .A2(inbar[147]), .ZN(n773bar);
  OR2_X1 U187 ( .A1(n771), .A2(n770), .ZN(n775) );
  AND2_X1 U187bar ( .A1(n771bar), .A2(n770bar), .ZN(n775bar);
  OR2_X1 U188 ( .A1(in[170]), .A2(in[156]), .ZN(n770) );
  AND2_X1 U188bar ( .A1(inbar[170]), .A2(inbar[156]), .ZN(n770bar);
  OR2_X1 U189 ( .A1(in[223]), .A2(in[190]), .ZN(n771) );
  AND2_X1 U189bar ( .A1(inbar[223]), .A2(inbar[190]), .ZN(n771bar);
  OR2_X1 U190 ( .A1(n769), .A2(n768), .ZN(n777) );
  AND2_X1 U190bar ( .A1(n769bar), .A2(n768bar), .ZN(n777bar);
  OR2_X1 U191 ( .A1(n767), .A2(n766), .ZN(n768) );
  AND2_X1 U191bar ( .A1(n767bar), .A2(n766bar), .ZN(n768bar);
  OR2_X1 U192 ( .A1(in[236]), .A2(in[230]), .ZN(n766) );
  AND2_X1 U192bar ( .A1(inbar[236]), .A2(inbar[230]), .ZN(n766bar);
  OR2_X1 U193 ( .A1(in[85]), .A2(in[240]), .ZN(n767) );
  AND2_X1 U193bar ( .A1(inbar[85]), .A2(inbar[240]), .ZN(n767bar);
  OR2_X1 U194 ( .A1(n765), .A2(n764), .ZN(n769) );
  AND2_X1 U194bar ( .A1(n765bar), .A2(n764bar), .ZN(n769bar);
  OR2_X1 U195 ( .A1(in_12), .A2(in[90]), .ZN(n764) );
  AND2_X1 U195bar ( .A1(in_12bar), .A2(inbar[90]), .ZN(n764bar);
  OR2_X1 U196 ( .A1(in_39), .A2(in_28), .ZN(n765) );
  AND2_X1 U196bar ( .A1(in_39bar), .A2(in_28bar), .ZN(n765bar);
  OR2_X1 U197 ( .A1(in[109]), .A2(n763), .ZN(n780) );
  AND2_X1 U197bar ( .A1(inbar[109]), .A2(n763bar), .ZN(n780bar);
  OR2_X1 U198 ( .A1(n762), .A2(n761), .ZN(n782) );
  AND2_X1 U198bar ( .A1(n762bar), .A2(n761bar), .ZN(n782bar);
  OR2_X1 U199 ( .A1(in[138]), .A2(in[129]), .ZN(n761) );
  AND2_X1 U199bar ( .A1(inbar[138]), .A2(inbar[129]), .ZN(n761bar);
  OR2_X1 U200 ( .A1(in[157]), .A2(n760), .ZN(n762) );
  AND2_X1 U200bar ( .A1(inbar[157]), .A2(n760bar), .ZN(n762bar);
  OR2_X1 U201 ( .A1(in[182]), .A2(in[167]), .ZN(n760) );
  AND2_X1 U201bar ( .A1(inbar[182]), .A2(inbar[167]), .ZN(n760bar);
  OR2_X1 U202 ( .A1(n759), .A2(n758), .ZN(n784) );
  AND2_X1 U202bar ( .A1(n759bar), .A2(n758bar), .ZN(n784bar);
  OR2_X1 U203 ( .A1(n757), .A2(n756), .ZN(n758) );
  AND2_X1 U203bar ( .A1(n757bar), .A2(n756bar), .ZN(n758bar);
  OR2_X1 U204 ( .A1(in[195]), .A2(in[184]), .ZN(n756) );
  AND2_X1 U204bar ( .A1(inbar[195]), .A2(inbar[184]), .ZN(n756bar);
  OR2_X1 U205 ( .A1(in[196]), .A2(n755), .ZN(n757) );
  AND2_X1 U205bar ( .A1(inbar[196]), .A2(n755bar), .ZN(n757bar);
  OR2_X1 U206 ( .A1(in[215]), .A2(in[209]), .ZN(n755) );
  AND2_X1 U206bar ( .A1(inbar[215]), .A2(inbar[209]), .ZN(n755bar);
  OR2_X1 U207 ( .A1(n754), .A2(n753), .ZN(n759) );
  AND2_X1 U207bar ( .A1(n754bar), .A2(n753bar), .ZN(n759bar);
  OR2_X1 U208 ( .A1(in[93]), .A2(in[233]), .ZN(n753) );
  AND2_X1 U208bar ( .A1(inbar[93]), .A2(inbar[233]), .ZN(n753bar);
  OR2_X1 U209 ( .A1(in_1), .A2(n752), .ZN(n754) );
  AND2_X1 U209bar ( .A1(in_1bar), .A2(n752bar), .ZN(n754bar);
  OR2_X1 U210 ( .A1(in_69), .A2(in_66), .ZN(n752) );
  AND2_X1 U210bar ( .A1(in_69bar), .A2(in_66bar), .ZN(n752bar);
  OR2_X1 U211 ( .A1(n966), .A2(n751), .ZN(n787) );
  AND2_X1 U211bar ( .A1(n966bar), .A2(n751bar), .ZN(n787bar);
  OR2_X1 U212 ( .A1(in[134]), .A2(n750), .ZN(n751) );
  AND2_X1 U212bar ( .A1(inbar[134]), .A2(n750bar), .ZN(n751bar);
  OR2_X1 U213 ( .A1(n749), .A2(n748), .ZN(n966) );
  AND2_X1 U213bar ( .A1(n749bar), .A2(n748bar), .ZN(n966bar);
  OR2_X1 U214 ( .A1(n747), .A2(n746), .ZN(n748) );
  AND2_X1 U214bar ( .A1(n747bar), .A2(n746bar), .ZN(n748bar);
  OR2_X1 U215 ( .A1(n745), .A2(n744), .ZN(n746) );
  AND2_X1 U215bar ( .A1(n745bar), .A2(n744bar), .ZN(n746bar);
  OR2_X1 U216 ( .A1(in[136]), .A2(in[121]), .ZN(n744) );
  AND2_X1 U216bar ( .A1(inbar[136]), .A2(inbar[121]), .ZN(n744bar);
  OR2_X1 U217 ( .A1(in[186]), .A2(in[174]), .ZN(n745) );
  AND2_X1 U217bar ( .A1(inbar[186]), .A2(inbar[174]), .ZN(n745bar);
  OR2_X1 U218 ( .A1(n743), .A2(n742), .ZN(n747) );
  AND2_X1 U218bar ( .A1(n743bar), .A2(n742bar), .ZN(n747bar);
  OR2_X1 U219 ( .A1(in[198]), .A2(in[197]), .ZN(n742) );
  AND2_X1 U219bar ( .A1(inbar[198]), .A2(inbar[197]), .ZN(n742bar);
  OR2_X1 U220 ( .A1(in[214]), .A2(in[199]), .ZN(n743) );
  AND2_X1 U220bar ( .A1(inbar[214]), .A2(inbar[199]), .ZN(n743bar);
  OR2_X1 U221 ( .A1(n741), .A2(n740), .ZN(n749) );
  AND2_X1 U221bar ( .A1(n741bar), .A2(n740bar), .ZN(n749bar);
  OR2_X1 U222 ( .A1(n739), .A2(n738), .ZN(n740) );
  AND2_X1 U222bar ( .A1(n739bar), .A2(n738bar), .ZN(n740bar);
  OR2_X1 U223 ( .A1(in[231]), .A2(in[220]), .ZN(n738) );
  AND2_X1 U223bar ( .A1(inbar[231]), .A2(inbar[220]), .ZN(n738bar);
  OR2_X1 U224 ( .A1(in_25), .A2(in[245]), .ZN(n739) );
  AND2_X1 U224bar ( .A1(in_25bar), .A2(inbar[245]), .ZN(n739bar);
  OR2_X1 U225 ( .A1(n737), .A2(n736), .ZN(n741) );
  AND2_X1 U225bar ( .A1(n737bar), .A2(n736bar), .ZN(n741bar);
  OR2_X1 U226 ( .A1(in_53), .A2(in_29), .ZN(n736) );
  AND2_X1 U226bar ( .A1(in_53bar), .A2(in_29bar), .ZN(n736bar);
  OR2_X1 U227 ( .A1(in_79), .A2(in_74), .ZN(n737) );
  AND2_X1 U227bar ( .A1(in_79bar), .A2(in_74bar), .ZN(n737bar);
  OR2_X1 U228 ( .A1(n735), .A2(n734), .ZN(n789) );
  AND2_X1 U228bar ( .A1(n735bar), .A2(n734bar), .ZN(n789bar);
  OR2_X1 U229 ( .A1(in[152]), .A2(in[140]), .ZN(n734) );
  AND2_X1 U229bar ( .A1(inbar[152]), .A2(inbar[140]), .ZN(n734bar);
  OR2_X1 U230 ( .A1(in[155]), .A2(n733), .ZN(n735) );
  AND2_X1 U230bar ( .A1(inbar[155]), .A2(n733bar), .ZN(n735bar);
  OR2_X1 U231 ( .A1(in[166]), .A2(in[165]), .ZN(n733) );
  AND2_X1 U231bar ( .A1(inbar[166]), .A2(inbar[165]), .ZN(n733bar);
  OR2_X1 U232 ( .A1(n732), .A2(n731), .ZN(n791) );
  AND2_X1 U232bar ( .A1(n732bar), .A2(n731bar), .ZN(n791bar);
  OR2_X1 U233 ( .A1(n730), .A2(n729), .ZN(n731) );
  AND2_X1 U233bar ( .A1(n730bar), .A2(n729bar), .ZN(n731bar);
  OR2_X1 U234 ( .A1(in[202]), .A2(in[185]), .ZN(n729) );
  AND2_X1 U234bar ( .A1(inbar[202]), .A2(inbar[185]), .ZN(n729bar);
  OR2_X1 U235 ( .A1(in[211]), .A2(n728), .ZN(n730) );
  AND2_X1 U235bar ( .A1(inbar[211]), .A2(n728bar), .ZN(n730bar);
  OR2_X1 U236 ( .A1(in[255]), .A2(in[253]), .ZN(n728) );
  AND2_X1 U236bar ( .A1(inbar[255]), .A2(inbar[253]), .ZN(n728bar);
  OR2_X1 U237 ( .A1(n727), .A2(n726), .ZN(n732) );
  AND2_X1 U237bar ( .A1(n727bar), .A2(n726bar), .ZN(n732bar);
  OR2_X1 U238 ( .A1(in_35), .A2(in_15), .ZN(n726) );
  AND2_X1 U238bar ( .A1(in_35bar), .A2(in_15bar), .ZN(n726bar);
  OR2_X1 U239 ( .A1(in_36), .A2(n725), .ZN(n727) );
  AND2_X1 U239bar ( .A1(in_36bar), .A2(n725bar), .ZN(n727bar);
  OR2_X1 U240 ( .A1(in_48), .A2(in_40), .ZN(n725) );
  AND2_X1 U240bar ( .A1(in_48bar), .A2(in_40bar), .ZN(n725bar);
  OR2_X1 U241 ( .A1(n724), .A2(n723), .ZN(out[1]) );
  AND2_X1 U241bar ( .A1(n724bar), .A2(n723bar), .ZN(outbar[1]);
  OR2_X1 U242 ( .A1(n722), .A2(n721), .ZN(n723) );
  AND2_X1 U242bar ( .A1(n722bar), .A2(n721bar), .ZN(n723bar);
  OR2_X1 U243 ( .A1(n720), .A2(n719), .ZN(n721) );
  AND2_X1 U243bar ( .A1(n720bar), .A2(n719bar), .ZN(n721bar);
  OR2_X1 U244 ( .A1(n921), .A2(n887), .ZN(n719) );
  AND2_X1 U244bar ( .A1(n921bar), .A2(n887bar), .ZN(n719bar);
  OR2_X1 U245 ( .A1(n718), .A2(n717), .ZN(n887) );
  AND2_X1 U245bar ( .A1(n718bar), .A2(n717bar), .ZN(n887bar);
  OR2_X1 U246 ( .A1(n716), .A2(n715), .ZN(n717) );
  AND2_X1 U246bar ( .A1(n716bar), .A2(n715bar), .ZN(n717bar);
  OR2_X1 U247 ( .A1(n714), .A2(n713), .ZN(n715) );
  AND2_X1 U247bar ( .A1(n714bar), .A2(n713bar), .ZN(n715bar);
  OR2_X1 U248 ( .A1(in[116]), .A2(in[110]), .ZN(n713) );
  AND2_X1 U248bar ( .A1(inbar[116]), .A2(inbar[110]), .ZN(n713bar);
  OR2_X1 U249 ( .A1(in[133]), .A2(in[130]), .ZN(n714) );
  AND2_X1 U249bar ( .A1(inbar[133]), .A2(inbar[130]), .ZN(n714bar);
  OR2_X1 U250 ( .A1(n712), .A2(n711), .ZN(n716) );
  AND2_X1 U250bar ( .A1(n712bar), .A2(n711bar), .ZN(n716bar);
  OR2_X1 U251 ( .A1(in[203]), .A2(in[135]), .ZN(n711) );
  AND2_X1 U251bar ( .A1(inbar[203]), .A2(inbar[135]), .ZN(n711bar);
  OR2_X1 U252 ( .A1(in[232]), .A2(in[223]), .ZN(n712) );
  AND2_X1 U252bar ( .A1(inbar[232]), .A2(inbar[223]), .ZN(n712bar);
  OR2_X1 U253 ( .A1(n710), .A2(n709), .ZN(n718) );
  AND2_X1 U253bar ( .A1(n710bar), .A2(n709bar), .ZN(n718bar);
  OR2_X1 U254 ( .A1(n708), .A2(n707), .ZN(n709) );
  AND2_X1 U254bar ( .A1(n708bar), .A2(n707bar), .ZN(n709bar);
  OR2_X1 U255 ( .A1(in[255]), .A2(in[233]), .ZN(n707) );
  AND2_X1 U255bar ( .A1(inbar[255]), .A2(inbar[233]), .ZN(n707bar);
  OR2_X1 U256 ( .A1(in_53), .A2(in_34), .ZN(n708) );
  AND2_X1 U256bar ( .A1(in_53bar), .A2(in_34bar), .ZN(n708bar);
  OR2_X1 U257 ( .A1(n706), .A2(n705), .ZN(n710) );
  AND2_X1 U257bar ( .A1(n706bar), .A2(n705bar), .ZN(n710bar);
  OR2_X1 U258 ( .A1(in_57), .A2(in_55), .ZN(n705) );
  AND2_X1 U258bar ( .A1(in_57bar), .A2(in_55bar), .ZN(n705bar);
  OR2_X1 U259 ( .A1(in_68), .A2(in_67), .ZN(n706) );
  AND2_X1 U259bar ( .A1(in_68bar), .A2(in_67bar), .ZN(n706bar);
  OR2_X1 U260 ( .A1(n704), .A2(n703), .ZN(n921) );
  AND2_X1 U260bar ( .A1(n704bar), .A2(n703bar), .ZN(n921bar);
  OR2_X1 U261 ( .A1(n702), .A2(n701), .ZN(n703) );
  AND2_X1 U261bar ( .A1(n702bar), .A2(n701bar), .ZN(n703bar);
  OR2_X1 U262 ( .A1(n700), .A2(n699), .ZN(n701) );
  AND2_X1 U262bar ( .A1(n700bar), .A2(n699bar), .ZN(n701bar);
  OR2_X1 U263 ( .A1(n944), .A2(n872), .ZN(n699) );
  AND2_X1 U263bar ( .A1(n944bar), .A2(n872bar), .ZN(n699bar);
  OR2_X1 U264 ( .A1(n698), .A2(n697), .ZN(n872) );
  AND2_X1 U264bar ( .A1(n698bar), .A2(n697bar), .ZN(n872bar);
  OR2_X1 U265 ( .A1(n696), .A2(n695), .ZN(n697) );
  AND2_X1 U265bar ( .A1(n696bar), .A2(n695bar), .ZN(n697bar);
  OR2_X1 U266 ( .A1(n694), .A2(n693), .ZN(n695) );
  AND2_X1 U266bar ( .A1(n694bar), .A2(n693bar), .ZN(n695bar);
  OR2_X1 U267 ( .A1(in[121]), .A2(in[102]), .ZN(n693) );
  AND2_X1 U267bar ( .A1(inbar[121]), .A2(inbar[102]), .ZN(n693bar);
  OR2_X1 U268 ( .A1(in[162]), .A2(in[161]), .ZN(n694) );
  AND2_X1 U268bar ( .A1(inbar[162]), .A2(inbar[161]), .ZN(n694bar);
  OR2_X1 U269 ( .A1(n692), .A2(n691), .ZN(n696) );
  AND2_X1 U269bar ( .A1(n692bar), .A2(n691bar), .ZN(n696bar);
  OR2_X1 U270 ( .A1(in[192]), .A2(in[178]), .ZN(n691) );
  AND2_X1 U270bar ( .A1(inbar[192]), .A2(inbar[178]), .ZN(n691bar);
  OR2_X1 U271 ( .A1(in[244]), .A2(in[209]), .ZN(n692) );
  AND2_X1 U271bar ( .A1(inbar[244]), .A2(inbar[209]), .ZN(n692bar);
  OR2_X1 U272 ( .A1(n690), .A2(n689), .ZN(n698) );
  AND2_X1 U272bar ( .A1(n690bar), .A2(n689bar), .ZN(n698bar);
  OR2_X1 U273 ( .A1(n688), .A2(n687), .ZN(n689) );
  AND2_X1 U273bar ( .A1(n688bar), .A2(n687bar), .ZN(n689bar);
  OR2_X1 U274 ( .A1(in[90]), .A2(in[254]), .ZN(n687) );
  AND2_X1 U274bar ( .A1(inbar[90]), .A2(inbar[254]), .ZN(n687bar);
  OR2_X1 U275 ( .A1(in_36), .A2(in_32), .ZN(n688) );
  AND2_X1 U275bar ( .A1(in_36bar), .A2(in_32bar), .ZN(n688bar);
  OR2_X1 U276 ( .A1(n686), .A2(n685), .ZN(n690) );
  AND2_X1 U276bar ( .A1(n686bar), .A2(n685bar), .ZN(n690bar);
  OR2_X1 U277 ( .A1(in_62), .A2(in_37), .ZN(n685) );
  AND2_X1 U277bar ( .A1(in_62bar), .A2(in_37bar), .ZN(n685bar);
  OR2_X1 U278 ( .A1(in_75), .A2(in_73), .ZN(n686) );
  AND2_X1 U278bar ( .A1(in_75bar), .A2(in_73bar), .ZN(n686bar);
  OR2_X1 U279 ( .A1(n684), .A2(n683), .ZN(n944) );
  AND2_X1 U279bar ( .A1(n684bar), .A2(n683bar), .ZN(n944bar);
  OR2_X1 U280 ( .A1(n682), .A2(n681), .ZN(n683) );
  AND2_X1 U280bar ( .A1(n682bar), .A2(n681bar), .ZN(n683bar);
  OR2_X1 U281 ( .A1(n680), .A2(n679), .ZN(n681) );
  AND2_X1 U281bar ( .A1(n680bar), .A2(n679bar), .ZN(n681bar);
  OR2_X1 U282 ( .A1(in[171]), .A2(in[153]), .ZN(n679) );
  AND2_X1 U282bar ( .A1(inbar[171]), .A2(inbar[153]), .ZN(n679bar);
  OR2_X1 U283 ( .A1(in[187]), .A2(in[176]), .ZN(n680) );
  AND2_X1 U283bar ( .A1(inbar[187]), .A2(inbar[176]), .ZN(n680bar);
  OR2_X1 U284 ( .A1(n678), .A2(n677), .ZN(n682) );
  AND2_X1 U284bar ( .A1(n678bar), .A2(n677bar), .ZN(n682bar);
  OR2_X1 U285 ( .A1(in[245]), .A2(in[211]), .ZN(n677) );
  AND2_X1 U285bar ( .A1(inbar[245]), .A2(inbar[211]), .ZN(n677bar);
  OR2_X1 U286 ( .A1(in[97]), .A2(in[88]), .ZN(n678) );
  AND2_X1 U286bar ( .A1(inbar[97]), .A2(inbar[88]), .ZN(n678bar);
  OR2_X1 U287 ( .A1(n676), .A2(n675), .ZN(n684) );
  AND2_X1 U287bar ( .A1(n676bar), .A2(n675bar), .ZN(n684bar);
  OR2_X1 U288 ( .A1(n674), .A2(n673), .ZN(n675) );
  AND2_X1 U288bar ( .A1(n674bar), .A2(n673bar), .ZN(n675bar);
  OR2_X1 U289 ( .A1(in_10), .A2(in_0), .ZN(n673) );
  AND2_X1 U289bar ( .A1(in_10bar), .A2(in_0bar), .ZN(n673bar);
  OR2_X1 U290 ( .A1(in_59), .A2(in_5), .ZN(n674) );
  AND2_X1 U290bar ( .A1(in_59bar), .A2(in_5bar), .ZN(n674bar);
  OR2_X1 U291 ( .A1(n672), .A2(n671), .ZN(n676) );
  AND2_X1 U291bar ( .A1(n672bar), .A2(n671bar), .ZN(n676bar);
  OR2_X1 U292 ( .A1(in_60), .A2(in_6), .ZN(n671) );
  AND2_X1 U292bar ( .A1(in_60bar), .A2(in_6bar), .ZN(n671bar);
  OR2_X1 U293 ( .A1(in_77), .A2(in_69), .ZN(n672) );
  AND2_X1 U293bar ( .A1(in_77bar), .A2(in_69bar), .ZN(n672bar);
  OR2_X1 U294 ( .A1(in[113]), .A2(n864), .ZN(n700) );
  AND2_X1 U294bar ( .A1(inbar[113]), .A2(n864bar), .ZN(n700bar);
  OR2_X1 U295 ( .A1(n670), .A2(n669), .ZN(n864) );
  AND2_X1 U295bar ( .A1(n670bar), .A2(n669bar), .ZN(n864bar);
  OR2_X1 U296 ( .A1(n668), .A2(n667), .ZN(n669) );
  AND2_X1 U296bar ( .A1(n668bar), .A2(n667bar), .ZN(n669bar);
  OR2_X1 U297 ( .A1(n666), .A2(n665), .ZN(n667) );
  AND2_X1 U297bar ( .A1(n666bar), .A2(n665bar), .ZN(n667bar);
  OR2_X1 U298 ( .A1(in[125]), .A2(in[107]), .ZN(n665) );
  AND2_X1 U298bar ( .A1(inbar[125]), .A2(inbar[107]), .ZN(n665bar);
  OR2_X1 U299 ( .A1(in[138]), .A2(in[126]), .ZN(n666) );
  AND2_X1 U299bar ( .A1(inbar[138]), .A2(inbar[126]), .ZN(n666bar);
  OR2_X1 U300 ( .A1(n664), .A2(n663), .ZN(n668) );
  AND2_X1 U300bar ( .A1(n664bar), .A2(n663bar), .ZN(n668bar);
  OR2_X1 U301 ( .A1(in[189]), .A2(in[143]), .ZN(n663) );
  AND2_X1 U301bar ( .A1(inbar[189]), .A2(inbar[143]), .ZN(n663bar);
  OR2_X1 U302 ( .A1(in[99]), .A2(in[214]), .ZN(n664) );
  AND2_X1 U302bar ( .A1(inbar[99]), .A2(inbar[214]), .ZN(n664bar);
  OR2_X1 U303 ( .A1(n662), .A2(n661), .ZN(n670) );
  AND2_X1 U303bar ( .A1(n662bar), .A2(n661bar), .ZN(n670bar);
  OR2_X1 U304 ( .A1(n660), .A2(n659), .ZN(n661) );
  AND2_X1 U304bar ( .A1(n660bar), .A2(n659bar), .ZN(n661bar);
  OR2_X1 U305 ( .A1(in_15), .A2(in_12), .ZN(n659) );
  AND2_X1 U305bar ( .A1(in_15bar), .A2(in_12bar), .ZN(n659bar);
  OR2_X1 U306 ( .A1(in_20), .A2(in_2), .ZN(n660) );
  AND2_X1 U306bar ( .A1(in_20bar), .A2(in_2bar), .ZN(n660bar);
  OR2_X1 U307 ( .A1(n658), .A2(n657), .ZN(n662) );
  AND2_X1 U307bar ( .A1(n658bar), .A2(n657bar), .ZN(n662bar);
  OR2_X1 U308 ( .A1(in_30), .A2(in_3), .ZN(n657) );
  AND2_X1 U308bar ( .A1(in_30bar), .A2(in_3bar), .ZN(n657bar);
  OR2_X1 U309 ( .A1(in_4), .A2(in_38), .ZN(n658) );
  AND2_X1 U309bar ( .A1(in_4bar), .A2(in_38bar), .ZN(n658bar);
  OR2_X1 U310 ( .A1(n656), .A2(n655), .ZN(n702) );
  AND2_X1 U310bar ( .A1(n656bar), .A2(n655bar), .ZN(n702bar);
  OR2_X1 U311 ( .A1(in[148]), .A2(in[137]), .ZN(n655) );
  AND2_X1 U311bar ( .A1(inbar[148]), .A2(inbar[137]), .ZN(n655bar);
  OR2_X1 U312 ( .A1(in[149]), .A2(n654), .ZN(n656) );
  AND2_X1 U312bar ( .A1(inbar[149]), .A2(n654bar), .ZN(n656bar);
  OR2_X1 U313 ( .A1(in[195]), .A2(in[190]), .ZN(n654) );
  AND2_X1 U313bar ( .A1(inbar[195]), .A2(inbar[190]), .ZN(n654bar);
  OR2_X1 U314 ( .A1(n653), .A2(n652), .ZN(n704) );
  AND2_X1 U314bar ( .A1(n653bar), .A2(n652bar), .ZN(n704bar);
  OR2_X1 U315 ( .A1(n651), .A2(n650), .ZN(n652) );
  AND2_X1 U315bar ( .A1(n651bar), .A2(n650bar), .ZN(n652bar);
  OR2_X1 U316 ( .A1(in[98]), .A2(in[197]), .ZN(n650) );
  AND2_X1 U316bar ( .A1(inbar[98]), .A2(inbar[197]), .ZN(n650bar);
  OR2_X1 U317 ( .A1(in_11), .A2(n649), .ZN(n651) );
  AND2_X1 U317bar ( .A1(in_11bar), .A2(n649bar), .ZN(n651bar);
  OR2_X1 U318 ( .A1(in_26), .A2(in_14), .ZN(n649) );
  AND2_X1 U318bar ( .A1(in_26bar), .A2(in_14bar), .ZN(n649bar);
  OR2_X1 U319 ( .A1(n648), .A2(n647), .ZN(n653) );
  AND2_X1 U319bar ( .A1(n648bar), .A2(n647bar), .ZN(n653bar);
  OR2_X1 U320 ( .A1(in_35), .A2(in_27), .ZN(n647) );
  AND2_X1 U320bar ( .A1(in_35bar), .A2(in_27bar), .ZN(n647bar);
  OR2_X1 U321 ( .A1(in_50), .A2(n646), .ZN(n648) );
  AND2_X1 U321bar ( .A1(in_50bar), .A2(n646bar), .ZN(n648bar);
  OR2_X1 U322 ( .A1(in_78), .A2(in_61), .ZN(n646) );
  AND2_X1 U322bar ( .A1(in_78bar), .A2(in_61bar), .ZN(n646bar);
  OR2_X1 U323 ( .A1(n942), .A2(n645), .ZN(n720) );
  AND2_X1 U323bar ( .A1(n942bar), .A2(n645bar), .ZN(n720bar);
  OR2_X1 U324 ( .A1(in[106]), .A2(n863), .ZN(n645) );
  AND2_X1 U324bar ( .A1(inbar[106]), .A2(n863bar), .ZN(n645bar);
  OR2_X1 U325 ( .A1(n644), .A2(n643), .ZN(n863) );
  AND2_X1 U325bar ( .A1(n644bar), .A2(n643bar), .ZN(n863bar);
  OR2_X1 U326 ( .A1(n642), .A2(n641), .ZN(n643) );
  AND2_X1 U326bar ( .A1(n642bar), .A2(n641bar), .ZN(n643bar);
  OR2_X1 U327 ( .A1(n640), .A2(n639), .ZN(n641) );
  AND2_X1 U327bar ( .A1(n640bar), .A2(n639bar), .ZN(n641bar);
  OR2_X1 U328 ( .A1(in[127]), .A2(in[122]), .ZN(n639) );
  AND2_X1 U328bar ( .A1(inbar[127]), .A2(inbar[122]), .ZN(n639bar);
  OR2_X1 U329 ( .A1(in[156]), .A2(in[132]), .ZN(n640) );
  AND2_X1 U329bar ( .A1(inbar[156]), .A2(inbar[132]), .ZN(n640bar);
  OR2_X1 U330 ( .A1(n638), .A2(n637), .ZN(n642) );
  AND2_X1 U330bar ( .A1(n638bar), .A2(n637bar), .ZN(n642bar);
  OR2_X1 U331 ( .A1(in[159]), .A2(in[157]), .ZN(n637) );
  AND2_X1 U331bar ( .A1(inbar[159]), .A2(inbar[157]), .ZN(n637bar);
  OR2_X1 U332 ( .A1(in[185]), .A2(in[169]), .ZN(n638) );
  AND2_X1 U332bar ( .A1(inbar[185]), .A2(inbar[169]), .ZN(n638bar);
  OR2_X1 U333 ( .A1(n636), .A2(n635), .ZN(n644) );
  AND2_X1 U333bar ( .A1(n636bar), .A2(n635bar), .ZN(n644bar);
  OR2_X1 U334 ( .A1(n634), .A2(n633), .ZN(n635) );
  AND2_X1 U334bar ( .A1(n634bar), .A2(n633bar), .ZN(n635bar);
  OR2_X1 U335 ( .A1(in[239]), .A2(in[218]), .ZN(n633) );
  AND2_X1 U335bar ( .A1(inbar[239]), .A2(inbar[218]), .ZN(n633bar);
  OR2_X1 U336 ( .A1(in_13), .A2(in[87]), .ZN(n634) );
  AND2_X1 U336bar ( .A1(in_13bar), .A2(inbar[87]), .ZN(n634bar);
  OR2_X1 U337 ( .A1(n632), .A2(n631), .ZN(n636) );
  AND2_X1 U337bar ( .A1(n632bar), .A2(n631bar), .ZN(n636bar);
  OR2_X1 U338 ( .A1(in_72), .A2(in_70), .ZN(n631) );
  AND2_X1 U338bar ( .A1(in_72bar), .A2(in_70bar), .ZN(n631bar);
  OR2_X1 U339 ( .A1(in_80), .A2(in_74), .ZN(n632) );
  AND2_X1 U339bar ( .A1(in_80bar), .A2(in_74bar), .ZN(n632bar);
  OR2_X1 U340 ( .A1(n630), .A2(n629), .ZN(n942) );
  AND2_X1 U340bar ( .A1(n630bar), .A2(n629bar), .ZN(n942bar);
  OR2_X1 U341 ( .A1(n628), .A2(n627), .ZN(n629) );
  AND2_X1 U341bar ( .A1(n628bar), .A2(n627bar), .ZN(n629bar);
  OR2_X1 U342 ( .A1(n626), .A2(n625), .ZN(n627) );
  AND2_X1 U342bar ( .A1(n626bar), .A2(n625bar), .ZN(n627bar);
  OR2_X1 U343 ( .A1(in[146]), .A2(in[100]), .ZN(n625) );
  AND2_X1 U343bar ( .A1(inbar[146]), .A2(inbar[100]), .ZN(n625bar);
  OR2_X1 U344 ( .A1(in[168]), .A2(in[152]), .ZN(n626) );
  AND2_X1 U344bar ( .A1(inbar[168]), .A2(inbar[152]), .ZN(n626bar);
  OR2_X1 U345 ( .A1(n624), .A2(n623), .ZN(n628) );
  AND2_X1 U345bar ( .A1(n624bar), .A2(n623bar), .ZN(n628bar);
  OR2_X1 U346 ( .A1(in[199]), .A2(in[182]), .ZN(n623) );
  AND2_X1 U346bar ( .A1(inbar[199]), .A2(inbar[182]), .ZN(n623bar);
  OR2_X1 U347 ( .A1(in[236]), .A2(in[204]), .ZN(n624) );
  AND2_X1 U347bar ( .A1(inbar[236]), .A2(inbar[204]), .ZN(n624bar);
  OR2_X1 U348 ( .A1(n622), .A2(n621), .ZN(n630) );
  AND2_X1 U348bar ( .A1(n622bar), .A2(n621bar), .ZN(n630bar);
  OR2_X1 U349 ( .A1(n620), .A2(n619), .ZN(n621) );
  AND2_X1 U349bar ( .A1(n620bar), .A2(n619bar), .ZN(n621bar);
  OR2_X1 U350 ( .A1(in[89]), .A2(in[246]), .ZN(n619) );
  AND2_X1 U350bar ( .A1(inbar[89]), .A2(inbar[246]), .ZN(n619bar);
  OR2_X1 U351 ( .A1(in[95]), .A2(in[92]), .ZN(n620) );
  AND2_X1 U351bar ( .A1(inbar[95]), .A2(inbar[92]), .ZN(n620bar);
  OR2_X1 U352 ( .A1(n618), .A2(n617), .ZN(n622) );
  AND2_X1 U352bar ( .A1(n618bar), .A2(n617bar), .ZN(n622bar);
  OR2_X1 U353 ( .A1(in_22), .A2(in_16), .ZN(n617) );
  AND2_X1 U353bar ( .A1(in_22bar), .A2(in_16bar), .ZN(n617bar);
  OR2_X1 U354 ( .A1(in_51), .A2(in_49), .ZN(n618) );
  AND2_X1 U354bar ( .A1(in_51bar), .A2(in_49bar), .ZN(n618bar);
  OR2_X1 U355 ( .A1(n616), .A2(n615), .ZN(n722) );
  AND2_X1 U355bar ( .A1(n616bar), .A2(n615bar), .ZN(n722bar);
  OR2_X1 U356 ( .A1(in[158]), .A2(in[115]), .ZN(n615) );
  AND2_X1 U356bar ( .A1(inbar[158]), .A2(inbar[115]), .ZN(n615bar);
  OR2_X1 U357 ( .A1(in[163]), .A2(n614), .ZN(n616) );
  AND2_X1 U357bar ( .A1(inbar[163]), .A2(n614bar), .ZN(n616bar);
  OR2_X1 U358 ( .A1(in[206]), .A2(in[165]), .ZN(n614) );
  AND2_X1 U358bar ( .A1(inbar[206]), .A2(inbar[165]), .ZN(n614bar);
  OR2_X1 U359 ( .A1(n613), .A2(n612), .ZN(n724) );
  AND2_X1 U359bar ( .A1(n613bar), .A2(n612bar), .ZN(n724bar);
  OR2_X1 U360 ( .A1(n611), .A2(n610), .ZN(n612) );
  AND2_X1 U360bar ( .A1(n611bar), .A2(n610bar), .ZN(n612bar);
  OR2_X1 U361 ( .A1(in[213]), .A2(in[207]), .ZN(n610) );
  AND2_X1 U361bar ( .A1(inbar[213]), .A2(inbar[207]), .ZN(n610bar);
  OR2_X1 U362 ( .A1(in[215]), .A2(n609), .ZN(n611) );
  AND2_X1 U362bar ( .A1(inbar[215]), .A2(n609bar), .ZN(n611bar);
  OR2_X1 U363 ( .A1(in[230]), .A2(in[220]), .ZN(n609) );
  AND2_X1 U363bar ( .A1(inbar[230]), .A2(inbar[220]), .ZN(n609bar);
  OR2_X1 U364 ( .A1(n608), .A2(n607), .ZN(n613) );
  AND2_X1 U364bar ( .A1(n608bar), .A2(n607bar), .ZN(n613bar);
  OR2_X1 U365 ( .A1(in[251]), .A2(in[234]), .ZN(n607) );
  AND2_X1 U365bar ( .A1(inbar[251]), .A2(inbar[234]), .ZN(n607bar);
  OR2_X1 U366 ( .A1(in_17), .A2(n606), .ZN(n608) );
  AND2_X1 U366bar ( .A1(in_17bar), .A2(n606bar), .ZN(n608bar);
  OR2_X1 U367 ( .A1(in_65), .A2(in_56), .ZN(n606) );
  AND2_X1 U367bar ( .A1(in_65bar), .A2(in_56bar), .ZN(n606bar);
  OR2_X1 U368 ( .A1(n605), .A2(n604), .ZN(out[0]) );
  AND2_X1 U368bar ( .A1(n605bar), .A2(n604bar), .ZN(outbar[0]);
  OR2_X1 U369 ( .A1(n603), .A2(n602), .ZN(n604) );
  AND2_X1 U369bar ( .A1(n603bar), .A2(n602bar), .ZN(n604bar);
  OR2_X1 U370 ( .A1(n601), .A2(n600), .ZN(n602) );
  AND2_X1 U370bar ( .A1(n601bar), .A2(n600bar), .ZN(n602bar);
  OR2_X1 U371 ( .A1(n820), .A2(n785), .ZN(n600) );
  AND2_X1 U371bar ( .A1(n820bar), .A2(n785bar), .ZN(n600bar);
  OR2_X1 U372 ( .A1(n599), .A2(n598), .ZN(n785) );
  AND2_X1 U372bar ( .A1(n599bar), .A2(n598bar), .ZN(n785bar);
  OR2_X1 U373 ( .A1(n597), .A2(n596), .ZN(n598) );
  AND2_X1 U373bar ( .A1(n597bar), .A2(n596bar), .ZN(n598bar);
  OR2_X1 U374 ( .A1(n595), .A2(n594), .ZN(n596) );
  AND2_X1 U374bar ( .A1(n595bar), .A2(n594bar), .ZN(n596bar);
  OR2_X1 U375 ( .A1(in[135]), .A2(in[104]), .ZN(n594) );
  AND2_X1 U375bar ( .A1(inbar[135]), .A2(inbar[104]), .ZN(n594bar);
  OR2_X1 U376 ( .A1(in[188]), .A2(in[178]), .ZN(n595) );
  AND2_X1 U376bar ( .A1(inbar[188]), .A2(inbar[178]), .ZN(n595bar);
  OR2_X1 U377 ( .A1(n593), .A2(n592), .ZN(n597) );
  AND2_X1 U377bar ( .A1(n593bar), .A2(n592bar), .ZN(n597bar);
  OR2_X1 U378 ( .A1(in[217]), .A2(in[194]), .ZN(n592) );
  AND2_X1 U378bar ( .A1(inbar[217]), .A2(inbar[194]), .ZN(n592bar);
  OR2_X1 U379 ( .A1(in[237]), .A2(in[218]), .ZN(n593) );
  AND2_X1 U379bar ( .A1(inbar[237]), .A2(inbar[218]), .ZN(n593bar);
  OR2_X1 U380 ( .A1(n591), .A2(n590), .ZN(n599) );
  AND2_X1 U380bar ( .A1(n591bar), .A2(n590bar), .ZN(n599bar);
  OR2_X1 U381 ( .A1(n589), .A2(n588), .ZN(n590) );
  AND2_X1 U381bar ( .A1(n589bar), .A2(n588bar), .ZN(n590bar);
  OR2_X1 U382 ( .A1(in_2), .A2(in_10), .ZN(n588) );
  AND2_X1 U382bar ( .A1(in_2bar), .A2(in_10bar), .ZN(n588bar);
  OR2_X1 U383 ( .A1(in_47), .A2(in_22), .ZN(n589) );
  AND2_X1 U383bar ( .A1(in_47bar), .A2(in_22bar), .ZN(n589bar);
  OR2_X1 U384 ( .A1(n587), .A2(n586), .ZN(n591) );
  AND2_X1 U384bar ( .A1(n587bar), .A2(n586bar), .ZN(n591bar);
  OR2_X1 U385 ( .A1(in_56), .A2(in_54), .ZN(n586) );
  AND2_X1 U385bar ( .A1(in_56bar), .A2(in_54bar), .ZN(n586bar);
  OR2_X1 U386 ( .A1(in_63), .A2(in_61), .ZN(n587) );
  AND2_X1 U386bar ( .A1(in_63bar), .A2(in_61bar), .ZN(n587bar);
  OR2_X1 U387 ( .A1(n585), .A2(n584), .ZN(n820) );
  AND2_X1 U387bar ( .A1(n585bar), .A2(n584bar), .ZN(n820bar);
  OR2_X1 U388 ( .A1(n583), .A2(n582), .ZN(n584) );
  AND2_X1 U388bar ( .A1(n583bar), .A2(n582bar), .ZN(n584bar);
  OR2_X1 U389 ( .A1(n581), .A2(n580), .ZN(n582) );
  AND2_X1 U389bar ( .A1(n581bar), .A2(n580bar), .ZN(n582bar);
  OR2_X1 U390 ( .A1(in[158]), .A2(in[142]), .ZN(n580) );
  AND2_X1 U390bar ( .A1(inbar[158]), .A2(inbar[142]), .ZN(n580bar);
  OR2_X1 U391 ( .A1(in[175]), .A2(in[164]), .ZN(n581) );
  AND2_X1 U391bar ( .A1(inbar[175]), .A2(inbar[164]), .ZN(n581bar);
  OR2_X1 U392 ( .A1(n579), .A2(n578), .ZN(n583) );
  AND2_X1 U392bar ( .A1(n579bar), .A2(n578bar), .ZN(n583bar);
  OR2_X1 U393 ( .A1(in[228]), .A2(in[204]), .ZN(n578) );
  AND2_X1 U393bar ( .A1(inbar[228]), .A2(inbar[204]), .ZN(n578bar);
  OR2_X1 U394 ( .A1(in[91]), .A2(in[87]), .ZN(n579) );
  AND2_X1 U394bar ( .A1(inbar[91]), .A2(inbar[87]), .ZN(n579bar);
  OR2_X1 U395 ( .A1(n577), .A2(n576), .ZN(n585) );
  AND2_X1 U395bar ( .A1(n577bar), .A2(n576bar), .ZN(n585bar);
  OR2_X1 U396 ( .A1(n575), .A2(n574), .ZN(n576) );
  AND2_X1 U396bar ( .A1(n575bar), .A2(n574bar), .ZN(n576bar);
  OR2_X1 U397 ( .A1(in_21), .A2(in_11), .ZN(n574) );
  AND2_X1 U397bar ( .A1(in_21bar), .A2(in_11bar), .ZN(n574bar);
  OR2_X1 U398 ( .A1(in_5), .A2(in_3), .ZN(n575) );
  AND2_X1 U398bar ( .A1(in_5bar), .A2(in_3bar), .ZN(n575bar);
  OR2_X1 U399 ( .A1(n573), .A2(n572), .ZN(n577) );
  AND2_X1 U399bar ( .A1(n573bar), .A2(n572bar), .ZN(n577bar);
  OR2_X1 U400 ( .A1(in_68), .A2(in_64), .ZN(n572) );
  AND2_X1 U400bar ( .A1(in_68bar), .A2(in_64bar), .ZN(n572bar);
  OR2_X1 U401 ( .A1(in_76), .A2(in_73), .ZN(n573) );
  AND2_X1 U401bar ( .A1(in_76bar), .A2(in_73bar), .ZN(n573bar);
  OR2_X1 U402 ( .A1(n778), .A2(n571), .ZN(n601) );
  AND2_X1 U402bar ( .A1(n778bar), .A2(n571bar), .ZN(n601bar);
  OR2_X1 U403 ( .A1(in[100]), .A2(n965), .ZN(n571) );
  AND2_X1 U403bar ( .A1(inbar[100]), .A2(n965bar), .ZN(n571bar);
  OR2_X1 U404 ( .A1(n570), .A2(n569), .ZN(n965) );
  AND2_X1 U404bar ( .A1(n570bar), .A2(n569bar), .ZN(n965bar);
  OR2_X1 U405 ( .A1(n568), .A2(n567), .ZN(n569) );
  AND2_X1 U405bar ( .A1(n568bar), .A2(n567bar), .ZN(n569bar);
  OR2_X1 U406 ( .A1(n566), .A2(n565), .ZN(n567) );
  AND2_X1 U406bar ( .A1(n566bar), .A2(n565bar), .ZN(n567bar);
  OR2_X1 U407 ( .A1(n817), .A2(n750), .ZN(n565) );
  AND2_X1 U407bar ( .A1(n817bar), .A2(n750bar), .ZN(n565bar);
  OR2_X1 U408 ( .A1(n564), .A2(n563), .ZN(n750) );
  AND2_X1 U408bar ( .A1(n564bar), .A2(n563bar), .ZN(n750bar);
  OR2_X1 U409 ( .A1(n562), .A2(n561), .ZN(n563) );
  AND2_X1 U409bar ( .A1(n562bar), .A2(n561bar), .ZN(n563bar);
  OR2_X1 U410 ( .A1(n560), .A2(n559), .ZN(n561) );
  AND2_X1 U410bar ( .A1(n560bar), .A2(n559bar), .ZN(n561bar);
  OR2_X1 U411 ( .A1(in[119]), .A2(in[103]), .ZN(n559) );
  AND2_X1 U411bar ( .A1(inbar[119]), .A2(inbar[103]), .ZN(n559bar);
  OR2_X1 U412 ( .A1(in[137]), .A2(in[133]), .ZN(n560) );
  AND2_X1 U412bar ( .A1(inbar[137]), .A2(inbar[133]), .ZN(n560bar);
  OR2_X1 U413 ( .A1(n558), .A2(n557), .ZN(n562) );
  AND2_X1 U413bar ( .A1(n558bar), .A2(n557bar), .ZN(n562bar);
  OR2_X1 U414 ( .A1(in[176]), .A2(in[173]), .ZN(n557) );
  AND2_X1 U414bar ( .A1(inbar[176]), .A2(inbar[173]), .ZN(n557bar);
  OR2_X1 U415 ( .A1(in[210]), .A2(in[181]), .ZN(n558) );
  AND2_X1 U415bar ( .A1(inbar[210]), .A2(inbar[181]), .ZN(n558bar);
  OR2_X1 U416 ( .A1(n556), .A2(n555), .ZN(n564) );
  AND2_X1 U416bar ( .A1(n556bar), .A2(n555bar), .ZN(n564bar);
  OR2_X1 U417 ( .A1(n554), .A2(n553), .ZN(n555) );
  AND2_X1 U417bar ( .A1(n554bar), .A2(n553bar), .ZN(n555bar);
  OR2_X1 U418 ( .A1(in_13), .A2(in[234]), .ZN(n553) );
  AND2_X1 U418bar ( .A1(in_13bar), .A2(inbar[234]), .ZN(n553bar);
  OR2_X1 U419 ( .A1(in_38), .A2(in_32), .ZN(n554) );
  AND2_X1 U419bar ( .A1(in_38bar), .A2(in_32bar), .ZN(n554bar);
  OR2_X1 U420 ( .A1(n552), .A2(n551), .ZN(n556) );
  AND2_X1 U420bar ( .A1(n552bar), .A2(n551bar), .ZN(n556bar);
  OR2_X1 U421 ( .A1(in_42), .A2(in_41), .ZN(n551) );
  AND2_X1 U421bar ( .A1(in_42bar), .A2(in_41bar), .ZN(n551bar);
  OR2_X1 U422 ( .A1(in_7), .A2(in_49), .ZN(n552) );
  AND2_X1 U422bar ( .A1(in_7bar), .A2(in_49bar), .ZN(n552bar);
  OR2_X1 U423 ( .A1(n550), .A2(n549), .ZN(n817) );
  AND2_X1 U423bar ( .A1(n550bar), .A2(n549bar), .ZN(n817bar);
  OR2_X1 U424 ( .A1(n548), .A2(n547), .ZN(n549) );
  AND2_X1 U424bar ( .A1(n548bar), .A2(n547bar), .ZN(n549bar);
  OR2_X1 U425 ( .A1(n546), .A2(n545), .ZN(n547) );
  AND2_X1 U425bar ( .A1(n546bar), .A2(n545bar), .ZN(n547bar);
  OR2_X1 U426 ( .A1(in[159]), .A2(in[105]), .ZN(n545) );
  AND2_X1 U426bar ( .A1(inbar[159]), .A2(inbar[105]), .ZN(n545bar);
  OR2_X1 U427 ( .A1(in[206]), .A2(in[183]), .ZN(n546) );
  AND2_X1 U427bar ( .A1(inbar[206]), .A2(inbar[183]), .ZN(n546bar);
  OR2_X1 U428 ( .A1(n544), .A2(n543), .ZN(n548) );
  AND2_X1 U428bar ( .A1(n544bar), .A2(n543bar), .ZN(n548bar);
  OR2_X1 U429 ( .A1(in[229]), .A2(in[219]), .ZN(n543) );
  AND2_X1 U429bar ( .A1(inbar[229]), .A2(inbar[219]), .ZN(n543bar);
  OR2_X1 U430 ( .A1(in[235]), .A2(in[232]), .ZN(n544) );
  AND2_X1 U430bar ( .A1(inbar[235]), .A2(inbar[232]), .ZN(n544bar);
  OR2_X1 U431 ( .A1(n542), .A2(n541), .ZN(n550) );
  AND2_X1 U431bar ( .A1(n542bar), .A2(n541bar), .ZN(n550bar);
  OR2_X1 U432 ( .A1(n540), .A2(n539), .ZN(n541) );
  AND2_X1 U432bar ( .A1(n540bar), .A2(n539bar), .ZN(n541bar);
  OR2_X1 U433 ( .A1(in[249]), .A2(in[242]), .ZN(n539) );
  AND2_X1 U433bar ( .A1(inbar[249]), .A2(inbar[242]), .ZN(n539bar);
  OR2_X1 U434 ( .A1(in[89]), .A2(in[254]), .ZN(n540) );
  AND2_X1 U434bar ( .A1(inbar[89]), .A2(inbar[254]), .ZN(n540bar);
  OR2_X1 U435 ( .A1(n538), .A2(n537), .ZN(n542) );
  AND2_X1 U435bar ( .A1(n538bar), .A2(n537bar), .ZN(n542bar);
  OR2_X1 U436 ( .A1(in_14), .A2(in[99]), .ZN(n537) );
  AND2_X1 U436bar ( .A1(in_14bar), .A2(inbar[99]), .ZN(n537bar);
  OR2_X1 U437 ( .A1(in_60), .A2(in_18), .ZN(n538) );
  AND2_X1 U437bar ( .A1(in_60bar), .A2(in_18bar), .ZN(n538bar);
  OR2_X1 U438 ( .A1(in[113]), .A2(n763), .ZN(n566) );
  AND2_X1 U438bar ( .A1(inbar[113]), .A2(n763bar), .ZN(n566bar);
  OR2_X1 U439 ( .A1(n536), .A2(n535), .ZN(n763) );
  AND2_X1 U439bar ( .A1(n536bar), .A2(n535bar), .ZN(n763bar);
  OR2_X1 U440 ( .A1(n534), .A2(n533), .ZN(n535) );
  AND2_X1 U440bar ( .A1(n534bar), .A2(n533bar), .ZN(n535bar);
  OR2_X1 U441 ( .A1(n532), .A2(n531), .ZN(n533) );
  AND2_X1 U441bar ( .A1(n532bar), .A2(n531bar), .ZN(n533bar);
  OR2_X1 U442 ( .A1(in[115]), .A2(in[110]), .ZN(n531) );
  AND2_X1 U442bar ( .A1(inbar[115]), .A2(inbar[110]), .ZN(n531bar);
  OR2_X1 U443 ( .A1(in[125]), .A2(in[117]), .ZN(n532) );
  AND2_X1 U443bar ( .A1(inbar[125]), .A2(inbar[117]), .ZN(n532bar);
  OR2_X1 U444 ( .A1(n530), .A2(n529), .ZN(n534) );
  AND2_X1 U444bar ( .A1(n530bar), .A2(n529bar), .ZN(n534bar);
  OR2_X1 U445 ( .A1(in[180]), .A2(in[128]), .ZN(n529) );
  AND2_X1 U445bar ( .A1(inbar[180]), .A2(inbar[128]), .ZN(n529bar);
  OR2_X1 U446 ( .A1(in[205]), .A2(in[201]), .ZN(n530) );
  AND2_X1 U446bar ( .A1(inbar[205]), .A2(inbar[201]), .ZN(n530bar);
  OR2_X1 U447 ( .A1(n528), .A2(n527), .ZN(n536) );
  AND2_X1 U447bar ( .A1(n528bar), .A2(n527bar), .ZN(n536bar);
  OR2_X1 U448 ( .A1(n526), .A2(n525), .ZN(n527) );
  AND2_X1 U448bar ( .A1(n526bar), .A2(n525bar), .ZN(n527bar);
  OR2_X1 U449 ( .A1(in[244]), .A2(in[239]), .ZN(n525) );
  AND2_X1 U449bar ( .A1(inbar[244]), .A2(inbar[239]), .ZN(n525bar);
  OR2_X1 U450 ( .A1(in[95]), .A2(in[83]), .ZN(n526) );
  AND2_X1 U450bar ( .A1(inbar[95]), .A2(inbar[83]), .ZN(n526bar);
  OR2_X1 U451 ( .A1(n524), .A2(n523), .ZN(n528) );
  AND2_X1 U451bar ( .A1(n524bar), .A2(n523bar), .ZN(n528bar);
  OR2_X1 U452 ( .A1(in_24), .A2(in[97]), .ZN(n523) );
  AND2_X1 U452bar ( .A1(in_24bar), .A2(inbar[97]), .ZN(n523bar);
  OR2_X1 U453 ( .A1(in_33), .A2(in_27), .ZN(n524) );
  AND2_X1 U453bar ( .A1(in_33bar), .A2(in_27bar), .ZN(n524bar);
  OR2_X1 U454 ( .A1(n522), .A2(n521), .ZN(n568) );
  AND2_X1 U454bar ( .A1(n522bar), .A2(n521bar), .ZN(n568bar);
  OR2_X1 U455 ( .A1(in[145]), .A2(in[126]), .ZN(n521) );
  AND2_X1 U455bar ( .A1(inbar[145]), .A2(inbar[126]), .ZN(n521bar);
  OR2_X1 U456 ( .A1(in[169]), .A2(n520), .ZN(n522) );
  AND2_X1 U456bar ( .A1(inbar[169]), .A2(n520bar), .ZN(n522bar);
  OR2_X1 U457 ( .A1(in[221]), .A2(in[172]), .ZN(n520) );
  AND2_X1 U457bar ( .A1(inbar[221]), .A2(inbar[172]), .ZN(n520bar);
  OR2_X1 U458 ( .A1(n519), .A2(n518), .ZN(n570) );
  AND2_X1 U458bar ( .A1(n519bar), .A2(n518bar), .ZN(n570bar);
  OR2_X1 U459 ( .A1(n517), .A2(n516), .ZN(n518) );
  AND2_X1 U459bar ( .A1(n517bar), .A2(n516bar), .ZN(n518bar);
  OR2_X1 U460 ( .A1(in[241]), .A2(in[224]), .ZN(n516) );
  AND2_X1 U460bar ( .A1(inbar[241]), .A2(inbar[224]), .ZN(n516bar);
  OR2_X1 U461 ( .A1(in[86]), .A2(n515), .ZN(n517) );
  AND2_X1 U461bar ( .A1(inbar[86]), .A2(n515bar), .ZN(n517bar);
  OR2_X1 U462 ( .A1(in_43), .A2(in_34), .ZN(n515) );
  AND2_X1 U462bar ( .A1(in_43bar), .A2(in_34bar), .ZN(n515bar);
  OR2_X1 U463 ( .A1(n514), .A2(n513), .ZN(n519) );
  AND2_X1 U463bar ( .A1(n514bar), .A2(n513bar), .ZN(n519bar);
  OR2_X1 U464 ( .A1(in_65), .A2(in_51), .ZN(n513) );
  AND2_X1 U464bar ( .A1(in_65bar), .A2(in_51bar), .ZN(n513bar);
  OR2_X1 U465 ( .A1(in_75), .A2(n512), .ZN(n514) );
  AND2_X1 U465bar ( .A1(in_75bar), .A2(n512bar), .ZN(n514bar);
  OR2_X1 U466 ( .A1(in_81), .A2(in_77), .ZN(n512) );
  AND2_X1 U466bar ( .A1(in_81bar), .A2(in_77bar), .ZN(n512bar);
  OR2_X1 U467 ( .A1(n511), .A2(n510), .ZN(n778) );
  AND2_X1 U467bar ( .A1(n511bar), .A2(n510bar), .ZN(n778bar);
  OR2_X1 U468 ( .A1(n509), .A2(n508), .ZN(n510) );
  AND2_X1 U468bar ( .A1(n509bar), .A2(n508bar), .ZN(n510bar);
  OR2_X1 U469 ( .A1(n507), .A2(n506), .ZN(n508) );
  AND2_X1 U469bar ( .A1(n507bar), .A2(n506bar), .ZN(n508bar);
  OR2_X1 U470 ( .A1(in[107]), .A2(in[101]), .ZN(n506) );
  AND2_X1 U470bar ( .A1(inbar[107]), .A2(inbar[101]), .ZN(n506bar);
  OR2_X1 U471 ( .A1(in[139]), .A2(in[132]), .ZN(n507) );
  AND2_X1 U471bar ( .A1(inbar[139]), .A2(inbar[132]), .ZN(n507bar);
  OR2_X1 U472 ( .A1(n505), .A2(n504), .ZN(n509) );
  AND2_X1 U472bar ( .A1(n505bar), .A2(n504bar), .ZN(n509bar);
  OR2_X1 U473 ( .A1(in[146]), .A2(in[141]), .ZN(n504) );
  AND2_X1 U473bar ( .A1(inbar[146]), .A2(inbar[141]), .ZN(n504bar);
  OR2_X1 U474 ( .A1(in[203]), .A2(in[179]), .ZN(n505) );
  AND2_X1 U474bar ( .A1(inbar[203]), .A2(inbar[179]), .ZN(n505bar);
  OR2_X1 U475 ( .A1(n503), .A2(n502), .ZN(n511) );
  AND2_X1 U475bar ( .A1(n503bar), .A2(n502bar), .ZN(n511bar);
  OR2_X1 U476 ( .A1(n501), .A2(n500), .ZN(n502) );
  AND2_X1 U476bar ( .A1(n501bar), .A2(n500bar), .ZN(n502bar);
  OR2_X1 U477 ( .A1(in[243]), .A2(in[222]), .ZN(n500) );
  AND2_X1 U477bar ( .A1(inbar[243]), .A2(inbar[222]), .ZN(n500bar);
  OR2_X1 U478 ( .A1(in[251]), .A2(in[250]), .ZN(n501) );
  AND2_X1 U478bar ( .A1(inbar[251]), .A2(inbar[250]), .ZN(n501bar);
  OR2_X1 U479 ( .A1(n499), .A2(n498), .ZN(n503) );
  AND2_X1 U479bar ( .A1(n499bar), .A2(n498bar), .ZN(n503bar);
  OR2_X1 U480 ( .A1(in_37), .A2(in_19), .ZN(n498) );
  AND2_X1 U480bar ( .A1(in_37bar), .A2(in_19bar), .ZN(n498bar);
  OR2_X1 U481 ( .A1(in_78), .A2(in_6), .ZN(n499) );
  AND2_X1 U481bar ( .A1(in_78bar), .A2(in_6bar), .ZN(n499bar);
  OR2_X1 U482 ( .A1(n497), .A2(n496), .ZN(n603) );
  AND2_X1 U482bar ( .A1(n497bar), .A2(n496bar), .ZN(n603bar);
  OR2_X1 U483 ( .A1(in[112]), .A2(in[102]), .ZN(n496) );
  AND2_X1 U483bar ( .A1(inbar[112]), .A2(inbar[102]), .ZN(n496bar);
  OR2_X1 U484 ( .A1(in[123]), .A2(n495), .ZN(n497) );
  AND2_X1 U484bar ( .A1(inbar[123]), .A2(n495bar), .ZN(n497bar);
  OR2_X1 U485 ( .A1(in[143]), .A2(in[130]), .ZN(n495) );
  AND2_X1 U485bar ( .A1(inbar[143]), .A2(inbar[130]), .ZN(n495bar);
  OR2_X1 U486 ( .A1(n494), .A2(n493), .ZN(n605) );
  AND2_X1 U486bar ( .A1(n494bar), .A2(n493bar), .ZN(n605bar);
  OR2_X1 U487 ( .A1(n492), .A2(n491), .ZN(n493) );
  AND2_X1 U487bar ( .A1(n492bar), .A2(n491bar), .ZN(n493bar);
  OR2_X1 U488 ( .A1(in[216]), .A2(in[213]), .ZN(n491) );
  AND2_X1 U488bar ( .A1(inbar[216]), .A2(inbar[213]), .ZN(n491bar);
  OR2_X1 U489 ( .A1(in[227]), .A2(n490), .ZN(n492) );
  AND2_X1 U489bar ( .A1(inbar[227]), .A2(n490bar), .ZN(n492bar);
  OR2_X1 U490 ( .A1(in_0), .A2(in[248]), .ZN(n490) );
  AND2_X1 U490bar ( .A1(in_0bar), .A2(inbar[248]), .ZN(n490bar);
  OR2_X1 U491 ( .A1(n489), .A2(n488), .ZN(n494) );
  AND2_X1 U491bar ( .A1(n489bar), .A2(n488bar), .ZN(n494bar);
  OR2_X1 U492 ( .A1(in_46), .A2(in_44), .ZN(n488) );
  AND2_X1 U492bar ( .A1(in_46bar), .A2(in_44bar), .ZN(n488bar);
  OR2_X1 U493 ( .A1(in_50), .A2(n487), .ZN(n489) );
  AND2_X1 U493bar ( .A1(in_50bar), .A2(n487bar), .ZN(n489bar);
  OR2_X1 U494 ( .A1(in_9), .A2(in_80), .ZN(n487) );
  AND2_X1 U494bar ( .A1(in_9bar), .A2(in_80bar), .ZN(n487bar);
endmodule




module sBox_13 ( in, out );
  input [7:0] in;
  //input_done

  output [7:0] out;
  //output_done

  wire   [255:0] decodeOut;
  //wire_done

  decode_13 dec ( .in(in), .out(decodeOut) );
  encode_13 enc ( .in(decodeOut), .out(out) );
endmodule


module CD2_53 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_54 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_55 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_56 ( a, b, y );
 input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD4_27 ( a, b, y );
  input [3:0] a;
  input [3:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  //input_done

  output [15:0] y;
  reg [15:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]);
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]);
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]);
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]);
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]);
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]);
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]);
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]);
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]);
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]);
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]);
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]);
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]);
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]);
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]);
endmodule




module CD4_28 ( a, b, y );
  input [3:0] a;
  input [3:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  //input_done

  output [15:0] y;
  reg [15:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]);
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]);
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]);
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]);
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]);
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]);
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]);
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]);
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]);
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]);
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]);
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]);
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]);
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]);
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]);
endmodule




module CD16_14 ( a, b, y );
  input [15:0] a;
  input [15:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign abar[8] = ~a[8];
  assign abar[9] = ~a[9];
  assign abar[10] = ~a[10];
  assign abar[11] = ~a[11];
  assign abar[12] = ~a[12];
  assign abar[13] = ~a[13];
  assign abar[14] = ~a[14];
  assign abar[15] = ~a[15];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign bbar[8] = ~b[8];
  assign bbar[9] = ~b[9];
  assign bbar[10] = ~b[10];
  assign bbar[11] = ~b[11];
  assign bbar[12] = ~b[12];
  assign bbar[13] = ~b[13];
  assign bbar[14] = ~b[14];
  assign bbar[15] = ~b[15];
  //input_done

  output [255:0] y;
  reg [255:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[9]), .A2(a[0]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[9]), .A2(abar[0]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[3]), .A2(a[6]), .ZN(y[99]) );
  OR2_X1 U2bar ( .A1(bbar[3]), .A2(abar[6]), .ZN(ybar[99]);
  AND2_X1 U3 ( .A1(b[2]), .A2(a[6]), .ZN(y[98]) );
  OR2_X1 U3bar ( .A1(bbar[2]), .A2(abar[6]), .ZN(ybar[98]);
  AND2_X1 U4 ( .A1(b[1]), .A2(a[6]), .ZN(y[97]) );
  OR2_X1 U4bar ( .A1(bbar[1]), .A2(abar[6]), .ZN(ybar[97]);
  AND2_X1 U5 ( .A1(b[0]), .A2(a[6]), .ZN(y[96]) );
  OR2_X1 U5bar ( .A1(bbar[0]), .A2(abar[6]), .ZN(ybar[96]);
  AND2_X1 U6 ( .A1(b[15]), .A2(a[5]), .ZN(y[95]) );
  OR2_X1 U6bar ( .A1(bbar[15]), .A2(abar[5]), .ZN(ybar[95]);
  AND2_X1 U7 ( .A1(b[14]), .A2(a[5]), .ZN(y[94]) );
  OR2_X1 U7bar ( .A1(bbar[14]), .A2(abar[5]), .ZN(ybar[94]);
  AND2_X1 U8 ( .A1(b[13]), .A2(a[5]), .ZN(y[93]) );
  OR2_X1 U8bar ( .A1(bbar[13]), .A2(abar[5]), .ZN(ybar[93]);
  AND2_X1 U9 ( .A1(b[12]), .A2(a[5]), .ZN(y[92]) );
  OR2_X1 U9bar ( .A1(bbar[12]), .A2(abar[5]), .ZN(ybar[92]);
  AND2_X1 U10 ( .A1(b[11]), .A2(a[5]), .ZN(y[91]) );
  OR2_X1 U10bar ( .A1(bbar[11]), .A2(abar[5]), .ZN(ybar[91]);
  AND2_X1 U11 ( .A1(b[10]), .A2(a[5]), .ZN(y[90]) );
  OR2_X1 U11bar ( .A1(bbar[10]), .A2(abar[5]), .ZN(ybar[90]);
  AND2_X1 U12 ( .A1(b[8]), .A2(a[0]), .ZN(y[8]) );
  OR2_X1 U12bar ( .A1(bbar[8]), .A2(abar[0]), .ZN(ybar[8]);
  AND2_X1 U13 ( .A1(a[5]), .A2(b[9]), .ZN(y[89]) );
  OR2_X1 U13bar ( .A1(abar[5]), .A2(bbar[9]), .ZN(ybar[89]);
  AND2_X1 U14 ( .A1(b[8]), .A2(a[5]), .ZN(y[88]) );
  OR2_X1 U14bar ( .A1(bbar[8]), .A2(abar[5]), .ZN(ybar[88]);
  AND2_X1 U15 ( .A1(b[7]), .A2(a[5]), .ZN(y[87]) );
  OR2_X1 U15bar ( .A1(bbar[7]), .A2(abar[5]), .ZN(ybar[87]);
  AND2_X1 U16 ( .A1(b[6]), .A2(a[5]), .ZN(y[86]) );
  OR2_X1 U16bar ( .A1(bbar[6]), .A2(abar[5]), .ZN(ybar[86]);
  AND2_X1 U17 ( .A1(b[5]), .A2(a[5]), .ZN(y[85]) );
  OR2_X1 U17bar ( .A1(bbar[5]), .A2(abar[5]), .ZN(ybar[85]);
  AND2_X1 U18 ( .A1(b[4]), .A2(a[5]), .ZN(y[84]) );
  OR2_X1 U18bar ( .A1(bbar[4]), .A2(abar[5]), .ZN(ybar[84]);
  AND2_X1 U19 ( .A1(a[5]), .A2(b[3]), .ZN(y[83]) );
  OR2_X1 U19bar ( .A1(abar[5]), .A2(bbar[3]), .ZN(ybar[83]);
  AND2_X1 U20 ( .A1(a[5]), .A2(b[2]), .ZN(y[82]) );
  OR2_X1 U20bar ( .A1(abar[5]), .A2(bbar[2]), .ZN(ybar[82]);
  AND2_X1 U21 ( .A1(a[5]), .A2(b[1]), .ZN(y[81]) );
  OR2_X1 U21bar ( .A1(abar[5]), .A2(bbar[1]), .ZN(ybar[81]);
  AND2_X1 U22 ( .A1(a[5]), .A2(b[0]), .ZN(y[80]) );
  OR2_X1 U22bar ( .A1(abar[5]), .A2(bbar[0]), .ZN(ybar[80]);
  AND2_X1 U23 ( .A1(b[7]), .A2(a[0]), .ZN(y[7]) );
  OR2_X1 U23bar ( .A1(bbar[7]), .A2(abar[0]), .ZN(ybar[7]);
  AND2_X1 U24 ( .A1(a[4]), .A2(b[15]), .ZN(y[79]) );
  OR2_X1 U24bar ( .A1(abar[4]), .A2(bbar[15]), .ZN(ybar[79]);
  AND2_X1 U25 ( .A1(a[4]), .A2(b[14]), .ZN(y[78]) );
  OR2_X1 U25bar ( .A1(abar[4]), .A2(bbar[14]), .ZN(ybar[78]);
  AND2_X1 U26 ( .A1(a[4]), .A2(b[13]), .ZN(y[77]) );
  OR2_X1 U26bar ( .A1(abar[4]), .A2(bbar[13]), .ZN(ybar[77]);
  AND2_X1 U27 ( .A1(a[4]), .A2(b[12]), .ZN(y[76]) );
  OR2_X1 U27bar ( .A1(abar[4]), .A2(bbar[12]), .ZN(ybar[76]);
  AND2_X1 U28 ( .A1(a[4]), .A2(b[11]), .ZN(y[75]) );
  OR2_X1 U28bar ( .A1(abar[4]), .A2(bbar[11]), .ZN(ybar[75]);
  AND2_X1 U29 ( .A1(a[4]), .A2(b[10]), .ZN(y[74]) );
  OR2_X1 U29bar ( .A1(abar[4]), .A2(bbar[10]), .ZN(ybar[74]);
  AND2_X1 U30 ( .A1(a[4]), .A2(b[9]), .ZN(y[73]) );
  OR2_X1 U30bar ( .A1(abar[4]), .A2(bbar[9]), .ZN(ybar[73]);
  AND2_X1 U31 ( .A1(a[4]), .A2(b[8]), .ZN(y[72]) );
  OR2_X1 U31bar ( .A1(abar[4]), .A2(bbar[8]), .ZN(ybar[72]);
  AND2_X1 U32 ( .A1(a[4]), .A2(b[7]), .ZN(y[71]) );
  OR2_X1 U32bar ( .A1(abar[4]), .A2(bbar[7]), .ZN(ybar[71]);
  AND2_X1 U33 ( .A1(a[4]), .A2(b[6]), .ZN(y[70]) );
  OR2_X1 U33bar ( .A1(abar[4]), .A2(bbar[6]), .ZN(ybar[70]);
  AND2_X1 U34 ( .A1(b[6]), .A2(a[0]), .ZN(y[6]) );
  OR2_X1 U34bar ( .A1(bbar[6]), .A2(abar[0]), .ZN(ybar[6]);
  AND2_X1 U35 ( .A1(a[4]), .A2(b[5]), .ZN(y[69]) );
  OR2_X1 U35bar ( .A1(abar[4]), .A2(bbar[5]), .ZN(ybar[69]);
  AND2_X1 U36 ( .A1(a[4]), .A2(b[4]), .ZN(y[68]) );
  OR2_X1 U36bar ( .A1(abar[4]), .A2(bbar[4]), .ZN(ybar[68]);
  AND2_X1 U37 ( .A1(a[4]), .A2(b[3]), .ZN(y[67]) );
  OR2_X1 U37bar ( .A1(abar[4]), .A2(bbar[3]), .ZN(ybar[67]);
  AND2_X1 U38 ( .A1(a[4]), .A2(b[2]), .ZN(y[66]) );
  OR2_X1 U38bar ( .A1(abar[4]), .A2(bbar[2]), .ZN(ybar[66]);
  AND2_X1 U39 ( .A1(a[4]), .A2(b[1]), .ZN(y[65]) );
  OR2_X1 U39bar ( .A1(abar[4]), .A2(bbar[1]), .ZN(ybar[65]);
  AND2_X1 U40 ( .A1(a[4]), .A2(b[0]), .ZN(y[64]) );
  OR2_X1 U40bar ( .A1(abar[4]), .A2(bbar[0]), .ZN(ybar[64]);
  AND2_X1 U41 ( .A1(a[3]), .A2(b[15]), .ZN(y[63]) );
  OR2_X1 U41bar ( .A1(abar[3]), .A2(bbar[15]), .ZN(ybar[63]);
  AND2_X1 U42 ( .A1(a[3]), .A2(b[14]), .ZN(y[62]) );
  OR2_X1 U42bar ( .A1(abar[3]), .A2(bbar[14]), .ZN(ybar[62]);
  AND2_X1 U43 ( .A1(a[3]), .A2(b[13]), .ZN(y[61]) );
  OR2_X1 U43bar ( .A1(abar[3]), .A2(bbar[13]), .ZN(ybar[61]);
  AND2_X1 U44 ( .A1(a[3]), .A2(b[12]), .ZN(y[60]) );
  OR2_X1 U44bar ( .A1(abar[3]), .A2(bbar[12]), .ZN(ybar[60]);
  AND2_X1 U45 ( .A1(b[5]), .A2(a[0]), .ZN(y[5]) );
  OR2_X1 U45bar ( .A1(bbar[5]), .A2(abar[0]), .ZN(ybar[5]);
  AND2_X1 U46 ( .A1(a[3]), .A2(b[11]), .ZN(y[59]) );
  OR2_X1 U46bar ( .A1(abar[3]), .A2(bbar[11]), .ZN(ybar[59]);
  AND2_X1 U47 ( .A1(a[3]), .A2(b[10]), .ZN(y[58]) );
  OR2_X1 U47bar ( .A1(abar[3]), .A2(bbar[10]), .ZN(ybar[58]);
  AND2_X1 U48 ( .A1(a[3]), .A2(b[9]), .ZN(y[57]) );
  OR2_X1 U48bar ( .A1(abar[3]), .A2(bbar[9]), .ZN(ybar[57]);
  AND2_X1 U49 ( .A1(a[3]), .A2(b[8]), .ZN(y[56]) );
  OR2_X1 U49bar ( .A1(abar[3]), .A2(bbar[8]), .ZN(ybar[56]);
  AND2_X1 U50 ( .A1(a[3]), .A2(b[7]), .ZN(y[55]) );
  OR2_X1 U50bar ( .A1(abar[3]), .A2(bbar[7]), .ZN(ybar[55]);
  AND2_X1 U51 ( .A1(a[3]), .A2(b[6]), .ZN(y[54]) );
  OR2_X1 U51bar ( .A1(abar[3]), .A2(bbar[6]), .ZN(ybar[54]);
  AND2_X1 U52 ( .A1(a[3]), .A2(b[5]), .ZN(y[53]) );
  OR2_X1 U52bar ( .A1(abar[3]), .A2(bbar[5]), .ZN(ybar[53]);
  AND2_X1 U53 ( .A1(a[3]), .A2(b[4]), .ZN(y[52]) );
  OR2_X1 U53bar ( .A1(abar[3]), .A2(bbar[4]), .ZN(ybar[52]);
  AND2_X1 U54 ( .A1(a[3]), .A2(b[3]), .ZN(y[51]) );
  OR2_X1 U54bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[51]);
  AND2_X1 U55 ( .A1(a[3]), .A2(b[2]), .ZN(y[50]) );
  OR2_X1 U55bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[50]);
  AND2_X1 U56 ( .A1(b[4]), .A2(a[0]), .ZN(y[4]) );
  OR2_X1 U56bar ( .A1(bbar[4]), .A2(abar[0]), .ZN(ybar[4]);
  AND2_X1 U57 ( .A1(a[3]), .A2(b[1]), .ZN(y[49]) );
  OR2_X1 U57bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[49]);
  AND2_X1 U58 ( .A1(a[3]), .A2(b[0]), .ZN(y[48]) );
  OR2_X1 U58bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[48]);
  AND2_X1 U59 ( .A1(a[2]), .A2(b[15]), .ZN(y[47]) );
  OR2_X1 U59bar ( .A1(abar[2]), .A2(bbar[15]), .ZN(ybar[47]);
  AND2_X1 U60 ( .A1(a[2]), .A2(b[14]), .ZN(y[46]) );
  OR2_X1 U60bar ( .A1(abar[2]), .A2(bbar[14]), .ZN(ybar[46]);
  AND2_X1 U61 ( .A1(a[2]), .A2(b[13]), .ZN(y[45]) );
  OR2_X1 U61bar ( .A1(abar[2]), .A2(bbar[13]), .ZN(ybar[45]);
  AND2_X1 U62 ( .A1(a[2]), .A2(b[12]), .ZN(y[44]) );
  OR2_X1 U62bar ( .A1(abar[2]), .A2(bbar[12]), .ZN(ybar[44]);
  AND2_X1 U63 ( .A1(a[2]), .A2(b[11]), .ZN(y[43]) );
  OR2_X1 U63bar ( .A1(abar[2]), .A2(bbar[11]), .ZN(ybar[43]);
  AND2_X1 U64 ( .A1(a[2]), .A2(b[10]), .ZN(y[42]) );
  OR2_X1 U64bar ( .A1(abar[2]), .A2(bbar[10]), .ZN(ybar[42]);
  AND2_X1 U65 ( .A1(a[2]), .A2(b[9]), .ZN(y[41]) );
  OR2_X1 U65bar ( .A1(abar[2]), .A2(bbar[9]), .ZN(ybar[41]);
  AND2_X1 U66 ( .A1(a[2]), .A2(b[8]), .ZN(y[40]) );
  OR2_X1 U66bar ( .A1(abar[2]), .A2(bbar[8]), .ZN(ybar[40]);
  AND2_X1 U67 ( .A1(b[3]), .A2(a[0]), .ZN(y[3]) );
  OR2_X1 U67bar ( .A1(bbar[3]), .A2(abar[0]), .ZN(ybar[3]);
  AND2_X1 U68 ( .A1(a[2]), .A2(b[7]), .ZN(y[39]) );
  OR2_X1 U68bar ( .A1(abar[2]), .A2(bbar[7]), .ZN(ybar[39]);
  AND2_X1 U69 ( .A1(a[2]), .A2(b[6]), .ZN(y[38]) );
  OR2_X1 U69bar ( .A1(abar[2]), .A2(bbar[6]), .ZN(ybar[38]);
  AND2_X1 U70 ( .A1(a[2]), .A2(b[5]), .ZN(y[37]) );
  OR2_X1 U70bar ( .A1(abar[2]), .A2(bbar[5]), .ZN(ybar[37]);
  AND2_X1 U71 ( .A1(a[2]), .A2(b[4]), .ZN(y[36]) );
  OR2_X1 U71bar ( .A1(abar[2]), .A2(bbar[4]), .ZN(ybar[36]);
  AND2_X1 U72 ( .A1(a[2]), .A2(b[3]), .ZN(y[35]) );
  OR2_X1 U72bar ( .A1(abar[2]), .A2(bbar[3]), .ZN(ybar[35]);
  AND2_X1 U73 ( .A1(a[2]), .A2(b[2]), .ZN(y[34]) );
  OR2_X1 U73bar ( .A1(abar[2]), .A2(bbar[2]), .ZN(ybar[34]);
  AND2_X1 U74 ( .A1(a[2]), .A2(b[1]), .ZN(y[33]) );
  OR2_X1 U74bar ( .A1(abar[2]), .A2(bbar[1]), .ZN(ybar[33]);
  AND2_X1 U75 ( .A1(a[2]), .A2(b[0]), .ZN(y[32]) );
  OR2_X1 U75bar ( .A1(abar[2]), .A2(bbar[0]), .ZN(ybar[32]);
  AND2_X1 U76 ( .A1(a[1]), .A2(b[15]), .ZN(y[31]) );
  OR2_X1 U76bar ( .A1(abar[1]), .A2(bbar[15]), .ZN(ybar[31]);
  AND2_X1 U77 ( .A1(a[1]), .A2(b[14]), .ZN(y[30]) );
  OR2_X1 U77bar ( .A1(abar[1]), .A2(bbar[14]), .ZN(ybar[30]);
  AND2_X1 U78 ( .A1(b[2]), .A2(a[0]), .ZN(y[2]) );
  OR2_X1 U78bar ( .A1(bbar[2]), .A2(abar[0]), .ZN(ybar[2]);
  AND2_X1 U79 ( .A1(a[1]), .A2(b[13]), .ZN(y[29]) );
  OR2_X1 U79bar ( .A1(abar[1]), .A2(bbar[13]), .ZN(ybar[29]);
  AND2_X1 U80 ( .A1(a[1]), .A2(b[12]), .ZN(y[28]) );
  OR2_X1 U80bar ( .A1(abar[1]), .A2(bbar[12]), .ZN(ybar[28]);
  AND2_X1 U81 ( .A1(a[1]), .A2(b[11]), .ZN(y[27]) );
  OR2_X1 U81bar ( .A1(abar[1]), .A2(bbar[11]), .ZN(ybar[27]);
  AND2_X1 U82 ( .A1(a[1]), .A2(b[10]), .ZN(y[26]) );
  OR2_X1 U82bar ( .A1(abar[1]), .A2(bbar[10]), .ZN(ybar[26]);
  AND2_X1 U83 ( .A1(a[1]), .A2(b[9]), .ZN(y[25]) );
  OR2_X1 U83bar ( .A1(abar[1]), .A2(bbar[9]), .ZN(ybar[25]);
  AND2_X1 U84 ( .A1(a[15]), .A2(b[15]), .ZN(y[255]) );
  OR2_X1 U84bar ( .A1(abar[15]), .A2(bbar[15]), .ZN(ybar[255]);
  AND2_X1 U85 ( .A1(a[15]), .A2(b[14]), .ZN(y[254]) );
  OR2_X1 U85bar ( .A1(abar[15]), .A2(bbar[14]), .ZN(ybar[254]);
  AND2_X1 U86 ( .A1(a[15]), .A2(b[13]), .ZN(y[253]) );
  OR2_X1 U86bar ( .A1(abar[15]), .A2(bbar[13]), .ZN(ybar[253]);
  AND2_X1 U87 ( .A1(a[15]), .A2(b[12]), .ZN(y[252]) );
  OR2_X1 U87bar ( .A1(abar[15]), .A2(bbar[12]), .ZN(ybar[252]);
  AND2_X1 U88 ( .A1(a[15]), .A2(b[11]), .ZN(y[251]) );
  OR2_X1 U88bar ( .A1(abar[15]), .A2(bbar[11]), .ZN(ybar[251]);
  AND2_X1 U89 ( .A1(a[15]), .A2(b[10]), .ZN(y[250]) );
  OR2_X1 U89bar ( .A1(abar[15]), .A2(bbar[10]), .ZN(ybar[250]);
  AND2_X1 U90 ( .A1(a[1]), .A2(b[8]), .ZN(y[24]) );
  OR2_X1 U90bar ( .A1(abar[1]), .A2(bbar[8]), .ZN(ybar[24]);
  AND2_X1 U91 ( .A1(a[15]), .A2(b[9]), .ZN(y[249]) );
  OR2_X1 U91bar ( .A1(abar[15]), .A2(bbar[9]), .ZN(ybar[249]);
  AND2_X1 U92 ( .A1(a[15]), .A2(b[8]), .ZN(y[248]) );
  OR2_X1 U92bar ( .A1(abar[15]), .A2(bbar[8]), .ZN(ybar[248]);
  AND2_X1 U93 ( .A1(a[15]), .A2(b[7]), .ZN(y[247]) );
  OR2_X1 U93bar ( .A1(abar[15]), .A2(bbar[7]), .ZN(ybar[247]);
  AND2_X1 U94 ( .A1(a[15]), .A2(b[6]), .ZN(y[246]) );
  OR2_X1 U94bar ( .A1(abar[15]), .A2(bbar[6]), .ZN(ybar[246]);
  AND2_X1 U95 ( .A1(a[15]), .A2(b[5]), .ZN(y[245]) );
  OR2_X1 U95bar ( .A1(abar[15]), .A2(bbar[5]), .ZN(ybar[245]);
  AND2_X1 U96 ( .A1(a[15]), .A2(b[4]), .ZN(y[244]) );
  OR2_X1 U96bar ( .A1(abar[15]), .A2(bbar[4]), .ZN(ybar[244]);
  AND2_X1 U97 ( .A1(a[15]), .A2(b[3]), .ZN(y[243]) );
  OR2_X1 U97bar ( .A1(abar[15]), .A2(bbar[3]), .ZN(ybar[243]);
  AND2_X1 U98 ( .A1(a[15]), .A2(b[2]), .ZN(y[242]) );
  OR2_X1 U98bar ( .A1(abar[15]), .A2(bbar[2]), .ZN(ybar[242]);
  AND2_X1 U99 ( .A1(a[15]), .A2(b[1]), .ZN(y[241]) );
  OR2_X1 U99bar ( .A1(abar[15]), .A2(bbar[1]), .ZN(ybar[241]);
  AND2_X1 U100 ( .A1(a[15]), .A2(b[0]), .ZN(y[240]) );
  OR2_X1 U100bar ( .A1(abar[15]), .A2(bbar[0]), .ZN(ybar[240]);
  AND2_X1 U101 ( .A1(a[1]), .A2(b[7]), .ZN(y[23]) );
  OR2_X1 U101bar ( .A1(abar[1]), .A2(bbar[7]), .ZN(ybar[23]);
  AND2_X1 U102 ( .A1(a[14]), .A2(b[15]), .ZN(y[239]) );
  OR2_X1 U102bar ( .A1(abar[14]), .A2(bbar[15]), .ZN(ybar[239]);
  AND2_X1 U103 ( .A1(a[14]), .A2(b[14]), .ZN(y[238]) );
  OR2_X1 U103bar ( .A1(abar[14]), .A2(bbar[14]), .ZN(ybar[238]);
  AND2_X1 U104 ( .A1(a[14]), .A2(b[13]), .ZN(y[237]) );
  OR2_X1 U104bar ( .A1(abar[14]), .A2(bbar[13]), .ZN(ybar[237]);
  AND2_X1 U105 ( .A1(a[14]), .A2(b[12]), .ZN(y[236]) );
  OR2_X1 U105bar ( .A1(abar[14]), .A2(bbar[12]), .ZN(ybar[236]);
  AND2_X1 U106 ( .A1(a[14]), .A2(b[11]), .ZN(y[235]) );
  OR2_X1 U106bar ( .A1(abar[14]), .A2(bbar[11]), .ZN(ybar[235]);
  AND2_X1 U107 ( .A1(a[14]), .A2(b[10]), .ZN(y[234]) );
  OR2_X1 U107bar ( .A1(abar[14]), .A2(bbar[10]), .ZN(ybar[234]);
  AND2_X1 U108 ( .A1(a[14]), .A2(b[9]), .ZN(y[233]) );
  OR2_X1 U108bar ( .A1(abar[14]), .A2(bbar[9]), .ZN(ybar[233]);
  AND2_X1 U109 ( .A1(a[14]), .A2(b[8]), .ZN(y[232]) );
  OR2_X1 U109bar ( .A1(abar[14]), .A2(bbar[8]), .ZN(ybar[232]);
  AND2_X1 U110 ( .A1(a[14]), .A2(b[7]), .ZN(y[231]) );
  OR2_X1 U110bar ( .A1(abar[14]), .A2(bbar[7]), .ZN(ybar[231]);
  AND2_X1 U111 ( .A1(a[14]), .A2(b[6]), .ZN(y[230]) );
  OR2_X1 U111bar ( .A1(abar[14]), .A2(bbar[6]), .ZN(ybar[230]);
  AND2_X1 U112 ( .A1(a[1]), .A2(b[6]), .ZN(y[22]) );
  OR2_X1 U112bar ( .A1(abar[1]), .A2(bbar[6]), .ZN(ybar[22]);
  AND2_X1 U113 ( .A1(a[14]), .A2(b[5]), .ZN(y[229]) );
  OR2_X1 U113bar ( .A1(abar[14]), .A2(bbar[5]), .ZN(ybar[229]);
  AND2_X1 U114 ( .A1(a[14]), .A2(b[4]), .ZN(y[228]) );
  OR2_X1 U114bar ( .A1(abar[14]), .A2(bbar[4]), .ZN(ybar[228]);
  AND2_X1 U115 ( .A1(a[14]), .A2(b[3]), .ZN(y[227]) );
  OR2_X1 U115bar ( .A1(abar[14]), .A2(bbar[3]), .ZN(ybar[227]);
  AND2_X1 U116 ( .A1(a[14]), .A2(b[2]), .ZN(y[226]) );
  OR2_X1 U116bar ( .A1(abar[14]), .A2(bbar[2]), .ZN(ybar[226]);
  AND2_X1 U117 ( .A1(a[14]), .A2(b[1]), .ZN(y[225]) );
  OR2_X1 U117bar ( .A1(abar[14]), .A2(bbar[1]), .ZN(ybar[225]);
  AND2_X1 U118 ( .A1(a[14]), .A2(b[0]), .ZN(y[224]) );
  OR2_X1 U118bar ( .A1(abar[14]), .A2(bbar[0]), .ZN(ybar[224]);
  AND2_X1 U119 ( .A1(a[13]), .A2(b[15]), .ZN(y[223]) );
  OR2_X1 U119bar ( .A1(abar[13]), .A2(bbar[15]), .ZN(ybar[223]);
  AND2_X1 U120 ( .A1(a[13]), .A2(b[14]), .ZN(y[222]) );
  OR2_X1 U120bar ( .A1(abar[13]), .A2(bbar[14]), .ZN(ybar[222]);
  AND2_X1 U121 ( .A1(a[13]), .A2(b[13]), .ZN(y[221]) );
  OR2_X1 U121bar ( .A1(abar[13]), .A2(bbar[13]), .ZN(ybar[221]);
  AND2_X1 U122 ( .A1(a[13]), .A2(b[12]), .ZN(y[220]) );
  OR2_X1 U122bar ( .A1(abar[13]), .A2(bbar[12]), .ZN(ybar[220]);
  AND2_X1 U123 ( .A1(a[1]), .A2(b[5]), .ZN(y[21]) );
  OR2_X1 U123bar ( .A1(abar[1]), .A2(bbar[5]), .ZN(ybar[21]);
  AND2_X1 U124 ( .A1(a[13]), .A2(b[11]), .ZN(y[219]) );
  OR2_X1 U124bar ( .A1(abar[13]), .A2(bbar[11]), .ZN(ybar[219]);
  AND2_X1 U125 ( .A1(a[13]), .A2(b[10]), .ZN(y[218]) );
  OR2_X1 U125bar ( .A1(abar[13]), .A2(bbar[10]), .ZN(ybar[218]);
  AND2_X1 U126 ( .A1(a[13]), .A2(b[9]), .ZN(y[217]) );
  OR2_X1 U126bar ( .A1(abar[13]), .A2(bbar[9]), .ZN(ybar[217]);
  AND2_X1 U127 ( .A1(a[13]), .A2(b[8]), .ZN(y[216]) );
  OR2_X1 U127bar ( .A1(abar[13]), .A2(bbar[8]), .ZN(ybar[216]);
  AND2_X1 U128 ( .A1(a[13]), .A2(b[7]), .ZN(y[215]) );
  OR2_X1 U128bar ( .A1(abar[13]), .A2(bbar[7]), .ZN(ybar[215]);
  AND2_X1 U129 ( .A1(a[13]), .A2(b[6]), .ZN(y[214]) );
  OR2_X1 U129bar ( .A1(abar[13]), .A2(bbar[6]), .ZN(ybar[214]);
  AND2_X1 U130 ( .A1(a[13]), .A2(b[5]), .ZN(y[213]) );
  OR2_X1 U130bar ( .A1(abar[13]), .A2(bbar[5]), .ZN(ybar[213]);
  AND2_X1 U131 ( .A1(a[13]), .A2(b[4]), .ZN(y[212]) );
  OR2_X1 U131bar ( .A1(abar[13]), .A2(bbar[4]), .ZN(ybar[212]);
  AND2_X1 U132 ( .A1(a[13]), .A2(b[3]), .ZN(y[211]) );
  OR2_X1 U132bar ( .A1(abar[13]), .A2(bbar[3]), .ZN(ybar[211]);
  AND2_X1 U133 ( .A1(a[13]), .A2(b[2]), .ZN(y[210]) );
  OR2_X1 U133bar ( .A1(abar[13]), .A2(bbar[2]), .ZN(ybar[210]);
  AND2_X1 U134 ( .A1(a[1]), .A2(b[4]), .ZN(y[20]) );
  OR2_X1 U134bar ( .A1(abar[1]), .A2(bbar[4]), .ZN(ybar[20]);
  AND2_X1 U135 ( .A1(a[13]), .A2(b[1]), .ZN(y[209]) );
  OR2_X1 U135bar ( .A1(abar[13]), .A2(bbar[1]), .ZN(ybar[209]);
  AND2_X1 U136 ( .A1(a[13]), .A2(b[0]), .ZN(y[208]) );
  OR2_X1 U136bar ( .A1(abar[13]), .A2(bbar[0]), .ZN(ybar[208]);
  AND2_X1 U137 ( .A1(a[12]), .A2(b[15]), .ZN(y[207]) );
  OR2_X1 U137bar ( .A1(abar[12]), .A2(bbar[15]), .ZN(ybar[207]);
  AND2_X1 U138 ( .A1(a[12]), .A2(b[14]), .ZN(y[206]) );
  OR2_X1 U138bar ( .A1(abar[12]), .A2(bbar[14]), .ZN(ybar[206]);
  AND2_X1 U139 ( .A1(a[12]), .A2(b[13]), .ZN(y[205]) );
  OR2_X1 U139bar ( .A1(abar[12]), .A2(bbar[13]), .ZN(ybar[205]);
  AND2_X1 U140 ( .A1(a[12]), .A2(b[12]), .ZN(y[204]) );
  OR2_X1 U140bar ( .A1(abar[12]), .A2(bbar[12]), .ZN(ybar[204]);
  AND2_X1 U141 ( .A1(a[12]), .A2(b[11]), .ZN(y[203]) );
  OR2_X1 U141bar ( .A1(abar[12]), .A2(bbar[11]), .ZN(ybar[203]);
  AND2_X1 U142 ( .A1(a[12]), .A2(b[10]), .ZN(y[202]) );
  OR2_X1 U142bar ( .A1(abar[12]), .A2(bbar[10]), .ZN(ybar[202]);
  AND2_X1 U143 ( .A1(a[12]), .A2(b[9]), .ZN(y[201]) );
  OR2_X1 U143bar ( .A1(abar[12]), .A2(bbar[9]), .ZN(ybar[201]);
  AND2_X1 U144 ( .A1(a[12]), .A2(b[8]), .ZN(y[200]) );
  OR2_X1 U144bar ( .A1(abar[12]), .A2(bbar[8]), .ZN(ybar[200]);
  AND2_X1 U145 ( .A1(b[1]), .A2(a[0]), .ZN(y[1]) );
  OR2_X1 U145bar ( .A1(bbar[1]), .A2(abar[0]), .ZN(ybar[1]);
  AND2_X1 U146 ( .A1(a[1]), .A2(b[3]), .ZN(y[19]) );
  OR2_X1 U146bar ( .A1(abar[1]), .A2(bbar[3]), .ZN(ybar[19]);
  AND2_X1 U147 ( .A1(a[12]), .A2(b[7]), .ZN(y[199]) );
  OR2_X1 U147bar ( .A1(abar[12]), .A2(bbar[7]), .ZN(ybar[199]);
  AND2_X1 U148 ( .A1(a[12]), .A2(b[6]), .ZN(y[198]) );
  OR2_X1 U148bar ( .A1(abar[12]), .A2(bbar[6]), .ZN(ybar[198]);
  AND2_X1 U149 ( .A1(a[12]), .A2(b[5]), .ZN(y[197]) );
  OR2_X1 U149bar ( .A1(abar[12]), .A2(bbar[5]), .ZN(ybar[197]);
  AND2_X1 U150 ( .A1(a[12]), .A2(b[4]), .ZN(y[196]) );
  OR2_X1 U150bar ( .A1(abar[12]), .A2(bbar[4]), .ZN(ybar[196]);
  AND2_X1 U151 ( .A1(a[12]), .A2(b[3]), .ZN(y[195]) );
  OR2_X1 U151bar ( .A1(abar[12]), .A2(bbar[3]), .ZN(ybar[195]);
  AND2_X1 U152 ( .A1(a[12]), .A2(b[2]), .ZN(y[194]) );
  OR2_X1 U152bar ( .A1(abar[12]), .A2(bbar[2]), .ZN(ybar[194]);
  AND2_X1 U153 ( .A1(a[12]), .A2(b[1]), .ZN(y[193]) );
  OR2_X1 U153bar ( .A1(abar[12]), .A2(bbar[1]), .ZN(ybar[193]);
  AND2_X1 U154 ( .A1(a[12]), .A2(b[0]), .ZN(y[192]) );
  OR2_X1 U154bar ( .A1(abar[12]), .A2(bbar[0]), .ZN(ybar[192]);
  AND2_X1 U155 ( .A1(a[11]), .A2(b[15]), .ZN(y[191]) );
  OR2_X1 U155bar ( .A1(abar[11]), .A2(bbar[15]), .ZN(ybar[191]);
  AND2_X1 U156 ( .A1(a[11]), .A2(b[14]), .ZN(y[190]) );
  OR2_X1 U156bar ( .A1(abar[11]), .A2(bbar[14]), .ZN(ybar[190]);
  AND2_X1 U157 ( .A1(a[1]), .A2(b[2]), .ZN(y[18]) );
  OR2_X1 U157bar ( .A1(abar[1]), .A2(bbar[2]), .ZN(ybar[18]);
  AND2_X1 U158 ( .A1(a[11]), .A2(b[13]), .ZN(y[189]) );
  OR2_X1 U158bar ( .A1(abar[11]), .A2(bbar[13]), .ZN(ybar[189]);
  AND2_X1 U159 ( .A1(a[11]), .A2(b[12]), .ZN(y[188]) );
  OR2_X1 U159bar ( .A1(abar[11]), .A2(bbar[12]), .ZN(ybar[188]);
  AND2_X1 U160 ( .A1(a[11]), .A2(b[11]), .ZN(y[187]) );
  OR2_X1 U160bar ( .A1(abar[11]), .A2(bbar[11]), .ZN(ybar[187]);
  AND2_X1 U161 ( .A1(a[11]), .A2(b[10]), .ZN(y[186]) );
  OR2_X1 U161bar ( .A1(abar[11]), .A2(bbar[10]), .ZN(ybar[186]);
  AND2_X1 U162 ( .A1(a[11]), .A2(b[9]), .ZN(y[185]) );
  OR2_X1 U162bar ( .A1(abar[11]), .A2(bbar[9]), .ZN(ybar[185]);
  AND2_X1 U163 ( .A1(a[11]), .A2(b[8]), .ZN(y[184]) );
  OR2_X1 U163bar ( .A1(abar[11]), .A2(bbar[8]), .ZN(ybar[184]);
  AND2_X1 U164 ( .A1(a[11]), .A2(b[7]), .ZN(y[183]) );
  OR2_X1 U164bar ( .A1(abar[11]), .A2(bbar[7]), .ZN(ybar[183]);
  AND2_X1 U165 ( .A1(a[11]), .A2(b[6]), .ZN(y[182]) );
  OR2_X1 U165bar ( .A1(abar[11]), .A2(bbar[6]), .ZN(ybar[182]);
  AND2_X1 U166 ( .A1(a[11]), .A2(b[5]), .ZN(y[181]) );
  OR2_X1 U166bar ( .A1(abar[11]), .A2(bbar[5]), .ZN(ybar[181]);
  AND2_X1 U167 ( .A1(a[11]), .A2(b[4]), .ZN(y[180]) );
  OR2_X1 U167bar ( .A1(abar[11]), .A2(bbar[4]), .ZN(ybar[180]);
  AND2_X1 U168 ( .A1(a[1]), .A2(b[1]), .ZN(y[17]) );
  OR2_X1 U168bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[17]);
  AND2_X1 U169 ( .A1(a[11]), .A2(b[3]), .ZN(y[179]) );
  OR2_X1 U169bar ( .A1(abar[11]), .A2(bbar[3]), .ZN(ybar[179]);
  AND2_X1 U170 ( .A1(a[11]), .A2(b[2]), .ZN(y[178]) );
  OR2_X1 U170bar ( .A1(abar[11]), .A2(bbar[2]), .ZN(ybar[178]);
  AND2_X1 U171 ( .A1(a[11]), .A2(b[1]), .ZN(y[177]) );
  OR2_X1 U171bar ( .A1(abar[11]), .A2(bbar[1]), .ZN(ybar[177]);
  AND2_X1 U172 ( .A1(a[11]), .A2(b[0]), .ZN(y[176]) );
  OR2_X1 U172bar ( .A1(abar[11]), .A2(bbar[0]), .ZN(ybar[176]);
  AND2_X1 U173 ( .A1(a[10]), .A2(b[15]), .ZN(y[175]) );
  OR2_X1 U173bar ( .A1(abar[10]), .A2(bbar[15]), .ZN(ybar[175]);
  AND2_X1 U174 ( .A1(a[10]), .A2(b[14]), .ZN(y[174]) );
  OR2_X1 U174bar ( .A1(abar[10]), .A2(bbar[14]), .ZN(ybar[174]);
  AND2_X1 U175 ( .A1(a[10]), .A2(b[13]), .ZN(y[173]) );
  OR2_X1 U175bar ( .A1(abar[10]), .A2(bbar[13]), .ZN(ybar[173]);
  AND2_X1 U176 ( .A1(a[10]), .A2(b[12]), .ZN(y[172]) );
  OR2_X1 U176bar ( .A1(abar[10]), .A2(bbar[12]), .ZN(ybar[172]);
  AND2_X1 U177 ( .A1(a[10]), .A2(b[11]), .ZN(y[171]) );
  OR2_X1 U177bar ( .A1(abar[10]), .A2(bbar[11]), .ZN(ybar[171]);
  AND2_X1 U178 ( .A1(a[10]), .A2(b[10]), .ZN(y[170]) );
  OR2_X1 U178bar ( .A1(abar[10]), .A2(bbar[10]), .ZN(ybar[170]);
  AND2_X1 U179 ( .A1(a[1]), .A2(b[0]), .ZN(y[16]) );
  OR2_X1 U179bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[16]);
  AND2_X1 U180 ( .A1(a[10]), .A2(b[9]), .ZN(y[169]) );
  OR2_X1 U180bar ( .A1(abar[10]), .A2(bbar[9]), .ZN(ybar[169]);
  AND2_X1 U181 ( .A1(a[10]), .A2(b[8]), .ZN(y[168]) );
  OR2_X1 U181bar ( .A1(abar[10]), .A2(bbar[8]), .ZN(ybar[168]);
  AND2_X1 U182 ( .A1(a[10]), .A2(b[7]), .ZN(y[167]) );
  OR2_X1 U182bar ( .A1(abar[10]), .A2(bbar[7]), .ZN(ybar[167]);
  AND2_X1 U183 ( .A1(a[10]), .A2(b[6]), .ZN(y[166]) );
  OR2_X1 U183bar ( .A1(abar[10]), .A2(bbar[6]), .ZN(ybar[166]);
  AND2_X1 U184 ( .A1(a[10]), .A2(b[5]), .ZN(y[165]) );
  OR2_X1 U184bar ( .A1(abar[10]), .A2(bbar[5]), .ZN(ybar[165]);
  AND2_X1 U185 ( .A1(a[10]), .A2(b[4]), .ZN(y[164]) );
  OR2_X1 U185bar ( .A1(abar[10]), .A2(bbar[4]), .ZN(ybar[164]);
  AND2_X1 U186 ( .A1(a[10]), .A2(b[3]), .ZN(y[163]) );
  OR2_X1 U186bar ( .A1(abar[10]), .A2(bbar[3]), .ZN(ybar[163]);
  AND2_X1 U187 ( .A1(a[10]), .A2(b[2]), .ZN(y[162]) );
  OR2_X1 U187bar ( .A1(abar[10]), .A2(bbar[2]), .ZN(ybar[162]);
  AND2_X1 U188 ( .A1(a[10]), .A2(b[1]), .ZN(y[161]) );
  OR2_X1 U188bar ( .A1(abar[10]), .A2(bbar[1]), .ZN(ybar[161]);
  AND2_X1 U189 ( .A1(a[10]), .A2(b[0]), .ZN(y[160]) );
  OR2_X1 U189bar ( .A1(abar[10]), .A2(bbar[0]), .ZN(ybar[160]);
  AND2_X1 U190 ( .A1(b[15]), .A2(a[0]), .ZN(y[15]) );
  OR2_X1 U190bar ( .A1(bbar[15]), .A2(abar[0]), .ZN(ybar[15]);
  AND2_X1 U191 ( .A1(a[9]), .A2(b[15]), .ZN(y[159]) );
  OR2_X1 U191bar ( .A1(abar[9]), .A2(bbar[15]), .ZN(ybar[159]);
  AND2_X1 U192 ( .A1(a[9]), .A2(b[14]), .ZN(y[158]) );
  OR2_X1 U192bar ( .A1(abar[9]), .A2(bbar[14]), .ZN(ybar[158]);
  AND2_X1 U193 ( .A1(a[9]), .A2(b[13]), .ZN(y[157]) );
  OR2_X1 U193bar ( .A1(abar[9]), .A2(bbar[13]), .ZN(ybar[157]);
  AND2_X1 U194 ( .A1(a[9]), .A2(b[12]), .ZN(y[156]) );
  OR2_X1 U194bar ( .A1(abar[9]), .A2(bbar[12]), .ZN(ybar[156]);
  AND2_X1 U195 ( .A1(a[9]), .A2(b[11]), .ZN(y[155]) );
  OR2_X1 U195bar ( .A1(abar[9]), .A2(bbar[11]), .ZN(ybar[155]);
  AND2_X1 U196 ( .A1(a[9]), .A2(b[10]), .ZN(y[154]) );
  OR2_X1 U196bar ( .A1(abar[9]), .A2(bbar[10]), .ZN(ybar[154]);
  AND2_X1 U197 ( .A1(a[9]), .A2(b[9]), .ZN(y[153]) );
  OR2_X1 U197bar ( .A1(abar[9]), .A2(bbar[9]), .ZN(ybar[153]);
  AND2_X1 U198 ( .A1(a[9]), .A2(b[8]), .ZN(y[152]) );
  OR2_X1 U198bar ( .A1(abar[9]), .A2(bbar[8]), .ZN(ybar[152]);
  AND2_X1 U199 ( .A1(a[9]), .A2(b[7]), .ZN(y[151]) );
  OR2_X1 U199bar ( .A1(abar[9]), .A2(bbar[7]), .ZN(ybar[151]);
  AND2_X1 U200 ( .A1(a[9]), .A2(b[6]), .ZN(y[150]) );
  OR2_X1 U200bar ( .A1(abar[9]), .A2(bbar[6]), .ZN(ybar[150]);
  AND2_X1 U201 ( .A1(b[14]), .A2(a[0]), .ZN(y[14]) );
  OR2_X1 U201bar ( .A1(bbar[14]), .A2(abar[0]), .ZN(ybar[14]);
  AND2_X1 U202 ( .A1(a[9]), .A2(b[5]), .ZN(y[149]) );
  OR2_X1 U202bar ( .A1(abar[9]), .A2(bbar[5]), .ZN(ybar[149]);
  AND2_X1 U203 ( .A1(a[9]), .A2(b[4]), .ZN(y[148]) );
  OR2_X1 U203bar ( .A1(abar[9]), .A2(bbar[4]), .ZN(ybar[148]);
  AND2_X1 U204 ( .A1(a[9]), .A2(b[3]), .ZN(y[147]) );
  OR2_X1 U204bar ( .A1(abar[9]), .A2(bbar[3]), .ZN(ybar[147]);
  AND2_X1 U205 ( .A1(a[9]), .A2(b[2]), .ZN(y[146]) );
  OR2_X1 U205bar ( .A1(abar[9]), .A2(bbar[2]), .ZN(ybar[146]);
  AND2_X1 U206 ( .A1(a[9]), .A2(b[1]), .ZN(y[145]) );
  OR2_X1 U206bar ( .A1(abar[9]), .A2(bbar[1]), .ZN(ybar[145]);
  AND2_X1 U207 ( .A1(a[9]), .A2(b[0]), .ZN(y[144]) );
  OR2_X1 U207bar ( .A1(abar[9]), .A2(bbar[0]), .ZN(ybar[144]);
  AND2_X1 U208 ( .A1(a[8]), .A2(b[15]), .ZN(y[143]) );
  OR2_X1 U208bar ( .A1(abar[8]), .A2(bbar[15]), .ZN(ybar[143]);
  AND2_X1 U209 ( .A1(a[8]), .A2(b[14]), .ZN(y[142]) );
  OR2_X1 U209bar ( .A1(abar[8]), .A2(bbar[14]), .ZN(ybar[142]);
  AND2_X1 U210 ( .A1(a[8]), .A2(b[13]), .ZN(y[141]) );
  OR2_X1 U210bar ( .A1(abar[8]), .A2(bbar[13]), .ZN(ybar[141]);
  AND2_X1 U211 ( .A1(a[8]), .A2(b[12]), .ZN(y[140]) );
  OR2_X1 U211bar ( .A1(abar[8]), .A2(bbar[12]), .ZN(ybar[140]);
  AND2_X1 U212 ( .A1(b[13]), .A2(a[0]), .ZN(y[13]) );
  OR2_X1 U212bar ( .A1(bbar[13]), .A2(abar[0]), .ZN(ybar[13]);
  AND2_X1 U213 ( .A1(a[8]), .A2(b[11]), .ZN(y[139]) );
  OR2_X1 U213bar ( .A1(abar[8]), .A2(bbar[11]), .ZN(ybar[139]);
  AND2_X1 U214 ( .A1(a[8]), .A2(b[10]), .ZN(y[138]) );
  OR2_X1 U214bar ( .A1(abar[8]), .A2(bbar[10]), .ZN(ybar[138]);
  AND2_X1 U215 ( .A1(a[8]), .A2(b[9]), .ZN(y[137]) );
  OR2_X1 U215bar ( .A1(abar[8]), .A2(bbar[9]), .ZN(ybar[137]);
  AND2_X1 U216 ( .A1(a[8]), .A2(b[8]), .ZN(y[136]) );
  OR2_X1 U216bar ( .A1(abar[8]), .A2(bbar[8]), .ZN(ybar[136]);
  AND2_X1 U217 ( .A1(a[8]), .A2(b[7]), .ZN(y[135]) );
  OR2_X1 U217bar ( .A1(abar[8]), .A2(bbar[7]), .ZN(ybar[135]);
  AND2_X1 U218 ( .A1(a[8]), .A2(b[6]), .ZN(y[134]) );
  OR2_X1 U218bar ( .A1(abar[8]), .A2(bbar[6]), .ZN(ybar[134]);
  AND2_X1 U219 ( .A1(a[8]), .A2(b[5]), .ZN(y[133]) );
  OR2_X1 U219bar ( .A1(abar[8]), .A2(bbar[5]), .ZN(ybar[133]);
  AND2_X1 U220 ( .A1(a[8]), .A2(b[4]), .ZN(y[132]) );
  OR2_X1 U220bar ( .A1(abar[8]), .A2(bbar[4]), .ZN(ybar[132]);
  AND2_X1 U221 ( .A1(a[8]), .A2(b[3]), .ZN(y[131]) );
  OR2_X1 U221bar ( .A1(abar[8]), .A2(bbar[3]), .ZN(ybar[131]);
  AND2_X1 U222 ( .A1(a[8]), .A2(b[2]), .ZN(y[130]) );
  OR2_X1 U222bar ( .A1(abar[8]), .A2(bbar[2]), .ZN(ybar[130]);
  AND2_X1 U223 ( .A1(b[12]), .A2(a[0]), .ZN(y[12]) );
  OR2_X1 U223bar ( .A1(bbar[12]), .A2(abar[0]), .ZN(ybar[12]);
  AND2_X1 U224 ( .A1(a[8]), .A2(b[1]), .ZN(y[129]) );
  OR2_X1 U224bar ( .A1(abar[8]), .A2(bbar[1]), .ZN(ybar[129]);
  AND2_X1 U225 ( .A1(a[8]), .A2(b[0]), .ZN(y[128]) );
  OR2_X1 U225bar ( .A1(abar[8]), .A2(bbar[0]), .ZN(ybar[128]);
  AND2_X1 U226 ( .A1(a[7]), .A2(b[15]), .ZN(y[127]) );
  OR2_X1 U226bar ( .A1(abar[7]), .A2(bbar[15]), .ZN(ybar[127]);
  AND2_X1 U227 ( .A1(a[7]), .A2(b[14]), .ZN(y[126]) );
  OR2_X1 U227bar ( .A1(abar[7]), .A2(bbar[14]), .ZN(ybar[126]);
  AND2_X1 U228 ( .A1(a[7]), .A2(b[13]), .ZN(y[125]) );
  OR2_X1 U228bar ( .A1(abar[7]), .A2(bbar[13]), .ZN(ybar[125]);
  AND2_X1 U229 ( .A1(a[7]), .A2(b[12]), .ZN(y[124]) );
  OR2_X1 U229bar ( .A1(abar[7]), .A2(bbar[12]), .ZN(ybar[124]);
  AND2_X1 U230 ( .A1(a[7]), .A2(b[11]), .ZN(y[123]) );
  OR2_X1 U230bar ( .A1(abar[7]), .A2(bbar[11]), .ZN(ybar[123]);
  AND2_X1 U231 ( .A1(a[7]), .A2(b[10]), .ZN(y[122]) );
  OR2_X1 U231bar ( .A1(abar[7]), .A2(bbar[10]), .ZN(ybar[122]);
  AND2_X1 U232 ( .A1(a[7]), .A2(b[9]), .ZN(y[121]) );
  OR2_X1 U232bar ( .A1(abar[7]), .A2(bbar[9]), .ZN(ybar[121]);
  AND2_X1 U233 ( .A1(a[7]), .A2(b[8]), .ZN(y[120]) );
  OR2_X1 U233bar ( .A1(abar[7]), .A2(bbar[8]), .ZN(ybar[120]);
  AND2_X1 U234 ( .A1(b[11]), .A2(a[0]), .ZN(y[11]) );
  OR2_X1 U234bar ( .A1(bbar[11]), .A2(abar[0]), .ZN(ybar[11]);
  AND2_X1 U235 ( .A1(a[7]), .A2(b[7]), .ZN(y[119]) );
  OR2_X1 U235bar ( .A1(abar[7]), .A2(bbar[7]), .ZN(ybar[119]);
  AND2_X1 U236 ( .A1(a[7]), .A2(b[6]), .ZN(y[118]) );
  OR2_X1 U236bar ( .A1(abar[7]), .A2(bbar[6]), .ZN(ybar[118]);
  AND2_X1 U237 ( .A1(a[7]), .A2(b[5]), .ZN(y[117]) );
  OR2_X1 U237bar ( .A1(abar[7]), .A2(bbar[5]), .ZN(ybar[117]);
  AND2_X1 U238 ( .A1(a[7]), .A2(b[4]), .ZN(y[116]) );
  OR2_X1 U238bar ( .A1(abar[7]), .A2(bbar[4]), .ZN(ybar[116]);
  AND2_X1 U239 ( .A1(a[7]), .A2(b[3]), .ZN(y[115]) );
  OR2_X1 U239bar ( .A1(abar[7]), .A2(bbar[3]), .ZN(ybar[115]);
  AND2_X1 U240 ( .A1(a[7]), .A2(b[2]), .ZN(y[114]) );
  OR2_X1 U240bar ( .A1(abar[7]), .A2(bbar[2]), .ZN(ybar[114]);
  AND2_X1 U241 ( .A1(a[7]), .A2(b[1]), .ZN(y[113]) );
  OR2_X1 U241bar ( .A1(abar[7]), .A2(bbar[1]), .ZN(ybar[113]);
  AND2_X1 U242 ( .A1(a[7]), .A2(b[0]), .ZN(y[112]) );
  OR2_X1 U242bar ( .A1(abar[7]), .A2(bbar[0]), .ZN(ybar[112]);
  AND2_X1 U243 ( .A1(b[15]), .A2(a[6]), .ZN(y[111]) );
  OR2_X1 U243bar ( .A1(bbar[15]), .A2(abar[6]), .ZN(ybar[111]);
  AND2_X1 U244 ( .A1(b[14]), .A2(a[6]), .ZN(y[110]) );
  OR2_X1 U244bar ( .A1(bbar[14]), .A2(abar[6]), .ZN(ybar[110]);
  AND2_X1 U245 ( .A1(b[10]), .A2(a[0]), .ZN(y[10]) );
  OR2_X1 U245bar ( .A1(bbar[10]), .A2(abar[0]), .ZN(ybar[10]);
  AND2_X1 U246 ( .A1(b[13]), .A2(a[6]), .ZN(y[109]) );
  OR2_X1 U246bar ( .A1(bbar[13]), .A2(abar[6]), .ZN(ybar[109]);
  AND2_X1 U247 ( .A1(b[12]), .A2(a[6]), .ZN(y[108]) );
  OR2_X1 U247bar ( .A1(bbar[12]), .A2(abar[6]), .ZN(ybar[108]);
  AND2_X1 U248 ( .A1(b[11]), .A2(a[6]), .ZN(y[107]) );
  OR2_X1 U248bar ( .A1(bbar[11]), .A2(abar[6]), .ZN(ybar[107]);
  AND2_X1 U249 ( .A1(b[10]), .A2(a[6]), .ZN(y[106]) );
  OR2_X1 U249bar ( .A1(bbar[10]), .A2(abar[6]), .ZN(ybar[106]);
  AND2_X1 U250 ( .A1(a[6]), .A2(b[9]), .ZN(y[105]) );
  OR2_X1 U250bar ( .A1(abar[6]), .A2(bbar[9]), .ZN(ybar[105]);
  AND2_X1 U251 ( .A1(b[8]), .A2(a[6]), .ZN(y[104]) );
  OR2_X1 U251bar ( .A1(bbar[8]), .A2(abar[6]), .ZN(ybar[104]);
  AND2_X1 U252 ( .A1(b[7]), .A2(a[6]), .ZN(y[103]) );
  OR2_X1 U252bar ( .A1(bbar[7]), .A2(abar[6]), .ZN(ybar[103]);
  AND2_X1 U253 ( .A1(b[6]), .A2(a[6]), .ZN(y[102]) );
  OR2_X1 U253bar ( .A1(bbar[6]), .A2(abar[6]), .ZN(ybar[102]);
  AND2_X1 U254 ( .A1(b[5]), .A2(a[6]), .ZN(y[101]) );
  OR2_X1 U254bar ( .A1(bbar[5]), .A2(abar[6]), .ZN(ybar[101]);
  AND2_X1 U255 ( .A1(b[4]), .A2(a[6]), .ZN(y[100]) );
  OR2_X1 U255bar ( .A1(bbar[4]), .A2(abar[6]), .ZN(ybar[100]);
  AND2_X1 U256 ( .A1(b[0]), .A2(a[0]), .ZN(y[0]) );
  OR2_X1 U256bar ( .A1(bbar[0]), .A2(abar[0]), .ZN(ybar[0]);
endmodule




module decode_14 ( in, out );
  input [7:0] in;
  //input_done

  output [255:0] out;
  //output_done

  wire   [15:0] level1;
  wire   [31:0] level2;
  //wire_done

  CD2_56 cd_l1_1 ( .a(in[1]), .b(in[0]), .y(level1[3:0]) );
  CD2_55 cd_l1_2 ( .a(in[3]), .b(in[2]), .y(level1[7:4]) );
  CD2_54 cd_l1_3 ( .a(in[5]), .b(in[4]), .y(level1[11:8]) );
  CD2_53 cd_l1_4 ( .a(in[7]), .b(in[6]), .y(level1[15:12]) );
  CD4_28 cd_l2_1 ( .a(level1[7:4]), .b(level1[3:0]), .y(level2[15:0]) );
  CD4_27 cd_l2_2 ( .a(level1[15:12]), .b(level1[11:8]), .y(level2[31:16]) );
  CD16_14 cd_l3 ( .a(level2[31:16]), .b(level2[15:0]), .y(out) );
endmodule


module encode_14 ( in, out );
  input [255:0] in;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
  assign inbar[8] = ~in[8];
  assign inbar[9] = ~in[9];
  assign inbar[10] = ~in[10];
  assign inbar[11] = ~in[11];
  assign inbar[12] = ~in[12];
  assign inbar[13] = ~in[13];
  assign inbar[14] = ~in[14];
  assign inbar[15] = ~in[15];
  assign inbar[16] = ~in[16];
  assign inbar[17] = ~in[17];
  assign inbar[18] = ~in[18];
  assign inbar[19] = ~in[19];
  assign inbar[20] = ~in[20];
  assign inbar[21] = ~in[21];
  assign inbar[22] = ~in[22];
  assign inbar[23] = ~in[23];
  assign inbar[24] = ~in[24];
  assign inbar[25] = ~in[25];
  assign inbar[26] = ~in[26];
  assign inbar[27] = ~in[27];
  assign inbar[28] = ~in[28];
  assign inbar[29] = ~in[29];
  assign inbar[30] = ~in[30];
  assign inbar[31] = ~in[31];
  assign inbar[32] = ~in[32];
  assign inbar[33] = ~in[33];
  assign inbar[34] = ~in[34];
  assign inbar[35] = ~in[35];
  assign inbar[36] = ~in[36];
  assign inbar[37] = ~in[37];
  assign inbar[38] = ~in[38];
  assign inbar[39] = ~in[39];
  assign inbar[40] = ~in[40];
  assign inbar[41] = ~in[41];
  assign inbar[42] = ~in[42];
  assign inbar[43] = ~in[43];
  assign inbar[44] = ~in[44];
  assign inbar[45] = ~in[45];
  assign inbar[46] = ~in[46];
  assign inbar[47] = ~in[47];
  assign inbar[48] = ~in[48];
  assign inbar[49] = ~in[49];
  assign inbar[50] = ~in[50];
  assign inbar[51] = ~in[51];
  assign inbar[52] = ~in[52];
  assign inbar[53] = ~in[53];
  assign inbar[54] = ~in[54];
  assign inbar[55] = ~in[55];
  assign inbar[56] = ~in[56];
  assign inbar[57] = ~in[57];
  assign inbar[58] = ~in[58];
  assign inbar[59] = ~in[59];
  assign inbar[60] = ~in[60];
  assign inbar[61] = ~in[61];
  assign inbar[62] = ~in[62];
  assign inbar[63] = ~in[63];
  assign inbar[64] = ~in[64];
  assign inbar[65] = ~in[65];
  assign inbar[66] = ~in[66];
  assign inbar[67] = ~in[67];
  assign inbar[68] = ~in[68];
  assign inbar[69] = ~in[69];
  assign inbar[70] = ~in[70];
  assign inbar[71] = ~in[71];
  assign inbar[72] = ~in[72];
  assign inbar[73] = ~in[73];
  assign inbar[74] = ~in[74];
  assign inbar[75] = ~in[75];
  assign inbar[76] = ~in[76];
  assign inbar[77] = ~in[77];
  assign inbar[78] = ~in[78];
  assign inbar[79] = ~in[79];
  assign inbar[80] = ~in[80];
  assign inbar[81] = ~in[81];
  assign inbar[82] = ~in[82];
  assign inbar[83] = ~in[83];
  assign inbar[84] = ~in[84];
  assign inbar[85] = ~in[85];
  assign inbar[86] = ~in[86];
  assign inbar[87] = ~in[87];
  assign inbar[88] = ~in[88];
  assign inbar[89] = ~in[89];
  assign inbar[90] = ~in[90];
  assign inbar[91] = ~in[91];
  assign inbar[92] = ~in[92];
  assign inbar[93] = ~in[93];
  assign inbar[94] = ~in[94];
  assign inbar[95] = ~in[95];
  assign inbar[96] = ~in[96];
  assign inbar[97] = ~in[97];
  assign inbar[98] = ~in[98];
  assign inbar[99] = ~in[99];
  assign inbar[100] = ~in[100];
  assign inbar[101] = ~in[101];
  assign inbar[102] = ~in[102];
  assign inbar[103] = ~in[103];
  assign inbar[104] = ~in[104];
  assign inbar[105] = ~in[105];
  assign inbar[106] = ~in[106];
  assign inbar[107] = ~in[107];
  assign inbar[108] = ~in[108];
  assign inbar[109] = ~in[109];
  assign inbar[110] = ~in[110];
  assign inbar[111] = ~in[111];
  assign inbar[112] = ~in[112];
  assign inbar[113] = ~in[113];
  assign inbar[114] = ~in[114];
  assign inbar[115] = ~in[115];
  assign inbar[116] = ~in[116];
  assign inbar[117] = ~in[117];
  assign inbar[118] = ~in[118];
  assign inbar[119] = ~in[119];
  assign inbar[120] = ~in[120];
  assign inbar[121] = ~in[121];
  assign inbar[122] = ~in[122];
  assign inbar[123] = ~in[123];
  assign inbar[124] = ~in[124];
  assign inbar[125] = ~in[125];
  assign inbar[126] = ~in[126];
  assign inbar[127] = ~in[127];
  assign inbar[128] = ~in[128];
  assign inbar[129] = ~in[129];
  assign inbar[130] = ~in[130];
  assign inbar[131] = ~in[131];
  assign inbar[132] = ~in[132];
  assign inbar[133] = ~in[133];
  assign inbar[134] = ~in[134];
  assign inbar[135] = ~in[135];
  assign inbar[136] = ~in[136];
  assign inbar[137] = ~in[137];
  assign inbar[138] = ~in[138];
  assign inbar[139] = ~in[139];
  assign inbar[140] = ~in[140];
  assign inbar[141] = ~in[141];
  assign inbar[142] = ~in[142];
  assign inbar[143] = ~in[143];
  assign inbar[144] = ~in[144];
  assign inbar[145] = ~in[145];
  assign inbar[146] = ~in[146];
  assign inbar[147] = ~in[147];
  assign inbar[148] = ~in[148];
  assign inbar[149] = ~in[149];
  assign inbar[150] = ~in[150];
  assign inbar[151] = ~in[151];
  assign inbar[152] = ~in[152];
  assign inbar[153] = ~in[153];
  assign inbar[154] = ~in[154];
  assign inbar[155] = ~in[155];
  assign inbar[156] = ~in[156];
  assign inbar[157] = ~in[157];
  assign inbar[158] = ~in[158];
  assign inbar[159] = ~in[159];
  assign inbar[160] = ~in[160];
  assign inbar[161] = ~in[161];
  assign inbar[162] = ~in[162];
  assign inbar[163] = ~in[163];
  assign inbar[164] = ~in[164];
  assign inbar[165] = ~in[165];
  assign inbar[166] = ~in[166];
  assign inbar[167] = ~in[167];
  assign inbar[168] = ~in[168];
  assign inbar[169] = ~in[169];
  assign inbar[170] = ~in[170];
  assign inbar[171] = ~in[171];
  assign inbar[172] = ~in[172];
  assign inbar[173] = ~in[173];
  assign inbar[174] = ~in[174];
  assign inbar[175] = ~in[175];
  assign inbar[176] = ~in[176];
  assign inbar[177] = ~in[177];
  assign inbar[178] = ~in[178];
  assign inbar[179] = ~in[179];
  assign inbar[180] = ~in[180];
  assign inbar[181] = ~in[181];
  assign inbar[182] = ~in[182];
  assign inbar[183] = ~in[183];
  assign inbar[184] = ~in[184];
  assign inbar[185] = ~in[185];
  assign inbar[186] = ~in[186];
  assign inbar[187] = ~in[187];
  assign inbar[188] = ~in[188];
  assign inbar[189] = ~in[189];
  assign inbar[190] = ~in[190];
  assign inbar[191] = ~in[191];
  assign inbar[192] = ~in[192];
  assign inbar[193] = ~in[193];
  assign inbar[194] = ~in[194];
  assign inbar[195] = ~in[195];
  assign inbar[196] = ~in[196];
  assign inbar[197] = ~in[197];
  assign inbar[198] = ~in[198];
  assign inbar[199] = ~in[199];
  assign inbar[200] = ~in[200];
  assign inbar[201] = ~in[201];
  assign inbar[202] = ~in[202];
  assign inbar[203] = ~in[203];
  assign inbar[204] = ~in[204];
  assign inbar[205] = ~in[205];
  assign inbar[206] = ~in[206];
  assign inbar[207] = ~in[207];
  assign inbar[208] = ~in[208];
  assign inbar[209] = ~in[209];
  assign inbar[210] = ~in[210];
  assign inbar[211] = ~in[211];
  assign inbar[212] = ~in[212];
  assign inbar[213] = ~in[213];
  assign inbar[214] = ~in[214];
  assign inbar[215] = ~in[215];
  assign inbar[216] = ~in[216];
  assign inbar[217] = ~in[217];
  assign inbar[218] = ~in[218];
  assign inbar[219] = ~in[219];
  assign inbar[220] = ~in[220];
  assign inbar[221] = ~in[221];
  assign inbar[222] = ~in[222];
  assign inbar[223] = ~in[223];
  assign inbar[224] = ~in[224];
  assign inbar[225] = ~in[225];
  assign inbar[226] = ~in[226];
  assign inbar[227] = ~in[227];
  assign inbar[228] = ~in[228];
  assign inbar[229] = ~in[229];
  assign inbar[230] = ~in[230];
  assign inbar[231] = ~in[231];
  assign inbar[232] = ~in[232];
  assign inbar[233] = ~in[233];
  assign inbar[234] = ~in[234];
  assign inbar[235] = ~in[235];
  assign inbar[236] = ~in[236];
  assign inbar[237] = ~in[237];
  assign inbar[238] = ~in[238];
  assign inbar[239] = ~in[239];
  assign inbar[240] = ~in[240];
  assign inbar[241] = ~in[241];
  assign inbar[242] = ~in[242];
  assign inbar[243] = ~in[243];
  assign inbar[244] = ~in[244];
  assign inbar[245] = ~in[245];
  assign inbar[246] = ~in[246];
  assign inbar[247] = ~in[247];
  assign inbar[248] = ~in[248];
  assign inbar[249] = ~in[249];
  assign inbar[250] = ~in[250];
  assign inbar[251] = ~in[251];
  assign inbar[252] = ~in[252];
  assign inbar[253] = ~in[253];
  assign inbar[254] = ~in[254];
  assign inbar[255] = ~in[255];
  //input_done

  output [7:0] out;
  reg [7:0] outbar;
  //output_done

  wire   in_81, in_80, in_79, in_78, in_77, in_76, in_75, in_74, in_73, in_72,
         in_71, in_70, in_69, in_68, in_67, in_66, in_65, in_64, in_63, in_62,
         in_61, in_60, in_59, in_58, in_57, in_56, in_55, in_54, in_53, in_52,
         in_51, in_50, in_49, in_48, in_47, in_46, in_45, in_44, in_43, in_42,
         in_41, in_40, in_39, in_38, in_37, in_36, in_35, in_34, in_33, in_32,
         in_31, in_30, in_29, in_28, in_27, in_26, in_25, in_24, in_23, in_22,
         in_21, in_20, in_19, in_18, in_17, in_16, in_15, in_14, in_13, in_12,
         in_11, in_10, in_9, in_8, in_7, in_6, in_5, in_4, in_3, in_2, in_1,
         in_0, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972;
  wire in_81bar, in_80bar, in_79bar, in_78bar, in_77bar, in_76bar, in_75bar, in_74bar, in_73bar, in_72bar, in_71bar, in_70bar, in_69bar, in_68bar, in_67bar, in_66bar, in_65bar, in_64bar, in_63bar, in_62bar, in_61bar, in_60bar, in_59bar, in_58bar, in_57bar, in_56bar, in_55bar, in_54bar, in_53bar, in_52bar, in_51bar, in_50bar, in_49bar, in_48bar, in_47bar, in_46bar, in_45bar, in_44bar, in_43bar, in_42bar, in_41bar, in_40bar, in_39bar, in_38bar, in_37bar, in_36bar, in_35bar, in_34bar, in_33bar, in_32bar, in_31bar, in_30bar, in_29bar, in_28bar, in_27bar, in_26bar, in_25bar, in_24bar, in_23bar, in_22bar, in_21bar, in_20bar, in_19bar, in_18bar, in_17bar, in_16bar, in_15bar, in_14bar, in_13bar, in_12bar, in_11bar, in_10bar, in_9bar, in_8bar, in_7bar, in_6bar, in_5bar, in_4bar, in_3bar, in_2bar, in_1bar, in_0bar, n487bar, n488bar, n489bar, n490bar, n491bar, n492bar, n493bar, n494bar, n495bar, n496bar, n497bar, n498bar, n499bar, n500bar, n501bar, n502bar, n503bar, n504bar, n505bar, n506bar, n507bar, n508bar, n509bar, n510bar, n511bar, n512bar, n513bar, n514bar, n515bar, n516bar, n517bar, n518bar, n519bar, n520bar, n521bar, n522bar, n523bar, n524bar, n525bar, n526bar, n527bar, n528bar, n529bar, n530bar, n531bar, n532bar, n533bar, n534bar, n535bar, n536bar, n537bar, n538bar, n539bar, n540bar, n541bar, n542bar, n543bar, n544bar, n545bar, n546bar, n547bar, n548bar, n549bar, n550bar, n551bar, n552bar, n553bar, n554bar, n555bar, n556bar, n557bar, n558bar, n559bar, n560bar, n561bar, n562bar, n563bar, n564bar, n565bar, n566bar, n567bar, n568bar, n569bar, n570bar, n571bar, n572bar, n573bar, n574bar, n575bar, n576bar, n577bar, n578bar, n579bar, n580bar, n581bar, n582bar, n583bar, n584bar, n585bar, n586bar, n587bar, n588bar, n589bar, n590bar, n591bar, n592bar, n593bar, n594bar, n595bar, n596bar, n597bar, n598bar, n599bar, n600bar, n601bar, n602bar, n603bar, n604bar, n605bar, n606bar, n607bar, n608bar, n609bar, n610bar, n611bar, n612bar, n613bar, n614bar, n615bar, n616bar, n617bar, n618bar, n619bar, n620bar, n621bar, n622bar, n623bar, n624bar, n625bar, n626bar, n627bar, n628bar, n629bar, n630bar, n631bar, n632bar, n633bar, n634bar, n635bar, n636bar, n637bar, n638bar, n639bar, n640bar, n641bar, n642bar, n643bar, n644bar, n645bar, n646bar, n647bar, n648bar, n649bar, n650bar, n651bar, n652bar, n653bar, n654bar, n655bar, n656bar, n657bar, n658bar, n659bar, n660bar, n661bar, n662bar, n663bar, n664bar, n665bar, n666bar, n667bar, n668bar, n669bar, n670bar, n671bar, n672bar, n673bar, n674bar, n675bar, n676bar, n677bar, n678bar, n679bar, n680bar, n681bar, n682bar, n683bar, n684bar, n685bar, n686bar, n687bar, n688bar, n689bar, n690bar, n691bar, n692bar, n693bar, n694bar, n695bar, n696bar, n697bar, n698bar, n699bar, n700bar, n701bar, n702bar, n703bar, n704bar, n705bar, n706bar, n707bar, n708bar, n709bar, n710bar, n711bar, n712bar, n713bar, n714bar, n715bar, n716bar, n717bar, n718bar, n719bar, n720bar, n721bar, n722bar, n723bar, n724bar, n725bar, n726bar, n727bar, n728bar, n729bar, n730bar, n731bar, n732bar, n733bar, n734bar, n735bar, n736bar, n737bar, n738bar, n739bar, n740bar, n741bar, n742bar, n743bar, n744bar, n745bar, n746bar, n747bar, n748bar, n749bar, n750bar, n751bar, n752bar, n753bar, n754bar, n755bar, n756bar, n757bar, n758bar, n759bar, n760bar, n761bar, n762bar, n763bar, n764bar, n765bar, n766bar, n767bar, n768bar, n769bar, n770bar, n771bar, n772bar, n773bar, n774bar, n775bar, n776bar, n777bar, n778bar, n779bar, n780bar, n781bar, n782bar, n783bar, n784bar, n785bar, n786bar, n787bar, n788bar, n789bar, n790bar, n791bar, n792bar, n793bar, n794bar, n795bar, n796bar, n797bar, n798bar, n799bar, n800bar, n801bar, n802bar, n803bar, n804bar, n805bar, n806bar, n807bar, n808bar, n809bar, n810bar, n811bar, n812bar, n813bar, n814bar, n815bar, n816bar, n817bar, n818bar, n819bar, n820bar, n821bar, n822bar, n823bar, n824bar, n825bar, n826bar, n827bar, n828bar, n829bar, n830bar, n831bar, n832bar, n833bar, n834bar, n835bar, n836bar, n837bar, n838bar, n839bar, n840bar, n841bar, n842bar, n843bar, n844bar, n845bar, n846bar, n847bar, n848bar, n849bar, n850bar, n851bar, n852bar, n853bar, n854bar, n855bar, n856bar, n857bar, n858bar, n859bar, n860bar, n861bar, n862bar, n863bar, n864bar, n865bar, n866bar, n867bar, n868bar, n869bar, n870bar, n871bar, n872bar, n873bar, n874bar, n875bar, n876bar, n877bar, n878bar, n879bar, n880bar, n881bar, n882bar, n883bar, n884bar, n885bar, n886bar, n887bar, n888bar, n889bar, n890bar, n891bar, n892bar, n893bar, n894bar, n895bar, n896bar, n897bar, n898bar, n899bar, n900bar, n901bar, n902bar, n903bar, n904bar, n905bar, n906bar, n907bar, n908bar, n909bar, n910bar, n911bar, n912bar, n913bar, n914bar, n915bar, n916bar, n917bar, n918bar, n919bar, n920bar, n921bar, n922bar, n923bar, n924bar, n925bar, n926bar, n927bar, n928bar, n929bar, n930bar, n931bar, n932bar, n933bar, n934bar, n935bar, n936bar, n937bar, n938bar, n939bar, n940bar, n941bar, n942bar, n943bar, n944bar, n945bar, n946bar, n947bar, n948bar, n949bar, n950bar, n951bar, n952bar, n953bar, n954bar, n955bar, n956bar, n957bar, n958bar, n959bar, n960bar, n961bar, n962bar, n963bar, n964bar, n965bar, n966bar, n967bar, n968bar, n969bar, n970bar, n971bar, n972bar;
  //wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];

  OR2_X1 U1 ( .A1(n972), .A2(n971), .ZN(out[7]) );
  AND2_X1 U1bar ( .A1(n972bar), .A2(n971bar), .ZN(outbar[7]);
  OR2_X1 U2 ( .A1(n970), .A2(n969), .ZN(n971) );
  AND2_X1 U2bar ( .A1(n970bar), .A2(n969bar), .ZN(n971bar);
  OR2_X1 U3 ( .A1(n968), .A2(n967), .ZN(n969) );
  AND2_X1 U3bar ( .A1(n968bar), .A2(n967bar), .ZN(n969bar);
  OR2_X1 U4 ( .A1(n966), .A2(n965), .ZN(n967) );
  AND2_X1 U4bar ( .A1(n966bar), .A2(n965bar), .ZN(n967bar);
  OR2_X1 U5 ( .A1(n964), .A2(n963), .ZN(n968) );
  AND2_X1 U5bar ( .A1(n964bar), .A2(n963bar), .ZN(n968bar);
  OR2_X1 U6 ( .A1(in[116]), .A2(n962), .ZN(n963) );
  AND2_X1 U6bar ( .A1(inbar[116]), .A2(n962bar), .ZN(n963bar);
  OR2_X1 U7 ( .A1(n961), .A2(n960), .ZN(n970) );
  AND2_X1 U7bar ( .A1(n961bar), .A2(n960bar), .ZN(n970bar);
  OR2_X1 U8 ( .A1(in[150]), .A2(in[127]), .ZN(n960) );
  AND2_X1 U8bar ( .A1(inbar[150]), .A2(inbar[127]), .ZN(n960bar);
  OR2_X1 U9 ( .A1(in[160]), .A2(n959), .ZN(n961) );
  AND2_X1 U9bar ( .A1(inbar[160]), .A2(n959bar), .ZN(n961bar);
  OR2_X1 U10 ( .A1(in[252]), .A2(in[168]), .ZN(n959) );
  AND2_X1 U10bar ( .A1(inbar[252]), .A2(inbar[168]), .ZN(n959bar);
  OR2_X1 U11 ( .A1(n958), .A2(n957), .ZN(n972) );
  AND2_X1 U11bar ( .A1(n958bar), .A2(n957bar), .ZN(n972bar);
  OR2_X1 U12 ( .A1(n956), .A2(n955), .ZN(n957) );
  AND2_X1 U12bar ( .A1(n956bar), .A2(n955bar), .ZN(n957bar);
  OR2_X1 U13 ( .A1(in_17), .A2(in[96]), .ZN(n955) );
  AND2_X1 U13bar ( .A1(in_17bar), .A2(inbar[96]), .ZN(n955bar);
  OR2_X1 U14 ( .A1(in_23), .A2(n954), .ZN(n956) );
  AND2_X1 U14bar ( .A1(in_23bar), .A2(n954bar), .ZN(n956bar);
  OR2_X1 U15 ( .A1(in_31), .A2(in_26), .ZN(n954) );
  AND2_X1 U15bar ( .A1(in_31bar), .A2(in_26bar), .ZN(n954bar);
  OR2_X1 U16 ( .A1(n953), .A2(n952), .ZN(n958) );
  AND2_X1 U16bar ( .A1(n953bar), .A2(n952bar), .ZN(n958bar);
  OR2_X1 U17 ( .A1(in_58), .A2(in_4), .ZN(n952) );
  AND2_X1 U17bar ( .A1(in_58bar), .A2(in_4bar), .ZN(n952bar);
  OR2_X1 U18 ( .A1(in_59), .A2(n951), .ZN(n953) );
  AND2_X1 U18bar ( .A1(in_59bar), .A2(n951bar), .ZN(n953bar);
  OR2_X1 U19 ( .A1(in_71), .A2(in_62), .ZN(n951) );
  AND2_X1 U19bar ( .A1(in_71bar), .A2(in_62bar), .ZN(n951bar);
  OR2_X1 U20 ( .A1(n950), .A2(n949), .ZN(out[6]) );
  AND2_X1 U20bar ( .A1(n950bar), .A2(n949bar), .ZN(outbar[6]);
  OR2_X1 U21 ( .A1(n948), .A2(n947), .ZN(n949) );
  AND2_X1 U21bar ( .A1(n948bar), .A2(n947bar), .ZN(n949bar);
  OR2_X1 U22 ( .A1(n946), .A2(n945), .ZN(n947) );
  AND2_X1 U22bar ( .A1(n946bar), .A2(n945bar), .ZN(n947bar);
  OR2_X1 U23 ( .A1(n944), .A2(n943), .ZN(n945) );
  AND2_X1 U23bar ( .A1(n944bar), .A2(n943bar), .ZN(n945bar);
  OR2_X1 U24 ( .A1(n942), .A2(n941), .ZN(n946) );
  AND2_X1 U24bar ( .A1(n942bar), .A2(n941bar), .ZN(n946bar);
  OR2_X1 U25 ( .A1(in[101]), .A2(n940), .ZN(n941) );
  AND2_X1 U25bar ( .A1(inbar[101]), .A2(n940bar), .ZN(n941bar);
  OR2_X1 U26 ( .A1(n939), .A2(n938), .ZN(n948) );
  AND2_X1 U26bar ( .A1(n939bar), .A2(n938bar), .ZN(n948bar);
  OR2_X1 U27 ( .A1(in[114]), .A2(in[104]), .ZN(n938) );
  AND2_X1 U27bar ( .A1(inbar[114]), .A2(inbar[104]), .ZN(n938bar);
  OR2_X1 U28 ( .A1(in[128]), .A2(n937), .ZN(n939) );
  AND2_X1 U28bar ( .A1(inbar[128]), .A2(n937bar), .ZN(n939bar);
  OR2_X1 U29 ( .A1(in[136]), .A2(in[134]), .ZN(n937) );
  AND2_X1 U29bar ( .A1(inbar[136]), .A2(inbar[134]), .ZN(n937bar);
  OR2_X1 U30 ( .A1(n936), .A2(n935), .ZN(n950) );
  AND2_X1 U30bar ( .A1(n936bar), .A2(n935bar), .ZN(n950bar);
  OR2_X1 U31 ( .A1(n934), .A2(n933), .ZN(n935) );
  AND2_X1 U31bar ( .A1(n934bar), .A2(n933bar), .ZN(n935bar);
  OR2_X1 U32 ( .A1(in[177]), .A2(in[164]), .ZN(n933) );
  AND2_X1 U32bar ( .A1(inbar[177]), .A2(inbar[164]), .ZN(n933bar);
  OR2_X1 U33 ( .A1(in[212]), .A2(n932), .ZN(n934) );
  AND2_X1 U33bar ( .A1(inbar[212]), .A2(n932bar), .ZN(n934bar);
  OR2_X1 U34 ( .A1(in[248]), .A2(in[221]), .ZN(n932) );
  AND2_X1 U34bar ( .A1(inbar[248]), .A2(inbar[221]), .ZN(n932bar);
  OR2_X1 U35 ( .A1(n931), .A2(n930), .ZN(n936) );
  AND2_X1 U35bar ( .A1(n931bar), .A2(n930bar), .ZN(n936bar);
  OR2_X1 U36 ( .A1(in_18), .A2(in[93]), .ZN(n930) );
  AND2_X1 U36bar ( .A1(in_18bar), .A2(inbar[93]), .ZN(n930bar);
  OR2_X1 U37 ( .A1(in_31), .A2(n929), .ZN(n931) );
  AND2_X1 U37bar ( .A1(in_31bar), .A2(n929bar), .ZN(n931bar);
  OR2_X1 U38 ( .A1(in_7), .A2(in_39), .ZN(n929) );
  AND2_X1 U38bar ( .A1(in_7bar), .A2(in_39bar), .ZN(n929bar);
  OR2_X1 U39 ( .A1(n928), .A2(n927), .ZN(out[5]) );
  AND2_X1 U39bar ( .A1(n928bar), .A2(n927bar), .ZN(outbar[5]);
  OR2_X1 U40 ( .A1(n926), .A2(n925), .ZN(n927) );
  AND2_X1 U40bar ( .A1(n926bar), .A2(n925bar), .ZN(n927bar);
  OR2_X1 U41 ( .A1(n924), .A2(n923), .ZN(n925) );
  AND2_X1 U41bar ( .A1(n924bar), .A2(n923bar), .ZN(n925bar);
  OR2_X1 U42 ( .A1(n922), .A2(n921), .ZN(n923) );
  AND2_X1 U42bar ( .A1(n922bar), .A2(n921bar), .ZN(n923bar);
  OR2_X1 U43 ( .A1(n940), .A2(n920), .ZN(n924) );
  AND2_X1 U43bar ( .A1(n940bar), .A2(n920bar), .ZN(n924bar);
  OR2_X1 U44 ( .A1(in[111]), .A2(n919), .ZN(n920) );
  AND2_X1 U44bar ( .A1(inbar[111]), .A2(n919bar), .ZN(n920bar);
  OR2_X1 U45 ( .A1(n918), .A2(n917), .ZN(n940) );
  AND2_X1 U45bar ( .A1(n918bar), .A2(n917bar), .ZN(n940bar);
  OR2_X1 U46 ( .A1(n916), .A2(n915), .ZN(n917) );
  AND2_X1 U46bar ( .A1(n916bar), .A2(n915bar), .ZN(n917bar);
  OR2_X1 U47 ( .A1(n914), .A2(n913), .ZN(n915) );
  AND2_X1 U47bar ( .A1(n914bar), .A2(n913bar), .ZN(n915bar);
  OR2_X1 U48 ( .A1(in[140]), .A2(in[131]), .ZN(n913) );
  AND2_X1 U48bar ( .A1(inbar[140]), .A2(inbar[131]), .ZN(n913bar);
  OR2_X1 U49 ( .A1(in[160]), .A2(in[144]), .ZN(n914) );
  AND2_X1 U49bar ( .A1(inbar[160]), .A2(inbar[144]), .ZN(n914bar);
  OR2_X1 U50 ( .A1(n912), .A2(n911), .ZN(n916) );
  AND2_X1 U50bar ( .A1(n912bar), .A2(n911bar), .ZN(n916bar);
  OR2_X1 U51 ( .A1(in[179]), .A2(in[174]), .ZN(n911) );
  AND2_X1 U51bar ( .A1(inbar[179]), .A2(inbar[174]), .ZN(n911bar);
  OR2_X1 U52 ( .A1(in[188]), .A2(in[184]), .ZN(n912) );
  AND2_X1 U52bar ( .A1(inbar[188]), .A2(inbar[184]), .ZN(n912bar);
  OR2_X1 U53 ( .A1(n910), .A2(n909), .ZN(n918) );
  AND2_X1 U53bar ( .A1(n910bar), .A2(n909bar), .ZN(n918bar);
  OR2_X1 U54 ( .A1(n908), .A2(n907), .ZN(n909) );
  AND2_X1 U54bar ( .A1(n908bar), .A2(n907bar), .ZN(n909bar);
  OR2_X1 U55 ( .A1(in[216]), .A2(in[200]), .ZN(n907) );
  AND2_X1 U55bar ( .A1(inbar[216]), .A2(inbar[200]), .ZN(n907bar);
  OR2_X1 U56 ( .A1(in[228]), .A2(in[224]), .ZN(n908) );
  AND2_X1 U56bar ( .A1(inbar[228]), .A2(inbar[224]), .ZN(n908bar);
  OR2_X1 U57 ( .A1(n906), .A2(n905), .ZN(n910) );
  AND2_X1 U57bar ( .A1(n906bar), .A2(n905bar), .ZN(n910bar);
  OR2_X1 U58 ( .A1(in[247]), .A2(in[235]), .ZN(n905) );
  AND2_X1 U58bar ( .A1(inbar[247]), .A2(inbar[235]), .ZN(n905bar);
  OR2_X1 U59 ( .A1(in_42), .A2(in[83]), .ZN(n906) );
  AND2_X1 U59bar ( .A1(in_42bar), .A2(inbar[83]), .ZN(n906bar);
  OR2_X1 U60 ( .A1(n904), .A2(n903), .ZN(n926) );
  AND2_X1 U60bar ( .A1(n904bar), .A2(n903bar), .ZN(n926bar);
  OR2_X1 U61 ( .A1(in[166]), .A2(in[123]), .ZN(n903) );
  AND2_X1 U61bar ( .A1(inbar[166]), .A2(inbar[123]), .ZN(n903bar);
  OR2_X1 U62 ( .A1(in[170]), .A2(n902), .ZN(n904) );
  AND2_X1 U62bar ( .A1(inbar[170]), .A2(n902bar), .ZN(n904bar);
  OR2_X1 U63 ( .A1(in[194]), .A2(in[183]), .ZN(n902) );
  AND2_X1 U63bar ( .A1(inbar[194]), .A2(inbar[183]), .ZN(n902bar);
  OR2_X1 U64 ( .A1(n901), .A2(n900), .ZN(n928) );
  AND2_X1 U64bar ( .A1(n901bar), .A2(n900bar), .ZN(n928bar);
  OR2_X1 U65 ( .A1(n899), .A2(n898), .ZN(n900) );
  AND2_X1 U65bar ( .A1(n899bar), .A2(n898bar), .ZN(n900bar);
  OR2_X1 U66 ( .A1(in[241]), .A2(in[238]), .ZN(n898) );
  AND2_X1 U66bar ( .A1(inbar[241]), .A2(inbar[238]), .ZN(n898bar);
  OR2_X1 U67 ( .A1(in[250]), .A2(n897), .ZN(n899) );
  AND2_X1 U67bar ( .A1(inbar[250]), .A2(n897bar), .ZN(n899bar);
  OR2_X1 U68 ( .A1(in_24), .A2(in[84]), .ZN(n897) );
  AND2_X1 U68bar ( .A1(in_24bar), .A2(inbar[84]), .ZN(n897bar);
  OR2_X1 U69 ( .A1(n896), .A2(n895), .ZN(n901) );
  AND2_X1 U69bar ( .A1(n896bar), .A2(n895bar), .ZN(n901bar);
  OR2_X1 U70 ( .A1(in_41), .A2(in_29), .ZN(n895) );
  AND2_X1 U70bar ( .A1(in_41bar), .A2(in_29bar), .ZN(n895bar);
  OR2_X1 U71 ( .A1(in_66), .A2(n894), .ZN(n896) );
  AND2_X1 U71bar ( .A1(in_66bar), .A2(n894bar), .ZN(n896bar);
  OR2_X1 U72 ( .A1(in_76), .A2(in_71), .ZN(n894) );
  AND2_X1 U72bar ( .A1(in_76bar), .A2(in_71bar), .ZN(n894bar);
  OR2_X1 U73 ( .A1(n893), .A2(n892), .ZN(out[4]) );
  AND2_X1 U73bar ( .A1(n893bar), .A2(n892bar), .ZN(outbar[4]);
  OR2_X1 U74 ( .A1(n891), .A2(n890), .ZN(n892) );
  AND2_X1 U74bar ( .A1(n891bar), .A2(n890bar), .ZN(n892bar);
  OR2_X1 U75 ( .A1(n889), .A2(n888), .ZN(n890) );
  AND2_X1 U75bar ( .A1(n889bar), .A2(n888bar), .ZN(n890bar);
  OR2_X1 U76 ( .A1(n922), .A2(n887), .ZN(n888) );
  AND2_X1 U76bar ( .A1(n922bar), .A2(n887bar), .ZN(n888bar);
  OR2_X1 U77 ( .A1(n886), .A2(n885), .ZN(n922) );
  AND2_X1 U77bar ( .A1(n886bar), .A2(n885bar), .ZN(n922bar);
  OR2_X1 U78 ( .A1(n884), .A2(n883), .ZN(n885) );
  AND2_X1 U78bar ( .A1(n884bar), .A2(n883bar), .ZN(n885bar);
  OR2_X1 U79 ( .A1(n882), .A2(n881), .ZN(n883) );
  AND2_X1 U79bar ( .A1(n882bar), .A2(n881bar), .ZN(n883bar);
  OR2_X1 U80 ( .A1(in[118]), .A2(in[109]), .ZN(n881) );
  AND2_X1 U80bar ( .A1(inbar[118]), .A2(inbar[109]), .ZN(n881bar);
  OR2_X1 U81 ( .A1(in[139]), .A2(in[120]), .ZN(n882) );
  AND2_X1 U81bar ( .A1(inbar[139]), .A2(inbar[120]), .ZN(n882bar);
  OR2_X1 U82 ( .A1(n880), .A2(n879), .ZN(n884) );
  AND2_X1 U82bar ( .A1(n880bar), .A2(n879bar), .ZN(n884bar);
  OR2_X1 U83 ( .A1(in[198]), .A2(in[154]), .ZN(n879) );
  AND2_X1 U83bar ( .A1(inbar[198]), .A2(inbar[154]), .ZN(n879bar);
  OR2_X1 U84 ( .A1(in[210]), .A2(in[205]), .ZN(n880) );
  AND2_X1 U84bar ( .A1(inbar[210]), .A2(inbar[205]), .ZN(n880bar);
  OR2_X1 U85 ( .A1(n878), .A2(n877), .ZN(n886) );
  AND2_X1 U85bar ( .A1(n878bar), .A2(n877bar), .ZN(n886bar);
  OR2_X1 U86 ( .A1(n876), .A2(n875), .ZN(n877) );
  AND2_X1 U86bar ( .A1(n876bar), .A2(n875bar), .ZN(n877bar);
  OR2_X1 U87 ( .A1(in[219]), .A2(in[217]), .ZN(n875) );
  AND2_X1 U87bar ( .A1(inbar[219]), .A2(inbar[217]), .ZN(n875bar);
  OR2_X1 U88 ( .A1(in[86]), .A2(in[252]), .ZN(n876) );
  AND2_X1 U88bar ( .A1(inbar[86]), .A2(inbar[252]), .ZN(n876bar);
  OR2_X1 U89 ( .A1(n874), .A2(n873), .ZN(n878) );
  AND2_X1 U89bar ( .A1(n874bar), .A2(n873bar), .ZN(n878bar);
  OR2_X1 U90 ( .A1(in_40), .A2(in[91]), .ZN(n873) );
  AND2_X1 U90bar ( .A1(in_40bar), .A2(inbar[91]), .ZN(n873bar);
  OR2_X1 U91 ( .A1(in_8), .A2(in_46), .ZN(n874) );
  AND2_X1 U91bar ( .A1(in_8bar), .A2(in_46bar), .ZN(n874bar);
  OR2_X1 U92 ( .A1(n872), .A2(n871), .ZN(n889) );
  AND2_X1 U92bar ( .A1(n872bar), .A2(n871bar), .ZN(n889bar);
  OR2_X1 U93 ( .A1(in[117]), .A2(n943), .ZN(n871) );
  AND2_X1 U93bar ( .A1(inbar[117]), .A2(n943bar), .ZN(n871bar);
  OR2_X1 U94 ( .A1(n870), .A2(n869), .ZN(n943) );
  AND2_X1 U94bar ( .A1(n870bar), .A2(n869bar), .ZN(n943bar);
  OR2_X1 U95 ( .A1(n868), .A2(n867), .ZN(n869) );
  AND2_X1 U95bar ( .A1(n868bar), .A2(n867bar), .ZN(n869bar);
  OR2_X1 U96 ( .A1(n866), .A2(n865), .ZN(n867) );
  AND2_X1 U96bar ( .A1(n866bar), .A2(n865bar), .ZN(n867bar);
  OR2_X1 U97 ( .A1(n864), .A2(n863), .ZN(n865) );
  AND2_X1 U97bar ( .A1(n864bar), .A2(n863bar), .ZN(n865bar);
  OR2_X1 U98 ( .A1(in[108]), .A2(n919), .ZN(n866) );
  AND2_X1 U98bar ( .A1(inbar[108]), .A2(n919bar), .ZN(n866bar);
  OR2_X1 U99 ( .A1(n862), .A2(n861), .ZN(n919) );
  AND2_X1 U99bar ( .A1(n862bar), .A2(n861bar), .ZN(n919bar);
  OR2_X1 U100 ( .A1(n860), .A2(n859), .ZN(n861) );
  AND2_X1 U100bar ( .A1(n860bar), .A2(n859bar), .ZN(n861bar);
  OR2_X1 U101 ( .A1(n858), .A2(n857), .ZN(n859) );
  AND2_X1 U101bar ( .A1(n858bar), .A2(n857bar), .ZN(n859bar);
  OR2_X1 U102 ( .A1(in[119]), .A2(in[105]), .ZN(n857) );
  AND2_X1 U102bar ( .A1(inbar[119]), .A2(inbar[105]), .ZN(n857bar);
  OR2_X1 U103 ( .A1(in[186]), .A2(in[175]), .ZN(n858) );
  AND2_X1 U103bar ( .A1(inbar[186]), .A2(inbar[175]), .ZN(n858bar);
  OR2_X1 U104 ( .A1(n856), .A2(n855), .ZN(n860) );
  AND2_X1 U104bar ( .A1(n856bar), .A2(n855bar), .ZN(n860bar);
  OR2_X1 U105 ( .A1(in[202]), .A2(in[193]), .ZN(n855) );
  AND2_X1 U105bar ( .A1(inbar[202]), .A2(inbar[193]), .ZN(n855bar);
  OR2_X1 U106 ( .A1(in[225]), .A2(in[208]), .ZN(n856) );
  AND2_X1 U106bar ( .A1(inbar[225]), .A2(inbar[208]), .ZN(n856bar);
  OR2_X1 U107 ( .A1(n854), .A2(n853), .ZN(n862) );
  AND2_X1 U107bar ( .A1(n854bar), .A2(n853bar), .ZN(n862bar);
  OR2_X1 U108 ( .A1(n852), .A2(n851), .ZN(n853) );
  AND2_X1 U108bar ( .A1(n852bar), .A2(n851bar), .ZN(n853bar);
  OR2_X1 U109 ( .A1(in_1), .A2(in[85]), .ZN(n851) );
  AND2_X1 U109bar ( .A1(in_1bar), .A2(inbar[85]), .ZN(n851bar);
  OR2_X1 U110 ( .A1(in_23), .A2(in_19), .ZN(n852) );
  AND2_X1 U110bar ( .A1(in_23bar), .A2(in_19bar), .ZN(n852bar);
  OR2_X1 U111 ( .A1(n850), .A2(n849), .ZN(n854) );
  AND2_X1 U111bar ( .A1(n850bar), .A2(n849bar), .ZN(n854bar);
  OR2_X1 U112 ( .A1(in_43), .A2(in_33), .ZN(n849) );
  AND2_X1 U112bar ( .A1(in_43bar), .A2(in_33bar), .ZN(n849bar);
  OR2_X1 U113 ( .A1(in_63), .A2(in_44), .ZN(n850) );
  AND2_X1 U113bar ( .A1(in_63bar), .A2(in_44bar), .ZN(n850bar);
  OR2_X1 U114 ( .A1(n848), .A2(n847), .ZN(n868) );
  AND2_X1 U114bar ( .A1(n848bar), .A2(n847bar), .ZN(n868bar);
  OR2_X1 U115 ( .A1(in[141]), .A2(in[112]), .ZN(n847) );
  AND2_X1 U115bar ( .A1(inbar[141]), .A2(inbar[112]), .ZN(n847bar);
  OR2_X1 U116 ( .A1(in[147]), .A2(n846), .ZN(n848) );
  AND2_X1 U116bar ( .A1(inbar[147]), .A2(n846bar), .ZN(n848bar);
  OR2_X1 U117 ( .A1(in[181]), .A2(in[167]), .ZN(n846) );
  AND2_X1 U117bar ( .A1(inbar[181]), .A2(inbar[167]), .ZN(n846bar);
  OR2_X1 U118 ( .A1(n845), .A2(n844), .ZN(n870) );
  AND2_X1 U118bar ( .A1(n845bar), .A2(n844bar), .ZN(n870bar);
  OR2_X1 U119 ( .A1(n843), .A2(n842), .ZN(n844) );
  AND2_X1 U119bar ( .A1(n843bar), .A2(n842bar), .ZN(n844bar);
  OR2_X1 U120 ( .A1(in[229]), .A2(in[201]), .ZN(n842) );
  AND2_X1 U120bar ( .A1(inbar[229]), .A2(inbar[201]), .ZN(n842bar);
  OR2_X1 U121 ( .A1(in[237]), .A2(n841), .ZN(n843) );
  AND2_X1 U121bar ( .A1(inbar[237]), .A2(n841bar), .ZN(n843bar);
  OR2_X1 U122 ( .A1(in[94]), .A2(in[253]), .ZN(n841) );
  AND2_X1 U122bar ( .A1(inbar[94]), .A2(inbar[253]), .ZN(n841bar);
  OR2_X1 U123 ( .A1(n840), .A2(n839), .ZN(n845) );
  AND2_X1 U123bar ( .A1(n840bar), .A2(n839bar), .ZN(n845bar);
  OR2_X1 U124 ( .A1(in_21), .A2(in[96]), .ZN(n839) );
  AND2_X1 U124bar ( .A1(in_21bar), .A2(inbar[96]), .ZN(n839bar);
  OR2_X1 U125 ( .A1(in_25), .A2(n838), .ZN(n840) );
  AND2_X1 U125bar ( .A1(in_25bar), .A2(n838bar), .ZN(n840bar);
  OR2_X1 U126 ( .A1(in_81), .A2(in_45), .ZN(n838) );
  AND2_X1 U126bar ( .A1(in_81bar), .A2(in_45bar), .ZN(n838bar);
  OR2_X1 U127 ( .A1(n837), .A2(n836), .ZN(n891) );
  AND2_X1 U127bar ( .A1(n837bar), .A2(n836bar), .ZN(n891bar);
  OR2_X1 U128 ( .A1(in[142]), .A2(in[124]), .ZN(n836) );
  AND2_X1 U128bar ( .A1(inbar[142]), .A2(inbar[124]), .ZN(n836bar);
  OR2_X1 U129 ( .A1(in[150]), .A2(n835), .ZN(n837) );
  AND2_X1 U129bar ( .A1(inbar[150]), .A2(n835bar), .ZN(n837bar);
  OR2_X1 U130 ( .A1(in[172]), .A2(in[155]), .ZN(n835) );
  AND2_X1 U130bar ( .A1(inbar[172]), .A2(inbar[155]), .ZN(n835bar);
  OR2_X1 U131 ( .A1(n834), .A2(n833), .ZN(n893) );
  AND2_X1 U131bar ( .A1(n834bar), .A2(n833bar), .ZN(n893bar);
  OR2_X1 U132 ( .A1(n832), .A2(n831), .ZN(n833) );
  AND2_X1 U132bar ( .A1(n832bar), .A2(n831bar), .ZN(n833bar);
  OR2_X1 U133 ( .A1(in[196]), .A2(in[173]), .ZN(n831) );
  AND2_X1 U133bar ( .A1(inbar[196]), .A2(inbar[173]), .ZN(n831bar);
  OR2_X1 U134 ( .A1(in[222]), .A2(n830), .ZN(n832) );
  AND2_X1 U134bar ( .A1(inbar[222]), .A2(n830bar), .ZN(n832bar);
  OR2_X1 U135 ( .A1(in[227]), .A2(in[226]), .ZN(n830) );
  AND2_X1 U135bar ( .A1(inbar[227]), .A2(inbar[226]), .ZN(n830bar);
  OR2_X1 U136 ( .A1(n829), .A2(n828), .ZN(n834) );
  AND2_X1 U136bar ( .A1(n829bar), .A2(n828bar), .ZN(n834bar);
  OR2_X1 U137 ( .A1(in[249]), .A2(in[231]), .ZN(n828) );
  AND2_X1 U137bar ( .A1(inbar[249]), .A2(inbar[231]), .ZN(n828bar);
  OR2_X1 U138 ( .A1(in_28), .A2(n827), .ZN(n829) );
  AND2_X1 U138bar ( .A1(in_28bar), .A2(n827bar), .ZN(n829bar);
  OR2_X1 U139 ( .A1(in_52), .A2(in_47), .ZN(n827) );
  AND2_X1 U139bar ( .A1(in_52bar), .A2(in_47bar), .ZN(n827bar);
  OR2_X1 U140 ( .A1(n826), .A2(n825), .ZN(out[3]) );
  AND2_X1 U140bar ( .A1(n826bar), .A2(n825bar), .ZN(outbar[3]);
  OR2_X1 U141 ( .A1(n824), .A2(n823), .ZN(n825) );
  AND2_X1 U141bar ( .A1(n824bar), .A2(n823bar), .ZN(n825bar);
  OR2_X1 U142 ( .A1(n822), .A2(n821), .ZN(n823) );
  AND2_X1 U142bar ( .A1(n822bar), .A2(n821bar), .ZN(n823bar);
  OR2_X1 U143 ( .A1(n820), .A2(n819), .ZN(n821) );
  AND2_X1 U143bar ( .A1(n820bar), .A2(n819bar), .ZN(n821bar);
  OR2_X1 U144 ( .A1(n964), .A2(n818), .ZN(n822) );
  AND2_X1 U144bar ( .A1(n964bar), .A2(n818bar), .ZN(n822bar);
  OR2_X1 U145 ( .A1(in[118]), .A2(n817), .ZN(n818) );
  AND2_X1 U145bar ( .A1(inbar[118]), .A2(n817bar), .ZN(n818bar);
  OR2_X1 U146 ( .A1(n816), .A2(n815), .ZN(n964) );
  AND2_X1 U146bar ( .A1(n816bar), .A2(n815bar), .ZN(n964bar);
  OR2_X1 U147 ( .A1(n814), .A2(n813), .ZN(n815) );
  AND2_X1 U147bar ( .A1(n814bar), .A2(n813bar), .ZN(n815bar);
  OR2_X1 U148 ( .A1(n812), .A2(n811), .ZN(n813) );
  AND2_X1 U148bar ( .A1(n812bar), .A2(n811bar), .ZN(n813bar);
  OR2_X1 U149 ( .A1(in[122]), .A2(in[111]), .ZN(n811) );
  AND2_X1 U149bar ( .A1(inbar[122]), .A2(inbar[111]), .ZN(n811bar);
  OR2_X1 U150 ( .A1(in[154]), .A2(in[151]), .ZN(n812) );
  AND2_X1 U150bar ( .A1(inbar[154]), .A2(inbar[151]), .ZN(n812bar);
  OR2_X1 U151 ( .A1(n810), .A2(n809), .ZN(n814) );
  AND2_X1 U151bar ( .A1(n810bar), .A2(n809bar), .ZN(n814bar);
  OR2_X1 U152 ( .A1(in[187]), .A2(in[177]), .ZN(n809) );
  AND2_X1 U152bar ( .A1(inbar[187]), .A2(inbar[177]), .ZN(n809bar);
  OR2_X1 U153 ( .A1(in[200]), .A2(in[192]), .ZN(n810) );
  AND2_X1 U153bar ( .A1(inbar[200]), .A2(inbar[192]), .ZN(n810bar);
  OR2_X1 U154 ( .A1(n808), .A2(n807), .ZN(n816) );
  AND2_X1 U154bar ( .A1(n808bar), .A2(n807bar), .ZN(n816bar);
  OR2_X1 U155 ( .A1(n806), .A2(n805), .ZN(n807) );
  AND2_X1 U155bar ( .A1(n806bar), .A2(n805bar), .ZN(n807bar);
  OR2_X1 U156 ( .A1(in[225]), .A2(in[207]), .ZN(n805) );
  AND2_X1 U156bar ( .A1(inbar[225]), .A2(inbar[207]), .ZN(n805bar);
  OR2_X1 U157 ( .A1(in[98]), .A2(in[226]), .ZN(n806) );
  AND2_X1 U157bar ( .A1(inbar[98]), .A2(inbar[226]), .ZN(n806bar);
  OR2_X1 U158 ( .A1(n804), .A2(n803), .ZN(n808) );
  AND2_X1 U158bar ( .A1(n804bar), .A2(n803bar), .ZN(n808bar);
  OR2_X1 U159 ( .A1(in_20), .A2(in_16), .ZN(n803) );
  AND2_X1 U159bar ( .A1(in_20bar), .A2(in_16bar), .ZN(n803bar);
  OR2_X1 U160 ( .A1(in_55), .A2(in_45), .ZN(n804) );
  AND2_X1 U160bar ( .A1(in_55bar), .A2(in_45bar), .ZN(n804bar);
  OR2_X1 U161 ( .A1(n802), .A2(n801), .ZN(n824) );
  AND2_X1 U161bar ( .A1(n802bar), .A2(n801bar), .ZN(n824bar);
  OR2_X1 U162 ( .A1(in[162]), .A2(in[149]), .ZN(n801) );
  AND2_X1 U162bar ( .A1(inbar[162]), .A2(inbar[149]), .ZN(n801bar);
  OR2_X1 U163 ( .A1(in[163]), .A2(n800), .ZN(n802) );
  AND2_X1 U163bar ( .A1(inbar[163]), .A2(n800bar), .ZN(n802bar);
  OR2_X1 U164 ( .A1(in[191]), .A2(in[189]), .ZN(n800) );
  AND2_X1 U164bar ( .A1(inbar[191]), .A2(inbar[189]), .ZN(n800bar);
  OR2_X1 U165 ( .A1(n799), .A2(n798), .ZN(n826) );
  AND2_X1 U165bar ( .A1(n799bar), .A2(n798bar), .ZN(n826bar);
  OR2_X1 U166 ( .A1(n797), .A2(n796), .ZN(n798) );
  AND2_X1 U166bar ( .A1(n797bar), .A2(n796bar), .ZN(n798bar);
  OR2_X1 U167 ( .A1(in[212]), .A2(in[193]), .ZN(n796) );
  AND2_X1 U167bar ( .A1(inbar[212]), .A2(inbar[193]), .ZN(n796bar);
  OR2_X1 U168 ( .A1(in[238]), .A2(n795), .ZN(n797) );
  AND2_X1 U168bar ( .A1(inbar[238]), .A2(n795bar), .ZN(n797bar);
  OR2_X1 U169 ( .A1(in[88]), .A2(in[247]), .ZN(n795) );
  AND2_X1 U169bar ( .A1(inbar[88]), .A2(inbar[247]), .ZN(n795bar);
  OR2_X1 U170 ( .A1(n794), .A2(n793), .ZN(n799) );
  AND2_X1 U170bar ( .A1(n794bar), .A2(n793bar), .ZN(n799bar);
  OR2_X1 U171 ( .A1(in[94]), .A2(in[92]), .ZN(n793) );
  AND2_X1 U171bar ( .A1(inbar[94]), .A2(inbar[92]), .ZN(n793bar);
  OR2_X1 U172 ( .A1(in_52), .A2(n792), .ZN(n794) );
  AND2_X1 U172bar ( .A1(in_52bar), .A2(n792bar), .ZN(n794bar);
  OR2_X1 U173 ( .A1(in_70), .A2(in_67), .ZN(n792) );
  AND2_X1 U173bar ( .A1(in_70bar), .A2(in_67bar), .ZN(n792bar);
  OR2_X1 U174 ( .A1(n791), .A2(n790), .ZN(out[2]) );
  AND2_X1 U174bar ( .A1(n791bar), .A2(n790bar), .ZN(outbar[2]);
  OR2_X1 U175 ( .A1(n789), .A2(n788), .ZN(n790) );
  AND2_X1 U175bar ( .A1(n789bar), .A2(n788bar), .ZN(n790bar);
  OR2_X1 U176 ( .A1(n787), .A2(n786), .ZN(n788) );
  AND2_X1 U176bar ( .A1(n787bar), .A2(n786bar), .ZN(n788bar);
  OR2_X1 U177 ( .A1(n819), .A2(n785), .ZN(n786) );
  AND2_X1 U177bar ( .A1(n819bar), .A2(n785bar), .ZN(n786bar);
  OR2_X1 U178 ( .A1(n784), .A2(n783), .ZN(n819) );
  AND2_X1 U178bar ( .A1(n784bar), .A2(n783bar), .ZN(n819bar);
  OR2_X1 U179 ( .A1(n782), .A2(n781), .ZN(n783) );
  AND2_X1 U179bar ( .A1(n782bar), .A2(n781bar), .ZN(n783bar);
  OR2_X1 U180 ( .A1(n780), .A2(n779), .ZN(n781) );
  AND2_X1 U180bar ( .A1(n780bar), .A2(n779bar), .ZN(n781bar);
  OR2_X1 U181 ( .A1(n962), .A2(n778), .ZN(n779) );
  AND2_X1 U181bar ( .A1(n962bar), .A2(n778bar), .ZN(n779bar);
  OR2_X1 U182 ( .A1(n777), .A2(n776), .ZN(n962) );
  AND2_X1 U182bar ( .A1(n777bar), .A2(n776bar), .ZN(n962bar);
  OR2_X1 U183 ( .A1(n775), .A2(n774), .ZN(n776) );
  AND2_X1 U183bar ( .A1(n775bar), .A2(n774bar), .ZN(n776bar);
  OR2_X1 U184 ( .A1(n773), .A2(n772), .ZN(n774) );
  AND2_X1 U184bar ( .A1(n773bar), .A2(n772bar), .ZN(n774bar);
  OR2_X1 U185 ( .A1(in[131]), .A2(in[120]), .ZN(n772) );
  AND2_X1 U185bar ( .A1(inbar[131]), .A2(inbar[120]), .ZN(n772bar);
  OR2_X1 U186 ( .A1(in[153]), .A2(in[147]), .ZN(n773) );
  AND2_X1 U186bar ( .A1(inbar[153]), .A2(inbar[147]), .ZN(n773bar);
  OR2_X1 U187 ( .A1(n771), .A2(n770), .ZN(n775) );
  AND2_X1 U187bar ( .A1(n771bar), .A2(n770bar), .ZN(n775bar);
  OR2_X1 U188 ( .A1(in[170]), .A2(in[156]), .ZN(n770) );
  AND2_X1 U188bar ( .A1(inbar[170]), .A2(inbar[156]), .ZN(n770bar);
  OR2_X1 U189 ( .A1(in[223]), .A2(in[190]), .ZN(n771) );
  AND2_X1 U189bar ( .A1(inbar[223]), .A2(inbar[190]), .ZN(n771bar);
  OR2_X1 U190 ( .A1(n769), .A2(n768), .ZN(n777) );
  AND2_X1 U190bar ( .A1(n769bar), .A2(n768bar), .ZN(n777bar);
  OR2_X1 U191 ( .A1(n767), .A2(n766), .ZN(n768) );
  AND2_X1 U191bar ( .A1(n767bar), .A2(n766bar), .ZN(n768bar);
  OR2_X1 U192 ( .A1(in[236]), .A2(in[230]), .ZN(n766) );
  AND2_X1 U192bar ( .A1(inbar[236]), .A2(inbar[230]), .ZN(n766bar);
  OR2_X1 U193 ( .A1(in[85]), .A2(in[240]), .ZN(n767) );
  AND2_X1 U193bar ( .A1(inbar[85]), .A2(inbar[240]), .ZN(n767bar);
  OR2_X1 U194 ( .A1(n765), .A2(n764), .ZN(n769) );
  AND2_X1 U194bar ( .A1(n765bar), .A2(n764bar), .ZN(n769bar);
  OR2_X1 U195 ( .A1(in_12), .A2(in[90]), .ZN(n764) );
  AND2_X1 U195bar ( .A1(in_12bar), .A2(inbar[90]), .ZN(n764bar);
  OR2_X1 U196 ( .A1(in_39), .A2(in_28), .ZN(n765) );
  AND2_X1 U196bar ( .A1(in_39bar), .A2(in_28bar), .ZN(n765bar);
  OR2_X1 U197 ( .A1(in[109]), .A2(n763), .ZN(n780) );
  AND2_X1 U197bar ( .A1(inbar[109]), .A2(n763bar), .ZN(n780bar);
  OR2_X1 U198 ( .A1(n762), .A2(n761), .ZN(n782) );
  AND2_X1 U198bar ( .A1(n762bar), .A2(n761bar), .ZN(n782bar);
  OR2_X1 U199 ( .A1(in[138]), .A2(in[129]), .ZN(n761) );
  AND2_X1 U199bar ( .A1(inbar[138]), .A2(inbar[129]), .ZN(n761bar);
  OR2_X1 U200 ( .A1(in[157]), .A2(n760), .ZN(n762) );
  AND2_X1 U200bar ( .A1(inbar[157]), .A2(n760bar), .ZN(n762bar);
  OR2_X1 U201 ( .A1(in[182]), .A2(in[167]), .ZN(n760) );
  AND2_X1 U201bar ( .A1(inbar[182]), .A2(inbar[167]), .ZN(n760bar);
  OR2_X1 U202 ( .A1(n759), .A2(n758), .ZN(n784) );
  AND2_X1 U202bar ( .A1(n759bar), .A2(n758bar), .ZN(n784bar);
  OR2_X1 U203 ( .A1(n757), .A2(n756), .ZN(n758) );
  AND2_X1 U203bar ( .A1(n757bar), .A2(n756bar), .ZN(n758bar);
  OR2_X1 U204 ( .A1(in[195]), .A2(in[184]), .ZN(n756) );
  AND2_X1 U204bar ( .A1(inbar[195]), .A2(inbar[184]), .ZN(n756bar);
  OR2_X1 U205 ( .A1(in[196]), .A2(n755), .ZN(n757) );
  AND2_X1 U205bar ( .A1(inbar[196]), .A2(n755bar), .ZN(n757bar);
  OR2_X1 U206 ( .A1(in[215]), .A2(in[209]), .ZN(n755) );
  AND2_X1 U206bar ( .A1(inbar[215]), .A2(inbar[209]), .ZN(n755bar);
  OR2_X1 U207 ( .A1(n754), .A2(n753), .ZN(n759) );
  AND2_X1 U207bar ( .A1(n754bar), .A2(n753bar), .ZN(n759bar);
  OR2_X1 U208 ( .A1(in[93]), .A2(in[233]), .ZN(n753) );
  AND2_X1 U208bar ( .A1(inbar[93]), .A2(inbar[233]), .ZN(n753bar);
  OR2_X1 U209 ( .A1(in_1), .A2(n752), .ZN(n754) );
  AND2_X1 U209bar ( .A1(in_1bar), .A2(n752bar), .ZN(n754bar);
  OR2_X1 U210 ( .A1(in_69), .A2(in_66), .ZN(n752) );
  AND2_X1 U210bar ( .A1(in_69bar), .A2(in_66bar), .ZN(n752bar);
  OR2_X1 U211 ( .A1(n966), .A2(n751), .ZN(n787) );
  AND2_X1 U211bar ( .A1(n966bar), .A2(n751bar), .ZN(n787bar);
  OR2_X1 U212 ( .A1(in[134]), .A2(n750), .ZN(n751) );
  AND2_X1 U212bar ( .A1(inbar[134]), .A2(n750bar), .ZN(n751bar);
  OR2_X1 U213 ( .A1(n749), .A2(n748), .ZN(n966) );
  AND2_X1 U213bar ( .A1(n749bar), .A2(n748bar), .ZN(n966bar);
  OR2_X1 U214 ( .A1(n747), .A2(n746), .ZN(n748) );
  AND2_X1 U214bar ( .A1(n747bar), .A2(n746bar), .ZN(n748bar);
  OR2_X1 U215 ( .A1(n745), .A2(n744), .ZN(n746) );
  AND2_X1 U215bar ( .A1(n745bar), .A2(n744bar), .ZN(n746bar);
  OR2_X1 U216 ( .A1(in[136]), .A2(in[121]), .ZN(n744) );
  AND2_X1 U216bar ( .A1(inbar[136]), .A2(inbar[121]), .ZN(n744bar);
  OR2_X1 U217 ( .A1(in[186]), .A2(in[174]), .ZN(n745) );
  AND2_X1 U217bar ( .A1(inbar[186]), .A2(inbar[174]), .ZN(n745bar);
  OR2_X1 U218 ( .A1(n743), .A2(n742), .ZN(n747) );
  AND2_X1 U218bar ( .A1(n743bar), .A2(n742bar), .ZN(n747bar);
  OR2_X1 U219 ( .A1(in[198]), .A2(in[197]), .ZN(n742) );
  AND2_X1 U219bar ( .A1(inbar[198]), .A2(inbar[197]), .ZN(n742bar);
  OR2_X1 U220 ( .A1(in[214]), .A2(in[199]), .ZN(n743) );
  AND2_X1 U220bar ( .A1(inbar[214]), .A2(inbar[199]), .ZN(n743bar);
  OR2_X1 U221 ( .A1(n741), .A2(n740), .ZN(n749) );
  AND2_X1 U221bar ( .A1(n741bar), .A2(n740bar), .ZN(n749bar);
  OR2_X1 U222 ( .A1(n739), .A2(n738), .ZN(n740) );
  AND2_X1 U222bar ( .A1(n739bar), .A2(n738bar), .ZN(n740bar);
  OR2_X1 U223 ( .A1(in[231]), .A2(in[220]), .ZN(n738) );
  AND2_X1 U223bar ( .A1(inbar[231]), .A2(inbar[220]), .ZN(n738bar);
  OR2_X1 U224 ( .A1(in_25), .A2(in[245]), .ZN(n739) );
  AND2_X1 U224bar ( .A1(in_25bar), .A2(inbar[245]), .ZN(n739bar);
  OR2_X1 U225 ( .A1(n737), .A2(n736), .ZN(n741) );
  AND2_X1 U225bar ( .A1(n737bar), .A2(n736bar), .ZN(n741bar);
  OR2_X1 U226 ( .A1(in_53), .A2(in_29), .ZN(n736) );
  AND2_X1 U226bar ( .A1(in_53bar), .A2(in_29bar), .ZN(n736bar);
  OR2_X1 U227 ( .A1(in_79), .A2(in_74), .ZN(n737) );
  AND2_X1 U227bar ( .A1(in_79bar), .A2(in_74bar), .ZN(n737bar);
  OR2_X1 U228 ( .A1(n735), .A2(n734), .ZN(n789) );
  AND2_X1 U228bar ( .A1(n735bar), .A2(n734bar), .ZN(n789bar);
  OR2_X1 U229 ( .A1(in[152]), .A2(in[140]), .ZN(n734) );
  AND2_X1 U229bar ( .A1(inbar[152]), .A2(inbar[140]), .ZN(n734bar);
  OR2_X1 U230 ( .A1(in[155]), .A2(n733), .ZN(n735) );
  AND2_X1 U230bar ( .A1(inbar[155]), .A2(n733bar), .ZN(n735bar);
  OR2_X1 U231 ( .A1(in[166]), .A2(in[165]), .ZN(n733) );
  AND2_X1 U231bar ( .A1(inbar[166]), .A2(inbar[165]), .ZN(n733bar);
  OR2_X1 U232 ( .A1(n732), .A2(n731), .ZN(n791) );
  AND2_X1 U232bar ( .A1(n732bar), .A2(n731bar), .ZN(n791bar);
  OR2_X1 U233 ( .A1(n730), .A2(n729), .ZN(n731) );
  AND2_X1 U233bar ( .A1(n730bar), .A2(n729bar), .ZN(n731bar);
  OR2_X1 U234 ( .A1(in[202]), .A2(in[185]), .ZN(n729) );
  AND2_X1 U234bar ( .A1(inbar[202]), .A2(inbar[185]), .ZN(n729bar);
  OR2_X1 U235 ( .A1(in[211]), .A2(n728), .ZN(n730) );
  AND2_X1 U235bar ( .A1(inbar[211]), .A2(n728bar), .ZN(n730bar);
  OR2_X1 U236 ( .A1(in[255]), .A2(in[253]), .ZN(n728) );
  AND2_X1 U236bar ( .A1(inbar[255]), .A2(inbar[253]), .ZN(n728bar);
  OR2_X1 U237 ( .A1(n727), .A2(n726), .ZN(n732) );
  AND2_X1 U237bar ( .A1(n727bar), .A2(n726bar), .ZN(n732bar);
  OR2_X1 U238 ( .A1(in_35), .A2(in_15), .ZN(n726) );
  AND2_X1 U238bar ( .A1(in_35bar), .A2(in_15bar), .ZN(n726bar);
  OR2_X1 U239 ( .A1(in_36), .A2(n725), .ZN(n727) );
  AND2_X1 U239bar ( .A1(in_36bar), .A2(n725bar), .ZN(n727bar);
  OR2_X1 U240 ( .A1(in_48), .A2(in_40), .ZN(n725) );
  AND2_X1 U240bar ( .A1(in_48bar), .A2(in_40bar), .ZN(n725bar);
  OR2_X1 U241 ( .A1(n724), .A2(n723), .ZN(out[1]) );
  AND2_X1 U241bar ( .A1(n724bar), .A2(n723bar), .ZN(outbar[1]);
  OR2_X1 U242 ( .A1(n722), .A2(n721), .ZN(n723) );
  AND2_X1 U242bar ( .A1(n722bar), .A2(n721bar), .ZN(n723bar);
  OR2_X1 U243 ( .A1(n720), .A2(n719), .ZN(n721) );
  AND2_X1 U243bar ( .A1(n720bar), .A2(n719bar), .ZN(n721bar);
  OR2_X1 U244 ( .A1(n921), .A2(n887), .ZN(n719) );
  AND2_X1 U244bar ( .A1(n921bar), .A2(n887bar), .ZN(n719bar);
  OR2_X1 U245 ( .A1(n718), .A2(n717), .ZN(n887) );
  AND2_X1 U245bar ( .A1(n718bar), .A2(n717bar), .ZN(n887bar);
  OR2_X1 U246 ( .A1(n716), .A2(n715), .ZN(n717) );
  AND2_X1 U246bar ( .A1(n716bar), .A2(n715bar), .ZN(n717bar);
  OR2_X1 U247 ( .A1(n714), .A2(n713), .ZN(n715) );
  AND2_X1 U247bar ( .A1(n714bar), .A2(n713bar), .ZN(n715bar);
  OR2_X1 U248 ( .A1(in[116]), .A2(in[110]), .ZN(n713) );
  AND2_X1 U248bar ( .A1(inbar[116]), .A2(inbar[110]), .ZN(n713bar);
  OR2_X1 U249 ( .A1(in[133]), .A2(in[130]), .ZN(n714) );
  AND2_X1 U249bar ( .A1(inbar[133]), .A2(inbar[130]), .ZN(n714bar);
  OR2_X1 U250 ( .A1(n712), .A2(n711), .ZN(n716) );
  AND2_X1 U250bar ( .A1(n712bar), .A2(n711bar), .ZN(n716bar);
  OR2_X1 U251 ( .A1(in[203]), .A2(in[135]), .ZN(n711) );
  AND2_X1 U251bar ( .A1(inbar[203]), .A2(inbar[135]), .ZN(n711bar);
  OR2_X1 U252 ( .A1(in[232]), .A2(in[223]), .ZN(n712) );
  AND2_X1 U252bar ( .A1(inbar[232]), .A2(inbar[223]), .ZN(n712bar);
  OR2_X1 U253 ( .A1(n710), .A2(n709), .ZN(n718) );
  AND2_X1 U253bar ( .A1(n710bar), .A2(n709bar), .ZN(n718bar);
  OR2_X1 U254 ( .A1(n708), .A2(n707), .ZN(n709) );
  AND2_X1 U254bar ( .A1(n708bar), .A2(n707bar), .ZN(n709bar);
  OR2_X1 U255 ( .A1(in[255]), .A2(in[233]), .ZN(n707) );
  AND2_X1 U255bar ( .A1(inbar[255]), .A2(inbar[233]), .ZN(n707bar);
  OR2_X1 U256 ( .A1(in_53), .A2(in_34), .ZN(n708) );
  AND2_X1 U256bar ( .A1(in_53bar), .A2(in_34bar), .ZN(n708bar);
  OR2_X1 U257 ( .A1(n706), .A2(n705), .ZN(n710) );
  AND2_X1 U257bar ( .A1(n706bar), .A2(n705bar), .ZN(n710bar);
  OR2_X1 U258 ( .A1(in_57), .A2(in_55), .ZN(n705) );
  AND2_X1 U258bar ( .A1(in_57bar), .A2(in_55bar), .ZN(n705bar);
  OR2_X1 U259 ( .A1(in_68), .A2(in_67), .ZN(n706) );
  AND2_X1 U259bar ( .A1(in_68bar), .A2(in_67bar), .ZN(n706bar);
  OR2_X1 U260 ( .A1(n704), .A2(n703), .ZN(n921) );
  AND2_X1 U260bar ( .A1(n704bar), .A2(n703bar), .ZN(n921bar);
  OR2_X1 U261 ( .A1(n702), .A2(n701), .ZN(n703) );
  AND2_X1 U261bar ( .A1(n702bar), .A2(n701bar), .ZN(n703bar);
  OR2_X1 U262 ( .A1(n700), .A2(n699), .ZN(n701) );
  AND2_X1 U262bar ( .A1(n700bar), .A2(n699bar), .ZN(n701bar);
  OR2_X1 U263 ( .A1(n944), .A2(n872), .ZN(n699) );
  AND2_X1 U263bar ( .A1(n944bar), .A2(n872bar), .ZN(n699bar);
  OR2_X1 U264 ( .A1(n698), .A2(n697), .ZN(n872) );
  AND2_X1 U264bar ( .A1(n698bar), .A2(n697bar), .ZN(n872bar);
  OR2_X1 U265 ( .A1(n696), .A2(n695), .ZN(n697) );
  AND2_X1 U265bar ( .A1(n696bar), .A2(n695bar), .ZN(n697bar);
  OR2_X1 U266 ( .A1(n694), .A2(n693), .ZN(n695) );
  AND2_X1 U266bar ( .A1(n694bar), .A2(n693bar), .ZN(n695bar);
  OR2_X1 U267 ( .A1(in[121]), .A2(in[102]), .ZN(n693) );
  AND2_X1 U267bar ( .A1(inbar[121]), .A2(inbar[102]), .ZN(n693bar);
  OR2_X1 U268 ( .A1(in[162]), .A2(in[161]), .ZN(n694) );
  AND2_X1 U268bar ( .A1(inbar[162]), .A2(inbar[161]), .ZN(n694bar);
  OR2_X1 U269 ( .A1(n692), .A2(n691), .ZN(n696) );
  AND2_X1 U269bar ( .A1(n692bar), .A2(n691bar), .ZN(n696bar);
  OR2_X1 U270 ( .A1(in[192]), .A2(in[178]), .ZN(n691) );
  AND2_X1 U270bar ( .A1(inbar[192]), .A2(inbar[178]), .ZN(n691bar);
  OR2_X1 U271 ( .A1(in[244]), .A2(in[209]), .ZN(n692) );
  AND2_X1 U271bar ( .A1(inbar[244]), .A2(inbar[209]), .ZN(n692bar);
  OR2_X1 U272 ( .A1(n690), .A2(n689), .ZN(n698) );
  AND2_X1 U272bar ( .A1(n690bar), .A2(n689bar), .ZN(n698bar);
  OR2_X1 U273 ( .A1(n688), .A2(n687), .ZN(n689) );
  AND2_X1 U273bar ( .A1(n688bar), .A2(n687bar), .ZN(n689bar);
  OR2_X1 U274 ( .A1(in[90]), .A2(in[254]), .ZN(n687) );
  AND2_X1 U274bar ( .A1(inbar[90]), .A2(inbar[254]), .ZN(n687bar);
  OR2_X1 U275 ( .A1(in_36), .A2(in_32), .ZN(n688) );
  AND2_X1 U275bar ( .A1(in_36bar), .A2(in_32bar), .ZN(n688bar);
  OR2_X1 U276 ( .A1(n686), .A2(n685), .ZN(n690) );
  AND2_X1 U276bar ( .A1(n686bar), .A2(n685bar), .ZN(n690bar);
  OR2_X1 U277 ( .A1(in_62), .A2(in_37), .ZN(n685) );
  AND2_X1 U277bar ( .A1(in_62bar), .A2(in_37bar), .ZN(n685bar);
  OR2_X1 U278 ( .A1(in_75), .A2(in_73), .ZN(n686) );
  AND2_X1 U278bar ( .A1(in_75bar), .A2(in_73bar), .ZN(n686bar);
  OR2_X1 U279 ( .A1(n684), .A2(n683), .ZN(n944) );
  AND2_X1 U279bar ( .A1(n684bar), .A2(n683bar), .ZN(n944bar);
  OR2_X1 U280 ( .A1(n682), .A2(n681), .ZN(n683) );
  AND2_X1 U280bar ( .A1(n682bar), .A2(n681bar), .ZN(n683bar);
  OR2_X1 U281 ( .A1(n680), .A2(n679), .ZN(n681) );
  AND2_X1 U281bar ( .A1(n680bar), .A2(n679bar), .ZN(n681bar);
  OR2_X1 U282 ( .A1(in[171]), .A2(in[153]), .ZN(n679) );
  AND2_X1 U282bar ( .A1(inbar[171]), .A2(inbar[153]), .ZN(n679bar);
  OR2_X1 U283 ( .A1(in[187]), .A2(in[176]), .ZN(n680) );
  AND2_X1 U283bar ( .A1(inbar[187]), .A2(inbar[176]), .ZN(n680bar);
  OR2_X1 U284 ( .A1(n678), .A2(n677), .ZN(n682) );
  AND2_X1 U284bar ( .A1(n678bar), .A2(n677bar), .ZN(n682bar);
  OR2_X1 U285 ( .A1(in[245]), .A2(in[211]), .ZN(n677) );
  AND2_X1 U285bar ( .A1(inbar[245]), .A2(inbar[211]), .ZN(n677bar);
  OR2_X1 U286 ( .A1(in[97]), .A2(in[88]), .ZN(n678) );
  AND2_X1 U286bar ( .A1(inbar[97]), .A2(inbar[88]), .ZN(n678bar);
  OR2_X1 U287 ( .A1(n676), .A2(n675), .ZN(n684) );
  AND2_X1 U287bar ( .A1(n676bar), .A2(n675bar), .ZN(n684bar);
  OR2_X1 U288 ( .A1(n674), .A2(n673), .ZN(n675) );
  AND2_X1 U288bar ( .A1(n674bar), .A2(n673bar), .ZN(n675bar);
  OR2_X1 U289 ( .A1(in_10), .A2(in_0), .ZN(n673) );
  AND2_X1 U289bar ( .A1(in_10bar), .A2(in_0bar), .ZN(n673bar);
  OR2_X1 U290 ( .A1(in_59), .A2(in_5), .ZN(n674) );
  AND2_X1 U290bar ( .A1(in_59bar), .A2(in_5bar), .ZN(n674bar);
  OR2_X1 U291 ( .A1(n672), .A2(n671), .ZN(n676) );
  AND2_X1 U291bar ( .A1(n672bar), .A2(n671bar), .ZN(n676bar);
  OR2_X1 U292 ( .A1(in_60), .A2(in_6), .ZN(n671) );
  AND2_X1 U292bar ( .A1(in_60bar), .A2(in_6bar), .ZN(n671bar);
  OR2_X1 U293 ( .A1(in_77), .A2(in_69), .ZN(n672) );
  AND2_X1 U293bar ( .A1(in_77bar), .A2(in_69bar), .ZN(n672bar);
  OR2_X1 U294 ( .A1(in[113]), .A2(n864), .ZN(n700) );
  AND2_X1 U294bar ( .A1(inbar[113]), .A2(n864bar), .ZN(n700bar);
  OR2_X1 U295 ( .A1(n670), .A2(n669), .ZN(n864) );
  AND2_X1 U295bar ( .A1(n670bar), .A2(n669bar), .ZN(n864bar);
  OR2_X1 U296 ( .A1(n668), .A2(n667), .ZN(n669) );
  AND2_X1 U296bar ( .A1(n668bar), .A2(n667bar), .ZN(n669bar);
  OR2_X1 U297 ( .A1(n666), .A2(n665), .ZN(n667) );
  AND2_X1 U297bar ( .A1(n666bar), .A2(n665bar), .ZN(n667bar);
  OR2_X1 U298 ( .A1(in[125]), .A2(in[107]), .ZN(n665) );
  AND2_X1 U298bar ( .A1(inbar[125]), .A2(inbar[107]), .ZN(n665bar);
  OR2_X1 U299 ( .A1(in[138]), .A2(in[126]), .ZN(n666) );
  AND2_X1 U299bar ( .A1(inbar[138]), .A2(inbar[126]), .ZN(n666bar);
  OR2_X1 U300 ( .A1(n664), .A2(n663), .ZN(n668) );
  AND2_X1 U300bar ( .A1(n664bar), .A2(n663bar), .ZN(n668bar);
  OR2_X1 U301 ( .A1(in[189]), .A2(in[143]), .ZN(n663) );
  AND2_X1 U301bar ( .A1(inbar[189]), .A2(inbar[143]), .ZN(n663bar);
  OR2_X1 U302 ( .A1(in[99]), .A2(in[214]), .ZN(n664) );
  AND2_X1 U302bar ( .A1(inbar[99]), .A2(inbar[214]), .ZN(n664bar);
  OR2_X1 U303 ( .A1(n662), .A2(n661), .ZN(n670) );
  AND2_X1 U303bar ( .A1(n662bar), .A2(n661bar), .ZN(n670bar);
  OR2_X1 U304 ( .A1(n660), .A2(n659), .ZN(n661) );
  AND2_X1 U304bar ( .A1(n660bar), .A2(n659bar), .ZN(n661bar);
  OR2_X1 U305 ( .A1(in_15), .A2(in_12), .ZN(n659) );
  AND2_X1 U305bar ( .A1(in_15bar), .A2(in_12bar), .ZN(n659bar);
  OR2_X1 U306 ( .A1(in_20), .A2(in_2), .ZN(n660) );
  AND2_X1 U306bar ( .A1(in_20bar), .A2(in_2bar), .ZN(n660bar);
  OR2_X1 U307 ( .A1(n658), .A2(n657), .ZN(n662) );
  AND2_X1 U307bar ( .A1(n658bar), .A2(n657bar), .ZN(n662bar);
  OR2_X1 U308 ( .A1(in_30), .A2(in_3), .ZN(n657) );
  AND2_X1 U308bar ( .A1(in_30bar), .A2(in_3bar), .ZN(n657bar);
  OR2_X1 U309 ( .A1(in_4), .A2(in_38), .ZN(n658) );
  AND2_X1 U309bar ( .A1(in_4bar), .A2(in_38bar), .ZN(n658bar);
  OR2_X1 U310 ( .A1(n656), .A2(n655), .ZN(n702) );
  AND2_X1 U310bar ( .A1(n656bar), .A2(n655bar), .ZN(n702bar);
  OR2_X1 U311 ( .A1(in[148]), .A2(in[137]), .ZN(n655) );
  AND2_X1 U311bar ( .A1(inbar[148]), .A2(inbar[137]), .ZN(n655bar);
  OR2_X1 U312 ( .A1(in[149]), .A2(n654), .ZN(n656) );
  AND2_X1 U312bar ( .A1(inbar[149]), .A2(n654bar), .ZN(n656bar);
  OR2_X1 U313 ( .A1(in[195]), .A2(in[190]), .ZN(n654) );
  AND2_X1 U313bar ( .A1(inbar[195]), .A2(inbar[190]), .ZN(n654bar);
  OR2_X1 U314 ( .A1(n653), .A2(n652), .ZN(n704) );
  AND2_X1 U314bar ( .A1(n653bar), .A2(n652bar), .ZN(n704bar);
  OR2_X1 U315 ( .A1(n651), .A2(n650), .ZN(n652) );
  AND2_X1 U315bar ( .A1(n651bar), .A2(n650bar), .ZN(n652bar);
  OR2_X1 U316 ( .A1(in[98]), .A2(in[197]), .ZN(n650) );
  AND2_X1 U316bar ( .A1(inbar[98]), .A2(inbar[197]), .ZN(n650bar);
  OR2_X1 U317 ( .A1(in_11), .A2(n649), .ZN(n651) );
  AND2_X1 U317bar ( .A1(in_11bar), .A2(n649bar), .ZN(n651bar);
  OR2_X1 U318 ( .A1(in_26), .A2(in_14), .ZN(n649) );
  AND2_X1 U318bar ( .A1(in_26bar), .A2(in_14bar), .ZN(n649bar);
  OR2_X1 U319 ( .A1(n648), .A2(n647), .ZN(n653) );
  AND2_X1 U319bar ( .A1(n648bar), .A2(n647bar), .ZN(n653bar);
  OR2_X1 U320 ( .A1(in_35), .A2(in_27), .ZN(n647) );
  AND2_X1 U320bar ( .A1(in_35bar), .A2(in_27bar), .ZN(n647bar);
  OR2_X1 U321 ( .A1(in_50), .A2(n646), .ZN(n648) );
  AND2_X1 U321bar ( .A1(in_50bar), .A2(n646bar), .ZN(n648bar);
  OR2_X1 U322 ( .A1(in_78), .A2(in_61), .ZN(n646) );
  AND2_X1 U322bar ( .A1(in_78bar), .A2(in_61bar), .ZN(n646bar);
  OR2_X1 U323 ( .A1(n942), .A2(n645), .ZN(n720) );
  AND2_X1 U323bar ( .A1(n942bar), .A2(n645bar), .ZN(n720bar);
  OR2_X1 U324 ( .A1(in[106]), .A2(n863), .ZN(n645) );
  AND2_X1 U324bar ( .A1(inbar[106]), .A2(n863bar), .ZN(n645bar);
  OR2_X1 U325 ( .A1(n644), .A2(n643), .ZN(n863) );
  AND2_X1 U325bar ( .A1(n644bar), .A2(n643bar), .ZN(n863bar);
  OR2_X1 U326 ( .A1(n642), .A2(n641), .ZN(n643) );
  AND2_X1 U326bar ( .A1(n642bar), .A2(n641bar), .ZN(n643bar);
  OR2_X1 U327 ( .A1(n640), .A2(n639), .ZN(n641) );
  AND2_X1 U327bar ( .A1(n640bar), .A2(n639bar), .ZN(n641bar);
  OR2_X1 U328 ( .A1(in[127]), .A2(in[122]), .ZN(n639) );
  AND2_X1 U328bar ( .A1(inbar[127]), .A2(inbar[122]), .ZN(n639bar);
  OR2_X1 U329 ( .A1(in[156]), .A2(in[132]), .ZN(n640) );
  AND2_X1 U329bar ( .A1(inbar[156]), .A2(inbar[132]), .ZN(n640bar);
  OR2_X1 U330 ( .A1(n638), .A2(n637), .ZN(n642) );
  AND2_X1 U330bar ( .A1(n638bar), .A2(n637bar), .ZN(n642bar);
  OR2_X1 U331 ( .A1(in[159]), .A2(in[157]), .ZN(n637) );
  AND2_X1 U331bar ( .A1(inbar[159]), .A2(inbar[157]), .ZN(n637bar);
  OR2_X1 U332 ( .A1(in[185]), .A2(in[169]), .ZN(n638) );
  AND2_X1 U332bar ( .A1(inbar[185]), .A2(inbar[169]), .ZN(n638bar);
  OR2_X1 U333 ( .A1(n636), .A2(n635), .ZN(n644) );
  AND2_X1 U333bar ( .A1(n636bar), .A2(n635bar), .ZN(n644bar);
  OR2_X1 U334 ( .A1(n634), .A2(n633), .ZN(n635) );
  AND2_X1 U334bar ( .A1(n634bar), .A2(n633bar), .ZN(n635bar);
  OR2_X1 U335 ( .A1(in[239]), .A2(in[218]), .ZN(n633) );
  AND2_X1 U335bar ( .A1(inbar[239]), .A2(inbar[218]), .ZN(n633bar);
  OR2_X1 U336 ( .A1(in_13), .A2(in[87]), .ZN(n634) );
  AND2_X1 U336bar ( .A1(in_13bar), .A2(inbar[87]), .ZN(n634bar);
  OR2_X1 U337 ( .A1(n632), .A2(n631), .ZN(n636) );
  AND2_X1 U337bar ( .A1(n632bar), .A2(n631bar), .ZN(n636bar);
  OR2_X1 U338 ( .A1(in_72), .A2(in_70), .ZN(n631) );
  AND2_X1 U338bar ( .A1(in_72bar), .A2(in_70bar), .ZN(n631bar);
  OR2_X1 U339 ( .A1(in_80), .A2(in_74), .ZN(n632) );
  AND2_X1 U339bar ( .A1(in_80bar), .A2(in_74bar), .ZN(n632bar);
  OR2_X1 U340 ( .A1(n630), .A2(n629), .ZN(n942) );
  AND2_X1 U340bar ( .A1(n630bar), .A2(n629bar), .ZN(n942bar);
  OR2_X1 U341 ( .A1(n628), .A2(n627), .ZN(n629) );
  AND2_X1 U341bar ( .A1(n628bar), .A2(n627bar), .ZN(n629bar);
  OR2_X1 U342 ( .A1(n626), .A2(n625), .ZN(n627) );
  AND2_X1 U342bar ( .A1(n626bar), .A2(n625bar), .ZN(n627bar);
  OR2_X1 U343 ( .A1(in[146]), .A2(in[100]), .ZN(n625) );
  AND2_X1 U343bar ( .A1(inbar[146]), .A2(inbar[100]), .ZN(n625bar);
  OR2_X1 U344 ( .A1(in[168]), .A2(in[152]), .ZN(n626) );
  AND2_X1 U344bar ( .A1(inbar[168]), .A2(inbar[152]), .ZN(n626bar);
  OR2_X1 U345 ( .A1(n624), .A2(n623), .ZN(n628) );
  AND2_X1 U345bar ( .A1(n624bar), .A2(n623bar), .ZN(n628bar);
  OR2_X1 U346 ( .A1(in[199]), .A2(in[182]), .ZN(n623) );
  AND2_X1 U346bar ( .A1(inbar[199]), .A2(inbar[182]), .ZN(n623bar);
  OR2_X1 U347 ( .A1(in[236]), .A2(in[204]), .ZN(n624) );
  AND2_X1 U347bar ( .A1(inbar[236]), .A2(inbar[204]), .ZN(n624bar);
  OR2_X1 U348 ( .A1(n622), .A2(n621), .ZN(n630) );
  AND2_X1 U348bar ( .A1(n622bar), .A2(n621bar), .ZN(n630bar);
  OR2_X1 U349 ( .A1(n620), .A2(n619), .ZN(n621) );
  AND2_X1 U349bar ( .A1(n620bar), .A2(n619bar), .ZN(n621bar);
  OR2_X1 U350 ( .A1(in[89]), .A2(in[246]), .ZN(n619) );
  AND2_X1 U350bar ( .A1(inbar[89]), .A2(inbar[246]), .ZN(n619bar);
  OR2_X1 U351 ( .A1(in[95]), .A2(in[92]), .ZN(n620) );
  AND2_X1 U351bar ( .A1(inbar[95]), .A2(inbar[92]), .ZN(n620bar);
  OR2_X1 U352 ( .A1(n618), .A2(n617), .ZN(n622) );
  AND2_X1 U352bar ( .A1(n618bar), .A2(n617bar), .ZN(n622bar);
  OR2_X1 U353 ( .A1(in_22), .A2(in_16), .ZN(n617) );
  AND2_X1 U353bar ( .A1(in_22bar), .A2(in_16bar), .ZN(n617bar);
  OR2_X1 U354 ( .A1(in_51), .A2(in_49), .ZN(n618) );
  AND2_X1 U354bar ( .A1(in_51bar), .A2(in_49bar), .ZN(n618bar);
  OR2_X1 U355 ( .A1(n616), .A2(n615), .ZN(n722) );
  AND2_X1 U355bar ( .A1(n616bar), .A2(n615bar), .ZN(n722bar);
  OR2_X1 U356 ( .A1(in[158]), .A2(in[115]), .ZN(n615) );
  AND2_X1 U356bar ( .A1(inbar[158]), .A2(inbar[115]), .ZN(n615bar);
  OR2_X1 U357 ( .A1(in[163]), .A2(n614), .ZN(n616) );
  AND2_X1 U357bar ( .A1(inbar[163]), .A2(n614bar), .ZN(n616bar);
  OR2_X1 U358 ( .A1(in[206]), .A2(in[165]), .ZN(n614) );
  AND2_X1 U358bar ( .A1(inbar[206]), .A2(inbar[165]), .ZN(n614bar);
  OR2_X1 U359 ( .A1(n613), .A2(n612), .ZN(n724) );
  AND2_X1 U359bar ( .A1(n613bar), .A2(n612bar), .ZN(n724bar);
  OR2_X1 U360 ( .A1(n611), .A2(n610), .ZN(n612) );
  AND2_X1 U360bar ( .A1(n611bar), .A2(n610bar), .ZN(n612bar);
  OR2_X1 U361 ( .A1(in[213]), .A2(in[207]), .ZN(n610) );
  AND2_X1 U361bar ( .A1(inbar[213]), .A2(inbar[207]), .ZN(n610bar);
  OR2_X1 U362 ( .A1(in[215]), .A2(n609), .ZN(n611) );
  AND2_X1 U362bar ( .A1(inbar[215]), .A2(n609bar), .ZN(n611bar);
  OR2_X1 U363 ( .A1(in[230]), .A2(in[220]), .ZN(n609) );
  AND2_X1 U363bar ( .A1(inbar[230]), .A2(inbar[220]), .ZN(n609bar);
  OR2_X1 U364 ( .A1(n608), .A2(n607), .ZN(n613) );
  AND2_X1 U364bar ( .A1(n608bar), .A2(n607bar), .ZN(n613bar);
  OR2_X1 U365 ( .A1(in[251]), .A2(in[234]), .ZN(n607) );
  AND2_X1 U365bar ( .A1(inbar[251]), .A2(inbar[234]), .ZN(n607bar);
  OR2_X1 U366 ( .A1(in_17), .A2(n606), .ZN(n608) );
  AND2_X1 U366bar ( .A1(in_17bar), .A2(n606bar), .ZN(n608bar);
  OR2_X1 U367 ( .A1(in_65), .A2(in_56), .ZN(n606) );
  AND2_X1 U367bar ( .A1(in_65bar), .A2(in_56bar), .ZN(n606bar);
  OR2_X1 U368 ( .A1(n605), .A2(n604), .ZN(out[0]) );
  AND2_X1 U368bar ( .A1(n605bar), .A2(n604bar), .ZN(outbar[0]);
  OR2_X1 U369 ( .A1(n603), .A2(n602), .ZN(n604) );
  AND2_X1 U369bar ( .A1(n603bar), .A2(n602bar), .ZN(n604bar);
  OR2_X1 U370 ( .A1(n601), .A2(n600), .ZN(n602) );
  AND2_X1 U370bar ( .A1(n601bar), .A2(n600bar), .ZN(n602bar);
  OR2_X1 U371 ( .A1(n820), .A2(n785), .ZN(n600) );
  AND2_X1 U371bar ( .A1(n820bar), .A2(n785bar), .ZN(n600bar);
  OR2_X1 U372 ( .A1(n599), .A2(n598), .ZN(n785) );
  AND2_X1 U372bar ( .A1(n599bar), .A2(n598bar), .ZN(n785bar);
  OR2_X1 U373 ( .A1(n597), .A2(n596), .ZN(n598) );
  AND2_X1 U373bar ( .A1(n597bar), .A2(n596bar), .ZN(n598bar);
  OR2_X1 U374 ( .A1(n595), .A2(n594), .ZN(n596) );
  AND2_X1 U374bar ( .A1(n595bar), .A2(n594bar), .ZN(n596bar);
  OR2_X1 U375 ( .A1(in[135]), .A2(in[104]), .ZN(n594) );
  AND2_X1 U375bar ( .A1(inbar[135]), .A2(inbar[104]), .ZN(n594bar);
  OR2_X1 U376 ( .A1(in[188]), .A2(in[178]), .ZN(n595) );
  AND2_X1 U376bar ( .A1(inbar[188]), .A2(inbar[178]), .ZN(n595bar);
  OR2_X1 U377 ( .A1(n593), .A2(n592), .ZN(n597) );
  AND2_X1 U377bar ( .A1(n593bar), .A2(n592bar), .ZN(n597bar);
  OR2_X1 U378 ( .A1(in[217]), .A2(in[194]), .ZN(n592) );
  AND2_X1 U378bar ( .A1(inbar[217]), .A2(inbar[194]), .ZN(n592bar);
  OR2_X1 U379 ( .A1(in[237]), .A2(in[218]), .ZN(n593) );
  AND2_X1 U379bar ( .A1(inbar[237]), .A2(inbar[218]), .ZN(n593bar);
  OR2_X1 U380 ( .A1(n591), .A2(n590), .ZN(n599) );
  AND2_X1 U380bar ( .A1(n591bar), .A2(n590bar), .ZN(n599bar);
  OR2_X1 U381 ( .A1(n589), .A2(n588), .ZN(n590) );
  AND2_X1 U381bar ( .A1(n589bar), .A2(n588bar), .ZN(n590bar);
  OR2_X1 U382 ( .A1(in_2), .A2(in_10), .ZN(n588) );
  AND2_X1 U382bar ( .A1(in_2bar), .A2(in_10bar), .ZN(n588bar);
  OR2_X1 U383 ( .A1(in_47), .A2(in_22), .ZN(n589) );
  AND2_X1 U383bar ( .A1(in_47bar), .A2(in_22bar), .ZN(n589bar);
  OR2_X1 U384 ( .A1(n587), .A2(n586), .ZN(n591) );
  AND2_X1 U384bar ( .A1(n587bar), .A2(n586bar), .ZN(n591bar);
  OR2_X1 U385 ( .A1(in_56), .A2(in_54), .ZN(n586) );
  AND2_X1 U385bar ( .A1(in_56bar), .A2(in_54bar), .ZN(n586bar);
  OR2_X1 U386 ( .A1(in_63), .A2(in_61), .ZN(n587) );
  AND2_X1 U386bar ( .A1(in_63bar), .A2(in_61bar), .ZN(n587bar);
  OR2_X1 U387 ( .A1(n585), .A2(n584), .ZN(n820) );
  AND2_X1 U387bar ( .A1(n585bar), .A2(n584bar), .ZN(n820bar);
  OR2_X1 U388 ( .A1(n583), .A2(n582), .ZN(n584) );
  AND2_X1 U388bar ( .A1(n583bar), .A2(n582bar), .ZN(n584bar);
  OR2_X1 U389 ( .A1(n581), .A2(n580), .ZN(n582) );
  AND2_X1 U389bar ( .A1(n581bar), .A2(n580bar), .ZN(n582bar);
  OR2_X1 U390 ( .A1(in[158]), .A2(in[142]), .ZN(n580) );
  AND2_X1 U390bar ( .A1(inbar[158]), .A2(inbar[142]), .ZN(n580bar);
  OR2_X1 U391 ( .A1(in[175]), .A2(in[164]), .ZN(n581) );
  AND2_X1 U391bar ( .A1(inbar[175]), .A2(inbar[164]), .ZN(n581bar);
  OR2_X1 U392 ( .A1(n579), .A2(n578), .ZN(n583) );
  AND2_X1 U392bar ( .A1(n579bar), .A2(n578bar), .ZN(n583bar);
  OR2_X1 U393 ( .A1(in[228]), .A2(in[204]), .ZN(n578) );
  AND2_X1 U393bar ( .A1(inbar[228]), .A2(inbar[204]), .ZN(n578bar);
  OR2_X1 U394 ( .A1(in[91]), .A2(in[87]), .ZN(n579) );
  AND2_X1 U394bar ( .A1(inbar[91]), .A2(inbar[87]), .ZN(n579bar);
  OR2_X1 U395 ( .A1(n577), .A2(n576), .ZN(n585) );
  AND2_X1 U395bar ( .A1(n577bar), .A2(n576bar), .ZN(n585bar);
  OR2_X1 U396 ( .A1(n575), .A2(n574), .ZN(n576) );
  AND2_X1 U396bar ( .A1(n575bar), .A2(n574bar), .ZN(n576bar);
  OR2_X1 U397 ( .A1(in_21), .A2(in_11), .ZN(n574) );
  AND2_X1 U397bar ( .A1(in_21bar), .A2(in_11bar), .ZN(n574bar);
  OR2_X1 U398 ( .A1(in_5), .A2(in_3), .ZN(n575) );
  AND2_X1 U398bar ( .A1(in_5bar), .A2(in_3bar), .ZN(n575bar);
  OR2_X1 U399 ( .A1(n573), .A2(n572), .ZN(n577) );
  AND2_X1 U399bar ( .A1(n573bar), .A2(n572bar), .ZN(n577bar);
  OR2_X1 U400 ( .A1(in_68), .A2(in_64), .ZN(n572) );
  AND2_X1 U400bar ( .A1(in_68bar), .A2(in_64bar), .ZN(n572bar);
  OR2_X1 U401 ( .A1(in_76), .A2(in_73), .ZN(n573) );
  AND2_X1 U401bar ( .A1(in_76bar), .A2(in_73bar), .ZN(n573bar);
  OR2_X1 U402 ( .A1(n778), .A2(n571), .ZN(n601) );
  AND2_X1 U402bar ( .A1(n778bar), .A2(n571bar), .ZN(n601bar);
  OR2_X1 U403 ( .A1(in[100]), .A2(n965), .ZN(n571) );
  AND2_X1 U403bar ( .A1(inbar[100]), .A2(n965bar), .ZN(n571bar);
  OR2_X1 U404 ( .A1(n570), .A2(n569), .ZN(n965) );
  AND2_X1 U404bar ( .A1(n570bar), .A2(n569bar), .ZN(n965bar);
  OR2_X1 U405 ( .A1(n568), .A2(n567), .ZN(n569) );
  AND2_X1 U405bar ( .A1(n568bar), .A2(n567bar), .ZN(n569bar);
  OR2_X1 U406 ( .A1(n566), .A2(n565), .ZN(n567) );
  AND2_X1 U406bar ( .A1(n566bar), .A2(n565bar), .ZN(n567bar);
  OR2_X1 U407 ( .A1(n817), .A2(n750), .ZN(n565) );
  AND2_X1 U407bar ( .A1(n817bar), .A2(n750bar), .ZN(n565bar);
  OR2_X1 U408 ( .A1(n564), .A2(n563), .ZN(n750) );
  AND2_X1 U408bar ( .A1(n564bar), .A2(n563bar), .ZN(n750bar);
  OR2_X1 U409 ( .A1(n562), .A2(n561), .ZN(n563) );
  AND2_X1 U409bar ( .A1(n562bar), .A2(n561bar), .ZN(n563bar);
  OR2_X1 U410 ( .A1(n560), .A2(n559), .ZN(n561) );
  AND2_X1 U410bar ( .A1(n560bar), .A2(n559bar), .ZN(n561bar);
  OR2_X1 U411 ( .A1(in[119]), .A2(in[103]), .ZN(n559) );
  AND2_X1 U411bar ( .A1(inbar[119]), .A2(inbar[103]), .ZN(n559bar);
  OR2_X1 U412 ( .A1(in[137]), .A2(in[133]), .ZN(n560) );
  AND2_X1 U412bar ( .A1(inbar[137]), .A2(inbar[133]), .ZN(n560bar);
  OR2_X1 U413 ( .A1(n558), .A2(n557), .ZN(n562) );
  AND2_X1 U413bar ( .A1(n558bar), .A2(n557bar), .ZN(n562bar);
  OR2_X1 U414 ( .A1(in[176]), .A2(in[173]), .ZN(n557) );
  AND2_X1 U414bar ( .A1(inbar[176]), .A2(inbar[173]), .ZN(n557bar);
  OR2_X1 U415 ( .A1(in[210]), .A2(in[181]), .ZN(n558) );
  AND2_X1 U415bar ( .A1(inbar[210]), .A2(inbar[181]), .ZN(n558bar);
  OR2_X1 U416 ( .A1(n556), .A2(n555), .ZN(n564) );
  AND2_X1 U416bar ( .A1(n556bar), .A2(n555bar), .ZN(n564bar);
  OR2_X1 U417 ( .A1(n554), .A2(n553), .ZN(n555) );
  AND2_X1 U417bar ( .A1(n554bar), .A2(n553bar), .ZN(n555bar);
  OR2_X1 U418 ( .A1(in_13), .A2(in[234]), .ZN(n553) );
  AND2_X1 U418bar ( .A1(in_13bar), .A2(inbar[234]), .ZN(n553bar);
  OR2_X1 U419 ( .A1(in_38), .A2(in_32), .ZN(n554) );
  AND2_X1 U419bar ( .A1(in_38bar), .A2(in_32bar), .ZN(n554bar);
  OR2_X1 U420 ( .A1(n552), .A2(n551), .ZN(n556) );
  AND2_X1 U420bar ( .A1(n552bar), .A2(n551bar), .ZN(n556bar);
  OR2_X1 U421 ( .A1(in_42), .A2(in_41), .ZN(n551) );
  AND2_X1 U421bar ( .A1(in_42bar), .A2(in_41bar), .ZN(n551bar);
  OR2_X1 U422 ( .A1(in_7), .A2(in_49), .ZN(n552) );
  AND2_X1 U422bar ( .A1(in_7bar), .A2(in_49bar), .ZN(n552bar);
  OR2_X1 U423 ( .A1(n550), .A2(n549), .ZN(n817) );
  AND2_X1 U423bar ( .A1(n550bar), .A2(n549bar), .ZN(n817bar);
  OR2_X1 U424 ( .A1(n548), .A2(n547), .ZN(n549) );
  AND2_X1 U424bar ( .A1(n548bar), .A2(n547bar), .ZN(n549bar);
  OR2_X1 U425 ( .A1(n546), .A2(n545), .ZN(n547) );
  AND2_X1 U425bar ( .A1(n546bar), .A2(n545bar), .ZN(n547bar);
  OR2_X1 U426 ( .A1(in[159]), .A2(in[105]), .ZN(n545) );
  AND2_X1 U426bar ( .A1(inbar[159]), .A2(inbar[105]), .ZN(n545bar);
  OR2_X1 U427 ( .A1(in[206]), .A2(in[183]), .ZN(n546) );
  AND2_X1 U427bar ( .A1(inbar[206]), .A2(inbar[183]), .ZN(n546bar);
  OR2_X1 U428 ( .A1(n544), .A2(n543), .ZN(n548) );
  AND2_X1 U428bar ( .A1(n544bar), .A2(n543bar), .ZN(n548bar);
  OR2_X1 U429 ( .A1(in[229]), .A2(in[219]), .ZN(n543) );
  AND2_X1 U429bar ( .A1(inbar[229]), .A2(inbar[219]), .ZN(n543bar);
  OR2_X1 U430 ( .A1(in[235]), .A2(in[232]), .ZN(n544) );
  AND2_X1 U430bar ( .A1(inbar[235]), .A2(inbar[232]), .ZN(n544bar);
  OR2_X1 U431 ( .A1(n542), .A2(n541), .ZN(n550) );
  AND2_X1 U431bar ( .A1(n542bar), .A2(n541bar), .ZN(n550bar);
  OR2_X1 U432 ( .A1(n540), .A2(n539), .ZN(n541) );
  AND2_X1 U432bar ( .A1(n540bar), .A2(n539bar), .ZN(n541bar);
  OR2_X1 U433 ( .A1(in[249]), .A2(in[242]), .ZN(n539) );
  AND2_X1 U433bar ( .A1(inbar[249]), .A2(inbar[242]), .ZN(n539bar);
  OR2_X1 U434 ( .A1(in[89]), .A2(in[254]), .ZN(n540) );
  AND2_X1 U434bar ( .A1(inbar[89]), .A2(inbar[254]), .ZN(n540bar);
  OR2_X1 U435 ( .A1(n538), .A2(n537), .ZN(n542) );
  AND2_X1 U435bar ( .A1(n538bar), .A2(n537bar), .ZN(n542bar);
  OR2_X1 U436 ( .A1(in_14), .A2(in[99]), .ZN(n537) );
  AND2_X1 U436bar ( .A1(in_14bar), .A2(inbar[99]), .ZN(n537bar);
  OR2_X1 U437 ( .A1(in_60), .A2(in_18), .ZN(n538) );
  AND2_X1 U437bar ( .A1(in_60bar), .A2(in_18bar), .ZN(n538bar);
  OR2_X1 U438 ( .A1(in[113]), .A2(n763), .ZN(n566) );
  AND2_X1 U438bar ( .A1(inbar[113]), .A2(n763bar), .ZN(n566bar);
  OR2_X1 U439 ( .A1(n536), .A2(n535), .ZN(n763) );
  AND2_X1 U439bar ( .A1(n536bar), .A2(n535bar), .ZN(n763bar);
  OR2_X1 U440 ( .A1(n534), .A2(n533), .ZN(n535) );
  AND2_X1 U440bar ( .A1(n534bar), .A2(n533bar), .ZN(n535bar);
  OR2_X1 U441 ( .A1(n532), .A2(n531), .ZN(n533) );
  AND2_X1 U441bar ( .A1(n532bar), .A2(n531bar), .ZN(n533bar);
  OR2_X1 U442 ( .A1(in[115]), .A2(in[110]), .ZN(n531) );
  AND2_X1 U442bar ( .A1(inbar[115]), .A2(inbar[110]), .ZN(n531bar);
  OR2_X1 U443 ( .A1(in[125]), .A2(in[117]), .ZN(n532) );
  AND2_X1 U443bar ( .A1(inbar[125]), .A2(inbar[117]), .ZN(n532bar);
  OR2_X1 U444 ( .A1(n530), .A2(n529), .ZN(n534) );
  AND2_X1 U444bar ( .A1(n530bar), .A2(n529bar), .ZN(n534bar);
  OR2_X1 U445 ( .A1(in[180]), .A2(in[128]), .ZN(n529) );
  AND2_X1 U445bar ( .A1(inbar[180]), .A2(inbar[128]), .ZN(n529bar);
  OR2_X1 U446 ( .A1(in[205]), .A2(in[201]), .ZN(n530) );
  AND2_X1 U446bar ( .A1(inbar[205]), .A2(inbar[201]), .ZN(n530bar);
  OR2_X1 U447 ( .A1(n528), .A2(n527), .ZN(n536) );
  AND2_X1 U447bar ( .A1(n528bar), .A2(n527bar), .ZN(n536bar);
  OR2_X1 U448 ( .A1(n526), .A2(n525), .ZN(n527) );
  AND2_X1 U448bar ( .A1(n526bar), .A2(n525bar), .ZN(n527bar);
  OR2_X1 U449 ( .A1(in[244]), .A2(in[239]), .ZN(n525) );
  AND2_X1 U449bar ( .A1(inbar[244]), .A2(inbar[239]), .ZN(n525bar);
  OR2_X1 U450 ( .A1(in[95]), .A2(in[83]), .ZN(n526) );
  AND2_X1 U450bar ( .A1(inbar[95]), .A2(inbar[83]), .ZN(n526bar);
  OR2_X1 U451 ( .A1(n524), .A2(n523), .ZN(n528) );
  AND2_X1 U451bar ( .A1(n524bar), .A2(n523bar), .ZN(n528bar);
  OR2_X1 U452 ( .A1(in_24), .A2(in[97]), .ZN(n523) );
  AND2_X1 U452bar ( .A1(in_24bar), .A2(inbar[97]), .ZN(n523bar);
  OR2_X1 U453 ( .A1(in_33), .A2(in_27), .ZN(n524) );
  AND2_X1 U453bar ( .A1(in_33bar), .A2(in_27bar), .ZN(n524bar);
  OR2_X1 U454 ( .A1(n522), .A2(n521), .ZN(n568) );
  AND2_X1 U454bar ( .A1(n522bar), .A2(n521bar), .ZN(n568bar);
  OR2_X1 U455 ( .A1(in[145]), .A2(in[126]), .ZN(n521) );
  AND2_X1 U455bar ( .A1(inbar[145]), .A2(inbar[126]), .ZN(n521bar);
  OR2_X1 U456 ( .A1(in[169]), .A2(n520), .ZN(n522) );
  AND2_X1 U456bar ( .A1(inbar[169]), .A2(n520bar), .ZN(n522bar);
  OR2_X1 U457 ( .A1(in[221]), .A2(in[172]), .ZN(n520) );
  AND2_X1 U457bar ( .A1(inbar[221]), .A2(inbar[172]), .ZN(n520bar);
  OR2_X1 U458 ( .A1(n519), .A2(n518), .ZN(n570) );
  AND2_X1 U458bar ( .A1(n519bar), .A2(n518bar), .ZN(n570bar);
  OR2_X1 U459 ( .A1(n517), .A2(n516), .ZN(n518) );
  AND2_X1 U459bar ( .A1(n517bar), .A2(n516bar), .ZN(n518bar);
  OR2_X1 U460 ( .A1(in[241]), .A2(in[224]), .ZN(n516) );
  AND2_X1 U460bar ( .A1(inbar[241]), .A2(inbar[224]), .ZN(n516bar);
  OR2_X1 U461 ( .A1(in[86]), .A2(n515), .ZN(n517) );
  AND2_X1 U461bar ( .A1(inbar[86]), .A2(n515bar), .ZN(n517bar);
  OR2_X1 U462 ( .A1(in_43), .A2(in_34), .ZN(n515) );
  AND2_X1 U462bar ( .A1(in_43bar), .A2(in_34bar), .ZN(n515bar);
  OR2_X1 U463 ( .A1(n514), .A2(n513), .ZN(n519) );
  AND2_X1 U463bar ( .A1(n514bar), .A2(n513bar), .ZN(n519bar);
  OR2_X1 U464 ( .A1(in_65), .A2(in_51), .ZN(n513) );
  AND2_X1 U464bar ( .A1(in_65bar), .A2(in_51bar), .ZN(n513bar);
  OR2_X1 U465 ( .A1(in_75), .A2(n512), .ZN(n514) );
  AND2_X1 U465bar ( .A1(in_75bar), .A2(n512bar), .ZN(n514bar);
  OR2_X1 U466 ( .A1(in_81), .A2(in_77), .ZN(n512) );
  AND2_X1 U466bar ( .A1(in_81bar), .A2(in_77bar), .ZN(n512bar);
  OR2_X1 U467 ( .A1(n511), .A2(n510), .ZN(n778) );
  AND2_X1 U467bar ( .A1(n511bar), .A2(n510bar), .ZN(n778bar);
  OR2_X1 U468 ( .A1(n509), .A2(n508), .ZN(n510) );
  AND2_X1 U468bar ( .A1(n509bar), .A2(n508bar), .ZN(n510bar);
  OR2_X1 U469 ( .A1(n507), .A2(n506), .ZN(n508) );
  AND2_X1 U469bar ( .A1(n507bar), .A2(n506bar), .ZN(n508bar);
  OR2_X1 U470 ( .A1(in[107]), .A2(in[101]), .ZN(n506) );
  AND2_X1 U470bar ( .A1(inbar[107]), .A2(inbar[101]), .ZN(n506bar);
  OR2_X1 U471 ( .A1(in[139]), .A2(in[132]), .ZN(n507) );
  AND2_X1 U471bar ( .A1(inbar[139]), .A2(inbar[132]), .ZN(n507bar);
  OR2_X1 U472 ( .A1(n505), .A2(n504), .ZN(n509) );
  AND2_X1 U472bar ( .A1(n505bar), .A2(n504bar), .ZN(n509bar);
  OR2_X1 U473 ( .A1(in[146]), .A2(in[141]), .ZN(n504) );
  AND2_X1 U473bar ( .A1(inbar[146]), .A2(inbar[141]), .ZN(n504bar);
  OR2_X1 U474 ( .A1(in[203]), .A2(in[179]), .ZN(n505) );
  AND2_X1 U474bar ( .A1(inbar[203]), .A2(inbar[179]), .ZN(n505bar);
  OR2_X1 U475 ( .A1(n503), .A2(n502), .ZN(n511) );
  AND2_X1 U475bar ( .A1(n503bar), .A2(n502bar), .ZN(n511bar);
  OR2_X1 U476 ( .A1(n501), .A2(n500), .ZN(n502) );
  AND2_X1 U476bar ( .A1(n501bar), .A2(n500bar), .ZN(n502bar);
  OR2_X1 U477 ( .A1(in[243]), .A2(in[222]), .ZN(n500) );
  AND2_X1 U477bar ( .A1(inbar[243]), .A2(inbar[222]), .ZN(n500bar);
  OR2_X1 U478 ( .A1(in[251]), .A2(in[250]), .ZN(n501) );
  AND2_X1 U478bar ( .A1(inbar[251]), .A2(inbar[250]), .ZN(n501bar);
  OR2_X1 U479 ( .A1(n499), .A2(n498), .ZN(n503) );
  AND2_X1 U479bar ( .A1(n499bar), .A2(n498bar), .ZN(n503bar);
  OR2_X1 U480 ( .A1(in_37), .A2(in_19), .ZN(n498) );
  AND2_X1 U480bar ( .A1(in_37bar), .A2(in_19bar), .ZN(n498bar);
  OR2_X1 U481 ( .A1(in_78), .A2(in_6), .ZN(n499) );
  AND2_X1 U481bar ( .A1(in_78bar), .A2(in_6bar), .ZN(n499bar);
  OR2_X1 U482 ( .A1(n497), .A2(n496), .ZN(n603) );
  AND2_X1 U482bar ( .A1(n497bar), .A2(n496bar), .ZN(n603bar);
  OR2_X1 U483 ( .A1(in[112]), .A2(in[102]), .ZN(n496) );
  AND2_X1 U483bar ( .A1(inbar[112]), .A2(inbar[102]), .ZN(n496bar);
  OR2_X1 U484 ( .A1(in[123]), .A2(n495), .ZN(n497) );
  AND2_X1 U484bar ( .A1(inbar[123]), .A2(n495bar), .ZN(n497bar);
  OR2_X1 U485 ( .A1(in[143]), .A2(in[130]), .ZN(n495) );
  AND2_X1 U485bar ( .A1(inbar[143]), .A2(inbar[130]), .ZN(n495bar);
  OR2_X1 U486 ( .A1(n494), .A2(n493), .ZN(n605) );
  AND2_X1 U486bar ( .A1(n494bar), .A2(n493bar), .ZN(n605bar);
  OR2_X1 U487 ( .A1(n492), .A2(n491), .ZN(n493) );
  AND2_X1 U487bar ( .A1(n492bar), .A2(n491bar), .ZN(n493bar);
  OR2_X1 U488 ( .A1(in[216]), .A2(in[213]), .ZN(n491) );
  AND2_X1 U488bar ( .A1(inbar[216]), .A2(inbar[213]), .ZN(n491bar);
  OR2_X1 U489 ( .A1(in[227]), .A2(n490), .ZN(n492) );
  AND2_X1 U489bar ( .A1(inbar[227]), .A2(n490bar), .ZN(n492bar);
  OR2_X1 U490 ( .A1(in_0), .A2(in[248]), .ZN(n490) );
  AND2_X1 U490bar ( .A1(in_0bar), .A2(inbar[248]), .ZN(n490bar);
  OR2_X1 U491 ( .A1(n489), .A2(n488), .ZN(n494) );
  AND2_X1 U491bar ( .A1(n489bar), .A2(n488bar), .ZN(n494bar);
  OR2_X1 U492 ( .A1(in_46), .A2(in_44), .ZN(n488) );
  AND2_X1 U492bar ( .A1(in_46bar), .A2(in_44bar), .ZN(n488bar);
  OR2_X1 U493 ( .A1(in_50), .A2(n487), .ZN(n489) );
  AND2_X1 U493bar ( .A1(in_50bar), .A2(n487bar), .ZN(n489bar);
  OR2_X1 U494 ( .A1(in_9), .A2(in_80), .ZN(n487) );
  AND2_X1 U494bar ( .A1(in_9bar), .A2(in_80bar), .ZN(n487bar);
endmodule




module sBox_14 ( in, out );
  input [7:0] in;
  //input_done

  output [7:0] out;
  //output_done

  wire   [255:0] decodeOut;
  //wire_done

  decode_14 dec ( .in(in), .out(decodeOut) );
  encode_14 enc ( .in(decodeOut), .out(out) );
endmodule


module CD2_57 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_58 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_59 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_60 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD4_29 ( a, b, y );
  input [3:0] a;
  input [3:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  //input_done

  output [15:0] y;
  reg [15:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]);
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]);
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]);
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]);
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]);
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]);
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]);
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]);
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]);
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]);
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]);
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]);
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]);
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]);
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]);
endmodule




module CD4_30 ( a, b, y );
  input [3:0] a;
  input [3:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  //input_done

  output [15:0] y;
  reg [15:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]);
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]);
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]);
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]);
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]);
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]);
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]);
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]);
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]);
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]);
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]);
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]);
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]);
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]);
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]);
endmodule




module CD16_15 ( a, b, y );
  input [15:0] a;
  input [15:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign abar[8] = ~a[8];
  assign abar[9] = ~a[9];
  assign abar[10] = ~a[10];
  assign abar[11] = ~a[11];
  assign abar[12] = ~a[12];
  assign abar[13] = ~a[13];
  assign abar[14] = ~a[14];
  assign abar[15] = ~a[15];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign bbar[8] = ~b[8];
  assign bbar[9] = ~b[9];
  assign bbar[10] = ~b[10];
  assign bbar[11] = ~b[11];
  assign bbar[12] = ~b[12];
  assign bbar[13] = ~b[13];
  assign bbar[14] = ~b[14];
  assign bbar[15] = ~b[15];
  //input_done

  output [255:0] y;
  reg [255:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[9]), .A2(a[0]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[9]), .A2(abar[0]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[3]), .A2(a[6]), .ZN(y[99]) );
  OR2_X1 U2bar ( .A1(bbar[3]), .A2(abar[6]), .ZN(ybar[99]);
  AND2_X1 U3 ( .A1(b[2]), .A2(a[6]), .ZN(y[98]) );
  OR2_X1 U3bar ( .A1(bbar[2]), .A2(abar[6]), .ZN(ybar[98]);
  AND2_X1 U4 ( .A1(b[1]), .A2(a[6]), .ZN(y[97]) );
  OR2_X1 U4bar ( .A1(bbar[1]), .A2(abar[6]), .ZN(ybar[97]);
  AND2_X1 U5 ( .A1(b[0]), .A2(a[6]), .ZN(y[96]) );
  OR2_X1 U5bar ( .A1(bbar[0]), .A2(abar[6]), .ZN(ybar[96]);
  AND2_X1 U6 ( .A1(b[15]), .A2(a[5]), .ZN(y[95]) );
  OR2_X1 U6bar ( .A1(bbar[15]), .A2(abar[5]), .ZN(ybar[95]);
  AND2_X1 U7 ( .A1(b[14]), .A2(a[5]), .ZN(y[94]) );
  OR2_X1 U7bar ( .A1(bbar[14]), .A2(abar[5]), .ZN(ybar[94]);
  AND2_X1 U8 ( .A1(b[13]), .A2(a[5]), .ZN(y[93]) );
  OR2_X1 U8bar ( .A1(bbar[13]), .A2(abar[5]), .ZN(ybar[93]);
  AND2_X1 U9 ( .A1(b[12]), .A2(a[5]), .ZN(y[92]) );
  OR2_X1 U9bar ( .A1(bbar[12]), .A2(abar[5]), .ZN(ybar[92]);
  AND2_X1 U10 ( .A1(b[11]), .A2(a[5]), .ZN(y[91]) );
  OR2_X1 U10bar ( .A1(bbar[11]), .A2(abar[5]), .ZN(ybar[91]);
  AND2_X1 U11 ( .A1(b[10]), .A2(a[5]), .ZN(y[90]) );
  OR2_X1 U11bar ( .A1(bbar[10]), .A2(abar[5]), .ZN(ybar[90]);
  AND2_X1 U12 ( .A1(b[8]), .A2(a[0]), .ZN(y[8]) );
  OR2_X1 U12bar ( .A1(bbar[8]), .A2(abar[0]), .ZN(ybar[8]);
  AND2_X1 U13 ( .A1(a[5]), .A2(b[9]), .ZN(y[89]) );
  OR2_X1 U13bar ( .A1(abar[5]), .A2(bbar[9]), .ZN(ybar[89]);
  AND2_X1 U14 ( .A1(b[8]), .A2(a[5]), .ZN(y[88]) );
  OR2_X1 U14bar ( .A1(bbar[8]), .A2(abar[5]), .ZN(ybar[88]);
  AND2_X1 U15 ( .A1(b[7]), .A2(a[5]), .ZN(y[87]) );
  OR2_X1 U15bar ( .A1(bbar[7]), .A2(abar[5]), .ZN(ybar[87]);
  AND2_X1 U16 ( .A1(b[6]), .A2(a[5]), .ZN(y[86]) );
  OR2_X1 U16bar ( .A1(bbar[6]), .A2(abar[5]), .ZN(ybar[86]);
  AND2_X1 U17 ( .A1(b[5]), .A2(a[5]), .ZN(y[85]) );
  OR2_X1 U17bar ( .A1(bbar[5]), .A2(abar[5]), .ZN(ybar[85]);
  AND2_X1 U18 ( .A1(b[4]), .A2(a[5]), .ZN(y[84]) );
  OR2_X1 U18bar ( .A1(bbar[4]), .A2(abar[5]), .ZN(ybar[84]);
  AND2_X1 U19 ( .A1(a[5]), .A2(b[3]), .ZN(y[83]) );
  OR2_X1 U19bar ( .A1(abar[5]), .A2(bbar[3]), .ZN(ybar[83]);
  AND2_X1 U20 ( .A1(a[5]), .A2(b[2]), .ZN(y[82]) );
  OR2_X1 U20bar ( .A1(abar[5]), .A2(bbar[2]), .ZN(ybar[82]);
  AND2_X1 U21 ( .A1(a[5]), .A2(b[1]), .ZN(y[81]) );
  OR2_X1 U21bar ( .A1(abar[5]), .A2(bbar[1]), .ZN(ybar[81]);
  AND2_X1 U22 ( .A1(a[5]), .A2(b[0]), .ZN(y[80]) );
  OR2_X1 U22bar ( .A1(abar[5]), .A2(bbar[0]), .ZN(ybar[80]);
  AND2_X1 U23 ( .A1(b[7]), .A2(a[0]), .ZN(y[7]) );
  OR2_X1 U23bar ( .A1(bbar[7]), .A2(abar[0]), .ZN(ybar[7]);
  AND2_X1 U24 ( .A1(a[4]), .A2(b[15]), .ZN(y[79]) );
  OR2_X1 U24bar ( .A1(abar[4]), .A2(bbar[15]), .ZN(ybar[79]);
  AND2_X1 U25 ( .A1(a[4]), .A2(b[14]), .ZN(y[78]) );
  OR2_X1 U25bar ( .A1(abar[4]), .A2(bbar[14]), .ZN(ybar[78]);
  AND2_X1 U26 ( .A1(a[4]), .A2(b[13]), .ZN(y[77]) );
  OR2_X1 U26bar ( .A1(abar[4]), .A2(bbar[13]), .ZN(ybar[77]);
  AND2_X1 U27 ( .A1(a[4]), .A2(b[12]), .ZN(y[76]) );
  OR2_X1 U27bar ( .A1(abar[4]), .A2(bbar[12]), .ZN(ybar[76]);
  AND2_X1 U28 ( .A1(a[4]), .A2(b[11]), .ZN(y[75]) );
  OR2_X1 U28bar ( .A1(abar[4]), .A2(bbar[11]), .ZN(ybar[75]);
  AND2_X1 U29 ( .A1(a[4]), .A2(b[10]), .ZN(y[74]) );
  OR2_X1 U29bar ( .A1(abar[4]), .A2(bbar[10]), .ZN(ybar[74]);
  AND2_X1 U30 ( .A1(a[4]), .A2(b[9]), .ZN(y[73]) );
  OR2_X1 U30bar ( .A1(abar[4]), .A2(bbar[9]), .ZN(ybar[73]);
  AND2_X1 U31 ( .A1(a[4]), .A2(b[8]), .ZN(y[72]) );
  OR2_X1 U31bar ( .A1(abar[4]), .A2(bbar[8]), .ZN(ybar[72]);
  AND2_X1 U32 ( .A1(a[4]), .A2(b[7]), .ZN(y[71]) );
  OR2_X1 U32bar ( .A1(abar[4]), .A2(bbar[7]), .ZN(ybar[71]);
  AND2_X1 U33 ( .A1(a[4]), .A2(b[6]), .ZN(y[70]) );
  OR2_X1 U33bar ( .A1(abar[4]), .A2(bbar[6]), .ZN(ybar[70]);
  AND2_X1 U34 ( .A1(b[6]), .A2(a[0]), .ZN(y[6]) );
  OR2_X1 U34bar ( .A1(bbar[6]), .A2(abar[0]), .ZN(ybar[6]);
  AND2_X1 U35 ( .A1(a[4]), .A2(b[5]), .ZN(y[69]) );
  OR2_X1 U35bar ( .A1(abar[4]), .A2(bbar[5]), .ZN(ybar[69]);
  AND2_X1 U36 ( .A1(a[4]), .A2(b[4]), .ZN(y[68]) );
  OR2_X1 U36bar ( .A1(abar[4]), .A2(bbar[4]), .ZN(ybar[68]);
  AND2_X1 U37 ( .A1(a[4]), .A2(b[3]), .ZN(y[67]) );
  OR2_X1 U37bar ( .A1(abar[4]), .A2(bbar[3]), .ZN(ybar[67]);
  AND2_X1 U38 ( .A1(a[4]), .A2(b[2]), .ZN(y[66]) );
  OR2_X1 U38bar ( .A1(abar[4]), .A2(bbar[2]), .ZN(ybar[66]);
  AND2_X1 U39 ( .A1(a[4]), .A2(b[1]), .ZN(y[65]) );
  OR2_X1 U39bar ( .A1(abar[4]), .A2(bbar[1]), .ZN(ybar[65]);
  AND2_X1 U40 ( .A1(a[4]), .A2(b[0]), .ZN(y[64]) );
  OR2_X1 U40bar ( .A1(abar[4]), .A2(bbar[0]), .ZN(ybar[64]);
  AND2_X1 U41 ( .A1(a[3]), .A2(b[15]), .ZN(y[63]) );
  OR2_X1 U41bar ( .A1(abar[3]), .A2(bbar[15]), .ZN(ybar[63]);
  AND2_X1 U42 ( .A1(a[3]), .A2(b[14]), .ZN(y[62]) );
  OR2_X1 U42bar ( .A1(abar[3]), .A2(bbar[14]), .ZN(ybar[62]);
  AND2_X1 U43 ( .A1(a[3]), .A2(b[13]), .ZN(y[61]) );
  OR2_X1 U43bar ( .A1(abar[3]), .A2(bbar[13]), .ZN(ybar[61]);
  AND2_X1 U44 ( .A1(a[3]), .A2(b[12]), .ZN(y[60]) );
  OR2_X1 U44bar ( .A1(abar[3]), .A2(bbar[12]), .ZN(ybar[60]);
  AND2_X1 U45 ( .A1(b[5]), .A2(a[0]), .ZN(y[5]) );
  OR2_X1 U45bar ( .A1(bbar[5]), .A2(abar[0]), .ZN(ybar[5]);
  AND2_X1 U46 ( .A1(a[3]), .A2(b[11]), .ZN(y[59]) );
  OR2_X1 U46bar ( .A1(abar[3]), .A2(bbar[11]), .ZN(ybar[59]);
  AND2_X1 U47 ( .A1(a[3]), .A2(b[10]), .ZN(y[58]) );
  OR2_X1 U47bar ( .A1(abar[3]), .A2(bbar[10]), .ZN(ybar[58]);
  AND2_X1 U48 ( .A1(a[3]), .A2(b[9]), .ZN(y[57]) );
  OR2_X1 U48bar ( .A1(abar[3]), .A2(bbar[9]), .ZN(ybar[57]);
  AND2_X1 U49 ( .A1(a[3]), .A2(b[8]), .ZN(y[56]) );
  OR2_X1 U49bar ( .A1(abar[3]), .A2(bbar[8]), .ZN(ybar[56]);
  AND2_X1 U50 ( .A1(a[3]), .A2(b[7]), .ZN(y[55]) );
  OR2_X1 U50bar ( .A1(abar[3]), .A2(bbar[7]), .ZN(ybar[55]);
  AND2_X1 U51 ( .A1(a[3]), .A2(b[6]), .ZN(y[54]) );
  OR2_X1 U51bar ( .A1(abar[3]), .A2(bbar[6]), .ZN(ybar[54]);
  AND2_X1 U52 ( .A1(a[3]), .A2(b[5]), .ZN(y[53]) );
  OR2_X1 U52bar ( .A1(abar[3]), .A2(bbar[5]), .ZN(ybar[53]);
  AND2_X1 U53 ( .A1(a[3]), .A2(b[4]), .ZN(y[52]) );
  OR2_X1 U53bar ( .A1(abar[3]), .A2(bbar[4]), .ZN(ybar[52]);
  AND2_X1 U54 ( .A1(a[3]), .A2(b[3]), .ZN(y[51]) );
  OR2_X1 U54bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[51]);
  AND2_X1 U55 ( .A1(a[3]), .A2(b[2]), .ZN(y[50]) );
  OR2_X1 U55bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[50]);
  AND2_X1 U56 ( .A1(b[4]), .A2(a[0]), .ZN(y[4]) );
  OR2_X1 U56bar ( .A1(bbar[4]), .A2(abar[0]), .ZN(ybar[4]);
  AND2_X1 U57 ( .A1(a[3]), .A2(b[1]), .ZN(y[49]) );
  OR2_X1 U57bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[49]);
  AND2_X1 U58 ( .A1(a[3]), .A2(b[0]), .ZN(y[48]) );
  OR2_X1 U58bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[48]);
  AND2_X1 U59 ( .A1(a[2]), .A2(b[15]), .ZN(y[47]) );
  OR2_X1 U59bar ( .A1(abar[2]), .A2(bbar[15]), .ZN(ybar[47]);
  AND2_X1 U60 ( .A1(a[2]), .A2(b[14]), .ZN(y[46]) );
  OR2_X1 U60bar ( .A1(abar[2]), .A2(bbar[14]), .ZN(ybar[46]);
  AND2_X1 U61 ( .A1(a[2]), .A2(b[13]), .ZN(y[45]) );
  OR2_X1 U61bar ( .A1(abar[2]), .A2(bbar[13]), .ZN(ybar[45]);
  AND2_X1 U62 ( .A1(a[2]), .A2(b[12]), .ZN(y[44]) );
  OR2_X1 U62bar ( .A1(abar[2]), .A2(bbar[12]), .ZN(ybar[44]);
  AND2_X1 U63 ( .A1(a[2]), .A2(b[11]), .ZN(y[43]) );
  OR2_X1 U63bar ( .A1(abar[2]), .A2(bbar[11]), .ZN(ybar[43]);
  AND2_X1 U64 ( .A1(a[2]), .A2(b[10]), .ZN(y[42]) );
  OR2_X1 U64bar ( .A1(abar[2]), .A2(bbar[10]), .ZN(ybar[42]);
  AND2_X1 U65 ( .A1(a[2]), .A2(b[9]), .ZN(y[41]) );
  OR2_X1 U65bar ( .A1(abar[2]), .A2(bbar[9]), .ZN(ybar[41]);
  AND2_X1 U66 ( .A1(a[2]), .A2(b[8]), .ZN(y[40]) );
  OR2_X1 U66bar ( .A1(abar[2]), .A2(bbar[8]), .ZN(ybar[40]);
  AND2_X1 U67 ( .A1(b[3]), .A2(a[0]), .ZN(y[3]) );
  OR2_X1 U67bar ( .A1(bbar[3]), .A2(abar[0]), .ZN(ybar[3]);
  AND2_X1 U68 ( .A1(a[2]), .A2(b[7]), .ZN(y[39]) );
  OR2_X1 U68bar ( .A1(abar[2]), .A2(bbar[7]), .ZN(ybar[39]);
  AND2_X1 U69 ( .A1(a[2]), .A2(b[6]), .ZN(y[38]) );
  OR2_X1 U69bar ( .A1(abar[2]), .A2(bbar[6]), .ZN(ybar[38]);
  AND2_X1 U70 ( .A1(a[2]), .A2(b[5]), .ZN(y[37]) );
  OR2_X1 U70bar ( .A1(abar[2]), .A2(bbar[5]), .ZN(ybar[37]);
  AND2_X1 U71 ( .A1(a[2]), .A2(b[4]), .ZN(y[36]) );
  OR2_X1 U71bar ( .A1(abar[2]), .A2(bbar[4]), .ZN(ybar[36]);
  AND2_X1 U72 ( .A1(a[2]), .A2(b[3]), .ZN(y[35]) );
  OR2_X1 U72bar ( .A1(abar[2]), .A2(bbar[3]), .ZN(ybar[35]);
  AND2_X1 U73 ( .A1(a[2]), .A2(b[2]), .ZN(y[34]) );
  OR2_X1 U73bar ( .A1(abar[2]), .A2(bbar[2]), .ZN(ybar[34]);
  AND2_X1 U74 ( .A1(a[2]), .A2(b[1]), .ZN(y[33]) );
  OR2_X1 U74bar ( .A1(abar[2]), .A2(bbar[1]), .ZN(ybar[33]);
  AND2_X1 U75 ( .A1(a[2]), .A2(b[0]), .ZN(y[32]) );
  OR2_X1 U75bar ( .A1(abar[2]), .A2(bbar[0]), .ZN(ybar[32]);
  AND2_X1 U76 ( .A1(a[1]), .A2(b[15]), .ZN(y[31]) );
  OR2_X1 U76bar ( .A1(abar[1]), .A2(bbar[15]), .ZN(ybar[31]);
  AND2_X1 U77 ( .A1(a[1]), .A2(b[14]), .ZN(y[30]) );
  OR2_X1 U77bar ( .A1(abar[1]), .A2(bbar[14]), .ZN(ybar[30]);
  AND2_X1 U78 ( .A1(b[2]), .A2(a[0]), .ZN(y[2]) );
  OR2_X1 U78bar ( .A1(bbar[2]), .A2(abar[0]), .ZN(ybar[2]);
  AND2_X1 U79 ( .A1(a[1]), .A2(b[13]), .ZN(y[29]) );
  OR2_X1 U79bar ( .A1(abar[1]), .A2(bbar[13]), .ZN(ybar[29]);
  AND2_X1 U80 ( .A1(a[1]), .A2(b[12]), .ZN(y[28]) );
  OR2_X1 U80bar ( .A1(abar[1]), .A2(bbar[12]), .ZN(ybar[28]);
  AND2_X1 U81 ( .A1(a[1]), .A2(b[11]), .ZN(y[27]) );
  OR2_X1 U81bar ( .A1(abar[1]), .A2(bbar[11]), .ZN(ybar[27]);
  AND2_X1 U82 ( .A1(a[1]), .A2(b[10]), .ZN(y[26]) );
  OR2_X1 U82bar ( .A1(abar[1]), .A2(bbar[10]), .ZN(ybar[26]);
  AND2_X1 U83 ( .A1(a[1]), .A2(b[9]), .ZN(y[25]) );
  OR2_X1 U83bar ( .A1(abar[1]), .A2(bbar[9]), .ZN(ybar[25]);
  AND2_X1 U84 ( .A1(a[15]), .A2(b[15]), .ZN(y[255]) );
  OR2_X1 U84bar ( .A1(abar[15]), .A2(bbar[15]), .ZN(ybar[255]);
  AND2_X1 U85 ( .A1(a[15]), .A2(b[14]), .ZN(y[254]) );
  OR2_X1 U85bar ( .A1(abar[15]), .A2(bbar[14]), .ZN(ybar[254]);
  AND2_X1 U86 ( .A1(a[15]), .A2(b[13]), .ZN(y[253]) );
  OR2_X1 U86bar ( .A1(abar[15]), .A2(bbar[13]), .ZN(ybar[253]);
  AND2_X1 U87 ( .A1(a[15]), .A2(b[12]), .ZN(y[252]) );
  OR2_X1 U87bar ( .A1(abar[15]), .A2(bbar[12]), .ZN(ybar[252]);
  AND2_X1 U88 ( .A1(a[15]), .A2(b[11]), .ZN(y[251]) );
  OR2_X1 U88bar ( .A1(abar[15]), .A2(bbar[11]), .ZN(ybar[251]);
  AND2_X1 U89 ( .A1(a[15]), .A2(b[10]), .ZN(y[250]) );
  OR2_X1 U89bar ( .A1(abar[15]), .A2(bbar[10]), .ZN(ybar[250]);
  AND2_X1 U90 ( .A1(a[1]), .A2(b[8]), .ZN(y[24]) );
  OR2_X1 U90bar ( .A1(abar[1]), .A2(bbar[8]), .ZN(ybar[24]);
  AND2_X1 U91 ( .A1(a[15]), .A2(b[9]), .ZN(y[249]) );
  OR2_X1 U91bar ( .A1(abar[15]), .A2(bbar[9]), .ZN(ybar[249]);
  AND2_X1 U92 ( .A1(a[15]), .A2(b[8]), .ZN(y[248]) );
  OR2_X1 U92bar ( .A1(abar[15]), .A2(bbar[8]), .ZN(ybar[248]);
  AND2_X1 U93 ( .A1(a[15]), .A2(b[7]), .ZN(y[247]) );
  OR2_X1 U93bar ( .A1(abar[15]), .A2(bbar[7]), .ZN(ybar[247]);
  AND2_X1 U94 ( .A1(a[15]), .A2(b[6]), .ZN(y[246]) );
  OR2_X1 U94bar ( .A1(abar[15]), .A2(bbar[6]), .ZN(ybar[246]);
  AND2_X1 U95 ( .A1(a[15]), .A2(b[5]), .ZN(y[245]) );
  OR2_X1 U95bar ( .A1(abar[15]), .A2(bbar[5]), .ZN(ybar[245]);
  AND2_X1 U96 ( .A1(a[15]), .A2(b[4]), .ZN(y[244]) );
  OR2_X1 U96bar ( .A1(abar[15]), .A2(bbar[4]), .ZN(ybar[244]);
  AND2_X1 U97 ( .A1(a[15]), .A2(b[3]), .ZN(y[243]) );
  OR2_X1 U97bar ( .A1(abar[15]), .A2(bbar[3]), .ZN(ybar[243]);
  AND2_X1 U98 ( .A1(a[15]), .A2(b[2]), .ZN(y[242]) );
  OR2_X1 U98bar ( .A1(abar[15]), .A2(bbar[2]), .ZN(ybar[242]);
  AND2_X1 U99 ( .A1(a[15]), .A2(b[1]), .ZN(y[241]) );
  OR2_X1 U99bar ( .A1(abar[15]), .A2(bbar[1]), .ZN(ybar[241]);
  AND2_X1 U100 ( .A1(a[15]), .A2(b[0]), .ZN(y[240]) );
  OR2_X1 U100bar ( .A1(abar[15]), .A2(bbar[0]), .ZN(ybar[240]);
  AND2_X1 U101 ( .A1(a[1]), .A2(b[7]), .ZN(y[23]) );
  OR2_X1 U101bar ( .A1(abar[1]), .A2(bbar[7]), .ZN(ybar[23]);
  AND2_X1 U102 ( .A1(a[14]), .A2(b[15]), .ZN(y[239]) );
  OR2_X1 U102bar ( .A1(abar[14]), .A2(bbar[15]), .ZN(ybar[239]);
  AND2_X1 U103 ( .A1(a[14]), .A2(b[14]), .ZN(y[238]) );
  OR2_X1 U103bar ( .A1(abar[14]), .A2(bbar[14]), .ZN(ybar[238]);
  AND2_X1 U104 ( .A1(a[14]), .A2(b[13]), .ZN(y[237]) );
  OR2_X1 U104bar ( .A1(abar[14]), .A2(bbar[13]), .ZN(ybar[237]);
  AND2_X1 U105 ( .A1(a[14]), .A2(b[12]), .ZN(y[236]) );
  OR2_X1 U105bar ( .A1(abar[14]), .A2(bbar[12]), .ZN(ybar[236]);
  AND2_X1 U106 ( .A1(a[14]), .A2(b[11]), .ZN(y[235]) );
  OR2_X1 U106bar ( .A1(abar[14]), .A2(bbar[11]), .ZN(ybar[235]);
  AND2_X1 U107 ( .A1(a[14]), .A2(b[10]), .ZN(y[234]) );
  OR2_X1 U107bar ( .A1(abar[14]), .A2(bbar[10]), .ZN(ybar[234]);
  AND2_X1 U108 ( .A1(a[14]), .A2(b[9]), .ZN(y[233]) );
  OR2_X1 U108bar ( .A1(abar[14]), .A2(bbar[9]), .ZN(ybar[233]);
  AND2_X1 U109 ( .A1(a[14]), .A2(b[8]), .ZN(y[232]) );
  OR2_X1 U109bar ( .A1(abar[14]), .A2(bbar[8]), .ZN(ybar[232]);
  AND2_X1 U110 ( .A1(a[14]), .A2(b[7]), .ZN(y[231]) );
  OR2_X1 U110bar ( .A1(abar[14]), .A2(bbar[7]), .ZN(ybar[231]);
  AND2_X1 U111 ( .A1(a[14]), .A2(b[6]), .ZN(y[230]) );
  OR2_X1 U111bar ( .A1(abar[14]), .A2(bbar[6]), .ZN(ybar[230]);
  AND2_X1 U112 ( .A1(a[1]), .A2(b[6]), .ZN(y[22]) );
  OR2_X1 U112bar ( .A1(abar[1]), .A2(bbar[6]), .ZN(ybar[22]);
  AND2_X1 U113 ( .A1(a[14]), .A2(b[5]), .ZN(y[229]) );
  OR2_X1 U113bar ( .A1(abar[14]), .A2(bbar[5]), .ZN(ybar[229]);
  AND2_X1 U114 ( .A1(a[14]), .A2(b[4]), .ZN(y[228]) );
  OR2_X1 U114bar ( .A1(abar[14]), .A2(bbar[4]), .ZN(ybar[228]);
  AND2_X1 U115 ( .A1(a[14]), .A2(b[3]), .ZN(y[227]) );
  OR2_X1 U115bar ( .A1(abar[14]), .A2(bbar[3]), .ZN(ybar[227]);
  AND2_X1 U116 ( .A1(a[14]), .A2(b[2]), .ZN(y[226]) );
  OR2_X1 U116bar ( .A1(abar[14]), .A2(bbar[2]), .ZN(ybar[226]);
  AND2_X1 U117 ( .A1(a[14]), .A2(b[1]), .ZN(y[225]) );
  OR2_X1 U117bar ( .A1(abar[14]), .A2(bbar[1]), .ZN(ybar[225]);
  AND2_X1 U118 ( .A1(a[14]), .A2(b[0]), .ZN(y[224]) );
  OR2_X1 U118bar ( .A1(abar[14]), .A2(bbar[0]), .ZN(ybar[224]);
  AND2_X1 U119 ( .A1(a[13]), .A2(b[15]), .ZN(y[223]) );
  OR2_X1 U119bar ( .A1(abar[13]), .A2(bbar[15]), .ZN(ybar[223]);
  AND2_X1 U120 ( .A1(a[13]), .A2(b[14]), .ZN(y[222]) );
  OR2_X1 U120bar ( .A1(abar[13]), .A2(bbar[14]), .ZN(ybar[222]);
  AND2_X1 U121 ( .A1(a[13]), .A2(b[13]), .ZN(y[221]) );
  OR2_X1 U121bar ( .A1(abar[13]), .A2(bbar[13]), .ZN(ybar[221]);
  AND2_X1 U122 ( .A1(a[13]), .A2(b[12]), .ZN(y[220]) );
  OR2_X1 U122bar ( .A1(abar[13]), .A2(bbar[12]), .ZN(ybar[220]);
  AND2_X1 U123 ( .A1(a[1]), .A2(b[5]), .ZN(y[21]) );
  OR2_X1 U123bar ( .A1(abar[1]), .A2(bbar[5]), .ZN(ybar[21]);
  AND2_X1 U124 ( .A1(a[13]), .A2(b[11]), .ZN(y[219]) );
  OR2_X1 U124bar ( .A1(abar[13]), .A2(bbar[11]), .ZN(ybar[219]);
  AND2_X1 U125 ( .A1(a[13]), .A2(b[10]), .ZN(y[218]) );
  OR2_X1 U125bar ( .A1(abar[13]), .A2(bbar[10]), .ZN(ybar[218]);
  AND2_X1 U126 ( .A1(a[13]), .A2(b[9]), .ZN(y[217]) );
  OR2_X1 U126bar ( .A1(abar[13]), .A2(bbar[9]), .ZN(ybar[217]);
  AND2_X1 U127 ( .A1(a[13]), .A2(b[8]), .ZN(y[216]) );
  OR2_X1 U127bar ( .A1(abar[13]), .A2(bbar[8]), .ZN(ybar[216]);
  AND2_X1 U128 ( .A1(a[13]), .A2(b[7]), .ZN(y[215]) );
  OR2_X1 U128bar ( .A1(abar[13]), .A2(bbar[7]), .ZN(ybar[215]);
  AND2_X1 U129 ( .A1(a[13]), .A2(b[6]), .ZN(y[214]) );
  OR2_X1 U129bar ( .A1(abar[13]), .A2(bbar[6]), .ZN(ybar[214]);
  AND2_X1 U130 ( .A1(a[13]), .A2(b[5]), .ZN(y[213]) );
  OR2_X1 U130bar ( .A1(abar[13]), .A2(bbar[5]), .ZN(ybar[213]);
  AND2_X1 U131 ( .A1(a[13]), .A2(b[4]), .ZN(y[212]) );
  OR2_X1 U131bar ( .A1(abar[13]), .A2(bbar[4]), .ZN(ybar[212]);
  AND2_X1 U132 ( .A1(a[13]), .A2(b[3]), .ZN(y[211]) );
  OR2_X1 U132bar ( .A1(abar[13]), .A2(bbar[3]), .ZN(ybar[211]);
  AND2_X1 U133 ( .A1(a[13]), .A2(b[2]), .ZN(y[210]) );
  OR2_X1 U133bar ( .A1(abar[13]), .A2(bbar[2]), .ZN(ybar[210]);
  AND2_X1 U134 ( .A1(a[1]), .A2(b[4]), .ZN(y[20]) );
  OR2_X1 U134bar ( .A1(abar[1]), .A2(bbar[4]), .ZN(ybar[20]);
  AND2_X1 U135 ( .A1(a[13]), .A2(b[1]), .ZN(y[209]) );
  OR2_X1 U135bar ( .A1(abar[13]), .A2(bbar[1]), .ZN(ybar[209]);
  AND2_X1 U136 ( .A1(a[13]), .A2(b[0]), .ZN(y[208]) );
  OR2_X1 U136bar ( .A1(abar[13]), .A2(bbar[0]), .ZN(ybar[208]);
  AND2_X1 U137 ( .A1(a[12]), .A2(b[15]), .ZN(y[207]) );
  OR2_X1 U137bar ( .A1(abar[12]), .A2(bbar[15]), .ZN(ybar[207]);
  AND2_X1 U138 ( .A1(a[12]), .A2(b[14]), .ZN(y[206]) );
  OR2_X1 U138bar ( .A1(abar[12]), .A2(bbar[14]), .ZN(ybar[206]);
  AND2_X1 U139 ( .A1(a[12]), .A2(b[13]), .ZN(y[205]) );
  OR2_X1 U139bar ( .A1(abar[12]), .A2(bbar[13]), .ZN(ybar[205]);
  AND2_X1 U140 ( .A1(a[12]), .A2(b[12]), .ZN(y[204]) );
  OR2_X1 U140bar ( .A1(abar[12]), .A2(bbar[12]), .ZN(ybar[204]);
  AND2_X1 U141 ( .A1(a[12]), .A2(b[11]), .ZN(y[203]) );
  OR2_X1 U141bar ( .A1(abar[12]), .A2(bbar[11]), .ZN(ybar[203]);
  AND2_X1 U142 ( .A1(a[12]), .A2(b[10]), .ZN(y[202]) );
  OR2_X1 U142bar ( .A1(abar[12]), .A2(bbar[10]), .ZN(ybar[202]);
  AND2_X1 U143 ( .A1(a[12]), .A2(b[9]), .ZN(y[201]) );
  OR2_X1 U143bar ( .A1(abar[12]), .A2(bbar[9]), .ZN(ybar[201]);
  AND2_X1 U144 ( .A1(a[12]), .A2(b[8]), .ZN(y[200]) );
  OR2_X1 U144bar ( .A1(abar[12]), .A2(bbar[8]), .ZN(ybar[200]);
  AND2_X1 U145 ( .A1(b[1]), .A2(a[0]), .ZN(y[1]) );
  OR2_X1 U145bar ( .A1(bbar[1]), .A2(abar[0]), .ZN(ybar[1]);
  AND2_X1 U146 ( .A1(a[1]), .A2(b[3]), .ZN(y[19]) );
  OR2_X1 U146bar ( .A1(abar[1]), .A2(bbar[3]), .ZN(ybar[19]);
  AND2_X1 U147 ( .A1(a[12]), .A2(b[7]), .ZN(y[199]) );
  OR2_X1 U147bar ( .A1(abar[12]), .A2(bbar[7]), .ZN(ybar[199]);
  AND2_X1 U148 ( .A1(a[12]), .A2(b[6]), .ZN(y[198]) );
  OR2_X1 U148bar ( .A1(abar[12]), .A2(bbar[6]), .ZN(ybar[198]);
  AND2_X1 U149 ( .A1(a[12]), .A2(b[5]), .ZN(y[197]) );
  OR2_X1 U149bar ( .A1(abar[12]), .A2(bbar[5]), .ZN(ybar[197]);
  AND2_X1 U150 ( .A1(a[12]), .A2(b[4]), .ZN(y[196]) );
  OR2_X1 U150bar ( .A1(abar[12]), .A2(bbar[4]), .ZN(ybar[196]);
  AND2_X1 U151 ( .A1(a[12]), .A2(b[3]), .ZN(y[195]) );
  OR2_X1 U151bar ( .A1(abar[12]), .A2(bbar[3]), .ZN(ybar[195]);
  AND2_X1 U152 ( .A1(a[12]), .A2(b[2]), .ZN(y[194]) );
  OR2_X1 U152bar ( .A1(abar[12]), .A2(bbar[2]), .ZN(ybar[194]);
  AND2_X1 U153 ( .A1(a[12]), .A2(b[1]), .ZN(y[193]) );
  OR2_X1 U153bar ( .A1(abar[12]), .A2(bbar[1]), .ZN(ybar[193]);
  AND2_X1 U154 ( .A1(a[12]), .A2(b[0]), .ZN(y[192]) );
  OR2_X1 U154bar ( .A1(abar[12]), .A2(bbar[0]), .ZN(ybar[192]);
  AND2_X1 U155 ( .A1(a[11]), .A2(b[15]), .ZN(y[191]) );
  OR2_X1 U155bar ( .A1(abar[11]), .A2(bbar[15]), .ZN(ybar[191]);
  AND2_X1 U156 ( .A1(a[11]), .A2(b[14]), .ZN(y[190]) );
  OR2_X1 U156bar ( .A1(abar[11]), .A2(bbar[14]), .ZN(ybar[190]);
  AND2_X1 U157 ( .A1(a[1]), .A2(b[2]), .ZN(y[18]) );
  OR2_X1 U157bar ( .A1(abar[1]), .A2(bbar[2]), .ZN(ybar[18]);
  AND2_X1 U158 ( .A1(a[11]), .A2(b[13]), .ZN(y[189]) );
  OR2_X1 U158bar ( .A1(abar[11]), .A2(bbar[13]), .ZN(ybar[189]);
  AND2_X1 U159 ( .A1(a[11]), .A2(b[12]), .ZN(y[188]) );
  OR2_X1 U159bar ( .A1(abar[11]), .A2(bbar[12]), .ZN(ybar[188]);
  AND2_X1 U160 ( .A1(a[11]), .A2(b[11]), .ZN(y[187]) );
  OR2_X1 U160bar ( .A1(abar[11]), .A2(bbar[11]), .ZN(ybar[187]);
  AND2_X1 U161 ( .A1(a[11]), .A2(b[10]), .ZN(y[186]) );
  OR2_X1 U161bar ( .A1(abar[11]), .A2(bbar[10]), .ZN(ybar[186]);
  AND2_X1 U162 ( .A1(a[11]), .A2(b[9]), .ZN(y[185]) );
  OR2_X1 U162bar ( .A1(abar[11]), .A2(bbar[9]), .ZN(ybar[185]);
  AND2_X1 U163 ( .A1(a[11]), .A2(b[8]), .ZN(y[184]) );
  OR2_X1 U163bar ( .A1(abar[11]), .A2(bbar[8]), .ZN(ybar[184]);
  AND2_X1 U164 ( .A1(a[11]), .A2(b[7]), .ZN(y[183]) );
  OR2_X1 U164bar ( .A1(abar[11]), .A2(bbar[7]), .ZN(ybar[183]);
  AND2_X1 U165 ( .A1(a[11]), .A2(b[6]), .ZN(y[182]) );
  OR2_X1 U165bar ( .A1(abar[11]), .A2(bbar[6]), .ZN(ybar[182]);
  AND2_X1 U166 ( .A1(a[11]), .A2(b[5]), .ZN(y[181]) );
  OR2_X1 U166bar ( .A1(abar[11]), .A2(bbar[5]), .ZN(ybar[181]);
  AND2_X1 U167 ( .A1(a[11]), .A2(b[4]), .ZN(y[180]) );
  OR2_X1 U167bar ( .A1(abar[11]), .A2(bbar[4]), .ZN(ybar[180]);
  AND2_X1 U168 ( .A1(a[1]), .A2(b[1]), .ZN(y[17]) );
  OR2_X1 U168bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[17]);
  AND2_X1 U169 ( .A1(a[11]), .A2(b[3]), .ZN(y[179]) );
  OR2_X1 U169bar ( .A1(abar[11]), .A2(bbar[3]), .ZN(ybar[179]);
  AND2_X1 U170 ( .A1(a[11]), .A2(b[2]), .ZN(y[178]) );
  OR2_X1 U170bar ( .A1(abar[11]), .A2(bbar[2]), .ZN(ybar[178]);
  AND2_X1 U171 ( .A1(a[11]), .A2(b[1]), .ZN(y[177]) );
  OR2_X1 U171bar ( .A1(abar[11]), .A2(bbar[1]), .ZN(ybar[177]);
  AND2_X1 U172 ( .A1(a[11]), .A2(b[0]), .ZN(y[176]) );
  OR2_X1 U172bar ( .A1(abar[11]), .A2(bbar[0]), .ZN(ybar[176]);
  AND2_X1 U173 ( .A1(a[10]), .A2(b[15]), .ZN(y[175]) );
  OR2_X1 U173bar ( .A1(abar[10]), .A2(bbar[15]), .ZN(ybar[175]);
  AND2_X1 U174 ( .A1(a[10]), .A2(b[14]), .ZN(y[174]) );
  OR2_X1 U174bar ( .A1(abar[10]), .A2(bbar[14]), .ZN(ybar[174]);
  AND2_X1 U175 ( .A1(a[10]), .A2(b[13]), .ZN(y[173]) );
  OR2_X1 U175bar ( .A1(abar[10]), .A2(bbar[13]), .ZN(ybar[173]);
  AND2_X1 U176 ( .A1(a[10]), .A2(b[12]), .ZN(y[172]) );
  OR2_X1 U176bar ( .A1(abar[10]), .A2(bbar[12]), .ZN(ybar[172]);
  AND2_X1 U177 ( .A1(a[10]), .A2(b[11]), .ZN(y[171]) );
  OR2_X1 U177bar ( .A1(abar[10]), .A2(bbar[11]), .ZN(ybar[171]);
  AND2_X1 U178 ( .A1(a[10]), .A2(b[10]), .ZN(y[170]) );
  OR2_X1 U178bar ( .A1(abar[10]), .A2(bbar[10]), .ZN(ybar[170]);
  AND2_X1 U179 ( .A1(a[1]), .A2(b[0]), .ZN(y[16]) );
  OR2_X1 U179bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[16]);
  AND2_X1 U180 ( .A1(a[10]), .A2(b[9]), .ZN(y[169]) );
  OR2_X1 U180bar ( .A1(abar[10]), .A2(bbar[9]), .ZN(ybar[169]);
  AND2_X1 U181 ( .A1(a[10]), .A2(b[8]), .ZN(y[168]) );
  OR2_X1 U181bar ( .A1(abar[10]), .A2(bbar[8]), .ZN(ybar[168]);
  AND2_X1 U182 ( .A1(a[10]), .A2(b[7]), .ZN(y[167]) );
  OR2_X1 U182bar ( .A1(abar[10]), .A2(bbar[7]), .ZN(ybar[167]);
  AND2_X1 U183 ( .A1(a[10]), .A2(b[6]), .ZN(y[166]) );
  OR2_X1 U183bar ( .A1(abar[10]), .A2(bbar[6]), .ZN(ybar[166]);
  AND2_X1 U184 ( .A1(a[10]), .A2(b[5]), .ZN(y[165]) );
  OR2_X1 U184bar ( .A1(abar[10]), .A2(bbar[5]), .ZN(ybar[165]);
  AND2_X1 U185 ( .A1(a[10]), .A2(b[4]), .ZN(y[164]) );
  OR2_X1 U185bar ( .A1(abar[10]), .A2(bbar[4]), .ZN(ybar[164]);
  AND2_X1 U186 ( .A1(a[10]), .A2(b[3]), .ZN(y[163]) );
  OR2_X1 U186bar ( .A1(abar[10]), .A2(bbar[3]), .ZN(ybar[163]);
  AND2_X1 U187 ( .A1(a[10]), .A2(b[2]), .ZN(y[162]) );
  OR2_X1 U187bar ( .A1(abar[10]), .A2(bbar[2]), .ZN(ybar[162]);
  AND2_X1 U188 ( .A1(a[10]), .A2(b[1]), .ZN(y[161]) );
  OR2_X1 U188bar ( .A1(abar[10]), .A2(bbar[1]), .ZN(ybar[161]);
  AND2_X1 U189 ( .A1(a[10]), .A2(b[0]), .ZN(y[160]) );
  OR2_X1 U189bar ( .A1(abar[10]), .A2(bbar[0]), .ZN(ybar[160]);
  AND2_X1 U190 ( .A1(b[15]), .A2(a[0]), .ZN(y[15]) );
  OR2_X1 U190bar ( .A1(bbar[15]), .A2(abar[0]), .ZN(ybar[15]);
  AND2_X1 U191 ( .A1(a[9]), .A2(b[15]), .ZN(y[159]) );
  OR2_X1 U191bar ( .A1(abar[9]), .A2(bbar[15]), .ZN(ybar[159]);
  AND2_X1 U192 ( .A1(a[9]), .A2(b[14]), .ZN(y[158]) );
  OR2_X1 U192bar ( .A1(abar[9]), .A2(bbar[14]), .ZN(ybar[158]);
  AND2_X1 U193 ( .A1(a[9]), .A2(b[13]), .ZN(y[157]) );
  OR2_X1 U193bar ( .A1(abar[9]), .A2(bbar[13]), .ZN(ybar[157]);
  AND2_X1 U194 ( .A1(a[9]), .A2(b[12]), .ZN(y[156]) );
  OR2_X1 U194bar ( .A1(abar[9]), .A2(bbar[12]), .ZN(ybar[156]);
  AND2_X1 U195 ( .A1(a[9]), .A2(b[11]), .ZN(y[155]) );
  OR2_X1 U195bar ( .A1(abar[9]), .A2(bbar[11]), .ZN(ybar[155]);
  AND2_X1 U196 ( .A1(a[9]), .A2(b[10]), .ZN(y[154]) );
  OR2_X1 U196bar ( .A1(abar[9]), .A2(bbar[10]), .ZN(ybar[154]);
  AND2_X1 U197 ( .A1(a[9]), .A2(b[9]), .ZN(y[153]) );
  OR2_X1 U197bar ( .A1(abar[9]), .A2(bbar[9]), .ZN(ybar[153]);
  AND2_X1 U198 ( .A1(a[9]), .A2(b[8]), .ZN(y[152]) );
  OR2_X1 U198bar ( .A1(abar[9]), .A2(bbar[8]), .ZN(ybar[152]);
  AND2_X1 U199 ( .A1(a[9]), .A2(b[7]), .ZN(y[151]) );
  OR2_X1 U199bar ( .A1(abar[9]), .A2(bbar[7]), .ZN(ybar[151]);
  AND2_X1 U200 ( .A1(a[9]), .A2(b[6]), .ZN(y[150]) );
  OR2_X1 U200bar ( .A1(abar[9]), .A2(bbar[6]), .ZN(ybar[150]);
  AND2_X1 U201 ( .A1(b[14]), .A2(a[0]), .ZN(y[14]) );
  OR2_X1 U201bar ( .A1(bbar[14]), .A2(abar[0]), .ZN(ybar[14]);
  AND2_X1 U202 ( .A1(a[9]), .A2(b[5]), .ZN(y[149]) );
  OR2_X1 U202bar ( .A1(abar[9]), .A2(bbar[5]), .ZN(ybar[149]);
  AND2_X1 U203 ( .A1(a[9]), .A2(b[4]), .ZN(y[148]) );
  OR2_X1 U203bar ( .A1(abar[9]), .A2(bbar[4]), .ZN(ybar[148]);
  AND2_X1 U204 ( .A1(a[9]), .A2(b[3]), .ZN(y[147]) );
  OR2_X1 U204bar ( .A1(abar[9]), .A2(bbar[3]), .ZN(ybar[147]);
  AND2_X1 U205 ( .A1(a[9]), .A2(b[2]), .ZN(y[146]) );
  OR2_X1 U205bar ( .A1(abar[9]), .A2(bbar[2]), .ZN(ybar[146]);
  AND2_X1 U206 ( .A1(a[9]), .A2(b[1]), .ZN(y[145]) );
  OR2_X1 U206bar ( .A1(abar[9]), .A2(bbar[1]), .ZN(ybar[145]);
  AND2_X1 U207 ( .A1(a[9]), .A2(b[0]), .ZN(y[144]) );
  OR2_X1 U207bar ( .A1(abar[9]), .A2(bbar[0]), .ZN(ybar[144]);
  AND2_X1 U208 ( .A1(a[8]), .A2(b[15]), .ZN(y[143]) );
  OR2_X1 U208bar ( .A1(abar[8]), .A2(bbar[15]), .ZN(ybar[143]);
  AND2_X1 U209 ( .A1(a[8]), .A2(b[14]), .ZN(y[142]) );
  OR2_X1 U209bar ( .A1(abar[8]), .A2(bbar[14]), .ZN(ybar[142]);
  AND2_X1 U210 ( .A1(a[8]), .A2(b[13]), .ZN(y[141]) );
  OR2_X1 U210bar ( .A1(abar[8]), .A2(bbar[13]), .ZN(ybar[141]);
  AND2_X1 U211 ( .A1(a[8]), .A2(b[12]), .ZN(y[140]) );
  OR2_X1 U211bar ( .A1(abar[8]), .A2(bbar[12]), .ZN(ybar[140]);
  AND2_X1 U212 ( .A1(b[13]), .A2(a[0]), .ZN(y[13]) );
  OR2_X1 U212bar ( .A1(bbar[13]), .A2(abar[0]), .ZN(ybar[13]);
  AND2_X1 U213 ( .A1(a[8]), .A2(b[11]), .ZN(y[139]) );
  OR2_X1 U213bar ( .A1(abar[8]), .A2(bbar[11]), .ZN(ybar[139]);
  AND2_X1 U214 ( .A1(a[8]), .A2(b[10]), .ZN(y[138]) );
  OR2_X1 U214bar ( .A1(abar[8]), .A2(bbar[10]), .ZN(ybar[138]);
  AND2_X1 U215 ( .A1(a[8]), .A2(b[9]), .ZN(y[137]) );
  OR2_X1 U215bar ( .A1(abar[8]), .A2(bbar[9]), .ZN(ybar[137]);
  AND2_X1 U216 ( .A1(a[8]), .A2(b[8]), .ZN(y[136]) );
  OR2_X1 U216bar ( .A1(abar[8]), .A2(bbar[8]), .ZN(ybar[136]);
  AND2_X1 U217 ( .A1(a[8]), .A2(b[7]), .ZN(y[135]) );
  OR2_X1 U217bar ( .A1(abar[8]), .A2(bbar[7]), .ZN(ybar[135]);
  AND2_X1 U218 ( .A1(a[8]), .A2(b[6]), .ZN(y[134]) );
  OR2_X1 U218bar ( .A1(abar[8]), .A2(bbar[6]), .ZN(ybar[134]);
  AND2_X1 U219 ( .A1(a[8]), .A2(b[5]), .ZN(y[133]) );
  OR2_X1 U219bar ( .A1(abar[8]), .A2(bbar[5]), .ZN(ybar[133]);
  AND2_X1 U220 ( .A1(a[8]), .A2(b[4]), .ZN(y[132]) );
  OR2_X1 U220bar ( .A1(abar[8]), .A2(bbar[4]), .ZN(ybar[132]);
  AND2_X1 U221 ( .A1(a[8]), .A2(b[3]), .ZN(y[131]) );
  OR2_X1 U221bar ( .A1(abar[8]), .A2(bbar[3]), .ZN(ybar[131]);
  AND2_X1 U222 ( .A1(a[8]), .A2(b[2]), .ZN(y[130]) );
  OR2_X1 U222bar ( .A1(abar[8]), .A2(bbar[2]), .ZN(ybar[130]);
  AND2_X1 U223 ( .A1(b[12]), .A2(a[0]), .ZN(y[12]) );
  OR2_X1 U223bar ( .A1(bbar[12]), .A2(abar[0]), .ZN(ybar[12]);
  AND2_X1 U224 ( .A1(a[8]), .A2(b[1]), .ZN(y[129]) );
  OR2_X1 U224bar ( .A1(abar[8]), .A2(bbar[1]), .ZN(ybar[129]);
  AND2_X1 U225 ( .A1(a[8]), .A2(b[0]), .ZN(y[128]) );
  OR2_X1 U225bar ( .A1(abar[8]), .A2(bbar[0]), .ZN(ybar[128]);
  AND2_X1 U226 ( .A1(a[7]), .A2(b[15]), .ZN(y[127]) );
  OR2_X1 U226bar ( .A1(abar[7]), .A2(bbar[15]), .ZN(ybar[127]);
  AND2_X1 U227 ( .A1(a[7]), .A2(b[14]), .ZN(y[126]) );
  OR2_X1 U227bar ( .A1(abar[7]), .A2(bbar[14]), .ZN(ybar[126]);
  AND2_X1 U228 ( .A1(a[7]), .A2(b[13]), .ZN(y[125]) );
  OR2_X1 U228bar ( .A1(abar[7]), .A2(bbar[13]), .ZN(ybar[125]);
  AND2_X1 U229 ( .A1(a[7]), .A2(b[12]), .ZN(y[124]) );
  OR2_X1 U229bar ( .A1(abar[7]), .A2(bbar[12]), .ZN(ybar[124]);
  AND2_X1 U230 ( .A1(a[7]), .A2(b[11]), .ZN(y[123]) );
  OR2_X1 U230bar ( .A1(abar[7]), .A2(bbar[11]), .ZN(ybar[123]);
  AND2_X1 U231 ( .A1(a[7]), .A2(b[10]), .ZN(y[122]) );
  OR2_X1 U231bar ( .A1(abar[7]), .A2(bbar[10]), .ZN(ybar[122]);
  AND2_X1 U232 ( .A1(a[7]), .A2(b[9]), .ZN(y[121]) );
  OR2_X1 U232bar ( .A1(abar[7]), .A2(bbar[9]), .ZN(ybar[121]);
  AND2_X1 U233 ( .A1(a[7]), .A2(b[8]), .ZN(y[120]) );
  OR2_X1 U233bar ( .A1(abar[7]), .A2(bbar[8]), .ZN(ybar[120]);
  AND2_X1 U234 ( .A1(b[11]), .A2(a[0]), .ZN(y[11]) );
  OR2_X1 U234bar ( .A1(bbar[11]), .A2(abar[0]), .ZN(ybar[11]);
  AND2_X1 U235 ( .A1(a[7]), .A2(b[7]), .ZN(y[119]) );
  OR2_X1 U235bar ( .A1(abar[7]), .A2(bbar[7]), .ZN(ybar[119]);
  AND2_X1 U236 ( .A1(a[7]), .A2(b[6]), .ZN(y[118]) );
  OR2_X1 U236bar ( .A1(abar[7]), .A2(bbar[6]), .ZN(ybar[118]);
  AND2_X1 U237 ( .A1(a[7]), .A2(b[5]), .ZN(y[117]) );
  OR2_X1 U237bar ( .A1(abar[7]), .A2(bbar[5]), .ZN(ybar[117]);
  AND2_X1 U238 ( .A1(a[7]), .A2(b[4]), .ZN(y[116]) );
  OR2_X1 U238bar ( .A1(abar[7]), .A2(bbar[4]), .ZN(ybar[116]);
  AND2_X1 U239 ( .A1(a[7]), .A2(b[3]), .ZN(y[115]) );
  OR2_X1 U239bar ( .A1(abar[7]), .A2(bbar[3]), .ZN(ybar[115]);
  AND2_X1 U240 ( .A1(a[7]), .A2(b[2]), .ZN(y[114]) );
  OR2_X1 U240bar ( .A1(abar[7]), .A2(bbar[2]), .ZN(ybar[114]);
  AND2_X1 U241 ( .A1(a[7]), .A2(b[1]), .ZN(y[113]) );
  OR2_X1 U241bar ( .A1(abar[7]), .A2(bbar[1]), .ZN(ybar[113]);
  AND2_X1 U242 ( .A1(a[7]), .A2(b[0]), .ZN(y[112]) );
  OR2_X1 U242bar ( .A1(abar[7]), .A2(bbar[0]), .ZN(ybar[112]);
  AND2_X1 U243 ( .A1(b[15]), .A2(a[6]), .ZN(y[111]) );
  OR2_X1 U243bar ( .A1(bbar[15]), .A2(abar[6]), .ZN(ybar[111]);
  AND2_X1 U244 ( .A1(b[14]), .A2(a[6]), .ZN(y[110]) );
  OR2_X1 U244bar ( .A1(bbar[14]), .A2(abar[6]), .ZN(ybar[110]);
  AND2_X1 U245 ( .A1(b[10]), .A2(a[0]), .ZN(y[10]) );
  OR2_X1 U245bar ( .A1(bbar[10]), .A2(abar[0]), .ZN(ybar[10]);
  AND2_X1 U246 ( .A1(b[13]), .A2(a[6]), .ZN(y[109]) );
  OR2_X1 U246bar ( .A1(bbar[13]), .A2(abar[6]), .ZN(ybar[109]);
  AND2_X1 U247 ( .A1(b[12]), .A2(a[6]), .ZN(y[108]) );
  OR2_X1 U247bar ( .A1(bbar[12]), .A2(abar[6]), .ZN(ybar[108]);
  AND2_X1 U248 ( .A1(b[11]), .A2(a[6]), .ZN(y[107]) );
  OR2_X1 U248bar ( .A1(bbar[11]), .A2(abar[6]), .ZN(ybar[107]);
  AND2_X1 U249 ( .A1(b[10]), .A2(a[6]), .ZN(y[106]) );
  OR2_X1 U249bar ( .A1(bbar[10]), .A2(abar[6]), .ZN(ybar[106]);
  AND2_X1 U250 ( .A1(a[6]), .A2(b[9]), .ZN(y[105]) );
  OR2_X1 U250bar ( .A1(abar[6]), .A2(bbar[9]), .ZN(ybar[105]);
  AND2_X1 U251 ( .A1(b[8]), .A2(a[6]), .ZN(y[104]) );
  OR2_X1 U251bar ( .A1(bbar[8]), .A2(abar[6]), .ZN(ybar[104]);
  AND2_X1 U252 ( .A1(b[7]), .A2(a[6]), .ZN(y[103]) );
  OR2_X1 U252bar ( .A1(bbar[7]), .A2(abar[6]), .ZN(ybar[103]);
  AND2_X1 U253 ( .A1(b[6]), .A2(a[6]), .ZN(y[102]) );
  OR2_X1 U253bar ( .A1(bbar[6]), .A2(abar[6]), .ZN(ybar[102]);
  AND2_X1 U254 ( .A1(b[5]), .A2(a[6]), .ZN(y[101]) );
  OR2_X1 U254bar ( .A1(bbar[5]), .A2(abar[6]), .ZN(ybar[101]);
  AND2_X1 U255 ( .A1(b[4]), .A2(a[6]), .ZN(y[100]) );
  OR2_X1 U255bar ( .A1(bbar[4]), .A2(abar[6]), .ZN(ybar[100]);
  AND2_X1 U256 ( .A1(b[0]), .A2(a[0]), .ZN(y[0]) );
  OR2_X1 U256bar ( .A1(bbar[0]), .A2(abar[0]), .ZN(ybar[0]);
endmodule




module decode_15 ( in, out );
  input [7:0] in;
  //input_done

  output [255:0] out;
  //output_done

  wire   [15:0] level1;
  wire   [31:0] level2;
  //wire_done

  CD2_60 cd_l1_1 ( .a(in[1]), .b(in[0]), .y(level1[3:0]) );
  CD2_59 cd_l1_2 ( .a(in[3]), .b(in[2]), .y(level1[7:4]) );
  CD2_58 cd_l1_3 ( .a(in[5]), .b(in[4]), .y(level1[11:8]) );
  CD2_57 cd_l1_4 ( .a(in[7]), .b(in[6]), .y(level1[15:12]) );
  CD4_30 cd_l2_1 ( .a(level1[7:4]), .b(level1[3:0]), .y(level2[15:0]) );
  CD4_29 cd_l2_2 ( .a(level1[15:12]), .b(level1[11:8]), .y(level2[31:16]) );
  CD16_15 cd_l3 ( .a(level2[31:16]), .b(level2[15:0]), .y(out) );
endmodule


module encode_15 ( in, out );
  input [255:0] in;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
  assign inbar[8] = ~in[8];
  assign inbar[9] = ~in[9];
  assign inbar[10] = ~in[10];
  assign inbar[11] = ~in[11];
  assign inbar[12] = ~in[12];
  assign inbar[13] = ~in[13];
  assign inbar[14] = ~in[14];
  assign inbar[15] = ~in[15];
  assign inbar[16] = ~in[16];
  assign inbar[17] = ~in[17];
  assign inbar[18] = ~in[18];
  assign inbar[19] = ~in[19];
  assign inbar[20] = ~in[20];
  assign inbar[21] = ~in[21];
  assign inbar[22] = ~in[22];
  assign inbar[23] = ~in[23];
  assign inbar[24] = ~in[24];
  assign inbar[25] = ~in[25];
  assign inbar[26] = ~in[26];
  assign inbar[27] = ~in[27];
  assign inbar[28] = ~in[28];
  assign inbar[29] = ~in[29];
  assign inbar[30] = ~in[30];
  assign inbar[31] = ~in[31];
  assign inbar[32] = ~in[32];
  assign inbar[33] = ~in[33];
  assign inbar[34] = ~in[34];
  assign inbar[35] = ~in[35];
  assign inbar[36] = ~in[36];
  assign inbar[37] = ~in[37];
  assign inbar[38] = ~in[38];
  assign inbar[39] = ~in[39];
  assign inbar[40] = ~in[40];
  assign inbar[41] = ~in[41];
  assign inbar[42] = ~in[42];
  assign inbar[43] = ~in[43];
  assign inbar[44] = ~in[44];
  assign inbar[45] = ~in[45];
  assign inbar[46] = ~in[46];
  assign inbar[47] = ~in[47];
  assign inbar[48] = ~in[48];
  assign inbar[49] = ~in[49];
  assign inbar[50] = ~in[50];
  assign inbar[51] = ~in[51];
  assign inbar[52] = ~in[52];
  assign inbar[53] = ~in[53];
  assign inbar[54] = ~in[54];
  assign inbar[55] = ~in[55];
  assign inbar[56] = ~in[56];
  assign inbar[57] = ~in[57];
  assign inbar[58] = ~in[58];
  assign inbar[59] = ~in[59];
  assign inbar[60] = ~in[60];
  assign inbar[61] = ~in[61];
  assign inbar[62] = ~in[62];
  assign inbar[63] = ~in[63];
  assign inbar[64] = ~in[64];
  assign inbar[65] = ~in[65];
  assign inbar[66] = ~in[66];
  assign inbar[67] = ~in[67];
  assign inbar[68] = ~in[68];
  assign inbar[69] = ~in[69];
  assign inbar[70] = ~in[70];
  assign inbar[71] = ~in[71];
  assign inbar[72] = ~in[72];
  assign inbar[73] = ~in[73];
  assign inbar[74] = ~in[74];
  assign inbar[75] = ~in[75];
  assign inbar[76] = ~in[76];
  assign inbar[77] = ~in[77];
  assign inbar[78] = ~in[78];
  assign inbar[79] = ~in[79];
  assign inbar[80] = ~in[80];
  assign inbar[81] = ~in[81];
  assign inbar[82] = ~in[82];
  assign inbar[83] = ~in[83];
  assign inbar[84] = ~in[84];
  assign inbar[85] = ~in[85];
  assign inbar[86] = ~in[86];
  assign inbar[87] = ~in[87];
  assign inbar[88] = ~in[88];
  assign inbar[89] = ~in[89];
  assign inbar[90] = ~in[90];
  assign inbar[91] = ~in[91];
  assign inbar[92] = ~in[92];
  assign inbar[93] = ~in[93];
  assign inbar[94] = ~in[94];
  assign inbar[95] = ~in[95];
  assign inbar[96] = ~in[96];
  assign inbar[97] = ~in[97];
  assign inbar[98] = ~in[98];
  assign inbar[99] = ~in[99];
  assign inbar[100] = ~in[100];
  assign inbar[101] = ~in[101];
  assign inbar[102] = ~in[102];
  assign inbar[103] = ~in[103];
  assign inbar[104] = ~in[104];
  assign inbar[105] = ~in[105];
  assign inbar[106] = ~in[106];
  assign inbar[107] = ~in[107];
  assign inbar[108] = ~in[108];
  assign inbar[109] = ~in[109];
  assign inbar[110] = ~in[110];
  assign inbar[111] = ~in[111];
  assign inbar[112] = ~in[112];
  assign inbar[113] = ~in[113];
  assign inbar[114] = ~in[114];
  assign inbar[115] = ~in[115];
  assign inbar[116] = ~in[116];
  assign inbar[117] = ~in[117];
  assign inbar[118] = ~in[118];
  assign inbar[119] = ~in[119];
  assign inbar[120] = ~in[120];
  assign inbar[121] = ~in[121];
  assign inbar[122] = ~in[122];
  assign inbar[123] = ~in[123];
  assign inbar[124] = ~in[124];
  assign inbar[125] = ~in[125];
  assign inbar[126] = ~in[126];
  assign inbar[127] = ~in[127];
  assign inbar[128] = ~in[128];
  assign inbar[129] = ~in[129];
  assign inbar[130] = ~in[130];
  assign inbar[131] = ~in[131];
  assign inbar[132] = ~in[132];
  assign inbar[133] = ~in[133];
  assign inbar[134] = ~in[134];
  assign inbar[135] = ~in[135];
  assign inbar[136] = ~in[136];
  assign inbar[137] = ~in[137];
  assign inbar[138] = ~in[138];
  assign inbar[139] = ~in[139];
  assign inbar[140] = ~in[140];
  assign inbar[141] = ~in[141];
  assign inbar[142] = ~in[142];
  assign inbar[143] = ~in[143];
  assign inbar[144] = ~in[144];
  assign inbar[145] = ~in[145];
  assign inbar[146] = ~in[146];
  assign inbar[147] = ~in[147];
  assign inbar[148] = ~in[148];
  assign inbar[149] = ~in[149];
  assign inbar[150] = ~in[150];
  assign inbar[151] = ~in[151];
  assign inbar[152] = ~in[152];
  assign inbar[153] = ~in[153];
  assign inbar[154] = ~in[154];
  assign inbar[155] = ~in[155];
  assign inbar[156] = ~in[156];
  assign inbar[157] = ~in[157];
  assign inbar[158] = ~in[158];
  assign inbar[159] = ~in[159];
  assign inbar[160] = ~in[160];
  assign inbar[161] = ~in[161];
  assign inbar[162] = ~in[162];
  assign inbar[163] = ~in[163];
  assign inbar[164] = ~in[164];
  assign inbar[165] = ~in[165];
  assign inbar[166] = ~in[166];
  assign inbar[167] = ~in[167];
  assign inbar[168] = ~in[168];
  assign inbar[169] = ~in[169];
  assign inbar[170] = ~in[170];
  assign inbar[171] = ~in[171];
  assign inbar[172] = ~in[172];
  assign inbar[173] = ~in[173];
  assign inbar[174] = ~in[174];
  assign inbar[175] = ~in[175];
  assign inbar[176] = ~in[176];
  assign inbar[177] = ~in[177];
  assign inbar[178] = ~in[178];
  assign inbar[179] = ~in[179];
  assign inbar[180] = ~in[180];
  assign inbar[181] = ~in[181];
  assign inbar[182] = ~in[182];
  assign inbar[183] = ~in[183];
  assign inbar[184] = ~in[184];
  assign inbar[185] = ~in[185];
  assign inbar[186] = ~in[186];
  assign inbar[187] = ~in[187];
  assign inbar[188] = ~in[188];
  assign inbar[189] = ~in[189];
  assign inbar[190] = ~in[190];
  assign inbar[191] = ~in[191];
  assign inbar[192] = ~in[192];
  assign inbar[193] = ~in[193];
  assign inbar[194] = ~in[194];
  assign inbar[195] = ~in[195];
  assign inbar[196] = ~in[196];
  assign inbar[197] = ~in[197];
  assign inbar[198] = ~in[198];
  assign inbar[199] = ~in[199];
  assign inbar[200] = ~in[200];
  assign inbar[201] = ~in[201];
  assign inbar[202] = ~in[202];
  assign inbar[203] = ~in[203];
  assign inbar[204] = ~in[204];
  assign inbar[205] = ~in[205];
  assign inbar[206] = ~in[206];
  assign inbar[207] = ~in[207];
  assign inbar[208] = ~in[208];
  assign inbar[209] = ~in[209];
  assign inbar[210] = ~in[210];
  assign inbar[211] = ~in[211];
  assign inbar[212] = ~in[212];
  assign inbar[213] = ~in[213];
  assign inbar[214] = ~in[214];
  assign inbar[215] = ~in[215];
  assign inbar[216] = ~in[216];
  assign inbar[217] = ~in[217];
  assign inbar[218] = ~in[218];
  assign inbar[219] = ~in[219];
  assign inbar[220] = ~in[220];
  assign inbar[221] = ~in[221];
  assign inbar[222] = ~in[222];
  assign inbar[223] = ~in[223];
  assign inbar[224] = ~in[224];
  assign inbar[225] = ~in[225];
  assign inbar[226] = ~in[226];
  assign inbar[227] = ~in[227];
  assign inbar[228] = ~in[228];
  assign inbar[229] = ~in[229];
  assign inbar[230] = ~in[230];
  assign inbar[231] = ~in[231];
  assign inbar[232] = ~in[232];
  assign inbar[233] = ~in[233];
  assign inbar[234] = ~in[234];
  assign inbar[235] = ~in[235];
  assign inbar[236] = ~in[236];
  assign inbar[237] = ~in[237];
  assign inbar[238] = ~in[238];
  assign inbar[239] = ~in[239];
  assign inbar[240] = ~in[240];
  assign inbar[241] = ~in[241];
  assign inbar[242] = ~in[242];
  assign inbar[243] = ~in[243];
  assign inbar[244] = ~in[244];
  assign inbar[245] = ~in[245];
  assign inbar[246] = ~in[246];
  assign inbar[247] = ~in[247];
  assign inbar[248] = ~in[248];
  assign inbar[249] = ~in[249];
  assign inbar[250] = ~in[250];
  assign inbar[251] = ~in[251];
  assign inbar[252] = ~in[252];
  assign inbar[253] = ~in[253];
  assign inbar[254] = ~in[254];
  assign inbar[255] = ~in[255];
  //input_done

  output [7:0] out;
  reg [7:0] outbar;
  //output_done

  wire   in_81, in_80, in_79, in_78, in_77, in_76, in_75, in_74, in_73, in_72,
         in_71, in_70, in_69, in_68, in_67, in_66, in_65, in_64, in_63, in_62,
         in_61, in_60, in_59, in_58, in_57, in_56, in_55, in_54, in_53, in_52,
         in_51, in_50, in_49, in_48, in_47, in_46, in_45, in_44, in_43, in_42,
         in_41, in_40, in_39, in_38, in_37, in_36, in_35, in_34, in_33, in_32,
         in_31, in_30, in_29, in_28, in_27, in_26, in_25, in_24, in_23, in_22,
         in_21, in_20, in_19, in_18, in_17, in_16, in_15, in_14, in_13, in_12,
         in_11, in_10, in_9, in_8, in_7, in_6, in_5, in_4, in_3, in_2, in_1,
         in_0, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972;
  wire in_81bar, in_80bar, in_79bar, in_78bar, in_77bar, in_76bar, in_75bar, in_74bar, in_73bar, in_72bar, in_71bar, in_70bar, in_69bar, in_68bar, in_67bar, in_66bar, in_65bar, in_64bar, in_63bar, in_62bar, in_61bar, in_60bar, in_59bar, in_58bar, in_57bar, in_56bar, in_55bar, in_54bar, in_53bar, in_52bar, in_51bar, in_50bar, in_49bar, in_48bar, in_47bar, in_46bar, in_45bar, in_44bar, in_43bar, in_42bar, in_41bar, in_40bar, in_39bar, in_38bar, in_37bar, in_36bar, in_35bar, in_34bar, in_33bar, in_32bar, in_31bar, in_30bar, in_29bar, in_28bar, in_27bar, in_26bar, in_25bar, in_24bar, in_23bar, in_22bar, in_21bar, in_20bar, in_19bar, in_18bar, in_17bar, in_16bar, in_15bar, in_14bar, in_13bar, in_12bar, in_11bar, in_10bar, in_9bar, in_8bar, in_7bar, in_6bar, in_5bar, in_4bar, in_3bar, in_2bar, in_1bar, in_0bar, n487bar, n488bar, n489bar, n490bar, n491bar, n492bar, n493bar, n494bar, n495bar, n496bar, n497bar, n498bar, n499bar, n500bar, n501bar, n502bar, n503bar, n504bar, n505bar, n506bar, n507bar, n508bar, n509bar, n510bar, n511bar, n512bar, n513bar, n514bar, n515bar, n516bar, n517bar, n518bar, n519bar, n520bar, n521bar, n522bar, n523bar, n524bar, n525bar, n526bar, n527bar, n528bar, n529bar, n530bar, n531bar, n532bar, n533bar, n534bar, n535bar, n536bar, n537bar, n538bar, n539bar, n540bar, n541bar, n542bar, n543bar, n544bar, n545bar, n546bar, n547bar, n548bar, n549bar, n550bar, n551bar, n552bar, n553bar, n554bar, n555bar, n556bar, n557bar, n558bar, n559bar, n560bar, n561bar, n562bar, n563bar, n564bar, n565bar, n566bar, n567bar, n568bar, n569bar, n570bar, n571bar, n572bar, n573bar, n574bar, n575bar, n576bar, n577bar, n578bar, n579bar, n580bar, n581bar, n582bar, n583bar, n584bar, n585bar, n586bar, n587bar, n588bar, n589bar, n590bar, n591bar, n592bar, n593bar, n594bar, n595bar, n596bar, n597bar, n598bar, n599bar, n600bar, n601bar, n602bar, n603bar, n604bar, n605bar, n606bar, n607bar, n608bar, n609bar, n610bar, n611bar, n612bar, n613bar, n614bar, n615bar, n616bar, n617bar, n618bar, n619bar, n620bar, n621bar, n622bar, n623bar, n624bar, n625bar, n626bar, n627bar, n628bar, n629bar, n630bar, n631bar, n632bar, n633bar, n634bar, n635bar, n636bar, n637bar, n638bar, n639bar, n640bar, n641bar, n642bar, n643bar, n644bar, n645bar, n646bar, n647bar, n648bar, n649bar, n650bar, n651bar, n652bar, n653bar, n654bar, n655bar, n656bar, n657bar, n658bar, n659bar, n660bar, n661bar, n662bar, n663bar, n664bar, n665bar, n666bar, n667bar, n668bar, n669bar, n670bar, n671bar, n672bar, n673bar, n674bar, n675bar, n676bar, n677bar, n678bar, n679bar, n680bar, n681bar, n682bar, n683bar, n684bar, n685bar, n686bar, n687bar, n688bar, n689bar, n690bar, n691bar, n692bar, n693bar, n694bar, n695bar, n696bar, n697bar, n698bar, n699bar, n700bar, n701bar, n702bar, n703bar, n704bar, n705bar, n706bar, n707bar, n708bar, n709bar, n710bar, n711bar, n712bar, n713bar, n714bar, n715bar, n716bar, n717bar, n718bar, n719bar, n720bar, n721bar, n722bar, n723bar, n724bar, n725bar, n726bar, n727bar, n728bar, n729bar, n730bar, n731bar, n732bar, n733bar, n734bar, n735bar, n736bar, n737bar, n738bar, n739bar, n740bar, n741bar, n742bar, n743bar, n744bar, n745bar, n746bar, n747bar, n748bar, n749bar, n750bar, n751bar, n752bar, n753bar, n754bar, n755bar, n756bar, n757bar, n758bar, n759bar, n760bar, n761bar, n762bar, n763bar, n764bar, n765bar, n766bar, n767bar, n768bar, n769bar, n770bar, n771bar, n772bar, n773bar, n774bar, n775bar, n776bar, n777bar, n778bar, n779bar, n780bar, n781bar, n782bar, n783bar, n784bar, n785bar, n786bar, n787bar, n788bar, n789bar, n790bar, n791bar, n792bar, n793bar, n794bar, n795bar, n796bar, n797bar, n798bar, n799bar, n800bar, n801bar, n802bar, n803bar, n804bar, n805bar, n806bar, n807bar, n808bar, n809bar, n810bar, n811bar, n812bar, n813bar, n814bar, n815bar, n816bar, n817bar, n818bar, n819bar, n820bar, n821bar, n822bar, n823bar, n824bar, n825bar, n826bar, n827bar, n828bar, n829bar, n830bar, n831bar, n832bar, n833bar, n834bar, n835bar, n836bar, n837bar, n838bar, n839bar, n840bar, n841bar, n842bar, n843bar, n844bar, n845bar, n846bar, n847bar, n848bar, n849bar, n850bar, n851bar, n852bar, n853bar, n854bar, n855bar, n856bar, n857bar, n858bar, n859bar, n860bar, n861bar, n862bar, n863bar, n864bar, n865bar, n866bar, n867bar, n868bar, n869bar, n870bar, n871bar, n872bar, n873bar, n874bar, n875bar, n876bar, n877bar, n878bar, n879bar, n880bar, n881bar, n882bar, n883bar, n884bar, n885bar, n886bar, n887bar, n888bar, n889bar, n890bar, n891bar, n892bar, n893bar, n894bar, n895bar, n896bar, n897bar, n898bar, n899bar, n900bar, n901bar, n902bar, n903bar, n904bar, n905bar, n906bar, n907bar, n908bar, n909bar, n910bar, n911bar, n912bar, n913bar, n914bar, n915bar, n916bar, n917bar, n918bar, n919bar, n920bar, n921bar, n922bar, n923bar, n924bar, n925bar, n926bar, n927bar, n928bar, n929bar, n930bar, n931bar, n932bar, n933bar, n934bar, n935bar, n936bar, n937bar, n938bar, n939bar, n940bar, n941bar, n942bar, n943bar, n944bar, n945bar, n946bar, n947bar, n948bar, n949bar, n950bar, n951bar, n952bar, n953bar, n954bar, n955bar, n956bar, n957bar, n958bar, n959bar, n960bar, n961bar, n962bar, n963bar, n964bar, n965bar, n966bar, n967bar, n968bar, n969bar, n970bar, n971bar, n972bar;
  //wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];

  OR2_X1 U1 ( .A1(n972), .A2(n971), .ZN(out[7]) );
  AND2_X1 U1bar ( .A1(n972bar), .A2(n971bar), .ZN(outbar[7]);
  OR2_X1 U2 ( .A1(n970), .A2(n969), .ZN(n971) );
  AND2_X1 U2bar ( .A1(n970bar), .A2(n969bar), .ZN(n971bar);
  OR2_X1 U3 ( .A1(n968), .A2(n967), .ZN(n969) );
  AND2_X1 U3bar ( .A1(n968bar), .A2(n967bar), .ZN(n969bar);
  OR2_X1 U4 ( .A1(n966), .A2(n965), .ZN(n967) );
  AND2_X1 U4bar ( .A1(n966bar), .A2(n965bar), .ZN(n967bar);
  OR2_X1 U5 ( .A1(n964), .A2(n963), .ZN(n968) );
  AND2_X1 U5bar ( .A1(n964bar), .A2(n963bar), .ZN(n968bar);
  OR2_X1 U6 ( .A1(in[116]), .A2(n962), .ZN(n963) );
  AND2_X1 U6bar ( .A1(inbar[116]), .A2(n962bar), .ZN(n963bar);
  OR2_X1 U7 ( .A1(n961), .A2(n960), .ZN(n970) );
  AND2_X1 U7bar ( .A1(n961bar), .A2(n960bar), .ZN(n970bar);
  OR2_X1 U8 ( .A1(in[150]), .A2(in[127]), .ZN(n960) );
  AND2_X1 U8bar ( .A1(inbar[150]), .A2(inbar[127]), .ZN(n960bar);
  OR2_X1 U9 ( .A1(in[160]), .A2(n959), .ZN(n961) );
  AND2_X1 U9bar ( .A1(inbar[160]), .A2(n959bar), .ZN(n961bar);
  OR2_X1 U10 ( .A1(in[252]), .A2(in[168]), .ZN(n959) );
  AND2_X1 U10bar ( .A1(inbar[252]), .A2(inbar[168]), .ZN(n959bar);
  OR2_X1 U11 ( .A1(n958), .A2(n957), .ZN(n972) );
  AND2_X1 U11bar ( .A1(n958bar), .A2(n957bar), .ZN(n972bar);
  OR2_X1 U12 ( .A1(n956), .A2(n955), .ZN(n957) );
  AND2_X1 U12bar ( .A1(n956bar), .A2(n955bar), .ZN(n957bar);
  OR2_X1 U13 ( .A1(in_17), .A2(in[96]), .ZN(n955) );
  AND2_X1 U13bar ( .A1(in_17bar), .A2(inbar[96]), .ZN(n955bar);
  OR2_X1 U14 ( .A1(in_23), .A2(n954), .ZN(n956) );
  AND2_X1 U14bar ( .A1(in_23bar), .A2(n954bar), .ZN(n956bar);
  OR2_X1 U15 ( .A1(in_31), .A2(in_26), .ZN(n954) );
  AND2_X1 U15bar ( .A1(in_31bar), .A2(in_26bar), .ZN(n954bar);
  OR2_X1 U16 ( .A1(n953), .A2(n952), .ZN(n958) );
  AND2_X1 U16bar ( .A1(n953bar), .A2(n952bar), .ZN(n958bar);
  OR2_X1 U17 ( .A1(in_58), .A2(in_4), .ZN(n952) );
  AND2_X1 U17bar ( .A1(in_58bar), .A2(in_4bar), .ZN(n952bar);
  OR2_X1 U18 ( .A1(in_59), .A2(n951), .ZN(n953) );
  AND2_X1 U18bar ( .A1(in_59bar), .A2(n951bar), .ZN(n953bar);
  OR2_X1 U19 ( .A1(in_71), .A2(in_62), .ZN(n951) );
  AND2_X1 U19bar ( .A1(in_71bar), .A2(in_62bar), .ZN(n951bar);
  OR2_X1 U20 ( .A1(n950), .A2(n949), .ZN(out[6]) );
  AND2_X1 U20bar ( .A1(n950bar), .A2(n949bar), .ZN(outbar[6]);
  OR2_X1 U21 ( .A1(n948), .A2(n947), .ZN(n949) );
  AND2_X1 U21bar ( .A1(n948bar), .A2(n947bar), .ZN(n949bar);
  OR2_X1 U22 ( .A1(n946), .A2(n945), .ZN(n947) );
  AND2_X1 U22bar ( .A1(n946bar), .A2(n945bar), .ZN(n947bar);
  OR2_X1 U23 ( .A1(n944), .A2(n943), .ZN(n945) );
  AND2_X1 U23bar ( .A1(n944bar), .A2(n943bar), .ZN(n945bar);
  OR2_X1 U24 ( .A1(n942), .A2(n941), .ZN(n946) );
  AND2_X1 U24bar ( .A1(n942bar), .A2(n941bar), .ZN(n946bar);
  OR2_X1 U25 ( .A1(in[101]), .A2(n940), .ZN(n941) );
  AND2_X1 U25bar ( .A1(inbar[101]), .A2(n940bar), .ZN(n941bar);
  OR2_X1 U26 ( .A1(n939), .A2(n938), .ZN(n948) );
  AND2_X1 U26bar ( .A1(n939bar), .A2(n938bar), .ZN(n948bar);
  OR2_X1 U27 ( .A1(in[114]), .A2(in[104]), .ZN(n938) );
  AND2_X1 U27bar ( .A1(inbar[114]), .A2(inbar[104]), .ZN(n938bar);
  OR2_X1 U28 ( .A1(in[128]), .A2(n937), .ZN(n939) );
  AND2_X1 U28bar ( .A1(inbar[128]), .A2(n937bar), .ZN(n939bar);
  OR2_X1 U29 ( .A1(in[136]), .A2(in[134]), .ZN(n937) );
  AND2_X1 U29bar ( .A1(inbar[136]), .A2(inbar[134]), .ZN(n937bar);
  OR2_X1 U30 ( .A1(n936), .A2(n935), .ZN(n950) );
  AND2_X1 U30bar ( .A1(n936bar), .A2(n935bar), .ZN(n950bar);
  OR2_X1 U31 ( .A1(n934), .A2(n933), .ZN(n935) );
  AND2_X1 U31bar ( .A1(n934bar), .A2(n933bar), .ZN(n935bar);
  OR2_X1 U32 ( .A1(in[177]), .A2(in[164]), .ZN(n933) );
  AND2_X1 U32bar ( .A1(inbar[177]), .A2(inbar[164]), .ZN(n933bar);
  OR2_X1 U33 ( .A1(in[212]), .A2(n932), .ZN(n934) );
  AND2_X1 U33bar ( .A1(inbar[212]), .A2(n932bar), .ZN(n934bar);
  OR2_X1 U34 ( .A1(in[248]), .A2(in[221]), .ZN(n932) );
  AND2_X1 U34bar ( .A1(inbar[248]), .A2(inbar[221]), .ZN(n932bar);
  OR2_X1 U35 ( .A1(n931), .A2(n930), .ZN(n936) );
  AND2_X1 U35bar ( .A1(n931bar), .A2(n930bar), .ZN(n936bar);
  OR2_X1 U36 ( .A1(in_18), .A2(in[93]), .ZN(n930) );
  AND2_X1 U36bar ( .A1(in_18bar), .A2(inbar[93]), .ZN(n930bar);
  OR2_X1 U37 ( .A1(in_31), .A2(n929), .ZN(n931) );
  AND2_X1 U37bar ( .A1(in_31bar), .A2(n929bar), .ZN(n931bar);
  OR2_X1 U38 ( .A1(in_7), .A2(in_39), .ZN(n929) );
  AND2_X1 U38bar ( .A1(in_7bar), .A2(in_39bar), .ZN(n929bar);
  OR2_X1 U39 ( .A1(n928), .A2(n927), .ZN(out[5]) );
  AND2_X1 U39bar ( .A1(n928bar), .A2(n927bar), .ZN(outbar[5]);
  OR2_X1 U40 ( .A1(n926), .A2(n925), .ZN(n927) );
  AND2_X1 U40bar ( .A1(n926bar), .A2(n925bar), .ZN(n927bar);
  OR2_X1 U41 ( .A1(n924), .A2(n923), .ZN(n925) );
  AND2_X1 U41bar ( .A1(n924bar), .A2(n923bar), .ZN(n925bar);
  OR2_X1 U42 ( .A1(n922), .A2(n921), .ZN(n923) );
  AND2_X1 U42bar ( .A1(n922bar), .A2(n921bar), .ZN(n923bar);
  OR2_X1 U43 ( .A1(n940), .A2(n920), .ZN(n924) );
  AND2_X1 U43bar ( .A1(n940bar), .A2(n920bar), .ZN(n924bar);
  OR2_X1 U44 ( .A1(in[111]), .A2(n919), .ZN(n920) );
  AND2_X1 U44bar ( .A1(inbar[111]), .A2(n919bar), .ZN(n920bar);
  OR2_X1 U45 ( .A1(n918), .A2(n917), .ZN(n940) );
  AND2_X1 U45bar ( .A1(n918bar), .A2(n917bar), .ZN(n940bar);
  OR2_X1 U46 ( .A1(n916), .A2(n915), .ZN(n917) );
  AND2_X1 U46bar ( .A1(n916bar), .A2(n915bar), .ZN(n917bar);
  OR2_X1 U47 ( .A1(n914), .A2(n913), .ZN(n915) );
  AND2_X1 U47bar ( .A1(n914bar), .A2(n913bar), .ZN(n915bar);
  OR2_X1 U48 ( .A1(in[140]), .A2(in[131]), .ZN(n913) );
  AND2_X1 U48bar ( .A1(inbar[140]), .A2(inbar[131]), .ZN(n913bar);
  OR2_X1 U49 ( .A1(in[160]), .A2(in[144]), .ZN(n914) );
  AND2_X1 U49bar ( .A1(inbar[160]), .A2(inbar[144]), .ZN(n914bar);
  OR2_X1 U50 ( .A1(n912), .A2(n911), .ZN(n916) );
  AND2_X1 U50bar ( .A1(n912bar), .A2(n911bar), .ZN(n916bar);
  OR2_X1 U51 ( .A1(in[179]), .A2(in[174]), .ZN(n911) );
  AND2_X1 U51bar ( .A1(inbar[179]), .A2(inbar[174]), .ZN(n911bar);
  OR2_X1 U52 ( .A1(in[188]), .A2(in[184]), .ZN(n912) );
  AND2_X1 U52bar ( .A1(inbar[188]), .A2(inbar[184]), .ZN(n912bar);
  OR2_X1 U53 ( .A1(n910), .A2(n909), .ZN(n918) );
  AND2_X1 U53bar ( .A1(n910bar), .A2(n909bar), .ZN(n918bar);
  OR2_X1 U54 ( .A1(n908), .A2(n907), .ZN(n909) );
  AND2_X1 U54bar ( .A1(n908bar), .A2(n907bar), .ZN(n909bar);
  OR2_X1 U55 ( .A1(in[216]), .A2(in[200]), .ZN(n907) );
  AND2_X1 U55bar ( .A1(inbar[216]), .A2(inbar[200]), .ZN(n907bar);
  OR2_X1 U56 ( .A1(in[228]), .A2(in[224]), .ZN(n908) );
  AND2_X1 U56bar ( .A1(inbar[228]), .A2(inbar[224]), .ZN(n908bar);
  OR2_X1 U57 ( .A1(n906), .A2(n905), .ZN(n910) );
  AND2_X1 U57bar ( .A1(n906bar), .A2(n905bar), .ZN(n910bar);
  OR2_X1 U58 ( .A1(in[247]), .A2(in[235]), .ZN(n905) );
  AND2_X1 U58bar ( .A1(inbar[247]), .A2(inbar[235]), .ZN(n905bar);
  OR2_X1 U59 ( .A1(in_42), .A2(in[83]), .ZN(n906) );
  AND2_X1 U59bar ( .A1(in_42bar), .A2(inbar[83]), .ZN(n906bar);
  OR2_X1 U60 ( .A1(n904), .A2(n903), .ZN(n926) );
  AND2_X1 U60bar ( .A1(n904bar), .A2(n903bar), .ZN(n926bar);
  OR2_X1 U61 ( .A1(in[166]), .A2(in[123]), .ZN(n903) );
  AND2_X1 U61bar ( .A1(inbar[166]), .A2(inbar[123]), .ZN(n903bar);
  OR2_X1 U62 ( .A1(in[170]), .A2(n902), .ZN(n904) );
  AND2_X1 U62bar ( .A1(inbar[170]), .A2(n902bar), .ZN(n904bar);
  OR2_X1 U63 ( .A1(in[194]), .A2(in[183]), .ZN(n902) );
  AND2_X1 U63bar ( .A1(inbar[194]), .A2(inbar[183]), .ZN(n902bar);
  OR2_X1 U64 ( .A1(n901), .A2(n900), .ZN(n928) );
  AND2_X1 U64bar ( .A1(n901bar), .A2(n900bar), .ZN(n928bar);
  OR2_X1 U65 ( .A1(n899), .A2(n898), .ZN(n900) );
  AND2_X1 U65bar ( .A1(n899bar), .A2(n898bar), .ZN(n900bar);
  OR2_X1 U66 ( .A1(in[241]), .A2(in[238]), .ZN(n898) );
  AND2_X1 U66bar ( .A1(inbar[241]), .A2(inbar[238]), .ZN(n898bar);
  OR2_X1 U67 ( .A1(in[250]), .A2(n897), .ZN(n899) );
  AND2_X1 U67bar ( .A1(inbar[250]), .A2(n897bar), .ZN(n899bar);
  OR2_X1 U68 ( .A1(in_24), .A2(in[84]), .ZN(n897) );
  AND2_X1 U68bar ( .A1(in_24bar), .A2(inbar[84]), .ZN(n897bar);
  OR2_X1 U69 ( .A1(n896), .A2(n895), .ZN(n901) );
  AND2_X1 U69bar ( .A1(n896bar), .A2(n895bar), .ZN(n901bar);
  OR2_X1 U70 ( .A1(in_41), .A2(in_29), .ZN(n895) );
  AND2_X1 U70bar ( .A1(in_41bar), .A2(in_29bar), .ZN(n895bar);
  OR2_X1 U71 ( .A1(in_66), .A2(n894), .ZN(n896) );
  AND2_X1 U71bar ( .A1(in_66bar), .A2(n894bar), .ZN(n896bar);
  OR2_X1 U72 ( .A1(in_76), .A2(in_71), .ZN(n894) );
  AND2_X1 U72bar ( .A1(in_76bar), .A2(in_71bar), .ZN(n894bar);
  OR2_X1 U73 ( .A1(n893), .A2(n892), .ZN(out[4]) );
  AND2_X1 U73bar ( .A1(n893bar), .A2(n892bar), .ZN(outbar[4]);
  OR2_X1 U74 ( .A1(n891), .A2(n890), .ZN(n892) );
  AND2_X1 U74bar ( .A1(n891bar), .A2(n890bar), .ZN(n892bar);
  OR2_X1 U75 ( .A1(n889), .A2(n888), .ZN(n890) );
  AND2_X1 U75bar ( .A1(n889bar), .A2(n888bar), .ZN(n890bar);
  OR2_X1 U76 ( .A1(n922), .A2(n887), .ZN(n888) );
  AND2_X1 U76bar ( .A1(n922bar), .A2(n887bar), .ZN(n888bar);
  OR2_X1 U77 ( .A1(n886), .A2(n885), .ZN(n922) );
  AND2_X1 U77bar ( .A1(n886bar), .A2(n885bar), .ZN(n922bar);
  OR2_X1 U78 ( .A1(n884), .A2(n883), .ZN(n885) );
  AND2_X1 U78bar ( .A1(n884bar), .A2(n883bar), .ZN(n885bar);
  OR2_X1 U79 ( .A1(n882), .A2(n881), .ZN(n883) );
  AND2_X1 U79bar ( .A1(n882bar), .A2(n881bar), .ZN(n883bar);
  OR2_X1 U80 ( .A1(in[118]), .A2(in[109]), .ZN(n881) );
  AND2_X1 U80bar ( .A1(inbar[118]), .A2(inbar[109]), .ZN(n881bar);
  OR2_X1 U81 ( .A1(in[139]), .A2(in[120]), .ZN(n882) );
  AND2_X1 U81bar ( .A1(inbar[139]), .A2(inbar[120]), .ZN(n882bar);
  OR2_X1 U82 ( .A1(n880), .A2(n879), .ZN(n884) );
  AND2_X1 U82bar ( .A1(n880bar), .A2(n879bar), .ZN(n884bar);
  OR2_X1 U83 ( .A1(in[198]), .A2(in[154]), .ZN(n879) );
  AND2_X1 U83bar ( .A1(inbar[198]), .A2(inbar[154]), .ZN(n879bar);
  OR2_X1 U84 ( .A1(in[210]), .A2(in[205]), .ZN(n880) );
  AND2_X1 U84bar ( .A1(inbar[210]), .A2(inbar[205]), .ZN(n880bar);
  OR2_X1 U85 ( .A1(n878), .A2(n877), .ZN(n886) );
  AND2_X1 U85bar ( .A1(n878bar), .A2(n877bar), .ZN(n886bar);
  OR2_X1 U86 ( .A1(n876), .A2(n875), .ZN(n877) );
  AND2_X1 U86bar ( .A1(n876bar), .A2(n875bar), .ZN(n877bar);
  OR2_X1 U87 ( .A1(in[219]), .A2(in[217]), .ZN(n875) );
  AND2_X1 U87bar ( .A1(inbar[219]), .A2(inbar[217]), .ZN(n875bar);
  OR2_X1 U88 ( .A1(in[86]), .A2(in[252]), .ZN(n876) );
  AND2_X1 U88bar ( .A1(inbar[86]), .A2(inbar[252]), .ZN(n876bar);
  OR2_X1 U89 ( .A1(n874), .A2(n873), .ZN(n878) );
  AND2_X1 U89bar ( .A1(n874bar), .A2(n873bar), .ZN(n878bar);
  OR2_X1 U90 ( .A1(in_40), .A2(in[91]), .ZN(n873) );
  AND2_X1 U90bar ( .A1(in_40bar), .A2(inbar[91]), .ZN(n873bar);
  OR2_X1 U91 ( .A1(in_8), .A2(in_46), .ZN(n874) );
  AND2_X1 U91bar ( .A1(in_8bar), .A2(in_46bar), .ZN(n874bar);
  OR2_X1 U92 ( .A1(n872), .A2(n871), .ZN(n889) );
  AND2_X1 U92bar ( .A1(n872bar), .A2(n871bar), .ZN(n889bar);
  OR2_X1 U93 ( .A1(in[117]), .A2(n943), .ZN(n871) );
  AND2_X1 U93bar ( .A1(inbar[117]), .A2(n943bar), .ZN(n871bar);
  OR2_X1 U94 ( .A1(n870), .A2(n869), .ZN(n943) );
  AND2_X1 U94bar ( .A1(n870bar), .A2(n869bar), .ZN(n943bar);
  OR2_X1 U95 ( .A1(n868), .A2(n867), .ZN(n869) );
  AND2_X1 U95bar ( .A1(n868bar), .A2(n867bar), .ZN(n869bar);
  OR2_X1 U96 ( .A1(n866), .A2(n865), .ZN(n867) );
  AND2_X1 U96bar ( .A1(n866bar), .A2(n865bar), .ZN(n867bar);
  OR2_X1 U97 ( .A1(n864), .A2(n863), .ZN(n865) );
  AND2_X1 U97bar ( .A1(n864bar), .A2(n863bar), .ZN(n865bar);
  OR2_X1 U98 ( .A1(in[108]), .A2(n919), .ZN(n866) );
  AND2_X1 U98bar ( .A1(inbar[108]), .A2(n919bar), .ZN(n866bar);
  OR2_X1 U99 ( .A1(n862), .A2(n861), .ZN(n919) );
  AND2_X1 U99bar ( .A1(n862bar), .A2(n861bar), .ZN(n919bar);
  OR2_X1 U100 ( .A1(n860), .A2(n859), .ZN(n861) );
  AND2_X1 U100bar ( .A1(n860bar), .A2(n859bar), .ZN(n861bar);
  OR2_X1 U101 ( .A1(n858), .A2(n857), .ZN(n859) );
  AND2_X1 U101bar ( .A1(n858bar), .A2(n857bar), .ZN(n859bar);
  OR2_X1 U102 ( .A1(in[119]), .A2(in[105]), .ZN(n857) );
  AND2_X1 U102bar ( .A1(inbar[119]), .A2(inbar[105]), .ZN(n857bar);
  OR2_X1 U103 ( .A1(in[186]), .A2(in[175]), .ZN(n858) );
  AND2_X1 U103bar ( .A1(inbar[186]), .A2(inbar[175]), .ZN(n858bar);
  OR2_X1 U104 ( .A1(n856), .A2(n855), .ZN(n860) );
  AND2_X1 U104bar ( .A1(n856bar), .A2(n855bar), .ZN(n860bar);
  OR2_X1 U105 ( .A1(in[202]), .A2(in[193]), .ZN(n855) );
  AND2_X1 U105bar ( .A1(inbar[202]), .A2(inbar[193]), .ZN(n855bar);
  OR2_X1 U106 ( .A1(in[225]), .A2(in[208]), .ZN(n856) );
  AND2_X1 U106bar ( .A1(inbar[225]), .A2(inbar[208]), .ZN(n856bar);
  OR2_X1 U107 ( .A1(n854), .A2(n853), .ZN(n862) );
  AND2_X1 U107bar ( .A1(n854bar), .A2(n853bar), .ZN(n862bar);
  OR2_X1 U108 ( .A1(n852), .A2(n851), .ZN(n853) );
  AND2_X1 U108bar ( .A1(n852bar), .A2(n851bar), .ZN(n853bar);
  OR2_X1 U109 ( .A1(in_1), .A2(in[85]), .ZN(n851) );
  AND2_X1 U109bar ( .A1(in_1bar), .A2(inbar[85]), .ZN(n851bar);
  OR2_X1 U110 ( .A1(in_23), .A2(in_19), .ZN(n852) );
  AND2_X1 U110bar ( .A1(in_23bar), .A2(in_19bar), .ZN(n852bar);
  OR2_X1 U111 ( .A1(n850), .A2(n849), .ZN(n854) );
  AND2_X1 U111bar ( .A1(n850bar), .A2(n849bar), .ZN(n854bar);
  OR2_X1 U112 ( .A1(in_43), .A2(in_33), .ZN(n849) );
  AND2_X1 U112bar ( .A1(in_43bar), .A2(in_33bar), .ZN(n849bar);
  OR2_X1 U113 ( .A1(in_63), .A2(in_44), .ZN(n850) );
  AND2_X1 U113bar ( .A1(in_63bar), .A2(in_44bar), .ZN(n850bar);
  OR2_X1 U114 ( .A1(n848), .A2(n847), .ZN(n868) );
  AND2_X1 U114bar ( .A1(n848bar), .A2(n847bar), .ZN(n868bar);
  OR2_X1 U115 ( .A1(in[141]), .A2(in[112]), .ZN(n847) );
  AND2_X1 U115bar ( .A1(inbar[141]), .A2(inbar[112]), .ZN(n847bar);
  OR2_X1 U116 ( .A1(in[147]), .A2(n846), .ZN(n848) );
  AND2_X1 U116bar ( .A1(inbar[147]), .A2(n846bar), .ZN(n848bar);
  OR2_X1 U117 ( .A1(in[181]), .A2(in[167]), .ZN(n846) );
  AND2_X1 U117bar ( .A1(inbar[181]), .A2(inbar[167]), .ZN(n846bar);
  OR2_X1 U118 ( .A1(n845), .A2(n844), .ZN(n870) );
  AND2_X1 U118bar ( .A1(n845bar), .A2(n844bar), .ZN(n870bar);
  OR2_X1 U119 ( .A1(n843), .A2(n842), .ZN(n844) );
  AND2_X1 U119bar ( .A1(n843bar), .A2(n842bar), .ZN(n844bar);
  OR2_X1 U120 ( .A1(in[229]), .A2(in[201]), .ZN(n842) );
  AND2_X1 U120bar ( .A1(inbar[229]), .A2(inbar[201]), .ZN(n842bar);
  OR2_X1 U121 ( .A1(in[237]), .A2(n841), .ZN(n843) );
  AND2_X1 U121bar ( .A1(inbar[237]), .A2(n841bar), .ZN(n843bar);
  OR2_X1 U122 ( .A1(in[94]), .A2(in[253]), .ZN(n841) );
  AND2_X1 U122bar ( .A1(inbar[94]), .A2(inbar[253]), .ZN(n841bar);
  OR2_X1 U123 ( .A1(n840), .A2(n839), .ZN(n845) );
  AND2_X1 U123bar ( .A1(n840bar), .A2(n839bar), .ZN(n845bar);
  OR2_X1 U124 ( .A1(in_21), .A2(in[96]), .ZN(n839) );
  AND2_X1 U124bar ( .A1(in_21bar), .A2(inbar[96]), .ZN(n839bar);
  OR2_X1 U125 ( .A1(in_25), .A2(n838), .ZN(n840) );
  AND2_X1 U125bar ( .A1(in_25bar), .A2(n838bar), .ZN(n840bar);
  OR2_X1 U126 ( .A1(in_81), .A2(in_45), .ZN(n838) );
  AND2_X1 U126bar ( .A1(in_81bar), .A2(in_45bar), .ZN(n838bar);
  OR2_X1 U127 ( .A1(n837), .A2(n836), .ZN(n891) );
  AND2_X1 U127bar ( .A1(n837bar), .A2(n836bar), .ZN(n891bar);
  OR2_X1 U128 ( .A1(in[142]), .A2(in[124]), .ZN(n836) );
  AND2_X1 U128bar ( .A1(inbar[142]), .A2(inbar[124]), .ZN(n836bar);
  OR2_X1 U129 ( .A1(in[150]), .A2(n835), .ZN(n837) );
  AND2_X1 U129bar ( .A1(inbar[150]), .A2(n835bar), .ZN(n837bar);
  OR2_X1 U130 ( .A1(in[172]), .A2(in[155]), .ZN(n835) );
  AND2_X1 U130bar ( .A1(inbar[172]), .A2(inbar[155]), .ZN(n835bar);
  OR2_X1 U131 ( .A1(n834), .A2(n833), .ZN(n893) );
  AND2_X1 U131bar ( .A1(n834bar), .A2(n833bar), .ZN(n893bar);
  OR2_X1 U132 ( .A1(n832), .A2(n831), .ZN(n833) );
  AND2_X1 U132bar ( .A1(n832bar), .A2(n831bar), .ZN(n833bar);
  OR2_X1 U133 ( .A1(in[196]), .A2(in[173]), .ZN(n831) );
  AND2_X1 U133bar ( .A1(inbar[196]), .A2(inbar[173]), .ZN(n831bar);
  OR2_X1 U134 ( .A1(in[222]), .A2(n830), .ZN(n832) );
  AND2_X1 U134bar ( .A1(inbar[222]), .A2(n830bar), .ZN(n832bar);
  OR2_X1 U135 ( .A1(in[227]), .A2(in[226]), .ZN(n830) );
  AND2_X1 U135bar ( .A1(inbar[227]), .A2(inbar[226]), .ZN(n830bar);
  OR2_X1 U136 ( .A1(n829), .A2(n828), .ZN(n834) );
  AND2_X1 U136bar ( .A1(n829bar), .A2(n828bar), .ZN(n834bar);
  OR2_X1 U137 ( .A1(in[249]), .A2(in[231]), .ZN(n828) );
  AND2_X1 U137bar ( .A1(inbar[249]), .A2(inbar[231]), .ZN(n828bar);
  OR2_X1 U138 ( .A1(in_28), .A2(n827), .ZN(n829) );
  AND2_X1 U138bar ( .A1(in_28bar), .A2(n827bar), .ZN(n829bar);
  OR2_X1 U139 ( .A1(in_52), .A2(in_47), .ZN(n827) );
  AND2_X1 U139bar ( .A1(in_52bar), .A2(in_47bar), .ZN(n827bar);
  OR2_X1 U140 ( .A1(n826), .A2(n825), .ZN(out[3]) );
  AND2_X1 U140bar ( .A1(n826bar), .A2(n825bar), .ZN(outbar[3]);
  OR2_X1 U141 ( .A1(n824), .A2(n823), .ZN(n825) );
  AND2_X1 U141bar ( .A1(n824bar), .A2(n823bar), .ZN(n825bar);
  OR2_X1 U142 ( .A1(n822), .A2(n821), .ZN(n823) );
  AND2_X1 U142bar ( .A1(n822bar), .A2(n821bar), .ZN(n823bar);
  OR2_X1 U143 ( .A1(n820), .A2(n819), .ZN(n821) );
  AND2_X1 U143bar ( .A1(n820bar), .A2(n819bar), .ZN(n821bar);
  OR2_X1 U144 ( .A1(n964), .A2(n818), .ZN(n822) );
  AND2_X1 U144bar ( .A1(n964bar), .A2(n818bar), .ZN(n822bar);
  OR2_X1 U145 ( .A1(in[118]), .A2(n817), .ZN(n818) );
  AND2_X1 U145bar ( .A1(inbar[118]), .A2(n817bar), .ZN(n818bar);
  OR2_X1 U146 ( .A1(n816), .A2(n815), .ZN(n964) );
  AND2_X1 U146bar ( .A1(n816bar), .A2(n815bar), .ZN(n964bar);
  OR2_X1 U147 ( .A1(n814), .A2(n813), .ZN(n815) );
  AND2_X1 U147bar ( .A1(n814bar), .A2(n813bar), .ZN(n815bar);
  OR2_X1 U148 ( .A1(n812), .A2(n811), .ZN(n813) );
  AND2_X1 U148bar ( .A1(n812bar), .A2(n811bar), .ZN(n813bar);
  OR2_X1 U149 ( .A1(in[122]), .A2(in[111]), .ZN(n811) );
  AND2_X1 U149bar ( .A1(inbar[122]), .A2(inbar[111]), .ZN(n811bar);
  OR2_X1 U150 ( .A1(in[154]), .A2(in[151]), .ZN(n812) );
  AND2_X1 U150bar ( .A1(inbar[154]), .A2(inbar[151]), .ZN(n812bar);
  OR2_X1 U151 ( .A1(n810), .A2(n809), .ZN(n814) );
  AND2_X1 U151bar ( .A1(n810bar), .A2(n809bar), .ZN(n814bar);
  OR2_X1 U152 ( .A1(in[187]), .A2(in[177]), .ZN(n809) );
  AND2_X1 U152bar ( .A1(inbar[187]), .A2(inbar[177]), .ZN(n809bar);
  OR2_X1 U153 ( .A1(in[200]), .A2(in[192]), .ZN(n810) );
  AND2_X1 U153bar ( .A1(inbar[200]), .A2(inbar[192]), .ZN(n810bar);
  OR2_X1 U154 ( .A1(n808), .A2(n807), .ZN(n816) );
  AND2_X1 U154bar ( .A1(n808bar), .A2(n807bar), .ZN(n816bar);
  OR2_X1 U155 ( .A1(n806), .A2(n805), .ZN(n807) );
  AND2_X1 U155bar ( .A1(n806bar), .A2(n805bar), .ZN(n807bar);
  OR2_X1 U156 ( .A1(in[225]), .A2(in[207]), .ZN(n805) );
  AND2_X1 U156bar ( .A1(inbar[225]), .A2(inbar[207]), .ZN(n805bar);
  OR2_X1 U157 ( .A1(in[98]), .A2(in[226]), .ZN(n806) );
  AND2_X1 U157bar ( .A1(inbar[98]), .A2(inbar[226]), .ZN(n806bar);
  OR2_X1 U158 ( .A1(n804), .A2(n803), .ZN(n808) );
  AND2_X1 U158bar ( .A1(n804bar), .A2(n803bar), .ZN(n808bar);
  OR2_X1 U159 ( .A1(in_20), .A2(in_16), .ZN(n803) );
  AND2_X1 U159bar ( .A1(in_20bar), .A2(in_16bar), .ZN(n803bar);
  OR2_X1 U160 ( .A1(in_55), .A2(in_45), .ZN(n804) );
  AND2_X1 U160bar ( .A1(in_55bar), .A2(in_45bar), .ZN(n804bar);
  OR2_X1 U161 ( .A1(n802), .A2(n801), .ZN(n824) );
  AND2_X1 U161bar ( .A1(n802bar), .A2(n801bar), .ZN(n824bar);
  OR2_X1 U162 ( .A1(in[162]), .A2(in[149]), .ZN(n801) );
  AND2_X1 U162bar ( .A1(inbar[162]), .A2(inbar[149]), .ZN(n801bar);
  OR2_X1 U163 ( .A1(in[163]), .A2(n800), .ZN(n802) );
  AND2_X1 U163bar ( .A1(inbar[163]), .A2(n800bar), .ZN(n802bar);
  OR2_X1 U164 ( .A1(in[191]), .A2(in[189]), .ZN(n800) );
  AND2_X1 U164bar ( .A1(inbar[191]), .A2(inbar[189]), .ZN(n800bar);
  OR2_X1 U165 ( .A1(n799), .A2(n798), .ZN(n826) );
  AND2_X1 U165bar ( .A1(n799bar), .A2(n798bar), .ZN(n826bar);
  OR2_X1 U166 ( .A1(n797), .A2(n796), .ZN(n798) );
  AND2_X1 U166bar ( .A1(n797bar), .A2(n796bar), .ZN(n798bar);
  OR2_X1 U167 ( .A1(in[212]), .A2(in[193]), .ZN(n796) );
  AND2_X1 U167bar ( .A1(inbar[212]), .A2(inbar[193]), .ZN(n796bar);
  OR2_X1 U168 ( .A1(in[238]), .A2(n795), .ZN(n797) );
  AND2_X1 U168bar ( .A1(inbar[238]), .A2(n795bar), .ZN(n797bar);
  OR2_X1 U169 ( .A1(in[88]), .A2(in[247]), .ZN(n795) );
  AND2_X1 U169bar ( .A1(inbar[88]), .A2(inbar[247]), .ZN(n795bar);
  OR2_X1 U170 ( .A1(n794), .A2(n793), .ZN(n799) );
  AND2_X1 U170bar ( .A1(n794bar), .A2(n793bar), .ZN(n799bar);
  OR2_X1 U171 ( .A1(in[94]), .A2(in[92]), .ZN(n793) );
  AND2_X1 U171bar ( .A1(inbar[94]), .A2(inbar[92]), .ZN(n793bar);
  OR2_X1 U172 ( .A1(in_52), .A2(n792), .ZN(n794) );
  AND2_X1 U172bar ( .A1(in_52bar), .A2(n792bar), .ZN(n794bar);
  OR2_X1 U173 ( .A1(in_70), .A2(in_67), .ZN(n792) );
  AND2_X1 U173bar ( .A1(in_70bar), .A2(in_67bar), .ZN(n792bar);
  OR2_X1 U174 ( .A1(n791), .A2(n790), .ZN(out[2]) );
  AND2_X1 U174bar ( .A1(n791bar), .A2(n790bar), .ZN(outbar[2]);
  OR2_X1 U175 ( .A1(n789), .A2(n788), .ZN(n790) );
  AND2_X1 U175bar ( .A1(n789bar), .A2(n788bar), .ZN(n790bar);
  OR2_X1 U176 ( .A1(n787), .A2(n786), .ZN(n788) );
  AND2_X1 U176bar ( .A1(n787bar), .A2(n786bar), .ZN(n788bar);
  OR2_X1 U177 ( .A1(n819), .A2(n785), .ZN(n786) );
  AND2_X1 U177bar ( .A1(n819bar), .A2(n785bar), .ZN(n786bar);
  OR2_X1 U178 ( .A1(n784), .A2(n783), .ZN(n819) );
  AND2_X1 U178bar ( .A1(n784bar), .A2(n783bar), .ZN(n819bar);
  OR2_X1 U179 ( .A1(n782), .A2(n781), .ZN(n783) );
  AND2_X1 U179bar ( .A1(n782bar), .A2(n781bar), .ZN(n783bar);
  OR2_X1 U180 ( .A1(n780), .A2(n779), .ZN(n781) );
  AND2_X1 U180bar ( .A1(n780bar), .A2(n779bar), .ZN(n781bar);
  OR2_X1 U181 ( .A1(n962), .A2(n778), .ZN(n779) );
  AND2_X1 U181bar ( .A1(n962bar), .A2(n778bar), .ZN(n779bar);
  OR2_X1 U182 ( .A1(n777), .A2(n776), .ZN(n962) );
  AND2_X1 U182bar ( .A1(n777bar), .A2(n776bar), .ZN(n962bar);
  OR2_X1 U183 ( .A1(n775), .A2(n774), .ZN(n776) );
  AND2_X1 U183bar ( .A1(n775bar), .A2(n774bar), .ZN(n776bar);
  OR2_X1 U184 ( .A1(n773), .A2(n772), .ZN(n774) );
  AND2_X1 U184bar ( .A1(n773bar), .A2(n772bar), .ZN(n774bar);
  OR2_X1 U185 ( .A1(in[131]), .A2(in[120]), .ZN(n772) );
  AND2_X1 U185bar ( .A1(inbar[131]), .A2(inbar[120]), .ZN(n772bar);
  OR2_X1 U186 ( .A1(in[153]), .A2(in[147]), .ZN(n773) );
  AND2_X1 U186bar ( .A1(inbar[153]), .A2(inbar[147]), .ZN(n773bar);
  OR2_X1 U187 ( .A1(n771), .A2(n770), .ZN(n775) );
  AND2_X1 U187bar ( .A1(n771bar), .A2(n770bar), .ZN(n775bar);
  OR2_X1 U188 ( .A1(in[170]), .A2(in[156]), .ZN(n770) );
  AND2_X1 U188bar ( .A1(inbar[170]), .A2(inbar[156]), .ZN(n770bar);
  OR2_X1 U189 ( .A1(in[223]), .A2(in[190]), .ZN(n771) );
  AND2_X1 U189bar ( .A1(inbar[223]), .A2(inbar[190]), .ZN(n771bar);
  OR2_X1 U190 ( .A1(n769), .A2(n768), .ZN(n777) );
  AND2_X1 U190bar ( .A1(n769bar), .A2(n768bar), .ZN(n777bar);
  OR2_X1 U191 ( .A1(n767), .A2(n766), .ZN(n768) );
  AND2_X1 U191bar ( .A1(n767bar), .A2(n766bar), .ZN(n768bar);
  OR2_X1 U192 ( .A1(in[236]), .A2(in[230]), .ZN(n766) );
  AND2_X1 U192bar ( .A1(inbar[236]), .A2(inbar[230]), .ZN(n766bar);
  OR2_X1 U193 ( .A1(in[85]), .A2(in[240]), .ZN(n767) );
  AND2_X1 U193bar ( .A1(inbar[85]), .A2(inbar[240]), .ZN(n767bar);
  OR2_X1 U194 ( .A1(n765), .A2(n764), .ZN(n769) );
  AND2_X1 U194bar ( .A1(n765bar), .A2(n764bar), .ZN(n769bar);
  OR2_X1 U195 ( .A1(in_12), .A2(in[90]), .ZN(n764) );
  AND2_X1 U195bar ( .A1(in_12bar), .A2(inbar[90]), .ZN(n764bar);
  OR2_X1 U196 ( .A1(in_39), .A2(in_28), .ZN(n765) );
  AND2_X1 U196bar ( .A1(in_39bar), .A2(in_28bar), .ZN(n765bar);
  OR2_X1 U197 ( .A1(in[109]), .A2(n763), .ZN(n780) );
  AND2_X1 U197bar ( .A1(inbar[109]), .A2(n763bar), .ZN(n780bar);
  OR2_X1 U198 ( .A1(n762), .A2(n761), .ZN(n782) );
  AND2_X1 U198bar ( .A1(n762bar), .A2(n761bar), .ZN(n782bar);
  OR2_X1 U199 ( .A1(in[138]), .A2(in[129]), .ZN(n761) );
  AND2_X1 U199bar ( .A1(inbar[138]), .A2(inbar[129]), .ZN(n761bar);
  OR2_X1 U200 ( .A1(in[157]), .A2(n760), .ZN(n762) );
  AND2_X1 U200bar ( .A1(inbar[157]), .A2(n760bar), .ZN(n762bar);
  OR2_X1 U201 ( .A1(in[182]), .A2(in[167]), .ZN(n760) );
  AND2_X1 U201bar ( .A1(inbar[182]), .A2(inbar[167]), .ZN(n760bar);
  OR2_X1 U202 ( .A1(n759), .A2(n758), .ZN(n784) );
  AND2_X1 U202bar ( .A1(n759bar), .A2(n758bar), .ZN(n784bar);
  OR2_X1 U203 ( .A1(n757), .A2(n756), .ZN(n758) );
  AND2_X1 U203bar ( .A1(n757bar), .A2(n756bar), .ZN(n758bar);
  OR2_X1 U204 ( .A1(in[195]), .A2(in[184]), .ZN(n756) );
  AND2_X1 U204bar ( .A1(inbar[195]), .A2(inbar[184]), .ZN(n756bar);
  OR2_X1 U205 ( .A1(in[196]), .A2(n755), .ZN(n757) );
  AND2_X1 U205bar ( .A1(inbar[196]), .A2(n755bar), .ZN(n757bar);
  OR2_X1 U206 ( .A1(in[215]), .A2(in[209]), .ZN(n755) );
  AND2_X1 U206bar ( .A1(inbar[215]), .A2(inbar[209]), .ZN(n755bar);
  OR2_X1 U207 ( .A1(n754), .A2(n753), .ZN(n759) );
  AND2_X1 U207bar ( .A1(n754bar), .A2(n753bar), .ZN(n759bar);
  OR2_X1 U208 ( .A1(in[93]), .A2(in[233]), .ZN(n753) );
  AND2_X1 U208bar ( .A1(inbar[93]), .A2(inbar[233]), .ZN(n753bar);
  OR2_X1 U209 ( .A1(in_1), .A2(n752), .ZN(n754) );
  AND2_X1 U209bar ( .A1(in_1bar), .A2(n752bar), .ZN(n754bar);
  OR2_X1 U210 ( .A1(in_69), .A2(in_66), .ZN(n752) );
  AND2_X1 U210bar ( .A1(in_69bar), .A2(in_66bar), .ZN(n752bar);
  OR2_X1 U211 ( .A1(n966), .A2(n751), .ZN(n787) );
  AND2_X1 U211bar ( .A1(n966bar), .A2(n751bar), .ZN(n787bar);
  OR2_X1 U212 ( .A1(in[134]), .A2(n750), .ZN(n751) );
  AND2_X1 U212bar ( .A1(inbar[134]), .A2(n750bar), .ZN(n751bar);
  OR2_X1 U213 ( .A1(n749), .A2(n748), .ZN(n966) );
  AND2_X1 U213bar ( .A1(n749bar), .A2(n748bar), .ZN(n966bar);
  OR2_X1 U214 ( .A1(n747), .A2(n746), .ZN(n748) );
  AND2_X1 U214bar ( .A1(n747bar), .A2(n746bar), .ZN(n748bar);
  OR2_X1 U215 ( .A1(n745), .A2(n744), .ZN(n746) );
  AND2_X1 U215bar ( .A1(n745bar), .A2(n744bar), .ZN(n746bar);
  OR2_X1 U216 ( .A1(in[136]), .A2(in[121]), .ZN(n744) );
  AND2_X1 U216bar ( .A1(inbar[136]), .A2(inbar[121]), .ZN(n744bar);
  OR2_X1 U217 ( .A1(in[186]), .A2(in[174]), .ZN(n745) );
  AND2_X1 U217bar ( .A1(inbar[186]), .A2(inbar[174]), .ZN(n745bar);
  OR2_X1 U218 ( .A1(n743), .A2(n742), .ZN(n747) );
  AND2_X1 U218bar ( .A1(n743bar), .A2(n742bar), .ZN(n747bar);
  OR2_X1 U219 ( .A1(in[198]), .A2(in[197]), .ZN(n742) );
  AND2_X1 U219bar ( .A1(inbar[198]), .A2(inbar[197]), .ZN(n742bar);
  OR2_X1 U220 ( .A1(in[214]), .A2(in[199]), .ZN(n743) );
  AND2_X1 U220bar ( .A1(inbar[214]), .A2(inbar[199]), .ZN(n743bar);
  OR2_X1 U221 ( .A1(n741), .A2(n740), .ZN(n749) );
  AND2_X1 U221bar ( .A1(n741bar), .A2(n740bar), .ZN(n749bar);
  OR2_X1 U222 ( .A1(n739), .A2(n738), .ZN(n740) );
  AND2_X1 U222bar ( .A1(n739bar), .A2(n738bar), .ZN(n740bar);
  OR2_X1 U223 ( .A1(in[231]), .A2(in[220]), .ZN(n738) );
  AND2_X1 U223bar ( .A1(inbar[231]), .A2(inbar[220]), .ZN(n738bar);
  OR2_X1 U224 ( .A1(in_25), .A2(in[245]), .ZN(n739) );
  AND2_X1 U224bar ( .A1(in_25bar), .A2(inbar[245]), .ZN(n739bar);
  OR2_X1 U225 ( .A1(n737), .A2(n736), .ZN(n741) );
  AND2_X1 U225bar ( .A1(n737bar), .A2(n736bar), .ZN(n741bar);
  OR2_X1 U226 ( .A1(in_53), .A2(in_29), .ZN(n736) );
  AND2_X1 U226bar ( .A1(in_53bar), .A2(in_29bar), .ZN(n736bar);
  OR2_X1 U227 ( .A1(in_79), .A2(in_74), .ZN(n737) );
  AND2_X1 U227bar ( .A1(in_79bar), .A2(in_74bar), .ZN(n737bar);
  OR2_X1 U228 ( .A1(n735), .A2(n734), .ZN(n789) );
  AND2_X1 U228bar ( .A1(n735bar), .A2(n734bar), .ZN(n789bar);
  OR2_X1 U229 ( .A1(in[152]), .A2(in[140]), .ZN(n734) );
  AND2_X1 U229bar ( .A1(inbar[152]), .A2(inbar[140]), .ZN(n734bar);
  OR2_X1 U230 ( .A1(in[155]), .A2(n733), .ZN(n735) );
  AND2_X1 U230bar ( .A1(inbar[155]), .A2(n733bar), .ZN(n735bar);
  OR2_X1 U231 ( .A1(in[166]), .A2(in[165]), .ZN(n733) );
  AND2_X1 U231bar ( .A1(inbar[166]), .A2(inbar[165]), .ZN(n733bar);
  OR2_X1 U232 ( .A1(n732), .A2(n731), .ZN(n791) );
  AND2_X1 U232bar ( .A1(n732bar), .A2(n731bar), .ZN(n791bar);
  OR2_X1 U233 ( .A1(n730), .A2(n729), .ZN(n731) );
  AND2_X1 U233bar ( .A1(n730bar), .A2(n729bar), .ZN(n731bar);
  OR2_X1 U234 ( .A1(in[202]), .A2(in[185]), .ZN(n729) );
  AND2_X1 U234bar ( .A1(inbar[202]), .A2(inbar[185]), .ZN(n729bar);
  OR2_X1 U235 ( .A1(in[211]), .A2(n728), .ZN(n730) );
  AND2_X1 U235bar ( .A1(inbar[211]), .A2(n728bar), .ZN(n730bar);
  OR2_X1 U236 ( .A1(in[255]), .A2(in[253]), .ZN(n728) );
  AND2_X1 U236bar ( .A1(inbar[255]), .A2(inbar[253]), .ZN(n728bar);
  OR2_X1 U237 ( .A1(n727), .A2(n726), .ZN(n732) );
  AND2_X1 U237bar ( .A1(n727bar), .A2(n726bar), .ZN(n732bar);
  OR2_X1 U238 ( .A1(in_35), .A2(in_15), .ZN(n726) );
  AND2_X1 U238bar ( .A1(in_35bar), .A2(in_15bar), .ZN(n726bar);
  OR2_X1 U239 ( .A1(in_36), .A2(n725), .ZN(n727) );
  AND2_X1 U239bar ( .A1(in_36bar), .A2(n725bar), .ZN(n727bar);
  OR2_X1 U240 ( .A1(in_48), .A2(in_40), .ZN(n725) );
  AND2_X1 U240bar ( .A1(in_48bar), .A2(in_40bar), .ZN(n725bar);
  OR2_X1 U241 ( .A1(n724), .A2(n723), .ZN(out[1]) );
  AND2_X1 U241bar ( .A1(n724bar), .A2(n723bar), .ZN(outbar[1]);
  OR2_X1 U242 ( .A1(n722), .A2(n721), .ZN(n723) );
  AND2_X1 U242bar ( .A1(n722bar), .A2(n721bar), .ZN(n723bar);
  OR2_X1 U243 ( .A1(n720), .A2(n719), .ZN(n721) );
  AND2_X1 U243bar ( .A1(n720bar), .A2(n719bar), .ZN(n721bar);
  OR2_X1 U244 ( .A1(n921), .A2(n887), .ZN(n719) );
  AND2_X1 U244bar ( .A1(n921bar), .A2(n887bar), .ZN(n719bar);
  OR2_X1 U245 ( .A1(n718), .A2(n717), .ZN(n887) );
  AND2_X1 U245bar ( .A1(n718bar), .A2(n717bar), .ZN(n887bar);
  OR2_X1 U246 ( .A1(n716), .A2(n715), .ZN(n717) );
  AND2_X1 U246bar ( .A1(n716bar), .A2(n715bar), .ZN(n717bar);
  OR2_X1 U247 ( .A1(n714), .A2(n713), .ZN(n715) );
  AND2_X1 U247bar ( .A1(n714bar), .A2(n713bar), .ZN(n715bar);
  OR2_X1 U248 ( .A1(in[116]), .A2(in[110]), .ZN(n713) );
  AND2_X1 U248bar ( .A1(inbar[116]), .A2(inbar[110]), .ZN(n713bar);
  OR2_X1 U249 ( .A1(in[133]), .A2(in[130]), .ZN(n714) );
  AND2_X1 U249bar ( .A1(inbar[133]), .A2(inbar[130]), .ZN(n714bar);
  OR2_X1 U250 ( .A1(n712), .A2(n711), .ZN(n716) );
  AND2_X1 U250bar ( .A1(n712bar), .A2(n711bar), .ZN(n716bar);
  OR2_X1 U251 ( .A1(in[203]), .A2(in[135]), .ZN(n711) );
  AND2_X1 U251bar ( .A1(inbar[203]), .A2(inbar[135]), .ZN(n711bar);
  OR2_X1 U252 ( .A1(in[232]), .A2(in[223]), .ZN(n712) );
  AND2_X1 U252bar ( .A1(inbar[232]), .A2(inbar[223]), .ZN(n712bar);
  OR2_X1 U253 ( .A1(n710), .A2(n709), .ZN(n718) );
  AND2_X1 U253bar ( .A1(n710bar), .A2(n709bar), .ZN(n718bar);
  OR2_X1 U254 ( .A1(n708), .A2(n707), .ZN(n709) );
  AND2_X1 U254bar ( .A1(n708bar), .A2(n707bar), .ZN(n709bar);
  OR2_X1 U255 ( .A1(in[255]), .A2(in[233]), .ZN(n707) );
  AND2_X1 U255bar ( .A1(inbar[255]), .A2(inbar[233]), .ZN(n707bar);
  OR2_X1 U256 ( .A1(in_53), .A2(in_34), .ZN(n708) );
  AND2_X1 U256bar ( .A1(in_53bar), .A2(in_34bar), .ZN(n708bar);
  OR2_X1 U257 ( .A1(n706), .A2(n705), .ZN(n710) );
  AND2_X1 U257bar ( .A1(n706bar), .A2(n705bar), .ZN(n710bar);
  OR2_X1 U258 ( .A1(in_57), .A2(in_55), .ZN(n705) );
  AND2_X1 U258bar ( .A1(in_57bar), .A2(in_55bar), .ZN(n705bar);
  OR2_X1 U259 ( .A1(in_68), .A2(in_67), .ZN(n706) );
  AND2_X1 U259bar ( .A1(in_68bar), .A2(in_67bar), .ZN(n706bar);
  OR2_X1 U260 ( .A1(n704), .A2(n703), .ZN(n921) );
  AND2_X1 U260bar ( .A1(n704bar), .A2(n703bar), .ZN(n921bar);
  OR2_X1 U261 ( .A1(n702), .A2(n701), .ZN(n703) );
  AND2_X1 U261bar ( .A1(n702bar), .A2(n701bar), .ZN(n703bar);
  OR2_X1 U262 ( .A1(n700), .A2(n699), .ZN(n701) );
  AND2_X1 U262bar ( .A1(n700bar), .A2(n699bar), .ZN(n701bar);
  OR2_X1 U263 ( .A1(n944), .A2(n872), .ZN(n699) );
  AND2_X1 U263bar ( .A1(n944bar), .A2(n872bar), .ZN(n699bar);
  OR2_X1 U264 ( .A1(n698), .A2(n697), .ZN(n872) );
  AND2_X1 U264bar ( .A1(n698bar), .A2(n697bar), .ZN(n872bar);
  OR2_X1 U265 ( .A1(n696), .A2(n695), .ZN(n697) );
  AND2_X1 U265bar ( .A1(n696bar), .A2(n695bar), .ZN(n697bar);
  OR2_X1 U266 ( .A1(n694), .A2(n693), .ZN(n695) );
  AND2_X1 U266bar ( .A1(n694bar), .A2(n693bar), .ZN(n695bar);
  OR2_X1 U267 ( .A1(in[121]), .A2(in[102]), .ZN(n693) );
  AND2_X1 U267bar ( .A1(inbar[121]), .A2(inbar[102]), .ZN(n693bar);
  OR2_X1 U268 ( .A1(in[162]), .A2(in[161]), .ZN(n694) );
  AND2_X1 U268bar ( .A1(inbar[162]), .A2(inbar[161]), .ZN(n694bar);
  OR2_X1 U269 ( .A1(n692), .A2(n691), .ZN(n696) );
  AND2_X1 U269bar ( .A1(n692bar), .A2(n691bar), .ZN(n696bar);
  OR2_X1 U270 ( .A1(in[192]), .A2(in[178]), .ZN(n691) );
  AND2_X1 U270bar ( .A1(inbar[192]), .A2(inbar[178]), .ZN(n691bar);
  OR2_X1 U271 ( .A1(in[244]), .A2(in[209]), .ZN(n692) );
  AND2_X1 U271bar ( .A1(inbar[244]), .A2(inbar[209]), .ZN(n692bar);
  OR2_X1 U272 ( .A1(n690), .A2(n689), .ZN(n698) );
  AND2_X1 U272bar ( .A1(n690bar), .A2(n689bar), .ZN(n698bar);
  OR2_X1 U273 ( .A1(n688), .A2(n687), .ZN(n689) );
  AND2_X1 U273bar ( .A1(n688bar), .A2(n687bar), .ZN(n689bar);
  OR2_X1 U274 ( .A1(in[90]), .A2(in[254]), .ZN(n687) );
  AND2_X1 U274bar ( .A1(inbar[90]), .A2(inbar[254]), .ZN(n687bar);
  OR2_X1 U275 ( .A1(in_36), .A2(in_32), .ZN(n688) );
  AND2_X1 U275bar ( .A1(in_36bar), .A2(in_32bar), .ZN(n688bar);
  OR2_X1 U276 ( .A1(n686), .A2(n685), .ZN(n690) );
  AND2_X1 U276bar ( .A1(n686bar), .A2(n685bar), .ZN(n690bar);
  OR2_X1 U277 ( .A1(in_62), .A2(in_37), .ZN(n685) );
  AND2_X1 U277bar ( .A1(in_62bar), .A2(in_37bar), .ZN(n685bar);
  OR2_X1 U278 ( .A1(in_75), .A2(in_73), .ZN(n686) );
  AND2_X1 U278bar ( .A1(in_75bar), .A2(in_73bar), .ZN(n686bar);
  OR2_X1 U279 ( .A1(n684), .A2(n683), .ZN(n944) );
  AND2_X1 U279bar ( .A1(n684bar), .A2(n683bar), .ZN(n944bar);
  OR2_X1 U280 ( .A1(n682), .A2(n681), .ZN(n683) );
  AND2_X1 U280bar ( .A1(n682bar), .A2(n681bar), .ZN(n683bar);
  OR2_X1 U281 ( .A1(n680), .A2(n679), .ZN(n681) );
  AND2_X1 U281bar ( .A1(n680bar), .A2(n679bar), .ZN(n681bar);
  OR2_X1 U282 ( .A1(in[171]), .A2(in[153]), .ZN(n679) );
  AND2_X1 U282bar ( .A1(inbar[171]), .A2(inbar[153]), .ZN(n679bar);
  OR2_X1 U283 ( .A1(in[187]), .A2(in[176]), .ZN(n680) );
  AND2_X1 U283bar ( .A1(inbar[187]), .A2(inbar[176]), .ZN(n680bar);
  OR2_X1 U284 ( .A1(n678), .A2(n677), .ZN(n682) );
  AND2_X1 U284bar ( .A1(n678bar), .A2(n677bar), .ZN(n682bar);
  OR2_X1 U285 ( .A1(in[245]), .A2(in[211]), .ZN(n677) );
  AND2_X1 U285bar ( .A1(inbar[245]), .A2(inbar[211]), .ZN(n677bar);
  OR2_X1 U286 ( .A1(in[97]), .A2(in[88]), .ZN(n678) );
  AND2_X1 U286bar ( .A1(inbar[97]), .A2(inbar[88]), .ZN(n678bar);
  OR2_X1 U287 ( .A1(n676), .A2(n675), .ZN(n684) );
  AND2_X1 U287bar ( .A1(n676bar), .A2(n675bar), .ZN(n684bar);
  OR2_X1 U288 ( .A1(n674), .A2(n673), .ZN(n675) );
  AND2_X1 U288bar ( .A1(n674bar), .A2(n673bar), .ZN(n675bar);
  OR2_X1 U289 ( .A1(in_10), .A2(in_0), .ZN(n673) );
  AND2_X1 U289bar ( .A1(in_10bar), .A2(in_0bar), .ZN(n673bar);
  OR2_X1 U290 ( .A1(in_59), .A2(in_5), .ZN(n674) );
  AND2_X1 U290bar ( .A1(in_59bar), .A2(in_5bar), .ZN(n674bar);
  OR2_X1 U291 ( .A1(n672), .A2(n671), .ZN(n676) );
  AND2_X1 U291bar ( .A1(n672bar), .A2(n671bar), .ZN(n676bar);
  OR2_X1 U292 ( .A1(in_60), .A2(in_6), .ZN(n671) );
  AND2_X1 U292bar ( .A1(in_60bar), .A2(in_6bar), .ZN(n671bar);
  OR2_X1 U293 ( .A1(in_77), .A2(in_69), .ZN(n672) );
  AND2_X1 U293bar ( .A1(in_77bar), .A2(in_69bar), .ZN(n672bar);
  OR2_X1 U294 ( .A1(in[113]), .A2(n864), .ZN(n700) );
  AND2_X1 U294bar ( .A1(inbar[113]), .A2(n864bar), .ZN(n700bar);
  OR2_X1 U295 ( .A1(n670), .A2(n669), .ZN(n864) );
  AND2_X1 U295bar ( .A1(n670bar), .A2(n669bar), .ZN(n864bar);
  OR2_X1 U296 ( .A1(n668), .A2(n667), .ZN(n669) );
  AND2_X1 U296bar ( .A1(n668bar), .A2(n667bar), .ZN(n669bar);
  OR2_X1 U297 ( .A1(n666), .A2(n665), .ZN(n667) );
  AND2_X1 U297bar ( .A1(n666bar), .A2(n665bar), .ZN(n667bar);
  OR2_X1 U298 ( .A1(in[125]), .A2(in[107]), .ZN(n665) );
  AND2_X1 U298bar ( .A1(inbar[125]), .A2(inbar[107]), .ZN(n665bar);
  OR2_X1 U299 ( .A1(in[138]), .A2(in[126]), .ZN(n666) );
  AND2_X1 U299bar ( .A1(inbar[138]), .A2(inbar[126]), .ZN(n666bar);
  OR2_X1 U300 ( .A1(n664), .A2(n663), .ZN(n668) );
  AND2_X1 U300bar ( .A1(n664bar), .A2(n663bar), .ZN(n668bar);
  OR2_X1 U301 ( .A1(in[189]), .A2(in[143]), .ZN(n663) );
  AND2_X1 U301bar ( .A1(inbar[189]), .A2(inbar[143]), .ZN(n663bar);
  OR2_X1 U302 ( .A1(in[99]), .A2(in[214]), .ZN(n664) );
  AND2_X1 U302bar ( .A1(inbar[99]), .A2(inbar[214]), .ZN(n664bar);
  OR2_X1 U303 ( .A1(n662), .A2(n661), .ZN(n670) );
  AND2_X1 U303bar ( .A1(n662bar), .A2(n661bar), .ZN(n670bar);
  OR2_X1 U304 ( .A1(n660), .A2(n659), .ZN(n661) );
  AND2_X1 U304bar ( .A1(n660bar), .A2(n659bar), .ZN(n661bar);
  OR2_X1 U305 ( .A1(in_15), .A2(in_12), .ZN(n659) );
  AND2_X1 U305bar ( .A1(in_15bar), .A2(in_12bar), .ZN(n659bar);
  OR2_X1 U306 ( .A1(in_20), .A2(in_2), .ZN(n660) );
  AND2_X1 U306bar ( .A1(in_20bar), .A2(in_2bar), .ZN(n660bar);
  OR2_X1 U307 ( .A1(n658), .A2(n657), .ZN(n662) );
  AND2_X1 U307bar ( .A1(n658bar), .A2(n657bar), .ZN(n662bar);
  OR2_X1 U308 ( .A1(in_30), .A2(in_3), .ZN(n657) );
  AND2_X1 U308bar ( .A1(in_30bar), .A2(in_3bar), .ZN(n657bar);
  OR2_X1 U309 ( .A1(in_4), .A2(in_38), .ZN(n658) );
  AND2_X1 U309bar ( .A1(in_4bar), .A2(in_38bar), .ZN(n658bar);
  OR2_X1 U310 ( .A1(n656), .A2(n655), .ZN(n702) );
  AND2_X1 U310bar ( .A1(n656bar), .A2(n655bar), .ZN(n702bar);
  OR2_X1 U311 ( .A1(in[148]), .A2(in[137]), .ZN(n655) );
  AND2_X1 U311bar ( .A1(inbar[148]), .A2(inbar[137]), .ZN(n655bar);
  OR2_X1 U312 ( .A1(in[149]), .A2(n654), .ZN(n656) );
  AND2_X1 U312bar ( .A1(inbar[149]), .A2(n654bar), .ZN(n656bar);
  OR2_X1 U313 ( .A1(in[195]), .A2(in[190]), .ZN(n654) );
  AND2_X1 U313bar ( .A1(inbar[195]), .A2(inbar[190]), .ZN(n654bar);
  OR2_X1 U314 ( .A1(n653), .A2(n652), .ZN(n704) );
  AND2_X1 U314bar ( .A1(n653bar), .A2(n652bar), .ZN(n704bar);
  OR2_X1 U315 ( .A1(n651), .A2(n650), .ZN(n652) );
  AND2_X1 U315bar ( .A1(n651bar), .A2(n650bar), .ZN(n652bar);
  OR2_X1 U316 ( .A1(in[98]), .A2(in[197]), .ZN(n650) );
  AND2_X1 U316bar ( .A1(inbar[98]), .A2(inbar[197]), .ZN(n650bar);
  OR2_X1 U317 ( .A1(in_11), .A2(n649), .ZN(n651) );
  AND2_X1 U317bar ( .A1(in_11bar), .A2(n649bar), .ZN(n651bar);
  OR2_X1 U318 ( .A1(in_26), .A2(in_14), .ZN(n649) );
  AND2_X1 U318bar ( .A1(in_26bar), .A2(in_14bar), .ZN(n649bar);
  OR2_X1 U319 ( .A1(n648), .A2(n647), .ZN(n653) );
  AND2_X1 U319bar ( .A1(n648bar), .A2(n647bar), .ZN(n653bar);
  OR2_X1 U320 ( .A1(in_35), .A2(in_27), .ZN(n647) );
  AND2_X1 U320bar ( .A1(in_35bar), .A2(in_27bar), .ZN(n647bar);
  OR2_X1 U321 ( .A1(in_50), .A2(n646), .ZN(n648) );
  AND2_X1 U321bar ( .A1(in_50bar), .A2(n646bar), .ZN(n648bar);
  OR2_X1 U322 ( .A1(in_78), .A2(in_61), .ZN(n646) );
  AND2_X1 U322bar ( .A1(in_78bar), .A2(in_61bar), .ZN(n646bar);
  OR2_X1 U323 ( .A1(n942), .A2(n645), .ZN(n720) );
  AND2_X1 U323bar ( .A1(n942bar), .A2(n645bar), .ZN(n720bar);
  OR2_X1 U324 ( .A1(in[106]), .A2(n863), .ZN(n645) );
  AND2_X1 U324bar ( .A1(inbar[106]), .A2(n863bar), .ZN(n645bar);
  OR2_X1 U325 ( .A1(n644), .A2(n643), .ZN(n863) );
  AND2_X1 U325bar ( .A1(n644bar), .A2(n643bar), .ZN(n863bar);
  OR2_X1 U326 ( .A1(n642), .A2(n641), .ZN(n643) );
  AND2_X1 U326bar ( .A1(n642bar), .A2(n641bar), .ZN(n643bar);
  OR2_X1 U327 ( .A1(n640), .A2(n639), .ZN(n641) );
  AND2_X1 U327bar ( .A1(n640bar), .A2(n639bar), .ZN(n641bar);
  OR2_X1 U328 ( .A1(in[127]), .A2(in[122]), .ZN(n639) );
  AND2_X1 U328bar ( .A1(inbar[127]), .A2(inbar[122]), .ZN(n639bar);
  OR2_X1 U329 ( .A1(in[156]), .A2(in[132]), .ZN(n640) );
  AND2_X1 U329bar ( .A1(inbar[156]), .A2(inbar[132]), .ZN(n640bar);
  OR2_X1 U330 ( .A1(n638), .A2(n637), .ZN(n642) );
  AND2_X1 U330bar ( .A1(n638bar), .A2(n637bar), .ZN(n642bar);
  OR2_X1 U331 ( .A1(in[159]), .A2(in[157]), .ZN(n637) );
  AND2_X1 U331bar ( .A1(inbar[159]), .A2(inbar[157]), .ZN(n637bar);
  OR2_X1 U332 ( .A1(in[185]), .A2(in[169]), .ZN(n638) );
  AND2_X1 U332bar ( .A1(inbar[185]), .A2(inbar[169]), .ZN(n638bar);
  OR2_X1 U333 ( .A1(n636), .A2(n635), .ZN(n644) );
  AND2_X1 U333bar ( .A1(n636bar), .A2(n635bar), .ZN(n644bar);
  OR2_X1 U334 ( .A1(n634), .A2(n633), .ZN(n635) );
  AND2_X1 U334bar ( .A1(n634bar), .A2(n633bar), .ZN(n635bar);
  OR2_X1 U335 ( .A1(in[239]), .A2(in[218]), .ZN(n633) );
  AND2_X1 U335bar ( .A1(inbar[239]), .A2(inbar[218]), .ZN(n633bar);
  OR2_X1 U336 ( .A1(in_13), .A2(in[87]), .ZN(n634) );
  AND2_X1 U336bar ( .A1(in_13bar), .A2(inbar[87]), .ZN(n634bar);
  OR2_X1 U337 ( .A1(n632), .A2(n631), .ZN(n636) );
  AND2_X1 U337bar ( .A1(n632bar), .A2(n631bar), .ZN(n636bar);
  OR2_X1 U338 ( .A1(in_72), .A2(in_70), .ZN(n631) );
  AND2_X1 U338bar ( .A1(in_72bar), .A2(in_70bar), .ZN(n631bar);
  OR2_X1 U339 ( .A1(in_80), .A2(in_74), .ZN(n632) );
  AND2_X1 U339bar ( .A1(in_80bar), .A2(in_74bar), .ZN(n632bar);
  OR2_X1 U340 ( .A1(n630), .A2(n629), .ZN(n942) );
  AND2_X1 U340bar ( .A1(n630bar), .A2(n629bar), .ZN(n942bar);
  OR2_X1 U341 ( .A1(n628), .A2(n627), .ZN(n629) );
  AND2_X1 U341bar ( .A1(n628bar), .A2(n627bar), .ZN(n629bar);
  OR2_X1 U342 ( .A1(n626), .A2(n625), .ZN(n627) );
  AND2_X1 U342bar ( .A1(n626bar), .A2(n625bar), .ZN(n627bar);
  OR2_X1 U343 ( .A1(in[146]), .A2(in[100]), .ZN(n625) );
  AND2_X1 U343bar ( .A1(inbar[146]), .A2(inbar[100]), .ZN(n625bar);
  OR2_X1 U344 ( .A1(in[168]), .A2(in[152]), .ZN(n626) );
  AND2_X1 U344bar ( .A1(inbar[168]), .A2(inbar[152]), .ZN(n626bar);
  OR2_X1 U345 ( .A1(n624), .A2(n623), .ZN(n628) );
  AND2_X1 U345bar ( .A1(n624bar), .A2(n623bar), .ZN(n628bar);
  OR2_X1 U346 ( .A1(in[199]), .A2(in[182]), .ZN(n623) );
  AND2_X1 U346bar ( .A1(inbar[199]), .A2(inbar[182]), .ZN(n623bar);
  OR2_X1 U347 ( .A1(in[236]), .A2(in[204]), .ZN(n624) );
  AND2_X1 U347bar ( .A1(inbar[236]), .A2(inbar[204]), .ZN(n624bar);
  OR2_X1 U348 ( .A1(n622), .A2(n621), .ZN(n630) );
  AND2_X1 U348bar ( .A1(n622bar), .A2(n621bar), .ZN(n630bar);
  OR2_X1 U349 ( .A1(n620), .A2(n619), .ZN(n621) );
  AND2_X1 U349bar ( .A1(n620bar), .A2(n619bar), .ZN(n621bar);
  OR2_X1 U350 ( .A1(in[89]), .A2(in[246]), .ZN(n619) );
  AND2_X1 U350bar ( .A1(inbar[89]), .A2(inbar[246]), .ZN(n619bar);
  OR2_X1 U351 ( .A1(in[95]), .A2(in[92]), .ZN(n620) );
  AND2_X1 U351bar ( .A1(inbar[95]), .A2(inbar[92]), .ZN(n620bar);
  OR2_X1 U352 ( .A1(n618), .A2(n617), .ZN(n622) );
  AND2_X1 U352bar ( .A1(n618bar), .A2(n617bar), .ZN(n622bar);
  OR2_X1 U353 ( .A1(in_22), .A2(in_16), .ZN(n617) );
  AND2_X1 U353bar ( .A1(in_22bar), .A2(in_16bar), .ZN(n617bar);
  OR2_X1 U354 ( .A1(in_51), .A2(in_49), .ZN(n618) );
  AND2_X1 U354bar ( .A1(in_51bar), .A2(in_49bar), .ZN(n618bar);
  OR2_X1 U355 ( .A1(n616), .A2(n615), .ZN(n722) );
  AND2_X1 U355bar ( .A1(n616bar), .A2(n615bar), .ZN(n722bar);
  OR2_X1 U356 ( .A1(in[158]), .A2(in[115]), .ZN(n615) );
  AND2_X1 U356bar ( .A1(inbar[158]), .A2(inbar[115]), .ZN(n615bar);
  OR2_X1 U357 ( .A1(in[163]), .A2(n614), .ZN(n616) );
  AND2_X1 U357bar ( .A1(inbar[163]), .A2(n614bar), .ZN(n616bar);
  OR2_X1 U358 ( .A1(in[206]), .A2(in[165]), .ZN(n614) );
  AND2_X1 U358bar ( .A1(inbar[206]), .A2(inbar[165]), .ZN(n614bar);
  OR2_X1 U359 ( .A1(n613), .A2(n612), .ZN(n724) );
  AND2_X1 U359bar ( .A1(n613bar), .A2(n612bar), .ZN(n724bar);
  OR2_X1 U360 ( .A1(n611), .A2(n610), .ZN(n612) );
  AND2_X1 U360bar ( .A1(n611bar), .A2(n610bar), .ZN(n612bar);
  OR2_X1 U361 ( .A1(in[213]), .A2(in[207]), .ZN(n610) );
  AND2_X1 U361bar ( .A1(inbar[213]), .A2(inbar[207]), .ZN(n610bar);
  OR2_X1 U362 ( .A1(in[215]), .A2(n609), .ZN(n611) );
  AND2_X1 U362bar ( .A1(inbar[215]), .A2(n609bar), .ZN(n611bar);
  OR2_X1 U363 ( .A1(in[230]), .A2(in[220]), .ZN(n609) );
  AND2_X1 U363bar ( .A1(inbar[230]), .A2(inbar[220]), .ZN(n609bar);
  OR2_X1 U364 ( .A1(n608), .A2(n607), .ZN(n613) );
  AND2_X1 U364bar ( .A1(n608bar), .A2(n607bar), .ZN(n613bar);
  OR2_X1 U365 ( .A1(in[251]), .A2(in[234]), .ZN(n607) );
  AND2_X1 U365bar ( .A1(inbar[251]), .A2(inbar[234]), .ZN(n607bar);
  OR2_X1 U366 ( .A1(in_17), .A2(n606), .ZN(n608) );
  AND2_X1 U366bar ( .A1(in_17bar), .A2(n606bar), .ZN(n608bar);
  OR2_X1 U367 ( .A1(in_65), .A2(in_56), .ZN(n606) );
  AND2_X1 U367bar ( .A1(in_65bar), .A2(in_56bar), .ZN(n606bar);
  OR2_X1 U368 ( .A1(n605), .A2(n604), .ZN(out[0]) );
  AND2_X1 U368bar ( .A1(n605bar), .A2(n604bar), .ZN(outbar[0]);
  OR2_X1 U369 ( .A1(n603), .A2(n602), .ZN(n604) );
  AND2_X1 U369bar ( .A1(n603bar), .A2(n602bar), .ZN(n604bar);
  OR2_X1 U370 ( .A1(n601), .A2(n600), .ZN(n602) );
  AND2_X1 U370bar ( .A1(n601bar), .A2(n600bar), .ZN(n602bar);
  OR2_X1 U371 ( .A1(n820), .A2(n785), .ZN(n600) );
  AND2_X1 U371bar ( .A1(n820bar), .A2(n785bar), .ZN(n600bar);
  OR2_X1 U372 ( .A1(n599), .A2(n598), .ZN(n785) );
  AND2_X1 U372bar ( .A1(n599bar), .A2(n598bar), .ZN(n785bar);
  OR2_X1 U373 ( .A1(n597), .A2(n596), .ZN(n598) );
  AND2_X1 U373bar ( .A1(n597bar), .A2(n596bar), .ZN(n598bar);
  OR2_X1 U374 ( .A1(n595), .A2(n594), .ZN(n596) );
  AND2_X1 U374bar ( .A1(n595bar), .A2(n594bar), .ZN(n596bar);
  OR2_X1 U375 ( .A1(in[135]), .A2(in[104]), .ZN(n594) );
  AND2_X1 U375bar ( .A1(inbar[135]), .A2(inbar[104]), .ZN(n594bar);
  OR2_X1 U376 ( .A1(in[188]), .A2(in[178]), .ZN(n595) );
  AND2_X1 U376bar ( .A1(inbar[188]), .A2(inbar[178]), .ZN(n595bar);
  OR2_X1 U377 ( .A1(n593), .A2(n592), .ZN(n597) );
  AND2_X1 U377bar ( .A1(n593bar), .A2(n592bar), .ZN(n597bar);
  OR2_X1 U378 ( .A1(in[217]), .A2(in[194]), .ZN(n592) );
  AND2_X1 U378bar ( .A1(inbar[217]), .A2(inbar[194]), .ZN(n592bar);
  OR2_X1 U379 ( .A1(in[237]), .A2(in[218]), .ZN(n593) );
  AND2_X1 U379bar ( .A1(inbar[237]), .A2(inbar[218]), .ZN(n593bar);
  OR2_X1 U380 ( .A1(n591), .A2(n590), .ZN(n599) );
  AND2_X1 U380bar ( .A1(n591bar), .A2(n590bar), .ZN(n599bar);
  OR2_X1 U381 ( .A1(n589), .A2(n588), .ZN(n590) );
  AND2_X1 U381bar ( .A1(n589bar), .A2(n588bar), .ZN(n590bar);
  OR2_X1 U382 ( .A1(in_2), .A2(in_10), .ZN(n588) );
  AND2_X1 U382bar ( .A1(in_2bar), .A2(in_10bar), .ZN(n588bar);
  OR2_X1 U383 ( .A1(in_47), .A2(in_22), .ZN(n589) );
  AND2_X1 U383bar ( .A1(in_47bar), .A2(in_22bar), .ZN(n589bar);
  OR2_X1 U384 ( .A1(n587), .A2(n586), .ZN(n591) );
  AND2_X1 U384bar ( .A1(n587bar), .A2(n586bar), .ZN(n591bar);
  OR2_X1 U385 ( .A1(in_56), .A2(in_54), .ZN(n586) );
  AND2_X1 U385bar ( .A1(in_56bar), .A2(in_54bar), .ZN(n586bar);
  OR2_X1 U386 ( .A1(in_63), .A2(in_61), .ZN(n587) );
  AND2_X1 U386bar ( .A1(in_63bar), .A2(in_61bar), .ZN(n587bar);
  OR2_X1 U387 ( .A1(n585), .A2(n584), .ZN(n820) );
  AND2_X1 U387bar ( .A1(n585bar), .A2(n584bar), .ZN(n820bar);
  OR2_X1 U388 ( .A1(n583), .A2(n582), .ZN(n584) );
  AND2_X1 U388bar ( .A1(n583bar), .A2(n582bar), .ZN(n584bar);
  OR2_X1 U389 ( .A1(n581), .A2(n580), .ZN(n582) );
  AND2_X1 U389bar ( .A1(n581bar), .A2(n580bar), .ZN(n582bar);
  OR2_X1 U390 ( .A1(in[158]), .A2(in[142]), .ZN(n580) );
  AND2_X1 U390bar ( .A1(inbar[158]), .A2(inbar[142]), .ZN(n580bar);
  OR2_X1 U391 ( .A1(in[175]), .A2(in[164]), .ZN(n581) );
  AND2_X1 U391bar ( .A1(inbar[175]), .A2(inbar[164]), .ZN(n581bar);
  OR2_X1 U392 ( .A1(n579), .A2(n578), .ZN(n583) );
  AND2_X1 U392bar ( .A1(n579bar), .A2(n578bar), .ZN(n583bar);
  OR2_X1 U393 ( .A1(in[228]), .A2(in[204]), .ZN(n578) );
  AND2_X1 U393bar ( .A1(inbar[228]), .A2(inbar[204]), .ZN(n578bar);
  OR2_X1 U394 ( .A1(in[91]), .A2(in[87]), .ZN(n579) );
  AND2_X1 U394bar ( .A1(inbar[91]), .A2(inbar[87]), .ZN(n579bar);
  OR2_X1 U395 ( .A1(n577), .A2(n576), .ZN(n585) );
  AND2_X1 U395bar ( .A1(n577bar), .A2(n576bar), .ZN(n585bar);
  OR2_X1 U396 ( .A1(n575), .A2(n574), .ZN(n576) );
  AND2_X1 U396bar ( .A1(n575bar), .A2(n574bar), .ZN(n576bar);
  OR2_X1 U397 ( .A1(in_21), .A2(in_11), .ZN(n574) );
  AND2_X1 U397bar ( .A1(in_21bar), .A2(in_11bar), .ZN(n574bar);
  OR2_X1 U398 ( .A1(in_5), .A2(in_3), .ZN(n575) );
  AND2_X1 U398bar ( .A1(in_5bar), .A2(in_3bar), .ZN(n575bar);
  OR2_X1 U399 ( .A1(n573), .A2(n572), .ZN(n577) );
  AND2_X1 U399bar ( .A1(n573bar), .A2(n572bar), .ZN(n577bar);
  OR2_X1 U400 ( .A1(in_68), .A2(in_64), .ZN(n572) );
  AND2_X1 U400bar ( .A1(in_68bar), .A2(in_64bar), .ZN(n572bar);
  OR2_X1 U401 ( .A1(in_76), .A2(in_73), .ZN(n573) );
  AND2_X1 U401bar ( .A1(in_76bar), .A2(in_73bar), .ZN(n573bar);
  OR2_X1 U402 ( .A1(n778), .A2(n571), .ZN(n601) );
  AND2_X1 U402bar ( .A1(n778bar), .A2(n571bar), .ZN(n601bar);
  OR2_X1 U403 ( .A1(in[100]), .A2(n965), .ZN(n571) );
  AND2_X1 U403bar ( .A1(inbar[100]), .A2(n965bar), .ZN(n571bar);
  OR2_X1 U404 ( .A1(n570), .A2(n569), .ZN(n965) );
  AND2_X1 U404bar ( .A1(n570bar), .A2(n569bar), .ZN(n965bar);
  OR2_X1 U405 ( .A1(n568), .A2(n567), .ZN(n569) );
  AND2_X1 U405bar ( .A1(n568bar), .A2(n567bar), .ZN(n569bar);
  OR2_X1 U406 ( .A1(n566), .A2(n565), .ZN(n567) );
  AND2_X1 U406bar ( .A1(n566bar), .A2(n565bar), .ZN(n567bar);
  OR2_X1 U407 ( .A1(n817), .A2(n750), .ZN(n565) );
  AND2_X1 U407bar ( .A1(n817bar), .A2(n750bar), .ZN(n565bar);
  OR2_X1 U408 ( .A1(n564), .A2(n563), .ZN(n750) );
  AND2_X1 U408bar ( .A1(n564bar), .A2(n563bar), .ZN(n750bar);
  OR2_X1 U409 ( .A1(n562), .A2(n561), .ZN(n563) );
  AND2_X1 U409bar ( .A1(n562bar), .A2(n561bar), .ZN(n563bar);
  OR2_X1 U410 ( .A1(n560), .A2(n559), .ZN(n561) );
  AND2_X1 U410bar ( .A1(n560bar), .A2(n559bar), .ZN(n561bar);
  OR2_X1 U411 ( .A1(in[119]), .A2(in[103]), .ZN(n559) );
  AND2_X1 U411bar ( .A1(inbar[119]), .A2(inbar[103]), .ZN(n559bar);
  OR2_X1 U412 ( .A1(in[137]), .A2(in[133]), .ZN(n560) );
  AND2_X1 U412bar ( .A1(inbar[137]), .A2(inbar[133]), .ZN(n560bar);
  OR2_X1 U413 ( .A1(n558), .A2(n557), .ZN(n562) );
  AND2_X1 U413bar ( .A1(n558bar), .A2(n557bar), .ZN(n562bar);
  OR2_X1 U414 ( .A1(in[176]), .A2(in[173]), .ZN(n557) );
  AND2_X1 U414bar ( .A1(inbar[176]), .A2(inbar[173]), .ZN(n557bar);
  OR2_X1 U415 ( .A1(in[210]), .A2(in[181]), .ZN(n558) );
  AND2_X1 U415bar ( .A1(inbar[210]), .A2(inbar[181]), .ZN(n558bar);
  OR2_X1 U416 ( .A1(n556), .A2(n555), .ZN(n564) );
  AND2_X1 U416bar ( .A1(n556bar), .A2(n555bar), .ZN(n564bar);
  OR2_X1 U417 ( .A1(n554), .A2(n553), .ZN(n555) );
  AND2_X1 U417bar ( .A1(n554bar), .A2(n553bar), .ZN(n555bar);
  OR2_X1 U418 ( .A1(in_13), .A2(in[234]), .ZN(n553) );
  AND2_X1 U418bar ( .A1(in_13bar), .A2(inbar[234]), .ZN(n553bar);
  OR2_X1 U419 ( .A1(in_38), .A2(in_32), .ZN(n554) );
  AND2_X1 U419bar ( .A1(in_38bar), .A2(in_32bar), .ZN(n554bar);
  OR2_X1 U420 ( .A1(n552), .A2(n551), .ZN(n556) );
  AND2_X1 U420bar ( .A1(n552bar), .A2(n551bar), .ZN(n556bar);
  OR2_X1 U421 ( .A1(in_42), .A2(in_41), .ZN(n551) );
  AND2_X1 U421bar ( .A1(in_42bar), .A2(in_41bar), .ZN(n551bar);
  OR2_X1 U422 ( .A1(in_7), .A2(in_49), .ZN(n552) );
  AND2_X1 U422bar ( .A1(in_7bar), .A2(in_49bar), .ZN(n552bar);
  OR2_X1 U423 ( .A1(n550), .A2(n549), .ZN(n817) );
  AND2_X1 U423bar ( .A1(n550bar), .A2(n549bar), .ZN(n817bar);
  OR2_X1 U424 ( .A1(n548), .A2(n547), .ZN(n549) );
  AND2_X1 U424bar ( .A1(n548bar), .A2(n547bar), .ZN(n549bar);
  OR2_X1 U425 ( .A1(n546), .A2(n545), .ZN(n547) );
  AND2_X1 U425bar ( .A1(n546bar), .A2(n545bar), .ZN(n547bar);
  OR2_X1 U426 ( .A1(in[159]), .A2(in[105]), .ZN(n545) );
  AND2_X1 U426bar ( .A1(inbar[159]), .A2(inbar[105]), .ZN(n545bar);
  OR2_X1 U427 ( .A1(in[206]), .A2(in[183]), .ZN(n546) );
  AND2_X1 U427bar ( .A1(inbar[206]), .A2(inbar[183]), .ZN(n546bar);
  OR2_X1 U428 ( .A1(n544), .A2(n543), .ZN(n548) );
  AND2_X1 U428bar ( .A1(n544bar), .A2(n543bar), .ZN(n548bar);
  OR2_X1 U429 ( .A1(in[229]), .A2(in[219]), .ZN(n543) );
  AND2_X1 U429bar ( .A1(inbar[229]), .A2(inbar[219]), .ZN(n543bar);
  OR2_X1 U430 ( .A1(in[235]), .A2(in[232]), .ZN(n544) );
  AND2_X1 U430bar ( .A1(inbar[235]), .A2(inbar[232]), .ZN(n544bar);
  OR2_X1 U431 ( .A1(n542), .A2(n541), .ZN(n550) );
  AND2_X1 U431bar ( .A1(n542bar), .A2(n541bar), .ZN(n550bar);
  OR2_X1 U432 ( .A1(n540), .A2(n539), .ZN(n541) );
  AND2_X1 U432bar ( .A1(n540bar), .A2(n539bar), .ZN(n541bar);
  OR2_X1 U433 ( .A1(in[249]), .A2(in[242]), .ZN(n539) );
  AND2_X1 U433bar ( .A1(inbar[249]), .A2(inbar[242]), .ZN(n539bar);
  OR2_X1 U434 ( .A1(in[89]), .A2(in[254]), .ZN(n540) );
  AND2_X1 U434bar ( .A1(inbar[89]), .A2(inbar[254]), .ZN(n540bar);
  OR2_X1 U435 ( .A1(n538), .A2(n537), .ZN(n542) );
  AND2_X1 U435bar ( .A1(n538bar), .A2(n537bar), .ZN(n542bar);
  OR2_X1 U436 ( .A1(in_14), .A2(in[99]), .ZN(n537) );
  AND2_X1 U436bar ( .A1(in_14bar), .A2(inbar[99]), .ZN(n537bar);
  OR2_X1 U437 ( .A1(in_60), .A2(in_18), .ZN(n538) );
  AND2_X1 U437bar ( .A1(in_60bar), .A2(in_18bar), .ZN(n538bar);
  OR2_X1 U438 ( .A1(in[113]), .A2(n763), .ZN(n566) );
  AND2_X1 U438bar ( .A1(inbar[113]), .A2(n763bar), .ZN(n566bar);
  OR2_X1 U439 ( .A1(n536), .A2(n535), .ZN(n763) );
  AND2_X1 U439bar ( .A1(n536bar), .A2(n535bar), .ZN(n763bar);
  OR2_X1 U440 ( .A1(n534), .A2(n533), .ZN(n535) );
  AND2_X1 U440bar ( .A1(n534bar), .A2(n533bar), .ZN(n535bar);
  OR2_X1 U441 ( .A1(n532), .A2(n531), .ZN(n533) );
  AND2_X1 U441bar ( .A1(n532bar), .A2(n531bar), .ZN(n533bar);
  OR2_X1 U442 ( .A1(in[115]), .A2(in[110]), .ZN(n531) );
  AND2_X1 U442bar ( .A1(inbar[115]), .A2(inbar[110]), .ZN(n531bar);
  OR2_X1 U443 ( .A1(in[125]), .A2(in[117]), .ZN(n532) );
  AND2_X1 U443bar ( .A1(inbar[125]), .A2(inbar[117]), .ZN(n532bar);
  OR2_X1 U444 ( .A1(n530), .A2(n529), .ZN(n534) );
  AND2_X1 U444bar ( .A1(n530bar), .A2(n529bar), .ZN(n534bar);
  OR2_X1 U445 ( .A1(in[180]), .A2(in[128]), .ZN(n529) );
  AND2_X1 U445bar ( .A1(inbar[180]), .A2(inbar[128]), .ZN(n529bar);
  OR2_X1 U446 ( .A1(in[205]), .A2(in[201]), .ZN(n530) );
  AND2_X1 U446bar ( .A1(inbar[205]), .A2(inbar[201]), .ZN(n530bar);
  OR2_X1 U447 ( .A1(n528), .A2(n527), .ZN(n536) );
  AND2_X1 U447bar ( .A1(n528bar), .A2(n527bar), .ZN(n536bar);
  OR2_X1 U448 ( .A1(n526), .A2(n525), .ZN(n527) );
  AND2_X1 U448bar ( .A1(n526bar), .A2(n525bar), .ZN(n527bar);
  OR2_X1 U449 ( .A1(in[244]), .A2(in[239]), .ZN(n525) );
  AND2_X1 U449bar ( .A1(inbar[244]), .A2(inbar[239]), .ZN(n525bar);
  OR2_X1 U450 ( .A1(in[95]), .A2(in[83]), .ZN(n526) );
  AND2_X1 U450bar ( .A1(inbar[95]), .A2(inbar[83]), .ZN(n526bar);
  OR2_X1 U451 ( .A1(n524), .A2(n523), .ZN(n528) );
  AND2_X1 U451bar ( .A1(n524bar), .A2(n523bar), .ZN(n528bar);
  OR2_X1 U452 ( .A1(in_24), .A2(in[97]), .ZN(n523) );
  AND2_X1 U452bar ( .A1(in_24bar), .A2(inbar[97]), .ZN(n523bar);
  OR2_X1 U453 ( .A1(in_33), .A2(in_27), .ZN(n524) );
  AND2_X1 U453bar ( .A1(in_33bar), .A2(in_27bar), .ZN(n524bar);
  OR2_X1 U454 ( .A1(n522), .A2(n521), .ZN(n568) );
  AND2_X1 U454bar ( .A1(n522bar), .A2(n521bar), .ZN(n568bar);
  OR2_X1 U455 ( .A1(in[145]), .A2(in[126]), .ZN(n521) );
  AND2_X1 U455bar ( .A1(inbar[145]), .A2(inbar[126]), .ZN(n521bar);
  OR2_X1 U456 ( .A1(in[169]), .A2(n520), .ZN(n522) );
  AND2_X1 U456bar ( .A1(inbar[169]), .A2(n520bar), .ZN(n522bar);
  OR2_X1 U457 ( .A1(in[221]), .A2(in[172]), .ZN(n520) );
  AND2_X1 U457bar ( .A1(inbar[221]), .A2(inbar[172]), .ZN(n520bar);
  OR2_X1 U458 ( .A1(n519), .A2(n518), .ZN(n570) );
  AND2_X1 U458bar ( .A1(n519bar), .A2(n518bar), .ZN(n570bar);
  OR2_X1 U459 ( .A1(n517), .A2(n516), .ZN(n518) );
  AND2_X1 U459bar ( .A1(n517bar), .A2(n516bar), .ZN(n518bar);
  OR2_X1 U460 ( .A1(in[241]), .A2(in[224]), .ZN(n516) );
  AND2_X1 U460bar ( .A1(inbar[241]), .A2(inbar[224]), .ZN(n516bar);
  OR2_X1 U461 ( .A1(in[86]), .A2(n515), .ZN(n517) );
  AND2_X1 U461bar ( .A1(inbar[86]), .A2(n515bar), .ZN(n517bar);
  OR2_X1 U462 ( .A1(in_43), .A2(in_34), .ZN(n515) );
  AND2_X1 U462bar ( .A1(in_43bar), .A2(in_34bar), .ZN(n515bar);
  OR2_X1 U463 ( .A1(n514), .A2(n513), .ZN(n519) );
  AND2_X1 U463bar ( .A1(n514bar), .A2(n513bar), .ZN(n519bar);
  OR2_X1 U464 ( .A1(in_65), .A2(in_51), .ZN(n513) );
  AND2_X1 U464bar ( .A1(in_65bar), .A2(in_51bar), .ZN(n513bar);
  OR2_X1 U465 ( .A1(in_75), .A2(n512), .ZN(n514) );
  AND2_X1 U465bar ( .A1(in_75bar), .A2(n512bar), .ZN(n514bar);
  OR2_X1 U466 ( .A1(in_81), .A2(in_77), .ZN(n512) );
  AND2_X1 U466bar ( .A1(in_81bar), .A2(in_77bar), .ZN(n512bar);
  OR2_X1 U467 ( .A1(n511), .A2(n510), .ZN(n778) );
  AND2_X1 U467bar ( .A1(n511bar), .A2(n510bar), .ZN(n778bar);
  OR2_X1 U468 ( .A1(n509), .A2(n508), .ZN(n510) );
  AND2_X1 U468bar ( .A1(n509bar), .A2(n508bar), .ZN(n510bar);
  OR2_X1 U469 ( .A1(n507), .A2(n506), .ZN(n508) );
  AND2_X1 U469bar ( .A1(n507bar), .A2(n506bar), .ZN(n508bar);
  OR2_X1 U470 ( .A1(in[107]), .A2(in[101]), .ZN(n506) );
  AND2_X1 U470bar ( .A1(inbar[107]), .A2(inbar[101]), .ZN(n506bar);
  OR2_X1 U471 ( .A1(in[139]), .A2(in[132]), .ZN(n507) );
  AND2_X1 U471bar ( .A1(inbar[139]), .A2(inbar[132]), .ZN(n507bar);
  OR2_X1 U472 ( .A1(n505), .A2(n504), .ZN(n509) );
  AND2_X1 U472bar ( .A1(n505bar), .A2(n504bar), .ZN(n509bar);
  OR2_X1 U473 ( .A1(in[146]), .A2(in[141]), .ZN(n504) );
  AND2_X1 U473bar ( .A1(inbar[146]), .A2(inbar[141]), .ZN(n504bar);
  OR2_X1 U474 ( .A1(in[203]), .A2(in[179]), .ZN(n505) );
  AND2_X1 U474bar ( .A1(inbar[203]), .A2(inbar[179]), .ZN(n505bar);
  OR2_X1 U475 ( .A1(n503), .A2(n502), .ZN(n511) );
  AND2_X1 U475bar ( .A1(n503bar), .A2(n502bar), .ZN(n511bar);
  OR2_X1 U476 ( .A1(n501), .A2(n500), .ZN(n502) );
  AND2_X1 U476bar ( .A1(n501bar), .A2(n500bar), .ZN(n502bar);
  OR2_X1 U477 ( .A1(in[243]), .A2(in[222]), .ZN(n500) );
  AND2_X1 U477bar ( .A1(inbar[243]), .A2(inbar[222]), .ZN(n500bar);
  OR2_X1 U478 ( .A1(in[251]), .A2(in[250]), .ZN(n501) );
  AND2_X1 U478bar ( .A1(inbar[251]), .A2(inbar[250]), .ZN(n501bar);
  OR2_X1 U479 ( .A1(n499), .A2(n498), .ZN(n503) );
  AND2_X1 U479bar ( .A1(n499bar), .A2(n498bar), .ZN(n503bar);
  OR2_X1 U480 ( .A1(in_37), .A2(in_19), .ZN(n498) );
  AND2_X1 U480bar ( .A1(in_37bar), .A2(in_19bar), .ZN(n498bar);
  OR2_X1 U481 ( .A1(in_78), .A2(in_6), .ZN(n499) );
  AND2_X1 U481bar ( .A1(in_78bar), .A2(in_6bar), .ZN(n499bar);
  OR2_X1 U482 ( .A1(n497), .A2(n496), .ZN(n603) );
  AND2_X1 U482bar ( .A1(n497bar), .A2(n496bar), .ZN(n603bar);
  OR2_X1 U483 ( .A1(in[112]), .A2(in[102]), .ZN(n496) );
  AND2_X1 U483bar ( .A1(inbar[112]), .A2(inbar[102]), .ZN(n496bar);
  OR2_X1 U484 ( .A1(in[123]), .A2(n495), .ZN(n497) );
  AND2_X1 U484bar ( .A1(inbar[123]), .A2(n495bar), .ZN(n497bar);
  OR2_X1 U485 ( .A1(in[143]), .A2(in[130]), .ZN(n495) );
  AND2_X1 U485bar ( .A1(inbar[143]), .A2(inbar[130]), .ZN(n495bar);
  OR2_X1 U486 ( .A1(n494), .A2(n493), .ZN(n605) );
  AND2_X1 U486bar ( .A1(n494bar), .A2(n493bar), .ZN(n605bar);
  OR2_X1 U487 ( .A1(n492), .A2(n491), .ZN(n493) );
  AND2_X1 U487bar ( .A1(n492bar), .A2(n491bar), .ZN(n493bar);
  OR2_X1 U488 ( .A1(in[216]), .A2(in[213]), .ZN(n491) );
  AND2_X1 U488bar ( .A1(inbar[216]), .A2(inbar[213]), .ZN(n491bar);
  OR2_X1 U489 ( .A1(in[227]), .A2(n490), .ZN(n492) );
  AND2_X1 U489bar ( .A1(inbar[227]), .A2(n490bar), .ZN(n492bar);
  OR2_X1 U490 ( .A1(in_0), .A2(in[248]), .ZN(n490) );
  AND2_X1 U490bar ( .A1(in_0bar), .A2(inbar[248]), .ZN(n490bar);
  OR2_X1 U491 ( .A1(n489), .A2(n488), .ZN(n494) );
  AND2_X1 U491bar ( .A1(n489bar), .A2(n488bar), .ZN(n494bar);
  OR2_X1 U492 ( .A1(in_46), .A2(in_44), .ZN(n488) );
  AND2_X1 U492bar ( .A1(in_46bar), .A2(in_44bar), .ZN(n488bar);
  OR2_X1 U493 ( .A1(in_50), .A2(n487), .ZN(n489) );
  AND2_X1 U493bar ( .A1(in_50bar), .A2(n487bar), .ZN(n489bar);
  OR2_X1 U494 ( .A1(in_9), .A2(in_80), .ZN(n487) );
  AND2_X1 U494bar ( .A1(in_9bar), .A2(in_80bar), .ZN(n487bar);
endmodule




module sBox_15 ( in, out );
  input [7:0] in;
  //input_done

  output [7:0] out;
  //output_done

  wire   [255:0] decodeOut;
  //wire_done

  decode_15 dec ( .in(in), .out(decodeOut) );
  encode_15 enc ( .in(decodeOut), .out(out) );
endmodule


module CD2_61 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_62 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_63 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_64 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD4_31 ( a, b, y );
  input [3:0] a;
  input [3:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  //input_done

  output [15:0] y;
  reg [15:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]);
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]);
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]);
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]);
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]);
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]);
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]);
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]);
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]);
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]);
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]);
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]);
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]);
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]);
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]);
endmodule




module CD4_32 ( a, b, y );
  input [3:0] a;
  input [3:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  //input_done

  output [15:0] y;
  reg [15:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]);
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]);
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]);
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]);
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]);
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]);
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]);
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]);
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]);
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]);
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]);
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]);
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]);
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]);
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]);
endmodule




module CD16_16 ( a, b, y );
  input [15:0] a;
  input [15:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign abar[8] = ~a[8];
  assign abar[9] = ~a[9];
  assign abar[10] = ~a[10];
  assign abar[11] = ~a[11];
  assign abar[12] = ~a[12];
  assign abar[13] = ~a[13];
  assign abar[14] = ~a[14];
  assign abar[15] = ~a[15];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign bbar[8] = ~b[8];
  assign bbar[9] = ~b[9];
  assign bbar[10] = ~b[10];
  assign bbar[11] = ~b[11];
  assign bbar[12] = ~b[12];
  assign bbar[13] = ~b[13];
  assign bbar[14] = ~b[14];
  assign bbar[15] = ~b[15];
  //input_done

  output [15:0] y;
  reg [15:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[9]), .A2(a[0]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[9]), .A2(abar[0]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[3]), .A2(a[6]), .ZN(y[99]) );
  OR2_X1 U2bar ( .A1(bbar[3]), .A2(abar[6]), .ZN(ybar[99]);
  AND2_X1 U3 ( .A1(b[2]), .A2(a[6]), .ZN(y[98]) );
  OR2_X1 U3bar ( .A1(bbar[2]), .A2(abar[6]), .ZN(ybar[98]);
  AND2_X1 U4 ( .A1(b[1]), .A2(a[6]), .ZN(y[97]) );
  OR2_X1 U4bar ( .A1(bbar[1]), .A2(abar[6]), .ZN(ybar[97]);
  AND2_X1 U5 ( .A1(b[0]), .A2(a[6]), .ZN(y[96]) );
  OR2_X1 U5bar ( .A1(bbar[0]), .A2(abar[6]), .ZN(ybar[96]);
  AND2_X1 U6 ( .A1(b[15]), .A2(a[5]), .ZN(y[95]) );
  OR2_X1 U6bar ( .A1(bbar[15]), .A2(abar[5]), .ZN(ybar[95]);
  AND2_X1 U7 ( .A1(b[14]), .A2(a[5]), .ZN(y[94]) );
  OR2_X1 U7bar ( .A1(bbar[14]), .A2(abar[5]), .ZN(ybar[94]);
  AND2_X1 U8 ( .A1(b[13]), .A2(a[5]), .ZN(y[93]) );
  OR2_X1 U8bar ( .A1(bbar[13]), .A2(abar[5]), .ZN(ybar[93]);
  AND2_X1 U9 ( .A1(b[12]), .A2(a[5]), .ZN(y[92]) );
  OR2_X1 U9bar ( .A1(bbar[12]), .A2(abar[5]), .ZN(ybar[92]);
  AND2_X1 U10 ( .A1(b[11]), .A2(a[5]), .ZN(y[91]) );
  OR2_X1 U10bar ( .A1(bbar[11]), .A2(abar[5]), .ZN(ybar[91]);
  AND2_X1 U11 ( .A1(b[10]), .A2(a[5]), .ZN(y[90]) );
  OR2_X1 U11bar ( .A1(bbar[10]), .A2(abar[5]), .ZN(ybar[90]);
  AND2_X1 U12 ( .A1(b[8]), .A2(a[0]), .ZN(y[8]) );
  OR2_X1 U12bar ( .A1(bbar[8]), .A2(abar[0]), .ZN(ybar[8]);
  AND2_X1 U13 ( .A1(a[5]), .A2(b[9]), .ZN(y[89]) );
  OR2_X1 U13bar ( .A1(abar[5]), .A2(bbar[9]), .ZN(ybar[89]);
  AND2_X1 U14 ( .A1(b[8]), .A2(a[5]), .ZN(y[88]) );
  OR2_X1 U14bar ( .A1(bbar[8]), .A2(abar[5]), .ZN(ybar[88]);
  AND2_X1 U15 ( .A1(b[7]), .A2(a[5]), .ZN(y[87]) );
  OR2_X1 U15bar ( .A1(bbar[7]), .A2(abar[5]), .ZN(ybar[87]);
  AND2_X1 U16 ( .A1(b[6]), .A2(a[5]), .ZN(y[86]) );
  OR2_X1 U16bar ( .A1(bbar[6]), .A2(abar[5]), .ZN(ybar[86]);
  AND2_X1 U17 ( .A1(b[5]), .A2(a[5]), .ZN(y[85]) );
  OR2_X1 U17bar ( .A1(bbar[5]), .A2(abar[5]), .ZN(ybar[85]);
  AND2_X1 U18 ( .A1(b[4]), .A2(a[5]), .ZN(y[84]) );
  OR2_X1 U18bar ( .A1(bbar[4]), .A2(abar[5]), .ZN(ybar[84]);
  AND2_X1 U19 ( .A1(a[5]), .A2(b[3]), .ZN(y[83]) );
  OR2_X1 U19bar ( .A1(abar[5]), .A2(bbar[3]), .ZN(ybar[83]);
  AND2_X1 U20 ( .A1(a[5]), .A2(b[2]), .ZN(y[82]) );
  OR2_X1 U20bar ( .A1(abar[5]), .A2(bbar[2]), .ZN(ybar[82]);
  AND2_X1 U21 ( .A1(a[5]), .A2(b[1]), .ZN(y[81]) );
  OR2_X1 U21bar ( .A1(abar[5]), .A2(bbar[1]), .ZN(ybar[81]);
  AND2_X1 U22 ( .A1(a[5]), .A2(b[0]), .ZN(y[80]) );
  OR2_X1 U22bar ( .A1(abar[5]), .A2(bbar[0]), .ZN(ybar[80]);
  AND2_X1 U23 ( .A1(b[7]), .A2(a[0]), .ZN(y[7]) );
  OR2_X1 U23bar ( .A1(bbar[7]), .A2(abar[0]), .ZN(ybar[7]);
  AND2_X1 U24 ( .A1(a[4]), .A2(b[15]), .ZN(y[79]) );
  OR2_X1 U24bar ( .A1(abar[4]), .A2(bbar[15]), .ZN(ybar[79]);
  AND2_X1 U25 ( .A1(a[4]), .A2(b[14]), .ZN(y[78]) );
  OR2_X1 U25bar ( .A1(abar[4]), .A2(bbar[14]), .ZN(ybar[78]);
  AND2_X1 U26 ( .A1(a[4]), .A2(b[13]), .ZN(y[77]) );
  OR2_X1 U26bar ( .A1(abar[4]), .A2(bbar[13]), .ZN(ybar[77]);
  AND2_X1 U27 ( .A1(a[4]), .A2(b[12]), .ZN(y[76]) );
  OR2_X1 U27bar ( .A1(abar[4]), .A2(bbar[12]), .ZN(ybar[76]);
  AND2_X1 U28 ( .A1(a[4]), .A2(b[11]), .ZN(y[75]) );
  OR2_X1 U28bar ( .A1(abar[4]), .A2(bbar[11]), .ZN(ybar[75]);
  AND2_X1 U29 ( .A1(a[4]), .A2(b[10]), .ZN(y[74]) );
  OR2_X1 U29bar ( .A1(abar[4]), .A2(bbar[10]), .ZN(ybar[74]);
  AND2_X1 U30 ( .A1(a[4]), .A2(b[9]), .ZN(y[73]) );
  OR2_X1 U30bar ( .A1(abar[4]), .A2(bbar[9]), .ZN(ybar[73]);
  AND2_X1 U31 ( .A1(a[4]), .A2(b[8]), .ZN(y[72]) );
  OR2_X1 U31bar ( .A1(abar[4]), .A2(bbar[8]), .ZN(ybar[72]);
  AND2_X1 U32 ( .A1(a[4]), .A2(b[7]), .ZN(y[71]) );
  OR2_X1 U32bar ( .A1(abar[4]), .A2(bbar[7]), .ZN(ybar[71]);
  AND2_X1 U33 ( .A1(a[4]), .A2(b[6]), .ZN(y[70]) );
  OR2_X1 U33bar ( .A1(abar[4]), .A2(bbar[6]), .ZN(ybar[70]);
  AND2_X1 U34 ( .A1(b[6]), .A2(a[0]), .ZN(y[6]) );
  OR2_X1 U34bar ( .A1(bbar[6]), .A2(abar[0]), .ZN(ybar[6]);
  AND2_X1 U35 ( .A1(a[4]), .A2(b[5]), .ZN(y[69]) );
  OR2_X1 U35bar ( .A1(abar[4]), .A2(bbar[5]), .ZN(ybar[69]);
  AND2_X1 U36 ( .A1(a[4]), .A2(b[4]), .ZN(y[68]) );
  OR2_X1 U36bar ( .A1(abar[4]), .A2(bbar[4]), .ZN(ybar[68]);
  AND2_X1 U37 ( .A1(a[4]), .A2(b[3]), .ZN(y[67]) );
  OR2_X1 U37bar ( .A1(abar[4]), .A2(bbar[3]), .ZN(ybar[67]);
  AND2_X1 U38 ( .A1(a[4]), .A2(b[2]), .ZN(y[66]) );
  OR2_X1 U38bar ( .A1(abar[4]), .A2(bbar[2]), .ZN(ybar[66]);
  AND2_X1 U39 ( .A1(a[4]), .A2(b[1]), .ZN(y[65]) );
  OR2_X1 U39bar ( .A1(abar[4]), .A2(bbar[1]), .ZN(ybar[65]);
  AND2_X1 U40 ( .A1(a[4]), .A2(b[0]), .ZN(y[64]) );
  OR2_X1 U40bar ( .A1(abar[4]), .A2(bbar[0]), .ZN(ybar[64]);
  AND2_X1 U41 ( .A1(a[3]), .A2(b[15]), .ZN(y[63]) );
  OR2_X1 U41bar ( .A1(abar[3]), .A2(bbar[15]), .ZN(ybar[63]);
  AND2_X1 U42 ( .A1(a[3]), .A2(b[14]), .ZN(y[62]) );
  OR2_X1 U42bar ( .A1(abar[3]), .A2(bbar[14]), .ZN(ybar[62]);
  AND2_X1 U43 ( .A1(a[3]), .A2(b[13]), .ZN(y[61]) );
  OR2_X1 U43bar ( .A1(abar[3]), .A2(bbar[13]), .ZN(ybar[61]);
  AND2_X1 U44 ( .A1(a[3]), .A2(b[12]), .ZN(y[60]) );
  OR2_X1 U44bar ( .A1(abar[3]), .A2(bbar[12]), .ZN(ybar[60]);
  AND2_X1 U45 ( .A1(b[5]), .A2(a[0]), .ZN(y[5]) );
  OR2_X1 U45bar ( .A1(bbar[5]), .A2(abar[0]), .ZN(ybar[5]);
  AND2_X1 U46 ( .A1(a[3]), .A2(b[11]), .ZN(y[59]) );
  OR2_X1 U46bar ( .A1(abar[3]), .A2(bbar[11]), .ZN(ybar[59]);
  AND2_X1 U47 ( .A1(a[3]), .A2(b[10]), .ZN(y[58]) );
  OR2_X1 U47bar ( .A1(abar[3]), .A2(bbar[10]), .ZN(ybar[58]);
  AND2_X1 U48 ( .A1(a[3]), .A2(b[9]), .ZN(y[57]) );
  OR2_X1 U48bar ( .A1(abar[3]), .A2(bbar[9]), .ZN(ybar[57]);
  AND2_X1 U49 ( .A1(a[3]), .A2(b[8]), .ZN(y[56]) );
  OR2_X1 U49bar ( .A1(abar[3]), .A2(bbar[8]), .ZN(ybar[56]);
  AND2_X1 U50 ( .A1(a[3]), .A2(b[7]), .ZN(y[55]) );
  OR2_X1 U50bar ( .A1(abar[3]), .A2(bbar[7]), .ZN(ybar[55]);
  AND2_X1 U51 ( .A1(a[3]), .A2(b[6]), .ZN(y[54]) );
  OR2_X1 U51bar ( .A1(abar[3]), .A2(bbar[6]), .ZN(ybar[54]);
  AND2_X1 U52 ( .A1(a[3]), .A2(b[5]), .ZN(y[53]) );
  OR2_X1 U52bar ( .A1(abar[3]), .A2(bbar[5]), .ZN(ybar[53]);
  AND2_X1 U53 ( .A1(a[3]), .A2(b[4]), .ZN(y[52]) );
  OR2_X1 U53bar ( .A1(abar[3]), .A2(bbar[4]), .ZN(ybar[52]);
  AND2_X1 U54 ( .A1(a[3]), .A2(b[3]), .ZN(y[51]) );
  OR2_X1 U54bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[51]);
  AND2_X1 U55 ( .A1(a[3]), .A2(b[2]), .ZN(y[50]) );
  OR2_X1 U55bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[50]);
  AND2_X1 U56 ( .A1(b[4]), .A2(a[0]), .ZN(y[4]) );
  OR2_X1 U56bar ( .A1(bbar[4]), .A2(abar[0]), .ZN(ybar[4]);
  AND2_X1 U57 ( .A1(a[3]), .A2(b[1]), .ZN(y[49]) );
  OR2_X1 U57bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[49]);
  AND2_X1 U58 ( .A1(a[3]), .A2(b[0]), .ZN(y[48]) );
  OR2_X1 U58bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[48]);
  AND2_X1 U59 ( .A1(a[2]), .A2(b[15]), .ZN(y[47]) );
  OR2_X1 U59bar ( .A1(abar[2]), .A2(bbar[15]), .ZN(ybar[47]);
  AND2_X1 U60 ( .A1(a[2]), .A2(b[14]), .ZN(y[46]) );
  OR2_X1 U60bar ( .A1(abar[2]), .A2(bbar[14]), .ZN(ybar[46]);
  AND2_X1 U61 ( .A1(a[2]), .A2(b[13]), .ZN(y[45]) );
  OR2_X1 U61bar ( .A1(abar[2]), .A2(bbar[13]), .ZN(ybar[45]);
  AND2_X1 U62 ( .A1(a[2]), .A2(b[12]), .ZN(y[44]) );
  OR2_X1 U62bar ( .A1(abar[2]), .A2(bbar[12]), .ZN(ybar[44]);
  AND2_X1 U63 ( .A1(a[2]), .A2(b[11]), .ZN(y[43]) );
  OR2_X1 U63bar ( .A1(abar[2]), .A2(bbar[11]), .ZN(ybar[43]);
  AND2_X1 U64 ( .A1(a[2]), .A2(b[10]), .ZN(y[42]) );
  OR2_X1 U64bar ( .A1(abar[2]), .A2(bbar[10]), .ZN(ybar[42]);
  AND2_X1 U65 ( .A1(a[2]), .A2(b[9]), .ZN(y[41]) );
  OR2_X1 U65bar ( .A1(abar[2]), .A2(bbar[9]), .ZN(ybar[41]);
  AND2_X1 U66 ( .A1(a[2]), .A2(b[8]), .ZN(y[40]) );
  OR2_X1 U66bar ( .A1(abar[2]), .A2(bbar[8]), .ZN(ybar[40]);
  AND2_X1 U67 ( .A1(b[3]), .A2(a[0]), .ZN(y[3]) );
  OR2_X1 U67bar ( .A1(bbar[3]), .A2(abar[0]), .ZN(ybar[3]);
  AND2_X1 U68 ( .A1(a[2]), .A2(b[7]), .ZN(y[39]) );
  OR2_X1 U68bar ( .A1(abar[2]), .A2(bbar[7]), .ZN(ybar[39]);
  AND2_X1 U69 ( .A1(a[2]), .A2(b[6]), .ZN(y[38]) );
  OR2_X1 U69bar ( .A1(abar[2]), .A2(bbar[6]), .ZN(ybar[38]);
  AND2_X1 U70 ( .A1(a[2]), .A2(b[5]), .ZN(y[37]) );
  OR2_X1 U70bar ( .A1(abar[2]), .A2(bbar[5]), .ZN(ybar[37]);
  AND2_X1 U71 ( .A1(a[2]), .A2(b[4]), .ZN(y[36]) );
  OR2_X1 U71bar ( .A1(abar[2]), .A2(bbar[4]), .ZN(ybar[36]);
  AND2_X1 U72 ( .A1(a[2]), .A2(b[3]), .ZN(y[35]) );
  OR2_X1 U72bar ( .A1(abar[2]), .A2(bbar[3]), .ZN(ybar[35]);
  AND2_X1 U73 ( .A1(a[2]), .A2(b[2]), .ZN(y[34]) );
  OR2_X1 U73bar ( .A1(abar[2]), .A2(bbar[2]), .ZN(ybar[34]);
  AND2_X1 U74 ( .A1(a[2]), .A2(b[1]), .ZN(y[33]) );
  OR2_X1 U74bar ( .A1(abar[2]), .A2(bbar[1]), .ZN(ybar[33]);
  AND2_X1 U75 ( .A1(a[2]), .A2(b[0]), .ZN(y[32]) );
  OR2_X1 U75bar ( .A1(abar[2]), .A2(bbar[0]), .ZN(ybar[32]);
  AND2_X1 U76 ( .A1(a[1]), .A2(b[15]), .ZN(y[31]) );
  OR2_X1 U76bar ( .A1(abar[1]), .A2(bbar[15]), .ZN(ybar[31]);
  AND2_X1 U77 ( .A1(a[1]), .A2(b[14]), .ZN(y[30]) );
  OR2_X1 U77bar ( .A1(abar[1]), .A2(bbar[14]), .ZN(ybar[30]);
  AND2_X1 U78 ( .A1(b[2]), .A2(a[0]), .ZN(y[2]) );
  OR2_X1 U78bar ( .A1(bbar[2]), .A2(abar[0]), .ZN(ybar[2]);
  AND2_X1 U79 ( .A1(a[1]), .A2(b[13]), .ZN(y[29]) );
  OR2_X1 U79bar ( .A1(abar[1]), .A2(bbar[13]), .ZN(ybar[29]);
  AND2_X1 U80 ( .A1(a[1]), .A2(b[12]), .ZN(y[28]) );
  OR2_X1 U80bar ( .A1(abar[1]), .A2(bbar[12]), .ZN(ybar[28]);
  AND2_X1 U81 ( .A1(a[1]), .A2(b[11]), .ZN(y[27]) );
  OR2_X1 U81bar ( .A1(abar[1]), .A2(bbar[11]), .ZN(ybar[27]);
  AND2_X1 U82 ( .A1(a[1]), .A2(b[10]), .ZN(y[26]) );
  OR2_X1 U82bar ( .A1(abar[1]), .A2(bbar[10]), .ZN(ybar[26]);
  AND2_X1 U83 ( .A1(a[1]), .A2(b[9]), .ZN(y[25]) );
  OR2_X1 U83bar ( .A1(abar[1]), .A2(bbar[9]), .ZN(ybar[25]);
  AND2_X1 U84 ( .A1(a[15]), .A2(b[15]), .ZN(y[255]) );
  OR2_X1 U84bar ( .A1(abar[15]), .A2(bbar[15]), .ZN(ybar[255]);
  AND2_X1 U85 ( .A1(a[15]), .A2(b[14]), .ZN(y[254]) );
  OR2_X1 U85bar ( .A1(abar[15]), .A2(bbar[14]), .ZN(ybar[254]);
  AND2_X1 U86 ( .A1(a[15]), .A2(b[13]), .ZN(y[253]) );
  OR2_X1 U86bar ( .A1(abar[15]), .A2(bbar[13]), .ZN(ybar[253]);
  AND2_X1 U87 ( .A1(a[15]), .A2(b[12]), .ZN(y[252]) );
  OR2_X1 U87bar ( .A1(abar[15]), .A2(bbar[12]), .ZN(ybar[252]);
  AND2_X1 U88 ( .A1(a[15]), .A2(b[11]), .ZN(y[251]) );
  OR2_X1 U88bar ( .A1(abar[15]), .A2(bbar[11]), .ZN(ybar[251]);
  AND2_X1 U89 ( .A1(a[15]), .A2(b[10]), .ZN(y[250]) );
  OR2_X1 U89bar ( .A1(abar[15]), .A2(bbar[10]), .ZN(ybar[250]);
  AND2_X1 U90 ( .A1(a[1]), .A2(b[8]), .ZN(y[24]) );
  OR2_X1 U90bar ( .A1(abar[1]), .A2(bbar[8]), .ZN(ybar[24]);
  AND2_X1 U91 ( .A1(a[15]), .A2(b[9]), .ZN(y[249]) );
  OR2_X1 U91bar ( .A1(abar[15]), .A2(bbar[9]), .ZN(ybar[249]);
  AND2_X1 U92 ( .A1(a[15]), .A2(b[8]), .ZN(y[248]) );
  OR2_X1 U92bar ( .A1(abar[15]), .A2(bbar[8]), .ZN(ybar[248]);
  AND2_X1 U93 ( .A1(a[15]), .A2(b[7]), .ZN(y[247]) );
  OR2_X1 U93bar ( .A1(abar[15]), .A2(bbar[7]), .ZN(ybar[247]);
  AND2_X1 U94 ( .A1(a[15]), .A2(b[6]), .ZN(y[246]) );
  OR2_X1 U94bar ( .A1(abar[15]), .A2(bbar[6]), .ZN(ybar[246]);
  AND2_X1 U95 ( .A1(a[15]), .A2(b[5]), .ZN(y[245]) );
  OR2_X1 U95bar ( .A1(abar[15]), .A2(bbar[5]), .ZN(ybar[245]);
  AND2_X1 U96 ( .A1(a[15]), .A2(b[4]), .ZN(y[244]) );
  OR2_X1 U96bar ( .A1(abar[15]), .A2(bbar[4]), .ZN(ybar[244]);
  AND2_X1 U97 ( .A1(a[15]), .A2(b[3]), .ZN(y[243]) );
  OR2_X1 U97bar ( .A1(abar[15]), .A2(bbar[3]), .ZN(ybar[243]);
  AND2_X1 U98 ( .A1(a[15]), .A2(b[2]), .ZN(y[242]) );
  OR2_X1 U98bar ( .A1(abar[15]), .A2(bbar[2]), .ZN(ybar[242]);
  AND2_X1 U99 ( .A1(a[15]), .A2(b[1]), .ZN(y[241]) );
  OR2_X1 U99bar ( .A1(abar[15]), .A2(bbar[1]), .ZN(ybar[241]);
  AND2_X1 U100 ( .A1(a[15]), .A2(b[0]), .ZN(y[240]) );
  OR2_X1 U100bar ( .A1(abar[15]), .A2(bbar[0]), .ZN(ybar[240]);
  AND2_X1 U101 ( .A1(a[1]), .A2(b[7]), .ZN(y[23]) );
  OR2_X1 U101bar ( .A1(abar[1]), .A2(bbar[7]), .ZN(ybar[23]);
  AND2_X1 U102 ( .A1(a[14]), .A2(b[15]), .ZN(y[239]) );
  OR2_X1 U102bar ( .A1(abar[14]), .A2(bbar[15]), .ZN(ybar[239]);
  AND2_X1 U103 ( .A1(a[14]), .A2(b[14]), .ZN(y[238]) );
  OR2_X1 U103bar ( .A1(abar[14]), .A2(bbar[14]), .ZN(ybar[238]);
  AND2_X1 U104 ( .A1(a[14]), .A2(b[13]), .ZN(y[237]) );
  OR2_X1 U104bar ( .A1(abar[14]), .A2(bbar[13]), .ZN(ybar[237]);
  AND2_X1 U105 ( .A1(a[14]), .A2(b[12]), .ZN(y[236]) );
  OR2_X1 U105bar ( .A1(abar[14]), .A2(bbar[12]), .ZN(ybar[236]);
  AND2_X1 U106 ( .A1(a[14]), .A2(b[11]), .ZN(y[235]) );
  OR2_X1 U106bar ( .A1(abar[14]), .A2(bbar[11]), .ZN(ybar[235]);
  AND2_X1 U107 ( .A1(a[14]), .A2(b[10]), .ZN(y[234]) );
  OR2_X1 U107bar ( .A1(abar[14]), .A2(bbar[10]), .ZN(ybar[234]);
  AND2_X1 U108 ( .A1(a[14]), .A2(b[9]), .ZN(y[233]) );
  OR2_X1 U108bar ( .A1(abar[14]), .A2(bbar[9]), .ZN(ybar[233]);
  AND2_X1 U109 ( .A1(a[14]), .A2(b[8]), .ZN(y[232]) );
  OR2_X1 U109bar ( .A1(abar[14]), .A2(bbar[8]), .ZN(ybar[232]);
  AND2_X1 U110 ( .A1(a[14]), .A2(b[7]), .ZN(y[231]) );
  OR2_X1 U110bar ( .A1(abar[14]), .A2(bbar[7]), .ZN(ybar[231]);
  AND2_X1 U111 ( .A1(a[14]), .A2(b[6]), .ZN(y[230]) );
  OR2_X1 U111bar ( .A1(abar[14]), .A2(bbar[6]), .ZN(ybar[230]);
  AND2_X1 U112 ( .A1(a[1]), .A2(b[6]), .ZN(y[22]) );
  OR2_X1 U112bar ( .A1(abar[1]), .A2(bbar[6]), .ZN(ybar[22]);
  AND2_X1 U113 ( .A1(a[14]), .A2(b[5]), .ZN(y[229]) );
  OR2_X1 U113bar ( .A1(abar[14]), .A2(bbar[5]), .ZN(ybar[229]);
  AND2_X1 U114 ( .A1(a[14]), .A2(b[4]), .ZN(y[228]) );
  OR2_X1 U114bar ( .A1(abar[14]), .A2(bbar[4]), .ZN(ybar[228]);
  AND2_X1 U115 ( .A1(a[14]), .A2(b[3]), .ZN(y[227]) );
  OR2_X1 U115bar ( .A1(abar[14]), .A2(bbar[3]), .ZN(ybar[227]);
  AND2_X1 U116 ( .A1(a[14]), .A2(b[2]), .ZN(y[226]) );
  OR2_X1 U116bar ( .A1(abar[14]), .A2(bbar[2]), .ZN(ybar[226]);
  AND2_X1 U117 ( .A1(a[14]), .A2(b[1]), .ZN(y[225]) );
  OR2_X1 U117bar ( .A1(abar[14]), .A2(bbar[1]), .ZN(ybar[225]);
  AND2_X1 U118 ( .A1(a[14]), .A2(b[0]), .ZN(y[224]) );
  OR2_X1 U118bar ( .A1(abar[14]), .A2(bbar[0]), .ZN(ybar[224]);
  AND2_X1 U119 ( .A1(a[13]), .A2(b[15]), .ZN(y[223]) );
  OR2_X1 U119bar ( .A1(abar[13]), .A2(bbar[15]), .ZN(ybar[223]);
  AND2_X1 U120 ( .A1(a[13]), .A2(b[14]), .ZN(y[222]) );
  OR2_X1 U120bar ( .A1(abar[13]), .A2(bbar[14]), .ZN(ybar[222]);
  AND2_X1 U121 ( .A1(a[13]), .A2(b[13]), .ZN(y[221]) );
  OR2_X1 U121bar ( .A1(abar[13]), .A2(bbar[13]), .ZN(ybar[221]);
  AND2_X1 U122 ( .A1(a[13]), .A2(b[12]), .ZN(y[220]) );
  OR2_X1 U122bar ( .A1(abar[13]), .A2(bbar[12]), .ZN(ybar[220]);
  AND2_X1 U123 ( .A1(a[1]), .A2(b[5]), .ZN(y[21]) );
  OR2_X1 U123bar ( .A1(abar[1]), .A2(bbar[5]), .ZN(ybar[21]);
  AND2_X1 U124 ( .A1(a[13]), .A2(b[11]), .ZN(y[219]) );
  OR2_X1 U124bar ( .A1(abar[13]), .A2(bbar[11]), .ZN(ybar[219]);
  AND2_X1 U125 ( .A1(a[13]), .A2(b[10]), .ZN(y[218]) );
  OR2_X1 U125bar ( .A1(abar[13]), .A2(bbar[10]), .ZN(ybar[218]);
  AND2_X1 U126 ( .A1(a[13]), .A2(b[9]), .ZN(y[217]) );
  OR2_X1 U126bar ( .A1(abar[13]), .A2(bbar[9]), .ZN(ybar[217]);
  AND2_X1 U127 ( .A1(a[13]), .A2(b[8]), .ZN(y[216]) );
  OR2_X1 U127bar ( .A1(abar[13]), .A2(bbar[8]), .ZN(ybar[216]);
  AND2_X1 U128 ( .A1(a[13]), .A2(b[7]), .ZN(y[215]) );
  OR2_X1 U128bar ( .A1(abar[13]), .A2(bbar[7]), .ZN(ybar[215]);
  AND2_X1 U129 ( .A1(a[13]), .A2(b[6]), .ZN(y[214]) );
  OR2_X1 U129bar ( .A1(abar[13]), .A2(bbar[6]), .ZN(ybar[214]);
  AND2_X1 U130 ( .A1(a[13]), .A2(b[5]), .ZN(y[213]) );
  OR2_X1 U130bar ( .A1(abar[13]), .A2(bbar[5]), .ZN(ybar[213]);
  AND2_X1 U131 ( .A1(a[13]), .A2(b[4]), .ZN(y[212]) );
  OR2_X1 U131bar ( .A1(abar[13]), .A2(bbar[4]), .ZN(ybar[212]);
  AND2_X1 U132 ( .A1(a[13]), .A2(b[3]), .ZN(y[211]) );
  OR2_X1 U132bar ( .A1(abar[13]), .A2(bbar[3]), .ZN(ybar[211]);
  AND2_X1 U133 ( .A1(a[13]), .A2(b[2]), .ZN(y[210]) );
  OR2_X1 U133bar ( .A1(abar[13]), .A2(bbar[2]), .ZN(ybar[210]);
  AND2_X1 U134 ( .A1(a[1]), .A2(b[4]), .ZN(y[20]) );
  OR2_X1 U134bar ( .A1(abar[1]), .A2(bbar[4]), .ZN(ybar[20]);
  AND2_X1 U135 ( .A1(a[13]), .A2(b[1]), .ZN(y[209]) );
  OR2_X1 U135bar ( .A1(abar[13]), .A2(bbar[1]), .ZN(ybar[209]);
  AND2_X1 U136 ( .A1(a[13]), .A2(b[0]), .ZN(y[208]) );
  OR2_X1 U136bar ( .A1(abar[13]), .A2(bbar[0]), .ZN(ybar[208]);
  AND2_X1 U137 ( .A1(a[12]), .A2(b[15]), .ZN(y[207]) );
  OR2_X1 U137bar ( .A1(abar[12]), .A2(bbar[15]), .ZN(ybar[207]);
  AND2_X1 U138 ( .A1(a[12]), .A2(b[14]), .ZN(y[206]) );
  OR2_X1 U138bar ( .A1(abar[12]), .A2(bbar[14]), .ZN(ybar[206]);
  AND2_X1 U139 ( .A1(a[12]), .A2(b[13]), .ZN(y[205]) );
  OR2_X1 U139bar ( .A1(abar[12]), .A2(bbar[13]), .ZN(ybar[205]);
  AND2_X1 U140 ( .A1(a[12]), .A2(b[12]), .ZN(y[204]) );
  OR2_X1 U140bar ( .A1(abar[12]), .A2(bbar[12]), .ZN(ybar[204]);
  AND2_X1 U141 ( .A1(a[12]), .A2(b[11]), .ZN(y[203]) );
  OR2_X1 U141bar ( .A1(abar[12]), .A2(bbar[11]), .ZN(ybar[203]);
  AND2_X1 U142 ( .A1(a[12]), .A2(b[10]), .ZN(y[202]) );
  OR2_X1 U142bar ( .A1(abar[12]), .A2(bbar[10]), .ZN(ybar[202]);
  AND2_X1 U143 ( .A1(a[12]), .A2(b[9]), .ZN(y[201]) );
  OR2_X1 U143bar ( .A1(abar[12]), .A2(bbar[9]), .ZN(ybar[201]);
  AND2_X1 U144 ( .A1(a[12]), .A2(b[8]), .ZN(y[200]) );
  OR2_X1 U144bar ( .A1(abar[12]), .A2(bbar[8]), .ZN(ybar[200]);
  AND2_X1 U145 ( .A1(b[1]), .A2(a[0]), .ZN(y[1]) );
  OR2_X1 U145bar ( .A1(bbar[1]), .A2(abar[0]), .ZN(ybar[1]);
  AND2_X1 U146 ( .A1(a[1]), .A2(b[3]), .ZN(y[19]) );
  OR2_X1 U146bar ( .A1(abar[1]), .A2(bbar[3]), .ZN(ybar[19]);
  AND2_X1 U147 ( .A1(a[12]), .A2(b[7]), .ZN(y[199]) );
  OR2_X1 U147bar ( .A1(abar[12]), .A2(bbar[7]), .ZN(ybar[199]);
  AND2_X1 U148 ( .A1(a[12]), .A2(b[6]), .ZN(y[198]) );
  OR2_X1 U148bar ( .A1(abar[12]), .A2(bbar[6]), .ZN(ybar[198]);
  AND2_X1 U149 ( .A1(a[12]), .A2(b[5]), .ZN(y[197]) );
  OR2_X1 U149bar ( .A1(abar[12]), .A2(bbar[5]), .ZN(ybar[197]);
  AND2_X1 U150 ( .A1(a[12]), .A2(b[4]), .ZN(y[196]) );
  OR2_X1 U150bar ( .A1(abar[12]), .A2(bbar[4]), .ZN(ybar[196]);
  AND2_X1 U151 ( .A1(a[12]), .A2(b[3]), .ZN(y[195]) );
  OR2_X1 U151bar ( .A1(abar[12]), .A2(bbar[3]), .ZN(ybar[195]);
  AND2_X1 U152 ( .A1(a[12]), .A2(b[2]), .ZN(y[194]) );
  OR2_X1 U152bar ( .A1(abar[12]), .A2(bbar[2]), .ZN(ybar[194]);
  AND2_X1 U153 ( .A1(a[12]), .A2(b[1]), .ZN(y[193]) );
  OR2_X1 U153bar ( .A1(abar[12]), .A2(bbar[1]), .ZN(ybar[193]);
  AND2_X1 U154 ( .A1(a[12]), .A2(b[0]), .ZN(y[192]) );
  OR2_X1 U154bar ( .A1(abar[12]), .A2(bbar[0]), .ZN(ybar[192]);
  AND2_X1 U155 ( .A1(a[11]), .A2(b[15]), .ZN(y[191]) );
  OR2_X1 U155bar ( .A1(abar[11]), .A2(bbar[15]), .ZN(ybar[191]);
  AND2_X1 U156 ( .A1(a[11]), .A2(b[14]), .ZN(y[190]) );
  OR2_X1 U156bar ( .A1(abar[11]), .A2(bbar[14]), .ZN(ybar[190]);
  AND2_X1 U157 ( .A1(a[1]), .A2(b[2]), .ZN(y[18]) );
  OR2_X1 U157bar ( .A1(abar[1]), .A2(bbar[2]), .ZN(ybar[18]);
  AND2_X1 U158 ( .A1(a[11]), .A2(b[13]), .ZN(y[189]) );
  OR2_X1 U158bar ( .A1(abar[11]), .A2(bbar[13]), .ZN(ybar[189]);
  AND2_X1 U159 ( .A1(a[11]), .A2(b[12]), .ZN(y[188]) );
  OR2_X1 U159bar ( .A1(abar[11]), .A2(bbar[12]), .ZN(ybar[188]);
  AND2_X1 U160 ( .A1(a[11]), .A2(b[11]), .ZN(y[187]) );
  OR2_X1 U160bar ( .A1(abar[11]), .A2(bbar[11]), .ZN(ybar[187]);
  AND2_X1 U161 ( .A1(a[11]), .A2(b[10]), .ZN(y[186]) );
  OR2_X1 U161bar ( .A1(abar[11]), .A2(bbar[10]), .ZN(ybar[186]);
  AND2_X1 U162 ( .A1(a[11]), .A2(b[9]), .ZN(y[185]) );
  OR2_X1 U162bar ( .A1(abar[11]), .A2(bbar[9]), .ZN(ybar[185]);
  AND2_X1 U163 ( .A1(a[11]), .A2(b[8]), .ZN(y[184]) );
  OR2_X1 U163bar ( .A1(abar[11]), .A2(bbar[8]), .ZN(ybar[184]);
  AND2_X1 U164 ( .A1(a[11]), .A2(b[7]), .ZN(y[183]) );
  OR2_X1 U164bar ( .A1(abar[11]), .A2(bbar[7]), .ZN(ybar[183]);
  AND2_X1 U165 ( .A1(a[11]), .A2(b[6]), .ZN(y[182]) );
  OR2_X1 U165bar ( .A1(abar[11]), .A2(bbar[6]), .ZN(ybar[182]);
  AND2_X1 U166 ( .A1(a[11]), .A2(b[5]), .ZN(y[181]) );
  OR2_X1 U166bar ( .A1(abar[11]), .A2(bbar[5]), .ZN(ybar[181]);
  AND2_X1 U167 ( .A1(a[11]), .A2(b[4]), .ZN(y[180]) );
  OR2_X1 U167bar ( .A1(abar[11]), .A2(bbar[4]), .ZN(ybar[180]);
  AND2_X1 U168 ( .A1(a[1]), .A2(b[1]), .ZN(y[17]) );
  OR2_X1 U168bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[17]);
  AND2_X1 U169 ( .A1(a[11]), .A2(b[3]), .ZN(y[179]) );
  OR2_X1 U169bar ( .A1(abar[11]), .A2(bbar[3]), .ZN(ybar[179]);
  AND2_X1 U170 ( .A1(a[11]), .A2(b[2]), .ZN(y[178]) );
  OR2_X1 U170bar ( .A1(abar[11]), .A2(bbar[2]), .ZN(ybar[178]);
  AND2_X1 U171 ( .A1(a[11]), .A2(b[1]), .ZN(y[177]) );
  OR2_X1 U171bar ( .A1(abar[11]), .A2(bbar[1]), .ZN(ybar[177]);
  AND2_X1 U172 ( .A1(a[11]), .A2(b[0]), .ZN(y[176]) );
  OR2_X1 U172bar ( .A1(abar[11]), .A2(bbar[0]), .ZN(ybar[176]);
  AND2_X1 U173 ( .A1(a[10]), .A2(b[15]), .ZN(y[175]) );
  OR2_X1 U173bar ( .A1(abar[10]), .A2(bbar[15]), .ZN(ybar[175]);
  AND2_X1 U174 ( .A1(a[10]), .A2(b[14]), .ZN(y[174]) );
  OR2_X1 U174bar ( .A1(abar[10]), .A2(bbar[14]), .ZN(ybar[174]);
  AND2_X1 U175 ( .A1(a[10]), .A2(b[13]), .ZN(y[173]) );
  OR2_X1 U175bar ( .A1(abar[10]), .A2(bbar[13]), .ZN(ybar[173]);
  AND2_X1 U176 ( .A1(a[10]), .A2(b[12]), .ZN(y[172]) );
  OR2_X1 U176bar ( .A1(abar[10]), .A2(bbar[12]), .ZN(ybar[172]);
  AND2_X1 U177 ( .A1(a[10]), .A2(b[11]), .ZN(y[171]) );
  OR2_X1 U177bar ( .A1(abar[10]), .A2(bbar[11]), .ZN(ybar[171]);
  AND2_X1 U178 ( .A1(a[10]), .A2(b[10]), .ZN(y[170]) );
  OR2_X1 U178bar ( .A1(abar[10]), .A2(bbar[10]), .ZN(ybar[170]);
  AND2_X1 U179 ( .A1(a[1]), .A2(b[0]), .ZN(y[16]) );
  OR2_X1 U179bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[16]);
  AND2_X1 U180 ( .A1(a[10]), .A2(b[9]), .ZN(y[169]) );
  OR2_X1 U180bar ( .A1(abar[10]), .A2(bbar[9]), .ZN(ybar[169]);
  AND2_X1 U181 ( .A1(a[10]), .A2(b[8]), .ZN(y[168]) );
  OR2_X1 U181bar ( .A1(abar[10]), .A2(bbar[8]), .ZN(ybar[168]);
  AND2_X1 U182 ( .A1(a[10]), .A2(b[7]), .ZN(y[167]) );
  OR2_X1 U182bar ( .A1(abar[10]), .A2(bbar[7]), .ZN(ybar[167]);
  AND2_X1 U183 ( .A1(a[10]), .A2(b[6]), .ZN(y[166]) );
  OR2_X1 U183bar ( .A1(abar[10]), .A2(bbar[6]), .ZN(ybar[166]);
  AND2_X1 U184 ( .A1(a[10]), .A2(b[5]), .ZN(y[165]) );
  OR2_X1 U184bar ( .A1(abar[10]), .A2(bbar[5]), .ZN(ybar[165]);
  AND2_X1 U185 ( .A1(a[10]), .A2(b[4]), .ZN(y[164]) );
  OR2_X1 U185bar ( .A1(abar[10]), .A2(bbar[4]), .ZN(ybar[164]);
  AND2_X1 U186 ( .A1(a[10]), .A2(b[3]), .ZN(y[163]) );
  OR2_X1 U186bar ( .A1(abar[10]), .A2(bbar[3]), .ZN(ybar[163]);
  AND2_X1 U187 ( .A1(a[10]), .A2(b[2]), .ZN(y[162]) );
  OR2_X1 U187bar ( .A1(abar[10]), .A2(bbar[2]), .ZN(ybar[162]);
  AND2_X1 U188 ( .A1(a[10]), .A2(b[1]), .ZN(y[161]) );
  OR2_X1 U188bar ( .A1(abar[10]), .A2(bbar[1]), .ZN(ybar[161]);
  AND2_X1 U189 ( .A1(a[10]), .A2(b[0]), .ZN(y[160]) );
  OR2_X1 U189bar ( .A1(abar[10]), .A2(bbar[0]), .ZN(ybar[160]);
  AND2_X1 U190 ( .A1(b[15]), .A2(a[0]), .ZN(y[15]) );
  OR2_X1 U190bar ( .A1(bbar[15]), .A2(abar[0]), .ZN(ybar[15]);
  AND2_X1 U191 ( .A1(a[9]), .A2(b[15]), .ZN(y[159]) );
  OR2_X1 U191bar ( .A1(abar[9]), .A2(bbar[15]), .ZN(ybar[159]);
  AND2_X1 U192 ( .A1(a[9]), .A2(b[14]), .ZN(y[158]) );
  OR2_X1 U192bar ( .A1(abar[9]), .A2(bbar[14]), .ZN(ybar[158]);
  AND2_X1 U193 ( .A1(a[9]), .A2(b[13]), .ZN(y[157]) );
  OR2_X1 U193bar ( .A1(abar[9]), .A2(bbar[13]), .ZN(ybar[157]);
  AND2_X1 U194 ( .A1(a[9]), .A2(b[12]), .ZN(y[156]) );
  OR2_X1 U194bar ( .A1(abar[9]), .A2(bbar[12]), .ZN(ybar[156]);
  AND2_X1 U195 ( .A1(a[9]), .A2(b[11]), .ZN(y[155]) );
  OR2_X1 U195bar ( .A1(abar[9]), .A2(bbar[11]), .ZN(ybar[155]);
  AND2_X1 U196 ( .A1(a[9]), .A2(b[10]), .ZN(y[154]) );
  OR2_X1 U196bar ( .A1(abar[9]), .A2(bbar[10]), .ZN(ybar[154]);
  AND2_X1 U197 ( .A1(a[9]), .A2(b[9]), .ZN(y[153]) );
  OR2_X1 U197bar ( .A1(abar[9]), .A2(bbar[9]), .ZN(ybar[153]);
  AND2_X1 U198 ( .A1(a[9]), .A2(b[8]), .ZN(y[152]) );
  OR2_X1 U198bar ( .A1(abar[9]), .A2(bbar[8]), .ZN(ybar[152]);
  AND2_X1 U199 ( .A1(a[9]), .A2(b[7]), .ZN(y[151]) );
  OR2_X1 U199bar ( .A1(abar[9]), .A2(bbar[7]), .ZN(ybar[151]);
  AND2_X1 U200 ( .A1(a[9]), .A2(b[6]), .ZN(y[150]) );
  OR2_X1 U200bar ( .A1(abar[9]), .A2(bbar[6]), .ZN(ybar[150]);
  AND2_X1 U201 ( .A1(b[14]), .A2(a[0]), .ZN(y[14]) );
  OR2_X1 U201bar ( .A1(bbar[14]), .A2(abar[0]), .ZN(ybar[14]);
  AND2_X1 U202 ( .A1(a[9]), .A2(b[5]), .ZN(y[149]) );
  OR2_X1 U202bar ( .A1(abar[9]), .A2(bbar[5]), .ZN(ybar[149]);
  AND2_X1 U203 ( .A1(a[9]), .A2(b[4]), .ZN(y[148]) );
  OR2_X1 U203bar ( .A1(abar[9]), .A2(bbar[4]), .ZN(ybar[148]);
  AND2_X1 U204 ( .A1(a[9]), .A2(b[3]), .ZN(y[147]) );
  OR2_X1 U204bar ( .A1(abar[9]), .A2(bbar[3]), .ZN(ybar[147]);
  AND2_X1 U205 ( .A1(a[9]), .A2(b[2]), .ZN(y[146]) );
  OR2_X1 U205bar ( .A1(abar[9]), .A2(bbar[2]), .ZN(ybar[146]);
  AND2_X1 U206 ( .A1(a[9]), .A2(b[1]), .ZN(y[145]) );
  OR2_X1 U206bar ( .A1(abar[9]), .A2(bbar[1]), .ZN(ybar[145]);
  AND2_X1 U207 ( .A1(a[9]), .A2(b[0]), .ZN(y[144]) );
  OR2_X1 U207bar ( .A1(abar[9]), .A2(bbar[0]), .ZN(ybar[144]);
  AND2_X1 U208 ( .A1(a[8]), .A2(b[15]), .ZN(y[143]) );
  OR2_X1 U208bar ( .A1(abar[8]), .A2(bbar[15]), .ZN(ybar[143]);
  AND2_X1 U209 ( .A1(a[8]), .A2(b[14]), .ZN(y[142]) );
  OR2_X1 U209bar ( .A1(abar[8]), .A2(bbar[14]), .ZN(ybar[142]);
  AND2_X1 U210 ( .A1(a[8]), .A2(b[13]), .ZN(y[141]) );
  OR2_X1 U210bar ( .A1(abar[8]), .A2(bbar[13]), .ZN(ybar[141]);
  AND2_X1 U211 ( .A1(a[8]), .A2(b[12]), .ZN(y[140]) );
  OR2_X1 U211bar ( .A1(abar[8]), .A2(bbar[12]), .ZN(ybar[140]);
  AND2_X1 U212 ( .A1(b[13]), .A2(a[0]), .ZN(y[13]) );
  OR2_X1 U212bar ( .A1(bbar[13]), .A2(abar[0]), .ZN(ybar[13]);
  AND2_X1 U213 ( .A1(a[8]), .A2(b[11]), .ZN(y[139]) );
  OR2_X1 U213bar ( .A1(abar[8]), .A2(bbar[11]), .ZN(ybar[139]);
  AND2_X1 U214 ( .A1(a[8]), .A2(b[10]), .ZN(y[138]) );
  OR2_X1 U214bar ( .A1(abar[8]), .A2(bbar[10]), .ZN(ybar[138]);
  AND2_X1 U215 ( .A1(a[8]), .A2(b[9]), .ZN(y[137]) );
  OR2_X1 U215bar ( .A1(abar[8]), .A2(bbar[9]), .ZN(ybar[137]);
  AND2_X1 U216 ( .A1(a[8]), .A2(b[8]), .ZN(y[136]) );
  OR2_X1 U216bar ( .A1(abar[8]), .A2(bbar[8]), .ZN(ybar[136]);
  AND2_X1 U217 ( .A1(a[8]), .A2(b[7]), .ZN(y[135]) );
  OR2_X1 U217bar ( .A1(abar[8]), .A2(bbar[7]), .ZN(ybar[135]);
  AND2_X1 U218 ( .A1(a[8]), .A2(b[6]), .ZN(y[134]) );
  OR2_X1 U218bar ( .A1(abar[8]), .A2(bbar[6]), .ZN(ybar[134]);
  AND2_X1 U219 ( .A1(a[8]), .A2(b[5]), .ZN(y[133]) );
  OR2_X1 U219bar ( .A1(abar[8]), .A2(bbar[5]), .ZN(ybar[133]);
  AND2_X1 U220 ( .A1(a[8]), .A2(b[4]), .ZN(y[132]) );
  OR2_X1 U220bar ( .A1(abar[8]), .A2(bbar[4]), .ZN(ybar[132]);
  AND2_X1 U221 ( .A1(a[8]), .A2(b[3]), .ZN(y[131]) );
  OR2_X1 U221bar ( .A1(abar[8]), .A2(bbar[3]), .ZN(ybar[131]);
  AND2_X1 U222 ( .A1(a[8]), .A2(b[2]), .ZN(y[130]) );
  OR2_X1 U222bar ( .A1(abar[8]), .A2(bbar[2]), .ZN(ybar[130]);
  AND2_X1 U223 ( .A1(b[12]), .A2(a[0]), .ZN(y[12]) );
  OR2_X1 U223bar ( .A1(bbar[12]), .A2(abar[0]), .ZN(ybar[12]);
  AND2_X1 U224 ( .A1(a[8]), .A2(b[1]), .ZN(y[129]) );
  OR2_X1 U224bar ( .A1(abar[8]), .A2(bbar[1]), .ZN(ybar[129]);
  AND2_X1 U225 ( .A1(a[8]), .A2(b[0]), .ZN(y[128]) );
  OR2_X1 U225bar ( .A1(abar[8]), .A2(bbar[0]), .ZN(ybar[128]);
  AND2_X1 U226 ( .A1(a[7]), .A2(b[15]), .ZN(y[127]) );
  OR2_X1 U226bar ( .A1(abar[7]), .A2(bbar[15]), .ZN(ybar[127]);
  AND2_X1 U227 ( .A1(a[7]), .A2(b[14]), .ZN(y[126]) );
  OR2_X1 U227bar ( .A1(abar[7]), .A2(bbar[14]), .ZN(ybar[126]);
  AND2_X1 U228 ( .A1(a[7]), .A2(b[13]), .ZN(y[125]) );
  OR2_X1 U228bar ( .A1(abar[7]), .A2(bbar[13]), .ZN(ybar[125]);
  AND2_X1 U229 ( .A1(a[7]), .A2(b[12]), .ZN(y[124]) );
  OR2_X1 U229bar ( .A1(abar[7]), .A2(bbar[12]), .ZN(ybar[124]);
  AND2_X1 U230 ( .A1(a[7]), .A2(b[11]), .ZN(y[123]) );
  OR2_X1 U230bar ( .A1(abar[7]), .A2(bbar[11]), .ZN(ybar[123]);
  AND2_X1 U231 ( .A1(a[7]), .A2(b[10]), .ZN(y[122]) );
  OR2_X1 U231bar ( .A1(abar[7]), .A2(bbar[10]), .ZN(ybar[122]);
  AND2_X1 U232 ( .A1(a[7]), .A2(b[9]), .ZN(y[121]) );
  OR2_X1 U232bar ( .A1(abar[7]), .A2(bbar[9]), .ZN(ybar[121]);
  AND2_X1 U233 ( .A1(a[7]), .A2(b[8]), .ZN(y[120]) );
  OR2_X1 U233bar ( .A1(abar[7]), .A2(bbar[8]), .ZN(ybar[120]);
  AND2_X1 U234 ( .A1(b[11]), .A2(a[0]), .ZN(y[11]) );
  OR2_X1 U234bar ( .A1(bbar[11]), .A2(abar[0]), .ZN(ybar[11]);
  AND2_X1 U235 ( .A1(a[7]), .A2(b[7]), .ZN(y[119]) );
  OR2_X1 U235bar ( .A1(abar[7]), .A2(bbar[7]), .ZN(ybar[119]);
  AND2_X1 U236 ( .A1(a[7]), .A2(b[6]), .ZN(y[118]) );
  OR2_X1 U236bar ( .A1(abar[7]), .A2(bbar[6]), .ZN(ybar[118]);
  AND2_X1 U237 ( .A1(a[7]), .A2(b[5]), .ZN(y[117]) );
  OR2_X1 U237bar ( .A1(abar[7]), .A2(bbar[5]), .ZN(ybar[117]);
  AND2_X1 U238 ( .A1(a[7]), .A2(b[4]), .ZN(y[116]) );
  OR2_X1 U238bar ( .A1(abar[7]), .A2(bbar[4]), .ZN(ybar[116]);
  AND2_X1 U239 ( .A1(a[7]), .A2(b[3]), .ZN(y[115]) );
  OR2_X1 U239bar ( .A1(abar[7]), .A2(bbar[3]), .ZN(ybar[115]);
  AND2_X1 U240 ( .A1(a[7]), .A2(b[2]), .ZN(y[114]) );
  OR2_X1 U240bar ( .A1(abar[7]), .A2(bbar[2]), .ZN(ybar[114]);
  AND2_X1 U241 ( .A1(a[7]), .A2(b[1]), .ZN(y[113]) );
  OR2_X1 U241bar ( .A1(abar[7]), .A2(bbar[1]), .ZN(ybar[113]);
  AND2_X1 U242 ( .A1(a[7]), .A2(b[0]), .ZN(y[112]) );
  OR2_X1 U242bar ( .A1(abar[7]), .A2(bbar[0]), .ZN(ybar[112]);
  AND2_X1 U243 ( .A1(b[15]), .A2(a[6]), .ZN(y[111]) );
  OR2_X1 U243bar ( .A1(bbar[15]), .A2(abar[6]), .ZN(ybar[111]);
  AND2_X1 U244 ( .A1(b[14]), .A2(a[6]), .ZN(y[110]) );
  OR2_X1 U244bar ( .A1(bbar[14]), .A2(abar[6]), .ZN(ybar[110]);
  AND2_X1 U245 ( .A1(b[10]), .A2(a[0]), .ZN(y[10]) );
  OR2_X1 U245bar ( .A1(bbar[10]), .A2(abar[0]), .ZN(ybar[10]);
  AND2_X1 U246 ( .A1(b[13]), .A2(a[6]), .ZN(y[109]) );
  OR2_X1 U246bar ( .A1(bbar[13]), .A2(abar[6]), .ZN(ybar[109]);
  AND2_X1 U247 ( .A1(b[12]), .A2(a[6]), .ZN(y[108]) );
  OR2_X1 U247bar ( .A1(bbar[12]), .A2(abar[6]), .ZN(ybar[108]);
  AND2_X1 U248 ( .A1(b[11]), .A2(a[6]), .ZN(y[107]) );
  OR2_X1 U248bar ( .A1(bbar[11]), .A2(abar[6]), .ZN(ybar[107]);
  AND2_X1 U249 ( .A1(b[10]), .A2(a[6]), .ZN(y[106]) );
  OR2_X1 U249bar ( .A1(bbar[10]), .A2(abar[6]), .ZN(ybar[106]);
  AND2_X1 U250 ( .A1(a[6]), .A2(b[9]), .ZN(y[105]) );
  OR2_X1 U250bar ( .A1(abar[6]), .A2(bbar[9]), .ZN(ybar[105]);
  AND2_X1 U251 ( .A1(b[8]), .A2(a[6]), .ZN(y[104]) );
  OR2_X1 U251bar ( .A1(bbar[8]), .A2(abar[6]), .ZN(ybar[104]);
  AND2_X1 U252 ( .A1(b[7]), .A2(a[6]), .ZN(y[103]) );
  OR2_X1 U252bar ( .A1(bbar[7]), .A2(abar[6]), .ZN(ybar[103]);
  AND2_X1 U253 ( .A1(b[6]), .A2(a[6]), .ZN(y[102]) );
  OR2_X1 U253bar ( .A1(bbar[6]), .A2(abar[6]), .ZN(ybar[102]);
  AND2_X1 U254 ( .A1(b[5]), .A2(a[6]), .ZN(y[101]) );
  OR2_X1 U254bar ( .A1(bbar[5]), .A2(abar[6]), .ZN(ybar[101]);
  AND2_X1 U255 ( .A1(b[4]), .A2(a[6]), .ZN(y[100]) );
  OR2_X1 U255bar ( .A1(bbar[4]), .A2(abar[6]), .ZN(ybar[100]);
  AND2_X1 U256 ( .A1(b[0]), .A2(a[0]), .ZN(y[0]) );
  OR2_X1 U256bar ( .A1(bbar[0]), .A2(abar[0]), .ZN(ybar[0]);
endmodule




module decode_16 ( in, out );
  input [7:0] in;
  //input_done

  output [255:0] out;
  //output_done

  wire   [15:0] level1;
  wire   [31:0] level2;
  //wire_done

  CD2_64 cd_l1_1 ( .a(in[1]), .b(in[0]), .y(level1[3:0]) );
  CD2_63 cd_l1_2 ( .a(in[3]), .b(in[2]), .y(level1[7:4]) );
  CD2_62 cd_l1_3 ( .a(in[5]), .b(in[4]), .y(level1[11:8]) );
  CD2_61 cd_l1_4 ( .a(in[7]), .b(in[6]), .y(level1[15:12]) );
  CD4_32 cd_l2_1 ( .a(level1[7:4]), .b(level1[3:0]), .y(level2[15:0]) );
  CD4_31 cd_l2_2 ( .a(level1[15:12]), .b(level1[11:8]), .y(level2[31:16]) );
  CD16_16 cd_l3 ( .a(level2[31:16]), .b(level2[15:0]), .y(out) );
endmodule


module encode_16 ( in, out );
  input [255:0] in;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
  assign inbar[8] = ~in[8];
  assign inbar[9] = ~in[9];
  assign inbar[10] = ~in[10];
  assign inbar[11] = ~in[11];
  assign inbar[12] = ~in[12];
  assign inbar[13] = ~in[13];
  assign inbar[14] = ~in[14];
  assign inbar[15] = ~in[15];
  assign inbar[16] = ~in[16];
  assign inbar[17] = ~in[17];
  assign inbar[18] = ~in[18];
  assign inbar[19] = ~in[19];
  assign inbar[20] = ~in[20];
  assign inbar[21] = ~in[21];
  assign inbar[22] = ~in[22];
  assign inbar[23] = ~in[23];
  assign inbar[24] = ~in[24];
  assign inbar[25] = ~in[25];
  assign inbar[26] = ~in[26];
  assign inbar[27] = ~in[27];
  assign inbar[28] = ~in[28];
  assign inbar[29] = ~in[29];
  assign inbar[30] = ~in[30];
  assign inbar[31] = ~in[31];
  assign inbar[32] = ~in[32];
  assign inbar[33] = ~in[33];
  assign inbar[34] = ~in[34];
  assign inbar[35] = ~in[35];
  assign inbar[36] = ~in[36];
  assign inbar[37] = ~in[37];
  assign inbar[38] = ~in[38];
  assign inbar[39] = ~in[39];
  assign inbar[40] = ~in[40];
  assign inbar[41] = ~in[41];
  assign inbar[42] = ~in[42];
  assign inbar[43] = ~in[43];
  assign inbar[44] = ~in[44];
  assign inbar[45] = ~in[45];
  assign inbar[46] = ~in[46];
  assign inbar[47] = ~in[47];
  assign inbar[48] = ~in[48];
  assign inbar[49] = ~in[49];
  assign inbar[50] = ~in[50];
  assign inbar[51] = ~in[51];
  assign inbar[52] = ~in[52];
  assign inbar[53] = ~in[53];
  assign inbar[54] = ~in[54];
  assign inbar[55] = ~in[55];
  assign inbar[56] = ~in[56];
  assign inbar[57] = ~in[57];
  assign inbar[58] = ~in[58];
  assign inbar[59] = ~in[59];
  assign inbar[60] = ~in[60];
  assign inbar[61] = ~in[61];
  assign inbar[62] = ~in[62];
  assign inbar[63] = ~in[63];
  assign inbar[64] = ~in[64];
  assign inbar[65] = ~in[65];
  assign inbar[66] = ~in[66];
  assign inbar[67] = ~in[67];
  assign inbar[68] = ~in[68];
  assign inbar[69] = ~in[69];
  assign inbar[70] = ~in[70];
  assign inbar[71] = ~in[71];
  assign inbar[72] = ~in[72];
  assign inbar[73] = ~in[73];
  assign inbar[74] = ~in[74];
  assign inbar[75] = ~in[75];
  assign inbar[76] = ~in[76];
  assign inbar[77] = ~in[77];
  assign inbar[78] = ~in[78];
  assign inbar[79] = ~in[79];
  assign inbar[80] = ~in[80];
  assign inbar[81] = ~in[81];
  assign inbar[82] = ~in[82];
  assign inbar[83] = ~in[83];
  assign inbar[84] = ~in[84];
  assign inbar[85] = ~in[85];
  assign inbar[86] = ~in[86];
  assign inbar[87] = ~in[87];
  assign inbar[88] = ~in[88];
  assign inbar[89] = ~in[89];
  assign inbar[90] = ~in[90];
  assign inbar[91] = ~in[91];
  assign inbar[92] = ~in[92];
  assign inbar[93] = ~in[93];
  assign inbar[94] = ~in[94];
  assign inbar[95] = ~in[95];
  assign inbar[96] = ~in[96];
  assign inbar[97] = ~in[97];
  assign inbar[98] = ~in[98];
  assign inbar[99] = ~in[99];
  assign inbar[100] = ~in[100];
  assign inbar[101] = ~in[101];
  assign inbar[102] = ~in[102];
  assign inbar[103] = ~in[103];
  assign inbar[104] = ~in[104];
  assign inbar[105] = ~in[105];
  assign inbar[106] = ~in[106];
  assign inbar[107] = ~in[107];
  assign inbar[108] = ~in[108];
  assign inbar[109] = ~in[109];
  assign inbar[110] = ~in[110];
  assign inbar[111] = ~in[111];
  assign inbar[112] = ~in[112];
  assign inbar[113] = ~in[113];
  assign inbar[114] = ~in[114];
  assign inbar[115] = ~in[115];
  assign inbar[116] = ~in[116];
  assign inbar[117] = ~in[117];
  assign inbar[118] = ~in[118];
  assign inbar[119] = ~in[119];
  assign inbar[120] = ~in[120];
  assign inbar[121] = ~in[121];
  assign inbar[122] = ~in[122];
  assign inbar[123] = ~in[123];
  assign inbar[124] = ~in[124];
  assign inbar[125] = ~in[125];
  assign inbar[126] = ~in[126];
  assign inbar[127] = ~in[127];
  assign inbar[128] = ~in[128];
  assign inbar[129] = ~in[129];
  assign inbar[130] = ~in[130];
  assign inbar[131] = ~in[131];
  assign inbar[132] = ~in[132];
  assign inbar[133] = ~in[133];
  assign inbar[134] = ~in[134];
  assign inbar[135] = ~in[135];
  assign inbar[136] = ~in[136];
  assign inbar[137] = ~in[137];
  assign inbar[138] = ~in[138];
  assign inbar[139] = ~in[139];
  assign inbar[140] = ~in[140];
  assign inbar[141] = ~in[141];
  assign inbar[142] = ~in[142];
  assign inbar[143] = ~in[143];
  assign inbar[144] = ~in[144];
  assign inbar[145] = ~in[145];
  assign inbar[146] = ~in[146];
  assign inbar[147] = ~in[147];
  assign inbar[148] = ~in[148];
  assign inbar[149] = ~in[149];
  assign inbar[150] = ~in[150];
  assign inbar[151] = ~in[151];
  assign inbar[152] = ~in[152];
  assign inbar[153] = ~in[153];
  assign inbar[154] = ~in[154];
  assign inbar[155] = ~in[155];
  assign inbar[156] = ~in[156];
  assign inbar[157] = ~in[157];
  assign inbar[158] = ~in[158];
  assign inbar[159] = ~in[159];
  assign inbar[160] = ~in[160];
  assign inbar[161] = ~in[161];
  assign inbar[162] = ~in[162];
  assign inbar[163] = ~in[163];
  assign inbar[164] = ~in[164];
  assign inbar[165] = ~in[165];
  assign inbar[166] = ~in[166];
  assign inbar[167] = ~in[167];
  assign inbar[168] = ~in[168];
  assign inbar[169] = ~in[169];
  assign inbar[170] = ~in[170];
  assign inbar[171] = ~in[171];
  assign inbar[172] = ~in[172];
  assign inbar[173] = ~in[173];
  assign inbar[174] = ~in[174];
  assign inbar[175] = ~in[175];
  assign inbar[176] = ~in[176];
  assign inbar[177] = ~in[177];
  assign inbar[178] = ~in[178];
  assign inbar[179] = ~in[179];
  assign inbar[180] = ~in[180];
  assign inbar[181] = ~in[181];
  assign inbar[182] = ~in[182];
  assign inbar[183] = ~in[183];
  assign inbar[184] = ~in[184];
  assign inbar[185] = ~in[185];
  assign inbar[186] = ~in[186];
  assign inbar[187] = ~in[187];
  assign inbar[188] = ~in[188];
  assign inbar[189] = ~in[189];
  assign inbar[190] = ~in[190];
  assign inbar[191] = ~in[191];
  assign inbar[192] = ~in[192];
  assign inbar[193] = ~in[193];
  assign inbar[194] = ~in[194];
  assign inbar[195] = ~in[195];
  assign inbar[196] = ~in[196];
  assign inbar[197] = ~in[197];
  assign inbar[198] = ~in[198];
  assign inbar[199] = ~in[199];
  assign inbar[200] = ~in[200];
  assign inbar[201] = ~in[201];
  assign inbar[202] = ~in[202];
  assign inbar[203] = ~in[203];
  assign inbar[204] = ~in[204];
  assign inbar[205] = ~in[205];
  assign inbar[206] = ~in[206];
  assign inbar[207] = ~in[207];
  assign inbar[208] = ~in[208];
  assign inbar[209] = ~in[209];
  assign inbar[210] = ~in[210];
  assign inbar[211] = ~in[211];
  assign inbar[212] = ~in[212];
  assign inbar[213] = ~in[213];
  assign inbar[214] = ~in[214];
  assign inbar[215] = ~in[215];
  assign inbar[216] = ~in[216];
  assign inbar[217] = ~in[217];
  assign inbar[218] = ~in[218];
  assign inbar[219] = ~in[219];
  assign inbar[220] = ~in[220];
  assign inbar[221] = ~in[221];
  assign inbar[222] = ~in[222];
  assign inbar[223] = ~in[223];
  assign inbar[224] = ~in[224];
  assign inbar[225] = ~in[225];
  assign inbar[226] = ~in[226];
  assign inbar[227] = ~in[227];
  assign inbar[228] = ~in[228];
  assign inbar[229] = ~in[229];
  assign inbar[230] = ~in[230];
  assign inbar[231] = ~in[231];
  assign inbar[232] = ~in[232];
  assign inbar[233] = ~in[233];
  assign inbar[234] = ~in[234];
  assign inbar[235] = ~in[235];
  assign inbar[236] = ~in[236];
  assign inbar[237] = ~in[237];
  assign inbar[238] = ~in[238];
  assign inbar[239] = ~in[239];
  assign inbar[240] = ~in[240];
  assign inbar[241] = ~in[241];
  assign inbar[242] = ~in[242];
  assign inbar[243] = ~in[243];
  assign inbar[244] = ~in[244];
  assign inbar[245] = ~in[245];
  assign inbar[246] = ~in[246];
  assign inbar[247] = ~in[247];
  assign inbar[248] = ~in[248];
  assign inbar[249] = ~in[249];
  assign inbar[250] = ~in[250];
  assign inbar[251] = ~in[251];
  assign inbar[252] = ~in[252];
  assign inbar[253] = ~in[253];
  assign inbar[254] = ~in[254];
  assign inbar[255] = ~in[255];
  //input_done

  output [7:0] out;
  reg [7:0] outbar;
  //output_done

  wire   in_81, in_80, in_79, in_78, in_77, in_76, in_75, in_74, in_73, in_72,
         in_71, in_70, in_69, in_68, in_67, in_66, in_65, in_64, in_63, in_62,
         in_61, in_60, in_59, in_58, in_57, in_56, in_55, in_54, in_53, in_52,
         in_51, in_50, in_49, in_48, in_47, in_46, in_45, in_44, in_43, in_42,
         in_41, in_40, in_39, in_38, in_37, in_36, in_35, in_34, in_33, in_32,
         in_31, in_30, in_29, in_28, in_27, in_26, in_25, in_24, in_23, in_22,
         in_21, in_20, in_19, in_18, in_17, in_16, in_15, in_14, in_13, in_12,
         in_11, in_10, in_9, in_8, in_7, in_6, in_5, in_4, in_3, in_2, in_1,
         in_0, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972;
  wire in_81bar, in_80bar, in_79bar, in_78bar, in_77bar, in_76bar, in_75bar, in_74bar, in_73bar, in_72bar, in_71bar, in_70bar, in_69bar, in_68bar, in_67bar, in_66bar, in_65bar, in_64bar, in_63bar, in_62bar, in_61bar, in_60bar, in_59bar, in_58bar, in_57bar, in_56bar, in_55bar, in_54bar, in_53bar, in_52bar, in_51bar, in_50bar, in_49bar, in_48bar, in_47bar, in_46bar, in_45bar, in_44bar, in_43bar, in_42bar, in_41bar, in_40bar, in_39bar, in_38bar, in_37bar, in_36bar, in_35bar, in_34bar, in_33bar, in_32bar, in_31bar, in_30bar, in_29bar, in_28bar, in_27bar, in_26bar, in_25bar, in_24bar, in_23bar, in_22bar, in_21bar, in_20bar, in_19bar, in_18bar, in_17bar, in_16bar, in_15bar, in_14bar, in_13bar, in_12bar, in_11bar, in_10bar, in_9bar, in_8bar, in_7bar, in_6bar, in_5bar, in_4bar, in_3bar, in_2bar, in_1bar, in_0bar, n487bar, n488bar, n489bar, n490bar, n491bar, n492bar, n493bar, n494bar, n495bar, n496bar, n497bar, n498bar, n499bar, n500bar, n501bar, n502bar, n503bar, n504bar, n505bar, n506bar, n507bar, n508bar, n509bar, n510bar, n511bar, n512bar, n513bar, n514bar, n515bar, n516bar, n517bar, n518bar, n519bar, n520bar, n521bar, n522bar, n523bar, n524bar, n525bar, n526bar, n527bar, n528bar, n529bar, n530bar, n531bar, n532bar, n533bar, n534bar, n535bar, n536bar, n537bar, n538bar, n539bar, n540bar, n541bar, n542bar, n543bar, n544bar, n545bar, n546bar, n547bar, n548bar, n549bar, n550bar, n551bar, n552bar, n553bar, n554bar, n555bar, n556bar, n557bar, n558bar, n559bar, n560bar, n561bar, n562bar, n563bar, n564bar, n565bar, n566bar, n567bar, n568bar, n569bar, n570bar, n571bar, n572bar, n573bar, n574bar, n575bar, n576bar, n577bar, n578bar, n579bar, n580bar, n581bar, n582bar, n583bar, n584bar, n585bar, n586bar, n587bar, n588bar, n589bar, n590bar, n591bar, n592bar, n593bar, n594bar, n595bar, n596bar, n597bar, n598bar, n599bar, n600bar, n601bar, n602bar, n603bar, n604bar, n605bar, n606bar, n607bar, n608bar, n609bar, n610bar, n611bar, n612bar, n613bar, n614bar, n615bar, n616bar, n617bar, n618bar, n619bar, n620bar, n621bar, n622bar, n623bar, n624bar, n625bar, n626bar, n627bar, n628bar, n629bar, n630bar, n631bar, n632bar, n633bar, n634bar, n635bar, n636bar, n637bar, n638bar, n639bar, n640bar, n641bar, n642bar, n643bar, n644bar, n645bar, n646bar, n647bar, n648bar, n649bar, n650bar, n651bar, n652bar, n653bar, n654bar, n655bar, n656bar, n657bar, n658bar, n659bar, n660bar, n661bar, n662bar, n663bar, n664bar, n665bar, n666bar, n667bar, n668bar, n669bar, n670bar, n671bar, n672bar, n673bar, n674bar, n675bar, n676bar, n677bar, n678bar, n679bar, n680bar, n681bar, n682bar, n683bar, n684bar, n685bar, n686bar, n687bar, n688bar, n689bar, n690bar, n691bar, n692bar, n693bar, n694bar, n695bar, n696bar, n697bar, n698bar, n699bar, n700bar, n701bar, n702bar, n703bar, n704bar, n705bar, n706bar, n707bar, n708bar, n709bar, n710bar, n711bar, n712bar, n713bar, n714bar, n715bar, n716bar, n717bar, n718bar, n719bar, n720bar, n721bar, n722bar, n723bar, n724bar, n725bar, n726bar, n727bar, n728bar, n729bar, n730bar, n731bar, n732bar, n733bar, n734bar, n735bar, n736bar, n737bar, n738bar, n739bar, n740bar, n741bar, n742bar, n743bar, n744bar, n745bar, n746bar, n747bar, n748bar, n749bar, n750bar, n751bar, n752bar, n753bar, n754bar, n755bar, n756bar, n757bar, n758bar, n759bar, n760bar, n761bar, n762bar, n763bar, n764bar, n765bar, n766bar, n767bar, n768bar, n769bar, n770bar, n771bar, n772bar, n773bar, n774bar, n775bar, n776bar, n777bar, n778bar, n779bar, n780bar, n781bar, n782bar, n783bar, n784bar, n785bar, n786bar, n787bar, n788bar, n789bar, n790bar, n791bar, n792bar, n793bar, n794bar, n795bar, n796bar, n797bar, n798bar, n799bar, n800bar, n801bar, n802bar, n803bar, n804bar, n805bar, n806bar, n807bar, n808bar, n809bar, n810bar, n811bar, n812bar, n813bar, n814bar, n815bar, n816bar, n817bar, n818bar, n819bar, n820bar, n821bar, n822bar, n823bar, n824bar, n825bar, n826bar, n827bar, n828bar, n829bar, n830bar, n831bar, n832bar, n833bar, n834bar, n835bar, n836bar, n837bar, n838bar, n839bar, n840bar, n841bar, n842bar, n843bar, n844bar, n845bar, n846bar, n847bar, n848bar, n849bar, n850bar, n851bar, n852bar, n853bar, n854bar, n855bar, n856bar, n857bar, n858bar, n859bar, n860bar, n861bar, n862bar, n863bar, n864bar, n865bar, n866bar, n867bar, n868bar, n869bar, n870bar, n871bar, n872bar, n873bar, n874bar, n875bar, n876bar, n877bar, n878bar, n879bar, n880bar, n881bar, n882bar, n883bar, n884bar, n885bar, n886bar, n887bar, n888bar, n889bar, n890bar, n891bar, n892bar, n893bar, n894bar, n895bar, n896bar, n897bar, n898bar, n899bar, n900bar, n901bar, n902bar, n903bar, n904bar, n905bar, n906bar, n907bar, n908bar, n909bar, n910bar, n911bar, n912bar, n913bar, n914bar, n915bar, n916bar, n917bar, n918bar, n919bar, n920bar, n921bar, n922bar, n923bar, n924bar, n925bar, n926bar, n927bar, n928bar, n929bar, n930bar, n931bar, n932bar, n933bar, n934bar, n935bar, n936bar, n937bar, n938bar, n939bar, n940bar, n941bar, n942bar, n943bar, n944bar, n945bar, n946bar, n947bar, n948bar, n949bar, n950bar, n951bar, n952bar, n953bar, n954bar, n955bar, n956bar, n957bar, n958bar, n959bar, n960bar, n961bar, n962bar, n963bar, n964bar, n965bar, n966bar, n967bar, n968bar, n969bar, n970bar, n971bar, n972bar;
  //wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];

  OR2_X1 U1 ( .A1(n972), .A2(n971), .ZN(out[7]) );
  AND2_X1 U1bar ( .A1(n972bar), .A2(n971bar), .ZN(outbar[7]);
  OR2_X1 U2 ( .A1(n970), .A2(n969), .ZN(n971) );
  AND2_X1 U2bar ( .A1(n970bar), .A2(n969bar), .ZN(n971bar);
  OR2_X1 U3 ( .A1(n968), .A2(n967), .ZN(n969) );
  AND2_X1 U3bar ( .A1(n968bar), .A2(n967bar), .ZN(n969bar);
  OR2_X1 U4 ( .A1(n966), .A2(n965), .ZN(n967) );
  AND2_X1 U4bar ( .A1(n966bar), .A2(n965bar), .ZN(n967bar);
  OR2_X1 U5 ( .A1(n964), .A2(n963), .ZN(n968) );
  AND2_X1 U5bar ( .A1(n964bar), .A2(n963bar), .ZN(n968bar);
  OR2_X1 U6 ( .A1(in[116]), .A2(n962), .ZN(n963) );
  AND2_X1 U6bar ( .A1(inbar[116]), .A2(n962bar), .ZN(n963bar);
  OR2_X1 U7 ( .A1(n961), .A2(n960), .ZN(n970) );
  AND2_X1 U7bar ( .A1(n961bar), .A2(n960bar), .ZN(n970bar);
  OR2_X1 U8 ( .A1(in[150]), .A2(in[127]), .ZN(n960) );
  AND2_X1 U8bar ( .A1(inbar[150]), .A2(inbar[127]), .ZN(n960bar);
  OR2_X1 U9 ( .A1(in[160]), .A2(n959), .ZN(n961) );
  AND2_X1 U9bar ( .A1(inbar[160]), .A2(n959bar), .ZN(n961bar);
  OR2_X1 U10 ( .A1(in[252]), .A2(in[168]), .ZN(n959) );
  AND2_X1 U10bar ( .A1(inbar[252]), .A2(inbar[168]), .ZN(n959bar);
  OR2_X1 U11 ( .A1(n958), .A2(n957), .ZN(n972) );
  AND2_X1 U11bar ( .A1(n958bar), .A2(n957bar), .ZN(n972bar);
  OR2_X1 U12 ( .A1(n956), .A2(n955), .ZN(n957) );
  AND2_X1 U12bar ( .A1(n956bar), .A2(n955bar), .ZN(n957bar);
  OR2_X1 U13 ( .A1(in_17), .A2(in[96]), .ZN(n955) );
  AND2_X1 U13bar ( .A1(in_17bar), .A2(inbar[96]), .ZN(n955bar);
  OR2_X1 U14 ( .A1(in_23), .A2(n954), .ZN(n956) );
  AND2_X1 U14bar ( .A1(in_23bar), .A2(n954bar), .ZN(n956bar);
  OR2_X1 U15 ( .A1(in_31), .A2(in_26), .ZN(n954) );
  AND2_X1 U15bar ( .A1(in_31bar), .A2(in_26bar), .ZN(n954bar);
  OR2_X1 U16 ( .A1(n953), .A2(n952), .ZN(n958) );
  AND2_X1 U16bar ( .A1(n953bar), .A2(n952bar), .ZN(n958bar);
  OR2_X1 U17 ( .A1(in_58), .A2(in_4), .ZN(n952) );
  AND2_X1 U17bar ( .A1(in_58bar), .A2(in_4bar), .ZN(n952bar);
  OR2_X1 U18 ( .A1(in_59), .A2(n951), .ZN(n953) );
  AND2_X1 U18bar ( .A1(in_59bar), .A2(n951bar), .ZN(n953bar);
  OR2_X1 U19 ( .A1(in_71), .A2(in_62), .ZN(n951) );
  AND2_X1 U19bar ( .A1(in_71bar), .A2(in_62bar), .ZN(n951bar);
  OR2_X1 U20 ( .A1(n950), .A2(n949), .ZN(out[6]) );
  AND2_X1 U20bar ( .A1(n950bar), .A2(n949bar), .ZN(outbar[6]);
  OR2_X1 U21 ( .A1(n948), .A2(n947), .ZN(n949) );
  AND2_X1 U21bar ( .A1(n948bar), .A2(n947bar), .ZN(n949bar);
  OR2_X1 U22 ( .A1(n946), .A2(n945), .ZN(n947) );
  AND2_X1 U22bar ( .A1(n946bar), .A2(n945bar), .ZN(n947bar);
  OR2_X1 U23 ( .A1(n944), .A2(n943), .ZN(n945) );
  AND2_X1 U23bar ( .A1(n944bar), .A2(n943bar), .ZN(n945bar);
  OR2_X1 U24 ( .A1(n942), .A2(n941), .ZN(n946) );
  AND2_X1 U24bar ( .A1(n942bar), .A2(n941bar), .ZN(n946bar);
  OR2_X1 U25 ( .A1(in[101]), .A2(n940), .ZN(n941) );
  AND2_X1 U25bar ( .A1(inbar[101]), .A2(n940bar), .ZN(n941bar);
  OR2_X1 U26 ( .A1(n939), .A2(n938), .ZN(n948) );
  AND2_X1 U26bar ( .A1(n939bar), .A2(n938bar), .ZN(n948bar);
  OR2_X1 U27 ( .A1(in[114]), .A2(in[104]), .ZN(n938) );
  AND2_X1 U27bar ( .A1(inbar[114]), .A2(inbar[104]), .ZN(n938bar);
  OR2_X1 U28 ( .A1(in[128]), .A2(n937), .ZN(n939) );
  AND2_X1 U28bar ( .A1(inbar[128]), .A2(n937bar), .ZN(n939bar);
  OR2_X1 U29 ( .A1(in[136]), .A2(in[134]), .ZN(n937) );
  AND2_X1 U29bar ( .A1(inbar[136]), .A2(inbar[134]), .ZN(n937bar);
  OR2_X1 U30 ( .A1(n936), .A2(n935), .ZN(n950) );
  AND2_X1 U30bar ( .A1(n936bar), .A2(n935bar), .ZN(n950bar);
  OR2_X1 U31 ( .A1(n934), .A2(n933), .ZN(n935) );
  AND2_X1 U31bar ( .A1(n934bar), .A2(n933bar), .ZN(n935bar);
  OR2_X1 U32 ( .A1(in[177]), .A2(in[164]), .ZN(n933) );
  AND2_X1 U32bar ( .A1(inbar[177]), .A2(inbar[164]), .ZN(n933bar);
  OR2_X1 U33 ( .A1(in[212]), .A2(n932), .ZN(n934) );
  AND2_X1 U33bar ( .A1(inbar[212]), .A2(n932bar), .ZN(n934bar);
  OR2_X1 U34 ( .A1(in[248]), .A2(in[221]), .ZN(n932) );
  AND2_X1 U34bar ( .A1(inbar[248]), .A2(inbar[221]), .ZN(n932bar);
  OR2_X1 U35 ( .A1(n931), .A2(n930), .ZN(n936) );
  AND2_X1 U35bar ( .A1(n931bar), .A2(n930bar), .ZN(n936bar);
  OR2_X1 U36 ( .A1(in_18), .A2(in[93]), .ZN(n930) );
  AND2_X1 U36bar ( .A1(in_18bar), .A2(inbar[93]), .ZN(n930bar);
  OR2_X1 U37 ( .A1(in_31), .A2(n929), .ZN(n931) );
  AND2_X1 U37bar ( .A1(in_31bar), .A2(n929bar), .ZN(n931bar);
  OR2_X1 U38 ( .A1(in_7), .A2(in_39), .ZN(n929) );
  AND2_X1 U38bar ( .A1(in_7bar), .A2(in_39bar), .ZN(n929bar);
  OR2_X1 U39 ( .A1(n928), .A2(n927), .ZN(out[5]) );
  AND2_X1 U39bar ( .A1(n928bar), .A2(n927bar), .ZN(outbar[5]);
  OR2_X1 U40 ( .A1(n926), .A2(n925), .ZN(n927) );
  AND2_X1 U40bar ( .A1(n926bar), .A2(n925bar), .ZN(n927bar);
  OR2_X1 U41 ( .A1(n924), .A2(n923), .ZN(n925) );
  AND2_X1 U41bar ( .A1(n924bar), .A2(n923bar), .ZN(n925bar);
  OR2_X1 U42 ( .A1(n922), .A2(n921), .ZN(n923) );
  AND2_X1 U42bar ( .A1(n922bar), .A2(n921bar), .ZN(n923bar);
  OR2_X1 U43 ( .A1(n940), .A2(n920), .ZN(n924) );
  AND2_X1 U43bar ( .A1(n940bar), .A2(n920bar), .ZN(n924bar);
  OR2_X1 U44 ( .A1(in[111]), .A2(n919), .ZN(n920) );
  AND2_X1 U44bar ( .A1(inbar[111]), .A2(n919bar), .ZN(n920bar);
  OR2_X1 U45 ( .A1(n918), .A2(n917), .ZN(n940) );
  AND2_X1 U45bar ( .A1(n918bar), .A2(n917bar), .ZN(n940bar);
  OR2_X1 U46 ( .A1(n916), .A2(n915), .ZN(n917) );
  AND2_X1 U46bar ( .A1(n916bar), .A2(n915bar), .ZN(n917bar);
  OR2_X1 U47 ( .A1(n914), .A2(n913), .ZN(n915) );
  AND2_X1 U47bar ( .A1(n914bar), .A2(n913bar), .ZN(n915bar);
  OR2_X1 U48 ( .A1(in[140]), .A2(in[131]), .ZN(n913) );
  AND2_X1 U48bar ( .A1(inbar[140]), .A2(inbar[131]), .ZN(n913bar);
  OR2_X1 U49 ( .A1(in[160]), .A2(in[144]), .ZN(n914) );
  AND2_X1 U49bar ( .A1(inbar[160]), .A2(inbar[144]), .ZN(n914bar);
  OR2_X1 U50 ( .A1(n912), .A2(n911), .ZN(n916) );
  AND2_X1 U50bar ( .A1(n912bar), .A2(n911bar), .ZN(n916bar);
  OR2_X1 U51 ( .A1(in[179]), .A2(in[174]), .ZN(n911) );
  AND2_X1 U51bar ( .A1(inbar[179]), .A2(inbar[174]), .ZN(n911bar);
  OR2_X1 U52 ( .A1(in[188]), .A2(in[184]), .ZN(n912) );
  AND2_X1 U52bar ( .A1(inbar[188]), .A2(inbar[184]), .ZN(n912bar);
  OR2_X1 U53 ( .A1(n910), .A2(n909), .ZN(n918) );
  AND2_X1 U53bar ( .A1(n910bar), .A2(n909bar), .ZN(n918bar);
  OR2_X1 U54 ( .A1(n908), .A2(n907), .ZN(n909) );
  AND2_X1 U54bar ( .A1(n908bar), .A2(n907bar), .ZN(n909bar);
  OR2_X1 U55 ( .A1(in[216]), .A2(in[200]), .ZN(n907) );
  AND2_X1 U55bar ( .A1(inbar[216]), .A2(inbar[200]), .ZN(n907bar);
  OR2_X1 U56 ( .A1(in[228]), .A2(in[224]), .ZN(n908) );
  AND2_X1 U56bar ( .A1(inbar[228]), .A2(inbar[224]), .ZN(n908bar);
  OR2_X1 U57 ( .A1(n906), .A2(n905), .ZN(n910) );
  AND2_X1 U57bar ( .A1(n906bar), .A2(n905bar), .ZN(n910bar);
  OR2_X1 U58 ( .A1(in[247]), .A2(in[235]), .ZN(n905) );
  AND2_X1 U58bar ( .A1(inbar[247]), .A2(inbar[235]), .ZN(n905bar);
  OR2_X1 U59 ( .A1(in_42), .A2(in[83]), .ZN(n906) );
  AND2_X1 U59bar ( .A1(in_42bar), .A2(inbar[83]), .ZN(n906bar);
  OR2_X1 U60 ( .A1(n904), .A2(n903), .ZN(n926) );
  AND2_X1 U60bar ( .A1(n904bar), .A2(n903bar), .ZN(n926bar);
  OR2_X1 U61 ( .A1(in[166]), .A2(in[123]), .ZN(n903) );
  AND2_X1 U61bar ( .A1(inbar[166]), .A2(inbar[123]), .ZN(n903bar);
  OR2_X1 U62 ( .A1(in[170]), .A2(n902), .ZN(n904) );
  AND2_X1 U62bar ( .A1(inbar[170]), .A2(n902bar), .ZN(n904bar);
  OR2_X1 U63 ( .A1(in[194]), .A2(in[183]), .ZN(n902) );
  AND2_X1 U63bar ( .A1(inbar[194]), .A2(inbar[183]), .ZN(n902bar);
  OR2_X1 U64 ( .A1(n901), .A2(n900), .ZN(n928) );
  AND2_X1 U64bar ( .A1(n901bar), .A2(n900bar), .ZN(n928bar);
  OR2_X1 U65 ( .A1(n899), .A2(n898), .ZN(n900) );
  AND2_X1 U65bar ( .A1(n899bar), .A2(n898bar), .ZN(n900bar);
  OR2_X1 U66 ( .A1(in[241]), .A2(in[238]), .ZN(n898) );
  AND2_X1 U66bar ( .A1(inbar[241]), .A2(inbar[238]), .ZN(n898bar);
  OR2_X1 U67 ( .A1(in[250]), .A2(n897), .ZN(n899) );
  AND2_X1 U67bar ( .A1(inbar[250]), .A2(n897bar), .ZN(n899bar);
  OR2_X1 U68 ( .A1(in_24), .A2(in[84]), .ZN(n897) );
  AND2_X1 U68bar ( .A1(in_24bar), .A2(inbar[84]), .ZN(n897bar);
  OR2_X1 U69 ( .A1(n896), .A2(n895), .ZN(n901) );
  AND2_X1 U69bar ( .A1(n896bar), .A2(n895bar), .ZN(n901bar);
  OR2_X1 U70 ( .A1(in_41), .A2(in_29), .ZN(n895) );
  AND2_X1 U70bar ( .A1(in_41bar), .A2(in_29bar), .ZN(n895bar);
  OR2_X1 U71 ( .A1(in_66), .A2(n894), .ZN(n896) );
  AND2_X1 U71bar ( .A1(in_66bar), .A2(n894bar), .ZN(n896bar);
  OR2_X1 U72 ( .A1(in_76), .A2(in_71), .ZN(n894) );
  AND2_X1 U72bar ( .A1(in_76bar), .A2(in_71bar), .ZN(n894bar);
  OR2_X1 U73 ( .A1(n893), .A2(n892), .ZN(out[4]) );
  AND2_X1 U73bar ( .A1(n893bar), .A2(n892bar), .ZN(outbar[4]);
  OR2_X1 U74 ( .A1(n891), .A2(n890), .ZN(n892) );
  AND2_X1 U74bar ( .A1(n891bar), .A2(n890bar), .ZN(n892bar);
  OR2_X1 U75 ( .A1(n889), .A2(n888), .ZN(n890) );
  AND2_X1 U75bar ( .A1(n889bar), .A2(n888bar), .ZN(n890bar);
  OR2_X1 U76 ( .A1(n922), .A2(n887), .ZN(n888) );
  AND2_X1 U76bar ( .A1(n922bar), .A2(n887bar), .ZN(n888bar);
  OR2_X1 U77 ( .A1(n886), .A2(n885), .ZN(n922) );
  AND2_X1 U77bar ( .A1(n886bar), .A2(n885bar), .ZN(n922bar);
  OR2_X1 U78 ( .A1(n884), .A2(n883), .ZN(n885) );
  AND2_X1 U78bar ( .A1(n884bar), .A2(n883bar), .ZN(n885bar);
  OR2_X1 U79 ( .A1(n882), .A2(n881), .ZN(n883) );
  AND2_X1 U79bar ( .A1(n882bar), .A2(n881bar), .ZN(n883bar);
  OR2_X1 U80 ( .A1(in[118]), .A2(in[109]), .ZN(n881) );
  AND2_X1 U80bar ( .A1(inbar[118]), .A2(inbar[109]), .ZN(n881bar);
  OR2_X1 U81 ( .A1(in[139]), .A2(in[120]), .ZN(n882) );
  AND2_X1 U81bar ( .A1(inbar[139]), .A2(inbar[120]), .ZN(n882bar);
  OR2_X1 U82 ( .A1(n880), .A2(n879), .ZN(n884) );
  AND2_X1 U82bar ( .A1(n880bar), .A2(n879bar), .ZN(n884bar);
  OR2_X1 U83 ( .A1(in[198]), .A2(in[154]), .ZN(n879) );
  AND2_X1 U83bar ( .A1(inbar[198]), .A2(inbar[154]), .ZN(n879bar);
  OR2_X1 U84 ( .A1(in[210]), .A2(in[205]), .ZN(n880) );
  AND2_X1 U84bar ( .A1(inbar[210]), .A2(inbar[205]), .ZN(n880bar);
  OR2_X1 U85 ( .A1(n878), .A2(n877), .ZN(n886) );
  AND2_X1 U85bar ( .A1(n878bar), .A2(n877bar), .ZN(n886bar);
  OR2_X1 U86 ( .A1(n876), .A2(n875), .ZN(n877) );
  AND2_X1 U86bar ( .A1(n876bar), .A2(n875bar), .ZN(n877bar);
  OR2_X1 U87 ( .A1(in[219]), .A2(in[217]), .ZN(n875) );
  AND2_X1 U87bar ( .A1(inbar[219]), .A2(inbar[217]), .ZN(n875bar);
  OR2_X1 U88 ( .A1(in[86]), .A2(in[252]), .ZN(n876) );
  AND2_X1 U88bar ( .A1(inbar[86]), .A2(inbar[252]), .ZN(n876bar);
  OR2_X1 U89 ( .A1(n874), .A2(n873), .ZN(n878) );
  AND2_X1 U89bar ( .A1(n874bar), .A2(n873bar), .ZN(n878bar);
  OR2_X1 U90 ( .A1(in_40), .A2(in[91]), .ZN(n873) );
  AND2_X1 U90bar ( .A1(in_40bar), .A2(inbar[91]), .ZN(n873bar);
  OR2_X1 U91 ( .A1(in_8), .A2(in_46), .ZN(n874) );
  AND2_X1 U91bar ( .A1(in_8bar), .A2(in_46bar), .ZN(n874bar);
  OR2_X1 U92 ( .A1(n872), .A2(n871), .ZN(n889) );
  AND2_X1 U92bar ( .A1(n872bar), .A2(n871bar), .ZN(n889bar);
  OR2_X1 U93 ( .A1(in[117]), .A2(n943), .ZN(n871) );
  AND2_X1 U93bar ( .A1(inbar[117]), .A2(n943bar), .ZN(n871bar);
  OR2_X1 U94 ( .A1(n870), .A2(n869), .ZN(n943) );
  AND2_X1 U94bar ( .A1(n870bar), .A2(n869bar), .ZN(n943bar);
  OR2_X1 U95 ( .A1(n868), .A2(n867), .ZN(n869) );
  AND2_X1 U95bar ( .A1(n868bar), .A2(n867bar), .ZN(n869bar);
  OR2_X1 U96 ( .A1(n866), .A2(n865), .ZN(n867) );
  AND2_X1 U96bar ( .A1(n866bar), .A2(n865bar), .ZN(n867bar);
  OR2_X1 U97 ( .A1(n864), .A2(n863), .ZN(n865) );
  AND2_X1 U97bar ( .A1(n864bar), .A2(n863bar), .ZN(n865bar);
  OR2_X1 U98 ( .A1(in[108]), .A2(n919), .ZN(n866) );
  AND2_X1 U98bar ( .A1(inbar[108]), .A2(n919bar), .ZN(n866bar);
  OR2_X1 U99 ( .A1(n862), .A2(n861), .ZN(n919) );
  AND2_X1 U99bar ( .A1(n862bar), .A2(n861bar), .ZN(n919bar);
  OR2_X1 U100 ( .A1(n860), .A2(n859), .ZN(n861) );
  AND2_X1 U100bar ( .A1(n860bar), .A2(n859bar), .ZN(n861bar);
  OR2_X1 U101 ( .A1(n858), .A2(n857), .ZN(n859) );
  AND2_X1 U101bar ( .A1(n858bar), .A2(n857bar), .ZN(n859bar);
  OR2_X1 U102 ( .A1(in[119]), .A2(in[105]), .ZN(n857) );
  AND2_X1 U102bar ( .A1(inbar[119]), .A2(inbar[105]), .ZN(n857bar);
  OR2_X1 U103 ( .A1(in[186]), .A2(in[175]), .ZN(n858) );
  AND2_X1 U103bar ( .A1(inbar[186]), .A2(inbar[175]), .ZN(n858bar);
  OR2_X1 U104 ( .A1(n856), .A2(n855), .ZN(n860) );
  AND2_X1 U104bar ( .A1(n856bar), .A2(n855bar), .ZN(n860bar);
  OR2_X1 U105 ( .A1(in[202]), .A2(in[193]), .ZN(n855) );
  AND2_X1 U105bar ( .A1(inbar[202]), .A2(inbar[193]), .ZN(n855bar);
  OR2_X1 U106 ( .A1(in[225]), .A2(in[208]), .ZN(n856) );
  AND2_X1 U106bar ( .A1(inbar[225]), .A2(inbar[208]), .ZN(n856bar);
  OR2_X1 U107 ( .A1(n854), .A2(n853), .ZN(n862) );
  AND2_X1 U107bar ( .A1(n854bar), .A2(n853bar), .ZN(n862bar);
  OR2_X1 U108 ( .A1(n852), .A2(n851), .ZN(n853) );
  AND2_X1 U108bar ( .A1(n852bar), .A2(n851bar), .ZN(n853bar);
  OR2_X1 U109 ( .A1(in_1), .A2(in[85]), .ZN(n851) );
  AND2_X1 U109bar ( .A1(in_1bar), .A2(inbar[85]), .ZN(n851bar);
  OR2_X1 U110 ( .A1(in_23), .A2(in_19), .ZN(n852) );
  AND2_X1 U110bar ( .A1(in_23bar), .A2(in_19bar), .ZN(n852bar);
  OR2_X1 U111 ( .A1(n850), .A2(n849), .ZN(n854) );
  AND2_X1 U111bar ( .A1(n850bar), .A2(n849bar), .ZN(n854bar);
  OR2_X1 U112 ( .A1(in_43), .A2(in_33), .ZN(n849) );
  AND2_X1 U112bar ( .A1(in_43bar), .A2(in_33bar), .ZN(n849bar);
  OR2_X1 U113 ( .A1(in_63), .A2(in_44), .ZN(n850) );
  AND2_X1 U113bar ( .A1(in_63bar), .A2(in_44bar), .ZN(n850bar);
  OR2_X1 U114 ( .A1(n848), .A2(n847), .ZN(n868) );
  AND2_X1 U114bar ( .A1(n848bar), .A2(n847bar), .ZN(n868bar);
  OR2_X1 U115 ( .A1(in[141]), .A2(in[112]), .ZN(n847) );
  AND2_X1 U115bar ( .A1(inbar[141]), .A2(inbar[112]), .ZN(n847bar);
  OR2_X1 U116 ( .A1(in[147]), .A2(n846), .ZN(n848) );
  AND2_X1 U116bar ( .A1(inbar[147]), .A2(n846bar), .ZN(n848bar);
  OR2_X1 U117 ( .A1(in[181]), .A2(in[167]), .ZN(n846) );
  AND2_X1 U117bar ( .A1(inbar[181]), .A2(inbar[167]), .ZN(n846bar);
  OR2_X1 U118 ( .A1(n845), .A2(n844), .ZN(n870) );
  AND2_X1 U118bar ( .A1(n845bar), .A2(n844bar), .ZN(n870bar);
  OR2_X1 U119 ( .A1(n843), .A2(n842), .ZN(n844) );
  AND2_X1 U119bar ( .A1(n843bar), .A2(n842bar), .ZN(n844bar);
  OR2_X1 U120 ( .A1(in[229]), .A2(in[201]), .ZN(n842) );
  AND2_X1 U120bar ( .A1(inbar[229]), .A2(inbar[201]), .ZN(n842bar);
  OR2_X1 U121 ( .A1(in[237]), .A2(n841), .ZN(n843) );
  AND2_X1 U121bar ( .A1(inbar[237]), .A2(n841bar), .ZN(n843bar);
  OR2_X1 U122 ( .A1(in[94]), .A2(in[253]), .ZN(n841) );
  AND2_X1 U122bar ( .A1(inbar[94]), .A2(inbar[253]), .ZN(n841bar);
  OR2_X1 U123 ( .A1(n840), .A2(n839), .ZN(n845) );
  AND2_X1 U123bar ( .A1(n840bar), .A2(n839bar), .ZN(n845bar);
  OR2_X1 U124 ( .A1(in_21), .A2(in[96]), .ZN(n839) );
  AND2_X1 U124bar ( .A1(in_21bar), .A2(inbar[96]), .ZN(n839bar);
  OR2_X1 U125 ( .A1(in_25), .A2(n838), .ZN(n840) );
  AND2_X1 U125bar ( .A1(in_25bar), .A2(n838bar), .ZN(n840bar);
  OR2_X1 U126 ( .A1(in_81), .A2(in_45), .ZN(n838) );
  AND2_X1 U126bar ( .A1(in_81bar), .A2(in_45bar), .ZN(n838bar);
  OR2_X1 U127 ( .A1(n837), .A2(n836), .ZN(n891) );
  AND2_X1 U127bar ( .A1(n837bar), .A2(n836bar), .ZN(n891bar);
  OR2_X1 U128 ( .A1(in[142]), .A2(in[124]), .ZN(n836) );
  AND2_X1 U128bar ( .A1(inbar[142]), .A2(inbar[124]), .ZN(n836bar);
  OR2_X1 U129 ( .A1(in[150]), .A2(n835), .ZN(n837) );
  AND2_X1 U129bar ( .A1(inbar[150]), .A2(n835bar), .ZN(n837bar);
  OR2_X1 U130 ( .A1(in[172]), .A2(in[155]), .ZN(n835) );
  AND2_X1 U130bar ( .A1(inbar[172]), .A2(inbar[155]), .ZN(n835bar);
  OR2_X1 U131 ( .A1(n834), .A2(n833), .ZN(n893) );
  AND2_X1 U131bar ( .A1(n834bar), .A2(n833bar), .ZN(n893bar);
  OR2_X1 U132 ( .A1(n832), .A2(n831), .ZN(n833) );
  AND2_X1 U132bar ( .A1(n832bar), .A2(n831bar), .ZN(n833bar);
  OR2_X1 U133 ( .A1(in[196]), .A2(in[173]), .ZN(n831) );
  AND2_X1 U133bar ( .A1(inbar[196]), .A2(inbar[173]), .ZN(n831bar);
  OR2_X1 U134 ( .A1(in[222]), .A2(n830), .ZN(n832) );
  AND2_X1 U134bar ( .A1(inbar[222]), .A2(n830bar), .ZN(n832bar);
  OR2_X1 U135 ( .A1(in[227]), .A2(in[226]), .ZN(n830) );
  AND2_X1 U135bar ( .A1(inbar[227]), .A2(inbar[226]), .ZN(n830bar);
  OR2_X1 U136 ( .A1(n829), .A2(n828), .ZN(n834) );
  AND2_X1 U136bar ( .A1(n829bar), .A2(n828bar), .ZN(n834bar);
  OR2_X1 U137 ( .A1(in[249]), .A2(in[231]), .ZN(n828) );
  AND2_X1 U137bar ( .A1(inbar[249]), .A2(inbar[231]), .ZN(n828bar);
  OR2_X1 U138 ( .A1(in_28), .A2(n827), .ZN(n829) );
  AND2_X1 U138bar ( .A1(in_28bar), .A2(n827bar), .ZN(n829bar);
  OR2_X1 U139 ( .A1(in_52), .A2(in_47), .ZN(n827) );
  AND2_X1 U139bar ( .A1(in_52bar), .A2(in_47bar), .ZN(n827bar);
  OR2_X1 U140 ( .A1(n826), .A2(n825), .ZN(out[3]) );
  AND2_X1 U140bar ( .A1(n826bar), .A2(n825bar), .ZN(outbar[3]);
  OR2_X1 U141 ( .A1(n824), .A2(n823), .ZN(n825) );
  AND2_X1 U141bar ( .A1(n824bar), .A2(n823bar), .ZN(n825bar);
  OR2_X1 U142 ( .A1(n822), .A2(n821), .ZN(n823) );
  AND2_X1 U142bar ( .A1(n822bar), .A2(n821bar), .ZN(n823bar);
  OR2_X1 U143 ( .A1(n820), .A2(n819), .ZN(n821) );
  AND2_X1 U143bar ( .A1(n820bar), .A2(n819bar), .ZN(n821bar);
  OR2_X1 U144 ( .A1(n964), .A2(n818), .ZN(n822) );
  AND2_X1 U144bar ( .A1(n964bar), .A2(n818bar), .ZN(n822bar);
  OR2_X1 U145 ( .A1(in[118]), .A2(n817), .ZN(n818) );
  AND2_X1 U145bar ( .A1(inbar[118]), .A2(n817bar), .ZN(n818bar);
  OR2_X1 U146 ( .A1(n816), .A2(n815), .ZN(n964) );
  AND2_X1 U146bar ( .A1(n816bar), .A2(n815bar), .ZN(n964bar);
  OR2_X1 U147 ( .A1(n814), .A2(n813), .ZN(n815) );
  AND2_X1 U147bar ( .A1(n814bar), .A2(n813bar), .ZN(n815bar);
  OR2_X1 U148 ( .A1(n812), .A2(n811), .ZN(n813) );
  AND2_X1 U148bar ( .A1(n812bar), .A2(n811bar), .ZN(n813bar);
  OR2_X1 U149 ( .A1(in[122]), .A2(in[111]), .ZN(n811) );
  AND2_X1 U149bar ( .A1(inbar[122]), .A2(inbar[111]), .ZN(n811bar);
  OR2_X1 U150 ( .A1(in[154]), .A2(in[151]), .ZN(n812) );
  AND2_X1 U150bar ( .A1(inbar[154]), .A2(inbar[151]), .ZN(n812bar);
  OR2_X1 U151 ( .A1(n810), .A2(n809), .ZN(n814) );
  AND2_X1 U151bar ( .A1(n810bar), .A2(n809bar), .ZN(n814bar);
  OR2_X1 U152 ( .A1(in[187]), .A2(in[177]), .ZN(n809) );
  AND2_X1 U152bar ( .A1(inbar[187]), .A2(inbar[177]), .ZN(n809bar);
  OR2_X1 U153 ( .A1(in[200]), .A2(in[192]), .ZN(n810) );
  AND2_X1 U153bar ( .A1(inbar[200]), .A2(inbar[192]), .ZN(n810bar);
  OR2_X1 U154 ( .A1(n808), .A2(n807), .ZN(n816) );
  AND2_X1 U154bar ( .A1(n808bar), .A2(n807bar), .ZN(n816bar);
  OR2_X1 U155 ( .A1(n806), .A2(n805), .ZN(n807) );
  AND2_X1 U155bar ( .A1(n806bar), .A2(n805bar), .ZN(n807bar);
  OR2_X1 U156 ( .A1(in[225]), .A2(in[207]), .ZN(n805) );
  AND2_X1 U156bar ( .A1(inbar[225]), .A2(inbar[207]), .ZN(n805bar);
  OR2_X1 U157 ( .A1(in[98]), .A2(in[226]), .ZN(n806) );
  AND2_X1 U157bar ( .A1(inbar[98]), .A2(inbar[226]), .ZN(n806bar);
  OR2_X1 U158 ( .A1(n804), .A2(n803), .ZN(n808) );
  AND2_X1 U158bar ( .A1(n804bar), .A2(n803bar), .ZN(n808bar);
  OR2_X1 U159 ( .A1(in_20), .A2(in_16), .ZN(n803) );
  AND2_X1 U159bar ( .A1(in_20bar), .A2(in_16bar), .ZN(n803bar);
  OR2_X1 U160 ( .A1(in_55), .A2(in_45), .ZN(n804) );
  AND2_X1 U160bar ( .A1(in_55bar), .A2(in_45bar), .ZN(n804bar);
  OR2_X1 U161 ( .A1(n802), .A2(n801), .ZN(n824) );
  AND2_X1 U161bar ( .A1(n802bar), .A2(n801bar), .ZN(n824bar);
  OR2_X1 U162 ( .A1(in[162]), .A2(in[149]), .ZN(n801) );
  AND2_X1 U162bar ( .A1(inbar[162]), .A2(inbar[149]), .ZN(n801bar);
  OR2_X1 U163 ( .A1(in[163]), .A2(n800), .ZN(n802) );
  AND2_X1 U163bar ( .A1(inbar[163]), .A2(n800bar), .ZN(n802bar);
  OR2_X1 U164 ( .A1(in[191]), .A2(in[189]), .ZN(n800) );
  AND2_X1 U164bar ( .A1(inbar[191]), .A2(inbar[189]), .ZN(n800bar);
  OR2_X1 U165 ( .A1(n799), .A2(n798), .ZN(n826) );
  AND2_X1 U165bar ( .A1(n799bar), .A2(n798bar), .ZN(n826bar);
  OR2_X1 U166 ( .A1(n797), .A2(n796), .ZN(n798) );
  AND2_X1 U166bar ( .A1(n797bar), .A2(n796bar), .ZN(n798bar);
  OR2_X1 U167 ( .A1(in[212]), .A2(in[193]), .ZN(n796) );
  AND2_X1 U167bar ( .A1(inbar[212]), .A2(inbar[193]), .ZN(n796bar);
  OR2_X1 U168 ( .A1(in[238]), .A2(n795), .ZN(n797) );
  AND2_X1 U168bar ( .A1(inbar[238]), .A2(n795bar), .ZN(n797bar);
  OR2_X1 U169 ( .A1(in[88]), .A2(in[247]), .ZN(n795) );
  AND2_X1 U169bar ( .A1(inbar[88]), .A2(inbar[247]), .ZN(n795bar);
  OR2_X1 U170 ( .A1(n794), .A2(n793), .ZN(n799) );
  AND2_X1 U170bar ( .A1(n794bar), .A2(n793bar), .ZN(n799bar);
  OR2_X1 U171 ( .A1(in[94]), .A2(in[92]), .ZN(n793) );
  AND2_X1 U171bar ( .A1(inbar[94]), .A2(inbar[92]), .ZN(n793bar);
  OR2_X1 U172 ( .A1(in_52), .A2(n792), .ZN(n794) );
  AND2_X1 U172bar ( .A1(in_52bar), .A2(n792bar), .ZN(n794bar);
  OR2_X1 U173 ( .A1(in_70), .A2(in_67), .ZN(n792) );
  AND2_X1 U173bar ( .A1(in_70bar), .A2(in_67bar), .ZN(n792bar);
  OR2_X1 U174 ( .A1(n791), .A2(n790), .ZN(out[2]) );
  AND2_X1 U174bar ( .A1(n791bar), .A2(n790bar), .ZN(outbar[2]);
  OR2_X1 U175 ( .A1(n789), .A2(n788), .ZN(n790) );
  AND2_X1 U175bar ( .A1(n789bar), .A2(n788bar), .ZN(n790bar);
  OR2_X1 U176 ( .A1(n787), .A2(n786), .ZN(n788) );
  AND2_X1 U176bar ( .A1(n787bar), .A2(n786bar), .ZN(n788bar);
  OR2_X1 U177 ( .A1(n819), .A2(n785), .ZN(n786) );
  AND2_X1 U177bar ( .A1(n819bar), .A2(n785bar), .ZN(n786bar);
  OR2_X1 U178 ( .A1(n784), .A2(n783), .ZN(n819) );
  AND2_X1 U178bar ( .A1(n784bar), .A2(n783bar), .ZN(n819bar);
  OR2_X1 U179 ( .A1(n782), .A2(n781), .ZN(n783) );
  AND2_X1 U179bar ( .A1(n782bar), .A2(n781bar), .ZN(n783bar);
  OR2_X1 U180 ( .A1(n780), .A2(n779), .ZN(n781) );
  AND2_X1 U180bar ( .A1(n780bar), .A2(n779bar), .ZN(n781bar);
  OR2_X1 U181 ( .A1(n962), .A2(n778), .ZN(n779) );
  AND2_X1 U181bar ( .A1(n962bar), .A2(n778bar), .ZN(n779bar);
  OR2_X1 U182 ( .A1(n777), .A2(n776), .ZN(n962) );
  AND2_X1 U182bar ( .A1(n777bar), .A2(n776bar), .ZN(n962bar);
  OR2_X1 U183 ( .A1(n775), .A2(n774), .ZN(n776) );
  AND2_X1 U183bar ( .A1(n775bar), .A2(n774bar), .ZN(n776bar);
  OR2_X1 U184 ( .A1(n773), .A2(n772), .ZN(n774) );
  AND2_X1 U184bar ( .A1(n773bar), .A2(n772bar), .ZN(n774bar);
  OR2_X1 U185 ( .A1(in[131]), .A2(in[120]), .ZN(n772) );
  AND2_X1 U185bar ( .A1(inbar[131]), .A2(inbar[120]), .ZN(n772bar);
  OR2_X1 U186 ( .A1(in[153]), .A2(in[147]), .ZN(n773) );
  AND2_X1 U186bar ( .A1(inbar[153]), .A2(inbar[147]), .ZN(n773bar);
  OR2_X1 U187 ( .A1(n771), .A2(n770), .ZN(n775) );
  AND2_X1 U187bar ( .A1(n771bar), .A2(n770bar), .ZN(n775bar);
  OR2_X1 U188 ( .A1(in[170]), .A2(in[156]), .ZN(n770) );
  AND2_X1 U188bar ( .A1(inbar[170]), .A2(inbar[156]), .ZN(n770bar);
  OR2_X1 U189 ( .A1(in[223]), .A2(in[190]), .ZN(n771) );
  AND2_X1 U189bar ( .A1(inbar[223]), .A2(inbar[190]), .ZN(n771bar);
  OR2_X1 U190 ( .A1(n769), .A2(n768), .ZN(n777) );
  AND2_X1 U190bar ( .A1(n769bar), .A2(n768bar), .ZN(n777bar);
  OR2_X1 U191 ( .A1(n767), .A2(n766), .ZN(n768) );
  AND2_X1 U191bar ( .A1(n767bar), .A2(n766bar), .ZN(n768bar);
  OR2_X1 U192 ( .A1(in[236]), .A2(in[230]), .ZN(n766) );
  AND2_X1 U192bar ( .A1(inbar[236]), .A2(inbar[230]), .ZN(n766bar);
  OR2_X1 U193 ( .A1(in[85]), .A2(in[240]), .ZN(n767) );
  AND2_X1 U193bar ( .A1(inbar[85]), .A2(inbar[240]), .ZN(n767bar);
  OR2_X1 U194 ( .A1(n765), .A2(n764), .ZN(n769) );
  AND2_X1 U194bar ( .A1(n765bar), .A2(n764bar), .ZN(n769bar);
  OR2_X1 U195 ( .A1(in_12), .A2(in[90]), .ZN(n764) );
  AND2_X1 U195bar ( .A1(in_12bar), .A2(inbar[90]), .ZN(n764bar);
  OR2_X1 U196 ( .A1(in_39), .A2(in_28), .ZN(n765) );
  AND2_X1 U196bar ( .A1(in_39bar), .A2(in_28bar), .ZN(n765bar);
  OR2_X1 U197 ( .A1(in[109]), .A2(n763), .ZN(n780) );
  AND2_X1 U197bar ( .A1(inbar[109]), .A2(n763bar), .ZN(n780bar);
  OR2_X1 U198 ( .A1(n762), .A2(n761), .ZN(n782) );
  AND2_X1 U198bar ( .A1(n762bar), .A2(n761bar), .ZN(n782bar);
  OR2_X1 U199 ( .A1(in[138]), .A2(in[129]), .ZN(n761) );
  AND2_X1 U199bar ( .A1(inbar[138]), .A2(inbar[129]), .ZN(n761bar);
  OR2_X1 U200 ( .A1(in[157]), .A2(n760), .ZN(n762) );
  AND2_X1 U200bar ( .A1(inbar[157]), .A2(n760bar), .ZN(n762bar);
  OR2_X1 U201 ( .A1(in[182]), .A2(in[167]), .ZN(n760) );
  AND2_X1 U201bar ( .A1(inbar[182]), .A2(inbar[167]), .ZN(n760bar);
  OR2_X1 U202 ( .A1(n759), .A2(n758), .ZN(n784) );
  AND2_X1 U202bar ( .A1(n759bar), .A2(n758bar), .ZN(n784bar);
  OR2_X1 U203 ( .A1(n757), .A2(n756), .ZN(n758) );
  AND2_X1 U203bar ( .A1(n757bar), .A2(n756bar), .ZN(n758bar);
  OR2_X1 U204 ( .A1(in[195]), .A2(in[184]), .ZN(n756) );
  AND2_X1 U204bar ( .A1(inbar[195]), .A2(inbar[184]), .ZN(n756bar);
  OR2_X1 U205 ( .A1(in[196]), .A2(n755), .ZN(n757) );
  AND2_X1 U205bar ( .A1(inbar[196]), .A2(n755bar), .ZN(n757bar);
  OR2_X1 U206 ( .A1(in[215]), .A2(in[209]), .ZN(n755) );
  AND2_X1 U206bar ( .A1(inbar[215]), .A2(inbar[209]), .ZN(n755bar);
  OR2_X1 U207 ( .A1(n754), .A2(n753), .ZN(n759) );
  AND2_X1 U207bar ( .A1(n754bar), .A2(n753bar), .ZN(n759bar);
  OR2_X1 U208 ( .A1(in[93]), .A2(in[233]), .ZN(n753) );
  AND2_X1 U208bar ( .A1(inbar[93]), .A2(inbar[233]), .ZN(n753bar);
  OR2_X1 U209 ( .A1(in_1), .A2(n752), .ZN(n754) );
  AND2_X1 U209bar ( .A1(in_1bar), .A2(n752bar), .ZN(n754bar);
  OR2_X1 U210 ( .A1(in_69), .A2(in_66), .ZN(n752) );
  AND2_X1 U210bar ( .A1(in_69bar), .A2(in_66bar), .ZN(n752bar);
  OR2_X1 U211 ( .A1(n966), .A2(n751), .ZN(n787) );
  AND2_X1 U211bar ( .A1(n966bar), .A2(n751bar), .ZN(n787bar);
  OR2_X1 U212 ( .A1(in[134]), .A2(n750), .ZN(n751) );
  AND2_X1 U212bar ( .A1(inbar[134]), .A2(n750bar), .ZN(n751bar);
  OR2_X1 U213 ( .A1(n749), .A2(n748), .ZN(n966) );
  AND2_X1 U213bar ( .A1(n749bar), .A2(n748bar), .ZN(n966bar);
  OR2_X1 U214 ( .A1(n747), .A2(n746), .ZN(n748) );
  AND2_X1 U214bar ( .A1(n747bar), .A2(n746bar), .ZN(n748bar);
  OR2_X1 U215 ( .A1(n745), .A2(n744), .ZN(n746) );
  AND2_X1 U215bar ( .A1(n745bar), .A2(n744bar), .ZN(n746bar);
  OR2_X1 U216 ( .A1(in[136]), .A2(in[121]), .ZN(n744) );
  AND2_X1 U216bar ( .A1(inbar[136]), .A2(inbar[121]), .ZN(n744bar);
  OR2_X1 U217 ( .A1(in[186]), .A2(in[174]), .ZN(n745) );
  AND2_X1 U217bar ( .A1(inbar[186]), .A2(inbar[174]), .ZN(n745bar);
  OR2_X1 U218 ( .A1(n743), .A2(n742), .ZN(n747) );
  AND2_X1 U218bar ( .A1(n743bar), .A2(n742bar), .ZN(n747bar);
  OR2_X1 U219 ( .A1(in[198]), .A2(in[197]), .ZN(n742) );
  AND2_X1 U219bar ( .A1(inbar[198]), .A2(inbar[197]), .ZN(n742bar);
  OR2_X1 U220 ( .A1(in[214]), .A2(in[199]), .ZN(n743) );
  AND2_X1 U220bar ( .A1(inbar[214]), .A2(inbar[199]), .ZN(n743bar);
  OR2_X1 U221 ( .A1(n741), .A2(n740), .ZN(n749) );
  AND2_X1 U221bar ( .A1(n741bar), .A2(n740bar), .ZN(n749bar);
  OR2_X1 U222 ( .A1(n739), .A2(n738), .ZN(n740) );
  AND2_X1 U222bar ( .A1(n739bar), .A2(n738bar), .ZN(n740bar);
  OR2_X1 U223 ( .A1(in[231]), .A2(in[220]), .ZN(n738) );
  AND2_X1 U223bar ( .A1(inbar[231]), .A2(inbar[220]), .ZN(n738bar);
  OR2_X1 U224 ( .A1(in_25), .A2(in[245]), .ZN(n739) );
  AND2_X1 U224bar ( .A1(in_25bar), .A2(inbar[245]), .ZN(n739bar);
  OR2_X1 U225 ( .A1(n737), .A2(n736), .ZN(n741) );
  AND2_X1 U225bar ( .A1(n737bar), .A2(n736bar), .ZN(n741bar);
  OR2_X1 U226 ( .A1(in_53), .A2(in_29), .ZN(n736) );
  AND2_X1 U226bar ( .A1(in_53bar), .A2(in_29bar), .ZN(n736bar);
  OR2_X1 U227 ( .A1(in_79), .A2(in_74), .ZN(n737) );
  AND2_X1 U227bar ( .A1(in_79bar), .A2(in_74bar), .ZN(n737bar);
  OR2_X1 U228 ( .A1(n735), .A2(n734), .ZN(n789) );
  AND2_X1 U228bar ( .A1(n735bar), .A2(n734bar), .ZN(n789bar);
  OR2_X1 U229 ( .A1(in[152]), .A2(in[140]), .ZN(n734) );
  AND2_X1 U229bar ( .A1(inbar[152]), .A2(inbar[140]), .ZN(n734bar);
  OR2_X1 U230 ( .A1(in[155]), .A2(n733), .ZN(n735) );
  AND2_X1 U230bar ( .A1(inbar[155]), .A2(n733bar), .ZN(n735bar);
  OR2_X1 U231 ( .A1(in[166]), .A2(in[165]), .ZN(n733) );
  AND2_X1 U231bar ( .A1(inbar[166]), .A2(inbar[165]), .ZN(n733bar);
  OR2_X1 U232 ( .A1(n732), .A2(n731), .ZN(n791) );
  AND2_X1 U232bar ( .A1(n732bar), .A2(n731bar), .ZN(n791bar);
  OR2_X1 U233 ( .A1(n730), .A2(n729), .ZN(n731) );
  AND2_X1 U233bar ( .A1(n730bar), .A2(n729bar), .ZN(n731bar);
  OR2_X1 U234 ( .A1(in[202]), .A2(in[185]), .ZN(n729) );
  AND2_X1 U234bar ( .A1(inbar[202]), .A2(inbar[185]), .ZN(n729bar);
  OR2_X1 U235 ( .A1(in[211]), .A2(n728), .ZN(n730) );
  AND2_X1 U235bar ( .A1(inbar[211]), .A2(n728bar), .ZN(n730bar);
  OR2_X1 U236 ( .A1(in[255]), .A2(in[253]), .ZN(n728) );
  AND2_X1 U236bar ( .A1(inbar[255]), .A2(inbar[253]), .ZN(n728bar);
  OR2_X1 U237 ( .A1(n727), .A2(n726), .ZN(n732) );
  AND2_X1 U237bar ( .A1(n727bar), .A2(n726bar), .ZN(n732bar);
  OR2_X1 U238 ( .A1(in_35), .A2(in_15), .ZN(n726) );
  AND2_X1 U238bar ( .A1(in_35bar), .A2(in_15bar), .ZN(n726bar);
  OR2_X1 U239 ( .A1(in_36), .A2(n725), .ZN(n727) );
  AND2_X1 U239bar ( .A1(in_36bar), .A2(n725bar), .ZN(n727bar);
  OR2_X1 U240 ( .A1(in_48), .A2(in_40), .ZN(n725) );
  AND2_X1 U240bar ( .A1(in_48bar), .A2(in_40bar), .ZN(n725bar);
  OR2_X1 U241 ( .A1(n724), .A2(n723), .ZN(out[1]) );
  AND2_X1 U241bar ( .A1(n724bar), .A2(n723bar), .ZN(outbar[1]);
  OR2_X1 U242 ( .A1(n722), .A2(n721), .ZN(n723) );
  AND2_X1 U242bar ( .A1(n722bar), .A2(n721bar), .ZN(n723bar);
  OR2_X1 U243 ( .A1(n720), .A2(n719), .ZN(n721) );
  AND2_X1 U243bar ( .A1(n720bar), .A2(n719bar), .ZN(n721bar);
  OR2_X1 U244 ( .A1(n921), .A2(n887), .ZN(n719) );
  AND2_X1 U244bar ( .A1(n921bar), .A2(n887bar), .ZN(n719bar);
  OR2_X1 U245 ( .A1(n718), .A2(n717), .ZN(n887) );
  AND2_X1 U245bar ( .A1(n718bar), .A2(n717bar), .ZN(n887bar);
  OR2_X1 U246 ( .A1(n716), .A2(n715), .ZN(n717) );
  AND2_X1 U246bar ( .A1(n716bar), .A2(n715bar), .ZN(n717bar);
  OR2_X1 U247 ( .A1(n714), .A2(n713), .ZN(n715) );
  AND2_X1 U247bar ( .A1(n714bar), .A2(n713bar), .ZN(n715bar);
  OR2_X1 U248 ( .A1(in[116]), .A2(in[110]), .ZN(n713) );
  AND2_X1 U248bar ( .A1(inbar[116]), .A2(inbar[110]), .ZN(n713bar);
  OR2_X1 U249 ( .A1(in[133]), .A2(in[130]), .ZN(n714) );
  AND2_X1 U249bar ( .A1(inbar[133]), .A2(inbar[130]), .ZN(n714bar);
  OR2_X1 U250 ( .A1(n712), .A2(n711), .ZN(n716) );
  AND2_X1 U250bar ( .A1(n712bar), .A2(n711bar), .ZN(n716bar);
  OR2_X1 U251 ( .A1(in[203]), .A2(in[135]), .ZN(n711) );
  AND2_X1 U251bar ( .A1(inbar[203]), .A2(inbar[135]), .ZN(n711bar);
  OR2_X1 U252 ( .A1(in[232]), .A2(in[223]), .ZN(n712) );
  AND2_X1 U252bar ( .A1(inbar[232]), .A2(inbar[223]), .ZN(n712bar);
  OR2_X1 U253 ( .A1(n710), .A2(n709), .ZN(n718) );
  AND2_X1 U253bar ( .A1(n710bar), .A2(n709bar), .ZN(n718bar);
  OR2_X1 U254 ( .A1(n708), .A2(n707), .ZN(n709) );
  AND2_X1 U254bar ( .A1(n708bar), .A2(n707bar), .ZN(n709bar);
  OR2_X1 U255 ( .A1(in[255]), .A2(in[233]), .ZN(n707) );
  AND2_X1 U255bar ( .A1(inbar[255]), .A2(inbar[233]), .ZN(n707bar);
  OR2_X1 U256 ( .A1(in_53), .A2(in_34), .ZN(n708) );
  AND2_X1 U256bar ( .A1(in_53bar), .A2(in_34bar), .ZN(n708bar);
  OR2_X1 U257 ( .A1(n706), .A2(n705), .ZN(n710) );
  AND2_X1 U257bar ( .A1(n706bar), .A2(n705bar), .ZN(n710bar);
  OR2_X1 U258 ( .A1(in_57), .A2(in_55), .ZN(n705) );
  AND2_X1 U258bar ( .A1(in_57bar), .A2(in_55bar), .ZN(n705bar);
  OR2_X1 U259 ( .A1(in_68), .A2(in_67), .ZN(n706) );
  AND2_X1 U259bar ( .A1(in_68bar), .A2(in_67bar), .ZN(n706bar);
  OR2_X1 U260 ( .A1(n704), .A2(n703), .ZN(n921) );
  AND2_X1 U260bar ( .A1(n704bar), .A2(n703bar), .ZN(n921bar);
  OR2_X1 U261 ( .A1(n702), .A2(n701), .ZN(n703) );
  AND2_X1 U261bar ( .A1(n702bar), .A2(n701bar), .ZN(n703bar);
  OR2_X1 U262 ( .A1(n700), .A2(n699), .ZN(n701) );
  AND2_X1 U262bar ( .A1(n700bar), .A2(n699bar), .ZN(n701bar);
  OR2_X1 U263 ( .A1(n944), .A2(n872), .ZN(n699) );
  AND2_X1 U263bar ( .A1(n944bar), .A2(n872bar), .ZN(n699bar);
  OR2_X1 U264 ( .A1(n698), .A2(n697), .ZN(n872) );
  AND2_X1 U264bar ( .A1(n698bar), .A2(n697bar), .ZN(n872bar);
  OR2_X1 U265 ( .A1(n696), .A2(n695), .ZN(n697) );
  AND2_X1 U265bar ( .A1(n696bar), .A2(n695bar), .ZN(n697bar);
  OR2_X1 U266 ( .A1(n694), .A2(n693), .ZN(n695) );
  AND2_X1 U266bar ( .A1(n694bar), .A2(n693bar), .ZN(n695bar);
  OR2_X1 U267 ( .A1(in[121]), .A2(in[102]), .ZN(n693) );
  AND2_X1 U267bar ( .A1(inbar[121]), .A2(inbar[102]), .ZN(n693bar);
  OR2_X1 U268 ( .A1(in[162]), .A2(in[161]), .ZN(n694) );
  AND2_X1 U268bar ( .A1(inbar[162]), .A2(inbar[161]), .ZN(n694bar);
  OR2_X1 U269 ( .A1(n692), .A2(n691), .ZN(n696) );
  AND2_X1 U269bar ( .A1(n692bar), .A2(n691bar), .ZN(n696bar);
  OR2_X1 U270 ( .A1(in[192]), .A2(in[178]), .ZN(n691) );
  AND2_X1 U270bar ( .A1(inbar[192]), .A2(inbar[178]), .ZN(n691bar);
  OR2_X1 U271 ( .A1(in[244]), .A2(in[209]), .ZN(n692) );
  AND2_X1 U271bar ( .A1(inbar[244]), .A2(inbar[209]), .ZN(n692bar);
  OR2_X1 U272 ( .A1(n690), .A2(n689), .ZN(n698) );
  AND2_X1 U272bar ( .A1(n690bar), .A2(n689bar), .ZN(n698bar);
  OR2_X1 U273 ( .A1(n688), .A2(n687), .ZN(n689) );
  AND2_X1 U273bar ( .A1(n688bar), .A2(n687bar), .ZN(n689bar);
  OR2_X1 U274 ( .A1(in[90]), .A2(in[254]), .ZN(n687) );
  AND2_X1 U274bar ( .A1(inbar[90]), .A2(inbar[254]), .ZN(n687bar);
  OR2_X1 U275 ( .A1(in_36), .A2(in_32), .ZN(n688) );
  AND2_X1 U275bar ( .A1(in_36bar), .A2(in_32bar), .ZN(n688bar);
  OR2_X1 U276 ( .A1(n686), .A2(n685), .ZN(n690) );
  AND2_X1 U276bar ( .A1(n686bar), .A2(n685bar), .ZN(n690bar);
  OR2_X1 U277 ( .A1(in_62), .A2(in_37), .ZN(n685) );
  AND2_X1 U277bar ( .A1(in_62bar), .A2(in_37bar), .ZN(n685bar);
  OR2_X1 U278 ( .A1(in_75), .A2(in_73), .ZN(n686) );
  AND2_X1 U278bar ( .A1(in_75bar), .A2(in_73bar), .ZN(n686bar);
  OR2_X1 U279 ( .A1(n684), .A2(n683), .ZN(n944) );
  AND2_X1 U279bar ( .A1(n684bar), .A2(n683bar), .ZN(n944bar);
  OR2_X1 U280 ( .A1(n682), .A2(n681), .ZN(n683) );
  AND2_X1 U280bar ( .A1(n682bar), .A2(n681bar), .ZN(n683bar);
  OR2_X1 U281 ( .A1(n680), .A2(n679), .ZN(n681) );
  AND2_X1 U281bar ( .A1(n680bar), .A2(n679bar), .ZN(n681bar);
  OR2_X1 U282 ( .A1(in[171]), .A2(in[153]), .ZN(n679) );
  AND2_X1 U282bar ( .A1(inbar[171]), .A2(inbar[153]), .ZN(n679bar);
  OR2_X1 U283 ( .A1(in[187]), .A2(in[176]), .ZN(n680) );
  AND2_X1 U283bar ( .A1(inbar[187]), .A2(inbar[176]), .ZN(n680bar);
  OR2_X1 U284 ( .A1(n678), .A2(n677), .ZN(n682) );
  AND2_X1 U284bar ( .A1(n678bar), .A2(n677bar), .ZN(n682bar);
  OR2_X1 U285 ( .A1(in[245]), .A2(in[211]), .ZN(n677) );
  AND2_X1 U285bar ( .A1(inbar[245]), .A2(inbar[211]), .ZN(n677bar);
  OR2_X1 U286 ( .A1(in[97]), .A2(in[88]), .ZN(n678) );
  AND2_X1 U286bar ( .A1(inbar[97]), .A2(inbar[88]), .ZN(n678bar);
  OR2_X1 U287 ( .A1(n676), .A2(n675), .ZN(n684) );
  AND2_X1 U287bar ( .A1(n676bar), .A2(n675bar), .ZN(n684bar);
  OR2_X1 U288 ( .A1(n674), .A2(n673), .ZN(n675) );
  AND2_X1 U288bar ( .A1(n674bar), .A2(n673bar), .ZN(n675bar);
  OR2_X1 U289 ( .A1(in_10), .A2(in_0), .ZN(n673) );
  AND2_X1 U289bar ( .A1(in_10bar), .A2(in_0bar), .ZN(n673bar);
  OR2_X1 U290 ( .A1(in_59), .A2(in_5), .ZN(n674) );
  AND2_X1 U290bar ( .A1(in_59bar), .A2(in_5bar), .ZN(n674bar);
  OR2_X1 U291 ( .A1(n672), .A2(n671), .ZN(n676) );
  AND2_X1 U291bar ( .A1(n672bar), .A2(n671bar), .ZN(n676bar);
  OR2_X1 U292 ( .A1(in_60), .A2(in_6), .ZN(n671) );
  AND2_X1 U292bar ( .A1(in_60bar), .A2(in_6bar), .ZN(n671bar);
  OR2_X1 U293 ( .A1(in_77), .A2(in_69), .ZN(n672) );
  AND2_X1 U293bar ( .A1(in_77bar), .A2(in_69bar), .ZN(n672bar);
  OR2_X1 U294 ( .A1(in[113]), .A2(n864), .ZN(n700) );
  AND2_X1 U294bar ( .A1(inbar[113]), .A2(n864bar), .ZN(n700bar);
  OR2_X1 U295 ( .A1(n670), .A2(n669), .ZN(n864) );
  AND2_X1 U295bar ( .A1(n670bar), .A2(n669bar), .ZN(n864bar);
  OR2_X1 U296 ( .A1(n668), .A2(n667), .ZN(n669) );
  AND2_X1 U296bar ( .A1(n668bar), .A2(n667bar), .ZN(n669bar);
  OR2_X1 U297 ( .A1(n666), .A2(n665), .ZN(n667) );
  AND2_X1 U297bar ( .A1(n666bar), .A2(n665bar), .ZN(n667bar);
  OR2_X1 U298 ( .A1(in[125]), .A2(in[107]), .ZN(n665) );
  AND2_X1 U298bar ( .A1(inbar[125]), .A2(inbar[107]), .ZN(n665bar);
  OR2_X1 U299 ( .A1(in[138]), .A2(in[126]), .ZN(n666) );
  AND2_X1 U299bar ( .A1(inbar[138]), .A2(inbar[126]), .ZN(n666bar);
  OR2_X1 U300 ( .A1(n664), .A2(n663), .ZN(n668) );
  AND2_X1 U300bar ( .A1(n664bar), .A2(n663bar), .ZN(n668bar);
  OR2_X1 U301 ( .A1(in[189]), .A2(in[143]), .ZN(n663) );
  AND2_X1 U301bar ( .A1(inbar[189]), .A2(inbar[143]), .ZN(n663bar);
  OR2_X1 U302 ( .A1(in[99]), .A2(in[214]), .ZN(n664) );
  AND2_X1 U302bar ( .A1(inbar[99]), .A2(inbar[214]), .ZN(n664bar);
  OR2_X1 U303 ( .A1(n662), .A2(n661), .ZN(n670) );
  AND2_X1 U303bar ( .A1(n662bar), .A2(n661bar), .ZN(n670bar);
  OR2_X1 U304 ( .A1(n660), .A2(n659), .ZN(n661) );
  AND2_X1 U304bar ( .A1(n660bar), .A2(n659bar), .ZN(n661bar);
  OR2_X1 U305 ( .A1(in_15), .A2(in_12), .ZN(n659) );
  AND2_X1 U305bar ( .A1(in_15bar), .A2(in_12bar), .ZN(n659bar);
  OR2_X1 U306 ( .A1(in_20), .A2(in_2), .ZN(n660) );
  AND2_X1 U306bar ( .A1(in_20bar), .A2(in_2bar), .ZN(n660bar);
  OR2_X1 U307 ( .A1(n658), .A2(n657), .ZN(n662) );
  AND2_X1 U307bar ( .A1(n658bar), .A2(n657bar), .ZN(n662bar);
  OR2_X1 U308 ( .A1(in_30), .A2(in_3), .ZN(n657) );
  AND2_X1 U308bar ( .A1(in_30bar), .A2(in_3bar), .ZN(n657bar);
  OR2_X1 U309 ( .A1(in_4), .A2(in_38), .ZN(n658) );
  AND2_X1 U309bar ( .A1(in_4bar), .A2(in_38bar), .ZN(n658bar);
  OR2_X1 U310 ( .A1(n656), .A2(n655), .ZN(n702) );
  AND2_X1 U310bar ( .A1(n656bar), .A2(n655bar), .ZN(n702bar);
  OR2_X1 U311 ( .A1(in[148]), .A2(in[137]), .ZN(n655) );
  AND2_X1 U311bar ( .A1(inbar[148]), .A2(inbar[137]), .ZN(n655bar);
  OR2_X1 U312 ( .A1(in[149]), .A2(n654), .ZN(n656) );
  AND2_X1 U312bar ( .A1(inbar[149]), .A2(n654bar), .ZN(n656bar);
  OR2_X1 U313 ( .A1(in[195]), .A2(in[190]), .ZN(n654) );
  AND2_X1 U313bar ( .A1(inbar[195]), .A2(inbar[190]), .ZN(n654bar);
  OR2_X1 U314 ( .A1(n653), .A2(n652), .ZN(n704) );
  AND2_X1 U314bar ( .A1(n653bar), .A2(n652bar), .ZN(n704bar);
  OR2_X1 U315 ( .A1(n651), .A2(n650), .ZN(n652) );
  AND2_X1 U315bar ( .A1(n651bar), .A2(n650bar), .ZN(n652bar);
  OR2_X1 U316 ( .A1(in[98]), .A2(in[197]), .ZN(n650) );
  AND2_X1 U316bar ( .A1(inbar[98]), .A2(inbar[197]), .ZN(n650bar);
  OR2_X1 U317 ( .A1(in_11), .A2(n649), .ZN(n651) );
  AND2_X1 U317bar ( .A1(in_11bar), .A2(n649bar), .ZN(n651bar);
  OR2_X1 U318 ( .A1(in_26), .A2(in_14), .ZN(n649) );
  AND2_X1 U318bar ( .A1(in_26bar), .A2(in_14bar), .ZN(n649bar);
  OR2_X1 U319 ( .A1(n648), .A2(n647), .ZN(n653) );
  AND2_X1 U319bar ( .A1(n648bar), .A2(n647bar), .ZN(n653bar);
  OR2_X1 U320 ( .A1(in_35), .A2(in_27), .ZN(n647) );
  AND2_X1 U320bar ( .A1(in_35bar), .A2(in_27bar), .ZN(n647bar);
  OR2_X1 U321 ( .A1(in_50), .A2(n646), .ZN(n648) );
  AND2_X1 U321bar ( .A1(in_50bar), .A2(n646bar), .ZN(n648bar);
  OR2_X1 U322 ( .A1(in_78), .A2(in_61), .ZN(n646) );
  AND2_X1 U322bar ( .A1(in_78bar), .A2(in_61bar), .ZN(n646bar);
  OR2_X1 U323 ( .A1(n942), .A2(n645), .ZN(n720) );
  AND2_X1 U323bar ( .A1(n942bar), .A2(n645bar), .ZN(n720bar);
  OR2_X1 U324 ( .A1(in[106]), .A2(n863), .ZN(n645) );
  AND2_X1 U324bar ( .A1(inbar[106]), .A2(n863bar), .ZN(n645bar);
  OR2_X1 U325 ( .A1(n644), .A2(n643), .ZN(n863) );
  AND2_X1 U325bar ( .A1(n644bar), .A2(n643bar), .ZN(n863bar);
  OR2_X1 U326 ( .A1(n642), .A2(n641), .ZN(n643) );
  AND2_X1 U326bar ( .A1(n642bar), .A2(n641bar), .ZN(n643bar);
  OR2_X1 U327 ( .A1(n640), .A2(n639), .ZN(n641) );
  AND2_X1 U327bar ( .A1(n640bar), .A2(n639bar), .ZN(n641bar);
  OR2_X1 U328 ( .A1(in[127]), .A2(in[122]), .ZN(n639) );
  AND2_X1 U328bar ( .A1(inbar[127]), .A2(inbar[122]), .ZN(n639bar);
  OR2_X1 U329 ( .A1(in[156]), .A2(in[132]), .ZN(n640) );
  AND2_X1 U329bar ( .A1(inbar[156]), .A2(inbar[132]), .ZN(n640bar);
  OR2_X1 U330 ( .A1(n638), .A2(n637), .ZN(n642) );
  AND2_X1 U330bar ( .A1(n638bar), .A2(n637bar), .ZN(n642bar);
  OR2_X1 U331 ( .A1(in[159]), .A2(in[157]), .ZN(n637) );
  AND2_X1 U331bar ( .A1(inbar[159]), .A2(inbar[157]), .ZN(n637bar);
  OR2_X1 U332 ( .A1(in[185]), .A2(in[169]), .ZN(n638) );
  AND2_X1 U332bar ( .A1(inbar[185]), .A2(inbar[169]), .ZN(n638bar);
  OR2_X1 U333 ( .A1(n636), .A2(n635), .ZN(n644) );
  AND2_X1 U333bar ( .A1(n636bar), .A2(n635bar), .ZN(n644bar);
  OR2_X1 U334 ( .A1(n634), .A2(n633), .ZN(n635) );
  AND2_X1 U334bar ( .A1(n634bar), .A2(n633bar), .ZN(n635bar);
  OR2_X1 U335 ( .A1(in[239]), .A2(in[218]), .ZN(n633) );
  AND2_X1 U335bar ( .A1(inbar[239]), .A2(inbar[218]), .ZN(n633bar);
  OR2_X1 U336 ( .A1(in_13), .A2(in[87]), .ZN(n634) );
  AND2_X1 U336bar ( .A1(in_13bar), .A2(inbar[87]), .ZN(n634bar);
  OR2_X1 U337 ( .A1(n632), .A2(n631), .ZN(n636) );
  AND2_X1 U337bar ( .A1(n632bar), .A2(n631bar), .ZN(n636bar);
  OR2_X1 U338 ( .A1(in_72), .A2(in_70), .ZN(n631) );
  AND2_X1 U338bar ( .A1(in_72bar), .A2(in_70bar), .ZN(n631bar);
  OR2_X1 U339 ( .A1(in_80), .A2(in_74), .ZN(n632) );
  AND2_X1 U339bar ( .A1(in_80bar), .A2(in_74bar), .ZN(n632bar);
  OR2_X1 U340 ( .A1(n630), .A2(n629), .ZN(n942) );
  AND2_X1 U340bar ( .A1(n630bar), .A2(n629bar), .ZN(n942bar);
  OR2_X1 U341 ( .A1(n628), .A2(n627), .ZN(n629) );
  AND2_X1 U341bar ( .A1(n628bar), .A2(n627bar), .ZN(n629bar);
  OR2_X1 U342 ( .A1(n626), .A2(n625), .ZN(n627) );
  AND2_X1 U342bar ( .A1(n626bar), .A2(n625bar), .ZN(n627bar);
  OR2_X1 U343 ( .A1(in[146]), .A2(in[100]), .ZN(n625) );
  AND2_X1 U343bar ( .A1(inbar[146]), .A2(inbar[100]), .ZN(n625bar);
  OR2_X1 U344 ( .A1(in[168]), .A2(in[152]), .ZN(n626) );
  AND2_X1 U344bar ( .A1(inbar[168]), .A2(inbar[152]), .ZN(n626bar);
  OR2_X1 U345 ( .A1(n624), .A2(n623), .ZN(n628) );
  AND2_X1 U345bar ( .A1(n624bar), .A2(n623bar), .ZN(n628bar);
  OR2_X1 U346 ( .A1(in[199]), .A2(in[182]), .ZN(n623) );
  AND2_X1 U346bar ( .A1(inbar[199]), .A2(inbar[182]), .ZN(n623bar);
  OR2_X1 U347 ( .A1(in[236]), .A2(in[204]), .ZN(n624) );
  AND2_X1 U347bar ( .A1(inbar[236]), .A2(inbar[204]), .ZN(n624bar);
  OR2_X1 U348 ( .A1(n622), .A2(n621), .ZN(n630) );
  AND2_X1 U348bar ( .A1(n622bar), .A2(n621bar), .ZN(n630bar);
  OR2_X1 U349 ( .A1(n620), .A2(n619), .ZN(n621) );
  AND2_X1 U349bar ( .A1(n620bar), .A2(n619bar), .ZN(n621bar);
  OR2_X1 U350 ( .A1(in[89]), .A2(in[246]), .ZN(n619) );
  AND2_X1 U350bar ( .A1(inbar[89]), .A2(inbar[246]), .ZN(n619bar);
  OR2_X1 U351 ( .A1(in[95]), .A2(in[92]), .ZN(n620) );
  AND2_X1 U351bar ( .A1(inbar[95]), .A2(inbar[92]), .ZN(n620bar);
  OR2_X1 U352 ( .A1(n618), .A2(n617), .ZN(n622) );
  AND2_X1 U352bar ( .A1(n618bar), .A2(n617bar), .ZN(n622bar);
  OR2_X1 U353 ( .A1(in_22), .A2(in_16), .ZN(n617) );
  AND2_X1 U353bar ( .A1(in_22bar), .A2(in_16bar), .ZN(n617bar);
  OR2_X1 U354 ( .A1(in_51), .A2(in_49), .ZN(n618) );
  AND2_X1 U354bar ( .A1(in_51bar), .A2(in_49bar), .ZN(n618bar);
  OR2_X1 U355 ( .A1(n616), .A2(n615), .ZN(n722) );
  AND2_X1 U355bar ( .A1(n616bar), .A2(n615bar), .ZN(n722bar);
  OR2_X1 U356 ( .A1(in[158]), .A2(in[115]), .ZN(n615) );
  AND2_X1 U356bar ( .A1(inbar[158]), .A2(inbar[115]), .ZN(n615bar);
  OR2_X1 U357 ( .A1(in[163]), .A2(n614), .ZN(n616) );
  AND2_X1 U357bar ( .A1(inbar[163]), .A2(n614bar), .ZN(n616bar);
  OR2_X1 U358 ( .A1(in[206]), .A2(in[165]), .ZN(n614) );
  AND2_X1 U358bar ( .A1(inbar[206]), .A2(inbar[165]), .ZN(n614bar);
  OR2_X1 U359 ( .A1(n613), .A2(n612), .ZN(n724) );
  AND2_X1 U359bar ( .A1(n613bar), .A2(n612bar), .ZN(n724bar);
  OR2_X1 U360 ( .A1(n611), .A2(n610), .ZN(n612) );
  AND2_X1 U360bar ( .A1(n611bar), .A2(n610bar), .ZN(n612bar);
  OR2_X1 U361 ( .A1(in[213]), .A2(in[207]), .ZN(n610) );
  AND2_X1 U361bar ( .A1(inbar[213]), .A2(inbar[207]), .ZN(n610bar);
  OR2_X1 U362 ( .A1(in[215]), .A2(n609), .ZN(n611) );
  AND2_X1 U362bar ( .A1(inbar[215]), .A2(n609bar), .ZN(n611bar);
  OR2_X1 U363 ( .A1(in[230]), .A2(in[220]), .ZN(n609) );
  AND2_X1 U363bar ( .A1(inbar[230]), .A2(inbar[220]), .ZN(n609bar);
  OR2_X1 U364 ( .A1(n608), .A2(n607), .ZN(n613) );
  AND2_X1 U364bar ( .A1(n608bar), .A2(n607bar), .ZN(n613bar);
  OR2_X1 U365 ( .A1(in[251]), .A2(in[234]), .ZN(n607) );
  AND2_X1 U365bar ( .A1(inbar[251]), .A2(inbar[234]), .ZN(n607bar);
  OR2_X1 U366 ( .A1(in_17), .A2(n606), .ZN(n608) );
  AND2_X1 U366bar ( .A1(in_17bar), .A2(n606bar), .ZN(n608bar);
  OR2_X1 U367 ( .A1(in_65), .A2(in_56), .ZN(n606) );
  AND2_X1 U367bar ( .A1(in_65bar), .A2(in_56bar), .ZN(n606bar);
  OR2_X1 U368 ( .A1(n605), .A2(n604), .ZN(out[0]) );
  AND2_X1 U368bar ( .A1(n605bar), .A2(n604bar), .ZN(outbar[0]);
  OR2_X1 U369 ( .A1(n603), .A2(n602), .ZN(n604) );
  AND2_X1 U369bar ( .A1(n603bar), .A2(n602bar), .ZN(n604bar);
  OR2_X1 U370 ( .A1(n601), .A2(n600), .ZN(n602) );
  AND2_X1 U370bar ( .A1(n601bar), .A2(n600bar), .ZN(n602bar);
  OR2_X1 U371 ( .A1(n820), .A2(n785), .ZN(n600) );
  AND2_X1 U371bar ( .A1(n820bar), .A2(n785bar), .ZN(n600bar);
  OR2_X1 U372 ( .A1(n599), .A2(n598), .ZN(n785) );
  AND2_X1 U372bar ( .A1(n599bar), .A2(n598bar), .ZN(n785bar);
  OR2_X1 U373 ( .A1(n597), .A2(n596), .ZN(n598) );
  AND2_X1 U373bar ( .A1(n597bar), .A2(n596bar), .ZN(n598bar);
  OR2_X1 U374 ( .A1(n595), .A2(n594), .ZN(n596) );
  AND2_X1 U374bar ( .A1(n595bar), .A2(n594bar), .ZN(n596bar);
  OR2_X1 U375 ( .A1(in[135]), .A2(in[104]), .ZN(n594) );
  AND2_X1 U375bar ( .A1(inbar[135]), .A2(inbar[104]), .ZN(n594bar);
  OR2_X1 U376 ( .A1(in[188]), .A2(in[178]), .ZN(n595) );
  AND2_X1 U376bar ( .A1(inbar[188]), .A2(inbar[178]), .ZN(n595bar);
  OR2_X1 U377 ( .A1(n593), .A2(n592), .ZN(n597) );
  AND2_X1 U377bar ( .A1(n593bar), .A2(n592bar), .ZN(n597bar);
  OR2_X1 U378 ( .A1(in[217]), .A2(in[194]), .ZN(n592) );
  AND2_X1 U378bar ( .A1(inbar[217]), .A2(inbar[194]), .ZN(n592bar);
  OR2_X1 U379 ( .A1(in[237]), .A2(in[218]), .ZN(n593) );
  AND2_X1 U379bar ( .A1(inbar[237]), .A2(inbar[218]), .ZN(n593bar);
  OR2_X1 U380 ( .A1(n591), .A2(n590), .ZN(n599) );
  AND2_X1 U380bar ( .A1(n591bar), .A2(n590bar), .ZN(n599bar);
  OR2_X1 U381 ( .A1(n589), .A2(n588), .ZN(n590) );
  AND2_X1 U381bar ( .A1(n589bar), .A2(n588bar), .ZN(n590bar);
  OR2_X1 U382 ( .A1(in_2), .A2(in_10), .ZN(n588) );
  AND2_X1 U382bar ( .A1(in_2bar), .A2(in_10bar), .ZN(n588bar);
  OR2_X1 U383 ( .A1(in_47), .A2(in_22), .ZN(n589) );
  AND2_X1 U383bar ( .A1(in_47bar), .A2(in_22bar), .ZN(n589bar);
  OR2_X1 U384 ( .A1(n587), .A2(n586), .ZN(n591) );
  AND2_X1 U384bar ( .A1(n587bar), .A2(n586bar), .ZN(n591bar);
  OR2_X1 U385 ( .A1(in_56), .A2(in_54), .ZN(n586) );
  AND2_X1 U385bar ( .A1(in_56bar), .A2(in_54bar), .ZN(n586bar);
  OR2_X1 U386 ( .A1(in_63), .A2(in_61), .ZN(n587) );
  AND2_X1 U386bar ( .A1(in_63bar), .A2(in_61bar), .ZN(n587bar);
  OR2_X1 U387 ( .A1(n585), .A2(n584), .ZN(n820) );
  AND2_X1 U387bar ( .A1(n585bar), .A2(n584bar), .ZN(n820bar);
  OR2_X1 U388 ( .A1(n583), .A2(n582), .ZN(n584) );
  AND2_X1 U388bar ( .A1(n583bar), .A2(n582bar), .ZN(n584bar);
  OR2_X1 U389 ( .A1(n581), .A2(n580), .ZN(n582) );
  AND2_X1 U389bar ( .A1(n581bar), .A2(n580bar), .ZN(n582bar);
  OR2_X1 U390 ( .A1(in[158]), .A2(in[142]), .ZN(n580) );
  AND2_X1 U390bar ( .A1(inbar[158]), .A2(inbar[142]), .ZN(n580bar);
  OR2_X1 U391 ( .A1(in[175]), .A2(in[164]), .ZN(n581) );
  AND2_X1 U391bar ( .A1(inbar[175]), .A2(inbar[164]), .ZN(n581bar);
  OR2_X1 U392 ( .A1(n579), .A2(n578), .ZN(n583) );
  AND2_X1 U392bar ( .A1(n579bar), .A2(n578bar), .ZN(n583bar);
  OR2_X1 U393 ( .A1(in[228]), .A2(in[204]), .ZN(n578) );
  AND2_X1 U393bar ( .A1(inbar[228]), .A2(inbar[204]), .ZN(n578bar);
  OR2_X1 U394 ( .A1(in[91]), .A2(in[87]), .ZN(n579) );
  AND2_X1 U394bar ( .A1(inbar[91]), .A2(inbar[87]), .ZN(n579bar);
  OR2_X1 U395 ( .A1(n577), .A2(n576), .ZN(n585) );
  AND2_X1 U395bar ( .A1(n577bar), .A2(n576bar), .ZN(n585bar);
  OR2_X1 U396 ( .A1(n575), .A2(n574), .ZN(n576) );
  AND2_X1 U396bar ( .A1(n575bar), .A2(n574bar), .ZN(n576bar);
  OR2_X1 U397 ( .A1(in_21), .A2(in_11), .ZN(n574) );
  AND2_X1 U397bar ( .A1(in_21bar), .A2(in_11bar), .ZN(n574bar);
  OR2_X1 U398 ( .A1(in_5), .A2(in_3), .ZN(n575) );
  AND2_X1 U398bar ( .A1(in_5bar), .A2(in_3bar), .ZN(n575bar);
  OR2_X1 U399 ( .A1(n573), .A2(n572), .ZN(n577) );
  AND2_X1 U399bar ( .A1(n573bar), .A2(n572bar), .ZN(n577bar);
  OR2_X1 U400 ( .A1(in_68), .A2(in_64), .ZN(n572) );
  AND2_X1 U400bar ( .A1(in_68bar), .A2(in_64bar), .ZN(n572bar);
  OR2_X1 U401 ( .A1(in_76), .A2(in_73), .ZN(n573) );
  AND2_X1 U401bar ( .A1(in_76bar), .A2(in_73bar), .ZN(n573bar);
  OR2_X1 U402 ( .A1(n778), .A2(n571), .ZN(n601) );
  AND2_X1 U402bar ( .A1(n778bar), .A2(n571bar), .ZN(n601bar);
  OR2_X1 U403 ( .A1(in[100]), .A2(n965), .ZN(n571) );
  AND2_X1 U403bar ( .A1(inbar[100]), .A2(n965bar), .ZN(n571bar);
  OR2_X1 U404 ( .A1(n570), .A2(n569), .ZN(n965) );
  AND2_X1 U404bar ( .A1(n570bar), .A2(n569bar), .ZN(n965bar);
  OR2_X1 U405 ( .A1(n568), .A2(n567), .ZN(n569) );
  AND2_X1 U405bar ( .A1(n568bar), .A2(n567bar), .ZN(n569bar);
  OR2_X1 U406 ( .A1(n566), .A2(n565), .ZN(n567) );
  AND2_X1 U406bar ( .A1(n566bar), .A2(n565bar), .ZN(n567bar);
  OR2_X1 U407 ( .A1(n817), .A2(n750), .ZN(n565) );
  AND2_X1 U407bar ( .A1(n817bar), .A2(n750bar), .ZN(n565bar);
  OR2_X1 U408 ( .A1(n564), .A2(n563), .ZN(n750) );
  AND2_X1 U408bar ( .A1(n564bar), .A2(n563bar), .ZN(n750bar);
  OR2_X1 U409 ( .A1(n562), .A2(n561), .ZN(n563) );
  AND2_X1 U409bar ( .A1(n562bar), .A2(n561bar), .ZN(n563bar);
  OR2_X1 U410 ( .A1(n560), .A2(n559), .ZN(n561) );
  AND2_X1 U410bar ( .A1(n560bar), .A2(n559bar), .ZN(n561bar);
  OR2_X1 U411 ( .A1(in[119]), .A2(in[103]), .ZN(n559) );
  AND2_X1 U411bar ( .A1(inbar[119]), .A2(inbar[103]), .ZN(n559bar);
  OR2_X1 U412 ( .A1(in[137]), .A2(in[133]), .ZN(n560) );
  AND2_X1 U412bar ( .A1(inbar[137]), .A2(inbar[133]), .ZN(n560bar);
  OR2_X1 U413 ( .A1(n558), .A2(n557), .ZN(n562) );
  AND2_X1 U413bar ( .A1(n558bar), .A2(n557bar), .ZN(n562bar);
  OR2_X1 U414 ( .A1(in[176]), .A2(in[173]), .ZN(n557) );
  AND2_X1 U414bar ( .A1(inbar[176]), .A2(inbar[173]), .ZN(n557bar);
  OR2_X1 U415 ( .A1(in[210]), .A2(in[181]), .ZN(n558) );
  AND2_X1 U415bar ( .A1(inbar[210]), .A2(inbar[181]), .ZN(n558bar);
  OR2_X1 U416 ( .A1(n556), .A2(n555), .ZN(n564) );
  AND2_X1 U416bar ( .A1(n556bar), .A2(n555bar), .ZN(n564bar);
  OR2_X1 U417 ( .A1(n554), .A2(n553), .ZN(n555) );
  AND2_X1 U417bar ( .A1(n554bar), .A2(n553bar), .ZN(n555bar);
  OR2_X1 U418 ( .A1(in_13), .A2(in[234]), .ZN(n553) );
  AND2_X1 U418bar ( .A1(in_13bar), .A2(inbar[234]), .ZN(n553bar);
  OR2_X1 U419 ( .A1(in_38), .A2(in_32), .ZN(n554) );
  AND2_X1 U419bar ( .A1(in_38bar), .A2(in_32bar), .ZN(n554bar);
  OR2_X1 U420 ( .A1(n552), .A2(n551), .ZN(n556) );
  AND2_X1 U420bar ( .A1(n552bar), .A2(n551bar), .ZN(n556bar);
  OR2_X1 U421 ( .A1(in_42), .A2(in_41), .ZN(n551) );
  AND2_X1 U421bar ( .A1(in_42bar), .A2(in_41bar), .ZN(n551bar);
  OR2_X1 U422 ( .A1(in_7), .A2(in_49), .ZN(n552) );
  AND2_X1 U422bar ( .A1(in_7bar), .A2(in_49bar), .ZN(n552bar);
  OR2_X1 U423 ( .A1(n550), .A2(n549), .ZN(n817) );
  AND2_X1 U423bar ( .A1(n550bar), .A2(n549bar), .ZN(n817bar);
  OR2_X1 U424 ( .A1(n548), .A2(n547), .ZN(n549) );
  AND2_X1 U424bar ( .A1(n548bar), .A2(n547bar), .ZN(n549bar);
  OR2_X1 U425 ( .A1(n546), .A2(n545), .ZN(n547) );
  AND2_X1 U425bar ( .A1(n546bar), .A2(n545bar), .ZN(n547bar);
  OR2_X1 U426 ( .A1(in[159]), .A2(in[105]), .ZN(n545) );
  AND2_X1 U426bar ( .A1(inbar[159]), .A2(inbar[105]), .ZN(n545bar);
  OR2_X1 U427 ( .A1(in[206]), .A2(in[183]), .ZN(n546) );
  AND2_X1 U427bar ( .A1(inbar[206]), .A2(inbar[183]), .ZN(n546bar);
  OR2_X1 U428 ( .A1(n544), .A2(n543), .ZN(n548) );
  AND2_X1 U428bar ( .A1(n544bar), .A2(n543bar), .ZN(n548bar);
  OR2_X1 U429 ( .A1(in[229]), .A2(in[219]), .ZN(n543) );
  AND2_X1 U429bar ( .A1(inbar[229]), .A2(inbar[219]), .ZN(n543bar);
  OR2_X1 U430 ( .A1(in[235]), .A2(in[232]), .ZN(n544) );
  AND2_X1 U430bar ( .A1(inbar[235]), .A2(inbar[232]), .ZN(n544bar);
  OR2_X1 U431 ( .A1(n542), .A2(n541), .ZN(n550) );
  AND2_X1 U431bar ( .A1(n542bar), .A2(n541bar), .ZN(n550bar);
  OR2_X1 U432 ( .A1(n540), .A2(n539), .ZN(n541) );
  AND2_X1 U432bar ( .A1(n540bar), .A2(n539bar), .ZN(n541bar);
  OR2_X1 U433 ( .A1(in[249]), .A2(in[242]), .ZN(n539) );
  AND2_X1 U433bar ( .A1(inbar[249]), .A2(inbar[242]), .ZN(n539bar);
  OR2_X1 U434 ( .A1(in[89]), .A2(in[254]), .ZN(n540) );
  AND2_X1 U434bar ( .A1(inbar[89]), .A2(inbar[254]), .ZN(n540bar);
  OR2_X1 U435 ( .A1(n538), .A2(n537), .ZN(n542) );
  AND2_X1 U435bar ( .A1(n538bar), .A2(n537bar), .ZN(n542bar);
  OR2_X1 U436 ( .A1(in_14), .A2(in[99]), .ZN(n537) );
  AND2_X1 U436bar ( .A1(in_14bar), .A2(inbar[99]), .ZN(n537bar);
  OR2_X1 U437 ( .A1(in_60), .A2(in_18), .ZN(n538) );
  AND2_X1 U437bar ( .A1(in_60bar), .A2(in_18bar), .ZN(n538bar);
  OR2_X1 U438 ( .A1(in[113]), .A2(n763), .ZN(n566) );
  AND2_X1 U438bar ( .A1(inbar[113]), .A2(n763bar), .ZN(n566bar);
  OR2_X1 U439 ( .A1(n536), .A2(n535), .ZN(n763) );
  AND2_X1 U439bar ( .A1(n536bar), .A2(n535bar), .ZN(n763bar);
  OR2_X1 U440 ( .A1(n534), .A2(n533), .ZN(n535) );
  AND2_X1 U440bar ( .A1(n534bar), .A2(n533bar), .ZN(n535bar);
  OR2_X1 U441 ( .A1(n532), .A2(n531), .ZN(n533) );
  AND2_X1 U441bar ( .A1(n532bar), .A2(n531bar), .ZN(n533bar);
  OR2_X1 U442 ( .A1(in[115]), .A2(in[110]), .ZN(n531) );
  AND2_X1 U442bar ( .A1(inbar[115]), .A2(inbar[110]), .ZN(n531bar);
  OR2_X1 U443 ( .A1(in[125]), .A2(in[117]), .ZN(n532) );
  AND2_X1 U443bar ( .A1(inbar[125]), .A2(inbar[117]), .ZN(n532bar);
  OR2_X1 U444 ( .A1(n530), .A2(n529), .ZN(n534) );
  AND2_X1 U444bar ( .A1(n530bar), .A2(n529bar), .ZN(n534bar);
  OR2_X1 U445 ( .A1(in[180]), .A2(in[128]), .ZN(n529) );
  AND2_X1 U445bar ( .A1(inbar[180]), .A2(inbar[128]), .ZN(n529bar);
  OR2_X1 U446 ( .A1(in[205]), .A2(in[201]), .ZN(n530) );
  AND2_X1 U446bar ( .A1(inbar[205]), .A2(inbar[201]), .ZN(n530bar);
  OR2_X1 U447 ( .A1(n528), .A2(n527), .ZN(n536) );
  AND2_X1 U447bar ( .A1(n528bar), .A2(n527bar), .ZN(n536bar);
  OR2_X1 U448 ( .A1(n526), .A2(n525), .ZN(n527) );
  AND2_X1 U448bar ( .A1(n526bar), .A2(n525bar), .ZN(n527bar);
  OR2_X1 U449 ( .A1(in[244]), .A2(in[239]), .ZN(n525) );
  AND2_X1 U449bar ( .A1(inbar[244]), .A2(inbar[239]), .ZN(n525bar);
  OR2_X1 U450 ( .A1(in[95]), .A2(in[83]), .ZN(n526) );
  AND2_X1 U450bar ( .A1(inbar[95]), .A2(inbar[83]), .ZN(n526bar);
  OR2_X1 U451 ( .A1(n524), .A2(n523), .ZN(n528) );
  AND2_X1 U451bar ( .A1(n524bar), .A2(n523bar), .ZN(n528bar);
  OR2_X1 U452 ( .A1(in_24), .A2(in[97]), .ZN(n523) );
  AND2_X1 U452bar ( .A1(in_24bar), .A2(inbar[97]), .ZN(n523bar);
  OR2_X1 U453 ( .A1(in_33), .A2(in_27), .ZN(n524) );
  AND2_X1 U453bar ( .A1(in_33bar), .A2(in_27bar), .ZN(n524bar);
  OR2_X1 U454 ( .A1(n522), .A2(n521), .ZN(n568) );
  AND2_X1 U454bar ( .A1(n522bar), .A2(n521bar), .ZN(n568bar);
  OR2_X1 U455 ( .A1(in[145]), .A2(in[126]), .ZN(n521) );
  AND2_X1 U455bar ( .A1(inbar[145]), .A2(inbar[126]), .ZN(n521bar);
  OR2_X1 U456 ( .A1(in[169]), .A2(n520), .ZN(n522) );
  AND2_X1 U456bar ( .A1(inbar[169]), .A2(n520bar), .ZN(n522bar);
  OR2_X1 U457 ( .A1(in[221]), .A2(in[172]), .ZN(n520) );
  AND2_X1 U457bar ( .A1(inbar[221]), .A2(inbar[172]), .ZN(n520bar);
  OR2_X1 U458 ( .A1(n519), .A2(n518), .ZN(n570) );
  AND2_X1 U458bar ( .A1(n519bar), .A2(n518bar), .ZN(n570bar);
  OR2_X1 U459 ( .A1(n517), .A2(n516), .ZN(n518) );
  AND2_X1 U459bar ( .A1(n517bar), .A2(n516bar), .ZN(n518bar);
  OR2_X1 U460 ( .A1(in[241]), .A2(in[224]), .ZN(n516) );
  AND2_X1 U460bar ( .A1(inbar[241]), .A2(inbar[224]), .ZN(n516bar);
  OR2_X1 U461 ( .A1(in[86]), .A2(n515), .ZN(n517) );
  AND2_X1 U461bar ( .A1(inbar[86]), .A2(n515bar), .ZN(n517bar);
  OR2_X1 U462 ( .A1(in_43), .A2(in_34), .ZN(n515) );
  AND2_X1 U462bar ( .A1(in_43bar), .A2(in_34bar), .ZN(n515bar);
  OR2_X1 U463 ( .A1(n514), .A2(n513), .ZN(n519) );
  AND2_X1 U463bar ( .A1(n514bar), .A2(n513bar), .ZN(n519bar);
  OR2_X1 U464 ( .A1(in_65), .A2(in_51), .ZN(n513) );
  AND2_X1 U464bar ( .A1(in_65bar), .A2(in_51bar), .ZN(n513bar);
  OR2_X1 U465 ( .A1(in_75), .A2(n512), .ZN(n514) );
  AND2_X1 U465bar ( .A1(in_75bar), .A2(n512bar), .ZN(n514bar);
  OR2_X1 U466 ( .A1(in_81), .A2(in_77), .ZN(n512) );
  AND2_X1 U466bar ( .A1(in_81bar), .A2(in_77bar), .ZN(n512bar);
  OR2_X1 U467 ( .A1(n511), .A2(n510), .ZN(n778) );
  AND2_X1 U467bar ( .A1(n511bar), .A2(n510bar), .ZN(n778bar);
  OR2_X1 U468 ( .A1(n509), .A2(n508), .ZN(n510) );
  AND2_X1 U468bar ( .A1(n509bar), .A2(n508bar), .ZN(n510bar);
  OR2_X1 U469 ( .A1(n507), .A2(n506), .ZN(n508) );
  AND2_X1 U469bar ( .A1(n507bar), .A2(n506bar), .ZN(n508bar);
  OR2_X1 U470 ( .A1(in[107]), .A2(in[101]), .ZN(n506) );
  AND2_X1 U470bar ( .A1(inbar[107]), .A2(inbar[101]), .ZN(n506bar);
  OR2_X1 U471 ( .A1(in[139]), .A2(in[132]), .ZN(n507) );
  AND2_X1 U471bar ( .A1(inbar[139]), .A2(inbar[132]), .ZN(n507bar);
  OR2_X1 U472 ( .A1(n505), .A2(n504), .ZN(n509) );
  AND2_X1 U472bar ( .A1(n505bar), .A2(n504bar), .ZN(n509bar);
  OR2_X1 U473 ( .A1(in[146]), .A2(in[141]), .ZN(n504) );
  AND2_X1 U473bar ( .A1(inbar[146]), .A2(inbar[141]), .ZN(n504bar);
  OR2_X1 U474 ( .A1(in[203]), .A2(in[179]), .ZN(n505) );
  AND2_X1 U474bar ( .A1(inbar[203]), .A2(inbar[179]), .ZN(n505bar);
  OR2_X1 U475 ( .A1(n503), .A2(n502), .ZN(n511) );
  AND2_X1 U475bar ( .A1(n503bar), .A2(n502bar), .ZN(n511bar);
  OR2_X1 U476 ( .A1(n501), .A2(n500), .ZN(n502) );
  AND2_X1 U476bar ( .A1(n501bar), .A2(n500bar), .ZN(n502bar);
  OR2_X1 U477 ( .A1(in[243]), .A2(in[222]), .ZN(n500) );
  AND2_X1 U477bar ( .A1(inbar[243]), .A2(inbar[222]), .ZN(n500bar);
  OR2_X1 U478 ( .A1(in[251]), .A2(in[250]), .ZN(n501) );
  AND2_X1 U478bar ( .A1(inbar[251]), .A2(inbar[250]), .ZN(n501bar);
  OR2_X1 U479 ( .A1(n499), .A2(n498), .ZN(n503) );
  AND2_X1 U479bar ( .A1(n499bar), .A2(n498bar), .ZN(n503bar);
  OR2_X1 U480 ( .A1(in_37), .A2(in_19), .ZN(n498) );
  AND2_X1 U480bar ( .A1(in_37bar), .A2(in_19bar), .ZN(n498bar);
  OR2_X1 U481 ( .A1(in_78), .A2(in_6), .ZN(n499) );
  AND2_X1 U481bar ( .A1(in_78bar), .A2(in_6bar), .ZN(n499bar);
  OR2_X1 U482 ( .A1(n497), .A2(n496), .ZN(n603) );
  AND2_X1 U482bar ( .A1(n497bar), .A2(n496bar), .ZN(n603bar);
  OR2_X1 U483 ( .A1(in[112]), .A2(in[102]), .ZN(n496) );
  AND2_X1 U483bar ( .A1(inbar[112]), .A2(inbar[102]), .ZN(n496bar);
  OR2_X1 U484 ( .A1(in[123]), .A2(n495), .ZN(n497) );
  AND2_X1 U484bar ( .A1(inbar[123]), .A2(n495bar), .ZN(n497bar);
  OR2_X1 U485 ( .A1(in[143]), .A2(in[130]), .ZN(n495) );
  AND2_X1 U485bar ( .A1(inbar[143]), .A2(inbar[130]), .ZN(n495bar);
  OR2_X1 U486 ( .A1(n494), .A2(n493), .ZN(n605) );
  AND2_X1 U486bar ( .A1(n494bar), .A2(n493bar), .ZN(n605bar);
  OR2_X1 U487 ( .A1(n492), .A2(n491), .ZN(n493) );
  AND2_X1 U487bar ( .A1(n492bar), .A2(n491bar), .ZN(n493bar);
  OR2_X1 U488 ( .A1(in[216]), .A2(in[213]), .ZN(n491) );
  AND2_X1 U488bar ( .A1(inbar[216]), .A2(inbar[213]), .ZN(n491bar);
  OR2_X1 U489 ( .A1(in[227]), .A2(n490), .ZN(n492) );
  AND2_X1 U489bar ( .A1(inbar[227]), .A2(n490bar), .ZN(n492bar);
  OR2_X1 U490 ( .A1(in_0), .A2(in[248]), .ZN(n490) );
  AND2_X1 U490bar ( .A1(in_0bar), .A2(inbar[248]), .ZN(n490bar);
  OR2_X1 U491 ( .A1(n489), .A2(n488), .ZN(n494) );
  AND2_X1 U491bar ( .A1(n489bar), .A2(n488bar), .ZN(n494bar);
  OR2_X1 U492 ( .A1(in_46), .A2(in_44), .ZN(n488) );
  AND2_X1 U492bar ( .A1(in_46bar), .A2(in_44bar), .ZN(n488bar);
  OR2_X1 U493 ( .A1(in_50), .A2(n487), .ZN(n489) );
  AND2_X1 U493bar ( .A1(in_50bar), .A2(n487bar), .ZN(n489bar);
  OR2_X1 U494 ( .A1(in_9), .A2(in_80), .ZN(n487) );
  AND2_X1 U494bar ( .A1(in_9bar), .A2(in_80bar), .ZN(n487bar);
endmodule




module sBox_16 ( in, out );
  input [7:0] in;
  //input_done

  output [7:0] out;
  //output_done

  wire   [255:0] decodeOut;
  //wire_done

  decode_16 dec ( .in(in), .out(decodeOut) );
  encode_16 enc ( .in(decodeOut), .out(out) );
endmodule


module CD2_65 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_66 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_67 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_68 ( a, b, y );
 input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD4_33 ( a, b, y );
  input [3:0] a;
  input [3:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  //input_done

  output [15:0] y;
  reg [15:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]);
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]);
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]);
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]);
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]);
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]);
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]);
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]);
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]);
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]);
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]);
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]);
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]);
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]);
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]);
endmodule




module CD4_34 ( a, b, y );
  input [3:0] a;
  input [3:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  //input_done

  output [15:0] y;
  reg [15:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]);
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]);
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]);
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]);
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]);
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]);
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]);
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]);
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]);
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]);
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]);
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]);
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]);
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]);
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]);
endmodule




module CD16_17 ( a, b, y );
  input [15:0] a;
  input [15:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign abar[8] = ~a[8];
  assign abar[9] = ~a[9];
  assign abar[10] = ~a[10];
  assign abar[11] = ~a[11];
  assign abar[12] = ~a[12];
  assign abar[13] = ~a[13];
  assign abar[14] = ~a[14];
  assign abar[15] = ~a[15];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign bbar[8] = ~b[8];
  assign bbar[9] = ~b[9];
  assign bbar[10] = ~b[10];
  assign bbar[11] = ~b[11];
  assign bbar[12] = ~b[12];
  assign bbar[13] = ~b[13];
  assign bbar[14] = ~b[14];
  assign bbar[15] = ~b[15];
  //input_done

  output [15:0] y;
  reg [15:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[9]), .A2(a[0]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[9]), .A2(abar[0]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[3]), .A2(a[6]), .ZN(y[99]) );
  OR2_X1 U2bar ( .A1(bbar[3]), .A2(abar[6]), .ZN(ybar[99]);
  AND2_X1 U3 ( .A1(b[2]), .A2(a[6]), .ZN(y[98]) );
  OR2_X1 U3bar ( .A1(bbar[2]), .A2(abar[6]), .ZN(ybar[98]);
  AND2_X1 U4 ( .A1(b[1]), .A2(a[6]), .ZN(y[97]) );
  OR2_X1 U4bar ( .A1(bbar[1]), .A2(abar[6]), .ZN(ybar[97]);
  AND2_X1 U5 ( .A1(b[0]), .A2(a[6]), .ZN(y[96]) );
  OR2_X1 U5bar ( .A1(bbar[0]), .A2(abar[6]), .ZN(ybar[96]);
  AND2_X1 U6 ( .A1(b[15]), .A2(a[5]), .ZN(y[95]) );
  OR2_X1 U6bar ( .A1(bbar[15]), .A2(abar[5]), .ZN(ybar[95]);
  AND2_X1 U7 ( .A1(b[14]), .A2(a[5]), .ZN(y[94]) );
  OR2_X1 U7bar ( .A1(bbar[14]), .A2(abar[5]), .ZN(ybar[94]);
  AND2_X1 U8 ( .A1(b[13]), .A2(a[5]), .ZN(y[93]) );
  OR2_X1 U8bar ( .A1(bbar[13]), .A2(abar[5]), .ZN(ybar[93]);
  AND2_X1 U9 ( .A1(b[12]), .A2(a[5]), .ZN(y[92]) );
  OR2_X1 U9bar ( .A1(bbar[12]), .A2(abar[5]), .ZN(ybar[92]);
  AND2_X1 U10 ( .A1(b[11]), .A2(a[5]), .ZN(y[91]) );
  OR2_X1 U10bar ( .A1(bbar[11]), .A2(abar[5]), .ZN(ybar[91]);
  AND2_X1 U11 ( .A1(b[10]), .A2(a[5]), .ZN(y[90]) );
  OR2_X1 U11bar ( .A1(bbar[10]), .A2(abar[5]), .ZN(ybar[90]);
  AND2_X1 U12 ( .A1(b[8]), .A2(a[0]), .ZN(y[8]) );
  OR2_X1 U12bar ( .A1(bbar[8]), .A2(abar[0]), .ZN(ybar[8]);
  AND2_X1 U13 ( .A1(a[5]), .A2(b[9]), .ZN(y[89]) );
  OR2_X1 U13bar ( .A1(abar[5]), .A2(bbar[9]), .ZN(ybar[89]);
  AND2_X1 U14 ( .A1(b[8]), .A2(a[5]), .ZN(y[88]) );
  OR2_X1 U14bar ( .A1(bbar[8]), .A2(abar[5]), .ZN(ybar[88]);
  AND2_X1 U15 ( .A1(b[7]), .A2(a[5]), .ZN(y[87]) );
  OR2_X1 U15bar ( .A1(bbar[7]), .A2(abar[5]), .ZN(ybar[87]);
  AND2_X1 U16 ( .A1(b[6]), .A2(a[5]), .ZN(y[86]) );
  OR2_X1 U16bar ( .A1(bbar[6]), .A2(abar[5]), .ZN(ybar[86]);
  AND2_X1 U17 ( .A1(b[5]), .A2(a[5]), .ZN(y[85]) );
  OR2_X1 U17bar ( .A1(bbar[5]), .A2(abar[5]), .ZN(ybar[85]);
  AND2_X1 U18 ( .A1(b[4]), .A2(a[5]), .ZN(y[84]) );
  OR2_X1 U18bar ( .A1(bbar[4]), .A2(abar[5]), .ZN(ybar[84]);
  AND2_X1 U19 ( .A1(a[5]), .A2(b[3]), .ZN(y[83]) );
  OR2_X1 U19bar ( .A1(abar[5]), .A2(bbar[3]), .ZN(ybar[83]);
  AND2_X1 U20 ( .A1(a[5]), .A2(b[2]), .ZN(y[82]) );
  OR2_X1 U20bar ( .A1(abar[5]), .A2(bbar[2]), .ZN(ybar[82]);
  AND2_X1 U21 ( .A1(a[5]), .A2(b[1]), .ZN(y[81]) );
  OR2_X1 U21bar ( .A1(abar[5]), .A2(bbar[1]), .ZN(ybar[81]);
  AND2_X1 U22 ( .A1(a[5]), .A2(b[0]), .ZN(y[80]) );
  OR2_X1 U22bar ( .A1(abar[5]), .A2(bbar[0]), .ZN(ybar[80]);
  AND2_X1 U23 ( .A1(b[7]), .A2(a[0]), .ZN(y[7]) );
  OR2_X1 U23bar ( .A1(bbar[7]), .A2(abar[0]), .ZN(ybar[7]);
  AND2_X1 U24 ( .A1(a[4]), .A2(b[15]), .ZN(y[79]) );
  OR2_X1 U24bar ( .A1(abar[4]), .A2(bbar[15]), .ZN(ybar[79]);
  AND2_X1 U25 ( .A1(a[4]), .A2(b[14]), .ZN(y[78]) );
  OR2_X1 U25bar ( .A1(abar[4]), .A2(bbar[14]), .ZN(ybar[78]);
  AND2_X1 U26 ( .A1(a[4]), .A2(b[13]), .ZN(y[77]) );
  OR2_X1 U26bar ( .A1(abar[4]), .A2(bbar[13]), .ZN(ybar[77]);
  AND2_X1 U27 ( .A1(a[4]), .A2(b[12]), .ZN(y[76]) );
  OR2_X1 U27bar ( .A1(abar[4]), .A2(bbar[12]), .ZN(ybar[76]);
  AND2_X1 U28 ( .A1(a[4]), .A2(b[11]), .ZN(y[75]) );
  OR2_X1 U28bar ( .A1(abar[4]), .A2(bbar[11]), .ZN(ybar[75]);
  AND2_X1 U29 ( .A1(a[4]), .A2(b[10]), .ZN(y[74]) );
  OR2_X1 U29bar ( .A1(abar[4]), .A2(bbar[10]), .ZN(ybar[74]);
  AND2_X1 U30 ( .A1(a[4]), .A2(b[9]), .ZN(y[73]) );
  OR2_X1 U30bar ( .A1(abar[4]), .A2(bbar[9]), .ZN(ybar[73]);
  AND2_X1 U31 ( .A1(a[4]), .A2(b[8]), .ZN(y[72]) );
  OR2_X1 U31bar ( .A1(abar[4]), .A2(bbar[8]), .ZN(ybar[72]);
  AND2_X1 U32 ( .A1(a[4]), .A2(b[7]), .ZN(y[71]) );
  OR2_X1 U32bar ( .A1(abar[4]), .A2(bbar[7]), .ZN(ybar[71]);
  AND2_X1 U33 ( .A1(a[4]), .A2(b[6]), .ZN(y[70]) );
  OR2_X1 U33bar ( .A1(abar[4]), .A2(bbar[6]), .ZN(ybar[70]);
  AND2_X1 U34 ( .A1(b[6]), .A2(a[0]), .ZN(y[6]) );
  OR2_X1 U34bar ( .A1(bbar[6]), .A2(abar[0]), .ZN(ybar[6]);
  AND2_X1 U35 ( .A1(a[4]), .A2(b[5]), .ZN(y[69]) );
  OR2_X1 U35bar ( .A1(abar[4]), .A2(bbar[5]), .ZN(ybar[69]);
  AND2_X1 U36 ( .A1(a[4]), .A2(b[4]), .ZN(y[68]) );
  OR2_X1 U36bar ( .A1(abar[4]), .A2(bbar[4]), .ZN(ybar[68]);
  AND2_X1 U37 ( .A1(a[4]), .A2(b[3]), .ZN(y[67]) );
  OR2_X1 U37bar ( .A1(abar[4]), .A2(bbar[3]), .ZN(ybar[67]);
  AND2_X1 U38 ( .A1(a[4]), .A2(b[2]), .ZN(y[66]) );
  OR2_X1 U38bar ( .A1(abar[4]), .A2(bbar[2]), .ZN(ybar[66]);
  AND2_X1 U39 ( .A1(a[4]), .A2(b[1]), .ZN(y[65]) );
  OR2_X1 U39bar ( .A1(abar[4]), .A2(bbar[1]), .ZN(ybar[65]);
  AND2_X1 U40 ( .A1(a[4]), .A2(b[0]), .ZN(y[64]) );
  OR2_X1 U40bar ( .A1(abar[4]), .A2(bbar[0]), .ZN(ybar[64]);
  AND2_X1 U41 ( .A1(a[3]), .A2(b[15]), .ZN(y[63]) );
  OR2_X1 U41bar ( .A1(abar[3]), .A2(bbar[15]), .ZN(ybar[63]);
  AND2_X1 U42 ( .A1(a[3]), .A2(b[14]), .ZN(y[62]) );
  OR2_X1 U42bar ( .A1(abar[3]), .A2(bbar[14]), .ZN(ybar[62]);
  AND2_X1 U43 ( .A1(a[3]), .A2(b[13]), .ZN(y[61]) );
  OR2_X1 U43bar ( .A1(abar[3]), .A2(bbar[13]), .ZN(ybar[61]);
  AND2_X1 U44 ( .A1(a[3]), .A2(b[12]), .ZN(y[60]) );
  OR2_X1 U44bar ( .A1(abar[3]), .A2(bbar[12]), .ZN(ybar[60]);
  AND2_X1 U45 ( .A1(b[5]), .A2(a[0]), .ZN(y[5]) );
  OR2_X1 U45bar ( .A1(bbar[5]), .A2(abar[0]), .ZN(ybar[5]);
  AND2_X1 U46 ( .A1(a[3]), .A2(b[11]), .ZN(y[59]) );
  OR2_X1 U46bar ( .A1(abar[3]), .A2(bbar[11]), .ZN(ybar[59]);
  AND2_X1 U47 ( .A1(a[3]), .A2(b[10]), .ZN(y[58]) );
  OR2_X1 U47bar ( .A1(abar[3]), .A2(bbar[10]), .ZN(ybar[58]);
  AND2_X1 U48 ( .A1(a[3]), .A2(b[9]), .ZN(y[57]) );
  OR2_X1 U48bar ( .A1(abar[3]), .A2(bbar[9]), .ZN(ybar[57]);
  AND2_X1 U49 ( .A1(a[3]), .A2(b[8]), .ZN(y[56]) );
  OR2_X1 U49bar ( .A1(abar[3]), .A2(bbar[8]), .ZN(ybar[56]);
  AND2_X1 U50 ( .A1(a[3]), .A2(b[7]), .ZN(y[55]) );
  OR2_X1 U50bar ( .A1(abar[3]), .A2(bbar[7]), .ZN(ybar[55]);
  AND2_X1 U51 ( .A1(a[3]), .A2(b[6]), .ZN(y[54]) );
  OR2_X1 U51bar ( .A1(abar[3]), .A2(bbar[6]), .ZN(ybar[54]);
  AND2_X1 U52 ( .A1(a[3]), .A2(b[5]), .ZN(y[53]) );
  OR2_X1 U52bar ( .A1(abar[3]), .A2(bbar[5]), .ZN(ybar[53]);
  AND2_X1 U53 ( .A1(a[3]), .A2(b[4]), .ZN(y[52]) );
  OR2_X1 U53bar ( .A1(abar[3]), .A2(bbar[4]), .ZN(ybar[52]);
  AND2_X1 U54 ( .A1(a[3]), .A2(b[3]), .ZN(y[51]) );
  OR2_X1 U54bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[51]);
  AND2_X1 U55 ( .A1(a[3]), .A2(b[2]), .ZN(y[50]) );
  OR2_X1 U55bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[50]);
  AND2_X1 U56 ( .A1(b[4]), .A2(a[0]), .ZN(y[4]) );
  OR2_X1 U56bar ( .A1(bbar[4]), .A2(abar[0]), .ZN(ybar[4]);
  AND2_X1 U57 ( .A1(a[3]), .A2(b[1]), .ZN(y[49]) );
  OR2_X1 U57bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[49]);
  AND2_X1 U58 ( .A1(a[3]), .A2(b[0]), .ZN(y[48]) );
  OR2_X1 U58bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[48]);
  AND2_X1 U59 ( .A1(a[2]), .A2(b[15]), .ZN(y[47]) );
  OR2_X1 U59bar ( .A1(abar[2]), .A2(bbar[15]), .ZN(ybar[47]);
  AND2_X1 U60 ( .A1(a[2]), .A2(b[14]), .ZN(y[46]) );
  OR2_X1 U60bar ( .A1(abar[2]), .A2(bbar[14]), .ZN(ybar[46]);
  AND2_X1 U61 ( .A1(a[2]), .A2(b[13]), .ZN(y[45]) );
  OR2_X1 U61bar ( .A1(abar[2]), .A2(bbar[13]), .ZN(ybar[45]);
  AND2_X1 U62 ( .A1(a[2]), .A2(b[12]), .ZN(y[44]) );
  OR2_X1 U62bar ( .A1(abar[2]), .A2(bbar[12]), .ZN(ybar[44]);
  AND2_X1 U63 ( .A1(a[2]), .A2(b[11]), .ZN(y[43]) );
  OR2_X1 U63bar ( .A1(abar[2]), .A2(bbar[11]), .ZN(ybar[43]);
  AND2_X1 U64 ( .A1(a[2]), .A2(b[10]), .ZN(y[42]) );
  OR2_X1 U64bar ( .A1(abar[2]), .A2(bbar[10]), .ZN(ybar[42]);
  AND2_X1 U65 ( .A1(a[2]), .A2(b[9]), .ZN(y[41]) );
  OR2_X1 U65bar ( .A1(abar[2]), .A2(bbar[9]), .ZN(ybar[41]);
  AND2_X1 U66 ( .A1(a[2]), .A2(b[8]), .ZN(y[40]) );
  OR2_X1 U66bar ( .A1(abar[2]), .A2(bbar[8]), .ZN(ybar[40]);
  AND2_X1 U67 ( .A1(b[3]), .A2(a[0]), .ZN(y[3]) );
  OR2_X1 U67bar ( .A1(bbar[3]), .A2(abar[0]), .ZN(ybar[3]);
  AND2_X1 U68 ( .A1(a[2]), .A2(b[7]), .ZN(y[39]) );
  OR2_X1 U68bar ( .A1(abar[2]), .A2(bbar[7]), .ZN(ybar[39]);
  AND2_X1 U69 ( .A1(a[2]), .A2(b[6]), .ZN(y[38]) );
  OR2_X1 U69bar ( .A1(abar[2]), .A2(bbar[6]), .ZN(ybar[38]);
  AND2_X1 U70 ( .A1(a[2]), .A2(b[5]), .ZN(y[37]) );
  OR2_X1 U70bar ( .A1(abar[2]), .A2(bbar[5]), .ZN(ybar[37]);
  AND2_X1 U71 ( .A1(a[2]), .A2(b[4]), .ZN(y[36]) );
  OR2_X1 U71bar ( .A1(abar[2]), .A2(bbar[4]), .ZN(ybar[36]);
  AND2_X1 U72 ( .A1(a[2]), .A2(b[3]), .ZN(y[35]) );
  OR2_X1 U72bar ( .A1(abar[2]), .A2(bbar[3]), .ZN(ybar[35]);
  AND2_X1 U73 ( .A1(a[2]), .A2(b[2]), .ZN(y[34]) );
  OR2_X1 U73bar ( .A1(abar[2]), .A2(bbar[2]), .ZN(ybar[34]);
  AND2_X1 U74 ( .A1(a[2]), .A2(b[1]), .ZN(y[33]) );
  OR2_X1 U74bar ( .A1(abar[2]), .A2(bbar[1]), .ZN(ybar[33]);
  AND2_X1 U75 ( .A1(a[2]), .A2(b[0]), .ZN(y[32]) );
  OR2_X1 U75bar ( .A1(abar[2]), .A2(bbar[0]), .ZN(ybar[32]);
  AND2_X1 U76 ( .A1(a[1]), .A2(b[15]), .ZN(y[31]) );
  OR2_X1 U76bar ( .A1(abar[1]), .A2(bbar[15]), .ZN(ybar[31]);
  AND2_X1 U77 ( .A1(a[1]), .A2(b[14]), .ZN(y[30]) );
  OR2_X1 U77bar ( .A1(abar[1]), .A2(bbar[14]), .ZN(ybar[30]);
  AND2_X1 U78 ( .A1(b[2]), .A2(a[0]), .ZN(y[2]) );
  OR2_X1 U78bar ( .A1(bbar[2]), .A2(abar[0]), .ZN(ybar[2]);
  AND2_X1 U79 ( .A1(a[1]), .A2(b[13]), .ZN(y[29]) );
  OR2_X1 U79bar ( .A1(abar[1]), .A2(bbar[13]), .ZN(ybar[29]);
  AND2_X1 U80 ( .A1(a[1]), .A2(b[12]), .ZN(y[28]) );
  OR2_X1 U80bar ( .A1(abar[1]), .A2(bbar[12]), .ZN(ybar[28]);
  AND2_X1 U81 ( .A1(a[1]), .A2(b[11]), .ZN(y[27]) );
  OR2_X1 U81bar ( .A1(abar[1]), .A2(bbar[11]), .ZN(ybar[27]);
  AND2_X1 U82 ( .A1(a[1]), .A2(b[10]), .ZN(y[26]) );
  OR2_X1 U82bar ( .A1(abar[1]), .A2(bbar[10]), .ZN(ybar[26]);
  AND2_X1 U83 ( .A1(a[1]), .A2(b[9]), .ZN(y[25]) );
  OR2_X1 U83bar ( .A1(abar[1]), .A2(bbar[9]), .ZN(ybar[25]);
  AND2_X1 U84 ( .A1(a[15]), .A2(b[15]), .ZN(y[255]) );
  OR2_X1 U84bar ( .A1(abar[15]), .A2(bbar[15]), .ZN(ybar[255]);
  AND2_X1 U85 ( .A1(a[15]), .A2(b[14]), .ZN(y[254]) );
  OR2_X1 U85bar ( .A1(abar[15]), .A2(bbar[14]), .ZN(ybar[254]);
  AND2_X1 U86 ( .A1(a[15]), .A2(b[13]), .ZN(y[253]) );
  OR2_X1 U86bar ( .A1(abar[15]), .A2(bbar[13]), .ZN(ybar[253]);
  AND2_X1 U87 ( .A1(a[15]), .A2(b[12]), .ZN(y[252]) );
  OR2_X1 U87bar ( .A1(abar[15]), .A2(bbar[12]), .ZN(ybar[252]);
  AND2_X1 U88 ( .A1(a[15]), .A2(b[11]), .ZN(y[251]) );
  OR2_X1 U88bar ( .A1(abar[15]), .A2(bbar[11]), .ZN(ybar[251]);
  AND2_X1 U89 ( .A1(a[15]), .A2(b[10]), .ZN(y[250]) );
  OR2_X1 U89bar ( .A1(abar[15]), .A2(bbar[10]), .ZN(ybar[250]);
  AND2_X1 U90 ( .A1(a[1]), .A2(b[8]), .ZN(y[24]) );
  OR2_X1 U90bar ( .A1(abar[1]), .A2(bbar[8]), .ZN(ybar[24]);
  AND2_X1 U91 ( .A1(a[15]), .A2(b[9]), .ZN(y[249]) );
  OR2_X1 U91bar ( .A1(abar[15]), .A2(bbar[9]), .ZN(ybar[249]);
  AND2_X1 U92 ( .A1(a[15]), .A2(b[8]), .ZN(y[248]) );
  OR2_X1 U92bar ( .A1(abar[15]), .A2(bbar[8]), .ZN(ybar[248]);
  AND2_X1 U93 ( .A1(a[15]), .A2(b[7]), .ZN(y[247]) );
  OR2_X1 U93bar ( .A1(abar[15]), .A2(bbar[7]), .ZN(ybar[247]);
  AND2_X1 U94 ( .A1(a[15]), .A2(b[6]), .ZN(y[246]) );
  OR2_X1 U94bar ( .A1(abar[15]), .A2(bbar[6]), .ZN(ybar[246]);
  AND2_X1 U95 ( .A1(a[15]), .A2(b[5]), .ZN(y[245]) );
  OR2_X1 U95bar ( .A1(abar[15]), .A2(bbar[5]), .ZN(ybar[245]);
  AND2_X1 U96 ( .A1(a[15]), .A2(b[4]), .ZN(y[244]) );
  OR2_X1 U96bar ( .A1(abar[15]), .A2(bbar[4]), .ZN(ybar[244]);
  AND2_X1 U97 ( .A1(a[15]), .A2(b[3]), .ZN(y[243]) );
  OR2_X1 U97bar ( .A1(abar[15]), .A2(bbar[3]), .ZN(ybar[243]);
  AND2_X1 U98 ( .A1(a[15]), .A2(b[2]), .ZN(y[242]) );
  OR2_X1 U98bar ( .A1(abar[15]), .A2(bbar[2]), .ZN(ybar[242]);
  AND2_X1 U99 ( .A1(a[15]), .A2(b[1]), .ZN(y[241]) );
  OR2_X1 U99bar ( .A1(abar[15]), .A2(bbar[1]), .ZN(ybar[241]);
  AND2_X1 U100 ( .A1(a[15]), .A2(b[0]), .ZN(y[240]) );
  OR2_X1 U100bar ( .A1(abar[15]), .A2(bbar[0]), .ZN(ybar[240]);
  AND2_X1 U101 ( .A1(a[1]), .A2(b[7]), .ZN(y[23]) );
  OR2_X1 U101bar ( .A1(abar[1]), .A2(bbar[7]), .ZN(ybar[23]);
  AND2_X1 U102 ( .A1(a[14]), .A2(b[15]), .ZN(y[239]) );
  OR2_X1 U102bar ( .A1(abar[14]), .A2(bbar[15]), .ZN(ybar[239]);
  AND2_X1 U103 ( .A1(a[14]), .A2(b[14]), .ZN(y[238]) );
  OR2_X1 U103bar ( .A1(abar[14]), .A2(bbar[14]), .ZN(ybar[238]);
  AND2_X1 U104 ( .A1(a[14]), .A2(b[13]), .ZN(y[237]) );
  OR2_X1 U104bar ( .A1(abar[14]), .A2(bbar[13]), .ZN(ybar[237]);
  AND2_X1 U105 ( .A1(a[14]), .A2(b[12]), .ZN(y[236]) );
  OR2_X1 U105bar ( .A1(abar[14]), .A2(bbar[12]), .ZN(ybar[236]);
  AND2_X1 U106 ( .A1(a[14]), .A2(b[11]), .ZN(y[235]) );
  OR2_X1 U106bar ( .A1(abar[14]), .A2(bbar[11]), .ZN(ybar[235]);
  AND2_X1 U107 ( .A1(a[14]), .A2(b[10]), .ZN(y[234]) );
  OR2_X1 U107bar ( .A1(abar[14]), .A2(bbar[10]), .ZN(ybar[234]);
  AND2_X1 U108 ( .A1(a[14]), .A2(b[9]), .ZN(y[233]) );
  OR2_X1 U108bar ( .A1(abar[14]), .A2(bbar[9]), .ZN(ybar[233]);
  AND2_X1 U109 ( .A1(a[14]), .A2(b[8]), .ZN(y[232]) );
  OR2_X1 U109bar ( .A1(abar[14]), .A2(bbar[8]), .ZN(ybar[232]);
  AND2_X1 U110 ( .A1(a[14]), .A2(b[7]), .ZN(y[231]) );
  OR2_X1 U110bar ( .A1(abar[14]), .A2(bbar[7]), .ZN(ybar[231]);
  AND2_X1 U111 ( .A1(a[14]), .A2(b[6]), .ZN(y[230]) );
  OR2_X1 U111bar ( .A1(abar[14]), .A2(bbar[6]), .ZN(ybar[230]);
  AND2_X1 U112 ( .A1(a[1]), .A2(b[6]), .ZN(y[22]) );
  OR2_X1 U112bar ( .A1(abar[1]), .A2(bbar[6]), .ZN(ybar[22]);
  AND2_X1 U113 ( .A1(a[14]), .A2(b[5]), .ZN(y[229]) );
  OR2_X1 U113bar ( .A1(abar[14]), .A2(bbar[5]), .ZN(ybar[229]);
  AND2_X1 U114 ( .A1(a[14]), .A2(b[4]), .ZN(y[228]) );
  OR2_X1 U114bar ( .A1(abar[14]), .A2(bbar[4]), .ZN(ybar[228]);
  AND2_X1 U115 ( .A1(a[14]), .A2(b[3]), .ZN(y[227]) );
  OR2_X1 U115bar ( .A1(abar[14]), .A2(bbar[3]), .ZN(ybar[227]);
  AND2_X1 U116 ( .A1(a[14]), .A2(b[2]), .ZN(y[226]) );
  OR2_X1 U116bar ( .A1(abar[14]), .A2(bbar[2]), .ZN(ybar[226]);
  AND2_X1 U117 ( .A1(a[14]), .A2(b[1]), .ZN(y[225]) );
  OR2_X1 U117bar ( .A1(abar[14]), .A2(bbar[1]), .ZN(ybar[225]);
  AND2_X1 U118 ( .A1(a[14]), .A2(b[0]), .ZN(y[224]) );
  OR2_X1 U118bar ( .A1(abar[14]), .A2(bbar[0]), .ZN(ybar[224]);
  AND2_X1 U119 ( .A1(a[13]), .A2(b[15]), .ZN(y[223]) );
  OR2_X1 U119bar ( .A1(abar[13]), .A2(bbar[15]), .ZN(ybar[223]);
  AND2_X1 U120 ( .A1(a[13]), .A2(b[14]), .ZN(y[222]) );
  OR2_X1 U120bar ( .A1(abar[13]), .A2(bbar[14]), .ZN(ybar[222]);
  AND2_X1 U121 ( .A1(a[13]), .A2(b[13]), .ZN(y[221]) );
  OR2_X1 U121bar ( .A1(abar[13]), .A2(bbar[13]), .ZN(ybar[221]);
  AND2_X1 U122 ( .A1(a[13]), .A2(b[12]), .ZN(y[220]) );
  OR2_X1 U122bar ( .A1(abar[13]), .A2(bbar[12]), .ZN(ybar[220]);
  AND2_X1 U123 ( .A1(a[1]), .A2(b[5]), .ZN(y[21]) );
  OR2_X1 U123bar ( .A1(abar[1]), .A2(bbar[5]), .ZN(ybar[21]);
  AND2_X1 U124 ( .A1(a[13]), .A2(b[11]), .ZN(y[219]) );
  OR2_X1 U124bar ( .A1(abar[13]), .A2(bbar[11]), .ZN(ybar[219]);
  AND2_X1 U125 ( .A1(a[13]), .A2(b[10]), .ZN(y[218]) );
  OR2_X1 U125bar ( .A1(abar[13]), .A2(bbar[10]), .ZN(ybar[218]);
  AND2_X1 U126 ( .A1(a[13]), .A2(b[9]), .ZN(y[217]) );
  OR2_X1 U126bar ( .A1(abar[13]), .A2(bbar[9]), .ZN(ybar[217]);
  AND2_X1 U127 ( .A1(a[13]), .A2(b[8]), .ZN(y[216]) );
  OR2_X1 U127bar ( .A1(abar[13]), .A2(bbar[8]), .ZN(ybar[216]);
  AND2_X1 U128 ( .A1(a[13]), .A2(b[7]), .ZN(y[215]) );
  OR2_X1 U128bar ( .A1(abar[13]), .A2(bbar[7]), .ZN(ybar[215]);
  AND2_X1 U129 ( .A1(a[13]), .A2(b[6]), .ZN(y[214]) );
  OR2_X1 U129bar ( .A1(abar[13]), .A2(bbar[6]), .ZN(ybar[214]);
  AND2_X1 U130 ( .A1(a[13]), .A2(b[5]), .ZN(y[213]) );
  OR2_X1 U130bar ( .A1(abar[13]), .A2(bbar[5]), .ZN(ybar[213]);
  AND2_X1 U131 ( .A1(a[13]), .A2(b[4]), .ZN(y[212]) );
  OR2_X1 U131bar ( .A1(abar[13]), .A2(bbar[4]), .ZN(ybar[212]);
  AND2_X1 U132 ( .A1(a[13]), .A2(b[3]), .ZN(y[211]) );
  OR2_X1 U132bar ( .A1(abar[13]), .A2(bbar[3]), .ZN(ybar[211]);
  AND2_X1 U133 ( .A1(a[13]), .A2(b[2]), .ZN(y[210]) );
  OR2_X1 U133bar ( .A1(abar[13]), .A2(bbar[2]), .ZN(ybar[210]);
  AND2_X1 U134 ( .A1(a[1]), .A2(b[4]), .ZN(y[20]) );
  OR2_X1 U134bar ( .A1(abar[1]), .A2(bbar[4]), .ZN(ybar[20]);
  AND2_X1 U135 ( .A1(a[13]), .A2(b[1]), .ZN(y[209]) );
  OR2_X1 U135bar ( .A1(abar[13]), .A2(bbar[1]), .ZN(ybar[209]);
  AND2_X1 U136 ( .A1(a[13]), .A2(b[0]), .ZN(y[208]) );
  OR2_X1 U136bar ( .A1(abar[13]), .A2(bbar[0]), .ZN(ybar[208]);
  AND2_X1 U137 ( .A1(a[12]), .A2(b[15]), .ZN(y[207]) );
  OR2_X1 U137bar ( .A1(abar[12]), .A2(bbar[15]), .ZN(ybar[207]);
  AND2_X1 U138 ( .A1(a[12]), .A2(b[14]), .ZN(y[206]) );
  OR2_X1 U138bar ( .A1(abar[12]), .A2(bbar[14]), .ZN(ybar[206]);
  AND2_X1 U139 ( .A1(a[12]), .A2(b[13]), .ZN(y[205]) );
  OR2_X1 U139bar ( .A1(abar[12]), .A2(bbar[13]), .ZN(ybar[205]);
  AND2_X1 U140 ( .A1(a[12]), .A2(b[12]), .ZN(y[204]) );
  OR2_X1 U140bar ( .A1(abar[12]), .A2(bbar[12]), .ZN(ybar[204]);
  AND2_X1 U141 ( .A1(a[12]), .A2(b[11]), .ZN(y[203]) );
  OR2_X1 U141bar ( .A1(abar[12]), .A2(bbar[11]), .ZN(ybar[203]);
  AND2_X1 U142 ( .A1(a[12]), .A2(b[10]), .ZN(y[202]) );
  OR2_X1 U142bar ( .A1(abar[12]), .A2(bbar[10]), .ZN(ybar[202]);
  AND2_X1 U143 ( .A1(a[12]), .A2(b[9]), .ZN(y[201]) );
  OR2_X1 U143bar ( .A1(abar[12]), .A2(bbar[9]), .ZN(ybar[201]);
  AND2_X1 U144 ( .A1(a[12]), .A2(b[8]), .ZN(y[200]) );
  OR2_X1 U144bar ( .A1(abar[12]), .A2(bbar[8]), .ZN(ybar[200]);
  AND2_X1 U145 ( .A1(b[1]), .A2(a[0]), .ZN(y[1]) );
  OR2_X1 U145bar ( .A1(bbar[1]), .A2(abar[0]), .ZN(ybar[1]);
  AND2_X1 U146 ( .A1(a[1]), .A2(b[3]), .ZN(y[19]) );
  OR2_X1 U146bar ( .A1(abar[1]), .A2(bbar[3]), .ZN(ybar[19]);
  AND2_X1 U147 ( .A1(a[12]), .A2(b[7]), .ZN(y[199]) );
  OR2_X1 U147bar ( .A1(abar[12]), .A2(bbar[7]), .ZN(ybar[199]);
  AND2_X1 U148 ( .A1(a[12]), .A2(b[6]), .ZN(y[198]) );
  OR2_X1 U148bar ( .A1(abar[12]), .A2(bbar[6]), .ZN(ybar[198]);
  AND2_X1 U149 ( .A1(a[12]), .A2(b[5]), .ZN(y[197]) );
  OR2_X1 U149bar ( .A1(abar[12]), .A2(bbar[5]), .ZN(ybar[197]);
  AND2_X1 U150 ( .A1(a[12]), .A2(b[4]), .ZN(y[196]) );
  OR2_X1 U150bar ( .A1(abar[12]), .A2(bbar[4]), .ZN(ybar[196]);
  AND2_X1 U151 ( .A1(a[12]), .A2(b[3]), .ZN(y[195]) );
  OR2_X1 U151bar ( .A1(abar[12]), .A2(bbar[3]), .ZN(ybar[195]);
  AND2_X1 U152 ( .A1(a[12]), .A2(b[2]), .ZN(y[194]) );
  OR2_X1 U152bar ( .A1(abar[12]), .A2(bbar[2]), .ZN(ybar[194]);
  AND2_X1 U153 ( .A1(a[12]), .A2(b[1]), .ZN(y[193]) );
  OR2_X1 U153bar ( .A1(abar[12]), .A2(bbar[1]), .ZN(ybar[193]);
  AND2_X1 U154 ( .A1(a[12]), .A2(b[0]), .ZN(y[192]) );
  OR2_X1 U154bar ( .A1(abar[12]), .A2(bbar[0]), .ZN(ybar[192]);
  AND2_X1 U155 ( .A1(a[11]), .A2(b[15]), .ZN(y[191]) );
  OR2_X1 U155bar ( .A1(abar[11]), .A2(bbar[15]), .ZN(ybar[191]);
  AND2_X1 U156 ( .A1(a[11]), .A2(b[14]), .ZN(y[190]) );
  OR2_X1 U156bar ( .A1(abar[11]), .A2(bbar[14]), .ZN(ybar[190]);
  AND2_X1 U157 ( .A1(a[1]), .A2(b[2]), .ZN(y[18]) );
  OR2_X1 U157bar ( .A1(abar[1]), .A2(bbar[2]), .ZN(ybar[18]);
  AND2_X1 U158 ( .A1(a[11]), .A2(b[13]), .ZN(y[189]) );
  OR2_X1 U158bar ( .A1(abar[11]), .A2(bbar[13]), .ZN(ybar[189]);
  AND2_X1 U159 ( .A1(a[11]), .A2(b[12]), .ZN(y[188]) );
  OR2_X1 U159bar ( .A1(abar[11]), .A2(bbar[12]), .ZN(ybar[188]);
  AND2_X1 U160 ( .A1(a[11]), .A2(b[11]), .ZN(y[187]) );
  OR2_X1 U160bar ( .A1(abar[11]), .A2(bbar[11]), .ZN(ybar[187]);
  AND2_X1 U161 ( .A1(a[11]), .A2(b[10]), .ZN(y[186]) );
  OR2_X1 U161bar ( .A1(abar[11]), .A2(bbar[10]), .ZN(ybar[186]);
  AND2_X1 U162 ( .A1(a[11]), .A2(b[9]), .ZN(y[185]) );
  OR2_X1 U162bar ( .A1(abar[11]), .A2(bbar[9]), .ZN(ybar[185]);
  AND2_X1 U163 ( .A1(a[11]), .A2(b[8]), .ZN(y[184]) );
  OR2_X1 U163bar ( .A1(abar[11]), .A2(bbar[8]), .ZN(ybar[184]);
  AND2_X1 U164 ( .A1(a[11]), .A2(b[7]), .ZN(y[183]) );
  OR2_X1 U164bar ( .A1(abar[11]), .A2(bbar[7]), .ZN(ybar[183]);
  AND2_X1 U165 ( .A1(a[11]), .A2(b[6]), .ZN(y[182]) );
  OR2_X1 U165bar ( .A1(abar[11]), .A2(bbar[6]), .ZN(ybar[182]);
  AND2_X1 U166 ( .A1(a[11]), .A2(b[5]), .ZN(y[181]) );
  OR2_X1 U166bar ( .A1(abar[11]), .A2(bbar[5]), .ZN(ybar[181]);
  AND2_X1 U167 ( .A1(a[11]), .A2(b[4]), .ZN(y[180]) );
  OR2_X1 U167bar ( .A1(abar[11]), .A2(bbar[4]), .ZN(ybar[180]);
  AND2_X1 U168 ( .A1(a[1]), .A2(b[1]), .ZN(y[17]) );
  OR2_X1 U168bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[17]);
  AND2_X1 U169 ( .A1(a[11]), .A2(b[3]), .ZN(y[179]) );
  OR2_X1 U169bar ( .A1(abar[11]), .A2(bbar[3]), .ZN(ybar[179]);
  AND2_X1 U170 ( .A1(a[11]), .A2(b[2]), .ZN(y[178]) );
  OR2_X1 U170bar ( .A1(abar[11]), .A2(bbar[2]), .ZN(ybar[178]);
  AND2_X1 U171 ( .A1(a[11]), .A2(b[1]), .ZN(y[177]) );
  OR2_X1 U171bar ( .A1(abar[11]), .A2(bbar[1]), .ZN(ybar[177]);
  AND2_X1 U172 ( .A1(a[11]), .A2(b[0]), .ZN(y[176]) );
  OR2_X1 U172bar ( .A1(abar[11]), .A2(bbar[0]), .ZN(ybar[176]);
  AND2_X1 U173 ( .A1(a[10]), .A2(b[15]), .ZN(y[175]) );
  OR2_X1 U173bar ( .A1(abar[10]), .A2(bbar[15]), .ZN(ybar[175]);
  AND2_X1 U174 ( .A1(a[10]), .A2(b[14]), .ZN(y[174]) );
  OR2_X1 U174bar ( .A1(abar[10]), .A2(bbar[14]), .ZN(ybar[174]);
  AND2_X1 U175 ( .A1(a[10]), .A2(b[13]), .ZN(y[173]) );
  OR2_X1 U175bar ( .A1(abar[10]), .A2(bbar[13]), .ZN(ybar[173]);
  AND2_X1 U176 ( .A1(a[10]), .A2(b[12]), .ZN(y[172]) );
  OR2_X1 U176bar ( .A1(abar[10]), .A2(bbar[12]), .ZN(ybar[172]);
  AND2_X1 U177 ( .A1(a[10]), .A2(b[11]), .ZN(y[171]) );
  OR2_X1 U177bar ( .A1(abar[10]), .A2(bbar[11]), .ZN(ybar[171]);
  AND2_X1 U178 ( .A1(a[10]), .A2(b[10]), .ZN(y[170]) );
  OR2_X1 U178bar ( .A1(abar[10]), .A2(bbar[10]), .ZN(ybar[170]);
  AND2_X1 U179 ( .A1(a[1]), .A2(b[0]), .ZN(y[16]) );
  OR2_X1 U179bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[16]);
  AND2_X1 U180 ( .A1(a[10]), .A2(b[9]), .ZN(y[169]) );
  OR2_X1 U180bar ( .A1(abar[10]), .A2(bbar[9]), .ZN(ybar[169]);
  AND2_X1 U181 ( .A1(a[10]), .A2(b[8]), .ZN(y[168]) );
  OR2_X1 U181bar ( .A1(abar[10]), .A2(bbar[8]), .ZN(ybar[168]);
  AND2_X1 U182 ( .A1(a[10]), .A2(b[7]), .ZN(y[167]) );
  OR2_X1 U182bar ( .A1(abar[10]), .A2(bbar[7]), .ZN(ybar[167]);
  AND2_X1 U183 ( .A1(a[10]), .A2(b[6]), .ZN(y[166]) );
  OR2_X1 U183bar ( .A1(abar[10]), .A2(bbar[6]), .ZN(ybar[166]);
  AND2_X1 U184 ( .A1(a[10]), .A2(b[5]), .ZN(y[165]) );
  OR2_X1 U184bar ( .A1(abar[10]), .A2(bbar[5]), .ZN(ybar[165]);
  AND2_X1 U185 ( .A1(a[10]), .A2(b[4]), .ZN(y[164]) );
  OR2_X1 U185bar ( .A1(abar[10]), .A2(bbar[4]), .ZN(ybar[164]);
  AND2_X1 U186 ( .A1(a[10]), .A2(b[3]), .ZN(y[163]) );
  OR2_X1 U186bar ( .A1(abar[10]), .A2(bbar[3]), .ZN(ybar[163]);
  AND2_X1 U187 ( .A1(a[10]), .A2(b[2]), .ZN(y[162]) );
  OR2_X1 U187bar ( .A1(abar[10]), .A2(bbar[2]), .ZN(ybar[162]);
  AND2_X1 U188 ( .A1(a[10]), .A2(b[1]), .ZN(y[161]) );
  OR2_X1 U188bar ( .A1(abar[10]), .A2(bbar[1]), .ZN(ybar[161]);
  AND2_X1 U189 ( .A1(a[10]), .A2(b[0]), .ZN(y[160]) );
  OR2_X1 U189bar ( .A1(abar[10]), .A2(bbar[0]), .ZN(ybar[160]);
  AND2_X1 U190 ( .A1(b[15]), .A2(a[0]), .ZN(y[15]) );
  OR2_X1 U190bar ( .A1(bbar[15]), .A2(abar[0]), .ZN(ybar[15]);
  AND2_X1 U191 ( .A1(a[9]), .A2(b[15]), .ZN(y[159]) );
  OR2_X1 U191bar ( .A1(abar[9]), .A2(bbar[15]), .ZN(ybar[159]);
  AND2_X1 U192 ( .A1(a[9]), .A2(b[14]), .ZN(y[158]) );
  OR2_X1 U192bar ( .A1(abar[9]), .A2(bbar[14]), .ZN(ybar[158]);
  AND2_X1 U193 ( .A1(a[9]), .A2(b[13]), .ZN(y[157]) );
  OR2_X1 U193bar ( .A1(abar[9]), .A2(bbar[13]), .ZN(ybar[157]);
  AND2_X1 U194 ( .A1(a[9]), .A2(b[12]), .ZN(y[156]) );
  OR2_X1 U194bar ( .A1(abar[9]), .A2(bbar[12]), .ZN(ybar[156]);
  AND2_X1 U195 ( .A1(a[9]), .A2(b[11]), .ZN(y[155]) );
  OR2_X1 U195bar ( .A1(abar[9]), .A2(bbar[11]), .ZN(ybar[155]);
  AND2_X1 U196 ( .A1(a[9]), .A2(b[10]), .ZN(y[154]) );
  OR2_X1 U196bar ( .A1(abar[9]), .A2(bbar[10]), .ZN(ybar[154]);
  AND2_X1 U197 ( .A1(a[9]), .A2(b[9]), .ZN(y[153]) );
  OR2_X1 U197bar ( .A1(abar[9]), .A2(bbar[9]), .ZN(ybar[153]);
  AND2_X1 U198 ( .A1(a[9]), .A2(b[8]), .ZN(y[152]) );
  OR2_X1 U198bar ( .A1(abar[9]), .A2(bbar[8]), .ZN(ybar[152]);
  AND2_X1 U199 ( .A1(a[9]), .A2(b[7]), .ZN(y[151]) );
  OR2_X1 U199bar ( .A1(abar[9]), .A2(bbar[7]), .ZN(ybar[151]);
  AND2_X1 U200 ( .A1(a[9]), .A2(b[6]), .ZN(y[150]) );
  OR2_X1 U200bar ( .A1(abar[9]), .A2(bbar[6]), .ZN(ybar[150]);
  AND2_X1 U201 ( .A1(b[14]), .A2(a[0]), .ZN(y[14]) );
  OR2_X1 U201bar ( .A1(bbar[14]), .A2(abar[0]), .ZN(ybar[14]);
  AND2_X1 U202 ( .A1(a[9]), .A2(b[5]), .ZN(y[149]) );
  OR2_X1 U202bar ( .A1(abar[9]), .A2(bbar[5]), .ZN(ybar[149]);
  AND2_X1 U203 ( .A1(a[9]), .A2(b[4]), .ZN(y[148]) );
  OR2_X1 U203bar ( .A1(abar[9]), .A2(bbar[4]), .ZN(ybar[148]);
  AND2_X1 U204 ( .A1(a[9]), .A2(b[3]), .ZN(y[147]) );
  OR2_X1 U204bar ( .A1(abar[9]), .A2(bbar[3]), .ZN(ybar[147]);
  AND2_X1 U205 ( .A1(a[9]), .A2(b[2]), .ZN(y[146]) );
  OR2_X1 U205bar ( .A1(abar[9]), .A2(bbar[2]), .ZN(ybar[146]);
  AND2_X1 U206 ( .A1(a[9]), .A2(b[1]), .ZN(y[145]) );
  OR2_X1 U206bar ( .A1(abar[9]), .A2(bbar[1]), .ZN(ybar[145]);
  AND2_X1 U207 ( .A1(a[9]), .A2(b[0]), .ZN(y[144]) );
  OR2_X1 U207bar ( .A1(abar[9]), .A2(bbar[0]), .ZN(ybar[144]);
  AND2_X1 U208 ( .A1(a[8]), .A2(b[15]), .ZN(y[143]) );
  OR2_X1 U208bar ( .A1(abar[8]), .A2(bbar[15]), .ZN(ybar[143]);
  AND2_X1 U209 ( .A1(a[8]), .A2(b[14]), .ZN(y[142]) );
  OR2_X1 U209bar ( .A1(abar[8]), .A2(bbar[14]), .ZN(ybar[142]);
  AND2_X1 U210 ( .A1(a[8]), .A2(b[13]), .ZN(y[141]) );
  OR2_X1 U210bar ( .A1(abar[8]), .A2(bbar[13]), .ZN(ybar[141]);
  AND2_X1 U211 ( .A1(a[8]), .A2(b[12]), .ZN(y[140]) );
  OR2_X1 U211bar ( .A1(abar[8]), .A2(bbar[12]), .ZN(ybar[140]);
  AND2_X1 U212 ( .A1(b[13]), .A2(a[0]), .ZN(y[13]) );
  OR2_X1 U212bar ( .A1(bbar[13]), .A2(abar[0]), .ZN(ybar[13]);
  AND2_X1 U213 ( .A1(a[8]), .A2(b[11]), .ZN(y[139]) );
  OR2_X1 U213bar ( .A1(abar[8]), .A2(bbar[11]), .ZN(ybar[139]);
  AND2_X1 U214 ( .A1(a[8]), .A2(b[10]), .ZN(y[138]) );
  OR2_X1 U214bar ( .A1(abar[8]), .A2(bbar[10]), .ZN(ybar[138]);
  AND2_X1 U215 ( .A1(a[8]), .A2(b[9]), .ZN(y[137]) );
  OR2_X1 U215bar ( .A1(abar[8]), .A2(bbar[9]), .ZN(ybar[137]);
  AND2_X1 U216 ( .A1(a[8]), .A2(b[8]), .ZN(y[136]) );
  OR2_X1 U216bar ( .A1(abar[8]), .A2(bbar[8]), .ZN(ybar[136]);
  AND2_X1 U217 ( .A1(a[8]), .A2(b[7]), .ZN(y[135]) );
  OR2_X1 U217bar ( .A1(abar[8]), .A2(bbar[7]), .ZN(ybar[135]);
  AND2_X1 U218 ( .A1(a[8]), .A2(b[6]), .ZN(y[134]) );
  OR2_X1 U218bar ( .A1(abar[8]), .A2(bbar[6]), .ZN(ybar[134]);
  AND2_X1 U219 ( .A1(a[8]), .A2(b[5]), .ZN(y[133]) );
  OR2_X1 U219bar ( .A1(abar[8]), .A2(bbar[5]), .ZN(ybar[133]);
  AND2_X1 U220 ( .A1(a[8]), .A2(b[4]), .ZN(y[132]) );
  OR2_X1 U220bar ( .A1(abar[8]), .A2(bbar[4]), .ZN(ybar[132]);
  AND2_X1 U221 ( .A1(a[8]), .A2(b[3]), .ZN(y[131]) );
  OR2_X1 U221bar ( .A1(abar[8]), .A2(bbar[3]), .ZN(ybar[131]);
  AND2_X1 U222 ( .A1(a[8]), .A2(b[2]), .ZN(y[130]) );
  OR2_X1 U222bar ( .A1(abar[8]), .A2(bbar[2]), .ZN(ybar[130]);
  AND2_X1 U223 ( .A1(b[12]), .A2(a[0]), .ZN(y[12]) );
  OR2_X1 U223bar ( .A1(bbar[12]), .A2(abar[0]), .ZN(ybar[12]);
  AND2_X1 U224 ( .A1(a[8]), .A2(b[1]), .ZN(y[129]) );
  OR2_X1 U224bar ( .A1(abar[8]), .A2(bbar[1]), .ZN(ybar[129]);
  AND2_X1 U225 ( .A1(a[8]), .A2(b[0]), .ZN(y[128]) );
  OR2_X1 U225bar ( .A1(abar[8]), .A2(bbar[0]), .ZN(ybar[128]);
  AND2_X1 U226 ( .A1(a[7]), .A2(b[15]), .ZN(y[127]) );
  OR2_X1 U226bar ( .A1(abar[7]), .A2(bbar[15]), .ZN(ybar[127]);
  AND2_X1 U227 ( .A1(a[7]), .A2(b[14]), .ZN(y[126]) );
  OR2_X1 U227bar ( .A1(abar[7]), .A2(bbar[14]), .ZN(ybar[126]);
  AND2_X1 U228 ( .A1(a[7]), .A2(b[13]), .ZN(y[125]) );
  OR2_X1 U228bar ( .A1(abar[7]), .A2(bbar[13]), .ZN(ybar[125]);
  AND2_X1 U229 ( .A1(a[7]), .A2(b[12]), .ZN(y[124]) );
  OR2_X1 U229bar ( .A1(abar[7]), .A2(bbar[12]), .ZN(ybar[124]);
  AND2_X1 U230 ( .A1(a[7]), .A2(b[11]), .ZN(y[123]) );
  OR2_X1 U230bar ( .A1(abar[7]), .A2(bbar[11]), .ZN(ybar[123]);
  AND2_X1 U231 ( .A1(a[7]), .A2(b[10]), .ZN(y[122]) );
  OR2_X1 U231bar ( .A1(abar[7]), .A2(bbar[10]), .ZN(ybar[122]);
  AND2_X1 U232 ( .A1(a[7]), .A2(b[9]), .ZN(y[121]) );
  OR2_X1 U232bar ( .A1(abar[7]), .A2(bbar[9]), .ZN(ybar[121]);
  AND2_X1 U233 ( .A1(a[7]), .A2(b[8]), .ZN(y[120]) );
  OR2_X1 U233bar ( .A1(abar[7]), .A2(bbar[8]), .ZN(ybar[120]);
  AND2_X1 U234 ( .A1(b[11]), .A2(a[0]), .ZN(y[11]) );
  OR2_X1 U234bar ( .A1(bbar[11]), .A2(abar[0]), .ZN(ybar[11]);
  AND2_X1 U235 ( .A1(a[7]), .A2(b[7]), .ZN(y[119]) );
  OR2_X1 U235bar ( .A1(abar[7]), .A2(bbar[7]), .ZN(ybar[119]);
  AND2_X1 U236 ( .A1(a[7]), .A2(b[6]), .ZN(y[118]) );
  OR2_X1 U236bar ( .A1(abar[7]), .A2(bbar[6]), .ZN(ybar[118]);
  AND2_X1 U237 ( .A1(a[7]), .A2(b[5]), .ZN(y[117]) );
  OR2_X1 U237bar ( .A1(abar[7]), .A2(bbar[5]), .ZN(ybar[117]);
  AND2_X1 U238 ( .A1(a[7]), .A2(b[4]), .ZN(y[116]) );
  OR2_X1 U238bar ( .A1(abar[7]), .A2(bbar[4]), .ZN(ybar[116]);
  AND2_X1 U239 ( .A1(a[7]), .A2(b[3]), .ZN(y[115]) );
  OR2_X1 U239bar ( .A1(abar[7]), .A2(bbar[3]), .ZN(ybar[115]);
  AND2_X1 U240 ( .A1(a[7]), .A2(b[2]), .ZN(y[114]) );
  OR2_X1 U240bar ( .A1(abar[7]), .A2(bbar[2]), .ZN(ybar[114]);
  AND2_X1 U241 ( .A1(a[7]), .A2(b[1]), .ZN(y[113]) );
  OR2_X1 U241bar ( .A1(abar[7]), .A2(bbar[1]), .ZN(ybar[113]);
  AND2_X1 U242 ( .A1(a[7]), .A2(b[0]), .ZN(y[112]) );
  OR2_X1 U242bar ( .A1(abar[7]), .A2(bbar[0]), .ZN(ybar[112]);
  AND2_X1 U243 ( .A1(b[15]), .A2(a[6]), .ZN(y[111]) );
  OR2_X1 U243bar ( .A1(bbar[15]), .A2(abar[6]), .ZN(ybar[111]);
  AND2_X1 U244 ( .A1(b[14]), .A2(a[6]), .ZN(y[110]) );
  OR2_X1 U244bar ( .A1(bbar[14]), .A2(abar[6]), .ZN(ybar[110]);
  AND2_X1 U245 ( .A1(b[10]), .A2(a[0]), .ZN(y[10]) );
  OR2_X1 U245bar ( .A1(bbar[10]), .A2(abar[0]), .ZN(ybar[10]);
  AND2_X1 U246 ( .A1(b[13]), .A2(a[6]), .ZN(y[109]) );
  OR2_X1 U246bar ( .A1(bbar[13]), .A2(abar[6]), .ZN(ybar[109]);
  AND2_X1 U247 ( .A1(b[12]), .A2(a[6]), .ZN(y[108]) );
  OR2_X1 U247bar ( .A1(bbar[12]), .A2(abar[6]), .ZN(ybar[108]);
  AND2_X1 U248 ( .A1(b[11]), .A2(a[6]), .ZN(y[107]) );
  OR2_X1 U248bar ( .A1(bbar[11]), .A2(abar[6]), .ZN(ybar[107]);
  AND2_X1 U249 ( .A1(b[10]), .A2(a[6]), .ZN(y[106]) );
  OR2_X1 U249bar ( .A1(bbar[10]), .A2(abar[6]), .ZN(ybar[106]);
  AND2_X1 U250 ( .A1(a[6]), .A2(b[9]), .ZN(y[105]) );
  OR2_X1 U250bar ( .A1(abar[6]), .A2(bbar[9]), .ZN(ybar[105]);
  AND2_X1 U251 ( .A1(b[8]), .A2(a[6]), .ZN(y[104]) );
  OR2_X1 U251bar ( .A1(bbar[8]), .A2(abar[6]), .ZN(ybar[104]);
  AND2_X1 U252 ( .A1(b[7]), .A2(a[6]), .ZN(y[103]) );
  OR2_X1 U252bar ( .A1(bbar[7]), .A2(abar[6]), .ZN(ybar[103]);
  AND2_X1 U253 ( .A1(b[6]), .A2(a[6]), .ZN(y[102]) );
  OR2_X1 U253bar ( .A1(bbar[6]), .A2(abar[6]), .ZN(ybar[102]);
  AND2_X1 U254 ( .A1(b[5]), .A2(a[6]), .ZN(y[101]) );
  OR2_X1 U254bar ( .A1(bbar[5]), .A2(abar[6]), .ZN(ybar[101]);
  AND2_X1 U255 ( .A1(b[4]), .A2(a[6]), .ZN(y[100]) );
  OR2_X1 U255bar ( .A1(bbar[4]), .A2(abar[6]), .ZN(ybar[100]);
  AND2_X1 U256 ( .A1(b[0]), .A2(a[0]), .ZN(y[0]) );
  OR2_X1 U256bar ( .A1(bbar[0]), .A2(abar[0]), .ZN(ybar[0]);
endmodule




module decode_17 ( in, out );
  input [7:0] in;
  //input_done

  output [255:0] out;
  //output_done

  wire   [15:0] level1;
  wire   [31:0] level2;
  //wire_done

  CD2_68 cd_l1_1 ( .a(in[1]), .b(in[0]), .y(level1[3:0]) );
  CD2_67 cd_l1_2 ( .a(in[3]), .b(in[2]), .y(level1[7:4]) );
  CD2_66 cd_l1_3 ( .a(in[5]), .b(in[4]), .y(level1[11:8]) );
  CD2_65 cd_l1_4 ( .a(in[7]), .b(in[6]), .y(level1[15:12]) );
  CD4_34 cd_l2_1 ( .a(level1[7:4]), .b(level1[3:0]), .y(level2[15:0]) );
  CD4_33 cd_l2_2 ( .a(level1[15:12]), .b(level1[11:8]), .y(level2[31:16]) );
  CD16_17 cd_l3 ( .a(level2[31:16]), .b(level2[15:0]), .y(out) );
endmodule


module encode_17 ( in, out );
  input [255:0] in;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
  assign inbar[8] = ~in[8];
  assign inbar[9] = ~in[9];
  assign inbar[10] = ~in[10];
  assign inbar[11] = ~in[11];
  assign inbar[12] = ~in[12];
  assign inbar[13] = ~in[13];
  assign inbar[14] = ~in[14];
  assign inbar[15] = ~in[15];
  assign inbar[16] = ~in[16];
  assign inbar[17] = ~in[17];
  assign inbar[18] = ~in[18];
  assign inbar[19] = ~in[19];
  assign inbar[20] = ~in[20];
  assign inbar[21] = ~in[21];
  assign inbar[22] = ~in[22];
  assign inbar[23] = ~in[23];
  assign inbar[24] = ~in[24];
  assign inbar[25] = ~in[25];
  assign inbar[26] = ~in[26];
  assign inbar[27] = ~in[27];
  assign inbar[28] = ~in[28];
  assign inbar[29] = ~in[29];
  assign inbar[30] = ~in[30];
  assign inbar[31] = ~in[31];
  assign inbar[32] = ~in[32];
  assign inbar[33] = ~in[33];
  assign inbar[34] = ~in[34];
  assign inbar[35] = ~in[35];
  assign inbar[36] = ~in[36];
  assign inbar[37] = ~in[37];
  assign inbar[38] = ~in[38];
  assign inbar[39] = ~in[39];
  assign inbar[40] = ~in[40];
  assign inbar[41] = ~in[41];
  assign inbar[42] = ~in[42];
  assign inbar[43] = ~in[43];
  assign inbar[44] = ~in[44];
  assign inbar[45] = ~in[45];
  assign inbar[46] = ~in[46];
  assign inbar[47] = ~in[47];
  assign inbar[48] = ~in[48];
  assign inbar[49] = ~in[49];
  assign inbar[50] = ~in[50];
  assign inbar[51] = ~in[51];
  assign inbar[52] = ~in[52];
  assign inbar[53] = ~in[53];
  assign inbar[54] = ~in[54];
  assign inbar[55] = ~in[55];
  assign inbar[56] = ~in[56];
  assign inbar[57] = ~in[57];
  assign inbar[58] = ~in[58];
  assign inbar[59] = ~in[59];
  assign inbar[60] = ~in[60];
  assign inbar[61] = ~in[61];
  assign inbar[62] = ~in[62];
  assign inbar[63] = ~in[63];
  assign inbar[64] = ~in[64];
  assign inbar[65] = ~in[65];
  assign inbar[66] = ~in[66];
  assign inbar[67] = ~in[67];
  assign inbar[68] = ~in[68];
  assign inbar[69] = ~in[69];
  assign inbar[70] = ~in[70];
  assign inbar[71] = ~in[71];
  assign inbar[72] = ~in[72];
  assign inbar[73] = ~in[73];
  assign inbar[74] = ~in[74];
  assign inbar[75] = ~in[75];
  assign inbar[76] = ~in[76];
  assign inbar[77] = ~in[77];
  assign inbar[78] = ~in[78];
  assign inbar[79] = ~in[79];
  assign inbar[80] = ~in[80];
  assign inbar[81] = ~in[81];
  assign inbar[82] = ~in[82];
  assign inbar[83] = ~in[83];
  assign inbar[84] = ~in[84];
  assign inbar[85] = ~in[85];
  assign inbar[86] = ~in[86];
  assign inbar[87] = ~in[87];
  assign inbar[88] = ~in[88];
  assign inbar[89] = ~in[89];
  assign inbar[90] = ~in[90];
  assign inbar[91] = ~in[91];
  assign inbar[92] = ~in[92];
  assign inbar[93] = ~in[93];
  assign inbar[94] = ~in[94];
  assign inbar[95] = ~in[95];
  assign inbar[96] = ~in[96];
  assign inbar[97] = ~in[97];
  assign inbar[98] = ~in[98];
  assign inbar[99] = ~in[99];
  assign inbar[100] = ~in[100];
  assign inbar[101] = ~in[101];
  assign inbar[102] = ~in[102];
  assign inbar[103] = ~in[103];
  assign inbar[104] = ~in[104];
  assign inbar[105] = ~in[105];
  assign inbar[106] = ~in[106];
  assign inbar[107] = ~in[107];
  assign inbar[108] = ~in[108];
  assign inbar[109] = ~in[109];
  assign inbar[110] = ~in[110];
  assign inbar[111] = ~in[111];
  assign inbar[112] = ~in[112];
  assign inbar[113] = ~in[113];
  assign inbar[114] = ~in[114];
  assign inbar[115] = ~in[115];
  assign inbar[116] = ~in[116];
  assign inbar[117] = ~in[117];
  assign inbar[118] = ~in[118];
  assign inbar[119] = ~in[119];
  assign inbar[120] = ~in[120];
  assign inbar[121] = ~in[121];
  assign inbar[122] = ~in[122];
  assign inbar[123] = ~in[123];
  assign inbar[124] = ~in[124];
  assign inbar[125] = ~in[125];
  assign inbar[126] = ~in[126];
  assign inbar[127] = ~in[127];
  assign inbar[128] = ~in[128];
  assign inbar[129] = ~in[129];
  assign inbar[130] = ~in[130];
  assign inbar[131] = ~in[131];
  assign inbar[132] = ~in[132];
  assign inbar[133] = ~in[133];
  assign inbar[134] = ~in[134];
  assign inbar[135] = ~in[135];
  assign inbar[136] = ~in[136];
  assign inbar[137] = ~in[137];
  assign inbar[138] = ~in[138];
  assign inbar[139] = ~in[139];
  assign inbar[140] = ~in[140];
  assign inbar[141] = ~in[141];
  assign inbar[142] = ~in[142];
  assign inbar[143] = ~in[143];
  assign inbar[144] = ~in[144];
  assign inbar[145] = ~in[145];
  assign inbar[146] = ~in[146];
  assign inbar[147] = ~in[147];
  assign inbar[148] = ~in[148];
  assign inbar[149] = ~in[149];
  assign inbar[150] = ~in[150];
  assign inbar[151] = ~in[151];
  assign inbar[152] = ~in[152];
  assign inbar[153] = ~in[153];
  assign inbar[154] = ~in[154];
  assign inbar[155] = ~in[155];
  assign inbar[156] = ~in[156];
  assign inbar[157] = ~in[157];
  assign inbar[158] = ~in[158];
  assign inbar[159] = ~in[159];
  assign inbar[160] = ~in[160];
  assign inbar[161] = ~in[161];
  assign inbar[162] = ~in[162];
  assign inbar[163] = ~in[163];
  assign inbar[164] = ~in[164];
  assign inbar[165] = ~in[165];
  assign inbar[166] = ~in[166];
  assign inbar[167] = ~in[167];
  assign inbar[168] = ~in[168];
  assign inbar[169] = ~in[169];
  assign inbar[170] = ~in[170];
  assign inbar[171] = ~in[171];
  assign inbar[172] = ~in[172];
  assign inbar[173] = ~in[173];
  assign inbar[174] = ~in[174];
  assign inbar[175] = ~in[175];
  assign inbar[176] = ~in[176];
  assign inbar[177] = ~in[177];
  assign inbar[178] = ~in[178];
  assign inbar[179] = ~in[179];
  assign inbar[180] = ~in[180];
  assign inbar[181] = ~in[181];
  assign inbar[182] = ~in[182];
  assign inbar[183] = ~in[183];
  assign inbar[184] = ~in[184];
  assign inbar[185] = ~in[185];
  assign inbar[186] = ~in[186];
  assign inbar[187] = ~in[187];
  assign inbar[188] = ~in[188];
  assign inbar[189] = ~in[189];
  assign inbar[190] = ~in[190];
  assign inbar[191] = ~in[191];
  assign inbar[192] = ~in[192];
  assign inbar[193] = ~in[193];
  assign inbar[194] = ~in[194];
  assign inbar[195] = ~in[195];
  assign inbar[196] = ~in[196];
  assign inbar[197] = ~in[197];
  assign inbar[198] = ~in[198];
  assign inbar[199] = ~in[199];
  assign inbar[200] = ~in[200];
  assign inbar[201] = ~in[201];
  assign inbar[202] = ~in[202];
  assign inbar[203] = ~in[203];
  assign inbar[204] = ~in[204];
  assign inbar[205] = ~in[205];
  assign inbar[206] = ~in[206];
  assign inbar[207] = ~in[207];
  assign inbar[208] = ~in[208];
  assign inbar[209] = ~in[209];
  assign inbar[210] = ~in[210];
  assign inbar[211] = ~in[211];
  assign inbar[212] = ~in[212];
  assign inbar[213] = ~in[213];
  assign inbar[214] = ~in[214];
  assign inbar[215] = ~in[215];
  assign inbar[216] = ~in[216];
  assign inbar[217] = ~in[217];
  assign inbar[218] = ~in[218];
  assign inbar[219] = ~in[219];
  assign inbar[220] = ~in[220];
  assign inbar[221] = ~in[221];
  assign inbar[222] = ~in[222];
  assign inbar[223] = ~in[223];
  assign inbar[224] = ~in[224];
  assign inbar[225] = ~in[225];
  assign inbar[226] = ~in[226];
  assign inbar[227] = ~in[227];
  assign inbar[228] = ~in[228];
  assign inbar[229] = ~in[229];
  assign inbar[230] = ~in[230];
  assign inbar[231] = ~in[231];
  assign inbar[232] = ~in[232];
  assign inbar[233] = ~in[233];
  assign inbar[234] = ~in[234];
  assign inbar[235] = ~in[235];
  assign inbar[236] = ~in[236];
  assign inbar[237] = ~in[237];
  assign inbar[238] = ~in[238];
  assign inbar[239] = ~in[239];
  assign inbar[240] = ~in[240];
  assign inbar[241] = ~in[241];
  assign inbar[242] = ~in[242];
  assign inbar[243] = ~in[243];
  assign inbar[244] = ~in[244];
  assign inbar[245] = ~in[245];
  assign inbar[246] = ~in[246];
  assign inbar[247] = ~in[247];
  assign inbar[248] = ~in[248];
  assign inbar[249] = ~in[249];
  assign inbar[250] = ~in[250];
  assign inbar[251] = ~in[251];
  assign inbar[252] = ~in[252];
  assign inbar[253] = ~in[253];
  assign inbar[254] = ~in[254];
  assign inbar[255] = ~in[255];
  //input_done

  output [7:0] out;
  reg [7:0] outbar;
  //output_done

  wire   in_81, in_80, in_79, in_78, in_77, in_76, in_75, in_74, in_73, in_72,
         in_71, in_70, in_69, in_68, in_67, in_66, in_65, in_64, in_63, in_62,
         in_61, in_60, in_59, in_58, in_57, in_56, in_55, in_54, in_53, in_52,
         in_51, in_50, in_49, in_48, in_47, in_46, in_45, in_44, in_43, in_42,
         in_41, in_40, in_39, in_38, in_37, in_36, in_35, in_34, in_33, in_32,
         in_31, in_30, in_29, in_28, in_27, in_26, in_25, in_24, in_23, in_22,
         in_21, in_20, in_19, in_18, in_17, in_16, in_15, in_14, in_13, in_12,
         in_11, in_10, in_9, in_8, in_7, in_6, in_5, in_4, in_3, in_2, in_1,
         in_0, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972;
  wire in_81bar, in_80bar, in_79bar, in_78bar, in_77bar, in_76bar, in_75bar, in_74bar, in_73bar, in_72bar, in_71bar, in_70bar, in_69bar, in_68bar, in_67bar, in_66bar, in_65bar, in_64bar, in_63bar, in_62bar, in_61bar, in_60bar, in_59bar, in_58bar, in_57bar, in_56bar, in_55bar, in_54bar, in_53bar, in_52bar, in_51bar, in_50bar, in_49bar, in_48bar, in_47bar, in_46bar, in_45bar, in_44bar, in_43bar, in_42bar, in_41bar, in_40bar, in_39bar, in_38bar, in_37bar, in_36bar, in_35bar, in_34bar, in_33bar, in_32bar, in_31bar, in_30bar, in_29bar, in_28bar, in_27bar, in_26bar, in_25bar, in_24bar, in_23bar, in_22bar, in_21bar, in_20bar, in_19bar, in_18bar, in_17bar, in_16bar, in_15bar, in_14bar, in_13bar, in_12bar, in_11bar, in_10bar, in_9bar, in_8bar, in_7bar, in_6bar, in_5bar, in_4bar, in_3bar, in_2bar, in_1bar, in_0bar, n487bar, n488bar, n489bar, n490bar, n491bar, n492bar, n493bar, n494bar, n495bar, n496bar, n497bar, n498bar, n499bar, n500bar, n501bar, n502bar, n503bar, n504bar, n505bar, n506bar, n507bar, n508bar, n509bar, n510bar, n511bar, n512bar, n513bar, n514bar, n515bar, n516bar, n517bar, n518bar, n519bar, n520bar, n521bar, n522bar, n523bar, n524bar, n525bar, n526bar, n527bar, n528bar, n529bar, n530bar, n531bar, n532bar, n533bar, n534bar, n535bar, n536bar, n537bar, n538bar, n539bar, n540bar, n541bar, n542bar, n543bar, n544bar, n545bar, n546bar, n547bar, n548bar, n549bar, n550bar, n551bar, n552bar, n553bar, n554bar, n555bar, n556bar, n557bar, n558bar, n559bar, n560bar, n561bar, n562bar, n563bar, n564bar, n565bar, n566bar, n567bar, n568bar, n569bar, n570bar, n571bar, n572bar, n573bar, n574bar, n575bar, n576bar, n577bar, n578bar, n579bar, n580bar, n581bar, n582bar, n583bar, n584bar, n585bar, n586bar, n587bar, n588bar, n589bar, n590bar, n591bar, n592bar, n593bar, n594bar, n595bar, n596bar, n597bar, n598bar, n599bar, n600bar, n601bar, n602bar, n603bar, n604bar, n605bar, n606bar, n607bar, n608bar, n609bar, n610bar, n611bar, n612bar, n613bar, n614bar, n615bar, n616bar, n617bar, n618bar, n619bar, n620bar, n621bar, n622bar, n623bar, n624bar, n625bar, n626bar, n627bar, n628bar, n629bar, n630bar, n631bar, n632bar, n633bar, n634bar, n635bar, n636bar, n637bar, n638bar, n639bar, n640bar, n641bar, n642bar, n643bar, n644bar, n645bar, n646bar, n647bar, n648bar, n649bar, n650bar, n651bar, n652bar, n653bar, n654bar, n655bar, n656bar, n657bar, n658bar, n659bar, n660bar, n661bar, n662bar, n663bar, n664bar, n665bar, n666bar, n667bar, n668bar, n669bar, n670bar, n671bar, n672bar, n673bar, n674bar, n675bar, n676bar, n677bar, n678bar, n679bar, n680bar, n681bar, n682bar, n683bar, n684bar, n685bar, n686bar, n687bar, n688bar, n689bar, n690bar, n691bar, n692bar, n693bar, n694bar, n695bar, n696bar, n697bar, n698bar, n699bar, n700bar, n701bar, n702bar, n703bar, n704bar, n705bar, n706bar, n707bar, n708bar, n709bar, n710bar, n711bar, n712bar, n713bar, n714bar, n715bar, n716bar, n717bar, n718bar, n719bar, n720bar, n721bar, n722bar, n723bar, n724bar, n725bar, n726bar, n727bar, n728bar, n729bar, n730bar, n731bar, n732bar, n733bar, n734bar, n735bar, n736bar, n737bar, n738bar, n739bar, n740bar, n741bar, n742bar, n743bar, n744bar, n745bar, n746bar, n747bar, n748bar, n749bar, n750bar, n751bar, n752bar, n753bar, n754bar, n755bar, n756bar, n757bar, n758bar, n759bar, n760bar, n761bar, n762bar, n763bar, n764bar, n765bar, n766bar, n767bar, n768bar, n769bar, n770bar, n771bar, n772bar, n773bar, n774bar, n775bar, n776bar, n777bar, n778bar, n779bar, n780bar, n781bar, n782bar, n783bar, n784bar, n785bar, n786bar, n787bar, n788bar, n789bar, n790bar, n791bar, n792bar, n793bar, n794bar, n795bar, n796bar, n797bar, n798bar, n799bar, n800bar, n801bar, n802bar, n803bar, n804bar, n805bar, n806bar, n807bar, n808bar, n809bar, n810bar, n811bar, n812bar, n813bar, n814bar, n815bar, n816bar, n817bar, n818bar, n819bar, n820bar, n821bar, n822bar, n823bar, n824bar, n825bar, n826bar, n827bar, n828bar, n829bar, n830bar, n831bar, n832bar, n833bar, n834bar, n835bar, n836bar, n837bar, n838bar, n839bar, n840bar, n841bar, n842bar, n843bar, n844bar, n845bar, n846bar, n847bar, n848bar, n849bar, n850bar, n851bar, n852bar, n853bar, n854bar, n855bar, n856bar, n857bar, n858bar, n859bar, n860bar, n861bar, n862bar, n863bar, n864bar, n865bar, n866bar, n867bar, n868bar, n869bar, n870bar, n871bar, n872bar, n873bar, n874bar, n875bar, n876bar, n877bar, n878bar, n879bar, n880bar, n881bar, n882bar, n883bar, n884bar, n885bar, n886bar, n887bar, n888bar, n889bar, n890bar, n891bar, n892bar, n893bar, n894bar, n895bar, n896bar, n897bar, n898bar, n899bar, n900bar, n901bar, n902bar, n903bar, n904bar, n905bar, n906bar, n907bar, n908bar, n909bar, n910bar, n911bar, n912bar, n913bar, n914bar, n915bar, n916bar, n917bar, n918bar, n919bar, n920bar, n921bar, n922bar, n923bar, n924bar, n925bar, n926bar, n927bar, n928bar, n929bar, n930bar, n931bar, n932bar, n933bar, n934bar, n935bar, n936bar, n937bar, n938bar, n939bar, n940bar, n941bar, n942bar, n943bar, n944bar, n945bar, n946bar, n947bar, n948bar, n949bar, n950bar, n951bar, n952bar, n953bar, n954bar, n955bar, n956bar, n957bar, n958bar, n959bar, n960bar, n961bar, n962bar, n963bar, n964bar, n965bar, n966bar, n967bar, n968bar, n969bar, n970bar, n971bar, n972bar;
  //wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];

  OR2_X1 U1 ( .A1(n972), .A2(n971), .ZN(out[7]) );
  AND2_X1 U1bar ( .A1(n972bar), .A2(n971bar), .ZN(outbar[7]);
  OR2_X1 U2 ( .A1(n970), .A2(n969), .ZN(n971) );
  AND2_X1 U2bar ( .A1(n970bar), .A2(n969bar), .ZN(n971bar);
  OR2_X1 U3 ( .A1(n968), .A2(n967), .ZN(n969) );
  AND2_X1 U3bar ( .A1(n968bar), .A2(n967bar), .ZN(n969bar);
  OR2_X1 U4 ( .A1(n966), .A2(n965), .ZN(n967) );
  AND2_X1 U4bar ( .A1(n966bar), .A2(n965bar), .ZN(n967bar);
  OR2_X1 U5 ( .A1(n964), .A2(n963), .ZN(n968) );
  AND2_X1 U5bar ( .A1(n964bar), .A2(n963bar), .ZN(n968bar);
  OR2_X1 U6 ( .A1(in[116]), .A2(n962), .ZN(n963) );
  AND2_X1 U6bar ( .A1(inbar[116]), .A2(n962bar), .ZN(n963bar);
  OR2_X1 U7 ( .A1(n961), .A2(n960), .ZN(n970) );
  AND2_X1 U7bar ( .A1(n961bar), .A2(n960bar), .ZN(n970bar);
  OR2_X1 U8 ( .A1(in[150]), .A2(in[127]), .ZN(n960) );
  AND2_X1 U8bar ( .A1(inbar[150]), .A2(inbar[127]), .ZN(n960bar);
  OR2_X1 U9 ( .A1(in[160]), .A2(n959), .ZN(n961) );
  AND2_X1 U9bar ( .A1(inbar[160]), .A2(n959bar), .ZN(n961bar);
  OR2_X1 U10 ( .A1(in[252]), .A2(in[168]), .ZN(n959) );
  AND2_X1 U10bar ( .A1(inbar[252]), .A2(inbar[168]), .ZN(n959bar);
  OR2_X1 U11 ( .A1(n958), .A2(n957), .ZN(n972) );
  AND2_X1 U11bar ( .A1(n958bar), .A2(n957bar), .ZN(n972bar);
  OR2_X1 U12 ( .A1(n956), .A2(n955), .ZN(n957) );
  AND2_X1 U12bar ( .A1(n956bar), .A2(n955bar), .ZN(n957bar);
  OR2_X1 U13 ( .A1(in_17), .A2(in[96]), .ZN(n955) );
  AND2_X1 U13bar ( .A1(in_17bar), .A2(inbar[96]), .ZN(n955bar);
  OR2_X1 U14 ( .A1(in_23), .A2(n954), .ZN(n956) );
  AND2_X1 U14bar ( .A1(in_23bar), .A2(n954bar), .ZN(n956bar);
  OR2_X1 U15 ( .A1(in_31), .A2(in_26), .ZN(n954) );
  AND2_X1 U15bar ( .A1(in_31bar), .A2(in_26bar), .ZN(n954bar);
  OR2_X1 U16 ( .A1(n953), .A2(n952), .ZN(n958) );
  AND2_X1 U16bar ( .A1(n953bar), .A2(n952bar), .ZN(n958bar);
  OR2_X1 U17 ( .A1(in_58), .A2(in_4), .ZN(n952) );
  AND2_X1 U17bar ( .A1(in_58bar), .A2(in_4bar), .ZN(n952bar);
  OR2_X1 U18 ( .A1(in_59), .A2(n951), .ZN(n953) );
  AND2_X1 U18bar ( .A1(in_59bar), .A2(n951bar), .ZN(n953bar);
  OR2_X1 U19 ( .A1(in_71), .A2(in_62), .ZN(n951) );
  AND2_X1 U19bar ( .A1(in_71bar), .A2(in_62bar), .ZN(n951bar);
  OR2_X1 U20 ( .A1(n950), .A2(n949), .ZN(out[6]) );
  AND2_X1 U20bar ( .A1(n950bar), .A2(n949bar), .ZN(outbar[6]);
  OR2_X1 U21 ( .A1(n948), .A2(n947), .ZN(n949) );
  AND2_X1 U21bar ( .A1(n948bar), .A2(n947bar), .ZN(n949bar);
  OR2_X1 U22 ( .A1(n946), .A2(n945), .ZN(n947) );
  AND2_X1 U22bar ( .A1(n946bar), .A2(n945bar), .ZN(n947bar);
  OR2_X1 U23 ( .A1(n944), .A2(n943), .ZN(n945) );
  AND2_X1 U23bar ( .A1(n944bar), .A2(n943bar), .ZN(n945bar);
  OR2_X1 U24 ( .A1(n942), .A2(n941), .ZN(n946) );
  AND2_X1 U24bar ( .A1(n942bar), .A2(n941bar), .ZN(n946bar);
  OR2_X1 U25 ( .A1(in[101]), .A2(n940), .ZN(n941) );
  AND2_X1 U25bar ( .A1(inbar[101]), .A2(n940bar), .ZN(n941bar);
  OR2_X1 U26 ( .A1(n939), .A2(n938), .ZN(n948) );
  AND2_X1 U26bar ( .A1(n939bar), .A2(n938bar), .ZN(n948bar);
  OR2_X1 U27 ( .A1(in[114]), .A2(in[104]), .ZN(n938) );
  AND2_X1 U27bar ( .A1(inbar[114]), .A2(inbar[104]), .ZN(n938bar);
  OR2_X1 U28 ( .A1(in[128]), .A2(n937), .ZN(n939) );
  AND2_X1 U28bar ( .A1(inbar[128]), .A2(n937bar), .ZN(n939bar);
  OR2_X1 U29 ( .A1(in[136]), .A2(in[134]), .ZN(n937) );
  AND2_X1 U29bar ( .A1(inbar[136]), .A2(inbar[134]), .ZN(n937bar);
  OR2_X1 U30 ( .A1(n936), .A2(n935), .ZN(n950) );
  AND2_X1 U30bar ( .A1(n936bar), .A2(n935bar), .ZN(n950bar);
  OR2_X1 U31 ( .A1(n934), .A2(n933), .ZN(n935) );
  AND2_X1 U31bar ( .A1(n934bar), .A2(n933bar), .ZN(n935bar);
  OR2_X1 U32 ( .A1(in[177]), .A2(in[164]), .ZN(n933) );
  AND2_X1 U32bar ( .A1(inbar[177]), .A2(inbar[164]), .ZN(n933bar);
  OR2_X1 U33 ( .A1(in[212]), .A2(n932), .ZN(n934) );
  AND2_X1 U33bar ( .A1(inbar[212]), .A2(n932bar), .ZN(n934bar);
  OR2_X1 U34 ( .A1(in[248]), .A2(in[221]), .ZN(n932) );
  AND2_X1 U34bar ( .A1(inbar[248]), .A2(inbar[221]), .ZN(n932bar);
  OR2_X1 U35 ( .A1(n931), .A2(n930), .ZN(n936) );
  AND2_X1 U35bar ( .A1(n931bar), .A2(n930bar), .ZN(n936bar);
  OR2_X1 U36 ( .A1(in_18), .A2(in[93]), .ZN(n930) );
  AND2_X1 U36bar ( .A1(in_18bar), .A2(inbar[93]), .ZN(n930bar);
  OR2_X1 U37 ( .A1(in_31), .A2(n929), .ZN(n931) );
  AND2_X1 U37bar ( .A1(in_31bar), .A2(n929bar), .ZN(n931bar);
  OR2_X1 U38 ( .A1(in_7), .A2(in_39), .ZN(n929) );
  AND2_X1 U38bar ( .A1(in_7bar), .A2(in_39bar), .ZN(n929bar);
  OR2_X1 U39 ( .A1(n928), .A2(n927), .ZN(out[5]) );
  AND2_X1 U39bar ( .A1(n928bar), .A2(n927bar), .ZN(outbar[5]);
  OR2_X1 U40 ( .A1(n926), .A2(n925), .ZN(n927) );
  AND2_X1 U40bar ( .A1(n926bar), .A2(n925bar), .ZN(n927bar);
  OR2_X1 U41 ( .A1(n924), .A2(n923), .ZN(n925) );
  AND2_X1 U41bar ( .A1(n924bar), .A2(n923bar), .ZN(n925bar);
  OR2_X1 U42 ( .A1(n922), .A2(n921), .ZN(n923) );
  AND2_X1 U42bar ( .A1(n922bar), .A2(n921bar), .ZN(n923bar);
  OR2_X1 U43 ( .A1(n940), .A2(n920), .ZN(n924) );
  AND2_X1 U43bar ( .A1(n940bar), .A2(n920bar), .ZN(n924bar);
  OR2_X1 U44 ( .A1(in[111]), .A2(n919), .ZN(n920) );
  AND2_X1 U44bar ( .A1(inbar[111]), .A2(n919bar), .ZN(n920bar);
  OR2_X1 U45 ( .A1(n918), .A2(n917), .ZN(n940) );
  AND2_X1 U45bar ( .A1(n918bar), .A2(n917bar), .ZN(n940bar);
  OR2_X1 U46 ( .A1(n916), .A2(n915), .ZN(n917) );
  AND2_X1 U46bar ( .A1(n916bar), .A2(n915bar), .ZN(n917bar);
  OR2_X1 U47 ( .A1(n914), .A2(n913), .ZN(n915) );
  AND2_X1 U47bar ( .A1(n914bar), .A2(n913bar), .ZN(n915bar);
  OR2_X1 U48 ( .A1(in[140]), .A2(in[131]), .ZN(n913) );
  AND2_X1 U48bar ( .A1(inbar[140]), .A2(inbar[131]), .ZN(n913bar);
  OR2_X1 U49 ( .A1(in[160]), .A2(in[144]), .ZN(n914) );
  AND2_X1 U49bar ( .A1(inbar[160]), .A2(inbar[144]), .ZN(n914bar);
  OR2_X1 U50 ( .A1(n912), .A2(n911), .ZN(n916) );
  AND2_X1 U50bar ( .A1(n912bar), .A2(n911bar), .ZN(n916bar);
  OR2_X1 U51 ( .A1(in[179]), .A2(in[174]), .ZN(n911) );
  AND2_X1 U51bar ( .A1(inbar[179]), .A2(inbar[174]), .ZN(n911bar);
  OR2_X1 U52 ( .A1(in[188]), .A2(in[184]), .ZN(n912) );
  AND2_X1 U52bar ( .A1(inbar[188]), .A2(inbar[184]), .ZN(n912bar);
  OR2_X1 U53 ( .A1(n910), .A2(n909), .ZN(n918) );
  AND2_X1 U53bar ( .A1(n910bar), .A2(n909bar), .ZN(n918bar);
  OR2_X1 U54 ( .A1(n908), .A2(n907), .ZN(n909) );
  AND2_X1 U54bar ( .A1(n908bar), .A2(n907bar), .ZN(n909bar);
  OR2_X1 U55 ( .A1(in[216]), .A2(in[200]), .ZN(n907) );
  AND2_X1 U55bar ( .A1(inbar[216]), .A2(inbar[200]), .ZN(n907bar);
  OR2_X1 U56 ( .A1(in[228]), .A2(in[224]), .ZN(n908) );
  AND2_X1 U56bar ( .A1(inbar[228]), .A2(inbar[224]), .ZN(n908bar);
  OR2_X1 U57 ( .A1(n906), .A2(n905), .ZN(n910) );
  AND2_X1 U57bar ( .A1(n906bar), .A2(n905bar), .ZN(n910bar);
  OR2_X1 U58 ( .A1(in[247]), .A2(in[235]), .ZN(n905) );
  AND2_X1 U58bar ( .A1(inbar[247]), .A2(inbar[235]), .ZN(n905bar);
  OR2_X1 U59 ( .A1(in_42), .A2(in[83]), .ZN(n906) );
  AND2_X1 U59bar ( .A1(in_42bar), .A2(inbar[83]), .ZN(n906bar);
  OR2_X1 U60 ( .A1(n904), .A2(n903), .ZN(n926) );
  AND2_X1 U60bar ( .A1(n904bar), .A2(n903bar), .ZN(n926bar);
  OR2_X1 U61 ( .A1(in[166]), .A2(in[123]), .ZN(n903) );
  AND2_X1 U61bar ( .A1(inbar[166]), .A2(inbar[123]), .ZN(n903bar);
  OR2_X1 U62 ( .A1(in[170]), .A2(n902), .ZN(n904) );
  AND2_X1 U62bar ( .A1(inbar[170]), .A2(n902bar), .ZN(n904bar);
  OR2_X1 U63 ( .A1(in[194]), .A2(in[183]), .ZN(n902) );
  AND2_X1 U63bar ( .A1(inbar[194]), .A2(inbar[183]), .ZN(n902bar);
  OR2_X1 U64 ( .A1(n901), .A2(n900), .ZN(n928) );
  AND2_X1 U64bar ( .A1(n901bar), .A2(n900bar), .ZN(n928bar);
  OR2_X1 U65 ( .A1(n899), .A2(n898), .ZN(n900) );
  AND2_X1 U65bar ( .A1(n899bar), .A2(n898bar), .ZN(n900bar);
  OR2_X1 U66 ( .A1(in[241]), .A2(in[238]), .ZN(n898) );
  AND2_X1 U66bar ( .A1(inbar[241]), .A2(inbar[238]), .ZN(n898bar);
  OR2_X1 U67 ( .A1(in[250]), .A2(n897), .ZN(n899) );
  AND2_X1 U67bar ( .A1(inbar[250]), .A2(n897bar), .ZN(n899bar);
  OR2_X1 U68 ( .A1(in_24), .A2(in[84]), .ZN(n897) );
  AND2_X1 U68bar ( .A1(in_24bar), .A2(inbar[84]), .ZN(n897bar);
  OR2_X1 U69 ( .A1(n896), .A2(n895), .ZN(n901) );
  AND2_X1 U69bar ( .A1(n896bar), .A2(n895bar), .ZN(n901bar);
  OR2_X1 U70 ( .A1(in_41), .A2(in_29), .ZN(n895) );
  AND2_X1 U70bar ( .A1(in_41bar), .A2(in_29bar), .ZN(n895bar);
  OR2_X1 U71 ( .A1(in_66), .A2(n894), .ZN(n896) );
  AND2_X1 U71bar ( .A1(in_66bar), .A2(n894bar), .ZN(n896bar);
  OR2_X1 U72 ( .A1(in_76), .A2(in_71), .ZN(n894) );
  AND2_X1 U72bar ( .A1(in_76bar), .A2(in_71bar), .ZN(n894bar);
  OR2_X1 U73 ( .A1(n893), .A2(n892), .ZN(out[4]) );
  AND2_X1 U73bar ( .A1(n893bar), .A2(n892bar), .ZN(outbar[4]);
  OR2_X1 U74 ( .A1(n891), .A2(n890), .ZN(n892) );
  AND2_X1 U74bar ( .A1(n891bar), .A2(n890bar), .ZN(n892bar);
  OR2_X1 U75 ( .A1(n889), .A2(n888), .ZN(n890) );
  AND2_X1 U75bar ( .A1(n889bar), .A2(n888bar), .ZN(n890bar);
  OR2_X1 U76 ( .A1(n922), .A2(n887), .ZN(n888) );
  AND2_X1 U76bar ( .A1(n922bar), .A2(n887bar), .ZN(n888bar);
  OR2_X1 U77 ( .A1(n886), .A2(n885), .ZN(n922) );
  AND2_X1 U77bar ( .A1(n886bar), .A2(n885bar), .ZN(n922bar);
  OR2_X1 U78 ( .A1(n884), .A2(n883), .ZN(n885) );
  AND2_X1 U78bar ( .A1(n884bar), .A2(n883bar), .ZN(n885bar);
  OR2_X1 U79 ( .A1(n882), .A2(n881), .ZN(n883) );
  AND2_X1 U79bar ( .A1(n882bar), .A2(n881bar), .ZN(n883bar);
  OR2_X1 U80 ( .A1(in[118]), .A2(in[109]), .ZN(n881) );
  AND2_X1 U80bar ( .A1(inbar[118]), .A2(inbar[109]), .ZN(n881bar);
  OR2_X1 U81 ( .A1(in[139]), .A2(in[120]), .ZN(n882) );
  AND2_X1 U81bar ( .A1(inbar[139]), .A2(inbar[120]), .ZN(n882bar);
  OR2_X1 U82 ( .A1(n880), .A2(n879), .ZN(n884) );
  AND2_X1 U82bar ( .A1(n880bar), .A2(n879bar), .ZN(n884bar);
  OR2_X1 U83 ( .A1(in[198]), .A2(in[154]), .ZN(n879) );
  AND2_X1 U83bar ( .A1(inbar[198]), .A2(inbar[154]), .ZN(n879bar);
  OR2_X1 U84 ( .A1(in[210]), .A2(in[205]), .ZN(n880) );
  AND2_X1 U84bar ( .A1(inbar[210]), .A2(inbar[205]), .ZN(n880bar);
  OR2_X1 U85 ( .A1(n878), .A2(n877), .ZN(n886) );
  AND2_X1 U85bar ( .A1(n878bar), .A2(n877bar), .ZN(n886bar);
  OR2_X1 U86 ( .A1(n876), .A2(n875), .ZN(n877) );
  AND2_X1 U86bar ( .A1(n876bar), .A2(n875bar), .ZN(n877bar);
  OR2_X1 U87 ( .A1(in[219]), .A2(in[217]), .ZN(n875) );
  AND2_X1 U87bar ( .A1(inbar[219]), .A2(inbar[217]), .ZN(n875bar);
  OR2_X1 U88 ( .A1(in[86]), .A2(in[252]), .ZN(n876) );
  AND2_X1 U88bar ( .A1(inbar[86]), .A2(inbar[252]), .ZN(n876bar);
  OR2_X1 U89 ( .A1(n874), .A2(n873), .ZN(n878) );
  AND2_X1 U89bar ( .A1(n874bar), .A2(n873bar), .ZN(n878bar);
  OR2_X1 U90 ( .A1(in_40), .A2(in[91]), .ZN(n873) );
  AND2_X1 U90bar ( .A1(in_40bar), .A2(inbar[91]), .ZN(n873bar);
  OR2_X1 U91 ( .A1(in_8), .A2(in_46), .ZN(n874) );
  AND2_X1 U91bar ( .A1(in_8bar), .A2(in_46bar), .ZN(n874bar);
  OR2_X1 U92 ( .A1(n872), .A2(n871), .ZN(n889) );
  AND2_X1 U92bar ( .A1(n872bar), .A2(n871bar), .ZN(n889bar);
  OR2_X1 U93 ( .A1(in[117]), .A2(n943), .ZN(n871) );
  AND2_X1 U93bar ( .A1(inbar[117]), .A2(n943bar), .ZN(n871bar);
  OR2_X1 U94 ( .A1(n870), .A2(n869), .ZN(n943) );
  AND2_X1 U94bar ( .A1(n870bar), .A2(n869bar), .ZN(n943bar);
  OR2_X1 U95 ( .A1(n868), .A2(n867), .ZN(n869) );
  AND2_X1 U95bar ( .A1(n868bar), .A2(n867bar), .ZN(n869bar);
  OR2_X1 U96 ( .A1(n866), .A2(n865), .ZN(n867) );
  AND2_X1 U96bar ( .A1(n866bar), .A2(n865bar), .ZN(n867bar);
  OR2_X1 U97 ( .A1(n864), .A2(n863), .ZN(n865) );
  AND2_X1 U97bar ( .A1(n864bar), .A2(n863bar), .ZN(n865bar);
  OR2_X1 U98 ( .A1(in[108]), .A2(n919), .ZN(n866) );
  AND2_X1 U98bar ( .A1(inbar[108]), .A2(n919bar), .ZN(n866bar);
  OR2_X1 U99 ( .A1(n862), .A2(n861), .ZN(n919) );
  AND2_X1 U99bar ( .A1(n862bar), .A2(n861bar), .ZN(n919bar);
  OR2_X1 U100 ( .A1(n860), .A2(n859), .ZN(n861) );
  AND2_X1 U100bar ( .A1(n860bar), .A2(n859bar), .ZN(n861bar);
  OR2_X1 U101 ( .A1(n858), .A2(n857), .ZN(n859) );
  AND2_X1 U101bar ( .A1(n858bar), .A2(n857bar), .ZN(n859bar);
  OR2_X1 U102 ( .A1(in[119]), .A2(in[105]), .ZN(n857) );
  AND2_X1 U102bar ( .A1(inbar[119]), .A2(inbar[105]), .ZN(n857bar);
  OR2_X1 U103 ( .A1(in[186]), .A2(in[175]), .ZN(n858) );
  AND2_X1 U103bar ( .A1(inbar[186]), .A2(inbar[175]), .ZN(n858bar);
  OR2_X1 U104 ( .A1(n856), .A2(n855), .ZN(n860) );
  AND2_X1 U104bar ( .A1(n856bar), .A2(n855bar), .ZN(n860bar);
  OR2_X1 U105 ( .A1(in[202]), .A2(in[193]), .ZN(n855) );
  AND2_X1 U105bar ( .A1(inbar[202]), .A2(inbar[193]), .ZN(n855bar);
  OR2_X1 U106 ( .A1(in[225]), .A2(in[208]), .ZN(n856) );
  AND2_X1 U106bar ( .A1(inbar[225]), .A2(inbar[208]), .ZN(n856bar);
  OR2_X1 U107 ( .A1(n854), .A2(n853), .ZN(n862) );
  AND2_X1 U107bar ( .A1(n854bar), .A2(n853bar), .ZN(n862bar);
  OR2_X1 U108 ( .A1(n852), .A2(n851), .ZN(n853) );
  AND2_X1 U108bar ( .A1(n852bar), .A2(n851bar), .ZN(n853bar);
  OR2_X1 U109 ( .A1(in_1), .A2(in[85]), .ZN(n851) );
  AND2_X1 U109bar ( .A1(in_1bar), .A2(inbar[85]), .ZN(n851bar);
  OR2_X1 U110 ( .A1(in_23), .A2(in_19), .ZN(n852) );
  AND2_X1 U110bar ( .A1(in_23bar), .A2(in_19bar), .ZN(n852bar);
  OR2_X1 U111 ( .A1(n850), .A2(n849), .ZN(n854) );
  AND2_X1 U111bar ( .A1(n850bar), .A2(n849bar), .ZN(n854bar);
  OR2_X1 U112 ( .A1(in_43), .A2(in_33), .ZN(n849) );
  AND2_X1 U112bar ( .A1(in_43bar), .A2(in_33bar), .ZN(n849bar);
  OR2_X1 U113 ( .A1(in_63), .A2(in_44), .ZN(n850) );
  AND2_X1 U113bar ( .A1(in_63bar), .A2(in_44bar), .ZN(n850bar);
  OR2_X1 U114 ( .A1(n848), .A2(n847), .ZN(n868) );
  AND2_X1 U114bar ( .A1(n848bar), .A2(n847bar), .ZN(n868bar);
  OR2_X1 U115 ( .A1(in[141]), .A2(in[112]), .ZN(n847) );
  AND2_X1 U115bar ( .A1(inbar[141]), .A2(inbar[112]), .ZN(n847bar);
  OR2_X1 U116 ( .A1(in[147]), .A2(n846), .ZN(n848) );
  AND2_X1 U116bar ( .A1(inbar[147]), .A2(n846bar), .ZN(n848bar);
  OR2_X1 U117 ( .A1(in[181]), .A2(in[167]), .ZN(n846) );
  AND2_X1 U117bar ( .A1(inbar[181]), .A2(inbar[167]), .ZN(n846bar);
  OR2_X1 U118 ( .A1(n845), .A2(n844), .ZN(n870) );
  AND2_X1 U118bar ( .A1(n845bar), .A2(n844bar), .ZN(n870bar);
  OR2_X1 U119 ( .A1(n843), .A2(n842), .ZN(n844) );
  AND2_X1 U119bar ( .A1(n843bar), .A2(n842bar), .ZN(n844bar);
  OR2_X1 U120 ( .A1(in[229]), .A2(in[201]), .ZN(n842) );
  AND2_X1 U120bar ( .A1(inbar[229]), .A2(inbar[201]), .ZN(n842bar);
  OR2_X1 U121 ( .A1(in[237]), .A2(n841), .ZN(n843) );
  AND2_X1 U121bar ( .A1(inbar[237]), .A2(n841bar), .ZN(n843bar);
  OR2_X1 U122 ( .A1(in[94]), .A2(in[253]), .ZN(n841) );
  AND2_X1 U122bar ( .A1(inbar[94]), .A2(inbar[253]), .ZN(n841bar);
  OR2_X1 U123 ( .A1(n840), .A2(n839), .ZN(n845) );
  AND2_X1 U123bar ( .A1(n840bar), .A2(n839bar), .ZN(n845bar);
  OR2_X1 U124 ( .A1(in_21), .A2(in[96]), .ZN(n839) );
  AND2_X1 U124bar ( .A1(in_21bar), .A2(inbar[96]), .ZN(n839bar);
  OR2_X1 U125 ( .A1(in_25), .A2(n838), .ZN(n840) );
  AND2_X1 U125bar ( .A1(in_25bar), .A2(n838bar), .ZN(n840bar);
  OR2_X1 U126 ( .A1(in_81), .A2(in_45), .ZN(n838) );
  AND2_X1 U126bar ( .A1(in_81bar), .A2(in_45bar), .ZN(n838bar);
  OR2_X1 U127 ( .A1(n837), .A2(n836), .ZN(n891) );
  AND2_X1 U127bar ( .A1(n837bar), .A2(n836bar), .ZN(n891bar);
  OR2_X1 U128 ( .A1(in[142]), .A2(in[124]), .ZN(n836) );
  AND2_X1 U128bar ( .A1(inbar[142]), .A2(inbar[124]), .ZN(n836bar);
  OR2_X1 U129 ( .A1(in[150]), .A2(n835), .ZN(n837) );
  AND2_X1 U129bar ( .A1(inbar[150]), .A2(n835bar), .ZN(n837bar);
  OR2_X1 U130 ( .A1(in[172]), .A2(in[155]), .ZN(n835) );
  AND2_X1 U130bar ( .A1(inbar[172]), .A2(inbar[155]), .ZN(n835bar);
  OR2_X1 U131 ( .A1(n834), .A2(n833), .ZN(n893) );
  AND2_X1 U131bar ( .A1(n834bar), .A2(n833bar), .ZN(n893bar);
  OR2_X1 U132 ( .A1(n832), .A2(n831), .ZN(n833) );
  AND2_X1 U132bar ( .A1(n832bar), .A2(n831bar), .ZN(n833bar);
  OR2_X1 U133 ( .A1(in[196]), .A2(in[173]), .ZN(n831) );
  AND2_X1 U133bar ( .A1(inbar[196]), .A2(inbar[173]), .ZN(n831bar);
  OR2_X1 U134 ( .A1(in[222]), .A2(n830), .ZN(n832) );
  AND2_X1 U134bar ( .A1(inbar[222]), .A2(n830bar), .ZN(n832bar);
  OR2_X1 U135 ( .A1(in[227]), .A2(in[226]), .ZN(n830) );
  AND2_X1 U135bar ( .A1(inbar[227]), .A2(inbar[226]), .ZN(n830bar);
  OR2_X1 U136 ( .A1(n829), .A2(n828), .ZN(n834) );
  AND2_X1 U136bar ( .A1(n829bar), .A2(n828bar), .ZN(n834bar);
  OR2_X1 U137 ( .A1(in[249]), .A2(in[231]), .ZN(n828) );
  AND2_X1 U137bar ( .A1(inbar[249]), .A2(inbar[231]), .ZN(n828bar);
  OR2_X1 U138 ( .A1(in_28), .A2(n827), .ZN(n829) );
  AND2_X1 U138bar ( .A1(in_28bar), .A2(n827bar), .ZN(n829bar);
  OR2_X1 U139 ( .A1(in_52), .A2(in_47), .ZN(n827) );
  AND2_X1 U139bar ( .A1(in_52bar), .A2(in_47bar), .ZN(n827bar);
  OR2_X1 U140 ( .A1(n826), .A2(n825), .ZN(out[3]) );
  AND2_X1 U140bar ( .A1(n826bar), .A2(n825bar), .ZN(outbar[3]);
  OR2_X1 U141 ( .A1(n824), .A2(n823), .ZN(n825) );
  AND2_X1 U141bar ( .A1(n824bar), .A2(n823bar), .ZN(n825bar);
  OR2_X1 U142 ( .A1(n822), .A2(n821), .ZN(n823) );
  AND2_X1 U142bar ( .A1(n822bar), .A2(n821bar), .ZN(n823bar);
  OR2_X1 U143 ( .A1(n820), .A2(n819), .ZN(n821) );
  AND2_X1 U143bar ( .A1(n820bar), .A2(n819bar), .ZN(n821bar);
  OR2_X1 U144 ( .A1(n964), .A2(n818), .ZN(n822) );
  AND2_X1 U144bar ( .A1(n964bar), .A2(n818bar), .ZN(n822bar);
  OR2_X1 U145 ( .A1(in[118]), .A2(n817), .ZN(n818) );
  AND2_X1 U145bar ( .A1(inbar[118]), .A2(n817bar), .ZN(n818bar);
  OR2_X1 U146 ( .A1(n816), .A2(n815), .ZN(n964) );
  AND2_X1 U146bar ( .A1(n816bar), .A2(n815bar), .ZN(n964bar);
  OR2_X1 U147 ( .A1(n814), .A2(n813), .ZN(n815) );
  AND2_X1 U147bar ( .A1(n814bar), .A2(n813bar), .ZN(n815bar);
  OR2_X1 U148 ( .A1(n812), .A2(n811), .ZN(n813) );
  AND2_X1 U148bar ( .A1(n812bar), .A2(n811bar), .ZN(n813bar);
  OR2_X1 U149 ( .A1(in[122]), .A2(in[111]), .ZN(n811) );
  AND2_X1 U149bar ( .A1(inbar[122]), .A2(inbar[111]), .ZN(n811bar);
  OR2_X1 U150 ( .A1(in[154]), .A2(in[151]), .ZN(n812) );
  AND2_X1 U150bar ( .A1(inbar[154]), .A2(inbar[151]), .ZN(n812bar);
  OR2_X1 U151 ( .A1(n810), .A2(n809), .ZN(n814) );
  AND2_X1 U151bar ( .A1(n810bar), .A2(n809bar), .ZN(n814bar);
  OR2_X1 U152 ( .A1(in[187]), .A2(in[177]), .ZN(n809) );
  AND2_X1 U152bar ( .A1(inbar[187]), .A2(inbar[177]), .ZN(n809bar);
  OR2_X1 U153 ( .A1(in[200]), .A2(in[192]), .ZN(n810) );
  AND2_X1 U153bar ( .A1(inbar[200]), .A2(inbar[192]), .ZN(n810bar);
  OR2_X1 U154 ( .A1(n808), .A2(n807), .ZN(n816) );
  AND2_X1 U154bar ( .A1(n808bar), .A2(n807bar), .ZN(n816bar);
  OR2_X1 U155 ( .A1(n806), .A2(n805), .ZN(n807) );
  AND2_X1 U155bar ( .A1(n806bar), .A2(n805bar), .ZN(n807bar);
  OR2_X1 U156 ( .A1(in[225]), .A2(in[207]), .ZN(n805) );
  AND2_X1 U156bar ( .A1(inbar[225]), .A2(inbar[207]), .ZN(n805bar);
  OR2_X1 U157 ( .A1(in[98]), .A2(in[226]), .ZN(n806) );
  AND2_X1 U157bar ( .A1(inbar[98]), .A2(inbar[226]), .ZN(n806bar);
  OR2_X1 U158 ( .A1(n804), .A2(n803), .ZN(n808) );
  AND2_X1 U158bar ( .A1(n804bar), .A2(n803bar), .ZN(n808bar);
  OR2_X1 U159 ( .A1(in_20), .A2(in_16), .ZN(n803) );
  AND2_X1 U159bar ( .A1(in_20bar), .A2(in_16bar), .ZN(n803bar);
  OR2_X1 U160 ( .A1(in_55), .A2(in_45), .ZN(n804) );
  AND2_X1 U160bar ( .A1(in_55bar), .A2(in_45bar), .ZN(n804bar);
  OR2_X1 U161 ( .A1(n802), .A2(n801), .ZN(n824) );
  AND2_X1 U161bar ( .A1(n802bar), .A2(n801bar), .ZN(n824bar);
  OR2_X1 U162 ( .A1(in[162]), .A2(in[149]), .ZN(n801) );
  AND2_X1 U162bar ( .A1(inbar[162]), .A2(inbar[149]), .ZN(n801bar);
  OR2_X1 U163 ( .A1(in[163]), .A2(n800), .ZN(n802) );
  AND2_X1 U163bar ( .A1(inbar[163]), .A2(n800bar), .ZN(n802bar);
  OR2_X1 U164 ( .A1(in[191]), .A2(in[189]), .ZN(n800) );
  AND2_X1 U164bar ( .A1(inbar[191]), .A2(inbar[189]), .ZN(n800bar);
  OR2_X1 U165 ( .A1(n799), .A2(n798), .ZN(n826) );
  AND2_X1 U165bar ( .A1(n799bar), .A2(n798bar), .ZN(n826bar);
  OR2_X1 U166 ( .A1(n797), .A2(n796), .ZN(n798) );
  AND2_X1 U166bar ( .A1(n797bar), .A2(n796bar), .ZN(n798bar);
  OR2_X1 U167 ( .A1(in[212]), .A2(in[193]), .ZN(n796) );
  AND2_X1 U167bar ( .A1(inbar[212]), .A2(inbar[193]), .ZN(n796bar);
  OR2_X1 U168 ( .A1(in[238]), .A2(n795), .ZN(n797) );
  AND2_X1 U168bar ( .A1(inbar[238]), .A2(n795bar), .ZN(n797bar);
  OR2_X1 U169 ( .A1(in[88]), .A2(in[247]), .ZN(n795) );
  AND2_X1 U169bar ( .A1(inbar[88]), .A2(inbar[247]), .ZN(n795bar);
  OR2_X1 U170 ( .A1(n794), .A2(n793), .ZN(n799) );
  AND2_X1 U170bar ( .A1(n794bar), .A2(n793bar), .ZN(n799bar);
  OR2_X1 U171 ( .A1(in[94]), .A2(in[92]), .ZN(n793) );
  AND2_X1 U171bar ( .A1(inbar[94]), .A2(inbar[92]), .ZN(n793bar);
  OR2_X1 U172 ( .A1(in_52), .A2(n792), .ZN(n794) );
  AND2_X1 U172bar ( .A1(in_52bar), .A2(n792bar), .ZN(n794bar);
  OR2_X1 U173 ( .A1(in_70), .A2(in_67), .ZN(n792) );
  AND2_X1 U173bar ( .A1(in_70bar), .A2(in_67bar), .ZN(n792bar);
  OR2_X1 U174 ( .A1(n791), .A2(n790), .ZN(out[2]) );
  AND2_X1 U174bar ( .A1(n791bar), .A2(n790bar), .ZN(outbar[2]);
  OR2_X1 U175 ( .A1(n789), .A2(n788), .ZN(n790) );
  AND2_X1 U175bar ( .A1(n789bar), .A2(n788bar), .ZN(n790bar);
  OR2_X1 U176 ( .A1(n787), .A2(n786), .ZN(n788) );
  AND2_X1 U176bar ( .A1(n787bar), .A2(n786bar), .ZN(n788bar);
  OR2_X1 U177 ( .A1(n819), .A2(n785), .ZN(n786) );
  AND2_X1 U177bar ( .A1(n819bar), .A2(n785bar), .ZN(n786bar);
  OR2_X1 U178 ( .A1(n784), .A2(n783), .ZN(n819) );
  AND2_X1 U178bar ( .A1(n784bar), .A2(n783bar), .ZN(n819bar);
  OR2_X1 U179 ( .A1(n782), .A2(n781), .ZN(n783) );
  AND2_X1 U179bar ( .A1(n782bar), .A2(n781bar), .ZN(n783bar);
  OR2_X1 U180 ( .A1(n780), .A2(n779), .ZN(n781) );
  AND2_X1 U180bar ( .A1(n780bar), .A2(n779bar), .ZN(n781bar);
  OR2_X1 U181 ( .A1(n962), .A2(n778), .ZN(n779) );
  AND2_X1 U181bar ( .A1(n962bar), .A2(n778bar), .ZN(n779bar);
  OR2_X1 U182 ( .A1(n777), .A2(n776), .ZN(n962) );
  AND2_X1 U182bar ( .A1(n777bar), .A2(n776bar), .ZN(n962bar);
  OR2_X1 U183 ( .A1(n775), .A2(n774), .ZN(n776) );
  AND2_X1 U183bar ( .A1(n775bar), .A2(n774bar), .ZN(n776bar);
  OR2_X1 U184 ( .A1(n773), .A2(n772), .ZN(n774) );
  AND2_X1 U184bar ( .A1(n773bar), .A2(n772bar), .ZN(n774bar);
  OR2_X1 U185 ( .A1(in[131]), .A2(in[120]), .ZN(n772) );
  AND2_X1 U185bar ( .A1(inbar[131]), .A2(inbar[120]), .ZN(n772bar);
  OR2_X1 U186 ( .A1(in[153]), .A2(in[147]), .ZN(n773) );
  AND2_X1 U186bar ( .A1(inbar[153]), .A2(inbar[147]), .ZN(n773bar);
  OR2_X1 U187 ( .A1(n771), .A2(n770), .ZN(n775) );
  AND2_X1 U187bar ( .A1(n771bar), .A2(n770bar), .ZN(n775bar);
  OR2_X1 U188 ( .A1(in[170]), .A2(in[156]), .ZN(n770) );
  AND2_X1 U188bar ( .A1(inbar[170]), .A2(inbar[156]), .ZN(n770bar);
  OR2_X1 U189 ( .A1(in[223]), .A2(in[190]), .ZN(n771) );
  AND2_X1 U189bar ( .A1(inbar[223]), .A2(inbar[190]), .ZN(n771bar);
  OR2_X1 U190 ( .A1(n769), .A2(n768), .ZN(n777) );
  AND2_X1 U190bar ( .A1(n769bar), .A2(n768bar), .ZN(n777bar);
  OR2_X1 U191 ( .A1(n767), .A2(n766), .ZN(n768) );
  AND2_X1 U191bar ( .A1(n767bar), .A2(n766bar), .ZN(n768bar);
  OR2_X1 U192 ( .A1(in[236]), .A2(in[230]), .ZN(n766) );
  AND2_X1 U192bar ( .A1(inbar[236]), .A2(inbar[230]), .ZN(n766bar);
  OR2_X1 U193 ( .A1(in[85]), .A2(in[240]), .ZN(n767) );
  AND2_X1 U193bar ( .A1(inbar[85]), .A2(inbar[240]), .ZN(n767bar);
  OR2_X1 U194 ( .A1(n765), .A2(n764), .ZN(n769) );
  AND2_X1 U194bar ( .A1(n765bar), .A2(n764bar), .ZN(n769bar);
  OR2_X1 U195 ( .A1(in_12), .A2(in[90]), .ZN(n764) );
  AND2_X1 U195bar ( .A1(in_12bar), .A2(inbar[90]), .ZN(n764bar);
  OR2_X1 U196 ( .A1(in_39), .A2(in_28), .ZN(n765) );
  AND2_X1 U196bar ( .A1(in_39bar), .A2(in_28bar), .ZN(n765bar);
  OR2_X1 U197 ( .A1(in[109]), .A2(n763), .ZN(n780) );
  AND2_X1 U197bar ( .A1(inbar[109]), .A2(n763bar), .ZN(n780bar);
  OR2_X1 U198 ( .A1(n762), .A2(n761), .ZN(n782) );
  AND2_X1 U198bar ( .A1(n762bar), .A2(n761bar), .ZN(n782bar);
  OR2_X1 U199 ( .A1(in[138]), .A2(in[129]), .ZN(n761) );
  AND2_X1 U199bar ( .A1(inbar[138]), .A2(inbar[129]), .ZN(n761bar);
  OR2_X1 U200 ( .A1(in[157]), .A2(n760), .ZN(n762) );
  AND2_X1 U200bar ( .A1(inbar[157]), .A2(n760bar), .ZN(n762bar);
  OR2_X1 U201 ( .A1(in[182]), .A2(in[167]), .ZN(n760) );
  AND2_X1 U201bar ( .A1(inbar[182]), .A2(inbar[167]), .ZN(n760bar);
  OR2_X1 U202 ( .A1(n759), .A2(n758), .ZN(n784) );
  AND2_X1 U202bar ( .A1(n759bar), .A2(n758bar), .ZN(n784bar);
  OR2_X1 U203 ( .A1(n757), .A2(n756), .ZN(n758) );
  AND2_X1 U203bar ( .A1(n757bar), .A2(n756bar), .ZN(n758bar);
  OR2_X1 U204 ( .A1(in[195]), .A2(in[184]), .ZN(n756) );
  AND2_X1 U204bar ( .A1(inbar[195]), .A2(inbar[184]), .ZN(n756bar);
  OR2_X1 U205 ( .A1(in[196]), .A2(n755), .ZN(n757) );
  AND2_X1 U205bar ( .A1(inbar[196]), .A2(n755bar), .ZN(n757bar);
  OR2_X1 U206 ( .A1(in[215]), .A2(in[209]), .ZN(n755) );
  AND2_X1 U206bar ( .A1(inbar[215]), .A2(inbar[209]), .ZN(n755bar);
  OR2_X1 U207 ( .A1(n754), .A2(n753), .ZN(n759) );
  AND2_X1 U207bar ( .A1(n754bar), .A2(n753bar), .ZN(n759bar);
  OR2_X1 U208 ( .A1(in[93]), .A2(in[233]), .ZN(n753) );
  AND2_X1 U208bar ( .A1(inbar[93]), .A2(inbar[233]), .ZN(n753bar);
  OR2_X1 U209 ( .A1(in_1), .A2(n752), .ZN(n754) );
  AND2_X1 U209bar ( .A1(in_1bar), .A2(n752bar), .ZN(n754bar);
  OR2_X1 U210 ( .A1(in_69), .A2(in_66), .ZN(n752) );
  AND2_X1 U210bar ( .A1(in_69bar), .A2(in_66bar), .ZN(n752bar);
  OR2_X1 U211 ( .A1(n966), .A2(n751), .ZN(n787) );
  AND2_X1 U211bar ( .A1(n966bar), .A2(n751bar), .ZN(n787bar);
  OR2_X1 U212 ( .A1(in[134]), .A2(n750), .ZN(n751) );
  AND2_X1 U212bar ( .A1(inbar[134]), .A2(n750bar), .ZN(n751bar);
  OR2_X1 U213 ( .A1(n749), .A2(n748), .ZN(n966) );
  AND2_X1 U213bar ( .A1(n749bar), .A2(n748bar), .ZN(n966bar);
  OR2_X1 U214 ( .A1(n747), .A2(n746), .ZN(n748) );
  AND2_X1 U214bar ( .A1(n747bar), .A2(n746bar), .ZN(n748bar);
  OR2_X1 U215 ( .A1(n745), .A2(n744), .ZN(n746) );
  AND2_X1 U215bar ( .A1(n745bar), .A2(n744bar), .ZN(n746bar);
  OR2_X1 U216 ( .A1(in[136]), .A2(in[121]), .ZN(n744) );
  AND2_X1 U216bar ( .A1(inbar[136]), .A2(inbar[121]), .ZN(n744bar);
  OR2_X1 U217 ( .A1(in[186]), .A2(in[174]), .ZN(n745) );
  AND2_X1 U217bar ( .A1(inbar[186]), .A2(inbar[174]), .ZN(n745bar);
  OR2_X1 U218 ( .A1(n743), .A2(n742), .ZN(n747) );
  AND2_X1 U218bar ( .A1(n743bar), .A2(n742bar), .ZN(n747bar);
  OR2_X1 U219 ( .A1(in[198]), .A2(in[197]), .ZN(n742) );
  AND2_X1 U219bar ( .A1(inbar[198]), .A2(inbar[197]), .ZN(n742bar);
  OR2_X1 U220 ( .A1(in[214]), .A2(in[199]), .ZN(n743) );
  AND2_X1 U220bar ( .A1(inbar[214]), .A2(inbar[199]), .ZN(n743bar);
  OR2_X1 U221 ( .A1(n741), .A2(n740), .ZN(n749) );
  AND2_X1 U221bar ( .A1(n741bar), .A2(n740bar), .ZN(n749bar);
  OR2_X1 U222 ( .A1(n739), .A2(n738), .ZN(n740) );
  AND2_X1 U222bar ( .A1(n739bar), .A2(n738bar), .ZN(n740bar);
  OR2_X1 U223 ( .A1(in[231]), .A2(in[220]), .ZN(n738) );
  AND2_X1 U223bar ( .A1(inbar[231]), .A2(inbar[220]), .ZN(n738bar);
  OR2_X1 U224 ( .A1(in_25), .A2(in[245]), .ZN(n739) );
  AND2_X1 U224bar ( .A1(in_25bar), .A2(inbar[245]), .ZN(n739bar);
  OR2_X1 U225 ( .A1(n737), .A2(n736), .ZN(n741) );
  AND2_X1 U225bar ( .A1(n737bar), .A2(n736bar), .ZN(n741bar);
  OR2_X1 U226 ( .A1(in_53), .A2(in_29), .ZN(n736) );
  AND2_X1 U226bar ( .A1(in_53bar), .A2(in_29bar), .ZN(n736bar);
  OR2_X1 U227 ( .A1(in_79), .A2(in_74), .ZN(n737) );
  AND2_X1 U227bar ( .A1(in_79bar), .A2(in_74bar), .ZN(n737bar);
  OR2_X1 U228 ( .A1(n735), .A2(n734), .ZN(n789) );
  AND2_X1 U228bar ( .A1(n735bar), .A2(n734bar), .ZN(n789bar);
  OR2_X1 U229 ( .A1(in[152]), .A2(in[140]), .ZN(n734) );
  AND2_X1 U229bar ( .A1(inbar[152]), .A2(inbar[140]), .ZN(n734bar);
  OR2_X1 U230 ( .A1(in[155]), .A2(n733), .ZN(n735) );
  AND2_X1 U230bar ( .A1(inbar[155]), .A2(n733bar), .ZN(n735bar);
  OR2_X1 U231 ( .A1(in[166]), .A2(in[165]), .ZN(n733) );
  AND2_X1 U231bar ( .A1(inbar[166]), .A2(inbar[165]), .ZN(n733bar);
  OR2_X1 U232 ( .A1(n732), .A2(n731), .ZN(n791) );
  AND2_X1 U232bar ( .A1(n732bar), .A2(n731bar), .ZN(n791bar);
  OR2_X1 U233 ( .A1(n730), .A2(n729), .ZN(n731) );
  AND2_X1 U233bar ( .A1(n730bar), .A2(n729bar), .ZN(n731bar);
  OR2_X1 U234 ( .A1(in[202]), .A2(in[185]), .ZN(n729) );
  AND2_X1 U234bar ( .A1(inbar[202]), .A2(inbar[185]), .ZN(n729bar);
  OR2_X1 U235 ( .A1(in[211]), .A2(n728), .ZN(n730) );
  AND2_X1 U235bar ( .A1(inbar[211]), .A2(n728bar), .ZN(n730bar);
  OR2_X1 U236 ( .A1(in[255]), .A2(in[253]), .ZN(n728) );
  AND2_X1 U236bar ( .A1(inbar[255]), .A2(inbar[253]), .ZN(n728bar);
  OR2_X1 U237 ( .A1(n727), .A2(n726), .ZN(n732) );
  AND2_X1 U237bar ( .A1(n727bar), .A2(n726bar), .ZN(n732bar);
  OR2_X1 U238 ( .A1(in_35), .A2(in_15), .ZN(n726) );
  AND2_X1 U238bar ( .A1(in_35bar), .A2(in_15bar), .ZN(n726bar);
  OR2_X1 U239 ( .A1(in_36), .A2(n725), .ZN(n727) );
  AND2_X1 U239bar ( .A1(in_36bar), .A2(n725bar), .ZN(n727bar);
  OR2_X1 U240 ( .A1(in_48), .A2(in_40), .ZN(n725) );
  AND2_X1 U240bar ( .A1(in_48bar), .A2(in_40bar), .ZN(n725bar);
  OR2_X1 U241 ( .A1(n724), .A2(n723), .ZN(out[1]) );
  AND2_X1 U241bar ( .A1(n724bar), .A2(n723bar), .ZN(outbar[1]);
  OR2_X1 U242 ( .A1(n722), .A2(n721), .ZN(n723) );
  AND2_X1 U242bar ( .A1(n722bar), .A2(n721bar), .ZN(n723bar);
  OR2_X1 U243 ( .A1(n720), .A2(n719), .ZN(n721) );
  AND2_X1 U243bar ( .A1(n720bar), .A2(n719bar), .ZN(n721bar);
  OR2_X1 U244 ( .A1(n921), .A2(n887), .ZN(n719) );
  AND2_X1 U244bar ( .A1(n921bar), .A2(n887bar), .ZN(n719bar);
  OR2_X1 U245 ( .A1(n718), .A2(n717), .ZN(n887) );
  AND2_X1 U245bar ( .A1(n718bar), .A2(n717bar), .ZN(n887bar);
  OR2_X1 U246 ( .A1(n716), .A2(n715), .ZN(n717) );
  AND2_X1 U246bar ( .A1(n716bar), .A2(n715bar), .ZN(n717bar);
  OR2_X1 U247 ( .A1(n714), .A2(n713), .ZN(n715) );
  AND2_X1 U247bar ( .A1(n714bar), .A2(n713bar), .ZN(n715bar);
  OR2_X1 U248 ( .A1(in[116]), .A2(in[110]), .ZN(n713) );
  AND2_X1 U248bar ( .A1(inbar[116]), .A2(inbar[110]), .ZN(n713bar);
  OR2_X1 U249 ( .A1(in[133]), .A2(in[130]), .ZN(n714) );
  AND2_X1 U249bar ( .A1(inbar[133]), .A2(inbar[130]), .ZN(n714bar);
  OR2_X1 U250 ( .A1(n712), .A2(n711), .ZN(n716) );
  AND2_X1 U250bar ( .A1(n712bar), .A2(n711bar), .ZN(n716bar);
  OR2_X1 U251 ( .A1(in[203]), .A2(in[135]), .ZN(n711) );
  AND2_X1 U251bar ( .A1(inbar[203]), .A2(inbar[135]), .ZN(n711bar);
  OR2_X1 U252 ( .A1(in[232]), .A2(in[223]), .ZN(n712) );
  AND2_X1 U252bar ( .A1(inbar[232]), .A2(inbar[223]), .ZN(n712bar);
  OR2_X1 U253 ( .A1(n710), .A2(n709), .ZN(n718) );
  AND2_X1 U253bar ( .A1(n710bar), .A2(n709bar), .ZN(n718bar);
  OR2_X1 U254 ( .A1(n708), .A2(n707), .ZN(n709) );
  AND2_X1 U254bar ( .A1(n708bar), .A2(n707bar), .ZN(n709bar);
  OR2_X1 U255 ( .A1(in[255]), .A2(in[233]), .ZN(n707) );
  AND2_X1 U255bar ( .A1(inbar[255]), .A2(inbar[233]), .ZN(n707bar);
  OR2_X1 U256 ( .A1(in_53), .A2(in_34), .ZN(n708) );
  AND2_X1 U256bar ( .A1(in_53bar), .A2(in_34bar), .ZN(n708bar);
  OR2_X1 U257 ( .A1(n706), .A2(n705), .ZN(n710) );
  AND2_X1 U257bar ( .A1(n706bar), .A2(n705bar), .ZN(n710bar);
  OR2_X1 U258 ( .A1(in_57), .A2(in_55), .ZN(n705) );
  AND2_X1 U258bar ( .A1(in_57bar), .A2(in_55bar), .ZN(n705bar);
  OR2_X1 U259 ( .A1(in_68), .A2(in_67), .ZN(n706) );
  AND2_X1 U259bar ( .A1(in_68bar), .A2(in_67bar), .ZN(n706bar);
  OR2_X1 U260 ( .A1(n704), .A2(n703), .ZN(n921) );
  AND2_X1 U260bar ( .A1(n704bar), .A2(n703bar), .ZN(n921bar);
  OR2_X1 U261 ( .A1(n702), .A2(n701), .ZN(n703) );
  AND2_X1 U261bar ( .A1(n702bar), .A2(n701bar), .ZN(n703bar);
  OR2_X1 U262 ( .A1(n700), .A2(n699), .ZN(n701) );
  AND2_X1 U262bar ( .A1(n700bar), .A2(n699bar), .ZN(n701bar);
  OR2_X1 U263 ( .A1(n944), .A2(n872), .ZN(n699) );
  AND2_X1 U263bar ( .A1(n944bar), .A2(n872bar), .ZN(n699bar);
  OR2_X1 U264 ( .A1(n698), .A2(n697), .ZN(n872) );
  AND2_X1 U264bar ( .A1(n698bar), .A2(n697bar), .ZN(n872bar);
  OR2_X1 U265 ( .A1(n696), .A2(n695), .ZN(n697) );
  AND2_X1 U265bar ( .A1(n696bar), .A2(n695bar), .ZN(n697bar);
  OR2_X1 U266 ( .A1(n694), .A2(n693), .ZN(n695) );
  AND2_X1 U266bar ( .A1(n694bar), .A2(n693bar), .ZN(n695bar);
  OR2_X1 U267 ( .A1(in[121]), .A2(in[102]), .ZN(n693) );
  AND2_X1 U267bar ( .A1(inbar[121]), .A2(inbar[102]), .ZN(n693bar);
  OR2_X1 U268 ( .A1(in[162]), .A2(in[161]), .ZN(n694) );
  AND2_X1 U268bar ( .A1(inbar[162]), .A2(inbar[161]), .ZN(n694bar);
  OR2_X1 U269 ( .A1(n692), .A2(n691), .ZN(n696) );
  AND2_X1 U269bar ( .A1(n692bar), .A2(n691bar), .ZN(n696bar);
  OR2_X1 U270 ( .A1(in[192]), .A2(in[178]), .ZN(n691) );
  AND2_X1 U270bar ( .A1(inbar[192]), .A2(inbar[178]), .ZN(n691bar);
  OR2_X1 U271 ( .A1(in[244]), .A2(in[209]), .ZN(n692) );
  AND2_X1 U271bar ( .A1(inbar[244]), .A2(inbar[209]), .ZN(n692bar);
  OR2_X1 U272 ( .A1(n690), .A2(n689), .ZN(n698) );
  AND2_X1 U272bar ( .A1(n690bar), .A2(n689bar), .ZN(n698bar);
  OR2_X1 U273 ( .A1(n688), .A2(n687), .ZN(n689) );
  AND2_X1 U273bar ( .A1(n688bar), .A2(n687bar), .ZN(n689bar);
  OR2_X1 U274 ( .A1(in[90]), .A2(in[254]), .ZN(n687) );
  AND2_X1 U274bar ( .A1(inbar[90]), .A2(inbar[254]), .ZN(n687bar);
  OR2_X1 U275 ( .A1(in_36), .A2(in_32), .ZN(n688) );
  AND2_X1 U275bar ( .A1(in_36bar), .A2(in_32bar), .ZN(n688bar);
  OR2_X1 U276 ( .A1(n686), .A2(n685), .ZN(n690) );
  AND2_X1 U276bar ( .A1(n686bar), .A2(n685bar), .ZN(n690bar);
  OR2_X1 U277 ( .A1(in_62), .A2(in_37), .ZN(n685) );
  AND2_X1 U277bar ( .A1(in_62bar), .A2(in_37bar), .ZN(n685bar);
  OR2_X1 U278 ( .A1(in_75), .A2(in_73), .ZN(n686) );
  AND2_X1 U278bar ( .A1(in_75bar), .A2(in_73bar), .ZN(n686bar);
  OR2_X1 U279 ( .A1(n684), .A2(n683), .ZN(n944) );
  AND2_X1 U279bar ( .A1(n684bar), .A2(n683bar), .ZN(n944bar);
  OR2_X1 U280 ( .A1(n682), .A2(n681), .ZN(n683) );
  AND2_X1 U280bar ( .A1(n682bar), .A2(n681bar), .ZN(n683bar);
  OR2_X1 U281 ( .A1(n680), .A2(n679), .ZN(n681) );
  AND2_X1 U281bar ( .A1(n680bar), .A2(n679bar), .ZN(n681bar);
  OR2_X1 U282 ( .A1(in[171]), .A2(in[153]), .ZN(n679) );
  AND2_X1 U282bar ( .A1(inbar[171]), .A2(inbar[153]), .ZN(n679bar);
  OR2_X1 U283 ( .A1(in[187]), .A2(in[176]), .ZN(n680) );
  AND2_X1 U283bar ( .A1(inbar[187]), .A2(inbar[176]), .ZN(n680bar);
  OR2_X1 U284 ( .A1(n678), .A2(n677), .ZN(n682) );
  AND2_X1 U284bar ( .A1(n678bar), .A2(n677bar), .ZN(n682bar);
  OR2_X1 U285 ( .A1(in[245]), .A2(in[211]), .ZN(n677) );
  AND2_X1 U285bar ( .A1(inbar[245]), .A2(inbar[211]), .ZN(n677bar);
  OR2_X1 U286 ( .A1(in[97]), .A2(in[88]), .ZN(n678) );
  AND2_X1 U286bar ( .A1(inbar[97]), .A2(inbar[88]), .ZN(n678bar);
  OR2_X1 U287 ( .A1(n676), .A2(n675), .ZN(n684) );
  AND2_X1 U287bar ( .A1(n676bar), .A2(n675bar), .ZN(n684bar);
  OR2_X1 U288 ( .A1(n674), .A2(n673), .ZN(n675) );
  AND2_X1 U288bar ( .A1(n674bar), .A2(n673bar), .ZN(n675bar);
  OR2_X1 U289 ( .A1(in_10), .A2(in_0), .ZN(n673) );
  AND2_X1 U289bar ( .A1(in_10bar), .A2(in_0bar), .ZN(n673bar);
  OR2_X1 U290 ( .A1(in_59), .A2(in_5), .ZN(n674) );
  AND2_X1 U290bar ( .A1(in_59bar), .A2(in_5bar), .ZN(n674bar);
  OR2_X1 U291 ( .A1(n672), .A2(n671), .ZN(n676) );
  AND2_X1 U291bar ( .A1(n672bar), .A2(n671bar), .ZN(n676bar);
  OR2_X1 U292 ( .A1(in_60), .A2(in_6), .ZN(n671) );
  AND2_X1 U292bar ( .A1(in_60bar), .A2(in_6bar), .ZN(n671bar);
  OR2_X1 U293 ( .A1(in_77), .A2(in_69), .ZN(n672) );
  AND2_X1 U293bar ( .A1(in_77bar), .A2(in_69bar), .ZN(n672bar);
  OR2_X1 U294 ( .A1(in[113]), .A2(n864), .ZN(n700) );
  AND2_X1 U294bar ( .A1(inbar[113]), .A2(n864bar), .ZN(n700bar);
  OR2_X1 U295 ( .A1(n670), .A2(n669), .ZN(n864) );
  AND2_X1 U295bar ( .A1(n670bar), .A2(n669bar), .ZN(n864bar);
  OR2_X1 U296 ( .A1(n668), .A2(n667), .ZN(n669) );
  AND2_X1 U296bar ( .A1(n668bar), .A2(n667bar), .ZN(n669bar);
  OR2_X1 U297 ( .A1(n666), .A2(n665), .ZN(n667) );
  AND2_X1 U297bar ( .A1(n666bar), .A2(n665bar), .ZN(n667bar);
  OR2_X1 U298 ( .A1(in[125]), .A2(in[107]), .ZN(n665) );
  AND2_X1 U298bar ( .A1(inbar[125]), .A2(inbar[107]), .ZN(n665bar);
  OR2_X1 U299 ( .A1(in[138]), .A2(in[126]), .ZN(n666) );
  AND2_X1 U299bar ( .A1(inbar[138]), .A2(inbar[126]), .ZN(n666bar);
  OR2_X1 U300 ( .A1(n664), .A2(n663), .ZN(n668) );
  AND2_X1 U300bar ( .A1(n664bar), .A2(n663bar), .ZN(n668bar);
  OR2_X1 U301 ( .A1(in[189]), .A2(in[143]), .ZN(n663) );
  AND2_X1 U301bar ( .A1(inbar[189]), .A2(inbar[143]), .ZN(n663bar);
  OR2_X1 U302 ( .A1(in[99]), .A2(in[214]), .ZN(n664) );
  AND2_X1 U302bar ( .A1(inbar[99]), .A2(inbar[214]), .ZN(n664bar);
  OR2_X1 U303 ( .A1(n662), .A2(n661), .ZN(n670) );
  AND2_X1 U303bar ( .A1(n662bar), .A2(n661bar), .ZN(n670bar);
  OR2_X1 U304 ( .A1(n660), .A2(n659), .ZN(n661) );
  AND2_X1 U304bar ( .A1(n660bar), .A2(n659bar), .ZN(n661bar);
  OR2_X1 U305 ( .A1(in_15), .A2(in_12), .ZN(n659) );
  AND2_X1 U305bar ( .A1(in_15bar), .A2(in_12bar), .ZN(n659bar);
  OR2_X1 U306 ( .A1(in_20), .A2(in_2), .ZN(n660) );
  AND2_X1 U306bar ( .A1(in_20bar), .A2(in_2bar), .ZN(n660bar);
  OR2_X1 U307 ( .A1(n658), .A2(n657), .ZN(n662) );
  AND2_X1 U307bar ( .A1(n658bar), .A2(n657bar), .ZN(n662bar);
  OR2_X1 U308 ( .A1(in_30), .A2(in_3), .ZN(n657) );
  AND2_X1 U308bar ( .A1(in_30bar), .A2(in_3bar), .ZN(n657bar);
  OR2_X1 U309 ( .A1(in_4), .A2(in_38), .ZN(n658) );
  AND2_X1 U309bar ( .A1(in_4bar), .A2(in_38bar), .ZN(n658bar);
  OR2_X1 U310 ( .A1(n656), .A2(n655), .ZN(n702) );
  AND2_X1 U310bar ( .A1(n656bar), .A2(n655bar), .ZN(n702bar);
  OR2_X1 U311 ( .A1(in[148]), .A2(in[137]), .ZN(n655) );
  AND2_X1 U311bar ( .A1(inbar[148]), .A2(inbar[137]), .ZN(n655bar);
  OR2_X1 U312 ( .A1(in[149]), .A2(n654), .ZN(n656) );
  AND2_X1 U312bar ( .A1(inbar[149]), .A2(n654bar), .ZN(n656bar);
  OR2_X1 U313 ( .A1(in[195]), .A2(in[190]), .ZN(n654) );
  AND2_X1 U313bar ( .A1(inbar[195]), .A2(inbar[190]), .ZN(n654bar);
  OR2_X1 U314 ( .A1(n653), .A2(n652), .ZN(n704) );
  AND2_X1 U314bar ( .A1(n653bar), .A2(n652bar), .ZN(n704bar);
  OR2_X1 U315 ( .A1(n651), .A2(n650), .ZN(n652) );
  AND2_X1 U315bar ( .A1(n651bar), .A2(n650bar), .ZN(n652bar);
  OR2_X1 U316 ( .A1(in[98]), .A2(in[197]), .ZN(n650) );
  AND2_X1 U316bar ( .A1(inbar[98]), .A2(inbar[197]), .ZN(n650bar);
  OR2_X1 U317 ( .A1(in_11), .A2(n649), .ZN(n651) );
  AND2_X1 U317bar ( .A1(in_11bar), .A2(n649bar), .ZN(n651bar);
  OR2_X1 U318 ( .A1(in_26), .A2(in_14), .ZN(n649) );
  AND2_X1 U318bar ( .A1(in_26bar), .A2(in_14bar), .ZN(n649bar);
  OR2_X1 U319 ( .A1(n648), .A2(n647), .ZN(n653) );
  AND2_X1 U319bar ( .A1(n648bar), .A2(n647bar), .ZN(n653bar);
  OR2_X1 U320 ( .A1(in_35), .A2(in_27), .ZN(n647) );
  AND2_X1 U320bar ( .A1(in_35bar), .A2(in_27bar), .ZN(n647bar);
  OR2_X1 U321 ( .A1(in_50), .A2(n646), .ZN(n648) );
  AND2_X1 U321bar ( .A1(in_50bar), .A2(n646bar), .ZN(n648bar);
  OR2_X1 U322 ( .A1(in_78), .A2(in_61), .ZN(n646) );
  AND2_X1 U322bar ( .A1(in_78bar), .A2(in_61bar), .ZN(n646bar);
  OR2_X1 U323 ( .A1(n942), .A2(n645), .ZN(n720) );
  AND2_X1 U323bar ( .A1(n942bar), .A2(n645bar), .ZN(n720bar);
  OR2_X1 U324 ( .A1(in[106]), .A2(n863), .ZN(n645) );
  AND2_X1 U324bar ( .A1(inbar[106]), .A2(n863bar), .ZN(n645bar);
  OR2_X1 U325 ( .A1(n644), .A2(n643), .ZN(n863) );
  AND2_X1 U325bar ( .A1(n644bar), .A2(n643bar), .ZN(n863bar);
  OR2_X1 U326 ( .A1(n642), .A2(n641), .ZN(n643) );
  AND2_X1 U326bar ( .A1(n642bar), .A2(n641bar), .ZN(n643bar);
  OR2_X1 U327 ( .A1(n640), .A2(n639), .ZN(n641) );
  AND2_X1 U327bar ( .A1(n640bar), .A2(n639bar), .ZN(n641bar);
  OR2_X1 U328 ( .A1(in[127]), .A2(in[122]), .ZN(n639) );
  AND2_X1 U328bar ( .A1(inbar[127]), .A2(inbar[122]), .ZN(n639bar);
  OR2_X1 U329 ( .A1(in[156]), .A2(in[132]), .ZN(n640) );
  AND2_X1 U329bar ( .A1(inbar[156]), .A2(inbar[132]), .ZN(n640bar);
  OR2_X1 U330 ( .A1(n638), .A2(n637), .ZN(n642) );
  AND2_X1 U330bar ( .A1(n638bar), .A2(n637bar), .ZN(n642bar);
  OR2_X1 U331 ( .A1(in[159]), .A2(in[157]), .ZN(n637) );
  AND2_X1 U331bar ( .A1(inbar[159]), .A2(inbar[157]), .ZN(n637bar);
  OR2_X1 U332 ( .A1(in[185]), .A2(in[169]), .ZN(n638) );
  AND2_X1 U332bar ( .A1(inbar[185]), .A2(inbar[169]), .ZN(n638bar);
  OR2_X1 U333 ( .A1(n636), .A2(n635), .ZN(n644) );
  AND2_X1 U333bar ( .A1(n636bar), .A2(n635bar), .ZN(n644bar);
  OR2_X1 U334 ( .A1(n634), .A2(n633), .ZN(n635) );
  AND2_X1 U334bar ( .A1(n634bar), .A2(n633bar), .ZN(n635bar);
  OR2_X1 U335 ( .A1(in[239]), .A2(in[218]), .ZN(n633) );
  AND2_X1 U335bar ( .A1(inbar[239]), .A2(inbar[218]), .ZN(n633bar);
  OR2_X1 U336 ( .A1(in_13), .A2(in[87]), .ZN(n634) );
  AND2_X1 U336bar ( .A1(in_13bar), .A2(inbar[87]), .ZN(n634bar);
  OR2_X1 U337 ( .A1(n632), .A2(n631), .ZN(n636) );
  AND2_X1 U337bar ( .A1(n632bar), .A2(n631bar), .ZN(n636bar);
  OR2_X1 U338 ( .A1(in_72), .A2(in_70), .ZN(n631) );
  AND2_X1 U338bar ( .A1(in_72bar), .A2(in_70bar), .ZN(n631bar);
  OR2_X1 U339 ( .A1(in_80), .A2(in_74), .ZN(n632) );
  AND2_X1 U339bar ( .A1(in_80bar), .A2(in_74bar), .ZN(n632bar);
  OR2_X1 U340 ( .A1(n630), .A2(n629), .ZN(n942) );
  AND2_X1 U340bar ( .A1(n630bar), .A2(n629bar), .ZN(n942bar);
  OR2_X1 U341 ( .A1(n628), .A2(n627), .ZN(n629) );
  AND2_X1 U341bar ( .A1(n628bar), .A2(n627bar), .ZN(n629bar);
  OR2_X1 U342 ( .A1(n626), .A2(n625), .ZN(n627) );
  AND2_X1 U342bar ( .A1(n626bar), .A2(n625bar), .ZN(n627bar);
  OR2_X1 U343 ( .A1(in[146]), .A2(in[100]), .ZN(n625) );
  AND2_X1 U343bar ( .A1(inbar[146]), .A2(inbar[100]), .ZN(n625bar);
  OR2_X1 U344 ( .A1(in[168]), .A2(in[152]), .ZN(n626) );
  AND2_X1 U344bar ( .A1(inbar[168]), .A2(inbar[152]), .ZN(n626bar);
  OR2_X1 U345 ( .A1(n624), .A2(n623), .ZN(n628) );
  AND2_X1 U345bar ( .A1(n624bar), .A2(n623bar), .ZN(n628bar);
  OR2_X1 U346 ( .A1(in[199]), .A2(in[182]), .ZN(n623) );
  AND2_X1 U346bar ( .A1(inbar[199]), .A2(inbar[182]), .ZN(n623bar);
  OR2_X1 U347 ( .A1(in[236]), .A2(in[204]), .ZN(n624) );
  AND2_X1 U347bar ( .A1(inbar[236]), .A2(inbar[204]), .ZN(n624bar);
  OR2_X1 U348 ( .A1(n622), .A2(n621), .ZN(n630) );
  AND2_X1 U348bar ( .A1(n622bar), .A2(n621bar), .ZN(n630bar);
  OR2_X1 U349 ( .A1(n620), .A2(n619), .ZN(n621) );
  AND2_X1 U349bar ( .A1(n620bar), .A2(n619bar), .ZN(n621bar);
  OR2_X1 U350 ( .A1(in[89]), .A2(in[246]), .ZN(n619) );
  AND2_X1 U350bar ( .A1(inbar[89]), .A2(inbar[246]), .ZN(n619bar);
  OR2_X1 U351 ( .A1(in[95]), .A2(in[92]), .ZN(n620) );
  AND2_X1 U351bar ( .A1(inbar[95]), .A2(inbar[92]), .ZN(n620bar);
  OR2_X1 U352 ( .A1(n618), .A2(n617), .ZN(n622) );
  AND2_X1 U352bar ( .A1(n618bar), .A2(n617bar), .ZN(n622bar);
  OR2_X1 U353 ( .A1(in_22), .A2(in_16), .ZN(n617) );
  AND2_X1 U353bar ( .A1(in_22bar), .A2(in_16bar), .ZN(n617bar);
  OR2_X1 U354 ( .A1(in_51), .A2(in_49), .ZN(n618) );
  AND2_X1 U354bar ( .A1(in_51bar), .A2(in_49bar), .ZN(n618bar);
  OR2_X1 U355 ( .A1(n616), .A2(n615), .ZN(n722) );
  AND2_X1 U355bar ( .A1(n616bar), .A2(n615bar), .ZN(n722bar);
  OR2_X1 U356 ( .A1(in[158]), .A2(in[115]), .ZN(n615) );
  AND2_X1 U356bar ( .A1(inbar[158]), .A2(inbar[115]), .ZN(n615bar);
  OR2_X1 U357 ( .A1(in[163]), .A2(n614), .ZN(n616) );
  AND2_X1 U357bar ( .A1(inbar[163]), .A2(n614bar), .ZN(n616bar);
  OR2_X1 U358 ( .A1(in[206]), .A2(in[165]), .ZN(n614) );
  AND2_X1 U358bar ( .A1(inbar[206]), .A2(inbar[165]), .ZN(n614bar);
  OR2_X1 U359 ( .A1(n613), .A2(n612), .ZN(n724) );
  AND2_X1 U359bar ( .A1(n613bar), .A2(n612bar), .ZN(n724bar);
  OR2_X1 U360 ( .A1(n611), .A2(n610), .ZN(n612) );
  AND2_X1 U360bar ( .A1(n611bar), .A2(n610bar), .ZN(n612bar);
  OR2_X1 U361 ( .A1(in[213]), .A2(in[207]), .ZN(n610) );
  AND2_X1 U361bar ( .A1(inbar[213]), .A2(inbar[207]), .ZN(n610bar);
  OR2_X1 U362 ( .A1(in[215]), .A2(n609), .ZN(n611) );
  AND2_X1 U362bar ( .A1(inbar[215]), .A2(n609bar), .ZN(n611bar);
  OR2_X1 U363 ( .A1(in[230]), .A2(in[220]), .ZN(n609) );
  AND2_X1 U363bar ( .A1(inbar[230]), .A2(inbar[220]), .ZN(n609bar);
  OR2_X1 U364 ( .A1(n608), .A2(n607), .ZN(n613) );
  AND2_X1 U364bar ( .A1(n608bar), .A2(n607bar), .ZN(n613bar);
  OR2_X1 U365 ( .A1(in[251]), .A2(in[234]), .ZN(n607) );
  AND2_X1 U365bar ( .A1(inbar[251]), .A2(inbar[234]), .ZN(n607bar);
  OR2_X1 U366 ( .A1(in_17), .A2(n606), .ZN(n608) );
  AND2_X1 U366bar ( .A1(in_17bar), .A2(n606bar), .ZN(n608bar);
  OR2_X1 U367 ( .A1(in_65), .A2(in_56), .ZN(n606) );
  AND2_X1 U367bar ( .A1(in_65bar), .A2(in_56bar), .ZN(n606bar);
  OR2_X1 U368 ( .A1(n605), .A2(n604), .ZN(out[0]) );
  AND2_X1 U368bar ( .A1(n605bar), .A2(n604bar), .ZN(outbar[0]);
  OR2_X1 U369 ( .A1(n603), .A2(n602), .ZN(n604) );
  AND2_X1 U369bar ( .A1(n603bar), .A2(n602bar), .ZN(n604bar);
  OR2_X1 U370 ( .A1(n601), .A2(n600), .ZN(n602) );
  AND2_X1 U370bar ( .A1(n601bar), .A2(n600bar), .ZN(n602bar);
  OR2_X1 U371 ( .A1(n820), .A2(n785), .ZN(n600) );
  AND2_X1 U371bar ( .A1(n820bar), .A2(n785bar), .ZN(n600bar);
  OR2_X1 U372 ( .A1(n599), .A2(n598), .ZN(n785) );
  AND2_X1 U372bar ( .A1(n599bar), .A2(n598bar), .ZN(n785bar);
  OR2_X1 U373 ( .A1(n597), .A2(n596), .ZN(n598) );
  AND2_X1 U373bar ( .A1(n597bar), .A2(n596bar), .ZN(n598bar);
  OR2_X1 U374 ( .A1(n595), .A2(n594), .ZN(n596) );
  AND2_X1 U374bar ( .A1(n595bar), .A2(n594bar), .ZN(n596bar);
  OR2_X1 U375 ( .A1(in[135]), .A2(in[104]), .ZN(n594) );
  AND2_X1 U375bar ( .A1(inbar[135]), .A2(inbar[104]), .ZN(n594bar);
  OR2_X1 U376 ( .A1(in[188]), .A2(in[178]), .ZN(n595) );
  AND2_X1 U376bar ( .A1(inbar[188]), .A2(inbar[178]), .ZN(n595bar);
  OR2_X1 U377 ( .A1(n593), .A2(n592), .ZN(n597) );
  AND2_X1 U377bar ( .A1(n593bar), .A2(n592bar), .ZN(n597bar);
  OR2_X1 U378 ( .A1(in[217]), .A2(in[194]), .ZN(n592) );
  AND2_X1 U378bar ( .A1(inbar[217]), .A2(inbar[194]), .ZN(n592bar);
  OR2_X1 U379 ( .A1(in[237]), .A2(in[218]), .ZN(n593) );
  AND2_X1 U379bar ( .A1(inbar[237]), .A2(inbar[218]), .ZN(n593bar);
  OR2_X1 U380 ( .A1(n591), .A2(n590), .ZN(n599) );
  AND2_X1 U380bar ( .A1(n591bar), .A2(n590bar), .ZN(n599bar);
  OR2_X1 U381 ( .A1(n589), .A2(n588), .ZN(n590) );
  AND2_X1 U381bar ( .A1(n589bar), .A2(n588bar), .ZN(n590bar);
  OR2_X1 U382 ( .A1(in_2), .A2(in_10), .ZN(n588) );
  AND2_X1 U382bar ( .A1(in_2bar), .A2(in_10bar), .ZN(n588bar);
  OR2_X1 U383 ( .A1(in_47), .A2(in_22), .ZN(n589) );
  AND2_X1 U383bar ( .A1(in_47bar), .A2(in_22bar), .ZN(n589bar);
  OR2_X1 U384 ( .A1(n587), .A2(n586), .ZN(n591) );
  AND2_X1 U384bar ( .A1(n587bar), .A2(n586bar), .ZN(n591bar);
  OR2_X1 U385 ( .A1(in_56), .A2(in_54), .ZN(n586) );
  AND2_X1 U385bar ( .A1(in_56bar), .A2(in_54bar), .ZN(n586bar);
  OR2_X1 U386 ( .A1(in_63), .A2(in_61), .ZN(n587) );
  AND2_X1 U386bar ( .A1(in_63bar), .A2(in_61bar), .ZN(n587bar);
  OR2_X1 U387 ( .A1(n585), .A2(n584), .ZN(n820) );
  AND2_X1 U387bar ( .A1(n585bar), .A2(n584bar), .ZN(n820bar);
  OR2_X1 U388 ( .A1(n583), .A2(n582), .ZN(n584) );
  AND2_X1 U388bar ( .A1(n583bar), .A2(n582bar), .ZN(n584bar);
  OR2_X1 U389 ( .A1(n581), .A2(n580), .ZN(n582) );
  AND2_X1 U389bar ( .A1(n581bar), .A2(n580bar), .ZN(n582bar);
  OR2_X1 U390 ( .A1(in[158]), .A2(in[142]), .ZN(n580) );
  AND2_X1 U390bar ( .A1(inbar[158]), .A2(inbar[142]), .ZN(n580bar);
  OR2_X1 U391 ( .A1(in[175]), .A2(in[164]), .ZN(n581) );
  AND2_X1 U391bar ( .A1(inbar[175]), .A2(inbar[164]), .ZN(n581bar);
  OR2_X1 U392 ( .A1(n579), .A2(n578), .ZN(n583) );
  AND2_X1 U392bar ( .A1(n579bar), .A2(n578bar), .ZN(n583bar);
  OR2_X1 U393 ( .A1(in[228]), .A2(in[204]), .ZN(n578) );
  AND2_X1 U393bar ( .A1(inbar[228]), .A2(inbar[204]), .ZN(n578bar);
  OR2_X1 U394 ( .A1(in[91]), .A2(in[87]), .ZN(n579) );
  AND2_X1 U394bar ( .A1(inbar[91]), .A2(inbar[87]), .ZN(n579bar);
  OR2_X1 U395 ( .A1(n577), .A2(n576), .ZN(n585) );
  AND2_X1 U395bar ( .A1(n577bar), .A2(n576bar), .ZN(n585bar);
  OR2_X1 U396 ( .A1(n575), .A2(n574), .ZN(n576) );
  AND2_X1 U396bar ( .A1(n575bar), .A2(n574bar), .ZN(n576bar);
  OR2_X1 U397 ( .A1(in_21), .A2(in_11), .ZN(n574) );
  AND2_X1 U397bar ( .A1(in_21bar), .A2(in_11bar), .ZN(n574bar);
  OR2_X1 U398 ( .A1(in_5), .A2(in_3), .ZN(n575) );
  AND2_X1 U398bar ( .A1(in_5bar), .A2(in_3bar), .ZN(n575bar);
  OR2_X1 U399 ( .A1(n573), .A2(n572), .ZN(n577) );
  AND2_X1 U399bar ( .A1(n573bar), .A2(n572bar), .ZN(n577bar);
  OR2_X1 U400 ( .A1(in_68), .A2(in_64), .ZN(n572) );
  AND2_X1 U400bar ( .A1(in_68bar), .A2(in_64bar), .ZN(n572bar);
  OR2_X1 U401 ( .A1(in_76), .A2(in_73), .ZN(n573) );
  AND2_X1 U401bar ( .A1(in_76bar), .A2(in_73bar), .ZN(n573bar);
  OR2_X1 U402 ( .A1(n778), .A2(n571), .ZN(n601) );
  AND2_X1 U402bar ( .A1(n778bar), .A2(n571bar), .ZN(n601bar);
  OR2_X1 U403 ( .A1(in[100]), .A2(n965), .ZN(n571) );
  AND2_X1 U403bar ( .A1(inbar[100]), .A2(n965bar), .ZN(n571bar);
  OR2_X1 U404 ( .A1(n570), .A2(n569), .ZN(n965) );
  AND2_X1 U404bar ( .A1(n570bar), .A2(n569bar), .ZN(n965bar);
  OR2_X1 U405 ( .A1(n568), .A2(n567), .ZN(n569) );
  AND2_X1 U405bar ( .A1(n568bar), .A2(n567bar), .ZN(n569bar);
  OR2_X1 U406 ( .A1(n566), .A2(n565), .ZN(n567) );
  AND2_X1 U406bar ( .A1(n566bar), .A2(n565bar), .ZN(n567bar);
  OR2_X1 U407 ( .A1(n817), .A2(n750), .ZN(n565) );
  AND2_X1 U407bar ( .A1(n817bar), .A2(n750bar), .ZN(n565bar);
  OR2_X1 U408 ( .A1(n564), .A2(n563), .ZN(n750) );
  AND2_X1 U408bar ( .A1(n564bar), .A2(n563bar), .ZN(n750bar);
  OR2_X1 U409 ( .A1(n562), .A2(n561), .ZN(n563) );
  AND2_X1 U409bar ( .A1(n562bar), .A2(n561bar), .ZN(n563bar);
  OR2_X1 U410 ( .A1(n560), .A2(n559), .ZN(n561) );
  AND2_X1 U410bar ( .A1(n560bar), .A2(n559bar), .ZN(n561bar);
  OR2_X1 U411 ( .A1(in[119]), .A2(in[103]), .ZN(n559) );
  AND2_X1 U411bar ( .A1(inbar[119]), .A2(inbar[103]), .ZN(n559bar);
  OR2_X1 U412 ( .A1(in[137]), .A2(in[133]), .ZN(n560) );
  AND2_X1 U412bar ( .A1(inbar[137]), .A2(inbar[133]), .ZN(n560bar);
  OR2_X1 U413 ( .A1(n558), .A2(n557), .ZN(n562) );
  AND2_X1 U413bar ( .A1(n558bar), .A2(n557bar), .ZN(n562bar);
  OR2_X1 U414 ( .A1(in[176]), .A2(in[173]), .ZN(n557) );
  AND2_X1 U414bar ( .A1(inbar[176]), .A2(inbar[173]), .ZN(n557bar);
  OR2_X1 U415 ( .A1(in[210]), .A2(in[181]), .ZN(n558) );
  AND2_X1 U415bar ( .A1(inbar[210]), .A2(inbar[181]), .ZN(n558bar);
  OR2_X1 U416 ( .A1(n556), .A2(n555), .ZN(n564) );
  AND2_X1 U416bar ( .A1(n556bar), .A2(n555bar), .ZN(n564bar);
  OR2_X1 U417 ( .A1(n554), .A2(n553), .ZN(n555) );
  AND2_X1 U417bar ( .A1(n554bar), .A2(n553bar), .ZN(n555bar);
  OR2_X1 U418 ( .A1(in_13), .A2(in[234]), .ZN(n553) );
  AND2_X1 U418bar ( .A1(in_13bar), .A2(inbar[234]), .ZN(n553bar);
  OR2_X1 U419 ( .A1(in_38), .A2(in_32), .ZN(n554) );
  AND2_X1 U419bar ( .A1(in_38bar), .A2(in_32bar), .ZN(n554bar);
  OR2_X1 U420 ( .A1(n552), .A2(n551), .ZN(n556) );
  AND2_X1 U420bar ( .A1(n552bar), .A2(n551bar), .ZN(n556bar);
  OR2_X1 U421 ( .A1(in_42), .A2(in_41), .ZN(n551) );
  AND2_X1 U421bar ( .A1(in_42bar), .A2(in_41bar), .ZN(n551bar);
  OR2_X1 U422 ( .A1(in_7), .A2(in_49), .ZN(n552) );
  AND2_X1 U422bar ( .A1(in_7bar), .A2(in_49bar), .ZN(n552bar);
  OR2_X1 U423 ( .A1(n550), .A2(n549), .ZN(n817) );
  AND2_X1 U423bar ( .A1(n550bar), .A2(n549bar), .ZN(n817bar);
  OR2_X1 U424 ( .A1(n548), .A2(n547), .ZN(n549) );
  AND2_X1 U424bar ( .A1(n548bar), .A2(n547bar), .ZN(n549bar);
  OR2_X1 U425 ( .A1(n546), .A2(n545), .ZN(n547) );
  AND2_X1 U425bar ( .A1(n546bar), .A2(n545bar), .ZN(n547bar);
  OR2_X1 U426 ( .A1(in[159]), .A2(in[105]), .ZN(n545) );
  AND2_X1 U426bar ( .A1(inbar[159]), .A2(inbar[105]), .ZN(n545bar);
  OR2_X1 U427 ( .A1(in[206]), .A2(in[183]), .ZN(n546) );
  AND2_X1 U427bar ( .A1(inbar[206]), .A2(inbar[183]), .ZN(n546bar);
  OR2_X1 U428 ( .A1(n544), .A2(n543), .ZN(n548) );
  AND2_X1 U428bar ( .A1(n544bar), .A2(n543bar), .ZN(n548bar);
  OR2_X1 U429 ( .A1(in[229]), .A2(in[219]), .ZN(n543) );
  AND2_X1 U429bar ( .A1(inbar[229]), .A2(inbar[219]), .ZN(n543bar);
  OR2_X1 U430 ( .A1(in[235]), .A2(in[232]), .ZN(n544) );
  AND2_X1 U430bar ( .A1(inbar[235]), .A2(inbar[232]), .ZN(n544bar);
  OR2_X1 U431 ( .A1(n542), .A2(n541), .ZN(n550) );
  AND2_X1 U431bar ( .A1(n542bar), .A2(n541bar), .ZN(n550bar);
  OR2_X1 U432 ( .A1(n540), .A2(n539), .ZN(n541) );
  AND2_X1 U432bar ( .A1(n540bar), .A2(n539bar), .ZN(n541bar);
  OR2_X1 U433 ( .A1(in[249]), .A2(in[242]), .ZN(n539) );
  AND2_X1 U433bar ( .A1(inbar[249]), .A2(inbar[242]), .ZN(n539bar);
  OR2_X1 U434 ( .A1(in[89]), .A2(in[254]), .ZN(n540) );
  AND2_X1 U434bar ( .A1(inbar[89]), .A2(inbar[254]), .ZN(n540bar);
  OR2_X1 U435 ( .A1(n538), .A2(n537), .ZN(n542) );
  AND2_X1 U435bar ( .A1(n538bar), .A2(n537bar), .ZN(n542bar);
  OR2_X1 U436 ( .A1(in_14), .A2(in[99]), .ZN(n537) );
  AND2_X1 U436bar ( .A1(in_14bar), .A2(inbar[99]), .ZN(n537bar);
  OR2_X1 U437 ( .A1(in_60), .A2(in_18), .ZN(n538) );
  AND2_X1 U437bar ( .A1(in_60bar), .A2(in_18bar), .ZN(n538bar);
  OR2_X1 U438 ( .A1(in[113]), .A2(n763), .ZN(n566) );
  AND2_X1 U438bar ( .A1(inbar[113]), .A2(n763bar), .ZN(n566bar);
  OR2_X1 U439 ( .A1(n536), .A2(n535), .ZN(n763) );
  AND2_X1 U439bar ( .A1(n536bar), .A2(n535bar), .ZN(n763bar);
  OR2_X1 U440 ( .A1(n534), .A2(n533), .ZN(n535) );
  AND2_X1 U440bar ( .A1(n534bar), .A2(n533bar), .ZN(n535bar);
  OR2_X1 U441 ( .A1(n532), .A2(n531), .ZN(n533) );
  AND2_X1 U441bar ( .A1(n532bar), .A2(n531bar), .ZN(n533bar);
  OR2_X1 U442 ( .A1(in[115]), .A2(in[110]), .ZN(n531) );
  AND2_X1 U442bar ( .A1(inbar[115]), .A2(inbar[110]), .ZN(n531bar);
  OR2_X1 U443 ( .A1(in[125]), .A2(in[117]), .ZN(n532) );
  AND2_X1 U443bar ( .A1(inbar[125]), .A2(inbar[117]), .ZN(n532bar);
  OR2_X1 U444 ( .A1(n530), .A2(n529), .ZN(n534) );
  AND2_X1 U444bar ( .A1(n530bar), .A2(n529bar), .ZN(n534bar);
  OR2_X1 U445 ( .A1(in[180]), .A2(in[128]), .ZN(n529) );
  AND2_X1 U445bar ( .A1(inbar[180]), .A2(inbar[128]), .ZN(n529bar);
  OR2_X1 U446 ( .A1(in[205]), .A2(in[201]), .ZN(n530) );
  AND2_X1 U446bar ( .A1(inbar[205]), .A2(inbar[201]), .ZN(n530bar);
  OR2_X1 U447 ( .A1(n528), .A2(n527), .ZN(n536) );
  AND2_X1 U447bar ( .A1(n528bar), .A2(n527bar), .ZN(n536bar);
  OR2_X1 U448 ( .A1(n526), .A2(n525), .ZN(n527) );
  AND2_X1 U448bar ( .A1(n526bar), .A2(n525bar), .ZN(n527bar);
  OR2_X1 U449 ( .A1(in[244]), .A2(in[239]), .ZN(n525) );
  AND2_X1 U449bar ( .A1(inbar[244]), .A2(inbar[239]), .ZN(n525bar);
  OR2_X1 U450 ( .A1(in[95]), .A2(in[83]), .ZN(n526) );
  AND2_X1 U450bar ( .A1(inbar[95]), .A2(inbar[83]), .ZN(n526bar);
  OR2_X1 U451 ( .A1(n524), .A2(n523), .ZN(n528) );
  AND2_X1 U451bar ( .A1(n524bar), .A2(n523bar), .ZN(n528bar);
  OR2_X1 U452 ( .A1(in_24), .A2(in[97]), .ZN(n523) );
  AND2_X1 U452bar ( .A1(in_24bar), .A2(inbar[97]), .ZN(n523bar);
  OR2_X1 U453 ( .A1(in_33), .A2(in_27), .ZN(n524) );
  AND2_X1 U453bar ( .A1(in_33bar), .A2(in_27bar), .ZN(n524bar);
  OR2_X1 U454 ( .A1(n522), .A2(n521), .ZN(n568) );
  AND2_X1 U454bar ( .A1(n522bar), .A2(n521bar), .ZN(n568bar);
  OR2_X1 U455 ( .A1(in[145]), .A2(in[126]), .ZN(n521) );
  AND2_X1 U455bar ( .A1(inbar[145]), .A2(inbar[126]), .ZN(n521bar);
  OR2_X1 U456 ( .A1(in[169]), .A2(n520), .ZN(n522) );
  AND2_X1 U456bar ( .A1(inbar[169]), .A2(n520bar), .ZN(n522bar);
  OR2_X1 U457 ( .A1(in[221]), .A2(in[172]), .ZN(n520) );
  AND2_X1 U457bar ( .A1(inbar[221]), .A2(inbar[172]), .ZN(n520bar);
  OR2_X1 U458 ( .A1(n519), .A2(n518), .ZN(n570) );
  AND2_X1 U458bar ( .A1(n519bar), .A2(n518bar), .ZN(n570bar);
  OR2_X1 U459 ( .A1(n517), .A2(n516), .ZN(n518) );
  AND2_X1 U459bar ( .A1(n517bar), .A2(n516bar), .ZN(n518bar);
  OR2_X1 U460 ( .A1(in[241]), .A2(in[224]), .ZN(n516) );
  AND2_X1 U460bar ( .A1(inbar[241]), .A2(inbar[224]), .ZN(n516bar);
  OR2_X1 U461 ( .A1(in[86]), .A2(n515), .ZN(n517) );
  AND2_X1 U461bar ( .A1(inbar[86]), .A2(n515bar), .ZN(n517bar);
  OR2_X1 U462 ( .A1(in_43), .A2(in_34), .ZN(n515) );
  AND2_X1 U462bar ( .A1(in_43bar), .A2(in_34bar), .ZN(n515bar);
  OR2_X1 U463 ( .A1(n514), .A2(n513), .ZN(n519) );
  AND2_X1 U463bar ( .A1(n514bar), .A2(n513bar), .ZN(n519bar);
  OR2_X1 U464 ( .A1(in_65), .A2(in_51), .ZN(n513) );
  AND2_X1 U464bar ( .A1(in_65bar), .A2(in_51bar), .ZN(n513bar);
  OR2_X1 U465 ( .A1(in_75), .A2(n512), .ZN(n514) );
  AND2_X1 U465bar ( .A1(in_75bar), .A2(n512bar), .ZN(n514bar);
  OR2_X1 U466 ( .A1(in_81), .A2(in_77), .ZN(n512) );
  AND2_X1 U466bar ( .A1(in_81bar), .A2(in_77bar), .ZN(n512bar);
  OR2_X1 U467 ( .A1(n511), .A2(n510), .ZN(n778) );
  AND2_X1 U467bar ( .A1(n511bar), .A2(n510bar), .ZN(n778bar);
  OR2_X1 U468 ( .A1(n509), .A2(n508), .ZN(n510) );
  AND2_X1 U468bar ( .A1(n509bar), .A2(n508bar), .ZN(n510bar);
  OR2_X1 U469 ( .A1(n507), .A2(n506), .ZN(n508) );
  AND2_X1 U469bar ( .A1(n507bar), .A2(n506bar), .ZN(n508bar);
  OR2_X1 U470 ( .A1(in[107]), .A2(in[101]), .ZN(n506) );
  AND2_X1 U470bar ( .A1(inbar[107]), .A2(inbar[101]), .ZN(n506bar);
  OR2_X1 U471 ( .A1(in[139]), .A2(in[132]), .ZN(n507) );
  AND2_X1 U471bar ( .A1(inbar[139]), .A2(inbar[132]), .ZN(n507bar);
  OR2_X1 U472 ( .A1(n505), .A2(n504), .ZN(n509) );
  AND2_X1 U472bar ( .A1(n505bar), .A2(n504bar), .ZN(n509bar);
  OR2_X1 U473 ( .A1(in[146]), .A2(in[141]), .ZN(n504) );
  AND2_X1 U473bar ( .A1(inbar[146]), .A2(inbar[141]), .ZN(n504bar);
  OR2_X1 U474 ( .A1(in[203]), .A2(in[179]), .ZN(n505) );
  AND2_X1 U474bar ( .A1(inbar[203]), .A2(inbar[179]), .ZN(n505bar);
  OR2_X1 U475 ( .A1(n503), .A2(n502), .ZN(n511) );
  AND2_X1 U475bar ( .A1(n503bar), .A2(n502bar), .ZN(n511bar);
  OR2_X1 U476 ( .A1(n501), .A2(n500), .ZN(n502) );
  AND2_X1 U476bar ( .A1(n501bar), .A2(n500bar), .ZN(n502bar);
  OR2_X1 U477 ( .A1(in[243]), .A2(in[222]), .ZN(n500) );
  AND2_X1 U477bar ( .A1(inbar[243]), .A2(inbar[222]), .ZN(n500bar);
  OR2_X1 U478 ( .A1(in[251]), .A2(in[250]), .ZN(n501) );
  AND2_X1 U478bar ( .A1(inbar[251]), .A2(inbar[250]), .ZN(n501bar);
  OR2_X1 U479 ( .A1(n499), .A2(n498), .ZN(n503) );
  AND2_X1 U479bar ( .A1(n499bar), .A2(n498bar), .ZN(n503bar);
  OR2_X1 U480 ( .A1(in_37), .A2(in_19), .ZN(n498) );
  AND2_X1 U480bar ( .A1(in_37bar), .A2(in_19bar), .ZN(n498bar);
  OR2_X1 U481 ( .A1(in_78), .A2(in_6), .ZN(n499) );
  AND2_X1 U481bar ( .A1(in_78bar), .A2(in_6bar), .ZN(n499bar);
  OR2_X1 U482 ( .A1(n497), .A2(n496), .ZN(n603) );
  AND2_X1 U482bar ( .A1(n497bar), .A2(n496bar), .ZN(n603bar);
  OR2_X1 U483 ( .A1(in[112]), .A2(in[102]), .ZN(n496) );
  AND2_X1 U483bar ( .A1(inbar[112]), .A2(inbar[102]), .ZN(n496bar);
  OR2_X1 U484 ( .A1(in[123]), .A2(n495), .ZN(n497) );
  AND2_X1 U484bar ( .A1(inbar[123]), .A2(n495bar), .ZN(n497bar);
  OR2_X1 U485 ( .A1(in[143]), .A2(in[130]), .ZN(n495) );
  AND2_X1 U485bar ( .A1(inbar[143]), .A2(inbar[130]), .ZN(n495bar);
  OR2_X1 U486 ( .A1(n494), .A2(n493), .ZN(n605) );
  AND2_X1 U486bar ( .A1(n494bar), .A2(n493bar), .ZN(n605bar);
  OR2_X1 U487 ( .A1(n492), .A2(n491), .ZN(n493) );
  AND2_X1 U487bar ( .A1(n492bar), .A2(n491bar), .ZN(n493bar);
  OR2_X1 U488 ( .A1(in[216]), .A2(in[213]), .ZN(n491) );
  AND2_X1 U488bar ( .A1(inbar[216]), .A2(inbar[213]), .ZN(n491bar);
  OR2_X1 U489 ( .A1(in[227]), .A2(n490), .ZN(n492) );
  AND2_X1 U489bar ( .A1(inbar[227]), .A2(n490bar), .ZN(n492bar);
  OR2_X1 U490 ( .A1(in_0), .A2(in[248]), .ZN(n490) );
  AND2_X1 U490bar ( .A1(in_0bar), .A2(inbar[248]), .ZN(n490bar);
  OR2_X1 U491 ( .A1(n489), .A2(n488), .ZN(n494) );
  AND2_X1 U491bar ( .A1(n489bar), .A2(n488bar), .ZN(n494bar);
  OR2_X1 U492 ( .A1(in_46), .A2(in_44), .ZN(n488) );
  AND2_X1 U492bar ( .A1(in_46bar), .A2(in_44bar), .ZN(n488bar);
  OR2_X1 U493 ( .A1(in_50), .A2(n487), .ZN(n489) );
  AND2_X1 U493bar ( .A1(in_50bar), .A2(n487bar), .ZN(n489bar);
  OR2_X1 U494 ( .A1(in_9), .A2(in_80), .ZN(n487) );
  AND2_X1 U494bar ( .A1(in_9bar), .A2(in_80bar), .ZN(n487bar);
endmodule




module sBox_17 ( in, out );
  input [7:0] in;
  //input_done

  output [7:0] out;
  //output_done

  wire   [255:0] decodeOut;
  //wire_done

  decode_17 dec ( .in(in), .out(decodeOut) );
  encode_17 enc ( .in(decodeOut), .out(out) );
endmodule


module CD2_69 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_70 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_71 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_72 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD4_35 ( a, b, y );
  input [3:0] a;
  input [3:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  //input_done

  output [15:0] y;
  reg [15:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]);
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]);
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]);
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]);
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]);
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]);
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]);
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]);
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]);
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]);
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]);
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]);
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]);
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]);
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]);
endmodule




module CD4_36 ( a, b, y );
  input [3:0] a;
  input [3:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  //input_done

  output [15:0] y;
  reg [15:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]);
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]);
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]);
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]);
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]);
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]);
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]);
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]);
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]);
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]);
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]);
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]);
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]);
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]);
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]);
endmodule




module CD16_18 ( a, b, y );
  input [15:0] a;
  input [15:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign abar[8] = ~a[8];
  assign abar[9] = ~a[9];
  assign abar[10] = ~a[10];
  assign abar[11] = ~a[11];
  assign abar[12] = ~a[12];
  assign abar[13] = ~a[13];
  assign abar[14] = ~a[14];
  assign abar[15] = ~a[15];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign bbar[8] = ~b[8];
  assign bbar[9] = ~b[9];
  assign bbar[10] = ~b[10];
  assign bbar[11] = ~b[11];
  assign bbar[12] = ~b[12];
  assign bbar[13] = ~b[13];
  assign bbar[14] = ~b[14];
  assign bbar[15] = ~b[15];
  //input_done

  output [15:0] y;
  reg [15:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[9]), .A2(a[0]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[9]), .A2(abar[0]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[3]), .A2(a[6]), .ZN(y[99]) );
  OR2_X1 U2bar ( .A1(bbar[3]), .A2(abar[6]), .ZN(ybar[99]);
  AND2_X1 U3 ( .A1(b[2]), .A2(a[6]), .ZN(y[98]) );
  OR2_X1 U3bar ( .A1(bbar[2]), .A2(abar[6]), .ZN(ybar[98]);
  AND2_X1 U4 ( .A1(b[1]), .A2(a[6]), .ZN(y[97]) );
  OR2_X1 U4bar ( .A1(bbar[1]), .A2(abar[6]), .ZN(ybar[97]);
  AND2_X1 U5 ( .A1(b[0]), .A2(a[6]), .ZN(y[96]) );
  OR2_X1 U5bar ( .A1(bbar[0]), .A2(abar[6]), .ZN(ybar[96]);
  AND2_X1 U6 ( .A1(b[15]), .A2(a[5]), .ZN(y[95]) );
  OR2_X1 U6bar ( .A1(bbar[15]), .A2(abar[5]), .ZN(ybar[95]);
  AND2_X1 U7 ( .A1(b[14]), .A2(a[5]), .ZN(y[94]) );
  OR2_X1 U7bar ( .A1(bbar[14]), .A2(abar[5]), .ZN(ybar[94]);
  AND2_X1 U8 ( .A1(b[13]), .A2(a[5]), .ZN(y[93]) );
  OR2_X1 U8bar ( .A1(bbar[13]), .A2(abar[5]), .ZN(ybar[93]);
  AND2_X1 U9 ( .A1(b[12]), .A2(a[5]), .ZN(y[92]) );
  OR2_X1 U9bar ( .A1(bbar[12]), .A2(abar[5]), .ZN(ybar[92]);
  AND2_X1 U10 ( .A1(b[11]), .A2(a[5]), .ZN(y[91]) );
  OR2_X1 U10bar ( .A1(bbar[11]), .A2(abar[5]), .ZN(ybar[91]);
  AND2_X1 U11 ( .A1(b[10]), .A2(a[5]), .ZN(y[90]) );
  OR2_X1 U11bar ( .A1(bbar[10]), .A2(abar[5]), .ZN(ybar[90]);
  AND2_X1 U12 ( .A1(b[8]), .A2(a[0]), .ZN(y[8]) );
  OR2_X1 U12bar ( .A1(bbar[8]), .A2(abar[0]), .ZN(ybar[8]);
  AND2_X1 U13 ( .A1(a[5]), .A2(b[9]), .ZN(y[89]) );
  OR2_X1 U13bar ( .A1(abar[5]), .A2(bbar[9]), .ZN(ybar[89]);
  AND2_X1 U14 ( .A1(b[8]), .A2(a[5]), .ZN(y[88]) );
  OR2_X1 U14bar ( .A1(bbar[8]), .A2(abar[5]), .ZN(ybar[88]);
  AND2_X1 U15 ( .A1(b[7]), .A2(a[5]), .ZN(y[87]) );
  OR2_X1 U15bar ( .A1(bbar[7]), .A2(abar[5]), .ZN(ybar[87]);
  AND2_X1 U16 ( .A1(b[6]), .A2(a[5]), .ZN(y[86]) );
  OR2_X1 U16bar ( .A1(bbar[6]), .A2(abar[5]), .ZN(ybar[86]);
  AND2_X1 U17 ( .A1(b[5]), .A2(a[5]), .ZN(y[85]) );
  OR2_X1 U17bar ( .A1(bbar[5]), .A2(abar[5]), .ZN(ybar[85]);
  AND2_X1 U18 ( .A1(b[4]), .A2(a[5]), .ZN(y[84]) );
  OR2_X1 U18bar ( .A1(bbar[4]), .A2(abar[5]), .ZN(ybar[84]);
  AND2_X1 U19 ( .A1(a[5]), .A2(b[3]), .ZN(y[83]) );
  OR2_X1 U19bar ( .A1(abar[5]), .A2(bbar[3]), .ZN(ybar[83]);
  AND2_X1 U20 ( .A1(a[5]), .A2(b[2]), .ZN(y[82]) );
  OR2_X1 U20bar ( .A1(abar[5]), .A2(bbar[2]), .ZN(ybar[82]);
  AND2_X1 U21 ( .A1(a[5]), .A2(b[1]), .ZN(y[81]) );
  OR2_X1 U21bar ( .A1(abar[5]), .A2(bbar[1]), .ZN(ybar[81]);
  AND2_X1 U22 ( .A1(a[5]), .A2(b[0]), .ZN(y[80]) );
  OR2_X1 U22bar ( .A1(abar[5]), .A2(bbar[0]), .ZN(ybar[80]);
  AND2_X1 U23 ( .A1(b[7]), .A2(a[0]), .ZN(y[7]) );
  OR2_X1 U23bar ( .A1(bbar[7]), .A2(abar[0]), .ZN(ybar[7]);
  AND2_X1 U24 ( .A1(a[4]), .A2(b[15]), .ZN(y[79]) );
  OR2_X1 U24bar ( .A1(abar[4]), .A2(bbar[15]), .ZN(ybar[79]);
  AND2_X1 U25 ( .A1(a[4]), .A2(b[14]), .ZN(y[78]) );
  OR2_X1 U25bar ( .A1(abar[4]), .A2(bbar[14]), .ZN(ybar[78]);
  AND2_X1 U26 ( .A1(a[4]), .A2(b[13]), .ZN(y[77]) );
  OR2_X1 U26bar ( .A1(abar[4]), .A2(bbar[13]), .ZN(ybar[77]);
  AND2_X1 U27 ( .A1(a[4]), .A2(b[12]), .ZN(y[76]) );
  OR2_X1 U27bar ( .A1(abar[4]), .A2(bbar[12]), .ZN(ybar[76]);
  AND2_X1 U28 ( .A1(a[4]), .A2(b[11]), .ZN(y[75]) );
  OR2_X1 U28bar ( .A1(abar[4]), .A2(bbar[11]), .ZN(ybar[75]);
  AND2_X1 U29 ( .A1(a[4]), .A2(b[10]), .ZN(y[74]) );
  OR2_X1 U29bar ( .A1(abar[4]), .A2(bbar[10]), .ZN(ybar[74]);
  AND2_X1 U30 ( .A1(a[4]), .A2(b[9]), .ZN(y[73]) );
  OR2_X1 U30bar ( .A1(abar[4]), .A2(bbar[9]), .ZN(ybar[73]);
  AND2_X1 U31 ( .A1(a[4]), .A2(b[8]), .ZN(y[72]) );
  OR2_X1 U31bar ( .A1(abar[4]), .A2(bbar[8]), .ZN(ybar[72]);
  AND2_X1 U32 ( .A1(a[4]), .A2(b[7]), .ZN(y[71]) );
  OR2_X1 U32bar ( .A1(abar[4]), .A2(bbar[7]), .ZN(ybar[71]);
  AND2_X1 U33 ( .A1(a[4]), .A2(b[6]), .ZN(y[70]) );
  OR2_X1 U33bar ( .A1(abar[4]), .A2(bbar[6]), .ZN(ybar[70]);
  AND2_X1 U34 ( .A1(b[6]), .A2(a[0]), .ZN(y[6]) );
  OR2_X1 U34bar ( .A1(bbar[6]), .A2(abar[0]), .ZN(ybar[6]);
  AND2_X1 U35 ( .A1(a[4]), .A2(b[5]), .ZN(y[69]) );
  OR2_X1 U35bar ( .A1(abar[4]), .A2(bbar[5]), .ZN(ybar[69]);
  AND2_X1 U36 ( .A1(a[4]), .A2(b[4]), .ZN(y[68]) );
  OR2_X1 U36bar ( .A1(abar[4]), .A2(bbar[4]), .ZN(ybar[68]);
  AND2_X1 U37 ( .A1(a[4]), .A2(b[3]), .ZN(y[67]) );
  OR2_X1 U37bar ( .A1(abar[4]), .A2(bbar[3]), .ZN(ybar[67]);
  AND2_X1 U38 ( .A1(a[4]), .A2(b[2]), .ZN(y[66]) );
  OR2_X1 U38bar ( .A1(abar[4]), .A2(bbar[2]), .ZN(ybar[66]);
  AND2_X1 U39 ( .A1(a[4]), .A2(b[1]), .ZN(y[65]) );
  OR2_X1 U39bar ( .A1(abar[4]), .A2(bbar[1]), .ZN(ybar[65]);
  AND2_X1 U40 ( .A1(a[4]), .A2(b[0]), .ZN(y[64]) );
  OR2_X1 U40bar ( .A1(abar[4]), .A2(bbar[0]), .ZN(ybar[64]);
  AND2_X1 U41 ( .A1(a[3]), .A2(b[15]), .ZN(y[63]) );
  OR2_X1 U41bar ( .A1(abar[3]), .A2(bbar[15]), .ZN(ybar[63]);
  AND2_X1 U42 ( .A1(a[3]), .A2(b[14]), .ZN(y[62]) );
  OR2_X1 U42bar ( .A1(abar[3]), .A2(bbar[14]), .ZN(ybar[62]);
  AND2_X1 U43 ( .A1(a[3]), .A2(b[13]), .ZN(y[61]) );
  OR2_X1 U43bar ( .A1(abar[3]), .A2(bbar[13]), .ZN(ybar[61]);
  AND2_X1 U44 ( .A1(a[3]), .A2(b[12]), .ZN(y[60]) );
  OR2_X1 U44bar ( .A1(abar[3]), .A2(bbar[12]), .ZN(ybar[60]);
  AND2_X1 U45 ( .A1(b[5]), .A2(a[0]), .ZN(y[5]) );
  OR2_X1 U45bar ( .A1(bbar[5]), .A2(abar[0]), .ZN(ybar[5]);
  AND2_X1 U46 ( .A1(a[3]), .A2(b[11]), .ZN(y[59]) );
  OR2_X1 U46bar ( .A1(abar[3]), .A2(bbar[11]), .ZN(ybar[59]);
  AND2_X1 U47 ( .A1(a[3]), .A2(b[10]), .ZN(y[58]) );
  OR2_X1 U47bar ( .A1(abar[3]), .A2(bbar[10]), .ZN(ybar[58]);
  AND2_X1 U48 ( .A1(a[3]), .A2(b[9]), .ZN(y[57]) );
  OR2_X1 U48bar ( .A1(abar[3]), .A2(bbar[9]), .ZN(ybar[57]);
  AND2_X1 U49 ( .A1(a[3]), .A2(b[8]), .ZN(y[56]) );
  OR2_X1 U49bar ( .A1(abar[3]), .A2(bbar[8]), .ZN(ybar[56]);
  AND2_X1 U50 ( .A1(a[3]), .A2(b[7]), .ZN(y[55]) );
  OR2_X1 U50bar ( .A1(abar[3]), .A2(bbar[7]), .ZN(ybar[55]);
  AND2_X1 U51 ( .A1(a[3]), .A2(b[6]), .ZN(y[54]) );
  OR2_X1 U51bar ( .A1(abar[3]), .A2(bbar[6]), .ZN(ybar[54]);
  AND2_X1 U52 ( .A1(a[3]), .A2(b[5]), .ZN(y[53]) );
  OR2_X1 U52bar ( .A1(abar[3]), .A2(bbar[5]), .ZN(ybar[53]);
  AND2_X1 U53 ( .A1(a[3]), .A2(b[4]), .ZN(y[52]) );
  OR2_X1 U53bar ( .A1(abar[3]), .A2(bbar[4]), .ZN(ybar[52]);
  AND2_X1 U54 ( .A1(a[3]), .A2(b[3]), .ZN(y[51]) );
  OR2_X1 U54bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[51]);
  AND2_X1 U55 ( .A1(a[3]), .A2(b[2]), .ZN(y[50]) );
  OR2_X1 U55bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[50]);
  AND2_X1 U56 ( .A1(b[4]), .A2(a[0]), .ZN(y[4]) );
  OR2_X1 U56bar ( .A1(bbar[4]), .A2(abar[0]), .ZN(ybar[4]);
  AND2_X1 U57 ( .A1(a[3]), .A2(b[1]), .ZN(y[49]) );
  OR2_X1 U57bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[49]);
  AND2_X1 U58 ( .A1(a[3]), .A2(b[0]), .ZN(y[48]) );
  OR2_X1 U58bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[48]);
  AND2_X1 U59 ( .A1(a[2]), .A2(b[15]), .ZN(y[47]) );
  OR2_X1 U59bar ( .A1(abar[2]), .A2(bbar[15]), .ZN(ybar[47]);
  AND2_X1 U60 ( .A1(a[2]), .A2(b[14]), .ZN(y[46]) );
  OR2_X1 U60bar ( .A1(abar[2]), .A2(bbar[14]), .ZN(ybar[46]);
  AND2_X1 U61 ( .A1(a[2]), .A2(b[13]), .ZN(y[45]) );
  OR2_X1 U61bar ( .A1(abar[2]), .A2(bbar[13]), .ZN(ybar[45]);
  AND2_X1 U62 ( .A1(a[2]), .A2(b[12]), .ZN(y[44]) );
  OR2_X1 U62bar ( .A1(abar[2]), .A2(bbar[12]), .ZN(ybar[44]);
  AND2_X1 U63 ( .A1(a[2]), .A2(b[11]), .ZN(y[43]) );
  OR2_X1 U63bar ( .A1(abar[2]), .A2(bbar[11]), .ZN(ybar[43]);
  AND2_X1 U64 ( .A1(a[2]), .A2(b[10]), .ZN(y[42]) );
  OR2_X1 U64bar ( .A1(abar[2]), .A2(bbar[10]), .ZN(ybar[42]);
  AND2_X1 U65 ( .A1(a[2]), .A2(b[9]), .ZN(y[41]) );
  OR2_X1 U65bar ( .A1(abar[2]), .A2(bbar[9]), .ZN(ybar[41]);
  AND2_X1 U66 ( .A1(a[2]), .A2(b[8]), .ZN(y[40]) );
  OR2_X1 U66bar ( .A1(abar[2]), .A2(bbar[8]), .ZN(ybar[40]);
  AND2_X1 U67 ( .A1(b[3]), .A2(a[0]), .ZN(y[3]) );
  OR2_X1 U67bar ( .A1(bbar[3]), .A2(abar[0]), .ZN(ybar[3]);
  AND2_X1 U68 ( .A1(a[2]), .A2(b[7]), .ZN(y[39]) );
  OR2_X1 U68bar ( .A1(abar[2]), .A2(bbar[7]), .ZN(ybar[39]);
  AND2_X1 U69 ( .A1(a[2]), .A2(b[6]), .ZN(y[38]) );
  OR2_X1 U69bar ( .A1(abar[2]), .A2(bbar[6]), .ZN(ybar[38]);
  AND2_X1 U70 ( .A1(a[2]), .A2(b[5]), .ZN(y[37]) );
  OR2_X1 U70bar ( .A1(abar[2]), .A2(bbar[5]), .ZN(ybar[37]);
  AND2_X1 U71 ( .A1(a[2]), .A2(b[4]), .ZN(y[36]) );
  OR2_X1 U71bar ( .A1(abar[2]), .A2(bbar[4]), .ZN(ybar[36]);
  AND2_X1 U72 ( .A1(a[2]), .A2(b[3]), .ZN(y[35]) );
  OR2_X1 U72bar ( .A1(abar[2]), .A2(bbar[3]), .ZN(ybar[35]);
  AND2_X1 U73 ( .A1(a[2]), .A2(b[2]), .ZN(y[34]) );
  OR2_X1 U73bar ( .A1(abar[2]), .A2(bbar[2]), .ZN(ybar[34]);
  AND2_X1 U74 ( .A1(a[2]), .A2(b[1]), .ZN(y[33]) );
  OR2_X1 U74bar ( .A1(abar[2]), .A2(bbar[1]), .ZN(ybar[33]);
  AND2_X1 U75 ( .A1(a[2]), .A2(b[0]), .ZN(y[32]) );
  OR2_X1 U75bar ( .A1(abar[2]), .A2(bbar[0]), .ZN(ybar[32]);
  AND2_X1 U76 ( .A1(a[1]), .A2(b[15]), .ZN(y[31]) );
  OR2_X1 U76bar ( .A1(abar[1]), .A2(bbar[15]), .ZN(ybar[31]);
  AND2_X1 U77 ( .A1(a[1]), .A2(b[14]), .ZN(y[30]) );
  OR2_X1 U77bar ( .A1(abar[1]), .A2(bbar[14]), .ZN(ybar[30]);
  AND2_X1 U78 ( .A1(b[2]), .A2(a[0]), .ZN(y[2]) );
  OR2_X1 U78bar ( .A1(bbar[2]), .A2(abar[0]), .ZN(ybar[2]);
  AND2_X1 U79 ( .A1(a[1]), .A2(b[13]), .ZN(y[29]) );
  OR2_X1 U79bar ( .A1(abar[1]), .A2(bbar[13]), .ZN(ybar[29]);
  AND2_X1 U80 ( .A1(a[1]), .A2(b[12]), .ZN(y[28]) );
  OR2_X1 U80bar ( .A1(abar[1]), .A2(bbar[12]), .ZN(ybar[28]);
  AND2_X1 U81 ( .A1(a[1]), .A2(b[11]), .ZN(y[27]) );
  OR2_X1 U81bar ( .A1(abar[1]), .A2(bbar[11]), .ZN(ybar[27]);
  AND2_X1 U82 ( .A1(a[1]), .A2(b[10]), .ZN(y[26]) );
  OR2_X1 U82bar ( .A1(abar[1]), .A2(bbar[10]), .ZN(ybar[26]);
  AND2_X1 U83 ( .A1(a[1]), .A2(b[9]), .ZN(y[25]) );
  OR2_X1 U83bar ( .A1(abar[1]), .A2(bbar[9]), .ZN(ybar[25]);
  AND2_X1 U84 ( .A1(a[15]), .A2(b[15]), .ZN(y[255]) );
  OR2_X1 U84bar ( .A1(abar[15]), .A2(bbar[15]), .ZN(ybar[255]);
  AND2_X1 U85 ( .A1(a[15]), .A2(b[14]), .ZN(y[254]) );
  OR2_X1 U85bar ( .A1(abar[15]), .A2(bbar[14]), .ZN(ybar[254]);
  AND2_X1 U86 ( .A1(a[15]), .A2(b[13]), .ZN(y[253]) );
  OR2_X1 U86bar ( .A1(abar[15]), .A2(bbar[13]), .ZN(ybar[253]);
  AND2_X1 U87 ( .A1(a[15]), .A2(b[12]), .ZN(y[252]) );
  OR2_X1 U87bar ( .A1(abar[15]), .A2(bbar[12]), .ZN(ybar[252]);
  AND2_X1 U88 ( .A1(a[15]), .A2(b[11]), .ZN(y[251]) );
  OR2_X1 U88bar ( .A1(abar[15]), .A2(bbar[11]), .ZN(ybar[251]);
  AND2_X1 U89 ( .A1(a[15]), .A2(b[10]), .ZN(y[250]) );
  OR2_X1 U89bar ( .A1(abar[15]), .A2(bbar[10]), .ZN(ybar[250]);
  AND2_X1 U90 ( .A1(a[1]), .A2(b[8]), .ZN(y[24]) );
  OR2_X1 U90bar ( .A1(abar[1]), .A2(bbar[8]), .ZN(ybar[24]);
  AND2_X1 U91 ( .A1(a[15]), .A2(b[9]), .ZN(y[249]) );
  OR2_X1 U91bar ( .A1(abar[15]), .A2(bbar[9]), .ZN(ybar[249]);
  AND2_X1 U92 ( .A1(a[15]), .A2(b[8]), .ZN(y[248]) );
  OR2_X1 U92bar ( .A1(abar[15]), .A2(bbar[8]), .ZN(ybar[248]);
  AND2_X1 U93 ( .A1(a[15]), .A2(b[7]), .ZN(y[247]) );
  OR2_X1 U93bar ( .A1(abar[15]), .A2(bbar[7]), .ZN(ybar[247]);
  AND2_X1 U94 ( .A1(a[15]), .A2(b[6]), .ZN(y[246]) );
  OR2_X1 U94bar ( .A1(abar[15]), .A2(bbar[6]), .ZN(ybar[246]);
  AND2_X1 U95 ( .A1(a[15]), .A2(b[5]), .ZN(y[245]) );
  OR2_X1 U95bar ( .A1(abar[15]), .A2(bbar[5]), .ZN(ybar[245]);
  AND2_X1 U96 ( .A1(a[15]), .A2(b[4]), .ZN(y[244]) );
  OR2_X1 U96bar ( .A1(abar[15]), .A2(bbar[4]), .ZN(ybar[244]);
  AND2_X1 U97 ( .A1(a[15]), .A2(b[3]), .ZN(y[243]) );
  OR2_X1 U97bar ( .A1(abar[15]), .A2(bbar[3]), .ZN(ybar[243]);
  AND2_X1 U98 ( .A1(a[15]), .A2(b[2]), .ZN(y[242]) );
  OR2_X1 U98bar ( .A1(abar[15]), .A2(bbar[2]), .ZN(ybar[242]);
  AND2_X1 U99 ( .A1(a[15]), .A2(b[1]), .ZN(y[241]) );
  OR2_X1 U99bar ( .A1(abar[15]), .A2(bbar[1]), .ZN(ybar[241]);
  AND2_X1 U100 ( .A1(a[15]), .A2(b[0]), .ZN(y[240]) );
  OR2_X1 U100bar ( .A1(abar[15]), .A2(bbar[0]), .ZN(ybar[240]);
  AND2_X1 U101 ( .A1(a[1]), .A2(b[7]), .ZN(y[23]) );
  OR2_X1 U101bar ( .A1(abar[1]), .A2(bbar[7]), .ZN(ybar[23]);
  AND2_X1 U102 ( .A1(a[14]), .A2(b[15]), .ZN(y[239]) );
  OR2_X1 U102bar ( .A1(abar[14]), .A2(bbar[15]), .ZN(ybar[239]);
  AND2_X1 U103 ( .A1(a[14]), .A2(b[14]), .ZN(y[238]) );
  OR2_X1 U103bar ( .A1(abar[14]), .A2(bbar[14]), .ZN(ybar[238]);
  AND2_X1 U104 ( .A1(a[14]), .A2(b[13]), .ZN(y[237]) );
  OR2_X1 U104bar ( .A1(abar[14]), .A2(bbar[13]), .ZN(ybar[237]);
  AND2_X1 U105 ( .A1(a[14]), .A2(b[12]), .ZN(y[236]) );
  OR2_X1 U105bar ( .A1(abar[14]), .A2(bbar[12]), .ZN(ybar[236]);
  AND2_X1 U106 ( .A1(a[14]), .A2(b[11]), .ZN(y[235]) );
  OR2_X1 U106bar ( .A1(abar[14]), .A2(bbar[11]), .ZN(ybar[235]);
  AND2_X1 U107 ( .A1(a[14]), .A2(b[10]), .ZN(y[234]) );
  OR2_X1 U107bar ( .A1(abar[14]), .A2(bbar[10]), .ZN(ybar[234]);
  AND2_X1 U108 ( .A1(a[14]), .A2(b[9]), .ZN(y[233]) );
  OR2_X1 U108bar ( .A1(abar[14]), .A2(bbar[9]), .ZN(ybar[233]);
  AND2_X1 U109 ( .A1(a[14]), .A2(b[8]), .ZN(y[232]) );
  OR2_X1 U109bar ( .A1(abar[14]), .A2(bbar[8]), .ZN(ybar[232]);
  AND2_X1 U110 ( .A1(a[14]), .A2(b[7]), .ZN(y[231]) );
  OR2_X1 U110bar ( .A1(abar[14]), .A2(bbar[7]), .ZN(ybar[231]);
  AND2_X1 U111 ( .A1(a[14]), .A2(b[6]), .ZN(y[230]) );
  OR2_X1 U111bar ( .A1(abar[14]), .A2(bbar[6]), .ZN(ybar[230]);
  AND2_X1 U112 ( .A1(a[1]), .A2(b[6]), .ZN(y[22]) );
  OR2_X1 U112bar ( .A1(abar[1]), .A2(bbar[6]), .ZN(ybar[22]);
  AND2_X1 U113 ( .A1(a[14]), .A2(b[5]), .ZN(y[229]) );
  OR2_X1 U113bar ( .A1(abar[14]), .A2(bbar[5]), .ZN(ybar[229]);
  AND2_X1 U114 ( .A1(a[14]), .A2(b[4]), .ZN(y[228]) );
  OR2_X1 U114bar ( .A1(abar[14]), .A2(bbar[4]), .ZN(ybar[228]);
  AND2_X1 U115 ( .A1(a[14]), .A2(b[3]), .ZN(y[227]) );
  OR2_X1 U115bar ( .A1(abar[14]), .A2(bbar[3]), .ZN(ybar[227]);
  AND2_X1 U116 ( .A1(a[14]), .A2(b[2]), .ZN(y[226]) );
  OR2_X1 U116bar ( .A1(abar[14]), .A2(bbar[2]), .ZN(ybar[226]);
  AND2_X1 U117 ( .A1(a[14]), .A2(b[1]), .ZN(y[225]) );
  OR2_X1 U117bar ( .A1(abar[14]), .A2(bbar[1]), .ZN(ybar[225]);
  AND2_X1 U118 ( .A1(a[14]), .A2(b[0]), .ZN(y[224]) );
  OR2_X1 U118bar ( .A1(abar[14]), .A2(bbar[0]), .ZN(ybar[224]);
  AND2_X1 U119 ( .A1(a[13]), .A2(b[15]), .ZN(y[223]) );
  OR2_X1 U119bar ( .A1(abar[13]), .A2(bbar[15]), .ZN(ybar[223]);
  AND2_X1 U120 ( .A1(a[13]), .A2(b[14]), .ZN(y[222]) );
  OR2_X1 U120bar ( .A1(abar[13]), .A2(bbar[14]), .ZN(ybar[222]);
  AND2_X1 U121 ( .A1(a[13]), .A2(b[13]), .ZN(y[221]) );
  OR2_X1 U121bar ( .A1(abar[13]), .A2(bbar[13]), .ZN(ybar[221]);
  AND2_X1 U122 ( .A1(a[13]), .A2(b[12]), .ZN(y[220]) );
  OR2_X1 U122bar ( .A1(abar[13]), .A2(bbar[12]), .ZN(ybar[220]);
  AND2_X1 U123 ( .A1(a[1]), .A2(b[5]), .ZN(y[21]) );
  OR2_X1 U123bar ( .A1(abar[1]), .A2(bbar[5]), .ZN(ybar[21]);
  AND2_X1 U124 ( .A1(a[13]), .A2(b[11]), .ZN(y[219]) );
  OR2_X1 U124bar ( .A1(abar[13]), .A2(bbar[11]), .ZN(ybar[219]);
  AND2_X1 U125 ( .A1(a[13]), .A2(b[10]), .ZN(y[218]) );
  OR2_X1 U125bar ( .A1(abar[13]), .A2(bbar[10]), .ZN(ybar[218]);
  AND2_X1 U126 ( .A1(a[13]), .A2(b[9]), .ZN(y[217]) );
  OR2_X1 U126bar ( .A1(abar[13]), .A2(bbar[9]), .ZN(ybar[217]);
  AND2_X1 U127 ( .A1(a[13]), .A2(b[8]), .ZN(y[216]) );
  OR2_X1 U127bar ( .A1(abar[13]), .A2(bbar[8]), .ZN(ybar[216]);
  AND2_X1 U128 ( .A1(a[13]), .A2(b[7]), .ZN(y[215]) );
  OR2_X1 U128bar ( .A1(abar[13]), .A2(bbar[7]), .ZN(ybar[215]);
  AND2_X1 U129 ( .A1(a[13]), .A2(b[6]), .ZN(y[214]) );
  OR2_X1 U129bar ( .A1(abar[13]), .A2(bbar[6]), .ZN(ybar[214]);
  AND2_X1 U130 ( .A1(a[13]), .A2(b[5]), .ZN(y[213]) );
  OR2_X1 U130bar ( .A1(abar[13]), .A2(bbar[5]), .ZN(ybar[213]);
  AND2_X1 U131 ( .A1(a[13]), .A2(b[4]), .ZN(y[212]) );
  OR2_X1 U131bar ( .A1(abar[13]), .A2(bbar[4]), .ZN(ybar[212]);
  AND2_X1 U132 ( .A1(a[13]), .A2(b[3]), .ZN(y[211]) );
  OR2_X1 U132bar ( .A1(abar[13]), .A2(bbar[3]), .ZN(ybar[211]);
  AND2_X1 U133 ( .A1(a[13]), .A2(b[2]), .ZN(y[210]) );
  OR2_X1 U133bar ( .A1(abar[13]), .A2(bbar[2]), .ZN(ybar[210]);
  AND2_X1 U134 ( .A1(a[1]), .A2(b[4]), .ZN(y[20]) );
  OR2_X1 U134bar ( .A1(abar[1]), .A2(bbar[4]), .ZN(ybar[20]);
  AND2_X1 U135 ( .A1(a[13]), .A2(b[1]), .ZN(y[209]) );
  OR2_X1 U135bar ( .A1(abar[13]), .A2(bbar[1]), .ZN(ybar[209]);
  AND2_X1 U136 ( .A1(a[13]), .A2(b[0]), .ZN(y[208]) );
  OR2_X1 U136bar ( .A1(abar[13]), .A2(bbar[0]), .ZN(ybar[208]);
  AND2_X1 U137 ( .A1(a[12]), .A2(b[15]), .ZN(y[207]) );
  OR2_X1 U137bar ( .A1(abar[12]), .A2(bbar[15]), .ZN(ybar[207]);
  AND2_X1 U138 ( .A1(a[12]), .A2(b[14]), .ZN(y[206]) );
  OR2_X1 U138bar ( .A1(abar[12]), .A2(bbar[14]), .ZN(ybar[206]);
  AND2_X1 U139 ( .A1(a[12]), .A2(b[13]), .ZN(y[205]) );
  OR2_X1 U139bar ( .A1(abar[12]), .A2(bbar[13]), .ZN(ybar[205]);
  AND2_X1 U140 ( .A1(a[12]), .A2(b[12]), .ZN(y[204]) );
  OR2_X1 U140bar ( .A1(abar[12]), .A2(bbar[12]), .ZN(ybar[204]);
  AND2_X1 U141 ( .A1(a[12]), .A2(b[11]), .ZN(y[203]) );
  OR2_X1 U141bar ( .A1(abar[12]), .A2(bbar[11]), .ZN(ybar[203]);
  AND2_X1 U142 ( .A1(a[12]), .A2(b[10]), .ZN(y[202]) );
  OR2_X1 U142bar ( .A1(abar[12]), .A2(bbar[10]), .ZN(ybar[202]);
  AND2_X1 U143 ( .A1(a[12]), .A2(b[9]), .ZN(y[201]) );
  OR2_X1 U143bar ( .A1(abar[12]), .A2(bbar[9]), .ZN(ybar[201]);
  AND2_X1 U144 ( .A1(a[12]), .A2(b[8]), .ZN(y[200]) );
  OR2_X1 U144bar ( .A1(abar[12]), .A2(bbar[8]), .ZN(ybar[200]);
  AND2_X1 U145 ( .A1(b[1]), .A2(a[0]), .ZN(y[1]) );
  OR2_X1 U145bar ( .A1(bbar[1]), .A2(abar[0]), .ZN(ybar[1]);
  AND2_X1 U146 ( .A1(a[1]), .A2(b[3]), .ZN(y[19]) );
  OR2_X1 U146bar ( .A1(abar[1]), .A2(bbar[3]), .ZN(ybar[19]);
  AND2_X1 U147 ( .A1(a[12]), .A2(b[7]), .ZN(y[199]) );
  OR2_X1 U147bar ( .A1(abar[12]), .A2(bbar[7]), .ZN(ybar[199]);
  AND2_X1 U148 ( .A1(a[12]), .A2(b[6]), .ZN(y[198]) );
  OR2_X1 U148bar ( .A1(abar[12]), .A2(bbar[6]), .ZN(ybar[198]);
  AND2_X1 U149 ( .A1(a[12]), .A2(b[5]), .ZN(y[197]) );
  OR2_X1 U149bar ( .A1(abar[12]), .A2(bbar[5]), .ZN(ybar[197]);
  AND2_X1 U150 ( .A1(a[12]), .A2(b[4]), .ZN(y[196]) );
  OR2_X1 U150bar ( .A1(abar[12]), .A2(bbar[4]), .ZN(ybar[196]);
  AND2_X1 U151 ( .A1(a[12]), .A2(b[3]), .ZN(y[195]) );
  OR2_X1 U151bar ( .A1(abar[12]), .A2(bbar[3]), .ZN(ybar[195]);
  AND2_X1 U152 ( .A1(a[12]), .A2(b[2]), .ZN(y[194]) );
  OR2_X1 U152bar ( .A1(abar[12]), .A2(bbar[2]), .ZN(ybar[194]);
  AND2_X1 U153 ( .A1(a[12]), .A2(b[1]), .ZN(y[193]) );
  OR2_X1 U153bar ( .A1(abar[12]), .A2(bbar[1]), .ZN(ybar[193]);
  AND2_X1 U154 ( .A1(a[12]), .A2(b[0]), .ZN(y[192]) );
  OR2_X1 U154bar ( .A1(abar[12]), .A2(bbar[0]), .ZN(ybar[192]);
  AND2_X1 U155 ( .A1(a[11]), .A2(b[15]), .ZN(y[191]) );
  OR2_X1 U155bar ( .A1(abar[11]), .A2(bbar[15]), .ZN(ybar[191]);
  AND2_X1 U156 ( .A1(a[11]), .A2(b[14]), .ZN(y[190]) );
  OR2_X1 U156bar ( .A1(abar[11]), .A2(bbar[14]), .ZN(ybar[190]);
  AND2_X1 U157 ( .A1(a[1]), .A2(b[2]), .ZN(y[18]) );
  OR2_X1 U157bar ( .A1(abar[1]), .A2(bbar[2]), .ZN(ybar[18]);
  AND2_X1 U158 ( .A1(a[11]), .A2(b[13]), .ZN(y[189]) );
  OR2_X1 U158bar ( .A1(abar[11]), .A2(bbar[13]), .ZN(ybar[189]);
  AND2_X1 U159 ( .A1(a[11]), .A2(b[12]), .ZN(y[188]) );
  OR2_X1 U159bar ( .A1(abar[11]), .A2(bbar[12]), .ZN(ybar[188]);
  AND2_X1 U160 ( .A1(a[11]), .A2(b[11]), .ZN(y[187]) );
  OR2_X1 U160bar ( .A1(abar[11]), .A2(bbar[11]), .ZN(ybar[187]);
  AND2_X1 U161 ( .A1(a[11]), .A2(b[10]), .ZN(y[186]) );
  OR2_X1 U161bar ( .A1(abar[11]), .A2(bbar[10]), .ZN(ybar[186]);
  AND2_X1 U162 ( .A1(a[11]), .A2(b[9]), .ZN(y[185]) );
  OR2_X1 U162bar ( .A1(abar[11]), .A2(bbar[9]), .ZN(ybar[185]);
  AND2_X1 U163 ( .A1(a[11]), .A2(b[8]), .ZN(y[184]) );
  OR2_X1 U163bar ( .A1(abar[11]), .A2(bbar[8]), .ZN(ybar[184]);
  AND2_X1 U164 ( .A1(a[11]), .A2(b[7]), .ZN(y[183]) );
  OR2_X1 U164bar ( .A1(abar[11]), .A2(bbar[7]), .ZN(ybar[183]);
  AND2_X1 U165 ( .A1(a[11]), .A2(b[6]), .ZN(y[182]) );
  OR2_X1 U165bar ( .A1(abar[11]), .A2(bbar[6]), .ZN(ybar[182]);
  AND2_X1 U166 ( .A1(a[11]), .A2(b[5]), .ZN(y[181]) );
  OR2_X1 U166bar ( .A1(abar[11]), .A2(bbar[5]), .ZN(ybar[181]);
  AND2_X1 U167 ( .A1(a[11]), .A2(b[4]), .ZN(y[180]) );
  OR2_X1 U167bar ( .A1(abar[11]), .A2(bbar[4]), .ZN(ybar[180]);
  AND2_X1 U168 ( .A1(a[1]), .A2(b[1]), .ZN(y[17]) );
  OR2_X1 U168bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[17]);
  AND2_X1 U169 ( .A1(a[11]), .A2(b[3]), .ZN(y[179]) );
  OR2_X1 U169bar ( .A1(abar[11]), .A2(bbar[3]), .ZN(ybar[179]);
  AND2_X1 U170 ( .A1(a[11]), .A2(b[2]), .ZN(y[178]) );
  OR2_X1 U170bar ( .A1(abar[11]), .A2(bbar[2]), .ZN(ybar[178]);
  AND2_X1 U171 ( .A1(a[11]), .A2(b[1]), .ZN(y[177]) );
  OR2_X1 U171bar ( .A1(abar[11]), .A2(bbar[1]), .ZN(ybar[177]);
  AND2_X1 U172 ( .A1(a[11]), .A2(b[0]), .ZN(y[176]) );
  OR2_X1 U172bar ( .A1(abar[11]), .A2(bbar[0]), .ZN(ybar[176]);
  AND2_X1 U173 ( .A1(a[10]), .A2(b[15]), .ZN(y[175]) );
  OR2_X1 U173bar ( .A1(abar[10]), .A2(bbar[15]), .ZN(ybar[175]);
  AND2_X1 U174 ( .A1(a[10]), .A2(b[14]), .ZN(y[174]) );
  OR2_X1 U174bar ( .A1(abar[10]), .A2(bbar[14]), .ZN(ybar[174]);
  AND2_X1 U175 ( .A1(a[10]), .A2(b[13]), .ZN(y[173]) );
  OR2_X1 U175bar ( .A1(abar[10]), .A2(bbar[13]), .ZN(ybar[173]);
  AND2_X1 U176 ( .A1(a[10]), .A2(b[12]), .ZN(y[172]) );
  OR2_X1 U176bar ( .A1(abar[10]), .A2(bbar[12]), .ZN(ybar[172]);
  AND2_X1 U177 ( .A1(a[10]), .A2(b[11]), .ZN(y[171]) );
  OR2_X1 U177bar ( .A1(abar[10]), .A2(bbar[11]), .ZN(ybar[171]);
  AND2_X1 U178 ( .A1(a[10]), .A2(b[10]), .ZN(y[170]) );
  OR2_X1 U178bar ( .A1(abar[10]), .A2(bbar[10]), .ZN(ybar[170]);
  AND2_X1 U179 ( .A1(a[1]), .A2(b[0]), .ZN(y[16]) );
  OR2_X1 U179bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[16]);
  AND2_X1 U180 ( .A1(a[10]), .A2(b[9]), .ZN(y[169]) );
  OR2_X1 U180bar ( .A1(abar[10]), .A2(bbar[9]), .ZN(ybar[169]);
  AND2_X1 U181 ( .A1(a[10]), .A2(b[8]), .ZN(y[168]) );
  OR2_X1 U181bar ( .A1(abar[10]), .A2(bbar[8]), .ZN(ybar[168]);
  AND2_X1 U182 ( .A1(a[10]), .A2(b[7]), .ZN(y[167]) );
  OR2_X1 U182bar ( .A1(abar[10]), .A2(bbar[7]), .ZN(ybar[167]);
  AND2_X1 U183 ( .A1(a[10]), .A2(b[6]), .ZN(y[166]) );
  OR2_X1 U183bar ( .A1(abar[10]), .A2(bbar[6]), .ZN(ybar[166]);
  AND2_X1 U184 ( .A1(a[10]), .A2(b[5]), .ZN(y[165]) );
  OR2_X1 U184bar ( .A1(abar[10]), .A2(bbar[5]), .ZN(ybar[165]);
  AND2_X1 U185 ( .A1(a[10]), .A2(b[4]), .ZN(y[164]) );
  OR2_X1 U185bar ( .A1(abar[10]), .A2(bbar[4]), .ZN(ybar[164]);
  AND2_X1 U186 ( .A1(a[10]), .A2(b[3]), .ZN(y[163]) );
  OR2_X1 U186bar ( .A1(abar[10]), .A2(bbar[3]), .ZN(ybar[163]);
  AND2_X1 U187 ( .A1(a[10]), .A2(b[2]), .ZN(y[162]) );
  OR2_X1 U187bar ( .A1(abar[10]), .A2(bbar[2]), .ZN(ybar[162]);
  AND2_X1 U188 ( .A1(a[10]), .A2(b[1]), .ZN(y[161]) );
  OR2_X1 U188bar ( .A1(abar[10]), .A2(bbar[1]), .ZN(ybar[161]);
  AND2_X1 U189 ( .A1(a[10]), .A2(b[0]), .ZN(y[160]) );
  OR2_X1 U189bar ( .A1(abar[10]), .A2(bbar[0]), .ZN(ybar[160]);
  AND2_X1 U190 ( .A1(b[15]), .A2(a[0]), .ZN(y[15]) );
  OR2_X1 U190bar ( .A1(bbar[15]), .A2(abar[0]), .ZN(ybar[15]);
  AND2_X1 U191 ( .A1(a[9]), .A2(b[15]), .ZN(y[159]) );
  OR2_X1 U191bar ( .A1(abar[9]), .A2(bbar[15]), .ZN(ybar[159]);
  AND2_X1 U192 ( .A1(a[9]), .A2(b[14]), .ZN(y[158]) );
  OR2_X1 U192bar ( .A1(abar[9]), .A2(bbar[14]), .ZN(ybar[158]);
  AND2_X1 U193 ( .A1(a[9]), .A2(b[13]), .ZN(y[157]) );
  OR2_X1 U193bar ( .A1(abar[9]), .A2(bbar[13]), .ZN(ybar[157]);
  AND2_X1 U194 ( .A1(a[9]), .A2(b[12]), .ZN(y[156]) );
  OR2_X1 U194bar ( .A1(abar[9]), .A2(bbar[12]), .ZN(ybar[156]);
  AND2_X1 U195 ( .A1(a[9]), .A2(b[11]), .ZN(y[155]) );
  OR2_X1 U195bar ( .A1(abar[9]), .A2(bbar[11]), .ZN(ybar[155]);
  AND2_X1 U196 ( .A1(a[9]), .A2(b[10]), .ZN(y[154]) );
  OR2_X1 U196bar ( .A1(abar[9]), .A2(bbar[10]), .ZN(ybar[154]);
  AND2_X1 U197 ( .A1(a[9]), .A2(b[9]), .ZN(y[153]) );
  OR2_X1 U197bar ( .A1(abar[9]), .A2(bbar[9]), .ZN(ybar[153]);
  AND2_X1 U198 ( .A1(a[9]), .A2(b[8]), .ZN(y[152]) );
  OR2_X1 U198bar ( .A1(abar[9]), .A2(bbar[8]), .ZN(ybar[152]);
  AND2_X1 U199 ( .A1(a[9]), .A2(b[7]), .ZN(y[151]) );
  OR2_X1 U199bar ( .A1(abar[9]), .A2(bbar[7]), .ZN(ybar[151]);
  AND2_X1 U200 ( .A1(a[9]), .A2(b[6]), .ZN(y[150]) );
  OR2_X1 U200bar ( .A1(abar[9]), .A2(bbar[6]), .ZN(ybar[150]);
  AND2_X1 U201 ( .A1(b[14]), .A2(a[0]), .ZN(y[14]) );
  OR2_X1 U201bar ( .A1(bbar[14]), .A2(abar[0]), .ZN(ybar[14]);
  AND2_X1 U202 ( .A1(a[9]), .A2(b[5]), .ZN(y[149]) );
  OR2_X1 U202bar ( .A1(abar[9]), .A2(bbar[5]), .ZN(ybar[149]);
  AND2_X1 U203 ( .A1(a[9]), .A2(b[4]), .ZN(y[148]) );
  OR2_X1 U203bar ( .A1(abar[9]), .A2(bbar[4]), .ZN(ybar[148]);
  AND2_X1 U204 ( .A1(a[9]), .A2(b[3]), .ZN(y[147]) );
  OR2_X1 U204bar ( .A1(abar[9]), .A2(bbar[3]), .ZN(ybar[147]);
  AND2_X1 U205 ( .A1(a[9]), .A2(b[2]), .ZN(y[146]) );
  OR2_X1 U205bar ( .A1(abar[9]), .A2(bbar[2]), .ZN(ybar[146]);
  AND2_X1 U206 ( .A1(a[9]), .A2(b[1]), .ZN(y[145]) );
  OR2_X1 U206bar ( .A1(abar[9]), .A2(bbar[1]), .ZN(ybar[145]);
  AND2_X1 U207 ( .A1(a[9]), .A2(b[0]), .ZN(y[144]) );
  OR2_X1 U207bar ( .A1(abar[9]), .A2(bbar[0]), .ZN(ybar[144]);
  AND2_X1 U208 ( .A1(a[8]), .A2(b[15]), .ZN(y[143]) );
  OR2_X1 U208bar ( .A1(abar[8]), .A2(bbar[15]), .ZN(ybar[143]);
  AND2_X1 U209 ( .A1(a[8]), .A2(b[14]), .ZN(y[142]) );
  OR2_X1 U209bar ( .A1(abar[8]), .A2(bbar[14]), .ZN(ybar[142]);
  AND2_X1 U210 ( .A1(a[8]), .A2(b[13]), .ZN(y[141]) );
  OR2_X1 U210bar ( .A1(abar[8]), .A2(bbar[13]), .ZN(ybar[141]);
  AND2_X1 U211 ( .A1(a[8]), .A2(b[12]), .ZN(y[140]) );
  OR2_X1 U211bar ( .A1(abar[8]), .A2(bbar[12]), .ZN(ybar[140]);
  AND2_X1 U212 ( .A1(b[13]), .A2(a[0]), .ZN(y[13]) );
  OR2_X1 U212bar ( .A1(bbar[13]), .A2(abar[0]), .ZN(ybar[13]);
  AND2_X1 U213 ( .A1(a[8]), .A2(b[11]), .ZN(y[139]) );
  OR2_X1 U213bar ( .A1(abar[8]), .A2(bbar[11]), .ZN(ybar[139]);
  AND2_X1 U214 ( .A1(a[8]), .A2(b[10]), .ZN(y[138]) );
  OR2_X1 U214bar ( .A1(abar[8]), .A2(bbar[10]), .ZN(ybar[138]);
  AND2_X1 U215 ( .A1(a[8]), .A2(b[9]), .ZN(y[137]) );
  OR2_X1 U215bar ( .A1(abar[8]), .A2(bbar[9]), .ZN(ybar[137]);
  AND2_X1 U216 ( .A1(a[8]), .A2(b[8]), .ZN(y[136]) );
  OR2_X1 U216bar ( .A1(abar[8]), .A2(bbar[8]), .ZN(ybar[136]);
  AND2_X1 U217 ( .A1(a[8]), .A2(b[7]), .ZN(y[135]) );
  OR2_X1 U217bar ( .A1(abar[8]), .A2(bbar[7]), .ZN(ybar[135]);
  AND2_X1 U218 ( .A1(a[8]), .A2(b[6]), .ZN(y[134]) );
  OR2_X1 U218bar ( .A1(abar[8]), .A2(bbar[6]), .ZN(ybar[134]);
  AND2_X1 U219 ( .A1(a[8]), .A2(b[5]), .ZN(y[133]) );
  OR2_X1 U219bar ( .A1(abar[8]), .A2(bbar[5]), .ZN(ybar[133]);
  AND2_X1 U220 ( .A1(a[8]), .A2(b[4]), .ZN(y[132]) );
  OR2_X1 U220bar ( .A1(abar[8]), .A2(bbar[4]), .ZN(ybar[132]);
  AND2_X1 U221 ( .A1(a[8]), .A2(b[3]), .ZN(y[131]) );
  OR2_X1 U221bar ( .A1(abar[8]), .A2(bbar[3]), .ZN(ybar[131]);
  AND2_X1 U222 ( .A1(a[8]), .A2(b[2]), .ZN(y[130]) );
  OR2_X1 U222bar ( .A1(abar[8]), .A2(bbar[2]), .ZN(ybar[130]);
  AND2_X1 U223 ( .A1(b[12]), .A2(a[0]), .ZN(y[12]) );
  OR2_X1 U223bar ( .A1(bbar[12]), .A2(abar[0]), .ZN(ybar[12]);
  AND2_X1 U224 ( .A1(a[8]), .A2(b[1]), .ZN(y[129]) );
  OR2_X1 U224bar ( .A1(abar[8]), .A2(bbar[1]), .ZN(ybar[129]);
  AND2_X1 U225 ( .A1(a[8]), .A2(b[0]), .ZN(y[128]) );
  OR2_X1 U225bar ( .A1(abar[8]), .A2(bbar[0]), .ZN(ybar[128]);
  AND2_X1 U226 ( .A1(a[7]), .A2(b[15]), .ZN(y[127]) );
  OR2_X1 U226bar ( .A1(abar[7]), .A2(bbar[15]), .ZN(ybar[127]);
  AND2_X1 U227 ( .A1(a[7]), .A2(b[14]), .ZN(y[126]) );
  OR2_X1 U227bar ( .A1(abar[7]), .A2(bbar[14]), .ZN(ybar[126]);
  AND2_X1 U228 ( .A1(a[7]), .A2(b[13]), .ZN(y[125]) );
  OR2_X1 U228bar ( .A1(abar[7]), .A2(bbar[13]), .ZN(ybar[125]);
  AND2_X1 U229 ( .A1(a[7]), .A2(b[12]), .ZN(y[124]) );
  OR2_X1 U229bar ( .A1(abar[7]), .A2(bbar[12]), .ZN(ybar[124]);
  AND2_X1 U230 ( .A1(a[7]), .A2(b[11]), .ZN(y[123]) );
  OR2_X1 U230bar ( .A1(abar[7]), .A2(bbar[11]), .ZN(ybar[123]);
  AND2_X1 U231 ( .A1(a[7]), .A2(b[10]), .ZN(y[122]) );
  OR2_X1 U231bar ( .A1(abar[7]), .A2(bbar[10]), .ZN(ybar[122]);
  AND2_X1 U232 ( .A1(a[7]), .A2(b[9]), .ZN(y[121]) );
  OR2_X1 U232bar ( .A1(abar[7]), .A2(bbar[9]), .ZN(ybar[121]);
  AND2_X1 U233 ( .A1(a[7]), .A2(b[8]), .ZN(y[120]) );
  OR2_X1 U233bar ( .A1(abar[7]), .A2(bbar[8]), .ZN(ybar[120]);
  AND2_X1 U234 ( .A1(b[11]), .A2(a[0]), .ZN(y[11]) );
  OR2_X1 U234bar ( .A1(bbar[11]), .A2(abar[0]), .ZN(ybar[11]);
  AND2_X1 U235 ( .A1(a[7]), .A2(b[7]), .ZN(y[119]) );
  OR2_X1 U235bar ( .A1(abar[7]), .A2(bbar[7]), .ZN(ybar[119]);
  AND2_X1 U236 ( .A1(a[7]), .A2(b[6]), .ZN(y[118]) );
  OR2_X1 U236bar ( .A1(abar[7]), .A2(bbar[6]), .ZN(ybar[118]);
  AND2_X1 U237 ( .A1(a[7]), .A2(b[5]), .ZN(y[117]) );
  OR2_X1 U237bar ( .A1(abar[7]), .A2(bbar[5]), .ZN(ybar[117]);
  AND2_X1 U238 ( .A1(a[7]), .A2(b[4]), .ZN(y[116]) );
  OR2_X1 U238bar ( .A1(abar[7]), .A2(bbar[4]), .ZN(ybar[116]);
  AND2_X1 U239 ( .A1(a[7]), .A2(b[3]), .ZN(y[115]) );
  OR2_X1 U239bar ( .A1(abar[7]), .A2(bbar[3]), .ZN(ybar[115]);
  AND2_X1 U240 ( .A1(a[7]), .A2(b[2]), .ZN(y[114]) );
  OR2_X1 U240bar ( .A1(abar[7]), .A2(bbar[2]), .ZN(ybar[114]);
  AND2_X1 U241 ( .A1(a[7]), .A2(b[1]), .ZN(y[113]) );
  OR2_X1 U241bar ( .A1(abar[7]), .A2(bbar[1]), .ZN(ybar[113]);
  AND2_X1 U242 ( .A1(a[7]), .A2(b[0]), .ZN(y[112]) );
  OR2_X1 U242bar ( .A1(abar[7]), .A2(bbar[0]), .ZN(ybar[112]);
  AND2_X1 U243 ( .A1(b[15]), .A2(a[6]), .ZN(y[111]) );
  OR2_X1 U243bar ( .A1(bbar[15]), .A2(abar[6]), .ZN(ybar[111]);
  AND2_X1 U244 ( .A1(b[14]), .A2(a[6]), .ZN(y[110]) );
  OR2_X1 U244bar ( .A1(bbar[14]), .A2(abar[6]), .ZN(ybar[110]);
  AND2_X1 U245 ( .A1(b[10]), .A2(a[0]), .ZN(y[10]) );
  OR2_X1 U245bar ( .A1(bbar[10]), .A2(abar[0]), .ZN(ybar[10]);
  AND2_X1 U246 ( .A1(b[13]), .A2(a[6]), .ZN(y[109]) );
  OR2_X1 U246bar ( .A1(bbar[13]), .A2(abar[6]), .ZN(ybar[109]);
  AND2_X1 U247 ( .A1(b[12]), .A2(a[6]), .ZN(y[108]) );
  OR2_X1 U247bar ( .A1(bbar[12]), .A2(abar[6]), .ZN(ybar[108]);
  AND2_X1 U248 ( .A1(b[11]), .A2(a[6]), .ZN(y[107]) );
  OR2_X1 U248bar ( .A1(bbar[11]), .A2(abar[6]), .ZN(ybar[107]);
  AND2_X1 U249 ( .A1(b[10]), .A2(a[6]), .ZN(y[106]) );
  OR2_X1 U249bar ( .A1(bbar[10]), .A2(abar[6]), .ZN(ybar[106]);
  AND2_X1 U250 ( .A1(a[6]), .A2(b[9]), .ZN(y[105]) );
  OR2_X1 U250bar ( .A1(abar[6]), .A2(bbar[9]), .ZN(ybar[105]);
  AND2_X1 U251 ( .A1(b[8]), .A2(a[6]), .ZN(y[104]) );
  OR2_X1 U251bar ( .A1(bbar[8]), .A2(abar[6]), .ZN(ybar[104]);
  AND2_X1 U252 ( .A1(b[7]), .A2(a[6]), .ZN(y[103]) );
  OR2_X1 U252bar ( .A1(bbar[7]), .A2(abar[6]), .ZN(ybar[103]);
  AND2_X1 U253 ( .A1(b[6]), .A2(a[6]), .ZN(y[102]) );
  OR2_X1 U253bar ( .A1(bbar[6]), .A2(abar[6]), .ZN(ybar[102]);
  AND2_X1 U254 ( .A1(b[5]), .A2(a[6]), .ZN(y[101]) );
  OR2_X1 U254bar ( .A1(bbar[5]), .A2(abar[6]), .ZN(ybar[101]);
  AND2_X1 U255 ( .A1(b[4]), .A2(a[6]), .ZN(y[100]) );
  OR2_X1 U255bar ( .A1(bbar[4]), .A2(abar[6]), .ZN(ybar[100]);
  AND2_X1 U256 ( .A1(b[0]), .A2(a[0]), .ZN(y[0]) );
  OR2_X1 U256bar ( .A1(bbar[0]), .A2(abar[0]), .ZN(ybar[0]);
endmodule




module decode_18 ( in, out );
  input [7:0] in;
  //input_done

  output [255:0] out;
  //output_done

  wire   [15:0] level1;
  wire   [31:0] level2;
  //wire_done

  CD2_72 cd_l1_1 ( .a(in[1]), .b(in[0]), .y(level1[3:0]) );
  CD2_71 cd_l1_2 ( .a(in[3]), .b(in[2]), .y(level1[7:4]) );
  CD2_70 cd_l1_3 ( .a(in[5]), .b(in[4]), .y(level1[11:8]) );
  CD2_69 cd_l1_4 ( .a(in[7]), .b(in[6]), .y(level1[15:12]) );
  CD4_36 cd_l2_1 ( .a(level1[7:4]), .b(level1[3:0]), .y(level2[15:0]) );
  CD4_35 cd_l2_2 ( .a(level1[15:12]), .b(level1[11:8]), .y(level2[31:16]) );
  CD16_18 cd_l3 ( .a(level2[31:16]), .b(level2[15:0]), .y(out) );
endmodule


module encode_18 ( in, out );
  input [255:0] in;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
  assign inbar[8] = ~in[8];
  assign inbar[9] = ~in[9];
  assign inbar[10] = ~in[10];
  assign inbar[11] = ~in[11];
  assign inbar[12] = ~in[12];
  assign inbar[13] = ~in[13];
  assign inbar[14] = ~in[14];
  assign inbar[15] = ~in[15];
  assign inbar[16] = ~in[16];
  assign inbar[17] = ~in[17];
  assign inbar[18] = ~in[18];
  assign inbar[19] = ~in[19];
  assign inbar[20] = ~in[20];
  assign inbar[21] = ~in[21];
  assign inbar[22] = ~in[22];
  assign inbar[23] = ~in[23];
  assign inbar[24] = ~in[24];
  assign inbar[25] = ~in[25];
  assign inbar[26] = ~in[26];
  assign inbar[27] = ~in[27];
  assign inbar[28] = ~in[28];
  assign inbar[29] = ~in[29];
  assign inbar[30] = ~in[30];
  assign inbar[31] = ~in[31];
  assign inbar[32] = ~in[32];
  assign inbar[33] = ~in[33];
  assign inbar[34] = ~in[34];
  assign inbar[35] = ~in[35];
  assign inbar[36] = ~in[36];
  assign inbar[37] = ~in[37];
  assign inbar[38] = ~in[38];
  assign inbar[39] = ~in[39];
  assign inbar[40] = ~in[40];
  assign inbar[41] = ~in[41];
  assign inbar[42] = ~in[42];
  assign inbar[43] = ~in[43];
  assign inbar[44] = ~in[44];
  assign inbar[45] = ~in[45];
  assign inbar[46] = ~in[46];
  assign inbar[47] = ~in[47];
  assign inbar[48] = ~in[48];
  assign inbar[49] = ~in[49];
  assign inbar[50] = ~in[50];
  assign inbar[51] = ~in[51];
  assign inbar[52] = ~in[52];
  assign inbar[53] = ~in[53];
  assign inbar[54] = ~in[54];
  assign inbar[55] = ~in[55];
  assign inbar[56] = ~in[56];
  assign inbar[57] = ~in[57];
  assign inbar[58] = ~in[58];
  assign inbar[59] = ~in[59];
  assign inbar[60] = ~in[60];
  assign inbar[61] = ~in[61];
  assign inbar[62] = ~in[62];
  assign inbar[63] = ~in[63];
  assign inbar[64] = ~in[64];
  assign inbar[65] = ~in[65];
  assign inbar[66] = ~in[66];
  assign inbar[67] = ~in[67];
  assign inbar[68] = ~in[68];
  assign inbar[69] = ~in[69];
  assign inbar[70] = ~in[70];
  assign inbar[71] = ~in[71];
  assign inbar[72] = ~in[72];
  assign inbar[73] = ~in[73];
  assign inbar[74] = ~in[74];
  assign inbar[75] = ~in[75];
  assign inbar[76] = ~in[76];
  assign inbar[77] = ~in[77];
  assign inbar[78] = ~in[78];
  assign inbar[79] = ~in[79];
  assign inbar[80] = ~in[80];
  assign inbar[81] = ~in[81];
  assign inbar[82] = ~in[82];
  assign inbar[83] = ~in[83];
  assign inbar[84] = ~in[84];
  assign inbar[85] = ~in[85];
  assign inbar[86] = ~in[86];
  assign inbar[87] = ~in[87];
  assign inbar[88] = ~in[88];
  assign inbar[89] = ~in[89];
  assign inbar[90] = ~in[90];
  assign inbar[91] = ~in[91];
  assign inbar[92] = ~in[92];
  assign inbar[93] = ~in[93];
  assign inbar[94] = ~in[94];
  assign inbar[95] = ~in[95];
  assign inbar[96] = ~in[96];
  assign inbar[97] = ~in[97];
  assign inbar[98] = ~in[98];
  assign inbar[99] = ~in[99];
  assign inbar[100] = ~in[100];
  assign inbar[101] = ~in[101];
  assign inbar[102] = ~in[102];
  assign inbar[103] = ~in[103];
  assign inbar[104] = ~in[104];
  assign inbar[105] = ~in[105];
  assign inbar[106] = ~in[106];
  assign inbar[107] = ~in[107];
  assign inbar[108] = ~in[108];
  assign inbar[109] = ~in[109];
  assign inbar[110] = ~in[110];
  assign inbar[111] = ~in[111];
  assign inbar[112] = ~in[112];
  assign inbar[113] = ~in[113];
  assign inbar[114] = ~in[114];
  assign inbar[115] = ~in[115];
  assign inbar[116] = ~in[116];
  assign inbar[117] = ~in[117];
  assign inbar[118] = ~in[118];
  assign inbar[119] = ~in[119];
  assign inbar[120] = ~in[120];
  assign inbar[121] = ~in[121];
  assign inbar[122] = ~in[122];
  assign inbar[123] = ~in[123];
  assign inbar[124] = ~in[124];
  assign inbar[125] = ~in[125];
  assign inbar[126] = ~in[126];
  assign inbar[127] = ~in[127];
  assign inbar[128] = ~in[128];
  assign inbar[129] = ~in[129];
  assign inbar[130] = ~in[130];
  assign inbar[131] = ~in[131];
  assign inbar[132] = ~in[132];
  assign inbar[133] = ~in[133];
  assign inbar[134] = ~in[134];
  assign inbar[135] = ~in[135];
  assign inbar[136] = ~in[136];
  assign inbar[137] = ~in[137];
  assign inbar[138] = ~in[138];
  assign inbar[139] = ~in[139];
  assign inbar[140] = ~in[140];
  assign inbar[141] = ~in[141];
  assign inbar[142] = ~in[142];
  assign inbar[143] = ~in[143];
  assign inbar[144] = ~in[144];
  assign inbar[145] = ~in[145];
  assign inbar[146] = ~in[146];
  assign inbar[147] = ~in[147];
  assign inbar[148] = ~in[148];
  assign inbar[149] = ~in[149];
  assign inbar[150] = ~in[150];
  assign inbar[151] = ~in[151];
  assign inbar[152] = ~in[152];
  assign inbar[153] = ~in[153];
  assign inbar[154] = ~in[154];
  assign inbar[155] = ~in[155];
  assign inbar[156] = ~in[156];
  assign inbar[157] = ~in[157];
  assign inbar[158] = ~in[158];
  assign inbar[159] = ~in[159];
  assign inbar[160] = ~in[160];
  assign inbar[161] = ~in[161];
  assign inbar[162] = ~in[162];
  assign inbar[163] = ~in[163];
  assign inbar[164] = ~in[164];
  assign inbar[165] = ~in[165];
  assign inbar[166] = ~in[166];
  assign inbar[167] = ~in[167];
  assign inbar[168] = ~in[168];
  assign inbar[169] = ~in[169];
  assign inbar[170] = ~in[170];
  assign inbar[171] = ~in[171];
  assign inbar[172] = ~in[172];
  assign inbar[173] = ~in[173];
  assign inbar[174] = ~in[174];
  assign inbar[175] = ~in[175];
  assign inbar[176] = ~in[176];
  assign inbar[177] = ~in[177];
  assign inbar[178] = ~in[178];
  assign inbar[179] = ~in[179];
  assign inbar[180] = ~in[180];
  assign inbar[181] = ~in[181];
  assign inbar[182] = ~in[182];
  assign inbar[183] = ~in[183];
  assign inbar[184] = ~in[184];
  assign inbar[185] = ~in[185];
  assign inbar[186] = ~in[186];
  assign inbar[187] = ~in[187];
  assign inbar[188] = ~in[188];
  assign inbar[189] = ~in[189];
  assign inbar[190] = ~in[190];
  assign inbar[191] = ~in[191];
  assign inbar[192] = ~in[192];
  assign inbar[193] = ~in[193];
  assign inbar[194] = ~in[194];
  assign inbar[195] = ~in[195];
  assign inbar[196] = ~in[196];
  assign inbar[197] = ~in[197];
  assign inbar[198] = ~in[198];
  assign inbar[199] = ~in[199];
  assign inbar[200] = ~in[200];
  assign inbar[201] = ~in[201];
  assign inbar[202] = ~in[202];
  assign inbar[203] = ~in[203];
  assign inbar[204] = ~in[204];
  assign inbar[205] = ~in[205];
  assign inbar[206] = ~in[206];
  assign inbar[207] = ~in[207];
  assign inbar[208] = ~in[208];
  assign inbar[209] = ~in[209];
  assign inbar[210] = ~in[210];
  assign inbar[211] = ~in[211];
  assign inbar[212] = ~in[212];
  assign inbar[213] = ~in[213];
  assign inbar[214] = ~in[214];
  assign inbar[215] = ~in[215];
  assign inbar[216] = ~in[216];
  assign inbar[217] = ~in[217];
  assign inbar[218] = ~in[218];
  assign inbar[219] = ~in[219];
  assign inbar[220] = ~in[220];
  assign inbar[221] = ~in[221];
  assign inbar[222] = ~in[222];
  assign inbar[223] = ~in[223];
  assign inbar[224] = ~in[224];
  assign inbar[225] = ~in[225];
  assign inbar[226] = ~in[226];
  assign inbar[227] = ~in[227];
  assign inbar[228] = ~in[228];
  assign inbar[229] = ~in[229];
  assign inbar[230] = ~in[230];
  assign inbar[231] = ~in[231];
  assign inbar[232] = ~in[232];
  assign inbar[233] = ~in[233];
  assign inbar[234] = ~in[234];
  assign inbar[235] = ~in[235];
  assign inbar[236] = ~in[236];
  assign inbar[237] = ~in[237];
  assign inbar[238] = ~in[238];
  assign inbar[239] = ~in[239];
  assign inbar[240] = ~in[240];
  assign inbar[241] = ~in[241];
  assign inbar[242] = ~in[242];
  assign inbar[243] = ~in[243];
  assign inbar[244] = ~in[244];
  assign inbar[245] = ~in[245];
  assign inbar[246] = ~in[246];
  assign inbar[247] = ~in[247];
  assign inbar[248] = ~in[248];
  assign inbar[249] = ~in[249];
  assign inbar[250] = ~in[250];
  assign inbar[251] = ~in[251];
  assign inbar[252] = ~in[252];
  assign inbar[253] = ~in[253];
  assign inbar[254] = ~in[254];
  assign inbar[255] = ~in[255];
  //input_done

  output [7:0] out;
  reg [7:0] outbar;
  //output_done

  wire   in_81, in_80, in_79, in_78, in_77, in_76, in_75, in_74, in_73, in_72,
         in_71, in_70, in_69, in_68, in_67, in_66, in_65, in_64, in_63, in_62,
         in_61, in_60, in_59, in_58, in_57, in_56, in_55, in_54, in_53, in_52,
         in_51, in_50, in_49, in_48, in_47, in_46, in_45, in_44, in_43, in_42,
         in_41, in_40, in_39, in_38, in_37, in_36, in_35, in_34, in_33, in_32,
         in_31, in_30, in_29, in_28, in_27, in_26, in_25, in_24, in_23, in_22,
         in_21, in_20, in_19, in_18, in_17, in_16, in_15, in_14, in_13, in_12,
         in_11, in_10, in_9, in_8, in_7, in_6, in_5, in_4, in_3, in_2, in_1,
         in_0, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972;
  wire in_81bar, in_80bar, in_79bar, in_78bar, in_77bar, in_76bar, in_75bar, in_74bar, in_73bar, in_72bar, in_71bar, in_70bar, in_69bar, in_68bar, in_67bar, in_66bar, in_65bar, in_64bar, in_63bar, in_62bar, in_61bar, in_60bar, in_59bar, in_58bar, in_57bar, in_56bar, in_55bar, in_54bar, in_53bar, in_52bar, in_51bar, in_50bar, in_49bar, in_48bar, in_47bar, in_46bar, in_45bar, in_44bar, in_43bar, in_42bar, in_41bar, in_40bar, in_39bar, in_38bar, in_37bar, in_36bar, in_35bar, in_34bar, in_33bar, in_32bar, in_31bar, in_30bar, in_29bar, in_28bar, in_27bar, in_26bar, in_25bar, in_24bar, in_23bar, in_22bar, in_21bar, in_20bar, in_19bar, in_18bar, in_17bar, in_16bar, in_15bar, in_14bar, in_13bar, in_12bar, in_11bar, in_10bar, in_9bar, in_8bar, in_7bar, in_6bar, in_5bar, in_4bar, in_3bar, in_2bar, in_1bar, in_0bar, n487bar, n488bar, n489bar, n490bar, n491bar, n492bar, n493bar, n494bar, n495bar, n496bar, n497bar, n498bar, n499bar, n500bar, n501bar, n502bar, n503bar, n504bar, n505bar, n506bar, n507bar, n508bar, n509bar, n510bar, n511bar, n512bar, n513bar, n514bar, n515bar, n516bar, n517bar, n518bar, n519bar, n520bar, n521bar, n522bar, n523bar, n524bar, n525bar, n526bar, n527bar, n528bar, n529bar, n530bar, n531bar, n532bar, n533bar, n534bar, n535bar, n536bar, n537bar, n538bar, n539bar, n540bar, n541bar, n542bar, n543bar, n544bar, n545bar, n546bar, n547bar, n548bar, n549bar, n550bar, n551bar, n552bar, n553bar, n554bar, n555bar, n556bar, n557bar, n558bar, n559bar, n560bar, n561bar, n562bar, n563bar, n564bar, n565bar, n566bar, n567bar, n568bar, n569bar, n570bar, n571bar, n572bar, n573bar, n574bar, n575bar, n576bar, n577bar, n578bar, n579bar, n580bar, n581bar, n582bar, n583bar, n584bar, n585bar, n586bar, n587bar, n588bar, n589bar, n590bar, n591bar, n592bar, n593bar, n594bar, n595bar, n596bar, n597bar, n598bar, n599bar, n600bar, n601bar, n602bar, n603bar, n604bar, n605bar, n606bar, n607bar, n608bar, n609bar, n610bar, n611bar, n612bar, n613bar, n614bar, n615bar, n616bar, n617bar, n618bar, n619bar, n620bar, n621bar, n622bar, n623bar, n624bar, n625bar, n626bar, n627bar, n628bar, n629bar, n630bar, n631bar, n632bar, n633bar, n634bar, n635bar, n636bar, n637bar, n638bar, n639bar, n640bar, n641bar, n642bar, n643bar, n644bar, n645bar, n646bar, n647bar, n648bar, n649bar, n650bar, n651bar, n652bar, n653bar, n654bar, n655bar, n656bar, n657bar, n658bar, n659bar, n660bar, n661bar, n662bar, n663bar, n664bar, n665bar, n666bar, n667bar, n668bar, n669bar, n670bar, n671bar, n672bar, n673bar, n674bar, n675bar, n676bar, n677bar, n678bar, n679bar, n680bar, n681bar, n682bar, n683bar, n684bar, n685bar, n686bar, n687bar, n688bar, n689bar, n690bar, n691bar, n692bar, n693bar, n694bar, n695bar, n696bar, n697bar, n698bar, n699bar, n700bar, n701bar, n702bar, n703bar, n704bar, n705bar, n706bar, n707bar, n708bar, n709bar, n710bar, n711bar, n712bar, n713bar, n714bar, n715bar, n716bar, n717bar, n718bar, n719bar, n720bar, n721bar, n722bar, n723bar, n724bar, n725bar, n726bar, n727bar, n728bar, n729bar, n730bar, n731bar, n732bar, n733bar, n734bar, n735bar, n736bar, n737bar, n738bar, n739bar, n740bar, n741bar, n742bar, n743bar, n744bar, n745bar, n746bar, n747bar, n748bar, n749bar, n750bar, n751bar, n752bar, n753bar, n754bar, n755bar, n756bar, n757bar, n758bar, n759bar, n760bar, n761bar, n762bar, n763bar, n764bar, n765bar, n766bar, n767bar, n768bar, n769bar, n770bar, n771bar, n772bar, n773bar, n774bar, n775bar, n776bar, n777bar, n778bar, n779bar, n780bar, n781bar, n782bar, n783bar, n784bar, n785bar, n786bar, n787bar, n788bar, n789bar, n790bar, n791bar, n792bar, n793bar, n794bar, n795bar, n796bar, n797bar, n798bar, n799bar, n800bar, n801bar, n802bar, n803bar, n804bar, n805bar, n806bar, n807bar, n808bar, n809bar, n810bar, n811bar, n812bar, n813bar, n814bar, n815bar, n816bar, n817bar, n818bar, n819bar, n820bar, n821bar, n822bar, n823bar, n824bar, n825bar, n826bar, n827bar, n828bar, n829bar, n830bar, n831bar, n832bar, n833bar, n834bar, n835bar, n836bar, n837bar, n838bar, n839bar, n840bar, n841bar, n842bar, n843bar, n844bar, n845bar, n846bar, n847bar, n848bar, n849bar, n850bar, n851bar, n852bar, n853bar, n854bar, n855bar, n856bar, n857bar, n858bar, n859bar, n860bar, n861bar, n862bar, n863bar, n864bar, n865bar, n866bar, n867bar, n868bar, n869bar, n870bar, n871bar, n872bar, n873bar, n874bar, n875bar, n876bar, n877bar, n878bar, n879bar, n880bar, n881bar, n882bar, n883bar, n884bar, n885bar, n886bar, n887bar, n888bar, n889bar, n890bar, n891bar, n892bar, n893bar, n894bar, n895bar, n896bar, n897bar, n898bar, n899bar, n900bar, n901bar, n902bar, n903bar, n904bar, n905bar, n906bar, n907bar, n908bar, n909bar, n910bar, n911bar, n912bar, n913bar, n914bar, n915bar, n916bar, n917bar, n918bar, n919bar, n920bar, n921bar, n922bar, n923bar, n924bar, n925bar, n926bar, n927bar, n928bar, n929bar, n930bar, n931bar, n932bar, n933bar, n934bar, n935bar, n936bar, n937bar, n938bar, n939bar, n940bar, n941bar, n942bar, n943bar, n944bar, n945bar, n946bar, n947bar, n948bar, n949bar, n950bar, n951bar, n952bar, n953bar, n954bar, n955bar, n956bar, n957bar, n958bar, n959bar, n960bar, n961bar, n962bar, n963bar, n964bar, n965bar, n966bar, n967bar, n968bar, n969bar, n970bar, n971bar, n972bar;
  //wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];

  OR2_X1 U1 ( .A1(n972), .A2(n971), .ZN(out[7]) );
  AND2_X1 U1bar ( .A1(n972bar), .A2(n971bar), .ZN(outbar[7]);
  OR2_X1 U2 ( .A1(n970), .A2(n969), .ZN(n971) );
  AND2_X1 U2bar ( .A1(n970bar), .A2(n969bar), .ZN(n971bar);
  OR2_X1 U3 ( .A1(n968), .A2(n967), .ZN(n969) );
  AND2_X1 U3bar ( .A1(n968bar), .A2(n967bar), .ZN(n969bar);
  OR2_X1 U4 ( .A1(n966), .A2(n965), .ZN(n967) );
  AND2_X1 U4bar ( .A1(n966bar), .A2(n965bar), .ZN(n967bar);
  OR2_X1 U5 ( .A1(n964), .A2(n963), .ZN(n968) );
  AND2_X1 U5bar ( .A1(n964bar), .A2(n963bar), .ZN(n968bar);
  OR2_X1 U6 ( .A1(in[116]), .A2(n962), .ZN(n963) );
  AND2_X1 U6bar ( .A1(inbar[116]), .A2(n962bar), .ZN(n963bar);
  OR2_X1 U7 ( .A1(n961), .A2(n960), .ZN(n970) );
  AND2_X1 U7bar ( .A1(n961bar), .A2(n960bar), .ZN(n970bar);
  OR2_X1 U8 ( .A1(in[150]), .A2(in[127]), .ZN(n960) );
  AND2_X1 U8bar ( .A1(inbar[150]), .A2(inbar[127]), .ZN(n960bar);
  OR2_X1 U9 ( .A1(in[160]), .A2(n959), .ZN(n961) );
  AND2_X1 U9bar ( .A1(inbar[160]), .A2(n959bar), .ZN(n961bar);
  OR2_X1 U10 ( .A1(in[252]), .A2(in[168]), .ZN(n959) );
  AND2_X1 U10bar ( .A1(inbar[252]), .A2(inbar[168]), .ZN(n959bar);
  OR2_X1 U11 ( .A1(n958), .A2(n957), .ZN(n972) );
  AND2_X1 U11bar ( .A1(n958bar), .A2(n957bar), .ZN(n972bar);
  OR2_X1 U12 ( .A1(n956), .A2(n955), .ZN(n957) );
  AND2_X1 U12bar ( .A1(n956bar), .A2(n955bar), .ZN(n957bar);
  OR2_X1 U13 ( .A1(in_17), .A2(in[96]), .ZN(n955) );
  AND2_X1 U13bar ( .A1(in_17bar), .A2(inbar[96]), .ZN(n955bar);
  OR2_X1 U14 ( .A1(in_23), .A2(n954), .ZN(n956) );
  AND2_X1 U14bar ( .A1(in_23bar), .A2(n954bar), .ZN(n956bar);
  OR2_X1 U15 ( .A1(in_31), .A2(in_26), .ZN(n954) );
  AND2_X1 U15bar ( .A1(in_31bar), .A2(in_26bar), .ZN(n954bar);
  OR2_X1 U16 ( .A1(n953), .A2(n952), .ZN(n958) );
  AND2_X1 U16bar ( .A1(n953bar), .A2(n952bar), .ZN(n958bar);
  OR2_X1 U17 ( .A1(in_58), .A2(in_4), .ZN(n952) );
  AND2_X1 U17bar ( .A1(in_58bar), .A2(in_4bar), .ZN(n952bar);
  OR2_X1 U18 ( .A1(in_59), .A2(n951), .ZN(n953) );
  AND2_X1 U18bar ( .A1(in_59bar), .A2(n951bar), .ZN(n953bar);
  OR2_X1 U19 ( .A1(in_71), .A2(in_62), .ZN(n951) );
  AND2_X1 U19bar ( .A1(in_71bar), .A2(in_62bar), .ZN(n951bar);
  OR2_X1 U20 ( .A1(n950), .A2(n949), .ZN(out[6]) );
  AND2_X1 U20bar ( .A1(n950bar), .A2(n949bar), .ZN(outbar[6]);
  OR2_X1 U21 ( .A1(n948), .A2(n947), .ZN(n949) );
  AND2_X1 U21bar ( .A1(n948bar), .A2(n947bar), .ZN(n949bar);
  OR2_X1 U22 ( .A1(n946), .A2(n945), .ZN(n947) );
  AND2_X1 U22bar ( .A1(n946bar), .A2(n945bar), .ZN(n947bar);
  OR2_X1 U23 ( .A1(n944), .A2(n943), .ZN(n945) );
  AND2_X1 U23bar ( .A1(n944bar), .A2(n943bar), .ZN(n945bar);
  OR2_X1 U24 ( .A1(n942), .A2(n941), .ZN(n946) );
  AND2_X1 U24bar ( .A1(n942bar), .A2(n941bar), .ZN(n946bar);
  OR2_X1 U25 ( .A1(in[101]), .A2(n940), .ZN(n941) );
  AND2_X1 U25bar ( .A1(inbar[101]), .A2(n940bar), .ZN(n941bar);
  OR2_X1 U26 ( .A1(n939), .A2(n938), .ZN(n948) );
  AND2_X1 U26bar ( .A1(n939bar), .A2(n938bar), .ZN(n948bar);
  OR2_X1 U27 ( .A1(in[114]), .A2(in[104]), .ZN(n938) );
  AND2_X1 U27bar ( .A1(inbar[114]), .A2(inbar[104]), .ZN(n938bar);
  OR2_X1 U28 ( .A1(in[128]), .A2(n937), .ZN(n939) );
  AND2_X1 U28bar ( .A1(inbar[128]), .A2(n937bar), .ZN(n939bar);
  OR2_X1 U29 ( .A1(in[136]), .A2(in[134]), .ZN(n937) );
  AND2_X1 U29bar ( .A1(inbar[136]), .A2(inbar[134]), .ZN(n937bar);
  OR2_X1 U30 ( .A1(n936), .A2(n935), .ZN(n950) );
  AND2_X1 U30bar ( .A1(n936bar), .A2(n935bar), .ZN(n950bar);
  OR2_X1 U31 ( .A1(n934), .A2(n933), .ZN(n935) );
  AND2_X1 U31bar ( .A1(n934bar), .A2(n933bar), .ZN(n935bar);
  OR2_X1 U32 ( .A1(in[177]), .A2(in[164]), .ZN(n933) );
  AND2_X1 U32bar ( .A1(inbar[177]), .A2(inbar[164]), .ZN(n933bar);
  OR2_X1 U33 ( .A1(in[212]), .A2(n932), .ZN(n934) );
  AND2_X1 U33bar ( .A1(inbar[212]), .A2(n932bar), .ZN(n934bar);
  OR2_X1 U34 ( .A1(in[248]), .A2(in[221]), .ZN(n932) );
  AND2_X1 U34bar ( .A1(inbar[248]), .A2(inbar[221]), .ZN(n932bar);
  OR2_X1 U35 ( .A1(n931), .A2(n930), .ZN(n936) );
  AND2_X1 U35bar ( .A1(n931bar), .A2(n930bar), .ZN(n936bar);
  OR2_X1 U36 ( .A1(in_18), .A2(in[93]), .ZN(n930) );
  AND2_X1 U36bar ( .A1(in_18bar), .A2(inbar[93]), .ZN(n930bar);
  OR2_X1 U37 ( .A1(in_31), .A2(n929), .ZN(n931) );
  AND2_X1 U37bar ( .A1(in_31bar), .A2(n929bar), .ZN(n931bar);
  OR2_X1 U38 ( .A1(in_7), .A2(in_39), .ZN(n929) );
  AND2_X1 U38bar ( .A1(in_7bar), .A2(in_39bar), .ZN(n929bar);
  OR2_X1 U39 ( .A1(n928), .A2(n927), .ZN(out[5]) );
  AND2_X1 U39bar ( .A1(n928bar), .A2(n927bar), .ZN(outbar[5]);
  OR2_X1 U40 ( .A1(n926), .A2(n925), .ZN(n927) );
  AND2_X1 U40bar ( .A1(n926bar), .A2(n925bar), .ZN(n927bar);
  OR2_X1 U41 ( .A1(n924), .A2(n923), .ZN(n925) );
  AND2_X1 U41bar ( .A1(n924bar), .A2(n923bar), .ZN(n925bar);
  OR2_X1 U42 ( .A1(n922), .A2(n921), .ZN(n923) );
  AND2_X1 U42bar ( .A1(n922bar), .A2(n921bar), .ZN(n923bar);
  OR2_X1 U43 ( .A1(n940), .A2(n920), .ZN(n924) );
  AND2_X1 U43bar ( .A1(n940bar), .A2(n920bar), .ZN(n924bar);
  OR2_X1 U44 ( .A1(in[111]), .A2(n919), .ZN(n920) );
  AND2_X1 U44bar ( .A1(inbar[111]), .A2(n919bar), .ZN(n920bar);
  OR2_X1 U45 ( .A1(n918), .A2(n917), .ZN(n940) );
  AND2_X1 U45bar ( .A1(n918bar), .A2(n917bar), .ZN(n940bar);
  OR2_X1 U46 ( .A1(n916), .A2(n915), .ZN(n917) );
  AND2_X1 U46bar ( .A1(n916bar), .A2(n915bar), .ZN(n917bar);
  OR2_X1 U47 ( .A1(n914), .A2(n913), .ZN(n915) );
  AND2_X1 U47bar ( .A1(n914bar), .A2(n913bar), .ZN(n915bar);
  OR2_X1 U48 ( .A1(in[140]), .A2(in[131]), .ZN(n913) );
  AND2_X1 U48bar ( .A1(inbar[140]), .A2(inbar[131]), .ZN(n913bar);
  OR2_X1 U49 ( .A1(in[160]), .A2(in[144]), .ZN(n914) );
  AND2_X1 U49bar ( .A1(inbar[160]), .A2(inbar[144]), .ZN(n914bar);
  OR2_X1 U50 ( .A1(n912), .A2(n911), .ZN(n916) );
  AND2_X1 U50bar ( .A1(n912bar), .A2(n911bar), .ZN(n916bar);
  OR2_X1 U51 ( .A1(in[179]), .A2(in[174]), .ZN(n911) );
  AND2_X1 U51bar ( .A1(inbar[179]), .A2(inbar[174]), .ZN(n911bar);
  OR2_X1 U52 ( .A1(in[188]), .A2(in[184]), .ZN(n912) );
  AND2_X1 U52bar ( .A1(inbar[188]), .A2(inbar[184]), .ZN(n912bar);
  OR2_X1 U53 ( .A1(n910), .A2(n909), .ZN(n918) );
  AND2_X1 U53bar ( .A1(n910bar), .A2(n909bar), .ZN(n918bar);
  OR2_X1 U54 ( .A1(n908), .A2(n907), .ZN(n909) );
  AND2_X1 U54bar ( .A1(n908bar), .A2(n907bar), .ZN(n909bar);
  OR2_X1 U55 ( .A1(in[216]), .A2(in[200]), .ZN(n907) );
  AND2_X1 U55bar ( .A1(inbar[216]), .A2(inbar[200]), .ZN(n907bar);
  OR2_X1 U56 ( .A1(in[228]), .A2(in[224]), .ZN(n908) );
  AND2_X1 U56bar ( .A1(inbar[228]), .A2(inbar[224]), .ZN(n908bar);
  OR2_X1 U57 ( .A1(n906), .A2(n905), .ZN(n910) );
  AND2_X1 U57bar ( .A1(n906bar), .A2(n905bar), .ZN(n910bar);
  OR2_X1 U58 ( .A1(in[247]), .A2(in[235]), .ZN(n905) );
  AND2_X1 U58bar ( .A1(inbar[247]), .A2(inbar[235]), .ZN(n905bar);
  OR2_X1 U59 ( .A1(in_42), .A2(in[83]), .ZN(n906) );
  AND2_X1 U59bar ( .A1(in_42bar), .A2(inbar[83]), .ZN(n906bar);
  OR2_X1 U60 ( .A1(n904), .A2(n903), .ZN(n926) );
  AND2_X1 U60bar ( .A1(n904bar), .A2(n903bar), .ZN(n926bar);
  OR2_X1 U61 ( .A1(in[166]), .A2(in[123]), .ZN(n903) );
  AND2_X1 U61bar ( .A1(inbar[166]), .A2(inbar[123]), .ZN(n903bar);
  OR2_X1 U62 ( .A1(in[170]), .A2(n902), .ZN(n904) );
  AND2_X1 U62bar ( .A1(inbar[170]), .A2(n902bar), .ZN(n904bar);
  OR2_X1 U63 ( .A1(in[194]), .A2(in[183]), .ZN(n902) );
  AND2_X1 U63bar ( .A1(inbar[194]), .A2(inbar[183]), .ZN(n902bar);
  OR2_X1 U64 ( .A1(n901), .A2(n900), .ZN(n928) );
  AND2_X1 U64bar ( .A1(n901bar), .A2(n900bar), .ZN(n928bar);
  OR2_X1 U65 ( .A1(n899), .A2(n898), .ZN(n900) );
  AND2_X1 U65bar ( .A1(n899bar), .A2(n898bar), .ZN(n900bar);
  OR2_X1 U66 ( .A1(in[241]), .A2(in[238]), .ZN(n898) );
  AND2_X1 U66bar ( .A1(inbar[241]), .A2(inbar[238]), .ZN(n898bar);
  OR2_X1 U67 ( .A1(in[250]), .A2(n897), .ZN(n899) );
  AND2_X1 U67bar ( .A1(inbar[250]), .A2(n897bar), .ZN(n899bar);
  OR2_X1 U68 ( .A1(in_24), .A2(in[84]), .ZN(n897) );
  AND2_X1 U68bar ( .A1(in_24bar), .A2(inbar[84]), .ZN(n897bar);
  OR2_X1 U69 ( .A1(n896), .A2(n895), .ZN(n901) );
  AND2_X1 U69bar ( .A1(n896bar), .A2(n895bar), .ZN(n901bar);
  OR2_X1 U70 ( .A1(in_41), .A2(in_29), .ZN(n895) );
  AND2_X1 U70bar ( .A1(in_41bar), .A2(in_29bar), .ZN(n895bar);
  OR2_X1 U71 ( .A1(in_66), .A2(n894), .ZN(n896) );
  AND2_X1 U71bar ( .A1(in_66bar), .A2(n894bar), .ZN(n896bar);
  OR2_X1 U72 ( .A1(in_76), .A2(in_71), .ZN(n894) );
  AND2_X1 U72bar ( .A1(in_76bar), .A2(in_71bar), .ZN(n894bar);
  OR2_X1 U73 ( .A1(n893), .A2(n892), .ZN(out[4]) );
  AND2_X1 U73bar ( .A1(n893bar), .A2(n892bar), .ZN(outbar[4]);
  OR2_X1 U74 ( .A1(n891), .A2(n890), .ZN(n892) );
  AND2_X1 U74bar ( .A1(n891bar), .A2(n890bar), .ZN(n892bar);
  OR2_X1 U75 ( .A1(n889), .A2(n888), .ZN(n890) );
  AND2_X1 U75bar ( .A1(n889bar), .A2(n888bar), .ZN(n890bar);
  OR2_X1 U76 ( .A1(n922), .A2(n887), .ZN(n888) );
  AND2_X1 U76bar ( .A1(n922bar), .A2(n887bar), .ZN(n888bar);
  OR2_X1 U77 ( .A1(n886), .A2(n885), .ZN(n922) );
  AND2_X1 U77bar ( .A1(n886bar), .A2(n885bar), .ZN(n922bar);
  OR2_X1 U78 ( .A1(n884), .A2(n883), .ZN(n885) );
  AND2_X1 U78bar ( .A1(n884bar), .A2(n883bar), .ZN(n885bar);
  OR2_X1 U79 ( .A1(n882), .A2(n881), .ZN(n883) );
  AND2_X1 U79bar ( .A1(n882bar), .A2(n881bar), .ZN(n883bar);
  OR2_X1 U80 ( .A1(in[118]), .A2(in[109]), .ZN(n881) );
  AND2_X1 U80bar ( .A1(inbar[118]), .A2(inbar[109]), .ZN(n881bar);
  OR2_X1 U81 ( .A1(in[139]), .A2(in[120]), .ZN(n882) );
  AND2_X1 U81bar ( .A1(inbar[139]), .A2(inbar[120]), .ZN(n882bar);
  OR2_X1 U82 ( .A1(n880), .A2(n879), .ZN(n884) );
  AND2_X1 U82bar ( .A1(n880bar), .A2(n879bar), .ZN(n884bar);
  OR2_X1 U83 ( .A1(in[198]), .A2(in[154]), .ZN(n879) );
  AND2_X1 U83bar ( .A1(inbar[198]), .A2(inbar[154]), .ZN(n879bar);
  OR2_X1 U84 ( .A1(in[210]), .A2(in[205]), .ZN(n880) );
  AND2_X1 U84bar ( .A1(inbar[210]), .A2(inbar[205]), .ZN(n880bar);
  OR2_X1 U85 ( .A1(n878), .A2(n877), .ZN(n886) );
  AND2_X1 U85bar ( .A1(n878bar), .A2(n877bar), .ZN(n886bar);
  OR2_X1 U86 ( .A1(n876), .A2(n875), .ZN(n877) );
  AND2_X1 U86bar ( .A1(n876bar), .A2(n875bar), .ZN(n877bar);
  OR2_X1 U87 ( .A1(in[219]), .A2(in[217]), .ZN(n875) );
  AND2_X1 U87bar ( .A1(inbar[219]), .A2(inbar[217]), .ZN(n875bar);
  OR2_X1 U88 ( .A1(in[86]), .A2(in[252]), .ZN(n876) );
  AND2_X1 U88bar ( .A1(inbar[86]), .A2(inbar[252]), .ZN(n876bar);
  OR2_X1 U89 ( .A1(n874), .A2(n873), .ZN(n878) );
  AND2_X1 U89bar ( .A1(n874bar), .A2(n873bar), .ZN(n878bar);
  OR2_X1 U90 ( .A1(in_40), .A2(in[91]), .ZN(n873) );
  AND2_X1 U90bar ( .A1(in_40bar), .A2(inbar[91]), .ZN(n873bar);
  OR2_X1 U91 ( .A1(in_8), .A2(in_46), .ZN(n874) );
  AND2_X1 U91bar ( .A1(in_8bar), .A2(in_46bar), .ZN(n874bar);
  OR2_X1 U92 ( .A1(n872), .A2(n871), .ZN(n889) );
  AND2_X1 U92bar ( .A1(n872bar), .A2(n871bar), .ZN(n889bar);
  OR2_X1 U93 ( .A1(in[117]), .A2(n943), .ZN(n871) );
  AND2_X1 U93bar ( .A1(inbar[117]), .A2(n943bar), .ZN(n871bar);
  OR2_X1 U94 ( .A1(n870), .A2(n869), .ZN(n943) );
  AND2_X1 U94bar ( .A1(n870bar), .A2(n869bar), .ZN(n943bar);
  OR2_X1 U95 ( .A1(n868), .A2(n867), .ZN(n869) );
  AND2_X1 U95bar ( .A1(n868bar), .A2(n867bar), .ZN(n869bar);
  OR2_X1 U96 ( .A1(n866), .A2(n865), .ZN(n867) );
  AND2_X1 U96bar ( .A1(n866bar), .A2(n865bar), .ZN(n867bar);
  OR2_X1 U97 ( .A1(n864), .A2(n863), .ZN(n865) );
  AND2_X1 U97bar ( .A1(n864bar), .A2(n863bar), .ZN(n865bar);
  OR2_X1 U98 ( .A1(in[108]), .A2(n919), .ZN(n866) );
  AND2_X1 U98bar ( .A1(inbar[108]), .A2(n919bar), .ZN(n866bar);
  OR2_X1 U99 ( .A1(n862), .A2(n861), .ZN(n919) );
  AND2_X1 U99bar ( .A1(n862bar), .A2(n861bar), .ZN(n919bar);
  OR2_X1 U100 ( .A1(n860), .A2(n859), .ZN(n861) );
  AND2_X1 U100bar ( .A1(n860bar), .A2(n859bar), .ZN(n861bar);
  OR2_X1 U101 ( .A1(n858), .A2(n857), .ZN(n859) );
  AND2_X1 U101bar ( .A1(n858bar), .A2(n857bar), .ZN(n859bar);
  OR2_X1 U102 ( .A1(in[119]), .A2(in[105]), .ZN(n857) );
  AND2_X1 U102bar ( .A1(inbar[119]), .A2(inbar[105]), .ZN(n857bar);
  OR2_X1 U103 ( .A1(in[186]), .A2(in[175]), .ZN(n858) );
  AND2_X1 U103bar ( .A1(inbar[186]), .A2(inbar[175]), .ZN(n858bar);
  OR2_X1 U104 ( .A1(n856), .A2(n855), .ZN(n860) );
  AND2_X1 U104bar ( .A1(n856bar), .A2(n855bar), .ZN(n860bar);
  OR2_X1 U105 ( .A1(in[202]), .A2(in[193]), .ZN(n855) );
  AND2_X1 U105bar ( .A1(inbar[202]), .A2(inbar[193]), .ZN(n855bar);
  OR2_X1 U106 ( .A1(in[225]), .A2(in[208]), .ZN(n856) );
  AND2_X1 U106bar ( .A1(inbar[225]), .A2(inbar[208]), .ZN(n856bar);
  OR2_X1 U107 ( .A1(n854), .A2(n853), .ZN(n862) );
  AND2_X1 U107bar ( .A1(n854bar), .A2(n853bar), .ZN(n862bar);
  OR2_X1 U108 ( .A1(n852), .A2(n851), .ZN(n853) );
  AND2_X1 U108bar ( .A1(n852bar), .A2(n851bar), .ZN(n853bar);
  OR2_X1 U109 ( .A1(in_1), .A2(in[85]), .ZN(n851) );
  AND2_X1 U109bar ( .A1(in_1bar), .A2(inbar[85]), .ZN(n851bar);
  OR2_X1 U110 ( .A1(in_23), .A2(in_19), .ZN(n852) );
  AND2_X1 U110bar ( .A1(in_23bar), .A2(in_19bar), .ZN(n852bar);
  OR2_X1 U111 ( .A1(n850), .A2(n849), .ZN(n854) );
  AND2_X1 U111bar ( .A1(n850bar), .A2(n849bar), .ZN(n854bar);
  OR2_X1 U112 ( .A1(in_43), .A2(in_33), .ZN(n849) );
  AND2_X1 U112bar ( .A1(in_43bar), .A2(in_33bar), .ZN(n849bar);
  OR2_X1 U113 ( .A1(in_63), .A2(in_44), .ZN(n850) );
  AND2_X1 U113bar ( .A1(in_63bar), .A2(in_44bar), .ZN(n850bar);
  OR2_X1 U114 ( .A1(n848), .A2(n847), .ZN(n868) );
  AND2_X1 U114bar ( .A1(n848bar), .A2(n847bar), .ZN(n868bar);
  OR2_X1 U115 ( .A1(in[141]), .A2(in[112]), .ZN(n847) );
  AND2_X1 U115bar ( .A1(inbar[141]), .A2(inbar[112]), .ZN(n847bar);
  OR2_X1 U116 ( .A1(in[147]), .A2(n846), .ZN(n848) );
  AND2_X1 U116bar ( .A1(inbar[147]), .A2(n846bar), .ZN(n848bar);
  OR2_X1 U117 ( .A1(in[181]), .A2(in[167]), .ZN(n846) );
  AND2_X1 U117bar ( .A1(inbar[181]), .A2(inbar[167]), .ZN(n846bar);
  OR2_X1 U118 ( .A1(n845), .A2(n844), .ZN(n870) );
  AND2_X1 U118bar ( .A1(n845bar), .A2(n844bar), .ZN(n870bar);
  OR2_X1 U119 ( .A1(n843), .A2(n842), .ZN(n844) );
  AND2_X1 U119bar ( .A1(n843bar), .A2(n842bar), .ZN(n844bar);
  OR2_X1 U120 ( .A1(in[229]), .A2(in[201]), .ZN(n842) );
  AND2_X1 U120bar ( .A1(inbar[229]), .A2(inbar[201]), .ZN(n842bar);
  OR2_X1 U121 ( .A1(in[237]), .A2(n841), .ZN(n843) );
  AND2_X1 U121bar ( .A1(inbar[237]), .A2(n841bar), .ZN(n843bar);
  OR2_X1 U122 ( .A1(in[94]), .A2(in[253]), .ZN(n841) );
  AND2_X1 U122bar ( .A1(inbar[94]), .A2(inbar[253]), .ZN(n841bar);
  OR2_X1 U123 ( .A1(n840), .A2(n839), .ZN(n845) );
  AND2_X1 U123bar ( .A1(n840bar), .A2(n839bar), .ZN(n845bar);
  OR2_X1 U124 ( .A1(in_21), .A2(in[96]), .ZN(n839) );
  AND2_X1 U124bar ( .A1(in_21bar), .A2(inbar[96]), .ZN(n839bar);
  OR2_X1 U125 ( .A1(in_25), .A2(n838), .ZN(n840) );
  AND2_X1 U125bar ( .A1(in_25bar), .A2(n838bar), .ZN(n840bar);
  OR2_X1 U126 ( .A1(in_81), .A2(in_45), .ZN(n838) );
  AND2_X1 U126bar ( .A1(in_81bar), .A2(in_45bar), .ZN(n838bar);
  OR2_X1 U127 ( .A1(n837), .A2(n836), .ZN(n891) );
  AND2_X1 U127bar ( .A1(n837bar), .A2(n836bar), .ZN(n891bar);
  OR2_X1 U128 ( .A1(in[142]), .A2(in[124]), .ZN(n836) );
  AND2_X1 U128bar ( .A1(inbar[142]), .A2(inbar[124]), .ZN(n836bar);
  OR2_X1 U129 ( .A1(in[150]), .A2(n835), .ZN(n837) );
  AND2_X1 U129bar ( .A1(inbar[150]), .A2(n835bar), .ZN(n837bar);
  OR2_X1 U130 ( .A1(in[172]), .A2(in[155]), .ZN(n835) );
  AND2_X1 U130bar ( .A1(inbar[172]), .A2(inbar[155]), .ZN(n835bar);
  OR2_X1 U131 ( .A1(n834), .A2(n833), .ZN(n893) );
  AND2_X1 U131bar ( .A1(n834bar), .A2(n833bar), .ZN(n893bar);
  OR2_X1 U132 ( .A1(n832), .A2(n831), .ZN(n833) );
  AND2_X1 U132bar ( .A1(n832bar), .A2(n831bar), .ZN(n833bar);
  OR2_X1 U133 ( .A1(in[196]), .A2(in[173]), .ZN(n831) );
  AND2_X1 U133bar ( .A1(inbar[196]), .A2(inbar[173]), .ZN(n831bar);
  OR2_X1 U134 ( .A1(in[222]), .A2(n830), .ZN(n832) );
  AND2_X1 U134bar ( .A1(inbar[222]), .A2(n830bar), .ZN(n832bar);
  OR2_X1 U135 ( .A1(in[227]), .A2(in[226]), .ZN(n830) );
  AND2_X1 U135bar ( .A1(inbar[227]), .A2(inbar[226]), .ZN(n830bar);
  OR2_X1 U136 ( .A1(n829), .A2(n828), .ZN(n834) );
  AND2_X1 U136bar ( .A1(n829bar), .A2(n828bar), .ZN(n834bar);
  OR2_X1 U137 ( .A1(in[249]), .A2(in[231]), .ZN(n828) );
  AND2_X1 U137bar ( .A1(inbar[249]), .A2(inbar[231]), .ZN(n828bar);
  OR2_X1 U138 ( .A1(in_28), .A2(n827), .ZN(n829) );
  AND2_X1 U138bar ( .A1(in_28bar), .A2(n827bar), .ZN(n829bar);
  OR2_X1 U139 ( .A1(in_52), .A2(in_47), .ZN(n827) );
  AND2_X1 U139bar ( .A1(in_52bar), .A2(in_47bar), .ZN(n827bar);
  OR2_X1 U140 ( .A1(n826), .A2(n825), .ZN(out[3]) );
  AND2_X1 U140bar ( .A1(n826bar), .A2(n825bar), .ZN(outbar[3]);
  OR2_X1 U141 ( .A1(n824), .A2(n823), .ZN(n825) );
  AND2_X1 U141bar ( .A1(n824bar), .A2(n823bar), .ZN(n825bar);
  OR2_X1 U142 ( .A1(n822), .A2(n821), .ZN(n823) );
  AND2_X1 U142bar ( .A1(n822bar), .A2(n821bar), .ZN(n823bar);
  OR2_X1 U143 ( .A1(n820), .A2(n819), .ZN(n821) );
  AND2_X1 U143bar ( .A1(n820bar), .A2(n819bar), .ZN(n821bar);
  OR2_X1 U144 ( .A1(n964), .A2(n818), .ZN(n822) );
  AND2_X1 U144bar ( .A1(n964bar), .A2(n818bar), .ZN(n822bar);
  OR2_X1 U145 ( .A1(in[118]), .A2(n817), .ZN(n818) );
  AND2_X1 U145bar ( .A1(inbar[118]), .A2(n817bar), .ZN(n818bar);
  OR2_X1 U146 ( .A1(n816), .A2(n815), .ZN(n964) );
  AND2_X1 U146bar ( .A1(n816bar), .A2(n815bar), .ZN(n964bar);
  OR2_X1 U147 ( .A1(n814), .A2(n813), .ZN(n815) );
  AND2_X1 U147bar ( .A1(n814bar), .A2(n813bar), .ZN(n815bar);
  OR2_X1 U148 ( .A1(n812), .A2(n811), .ZN(n813) );
  AND2_X1 U148bar ( .A1(n812bar), .A2(n811bar), .ZN(n813bar);
  OR2_X1 U149 ( .A1(in[122]), .A2(in[111]), .ZN(n811) );
  AND2_X1 U149bar ( .A1(inbar[122]), .A2(inbar[111]), .ZN(n811bar);
  OR2_X1 U150 ( .A1(in[154]), .A2(in[151]), .ZN(n812) );
  AND2_X1 U150bar ( .A1(inbar[154]), .A2(inbar[151]), .ZN(n812bar);
  OR2_X1 U151 ( .A1(n810), .A2(n809), .ZN(n814) );
  AND2_X1 U151bar ( .A1(n810bar), .A2(n809bar), .ZN(n814bar);
  OR2_X1 U152 ( .A1(in[187]), .A2(in[177]), .ZN(n809) );
  AND2_X1 U152bar ( .A1(inbar[187]), .A2(inbar[177]), .ZN(n809bar);
  OR2_X1 U153 ( .A1(in[200]), .A2(in[192]), .ZN(n810) );
  AND2_X1 U153bar ( .A1(inbar[200]), .A2(inbar[192]), .ZN(n810bar);
  OR2_X1 U154 ( .A1(n808), .A2(n807), .ZN(n816) );
  AND2_X1 U154bar ( .A1(n808bar), .A2(n807bar), .ZN(n816bar);
  OR2_X1 U155 ( .A1(n806), .A2(n805), .ZN(n807) );
  AND2_X1 U155bar ( .A1(n806bar), .A2(n805bar), .ZN(n807bar);
  OR2_X1 U156 ( .A1(in[225]), .A2(in[207]), .ZN(n805) );
  AND2_X1 U156bar ( .A1(inbar[225]), .A2(inbar[207]), .ZN(n805bar);
  OR2_X1 U157 ( .A1(in[98]), .A2(in[226]), .ZN(n806) );
  AND2_X1 U157bar ( .A1(inbar[98]), .A2(inbar[226]), .ZN(n806bar);
  OR2_X1 U158 ( .A1(n804), .A2(n803), .ZN(n808) );
  AND2_X1 U158bar ( .A1(n804bar), .A2(n803bar), .ZN(n808bar);
  OR2_X1 U159 ( .A1(in_20), .A2(in_16), .ZN(n803) );
  AND2_X1 U159bar ( .A1(in_20bar), .A2(in_16bar), .ZN(n803bar);
  OR2_X1 U160 ( .A1(in_55), .A2(in_45), .ZN(n804) );
  AND2_X1 U160bar ( .A1(in_55bar), .A2(in_45bar), .ZN(n804bar);
  OR2_X1 U161 ( .A1(n802), .A2(n801), .ZN(n824) );
  AND2_X1 U161bar ( .A1(n802bar), .A2(n801bar), .ZN(n824bar);
  OR2_X1 U162 ( .A1(in[162]), .A2(in[149]), .ZN(n801) );
  AND2_X1 U162bar ( .A1(inbar[162]), .A2(inbar[149]), .ZN(n801bar);
  OR2_X1 U163 ( .A1(in[163]), .A2(n800), .ZN(n802) );
  AND2_X1 U163bar ( .A1(inbar[163]), .A2(n800bar), .ZN(n802bar);
  OR2_X1 U164 ( .A1(in[191]), .A2(in[189]), .ZN(n800) );
  AND2_X1 U164bar ( .A1(inbar[191]), .A2(inbar[189]), .ZN(n800bar);
  OR2_X1 U165 ( .A1(n799), .A2(n798), .ZN(n826) );
  AND2_X1 U165bar ( .A1(n799bar), .A2(n798bar), .ZN(n826bar);
  OR2_X1 U166 ( .A1(n797), .A2(n796), .ZN(n798) );
  AND2_X1 U166bar ( .A1(n797bar), .A2(n796bar), .ZN(n798bar);
  OR2_X1 U167 ( .A1(in[212]), .A2(in[193]), .ZN(n796) );
  AND2_X1 U167bar ( .A1(inbar[212]), .A2(inbar[193]), .ZN(n796bar);
  OR2_X1 U168 ( .A1(in[238]), .A2(n795), .ZN(n797) );
  AND2_X1 U168bar ( .A1(inbar[238]), .A2(n795bar), .ZN(n797bar);
  OR2_X1 U169 ( .A1(in[88]), .A2(in[247]), .ZN(n795) );
  AND2_X1 U169bar ( .A1(inbar[88]), .A2(inbar[247]), .ZN(n795bar);
  OR2_X1 U170 ( .A1(n794), .A2(n793), .ZN(n799) );
  AND2_X1 U170bar ( .A1(n794bar), .A2(n793bar), .ZN(n799bar);
  OR2_X1 U171 ( .A1(in[94]), .A2(in[92]), .ZN(n793) );
  AND2_X1 U171bar ( .A1(inbar[94]), .A2(inbar[92]), .ZN(n793bar);
  OR2_X1 U172 ( .A1(in_52), .A2(n792), .ZN(n794) );
  AND2_X1 U172bar ( .A1(in_52bar), .A2(n792bar), .ZN(n794bar);
  OR2_X1 U173 ( .A1(in_70), .A2(in_67), .ZN(n792) );
  AND2_X1 U173bar ( .A1(in_70bar), .A2(in_67bar), .ZN(n792bar);
  OR2_X1 U174 ( .A1(n791), .A2(n790), .ZN(out[2]) );
  AND2_X1 U174bar ( .A1(n791bar), .A2(n790bar), .ZN(outbar[2]);
  OR2_X1 U175 ( .A1(n789), .A2(n788), .ZN(n790) );
  AND2_X1 U175bar ( .A1(n789bar), .A2(n788bar), .ZN(n790bar);
  OR2_X1 U176 ( .A1(n787), .A2(n786), .ZN(n788) );
  AND2_X1 U176bar ( .A1(n787bar), .A2(n786bar), .ZN(n788bar);
  OR2_X1 U177 ( .A1(n819), .A2(n785), .ZN(n786) );
  AND2_X1 U177bar ( .A1(n819bar), .A2(n785bar), .ZN(n786bar);
  OR2_X1 U178 ( .A1(n784), .A2(n783), .ZN(n819) );
  AND2_X1 U178bar ( .A1(n784bar), .A2(n783bar), .ZN(n819bar);
  OR2_X1 U179 ( .A1(n782), .A2(n781), .ZN(n783) );
  AND2_X1 U179bar ( .A1(n782bar), .A2(n781bar), .ZN(n783bar);
  OR2_X1 U180 ( .A1(n780), .A2(n779), .ZN(n781) );
  AND2_X1 U180bar ( .A1(n780bar), .A2(n779bar), .ZN(n781bar);
  OR2_X1 U181 ( .A1(n962), .A2(n778), .ZN(n779) );
  AND2_X1 U181bar ( .A1(n962bar), .A2(n778bar), .ZN(n779bar);
  OR2_X1 U182 ( .A1(n777), .A2(n776), .ZN(n962) );
  AND2_X1 U182bar ( .A1(n777bar), .A2(n776bar), .ZN(n962bar);
  OR2_X1 U183 ( .A1(n775), .A2(n774), .ZN(n776) );
  AND2_X1 U183bar ( .A1(n775bar), .A2(n774bar), .ZN(n776bar);
  OR2_X1 U184 ( .A1(n773), .A2(n772), .ZN(n774) );
  AND2_X1 U184bar ( .A1(n773bar), .A2(n772bar), .ZN(n774bar);
  OR2_X1 U185 ( .A1(in[131]), .A2(in[120]), .ZN(n772) );
  AND2_X1 U185bar ( .A1(inbar[131]), .A2(inbar[120]), .ZN(n772bar);
  OR2_X1 U186 ( .A1(in[153]), .A2(in[147]), .ZN(n773) );
  AND2_X1 U186bar ( .A1(inbar[153]), .A2(inbar[147]), .ZN(n773bar);
  OR2_X1 U187 ( .A1(n771), .A2(n770), .ZN(n775) );
  AND2_X1 U187bar ( .A1(n771bar), .A2(n770bar), .ZN(n775bar);
  OR2_X1 U188 ( .A1(in[170]), .A2(in[156]), .ZN(n770) );
  AND2_X1 U188bar ( .A1(inbar[170]), .A2(inbar[156]), .ZN(n770bar);
  OR2_X1 U189 ( .A1(in[223]), .A2(in[190]), .ZN(n771) );
  AND2_X1 U189bar ( .A1(inbar[223]), .A2(inbar[190]), .ZN(n771bar);
  OR2_X1 U190 ( .A1(n769), .A2(n768), .ZN(n777) );
  AND2_X1 U190bar ( .A1(n769bar), .A2(n768bar), .ZN(n777bar);
  OR2_X1 U191 ( .A1(n767), .A2(n766), .ZN(n768) );
  AND2_X1 U191bar ( .A1(n767bar), .A2(n766bar), .ZN(n768bar);
  OR2_X1 U192 ( .A1(in[236]), .A2(in[230]), .ZN(n766) );
  AND2_X1 U192bar ( .A1(inbar[236]), .A2(inbar[230]), .ZN(n766bar);
  OR2_X1 U193 ( .A1(in[85]), .A2(in[240]), .ZN(n767) );
  AND2_X1 U193bar ( .A1(inbar[85]), .A2(inbar[240]), .ZN(n767bar);
  OR2_X1 U194 ( .A1(n765), .A2(n764), .ZN(n769) );
  AND2_X1 U194bar ( .A1(n765bar), .A2(n764bar), .ZN(n769bar);
  OR2_X1 U195 ( .A1(in_12), .A2(in[90]), .ZN(n764) );
  AND2_X1 U195bar ( .A1(in_12bar), .A2(inbar[90]), .ZN(n764bar);
  OR2_X1 U196 ( .A1(in_39), .A2(in_28), .ZN(n765) );
  AND2_X1 U196bar ( .A1(in_39bar), .A2(in_28bar), .ZN(n765bar);
  OR2_X1 U197 ( .A1(in[109]), .A2(n763), .ZN(n780) );
  AND2_X1 U197bar ( .A1(inbar[109]), .A2(n763bar), .ZN(n780bar);
  OR2_X1 U198 ( .A1(n762), .A2(n761), .ZN(n782) );
  AND2_X1 U198bar ( .A1(n762bar), .A2(n761bar), .ZN(n782bar);
  OR2_X1 U199 ( .A1(in[138]), .A2(in[129]), .ZN(n761) );
  AND2_X1 U199bar ( .A1(inbar[138]), .A2(inbar[129]), .ZN(n761bar);
  OR2_X1 U200 ( .A1(in[157]), .A2(n760), .ZN(n762) );
  AND2_X1 U200bar ( .A1(inbar[157]), .A2(n760bar), .ZN(n762bar);
  OR2_X1 U201 ( .A1(in[182]), .A2(in[167]), .ZN(n760) );
  AND2_X1 U201bar ( .A1(inbar[182]), .A2(inbar[167]), .ZN(n760bar);
  OR2_X1 U202 ( .A1(n759), .A2(n758), .ZN(n784) );
  AND2_X1 U202bar ( .A1(n759bar), .A2(n758bar), .ZN(n784bar);
  OR2_X1 U203 ( .A1(n757), .A2(n756), .ZN(n758) );
  AND2_X1 U203bar ( .A1(n757bar), .A2(n756bar), .ZN(n758bar);
  OR2_X1 U204 ( .A1(in[195]), .A2(in[184]), .ZN(n756) );
  AND2_X1 U204bar ( .A1(inbar[195]), .A2(inbar[184]), .ZN(n756bar);
  OR2_X1 U205 ( .A1(in[196]), .A2(n755), .ZN(n757) );
  AND2_X1 U205bar ( .A1(inbar[196]), .A2(n755bar), .ZN(n757bar);
  OR2_X1 U206 ( .A1(in[215]), .A2(in[209]), .ZN(n755) );
  AND2_X1 U206bar ( .A1(inbar[215]), .A2(inbar[209]), .ZN(n755bar);
  OR2_X1 U207 ( .A1(n754), .A2(n753), .ZN(n759) );
  AND2_X1 U207bar ( .A1(n754bar), .A2(n753bar), .ZN(n759bar);
  OR2_X1 U208 ( .A1(in[93]), .A2(in[233]), .ZN(n753) );
  AND2_X1 U208bar ( .A1(inbar[93]), .A2(inbar[233]), .ZN(n753bar);
  OR2_X1 U209 ( .A1(in_1), .A2(n752), .ZN(n754) );
  AND2_X1 U209bar ( .A1(in_1bar), .A2(n752bar), .ZN(n754bar);
  OR2_X1 U210 ( .A1(in_69), .A2(in_66), .ZN(n752) );
  AND2_X1 U210bar ( .A1(in_69bar), .A2(in_66bar), .ZN(n752bar);
  OR2_X1 U211 ( .A1(n966), .A2(n751), .ZN(n787) );
  AND2_X1 U211bar ( .A1(n966bar), .A2(n751bar), .ZN(n787bar);
  OR2_X1 U212 ( .A1(in[134]), .A2(n750), .ZN(n751) );
  AND2_X1 U212bar ( .A1(inbar[134]), .A2(n750bar), .ZN(n751bar);
  OR2_X1 U213 ( .A1(n749), .A2(n748), .ZN(n966) );
  AND2_X1 U213bar ( .A1(n749bar), .A2(n748bar), .ZN(n966bar);
  OR2_X1 U214 ( .A1(n747), .A2(n746), .ZN(n748) );
  AND2_X1 U214bar ( .A1(n747bar), .A2(n746bar), .ZN(n748bar);
  OR2_X1 U215 ( .A1(n745), .A2(n744), .ZN(n746) );
  AND2_X1 U215bar ( .A1(n745bar), .A2(n744bar), .ZN(n746bar);
  OR2_X1 U216 ( .A1(in[136]), .A2(in[121]), .ZN(n744) );
  AND2_X1 U216bar ( .A1(inbar[136]), .A2(inbar[121]), .ZN(n744bar);
  OR2_X1 U217 ( .A1(in[186]), .A2(in[174]), .ZN(n745) );
  AND2_X1 U217bar ( .A1(inbar[186]), .A2(inbar[174]), .ZN(n745bar);
  OR2_X1 U218 ( .A1(n743), .A2(n742), .ZN(n747) );
  AND2_X1 U218bar ( .A1(n743bar), .A2(n742bar), .ZN(n747bar);
  OR2_X1 U219 ( .A1(in[198]), .A2(in[197]), .ZN(n742) );
  AND2_X1 U219bar ( .A1(inbar[198]), .A2(inbar[197]), .ZN(n742bar);
  OR2_X1 U220 ( .A1(in[214]), .A2(in[199]), .ZN(n743) );
  AND2_X1 U220bar ( .A1(inbar[214]), .A2(inbar[199]), .ZN(n743bar);
  OR2_X1 U221 ( .A1(n741), .A2(n740), .ZN(n749) );
  AND2_X1 U221bar ( .A1(n741bar), .A2(n740bar), .ZN(n749bar);
  OR2_X1 U222 ( .A1(n739), .A2(n738), .ZN(n740) );
  AND2_X1 U222bar ( .A1(n739bar), .A2(n738bar), .ZN(n740bar);
  OR2_X1 U223 ( .A1(in[231]), .A2(in[220]), .ZN(n738) );
  AND2_X1 U223bar ( .A1(inbar[231]), .A2(inbar[220]), .ZN(n738bar);
  OR2_X1 U224 ( .A1(in_25), .A2(in[245]), .ZN(n739) );
  AND2_X1 U224bar ( .A1(in_25bar), .A2(inbar[245]), .ZN(n739bar);
  OR2_X1 U225 ( .A1(n737), .A2(n736), .ZN(n741) );
  AND2_X1 U225bar ( .A1(n737bar), .A2(n736bar), .ZN(n741bar);
  OR2_X1 U226 ( .A1(in_53), .A2(in_29), .ZN(n736) );
  AND2_X1 U226bar ( .A1(in_53bar), .A2(in_29bar), .ZN(n736bar);
  OR2_X1 U227 ( .A1(in_79), .A2(in_74), .ZN(n737) );
  AND2_X1 U227bar ( .A1(in_79bar), .A2(in_74bar), .ZN(n737bar);
  OR2_X1 U228 ( .A1(n735), .A2(n734), .ZN(n789) );
  AND2_X1 U228bar ( .A1(n735bar), .A2(n734bar), .ZN(n789bar);
  OR2_X1 U229 ( .A1(in[152]), .A2(in[140]), .ZN(n734) );
  AND2_X1 U229bar ( .A1(inbar[152]), .A2(inbar[140]), .ZN(n734bar);
  OR2_X1 U230 ( .A1(in[155]), .A2(n733), .ZN(n735) );
  AND2_X1 U230bar ( .A1(inbar[155]), .A2(n733bar), .ZN(n735bar);
  OR2_X1 U231 ( .A1(in[166]), .A2(in[165]), .ZN(n733) );
  AND2_X1 U231bar ( .A1(inbar[166]), .A2(inbar[165]), .ZN(n733bar);
  OR2_X1 U232 ( .A1(n732), .A2(n731), .ZN(n791) );
  AND2_X1 U232bar ( .A1(n732bar), .A2(n731bar), .ZN(n791bar);
  OR2_X1 U233 ( .A1(n730), .A2(n729), .ZN(n731) );
  AND2_X1 U233bar ( .A1(n730bar), .A2(n729bar), .ZN(n731bar);
  OR2_X1 U234 ( .A1(in[202]), .A2(in[185]), .ZN(n729) );
  AND2_X1 U234bar ( .A1(inbar[202]), .A2(inbar[185]), .ZN(n729bar);
  OR2_X1 U235 ( .A1(in[211]), .A2(n728), .ZN(n730) );
  AND2_X1 U235bar ( .A1(inbar[211]), .A2(n728bar), .ZN(n730bar);
  OR2_X1 U236 ( .A1(in[255]), .A2(in[253]), .ZN(n728) );
  AND2_X1 U236bar ( .A1(inbar[255]), .A2(inbar[253]), .ZN(n728bar);
  OR2_X1 U237 ( .A1(n727), .A2(n726), .ZN(n732) );
  AND2_X1 U237bar ( .A1(n727bar), .A2(n726bar), .ZN(n732bar);
  OR2_X1 U238 ( .A1(in_35), .A2(in_15), .ZN(n726) );
  AND2_X1 U238bar ( .A1(in_35bar), .A2(in_15bar), .ZN(n726bar);
  OR2_X1 U239 ( .A1(in_36), .A2(n725), .ZN(n727) );
  AND2_X1 U239bar ( .A1(in_36bar), .A2(n725bar), .ZN(n727bar);
  OR2_X1 U240 ( .A1(in_48), .A2(in_40), .ZN(n725) );
  AND2_X1 U240bar ( .A1(in_48bar), .A2(in_40bar), .ZN(n725bar);
  OR2_X1 U241 ( .A1(n724), .A2(n723), .ZN(out[1]) );
  AND2_X1 U241bar ( .A1(n724bar), .A2(n723bar), .ZN(outbar[1]);
  OR2_X1 U242 ( .A1(n722), .A2(n721), .ZN(n723) );
  AND2_X1 U242bar ( .A1(n722bar), .A2(n721bar), .ZN(n723bar);
  OR2_X1 U243 ( .A1(n720), .A2(n719), .ZN(n721) );
  AND2_X1 U243bar ( .A1(n720bar), .A2(n719bar), .ZN(n721bar);
  OR2_X1 U244 ( .A1(n921), .A2(n887), .ZN(n719) );
  AND2_X1 U244bar ( .A1(n921bar), .A2(n887bar), .ZN(n719bar);
  OR2_X1 U245 ( .A1(n718), .A2(n717), .ZN(n887) );
  AND2_X1 U245bar ( .A1(n718bar), .A2(n717bar), .ZN(n887bar);
  OR2_X1 U246 ( .A1(n716), .A2(n715), .ZN(n717) );
  AND2_X1 U246bar ( .A1(n716bar), .A2(n715bar), .ZN(n717bar);
  OR2_X1 U247 ( .A1(n714), .A2(n713), .ZN(n715) );
  AND2_X1 U247bar ( .A1(n714bar), .A2(n713bar), .ZN(n715bar);
  OR2_X1 U248 ( .A1(in[116]), .A2(in[110]), .ZN(n713) );
  AND2_X1 U248bar ( .A1(inbar[116]), .A2(inbar[110]), .ZN(n713bar);
  OR2_X1 U249 ( .A1(in[133]), .A2(in[130]), .ZN(n714) );
  AND2_X1 U249bar ( .A1(inbar[133]), .A2(inbar[130]), .ZN(n714bar);
  OR2_X1 U250 ( .A1(n712), .A2(n711), .ZN(n716) );
  AND2_X1 U250bar ( .A1(n712bar), .A2(n711bar), .ZN(n716bar);
  OR2_X1 U251 ( .A1(in[203]), .A2(in[135]), .ZN(n711) );
  AND2_X1 U251bar ( .A1(inbar[203]), .A2(inbar[135]), .ZN(n711bar);
  OR2_X1 U252 ( .A1(in[232]), .A2(in[223]), .ZN(n712) );
  AND2_X1 U252bar ( .A1(inbar[232]), .A2(inbar[223]), .ZN(n712bar);
  OR2_X1 U253 ( .A1(n710), .A2(n709), .ZN(n718) );
  AND2_X1 U253bar ( .A1(n710bar), .A2(n709bar), .ZN(n718bar);
  OR2_X1 U254 ( .A1(n708), .A2(n707), .ZN(n709) );
  AND2_X1 U254bar ( .A1(n708bar), .A2(n707bar), .ZN(n709bar);
  OR2_X1 U255 ( .A1(in[255]), .A2(in[233]), .ZN(n707) );
  AND2_X1 U255bar ( .A1(inbar[255]), .A2(inbar[233]), .ZN(n707bar);
  OR2_X1 U256 ( .A1(in_53), .A2(in_34), .ZN(n708) );
  AND2_X1 U256bar ( .A1(in_53bar), .A2(in_34bar), .ZN(n708bar);
  OR2_X1 U257 ( .A1(n706), .A2(n705), .ZN(n710) );
  AND2_X1 U257bar ( .A1(n706bar), .A2(n705bar), .ZN(n710bar);
  OR2_X1 U258 ( .A1(in_57), .A2(in_55), .ZN(n705) );
  AND2_X1 U258bar ( .A1(in_57bar), .A2(in_55bar), .ZN(n705bar);
  OR2_X1 U259 ( .A1(in_68), .A2(in_67), .ZN(n706) );
  AND2_X1 U259bar ( .A1(in_68bar), .A2(in_67bar), .ZN(n706bar);
  OR2_X1 U260 ( .A1(n704), .A2(n703), .ZN(n921) );
  AND2_X1 U260bar ( .A1(n704bar), .A2(n703bar), .ZN(n921bar);
  OR2_X1 U261 ( .A1(n702), .A2(n701), .ZN(n703) );
  AND2_X1 U261bar ( .A1(n702bar), .A2(n701bar), .ZN(n703bar);
  OR2_X1 U262 ( .A1(n700), .A2(n699), .ZN(n701) );
  AND2_X1 U262bar ( .A1(n700bar), .A2(n699bar), .ZN(n701bar);
  OR2_X1 U263 ( .A1(n944), .A2(n872), .ZN(n699) );
  AND2_X1 U263bar ( .A1(n944bar), .A2(n872bar), .ZN(n699bar);
  OR2_X1 U264 ( .A1(n698), .A2(n697), .ZN(n872) );
  AND2_X1 U264bar ( .A1(n698bar), .A2(n697bar), .ZN(n872bar);
  OR2_X1 U265 ( .A1(n696), .A2(n695), .ZN(n697) );
  AND2_X1 U265bar ( .A1(n696bar), .A2(n695bar), .ZN(n697bar);
  OR2_X1 U266 ( .A1(n694), .A2(n693), .ZN(n695) );
  AND2_X1 U266bar ( .A1(n694bar), .A2(n693bar), .ZN(n695bar);
  OR2_X1 U267 ( .A1(in[121]), .A2(in[102]), .ZN(n693) );
  AND2_X1 U267bar ( .A1(inbar[121]), .A2(inbar[102]), .ZN(n693bar);
  OR2_X1 U268 ( .A1(in[162]), .A2(in[161]), .ZN(n694) );
  AND2_X1 U268bar ( .A1(inbar[162]), .A2(inbar[161]), .ZN(n694bar);
  OR2_X1 U269 ( .A1(n692), .A2(n691), .ZN(n696) );
  AND2_X1 U269bar ( .A1(n692bar), .A2(n691bar), .ZN(n696bar);
  OR2_X1 U270 ( .A1(in[192]), .A2(in[178]), .ZN(n691) );
  AND2_X1 U270bar ( .A1(inbar[192]), .A2(inbar[178]), .ZN(n691bar);
  OR2_X1 U271 ( .A1(in[244]), .A2(in[209]), .ZN(n692) );
  AND2_X1 U271bar ( .A1(inbar[244]), .A2(inbar[209]), .ZN(n692bar);
  OR2_X1 U272 ( .A1(n690), .A2(n689), .ZN(n698) );
  AND2_X1 U272bar ( .A1(n690bar), .A2(n689bar), .ZN(n698bar);
  OR2_X1 U273 ( .A1(n688), .A2(n687), .ZN(n689) );
  AND2_X1 U273bar ( .A1(n688bar), .A2(n687bar), .ZN(n689bar);
  OR2_X1 U274 ( .A1(in[90]), .A2(in[254]), .ZN(n687) );
  AND2_X1 U274bar ( .A1(inbar[90]), .A2(inbar[254]), .ZN(n687bar);
  OR2_X1 U275 ( .A1(in_36), .A2(in_32), .ZN(n688) );
  AND2_X1 U275bar ( .A1(in_36bar), .A2(in_32bar), .ZN(n688bar);
  OR2_X1 U276 ( .A1(n686), .A2(n685), .ZN(n690) );
  AND2_X1 U276bar ( .A1(n686bar), .A2(n685bar), .ZN(n690bar);
  OR2_X1 U277 ( .A1(in_62), .A2(in_37), .ZN(n685) );
  AND2_X1 U277bar ( .A1(in_62bar), .A2(in_37bar), .ZN(n685bar);
  OR2_X1 U278 ( .A1(in_75), .A2(in_73), .ZN(n686) );
  AND2_X1 U278bar ( .A1(in_75bar), .A2(in_73bar), .ZN(n686bar);
  OR2_X1 U279 ( .A1(n684), .A2(n683), .ZN(n944) );
  AND2_X1 U279bar ( .A1(n684bar), .A2(n683bar), .ZN(n944bar);
  OR2_X1 U280 ( .A1(n682), .A2(n681), .ZN(n683) );
  AND2_X1 U280bar ( .A1(n682bar), .A2(n681bar), .ZN(n683bar);
  OR2_X1 U281 ( .A1(n680), .A2(n679), .ZN(n681) );
  AND2_X1 U281bar ( .A1(n680bar), .A2(n679bar), .ZN(n681bar);
  OR2_X1 U282 ( .A1(in[171]), .A2(in[153]), .ZN(n679) );
  AND2_X1 U282bar ( .A1(inbar[171]), .A2(inbar[153]), .ZN(n679bar);
  OR2_X1 U283 ( .A1(in[187]), .A2(in[176]), .ZN(n680) );
  AND2_X1 U283bar ( .A1(inbar[187]), .A2(inbar[176]), .ZN(n680bar);
  OR2_X1 U284 ( .A1(n678), .A2(n677), .ZN(n682) );
  AND2_X1 U284bar ( .A1(n678bar), .A2(n677bar), .ZN(n682bar);
  OR2_X1 U285 ( .A1(in[245]), .A2(in[211]), .ZN(n677) );
  AND2_X1 U285bar ( .A1(inbar[245]), .A2(inbar[211]), .ZN(n677bar);
  OR2_X1 U286 ( .A1(in[97]), .A2(in[88]), .ZN(n678) );
  AND2_X1 U286bar ( .A1(inbar[97]), .A2(inbar[88]), .ZN(n678bar);
  OR2_X1 U287 ( .A1(n676), .A2(n675), .ZN(n684) );
  AND2_X1 U287bar ( .A1(n676bar), .A2(n675bar), .ZN(n684bar);
  OR2_X1 U288 ( .A1(n674), .A2(n673), .ZN(n675) );
  AND2_X1 U288bar ( .A1(n674bar), .A2(n673bar), .ZN(n675bar);
  OR2_X1 U289 ( .A1(in_10), .A2(in_0), .ZN(n673) );
  AND2_X1 U289bar ( .A1(in_10bar), .A2(in_0bar), .ZN(n673bar);
  OR2_X1 U290 ( .A1(in_59), .A2(in_5), .ZN(n674) );
  AND2_X1 U290bar ( .A1(in_59bar), .A2(in_5bar), .ZN(n674bar);
  OR2_X1 U291 ( .A1(n672), .A2(n671), .ZN(n676) );
  AND2_X1 U291bar ( .A1(n672bar), .A2(n671bar), .ZN(n676bar);
  OR2_X1 U292 ( .A1(in_60), .A2(in_6), .ZN(n671) );
  AND2_X1 U292bar ( .A1(in_60bar), .A2(in_6bar), .ZN(n671bar);
  OR2_X1 U293 ( .A1(in_77), .A2(in_69), .ZN(n672) );
  AND2_X1 U293bar ( .A1(in_77bar), .A2(in_69bar), .ZN(n672bar);
  OR2_X1 U294 ( .A1(in[113]), .A2(n864), .ZN(n700) );
  AND2_X1 U294bar ( .A1(inbar[113]), .A2(n864bar), .ZN(n700bar);
  OR2_X1 U295 ( .A1(n670), .A2(n669), .ZN(n864) );
  AND2_X1 U295bar ( .A1(n670bar), .A2(n669bar), .ZN(n864bar);
  OR2_X1 U296 ( .A1(n668), .A2(n667), .ZN(n669) );
  AND2_X1 U296bar ( .A1(n668bar), .A2(n667bar), .ZN(n669bar);
  OR2_X1 U297 ( .A1(n666), .A2(n665), .ZN(n667) );
  AND2_X1 U297bar ( .A1(n666bar), .A2(n665bar), .ZN(n667bar);
  OR2_X1 U298 ( .A1(in[125]), .A2(in[107]), .ZN(n665) );
  AND2_X1 U298bar ( .A1(inbar[125]), .A2(inbar[107]), .ZN(n665bar);
  OR2_X1 U299 ( .A1(in[138]), .A2(in[126]), .ZN(n666) );
  AND2_X1 U299bar ( .A1(inbar[138]), .A2(inbar[126]), .ZN(n666bar);
  OR2_X1 U300 ( .A1(n664), .A2(n663), .ZN(n668) );
  AND2_X1 U300bar ( .A1(n664bar), .A2(n663bar), .ZN(n668bar);
  OR2_X1 U301 ( .A1(in[189]), .A2(in[143]), .ZN(n663) );
  AND2_X1 U301bar ( .A1(inbar[189]), .A2(inbar[143]), .ZN(n663bar);
  OR2_X1 U302 ( .A1(in[99]), .A2(in[214]), .ZN(n664) );
  AND2_X1 U302bar ( .A1(inbar[99]), .A2(inbar[214]), .ZN(n664bar);
  OR2_X1 U303 ( .A1(n662), .A2(n661), .ZN(n670) );
  AND2_X1 U303bar ( .A1(n662bar), .A2(n661bar), .ZN(n670bar);
  OR2_X1 U304 ( .A1(n660), .A2(n659), .ZN(n661) );
  AND2_X1 U304bar ( .A1(n660bar), .A2(n659bar), .ZN(n661bar);
  OR2_X1 U305 ( .A1(in_15), .A2(in_12), .ZN(n659) );
  AND2_X1 U305bar ( .A1(in_15bar), .A2(in_12bar), .ZN(n659bar);
  OR2_X1 U306 ( .A1(in_20), .A2(in_2), .ZN(n660) );
  AND2_X1 U306bar ( .A1(in_20bar), .A2(in_2bar), .ZN(n660bar);
  OR2_X1 U307 ( .A1(n658), .A2(n657), .ZN(n662) );
  AND2_X1 U307bar ( .A1(n658bar), .A2(n657bar), .ZN(n662bar);
  OR2_X1 U308 ( .A1(in_30), .A2(in_3), .ZN(n657) );
  AND2_X1 U308bar ( .A1(in_30bar), .A2(in_3bar), .ZN(n657bar);
  OR2_X1 U309 ( .A1(in_4), .A2(in_38), .ZN(n658) );
  AND2_X1 U309bar ( .A1(in_4bar), .A2(in_38bar), .ZN(n658bar);
  OR2_X1 U310 ( .A1(n656), .A2(n655), .ZN(n702) );
  AND2_X1 U310bar ( .A1(n656bar), .A2(n655bar), .ZN(n702bar);
  OR2_X1 U311 ( .A1(in[148]), .A2(in[137]), .ZN(n655) );
  AND2_X1 U311bar ( .A1(inbar[148]), .A2(inbar[137]), .ZN(n655bar);
  OR2_X1 U312 ( .A1(in[149]), .A2(n654), .ZN(n656) );
  AND2_X1 U312bar ( .A1(inbar[149]), .A2(n654bar), .ZN(n656bar);
  OR2_X1 U313 ( .A1(in[195]), .A2(in[190]), .ZN(n654) );
  AND2_X1 U313bar ( .A1(inbar[195]), .A2(inbar[190]), .ZN(n654bar);
  OR2_X1 U314 ( .A1(n653), .A2(n652), .ZN(n704) );
  AND2_X1 U314bar ( .A1(n653bar), .A2(n652bar), .ZN(n704bar);
  OR2_X1 U315 ( .A1(n651), .A2(n650), .ZN(n652) );
  AND2_X1 U315bar ( .A1(n651bar), .A2(n650bar), .ZN(n652bar);
  OR2_X1 U316 ( .A1(in[98]), .A2(in[197]), .ZN(n650) );
  AND2_X1 U316bar ( .A1(inbar[98]), .A2(inbar[197]), .ZN(n650bar);
  OR2_X1 U317 ( .A1(in_11), .A2(n649), .ZN(n651) );
  AND2_X1 U317bar ( .A1(in_11bar), .A2(n649bar), .ZN(n651bar);
  OR2_X1 U318 ( .A1(in_26), .A2(in_14), .ZN(n649) );
  AND2_X1 U318bar ( .A1(in_26bar), .A2(in_14bar), .ZN(n649bar);
  OR2_X1 U319 ( .A1(n648), .A2(n647), .ZN(n653) );
  AND2_X1 U319bar ( .A1(n648bar), .A2(n647bar), .ZN(n653bar);
  OR2_X1 U320 ( .A1(in_35), .A2(in_27), .ZN(n647) );
  AND2_X1 U320bar ( .A1(in_35bar), .A2(in_27bar), .ZN(n647bar);
  OR2_X1 U321 ( .A1(in_50), .A2(n646), .ZN(n648) );
  AND2_X1 U321bar ( .A1(in_50bar), .A2(n646bar), .ZN(n648bar);
  OR2_X1 U322 ( .A1(in_78), .A2(in_61), .ZN(n646) );
  AND2_X1 U322bar ( .A1(in_78bar), .A2(in_61bar), .ZN(n646bar);
  OR2_X1 U323 ( .A1(n942), .A2(n645), .ZN(n720) );
  AND2_X1 U323bar ( .A1(n942bar), .A2(n645bar), .ZN(n720bar);
  OR2_X1 U324 ( .A1(in[106]), .A2(n863), .ZN(n645) );
  AND2_X1 U324bar ( .A1(inbar[106]), .A2(n863bar), .ZN(n645bar);
  OR2_X1 U325 ( .A1(n644), .A2(n643), .ZN(n863) );
  AND2_X1 U325bar ( .A1(n644bar), .A2(n643bar), .ZN(n863bar);
  OR2_X1 U326 ( .A1(n642), .A2(n641), .ZN(n643) );
  AND2_X1 U326bar ( .A1(n642bar), .A2(n641bar), .ZN(n643bar);
  OR2_X1 U327 ( .A1(n640), .A2(n639), .ZN(n641) );
  AND2_X1 U327bar ( .A1(n640bar), .A2(n639bar), .ZN(n641bar);
  OR2_X1 U328 ( .A1(in[127]), .A2(in[122]), .ZN(n639) );
  AND2_X1 U328bar ( .A1(inbar[127]), .A2(inbar[122]), .ZN(n639bar);
  OR2_X1 U329 ( .A1(in[156]), .A2(in[132]), .ZN(n640) );
  AND2_X1 U329bar ( .A1(inbar[156]), .A2(inbar[132]), .ZN(n640bar);
  OR2_X1 U330 ( .A1(n638), .A2(n637), .ZN(n642) );
  AND2_X1 U330bar ( .A1(n638bar), .A2(n637bar), .ZN(n642bar);
  OR2_X1 U331 ( .A1(in[159]), .A2(in[157]), .ZN(n637) );
  AND2_X1 U331bar ( .A1(inbar[159]), .A2(inbar[157]), .ZN(n637bar);
  OR2_X1 U332 ( .A1(in[185]), .A2(in[169]), .ZN(n638) );
  AND2_X1 U332bar ( .A1(inbar[185]), .A2(inbar[169]), .ZN(n638bar);
  OR2_X1 U333 ( .A1(n636), .A2(n635), .ZN(n644) );
  AND2_X1 U333bar ( .A1(n636bar), .A2(n635bar), .ZN(n644bar);
  OR2_X1 U334 ( .A1(n634), .A2(n633), .ZN(n635) );
  AND2_X1 U334bar ( .A1(n634bar), .A2(n633bar), .ZN(n635bar);
  OR2_X1 U335 ( .A1(in[239]), .A2(in[218]), .ZN(n633) );
  AND2_X1 U335bar ( .A1(inbar[239]), .A2(inbar[218]), .ZN(n633bar);
  OR2_X1 U336 ( .A1(in_13), .A2(in[87]), .ZN(n634) );
  AND2_X1 U336bar ( .A1(in_13bar), .A2(inbar[87]), .ZN(n634bar);
  OR2_X1 U337 ( .A1(n632), .A2(n631), .ZN(n636) );
  AND2_X1 U337bar ( .A1(n632bar), .A2(n631bar), .ZN(n636bar);
  OR2_X1 U338 ( .A1(in_72), .A2(in_70), .ZN(n631) );
  AND2_X1 U338bar ( .A1(in_72bar), .A2(in_70bar), .ZN(n631bar);
  OR2_X1 U339 ( .A1(in_80), .A2(in_74), .ZN(n632) );
  AND2_X1 U339bar ( .A1(in_80bar), .A2(in_74bar), .ZN(n632bar);
  OR2_X1 U340 ( .A1(n630), .A2(n629), .ZN(n942) );
  AND2_X1 U340bar ( .A1(n630bar), .A2(n629bar), .ZN(n942bar);
  OR2_X1 U341 ( .A1(n628), .A2(n627), .ZN(n629) );
  AND2_X1 U341bar ( .A1(n628bar), .A2(n627bar), .ZN(n629bar);
  OR2_X1 U342 ( .A1(n626), .A2(n625), .ZN(n627) );
  AND2_X1 U342bar ( .A1(n626bar), .A2(n625bar), .ZN(n627bar);
  OR2_X1 U343 ( .A1(in[146]), .A2(in[100]), .ZN(n625) );
  AND2_X1 U343bar ( .A1(inbar[146]), .A2(inbar[100]), .ZN(n625bar);
  OR2_X1 U344 ( .A1(in[168]), .A2(in[152]), .ZN(n626) );
  AND2_X1 U344bar ( .A1(inbar[168]), .A2(inbar[152]), .ZN(n626bar);
  OR2_X1 U345 ( .A1(n624), .A2(n623), .ZN(n628) );
  AND2_X1 U345bar ( .A1(n624bar), .A2(n623bar), .ZN(n628bar);
  OR2_X1 U346 ( .A1(in[199]), .A2(in[182]), .ZN(n623) );
  AND2_X1 U346bar ( .A1(inbar[199]), .A2(inbar[182]), .ZN(n623bar);
  OR2_X1 U347 ( .A1(in[236]), .A2(in[204]), .ZN(n624) );
  AND2_X1 U347bar ( .A1(inbar[236]), .A2(inbar[204]), .ZN(n624bar);
  OR2_X1 U348 ( .A1(n622), .A2(n621), .ZN(n630) );
  AND2_X1 U348bar ( .A1(n622bar), .A2(n621bar), .ZN(n630bar);
  OR2_X1 U349 ( .A1(n620), .A2(n619), .ZN(n621) );
  AND2_X1 U349bar ( .A1(n620bar), .A2(n619bar), .ZN(n621bar);
  OR2_X1 U350 ( .A1(in[89]), .A2(in[246]), .ZN(n619) );
  AND2_X1 U350bar ( .A1(inbar[89]), .A2(inbar[246]), .ZN(n619bar);
  OR2_X1 U351 ( .A1(in[95]), .A2(in[92]), .ZN(n620) );
  AND2_X1 U351bar ( .A1(inbar[95]), .A2(inbar[92]), .ZN(n620bar);
  OR2_X1 U352 ( .A1(n618), .A2(n617), .ZN(n622) );
  AND2_X1 U352bar ( .A1(n618bar), .A2(n617bar), .ZN(n622bar);
  OR2_X1 U353 ( .A1(in_22), .A2(in_16), .ZN(n617) );
  AND2_X1 U353bar ( .A1(in_22bar), .A2(in_16bar), .ZN(n617bar);
  OR2_X1 U354 ( .A1(in_51), .A2(in_49), .ZN(n618) );
  AND2_X1 U354bar ( .A1(in_51bar), .A2(in_49bar), .ZN(n618bar);
  OR2_X1 U355 ( .A1(n616), .A2(n615), .ZN(n722) );
  AND2_X1 U355bar ( .A1(n616bar), .A2(n615bar), .ZN(n722bar);
  OR2_X1 U356 ( .A1(in[158]), .A2(in[115]), .ZN(n615) );
  AND2_X1 U356bar ( .A1(inbar[158]), .A2(inbar[115]), .ZN(n615bar);
  OR2_X1 U357 ( .A1(in[163]), .A2(n614), .ZN(n616) );
  AND2_X1 U357bar ( .A1(inbar[163]), .A2(n614bar), .ZN(n616bar);
  OR2_X1 U358 ( .A1(in[206]), .A2(in[165]), .ZN(n614) );
  AND2_X1 U358bar ( .A1(inbar[206]), .A2(inbar[165]), .ZN(n614bar);
  OR2_X1 U359 ( .A1(n613), .A2(n612), .ZN(n724) );
  AND2_X1 U359bar ( .A1(n613bar), .A2(n612bar), .ZN(n724bar);
  OR2_X1 U360 ( .A1(n611), .A2(n610), .ZN(n612) );
  AND2_X1 U360bar ( .A1(n611bar), .A2(n610bar), .ZN(n612bar);
  OR2_X1 U361 ( .A1(in[213]), .A2(in[207]), .ZN(n610) );
  AND2_X1 U361bar ( .A1(inbar[213]), .A2(inbar[207]), .ZN(n610bar);
  OR2_X1 U362 ( .A1(in[215]), .A2(n609), .ZN(n611) );
  AND2_X1 U362bar ( .A1(inbar[215]), .A2(n609bar), .ZN(n611bar);
  OR2_X1 U363 ( .A1(in[230]), .A2(in[220]), .ZN(n609) );
  AND2_X1 U363bar ( .A1(inbar[230]), .A2(inbar[220]), .ZN(n609bar);
  OR2_X1 U364 ( .A1(n608), .A2(n607), .ZN(n613) );
  AND2_X1 U364bar ( .A1(n608bar), .A2(n607bar), .ZN(n613bar);
  OR2_X1 U365 ( .A1(in[251]), .A2(in[234]), .ZN(n607) );
  AND2_X1 U365bar ( .A1(inbar[251]), .A2(inbar[234]), .ZN(n607bar);
  OR2_X1 U366 ( .A1(in_17), .A2(n606), .ZN(n608) );
  AND2_X1 U366bar ( .A1(in_17bar), .A2(n606bar), .ZN(n608bar);
  OR2_X1 U367 ( .A1(in_65), .A2(in_56), .ZN(n606) );
  AND2_X1 U367bar ( .A1(in_65bar), .A2(in_56bar), .ZN(n606bar);
  OR2_X1 U368 ( .A1(n605), .A2(n604), .ZN(out[0]) );
  AND2_X1 U368bar ( .A1(n605bar), .A2(n604bar), .ZN(outbar[0]);
  OR2_X1 U369 ( .A1(n603), .A2(n602), .ZN(n604) );
  AND2_X1 U369bar ( .A1(n603bar), .A2(n602bar), .ZN(n604bar);
  OR2_X1 U370 ( .A1(n601), .A2(n600), .ZN(n602) );
  AND2_X1 U370bar ( .A1(n601bar), .A2(n600bar), .ZN(n602bar);
  OR2_X1 U371 ( .A1(n820), .A2(n785), .ZN(n600) );
  AND2_X1 U371bar ( .A1(n820bar), .A2(n785bar), .ZN(n600bar);
  OR2_X1 U372 ( .A1(n599), .A2(n598), .ZN(n785) );
  AND2_X1 U372bar ( .A1(n599bar), .A2(n598bar), .ZN(n785bar);
  OR2_X1 U373 ( .A1(n597), .A2(n596), .ZN(n598) );
  AND2_X1 U373bar ( .A1(n597bar), .A2(n596bar), .ZN(n598bar);
  OR2_X1 U374 ( .A1(n595), .A2(n594), .ZN(n596) );
  AND2_X1 U374bar ( .A1(n595bar), .A2(n594bar), .ZN(n596bar);
  OR2_X1 U375 ( .A1(in[135]), .A2(in[104]), .ZN(n594) );
  AND2_X1 U375bar ( .A1(inbar[135]), .A2(inbar[104]), .ZN(n594bar);
  OR2_X1 U376 ( .A1(in[188]), .A2(in[178]), .ZN(n595) );
  AND2_X1 U376bar ( .A1(inbar[188]), .A2(inbar[178]), .ZN(n595bar);
  OR2_X1 U377 ( .A1(n593), .A2(n592), .ZN(n597) );
  AND2_X1 U377bar ( .A1(n593bar), .A2(n592bar), .ZN(n597bar);
  OR2_X1 U378 ( .A1(in[217]), .A2(in[194]), .ZN(n592) );
  AND2_X1 U378bar ( .A1(inbar[217]), .A2(inbar[194]), .ZN(n592bar);
  OR2_X1 U379 ( .A1(in[237]), .A2(in[218]), .ZN(n593) );
  AND2_X1 U379bar ( .A1(inbar[237]), .A2(inbar[218]), .ZN(n593bar);
  OR2_X1 U380 ( .A1(n591), .A2(n590), .ZN(n599) );
  AND2_X1 U380bar ( .A1(n591bar), .A2(n590bar), .ZN(n599bar);
  OR2_X1 U381 ( .A1(n589), .A2(n588), .ZN(n590) );
  AND2_X1 U381bar ( .A1(n589bar), .A2(n588bar), .ZN(n590bar);
  OR2_X1 U382 ( .A1(in_2), .A2(in_10), .ZN(n588) );
  AND2_X1 U382bar ( .A1(in_2bar), .A2(in_10bar), .ZN(n588bar);
  OR2_X1 U383 ( .A1(in_47), .A2(in_22), .ZN(n589) );
  AND2_X1 U383bar ( .A1(in_47bar), .A2(in_22bar), .ZN(n589bar);
  OR2_X1 U384 ( .A1(n587), .A2(n586), .ZN(n591) );
  AND2_X1 U384bar ( .A1(n587bar), .A2(n586bar), .ZN(n591bar);
  OR2_X1 U385 ( .A1(in_56), .A2(in_54), .ZN(n586) );
  AND2_X1 U385bar ( .A1(in_56bar), .A2(in_54bar), .ZN(n586bar);
  OR2_X1 U386 ( .A1(in_63), .A2(in_61), .ZN(n587) );
  AND2_X1 U386bar ( .A1(in_63bar), .A2(in_61bar), .ZN(n587bar);
  OR2_X1 U387 ( .A1(n585), .A2(n584), .ZN(n820) );
  AND2_X1 U387bar ( .A1(n585bar), .A2(n584bar), .ZN(n820bar);
  OR2_X1 U388 ( .A1(n583), .A2(n582), .ZN(n584) );
  AND2_X1 U388bar ( .A1(n583bar), .A2(n582bar), .ZN(n584bar);
  OR2_X1 U389 ( .A1(n581), .A2(n580), .ZN(n582) );
  AND2_X1 U389bar ( .A1(n581bar), .A2(n580bar), .ZN(n582bar);
  OR2_X1 U390 ( .A1(in[158]), .A2(in[142]), .ZN(n580) );
  AND2_X1 U390bar ( .A1(inbar[158]), .A2(inbar[142]), .ZN(n580bar);
  OR2_X1 U391 ( .A1(in[175]), .A2(in[164]), .ZN(n581) );
  AND2_X1 U391bar ( .A1(inbar[175]), .A2(inbar[164]), .ZN(n581bar);
  OR2_X1 U392 ( .A1(n579), .A2(n578), .ZN(n583) );
  AND2_X1 U392bar ( .A1(n579bar), .A2(n578bar), .ZN(n583bar);
  OR2_X1 U393 ( .A1(in[228]), .A2(in[204]), .ZN(n578) );
  AND2_X1 U393bar ( .A1(inbar[228]), .A2(inbar[204]), .ZN(n578bar);
  OR2_X1 U394 ( .A1(in[91]), .A2(in[87]), .ZN(n579) );
  AND2_X1 U394bar ( .A1(inbar[91]), .A2(inbar[87]), .ZN(n579bar);
  OR2_X1 U395 ( .A1(n577), .A2(n576), .ZN(n585) );
  AND2_X1 U395bar ( .A1(n577bar), .A2(n576bar), .ZN(n585bar);
  OR2_X1 U396 ( .A1(n575), .A2(n574), .ZN(n576) );
  AND2_X1 U396bar ( .A1(n575bar), .A2(n574bar), .ZN(n576bar);
  OR2_X1 U397 ( .A1(in_21), .A2(in_11), .ZN(n574) );
  AND2_X1 U397bar ( .A1(in_21bar), .A2(in_11bar), .ZN(n574bar);
  OR2_X1 U398 ( .A1(in_5), .A2(in_3), .ZN(n575) );
  AND2_X1 U398bar ( .A1(in_5bar), .A2(in_3bar), .ZN(n575bar);
  OR2_X1 U399 ( .A1(n573), .A2(n572), .ZN(n577) );
  AND2_X1 U399bar ( .A1(n573bar), .A2(n572bar), .ZN(n577bar);
  OR2_X1 U400 ( .A1(in_68), .A2(in_64), .ZN(n572) );
  AND2_X1 U400bar ( .A1(in_68bar), .A2(in_64bar), .ZN(n572bar);
  OR2_X1 U401 ( .A1(in_76), .A2(in_73), .ZN(n573) );
  AND2_X1 U401bar ( .A1(in_76bar), .A2(in_73bar), .ZN(n573bar);
  OR2_X1 U402 ( .A1(n778), .A2(n571), .ZN(n601) );
  AND2_X1 U402bar ( .A1(n778bar), .A2(n571bar), .ZN(n601bar);
  OR2_X1 U403 ( .A1(in[100]), .A2(n965), .ZN(n571) );
  AND2_X1 U403bar ( .A1(inbar[100]), .A2(n965bar), .ZN(n571bar);
  OR2_X1 U404 ( .A1(n570), .A2(n569), .ZN(n965) );
  AND2_X1 U404bar ( .A1(n570bar), .A2(n569bar), .ZN(n965bar);
  OR2_X1 U405 ( .A1(n568), .A2(n567), .ZN(n569) );
  AND2_X1 U405bar ( .A1(n568bar), .A2(n567bar), .ZN(n569bar);
  OR2_X1 U406 ( .A1(n566), .A2(n565), .ZN(n567) );
  AND2_X1 U406bar ( .A1(n566bar), .A2(n565bar), .ZN(n567bar);
  OR2_X1 U407 ( .A1(n817), .A2(n750), .ZN(n565) );
  AND2_X1 U407bar ( .A1(n817bar), .A2(n750bar), .ZN(n565bar);
  OR2_X1 U408 ( .A1(n564), .A2(n563), .ZN(n750) );
  AND2_X1 U408bar ( .A1(n564bar), .A2(n563bar), .ZN(n750bar);
  OR2_X1 U409 ( .A1(n562), .A2(n561), .ZN(n563) );
  AND2_X1 U409bar ( .A1(n562bar), .A2(n561bar), .ZN(n563bar);
  OR2_X1 U410 ( .A1(n560), .A2(n559), .ZN(n561) );
  AND2_X1 U410bar ( .A1(n560bar), .A2(n559bar), .ZN(n561bar);
  OR2_X1 U411 ( .A1(in[119]), .A2(in[103]), .ZN(n559) );
  AND2_X1 U411bar ( .A1(inbar[119]), .A2(inbar[103]), .ZN(n559bar);
  OR2_X1 U412 ( .A1(in[137]), .A2(in[133]), .ZN(n560) );
  AND2_X1 U412bar ( .A1(inbar[137]), .A2(inbar[133]), .ZN(n560bar);
  OR2_X1 U413 ( .A1(n558), .A2(n557), .ZN(n562) );
  AND2_X1 U413bar ( .A1(n558bar), .A2(n557bar), .ZN(n562bar);
  OR2_X1 U414 ( .A1(in[176]), .A2(in[173]), .ZN(n557) );
  AND2_X1 U414bar ( .A1(inbar[176]), .A2(inbar[173]), .ZN(n557bar);
  OR2_X1 U415 ( .A1(in[210]), .A2(in[181]), .ZN(n558) );
  AND2_X1 U415bar ( .A1(inbar[210]), .A2(inbar[181]), .ZN(n558bar);
  OR2_X1 U416 ( .A1(n556), .A2(n555), .ZN(n564) );
  AND2_X1 U416bar ( .A1(n556bar), .A2(n555bar), .ZN(n564bar);
  OR2_X1 U417 ( .A1(n554), .A2(n553), .ZN(n555) );
  AND2_X1 U417bar ( .A1(n554bar), .A2(n553bar), .ZN(n555bar);
  OR2_X1 U418 ( .A1(in_13), .A2(in[234]), .ZN(n553) );
  AND2_X1 U418bar ( .A1(in_13bar), .A2(inbar[234]), .ZN(n553bar);
  OR2_X1 U419 ( .A1(in_38), .A2(in_32), .ZN(n554) );
  AND2_X1 U419bar ( .A1(in_38bar), .A2(in_32bar), .ZN(n554bar);
  OR2_X1 U420 ( .A1(n552), .A2(n551), .ZN(n556) );
  AND2_X1 U420bar ( .A1(n552bar), .A2(n551bar), .ZN(n556bar);
  OR2_X1 U421 ( .A1(in_42), .A2(in_41), .ZN(n551) );
  AND2_X1 U421bar ( .A1(in_42bar), .A2(in_41bar), .ZN(n551bar);
  OR2_X1 U422 ( .A1(in_7), .A2(in_49), .ZN(n552) );
  AND2_X1 U422bar ( .A1(in_7bar), .A2(in_49bar), .ZN(n552bar);
  OR2_X1 U423 ( .A1(n550), .A2(n549), .ZN(n817) );
  AND2_X1 U423bar ( .A1(n550bar), .A2(n549bar), .ZN(n817bar);
  OR2_X1 U424 ( .A1(n548), .A2(n547), .ZN(n549) );
  AND2_X1 U424bar ( .A1(n548bar), .A2(n547bar), .ZN(n549bar);
  OR2_X1 U425 ( .A1(n546), .A2(n545), .ZN(n547) );
  AND2_X1 U425bar ( .A1(n546bar), .A2(n545bar), .ZN(n547bar);
  OR2_X1 U426 ( .A1(in[159]), .A2(in[105]), .ZN(n545) );
  AND2_X1 U426bar ( .A1(inbar[159]), .A2(inbar[105]), .ZN(n545bar);
  OR2_X1 U427 ( .A1(in[206]), .A2(in[183]), .ZN(n546) );
  AND2_X1 U427bar ( .A1(inbar[206]), .A2(inbar[183]), .ZN(n546bar);
  OR2_X1 U428 ( .A1(n544), .A2(n543), .ZN(n548) );
  AND2_X1 U428bar ( .A1(n544bar), .A2(n543bar), .ZN(n548bar);
  OR2_X1 U429 ( .A1(in[229]), .A2(in[219]), .ZN(n543) );
  AND2_X1 U429bar ( .A1(inbar[229]), .A2(inbar[219]), .ZN(n543bar);
  OR2_X1 U430 ( .A1(in[235]), .A2(in[232]), .ZN(n544) );
  AND2_X1 U430bar ( .A1(inbar[235]), .A2(inbar[232]), .ZN(n544bar);
  OR2_X1 U431 ( .A1(n542), .A2(n541), .ZN(n550) );
  AND2_X1 U431bar ( .A1(n542bar), .A2(n541bar), .ZN(n550bar);
  OR2_X1 U432 ( .A1(n540), .A2(n539), .ZN(n541) );
  AND2_X1 U432bar ( .A1(n540bar), .A2(n539bar), .ZN(n541bar);
  OR2_X1 U433 ( .A1(in[249]), .A2(in[242]), .ZN(n539) );
  AND2_X1 U433bar ( .A1(inbar[249]), .A2(inbar[242]), .ZN(n539bar);
  OR2_X1 U434 ( .A1(in[89]), .A2(in[254]), .ZN(n540) );
  AND2_X1 U434bar ( .A1(inbar[89]), .A2(inbar[254]), .ZN(n540bar);
  OR2_X1 U435 ( .A1(n538), .A2(n537), .ZN(n542) );
  AND2_X1 U435bar ( .A1(n538bar), .A2(n537bar), .ZN(n542bar);
  OR2_X1 U436 ( .A1(in_14), .A2(in[99]), .ZN(n537) );
  AND2_X1 U436bar ( .A1(in_14bar), .A2(inbar[99]), .ZN(n537bar);
  OR2_X1 U437 ( .A1(in_60), .A2(in_18), .ZN(n538) );
  AND2_X1 U437bar ( .A1(in_60bar), .A2(in_18bar), .ZN(n538bar);
  OR2_X1 U438 ( .A1(in[113]), .A2(n763), .ZN(n566) );
  AND2_X1 U438bar ( .A1(inbar[113]), .A2(n763bar), .ZN(n566bar);
  OR2_X1 U439 ( .A1(n536), .A2(n535), .ZN(n763) );
  AND2_X1 U439bar ( .A1(n536bar), .A2(n535bar), .ZN(n763bar);
  OR2_X1 U440 ( .A1(n534), .A2(n533), .ZN(n535) );
  AND2_X1 U440bar ( .A1(n534bar), .A2(n533bar), .ZN(n535bar);
  OR2_X1 U441 ( .A1(n532), .A2(n531), .ZN(n533) );
  AND2_X1 U441bar ( .A1(n532bar), .A2(n531bar), .ZN(n533bar);
  OR2_X1 U442 ( .A1(in[115]), .A2(in[110]), .ZN(n531) );
  AND2_X1 U442bar ( .A1(inbar[115]), .A2(inbar[110]), .ZN(n531bar);
  OR2_X1 U443 ( .A1(in[125]), .A2(in[117]), .ZN(n532) );
  AND2_X1 U443bar ( .A1(inbar[125]), .A2(inbar[117]), .ZN(n532bar);
  OR2_X1 U444 ( .A1(n530), .A2(n529), .ZN(n534) );
  AND2_X1 U444bar ( .A1(n530bar), .A2(n529bar), .ZN(n534bar);
  OR2_X1 U445 ( .A1(in[180]), .A2(in[128]), .ZN(n529) );
  AND2_X1 U445bar ( .A1(inbar[180]), .A2(inbar[128]), .ZN(n529bar);
  OR2_X1 U446 ( .A1(in[205]), .A2(in[201]), .ZN(n530) );
  AND2_X1 U446bar ( .A1(inbar[205]), .A2(inbar[201]), .ZN(n530bar);
  OR2_X1 U447 ( .A1(n528), .A2(n527), .ZN(n536) );
  AND2_X1 U447bar ( .A1(n528bar), .A2(n527bar), .ZN(n536bar);
  OR2_X1 U448 ( .A1(n526), .A2(n525), .ZN(n527) );
  AND2_X1 U448bar ( .A1(n526bar), .A2(n525bar), .ZN(n527bar);
  OR2_X1 U449 ( .A1(in[244]), .A2(in[239]), .ZN(n525) );
  AND2_X1 U449bar ( .A1(inbar[244]), .A2(inbar[239]), .ZN(n525bar);
  OR2_X1 U450 ( .A1(in[95]), .A2(in[83]), .ZN(n526) );
  AND2_X1 U450bar ( .A1(inbar[95]), .A2(inbar[83]), .ZN(n526bar);
  OR2_X1 U451 ( .A1(n524), .A2(n523), .ZN(n528) );
  AND2_X1 U451bar ( .A1(n524bar), .A2(n523bar), .ZN(n528bar);
  OR2_X1 U452 ( .A1(in_24), .A2(in[97]), .ZN(n523) );
  AND2_X1 U452bar ( .A1(in_24bar), .A2(inbar[97]), .ZN(n523bar);
  OR2_X1 U453 ( .A1(in_33), .A2(in_27), .ZN(n524) );
  AND2_X1 U453bar ( .A1(in_33bar), .A2(in_27bar), .ZN(n524bar);
  OR2_X1 U454 ( .A1(n522), .A2(n521), .ZN(n568) );
  AND2_X1 U454bar ( .A1(n522bar), .A2(n521bar), .ZN(n568bar);
  OR2_X1 U455 ( .A1(in[145]), .A2(in[126]), .ZN(n521) );
  AND2_X1 U455bar ( .A1(inbar[145]), .A2(inbar[126]), .ZN(n521bar);
  OR2_X1 U456 ( .A1(in[169]), .A2(n520), .ZN(n522) );
  AND2_X1 U456bar ( .A1(inbar[169]), .A2(n520bar), .ZN(n522bar);
  OR2_X1 U457 ( .A1(in[221]), .A2(in[172]), .ZN(n520) );
  AND2_X1 U457bar ( .A1(inbar[221]), .A2(inbar[172]), .ZN(n520bar);
  OR2_X1 U458 ( .A1(n519), .A2(n518), .ZN(n570) );
  AND2_X1 U458bar ( .A1(n519bar), .A2(n518bar), .ZN(n570bar);
  OR2_X1 U459 ( .A1(n517), .A2(n516), .ZN(n518) );
  AND2_X1 U459bar ( .A1(n517bar), .A2(n516bar), .ZN(n518bar);
  OR2_X1 U460 ( .A1(in[241]), .A2(in[224]), .ZN(n516) );
  AND2_X1 U460bar ( .A1(inbar[241]), .A2(inbar[224]), .ZN(n516bar);
  OR2_X1 U461 ( .A1(in[86]), .A2(n515), .ZN(n517) );
  AND2_X1 U461bar ( .A1(inbar[86]), .A2(n515bar), .ZN(n517bar);
  OR2_X1 U462 ( .A1(in_43), .A2(in_34), .ZN(n515) );
  AND2_X1 U462bar ( .A1(in_43bar), .A2(in_34bar), .ZN(n515bar);
  OR2_X1 U463 ( .A1(n514), .A2(n513), .ZN(n519) );
  AND2_X1 U463bar ( .A1(n514bar), .A2(n513bar), .ZN(n519bar);
  OR2_X1 U464 ( .A1(in_65), .A2(in_51), .ZN(n513) );
  AND2_X1 U464bar ( .A1(in_65bar), .A2(in_51bar), .ZN(n513bar);
  OR2_X1 U465 ( .A1(in_75), .A2(n512), .ZN(n514) );
  AND2_X1 U465bar ( .A1(in_75bar), .A2(n512bar), .ZN(n514bar);
  OR2_X1 U466 ( .A1(in_81), .A2(in_77), .ZN(n512) );
  AND2_X1 U466bar ( .A1(in_81bar), .A2(in_77bar), .ZN(n512bar);
  OR2_X1 U467 ( .A1(n511), .A2(n510), .ZN(n778) );
  AND2_X1 U467bar ( .A1(n511bar), .A2(n510bar), .ZN(n778bar);
  OR2_X1 U468 ( .A1(n509), .A2(n508), .ZN(n510) );
  AND2_X1 U468bar ( .A1(n509bar), .A2(n508bar), .ZN(n510bar);
  OR2_X1 U469 ( .A1(n507), .A2(n506), .ZN(n508) );
  AND2_X1 U469bar ( .A1(n507bar), .A2(n506bar), .ZN(n508bar);
  OR2_X1 U470 ( .A1(in[107]), .A2(in[101]), .ZN(n506) );
  AND2_X1 U470bar ( .A1(inbar[107]), .A2(inbar[101]), .ZN(n506bar);
  OR2_X1 U471 ( .A1(in[139]), .A2(in[132]), .ZN(n507) );
  AND2_X1 U471bar ( .A1(inbar[139]), .A2(inbar[132]), .ZN(n507bar);
  OR2_X1 U472 ( .A1(n505), .A2(n504), .ZN(n509) );
  AND2_X1 U472bar ( .A1(n505bar), .A2(n504bar), .ZN(n509bar);
  OR2_X1 U473 ( .A1(in[146]), .A2(in[141]), .ZN(n504) );
  AND2_X1 U473bar ( .A1(inbar[146]), .A2(inbar[141]), .ZN(n504bar);
  OR2_X1 U474 ( .A1(in[203]), .A2(in[179]), .ZN(n505) );
  AND2_X1 U474bar ( .A1(inbar[203]), .A2(inbar[179]), .ZN(n505bar);
  OR2_X1 U475 ( .A1(n503), .A2(n502), .ZN(n511) );
  AND2_X1 U475bar ( .A1(n503bar), .A2(n502bar), .ZN(n511bar);
  OR2_X1 U476 ( .A1(n501), .A2(n500), .ZN(n502) );
  AND2_X1 U476bar ( .A1(n501bar), .A2(n500bar), .ZN(n502bar);
  OR2_X1 U477 ( .A1(in[243]), .A2(in[222]), .ZN(n500) );
  AND2_X1 U477bar ( .A1(inbar[243]), .A2(inbar[222]), .ZN(n500bar);
  OR2_X1 U478 ( .A1(in[251]), .A2(in[250]), .ZN(n501) );
  AND2_X1 U478bar ( .A1(inbar[251]), .A2(inbar[250]), .ZN(n501bar);
  OR2_X1 U479 ( .A1(n499), .A2(n498), .ZN(n503) );
  AND2_X1 U479bar ( .A1(n499bar), .A2(n498bar), .ZN(n503bar);
  OR2_X1 U480 ( .A1(in_37), .A2(in_19), .ZN(n498) );
  AND2_X1 U480bar ( .A1(in_37bar), .A2(in_19bar), .ZN(n498bar);
  OR2_X1 U481 ( .A1(in_78), .A2(in_6), .ZN(n499) );
  AND2_X1 U481bar ( .A1(in_78bar), .A2(in_6bar), .ZN(n499bar);
  OR2_X1 U482 ( .A1(n497), .A2(n496), .ZN(n603) );
  AND2_X1 U482bar ( .A1(n497bar), .A2(n496bar), .ZN(n603bar);
  OR2_X1 U483 ( .A1(in[112]), .A2(in[102]), .ZN(n496) );
  AND2_X1 U483bar ( .A1(inbar[112]), .A2(inbar[102]), .ZN(n496bar);
  OR2_X1 U484 ( .A1(in[123]), .A2(n495), .ZN(n497) );
  AND2_X1 U484bar ( .A1(inbar[123]), .A2(n495bar), .ZN(n497bar);
  OR2_X1 U485 ( .A1(in[143]), .A2(in[130]), .ZN(n495) );
  AND2_X1 U485bar ( .A1(inbar[143]), .A2(inbar[130]), .ZN(n495bar);
  OR2_X1 U486 ( .A1(n494), .A2(n493), .ZN(n605) );
  AND2_X1 U486bar ( .A1(n494bar), .A2(n493bar), .ZN(n605bar);
  OR2_X1 U487 ( .A1(n492), .A2(n491), .ZN(n493) );
  AND2_X1 U487bar ( .A1(n492bar), .A2(n491bar), .ZN(n493bar);
  OR2_X1 U488 ( .A1(in[216]), .A2(in[213]), .ZN(n491) );
  AND2_X1 U488bar ( .A1(inbar[216]), .A2(inbar[213]), .ZN(n491bar);
  OR2_X1 U489 ( .A1(in[227]), .A2(n490), .ZN(n492) );
  AND2_X1 U489bar ( .A1(inbar[227]), .A2(n490bar), .ZN(n492bar);
  OR2_X1 U490 ( .A1(in_0), .A2(in[248]), .ZN(n490) );
  AND2_X1 U490bar ( .A1(in_0bar), .A2(inbar[248]), .ZN(n490bar);
  OR2_X1 U491 ( .A1(n489), .A2(n488), .ZN(n494) );
  AND2_X1 U491bar ( .A1(n489bar), .A2(n488bar), .ZN(n494bar);
  OR2_X1 U492 ( .A1(in_46), .A2(in_44), .ZN(n488) );
  AND2_X1 U492bar ( .A1(in_46bar), .A2(in_44bar), .ZN(n488bar);
  OR2_X1 U493 ( .A1(in_50), .A2(n487), .ZN(n489) );
  AND2_X1 U493bar ( .A1(in_50bar), .A2(n487bar), .ZN(n489bar);
  OR2_X1 U494 ( .A1(in_9), .A2(in_80), .ZN(n487) );
  AND2_X1 U494bar ( .A1(in_9bar), .A2(in_80bar), .ZN(n487bar);
endmodule




module sBox_18 ( in, out );
  input [7:0] in;
  //input_done

  output [7:0] out;
  //output_done

  wire   [255:0] decodeOut;
  //wire_done

  decode_18 dec ( .in(in), .out(decodeOut) );
  encode_18 enc ( .in(decodeOut), .out(out) );
endmodule


module CD2_73 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_74 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_75 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD2_76 ( a, b, y );
  input a, b;
  assign abar = ~a;
  assign bbar = ~b;
  //input_done

  output [3:0] y;
  reg [3:0] ybar;
  //output_done
  
  wire   n3, n4;
  wire n3bar, n4bar;
  //wire_done

  assign n4bar = a;
  assign n4 = abar;
  assign n3bar = b;
  assign n3 = bbar;
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(y[3]) );
  OR2_X1 U3bar ( .A1(bbar), .A2(abar), .ZN(ybar[3]);
  AND2_X1 U4 ( .A1(a), .A2(n3), .ZN(y[2]) );
  OR2_X1 U4bar ( .A1(abar), .A2(n3bar), .ZN(ybar[2]);
  AND2_X1 U5 ( .A1(b), .A2(n4), .ZN(y[1]) );
  OR2_X1 U5bar ( .A1(bbar), .A2(n4bar), .ZN(ybar[1]);
  AND2_X1 U6 ( .A1(n4), .A2(n3), .ZN(y[0]) );
  OR2_X1 U6bar ( .A1(n4bar), .A2(n3bar), .ZN(ybar[0]);
endmodule




module CD4_37 ( a, b, y );
  input [3:0] a;
  input [3:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  //input_done

  output [15:0] y;
  reg [15:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]);
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]);
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]);
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]);
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]);
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]);
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]);
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]);
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]);
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]);
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]);
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]);
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]);
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]);
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]);
endmodule




module CD4_38 ( a, b, y );
  input [3:0] a;
  input [3:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  //input_done

  output [15:0] y;
  reg [15:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[1]), .A2(a[2]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[1]), .A2(abar[2]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[0]), .A2(a[2]), .ZN(y[8]) );
  OR2_X1 U2bar ( .A1(bbar[0]), .A2(abar[2]), .ZN(ybar[8]);
  AND2_X1 U3 ( .A1(b[3]), .A2(a[1]), .ZN(y[7]) );
  OR2_X1 U3bar ( .A1(bbar[3]), .A2(abar[1]), .ZN(ybar[7]);
  AND2_X1 U4 ( .A1(b[2]), .A2(a[1]), .ZN(y[6]) );
  OR2_X1 U4bar ( .A1(bbar[2]), .A2(abar[1]), .ZN(ybar[6]);
  AND2_X1 U5 ( .A1(a[1]), .A2(b[1]), .ZN(y[5]) );
  OR2_X1 U5bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[5]);
  AND2_X1 U6 ( .A1(a[1]), .A2(b[0]), .ZN(y[4]) );
  OR2_X1 U6bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[4]);
  AND2_X1 U7 ( .A1(a[0]), .A2(b[3]), .ZN(y[3]) );
  OR2_X1 U7bar ( .A1(abar[0]), .A2(bbar[3]), .ZN(ybar[3]);
  AND2_X1 U8 ( .A1(a[0]), .A2(b[2]), .ZN(y[2]) );
  OR2_X1 U8bar ( .A1(abar[0]), .A2(bbar[2]), .ZN(ybar[2]);
  AND2_X1 U9 ( .A1(a[0]), .A2(b[1]), .ZN(y[1]) );
  OR2_X1 U9bar ( .A1(abar[0]), .A2(bbar[1]), .ZN(ybar[1]);
  AND2_X1 U10 ( .A1(a[3]), .A2(b[3]), .ZN(y[15]) );
  OR2_X1 U10bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[15]);
  AND2_X1 U11 ( .A1(a[3]), .A2(b[2]), .ZN(y[14]) );
  OR2_X1 U11bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[14]);
  AND2_X1 U12 ( .A1(a[3]), .A2(b[1]), .ZN(y[13]) );
  OR2_X1 U12bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[13]);
  AND2_X1 U13 ( .A1(a[3]), .A2(b[0]), .ZN(y[12]) );
  OR2_X1 U13bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[12]);
  AND2_X1 U14 ( .A1(b[3]), .A2(a[2]), .ZN(y[11]) );
  OR2_X1 U14bar ( .A1(bbar[3]), .A2(abar[2]), .ZN(ybar[11]);
  AND2_X1 U15 ( .A1(b[2]), .A2(a[2]), .ZN(y[10]) );
  OR2_X1 U15bar ( .A1(bbar[2]), .A2(abar[2]), .ZN(ybar[10]);
  AND2_X1 U16 ( .A1(a[0]), .A2(b[0]), .ZN(y[0]) );
  OR2_X1 U16bar ( .A1(abar[0]), .A2(bbar[0]), .ZN(ybar[0]);
endmodule




module CD16_19 ( a, b, y );
  input [15:0] a;
  input [15:0] b;
  assign abar[0] = ~a[0];
  assign abar[1] = ~a[1];
  assign abar[2] = ~a[2];
  assign abar[3] = ~a[3];
  assign abar[4] = ~a[4];
  assign abar[5] = ~a[5];
  assign abar[6] = ~a[6];
  assign abar[7] = ~a[7];
  assign abar[8] = ~a[8];
  assign abar[9] = ~a[9];
  assign abar[10] = ~a[10];
  assign abar[11] = ~a[11];
  assign abar[12] = ~a[12];
  assign abar[13] = ~a[13];
  assign abar[14] = ~a[14];
  assign abar[15] = ~a[15];
  assign bbar[0] = ~b[0];
  assign bbar[1] = ~b[1];
  assign bbar[2] = ~b[2];
  assign bbar[3] = ~b[3];
  assign bbar[4] = ~b[4];
  assign bbar[5] = ~b[5];
  assign bbar[6] = ~b[6];
  assign bbar[7] = ~b[7];
  assign bbar[8] = ~b[8];
  assign bbar[9] = ~b[9];
  assign bbar[10] = ~b[10];
  assign bbar[11] = ~b[11];
  assign bbar[12] = ~b[12];
  assign bbar[13] = ~b[13];
  assign bbar[14] = ~b[14];
  assign bbar[15] = ~b[15];
  //input_done

  output [15:0] y;
  reg [15:0] ybar;
  //output_done



  AND2_X1 U1 ( .A1(b[9]), .A2(a[0]), .ZN(y[9]) );
  OR2_X1 U1bar ( .A1(bbar[9]), .A2(abar[0]), .ZN(ybar[9]);
  AND2_X1 U2 ( .A1(b[3]), .A2(a[6]), .ZN(y[99]) );
  OR2_X1 U2bar ( .A1(bbar[3]), .A2(abar[6]), .ZN(ybar[99]);
  AND2_X1 U3 ( .A1(b[2]), .A2(a[6]), .ZN(y[98]) );
  OR2_X1 U3bar ( .A1(bbar[2]), .A2(abar[6]), .ZN(ybar[98]);
  AND2_X1 U4 ( .A1(b[1]), .A2(a[6]), .ZN(y[97]) );
  OR2_X1 U4bar ( .A1(bbar[1]), .A2(abar[6]), .ZN(ybar[97]);
  AND2_X1 U5 ( .A1(b[0]), .A2(a[6]), .ZN(y[96]) );
  OR2_X1 U5bar ( .A1(bbar[0]), .A2(abar[6]), .ZN(ybar[96]);
  AND2_X1 U6 ( .A1(b[15]), .A2(a[5]), .ZN(y[95]) );
  OR2_X1 U6bar ( .A1(bbar[15]), .A2(abar[5]), .ZN(ybar[95]);
  AND2_X1 U7 ( .A1(b[14]), .A2(a[5]), .ZN(y[94]) );
  OR2_X1 U7bar ( .A1(bbar[14]), .A2(abar[5]), .ZN(ybar[94]);
  AND2_X1 U8 ( .A1(b[13]), .A2(a[5]), .ZN(y[93]) );
  OR2_X1 U8bar ( .A1(bbar[13]), .A2(abar[5]), .ZN(ybar[93]);
  AND2_X1 U9 ( .A1(b[12]), .A2(a[5]), .ZN(y[92]) );
  OR2_X1 U9bar ( .A1(bbar[12]), .A2(abar[5]), .ZN(ybar[92]);
  AND2_X1 U10 ( .A1(b[11]), .A2(a[5]), .ZN(y[91]) );
  OR2_X1 U10bar ( .A1(bbar[11]), .A2(abar[5]), .ZN(ybar[91]);
  AND2_X1 U11 ( .A1(b[10]), .A2(a[5]), .ZN(y[90]) );
  OR2_X1 U11bar ( .A1(bbar[10]), .A2(abar[5]), .ZN(ybar[90]);
  AND2_X1 U12 ( .A1(b[8]), .A2(a[0]), .ZN(y[8]) );
  OR2_X1 U12bar ( .A1(bbar[8]), .A2(abar[0]), .ZN(ybar[8]);
  AND2_X1 U13 ( .A1(a[5]), .A2(b[9]), .ZN(y[89]) );
  OR2_X1 U13bar ( .A1(abar[5]), .A2(bbar[9]), .ZN(ybar[89]);
  AND2_X1 U14 ( .A1(b[8]), .A2(a[5]), .ZN(y[88]) );
  OR2_X1 U14bar ( .A1(bbar[8]), .A2(abar[5]), .ZN(ybar[88]);
  AND2_X1 U15 ( .A1(b[7]), .A2(a[5]), .ZN(y[87]) );
  OR2_X1 U15bar ( .A1(bbar[7]), .A2(abar[5]), .ZN(ybar[87]);
  AND2_X1 U16 ( .A1(b[6]), .A2(a[5]), .ZN(y[86]) );
  OR2_X1 U16bar ( .A1(bbar[6]), .A2(abar[5]), .ZN(ybar[86]);
  AND2_X1 U17 ( .A1(b[5]), .A2(a[5]), .ZN(y[85]) );
  OR2_X1 U17bar ( .A1(bbar[5]), .A2(abar[5]), .ZN(ybar[85]);
  AND2_X1 U18 ( .A1(b[4]), .A2(a[5]), .ZN(y[84]) );
  OR2_X1 U18bar ( .A1(bbar[4]), .A2(abar[5]), .ZN(ybar[84]);
  AND2_X1 U19 ( .A1(a[5]), .A2(b[3]), .ZN(y[83]) );
  OR2_X1 U19bar ( .A1(abar[5]), .A2(bbar[3]), .ZN(ybar[83]);
  AND2_X1 U20 ( .A1(a[5]), .A2(b[2]), .ZN(y[82]) );
  OR2_X1 U20bar ( .A1(abar[5]), .A2(bbar[2]), .ZN(ybar[82]);
  AND2_X1 U21 ( .A1(a[5]), .A2(b[1]), .ZN(y[81]) );
  OR2_X1 U21bar ( .A1(abar[5]), .A2(bbar[1]), .ZN(ybar[81]);
  AND2_X1 U22 ( .A1(a[5]), .A2(b[0]), .ZN(y[80]) );
  OR2_X1 U22bar ( .A1(abar[5]), .A2(bbar[0]), .ZN(ybar[80]);
  AND2_X1 U23 ( .A1(b[7]), .A2(a[0]), .ZN(y[7]) );
  OR2_X1 U23bar ( .A1(bbar[7]), .A2(abar[0]), .ZN(ybar[7]);
  AND2_X1 U24 ( .A1(a[4]), .A2(b[15]), .ZN(y[79]) );
  OR2_X1 U24bar ( .A1(abar[4]), .A2(bbar[15]), .ZN(ybar[79]);
  AND2_X1 U25 ( .A1(a[4]), .A2(b[14]), .ZN(y[78]) );
  OR2_X1 U25bar ( .A1(abar[4]), .A2(bbar[14]), .ZN(ybar[78]);
  AND2_X1 U26 ( .A1(a[4]), .A2(b[13]), .ZN(y[77]) );
  OR2_X1 U26bar ( .A1(abar[4]), .A2(bbar[13]), .ZN(ybar[77]);
  AND2_X1 U27 ( .A1(a[4]), .A2(b[12]), .ZN(y[76]) );
  OR2_X1 U27bar ( .A1(abar[4]), .A2(bbar[12]), .ZN(ybar[76]);
  AND2_X1 U28 ( .A1(a[4]), .A2(b[11]), .ZN(y[75]) );
  OR2_X1 U28bar ( .A1(abar[4]), .A2(bbar[11]), .ZN(ybar[75]);
  AND2_X1 U29 ( .A1(a[4]), .A2(b[10]), .ZN(y[74]) );
  OR2_X1 U29bar ( .A1(abar[4]), .A2(bbar[10]), .ZN(ybar[74]);
  AND2_X1 U30 ( .A1(a[4]), .A2(b[9]), .ZN(y[73]) );
  OR2_X1 U30bar ( .A1(abar[4]), .A2(bbar[9]), .ZN(ybar[73]);
  AND2_X1 U31 ( .A1(a[4]), .A2(b[8]), .ZN(y[72]) );
  OR2_X1 U31bar ( .A1(abar[4]), .A2(bbar[8]), .ZN(ybar[72]);
  AND2_X1 U32 ( .A1(a[4]), .A2(b[7]), .ZN(y[71]) );
  OR2_X1 U32bar ( .A1(abar[4]), .A2(bbar[7]), .ZN(ybar[71]);
  AND2_X1 U33 ( .A1(a[4]), .A2(b[6]), .ZN(y[70]) );
  OR2_X1 U33bar ( .A1(abar[4]), .A2(bbar[6]), .ZN(ybar[70]);
  AND2_X1 U34 ( .A1(b[6]), .A2(a[0]), .ZN(y[6]) );
  OR2_X1 U34bar ( .A1(bbar[6]), .A2(abar[0]), .ZN(ybar[6]);
  AND2_X1 U35 ( .A1(a[4]), .A2(b[5]), .ZN(y[69]) );
  OR2_X1 U35bar ( .A1(abar[4]), .A2(bbar[5]), .ZN(ybar[69]);
  AND2_X1 U36 ( .A1(a[4]), .A2(b[4]), .ZN(y[68]) );
  OR2_X1 U36bar ( .A1(abar[4]), .A2(bbar[4]), .ZN(ybar[68]);
  AND2_X1 U37 ( .A1(a[4]), .A2(b[3]), .ZN(y[67]) );
  OR2_X1 U37bar ( .A1(abar[4]), .A2(bbar[3]), .ZN(ybar[67]);
  AND2_X1 U38 ( .A1(a[4]), .A2(b[2]), .ZN(y[66]) );
  OR2_X1 U38bar ( .A1(abar[4]), .A2(bbar[2]), .ZN(ybar[66]);
  AND2_X1 U39 ( .A1(a[4]), .A2(b[1]), .ZN(y[65]) );
  OR2_X1 U39bar ( .A1(abar[4]), .A2(bbar[1]), .ZN(ybar[65]);
  AND2_X1 U40 ( .A1(a[4]), .A2(b[0]), .ZN(y[64]) );
  OR2_X1 U40bar ( .A1(abar[4]), .A2(bbar[0]), .ZN(ybar[64]);
  AND2_X1 U41 ( .A1(a[3]), .A2(b[15]), .ZN(y[63]) );
  OR2_X1 U41bar ( .A1(abar[3]), .A2(bbar[15]), .ZN(ybar[63]);
  AND2_X1 U42 ( .A1(a[3]), .A2(b[14]), .ZN(y[62]) );
  OR2_X1 U42bar ( .A1(abar[3]), .A2(bbar[14]), .ZN(ybar[62]);
  AND2_X1 U43 ( .A1(a[3]), .A2(b[13]), .ZN(y[61]) );
  OR2_X1 U43bar ( .A1(abar[3]), .A2(bbar[13]), .ZN(ybar[61]);
  AND2_X1 U44 ( .A1(a[3]), .A2(b[12]), .ZN(y[60]) );
  OR2_X1 U44bar ( .A1(abar[3]), .A2(bbar[12]), .ZN(ybar[60]);
  AND2_X1 U45 ( .A1(b[5]), .A2(a[0]), .ZN(y[5]) );
  OR2_X1 U45bar ( .A1(bbar[5]), .A2(abar[0]), .ZN(ybar[5]);
  AND2_X1 U46 ( .A1(a[3]), .A2(b[11]), .ZN(y[59]) );
  OR2_X1 U46bar ( .A1(abar[3]), .A2(bbar[11]), .ZN(ybar[59]);
  AND2_X1 U47 ( .A1(a[3]), .A2(b[10]), .ZN(y[58]) );
  OR2_X1 U47bar ( .A1(abar[3]), .A2(bbar[10]), .ZN(ybar[58]);
  AND2_X1 U48 ( .A1(a[3]), .A2(b[9]), .ZN(y[57]) );
  OR2_X1 U48bar ( .A1(abar[3]), .A2(bbar[9]), .ZN(ybar[57]);
  AND2_X1 U49 ( .A1(a[3]), .A2(b[8]), .ZN(y[56]) );
  OR2_X1 U49bar ( .A1(abar[3]), .A2(bbar[8]), .ZN(ybar[56]);
  AND2_X1 U50 ( .A1(a[3]), .A2(b[7]), .ZN(y[55]) );
  OR2_X1 U50bar ( .A1(abar[3]), .A2(bbar[7]), .ZN(ybar[55]);
  AND2_X1 U51 ( .A1(a[3]), .A2(b[6]), .ZN(y[54]) );
  OR2_X1 U51bar ( .A1(abar[3]), .A2(bbar[6]), .ZN(ybar[54]);
  AND2_X1 U52 ( .A1(a[3]), .A2(b[5]), .ZN(y[53]) );
  OR2_X1 U52bar ( .A1(abar[3]), .A2(bbar[5]), .ZN(ybar[53]);
  AND2_X1 U53 ( .A1(a[3]), .A2(b[4]), .ZN(y[52]) );
  OR2_X1 U53bar ( .A1(abar[3]), .A2(bbar[4]), .ZN(ybar[52]);
  AND2_X1 U54 ( .A1(a[3]), .A2(b[3]), .ZN(y[51]) );
  OR2_X1 U54bar ( .A1(abar[3]), .A2(bbar[3]), .ZN(ybar[51]);
  AND2_X1 U55 ( .A1(a[3]), .A2(b[2]), .ZN(y[50]) );
  OR2_X1 U55bar ( .A1(abar[3]), .A2(bbar[2]), .ZN(ybar[50]);
  AND2_X1 U56 ( .A1(b[4]), .A2(a[0]), .ZN(y[4]) );
  OR2_X1 U56bar ( .A1(bbar[4]), .A2(abar[0]), .ZN(ybar[4]);
  AND2_X1 U57 ( .A1(a[3]), .A2(b[1]), .ZN(y[49]) );
  OR2_X1 U57bar ( .A1(abar[3]), .A2(bbar[1]), .ZN(ybar[49]);
  AND2_X1 U58 ( .A1(a[3]), .A2(b[0]), .ZN(y[48]) );
  OR2_X1 U58bar ( .A1(abar[3]), .A2(bbar[0]), .ZN(ybar[48]);
  AND2_X1 U59 ( .A1(a[2]), .A2(b[15]), .ZN(y[47]) );
  OR2_X1 U59bar ( .A1(abar[2]), .A2(bbar[15]), .ZN(ybar[47]);
  AND2_X1 U60 ( .A1(a[2]), .A2(b[14]), .ZN(y[46]) );
  OR2_X1 U60bar ( .A1(abar[2]), .A2(bbar[14]), .ZN(ybar[46]);
  AND2_X1 U61 ( .A1(a[2]), .A2(b[13]), .ZN(y[45]) );
  OR2_X1 U61bar ( .A1(abar[2]), .A2(bbar[13]), .ZN(ybar[45]);
  AND2_X1 U62 ( .A1(a[2]), .A2(b[12]), .ZN(y[44]) );
  OR2_X1 U62bar ( .A1(abar[2]), .A2(bbar[12]), .ZN(ybar[44]);
  AND2_X1 U63 ( .A1(a[2]), .A2(b[11]), .ZN(y[43]) );
  OR2_X1 U63bar ( .A1(abar[2]), .A2(bbar[11]), .ZN(ybar[43]);
  AND2_X1 U64 ( .A1(a[2]), .A2(b[10]), .ZN(y[42]) );
  OR2_X1 U64bar ( .A1(abar[2]), .A2(bbar[10]), .ZN(ybar[42]);
  AND2_X1 U65 ( .A1(a[2]), .A2(b[9]), .ZN(y[41]) );
  OR2_X1 U65bar ( .A1(abar[2]), .A2(bbar[9]), .ZN(ybar[41]);
  AND2_X1 U66 ( .A1(a[2]), .A2(b[8]), .ZN(y[40]) );
  OR2_X1 U66bar ( .A1(abar[2]), .A2(bbar[8]), .ZN(ybar[40]);
  AND2_X1 U67 ( .A1(b[3]), .A2(a[0]), .ZN(y[3]) );
  OR2_X1 U67bar ( .A1(bbar[3]), .A2(abar[0]), .ZN(ybar[3]);
  AND2_X1 U68 ( .A1(a[2]), .A2(b[7]), .ZN(y[39]) );
  OR2_X1 U68bar ( .A1(abar[2]), .A2(bbar[7]), .ZN(ybar[39]);
  AND2_X1 U69 ( .A1(a[2]), .A2(b[6]), .ZN(y[38]) );
  OR2_X1 U69bar ( .A1(abar[2]), .A2(bbar[6]), .ZN(ybar[38]);
  AND2_X1 U70 ( .A1(a[2]), .A2(b[5]), .ZN(y[37]) );
  OR2_X1 U70bar ( .A1(abar[2]), .A2(bbar[5]), .ZN(ybar[37]);
  AND2_X1 U71 ( .A1(a[2]), .A2(b[4]), .ZN(y[36]) );
  OR2_X1 U71bar ( .A1(abar[2]), .A2(bbar[4]), .ZN(ybar[36]);
  AND2_X1 U72 ( .A1(a[2]), .A2(b[3]), .ZN(y[35]) );
  OR2_X1 U72bar ( .A1(abar[2]), .A2(bbar[3]), .ZN(ybar[35]);
  AND2_X1 U73 ( .A1(a[2]), .A2(b[2]), .ZN(y[34]) );
  OR2_X1 U73bar ( .A1(abar[2]), .A2(bbar[2]), .ZN(ybar[34]);
  AND2_X1 U74 ( .A1(a[2]), .A2(b[1]), .ZN(y[33]) );
  OR2_X1 U74bar ( .A1(abar[2]), .A2(bbar[1]), .ZN(ybar[33]);
  AND2_X1 U75 ( .A1(a[2]), .A2(b[0]), .ZN(y[32]) );
  OR2_X1 U75bar ( .A1(abar[2]), .A2(bbar[0]), .ZN(ybar[32]);
  AND2_X1 U76 ( .A1(a[1]), .A2(b[15]), .ZN(y[31]) );
  OR2_X1 U76bar ( .A1(abar[1]), .A2(bbar[15]), .ZN(ybar[31]);
  AND2_X1 U77 ( .A1(a[1]), .A2(b[14]), .ZN(y[30]) );
  OR2_X1 U77bar ( .A1(abar[1]), .A2(bbar[14]), .ZN(ybar[30]);
  AND2_X1 U78 ( .A1(b[2]), .A2(a[0]), .ZN(y[2]) );
  OR2_X1 U78bar ( .A1(bbar[2]), .A2(abar[0]), .ZN(ybar[2]);
  AND2_X1 U79 ( .A1(a[1]), .A2(b[13]), .ZN(y[29]) );
  OR2_X1 U79bar ( .A1(abar[1]), .A2(bbar[13]), .ZN(ybar[29]);
  AND2_X1 U80 ( .A1(a[1]), .A2(b[12]), .ZN(y[28]) );
  OR2_X1 U80bar ( .A1(abar[1]), .A2(bbar[12]), .ZN(ybar[28]);
  AND2_X1 U81 ( .A1(a[1]), .A2(b[11]), .ZN(y[27]) );
  OR2_X1 U81bar ( .A1(abar[1]), .A2(bbar[11]), .ZN(ybar[27]);
  AND2_X1 U82 ( .A1(a[1]), .A2(b[10]), .ZN(y[26]) );
  OR2_X1 U82bar ( .A1(abar[1]), .A2(bbar[10]), .ZN(ybar[26]);
  AND2_X1 U83 ( .A1(a[1]), .A2(b[9]), .ZN(y[25]) );
  OR2_X1 U83bar ( .A1(abar[1]), .A2(bbar[9]), .ZN(ybar[25]);
  AND2_X1 U84 ( .A1(a[15]), .A2(b[15]), .ZN(y[255]) );
  OR2_X1 U84bar ( .A1(abar[15]), .A2(bbar[15]), .ZN(ybar[255]);
  AND2_X1 U85 ( .A1(a[15]), .A2(b[14]), .ZN(y[254]) );
  OR2_X1 U85bar ( .A1(abar[15]), .A2(bbar[14]), .ZN(ybar[254]);
  AND2_X1 U86 ( .A1(a[15]), .A2(b[13]), .ZN(y[253]) );
  OR2_X1 U86bar ( .A1(abar[15]), .A2(bbar[13]), .ZN(ybar[253]);
  AND2_X1 U87 ( .A1(a[15]), .A2(b[12]), .ZN(y[252]) );
  OR2_X1 U87bar ( .A1(abar[15]), .A2(bbar[12]), .ZN(ybar[252]);
  AND2_X1 U88 ( .A1(a[15]), .A2(b[11]), .ZN(y[251]) );
  OR2_X1 U88bar ( .A1(abar[15]), .A2(bbar[11]), .ZN(ybar[251]);
  AND2_X1 U89 ( .A1(a[15]), .A2(b[10]), .ZN(y[250]) );
  OR2_X1 U89bar ( .A1(abar[15]), .A2(bbar[10]), .ZN(ybar[250]);
  AND2_X1 U90 ( .A1(a[1]), .A2(b[8]), .ZN(y[24]) );
  OR2_X1 U90bar ( .A1(abar[1]), .A2(bbar[8]), .ZN(ybar[24]);
  AND2_X1 U91 ( .A1(a[15]), .A2(b[9]), .ZN(y[249]) );
  OR2_X1 U91bar ( .A1(abar[15]), .A2(bbar[9]), .ZN(ybar[249]);
  AND2_X1 U92 ( .A1(a[15]), .A2(b[8]), .ZN(y[248]) );
  OR2_X1 U92bar ( .A1(abar[15]), .A2(bbar[8]), .ZN(ybar[248]);
  AND2_X1 U93 ( .A1(a[15]), .A2(b[7]), .ZN(y[247]) );
  OR2_X1 U93bar ( .A1(abar[15]), .A2(bbar[7]), .ZN(ybar[247]);
  AND2_X1 U94 ( .A1(a[15]), .A2(b[6]), .ZN(y[246]) );
  OR2_X1 U94bar ( .A1(abar[15]), .A2(bbar[6]), .ZN(ybar[246]);
  AND2_X1 U95 ( .A1(a[15]), .A2(b[5]), .ZN(y[245]) );
  OR2_X1 U95bar ( .A1(abar[15]), .A2(bbar[5]), .ZN(ybar[245]);
  AND2_X1 U96 ( .A1(a[15]), .A2(b[4]), .ZN(y[244]) );
  OR2_X1 U96bar ( .A1(abar[15]), .A2(bbar[4]), .ZN(ybar[244]);
  AND2_X1 U97 ( .A1(a[15]), .A2(b[3]), .ZN(y[243]) );
  OR2_X1 U97bar ( .A1(abar[15]), .A2(bbar[3]), .ZN(ybar[243]);
  AND2_X1 U98 ( .A1(a[15]), .A2(b[2]), .ZN(y[242]) );
  OR2_X1 U98bar ( .A1(abar[15]), .A2(bbar[2]), .ZN(ybar[242]);
  AND2_X1 U99 ( .A1(a[15]), .A2(b[1]), .ZN(y[241]) );
  OR2_X1 U99bar ( .A1(abar[15]), .A2(bbar[1]), .ZN(ybar[241]);
  AND2_X1 U100 ( .A1(a[15]), .A2(b[0]), .ZN(y[240]) );
  OR2_X1 U100bar ( .A1(abar[15]), .A2(bbar[0]), .ZN(ybar[240]);
  AND2_X1 U101 ( .A1(a[1]), .A2(b[7]), .ZN(y[23]) );
  OR2_X1 U101bar ( .A1(abar[1]), .A2(bbar[7]), .ZN(ybar[23]);
  AND2_X1 U102 ( .A1(a[14]), .A2(b[15]), .ZN(y[239]) );
  OR2_X1 U102bar ( .A1(abar[14]), .A2(bbar[15]), .ZN(ybar[239]);
  AND2_X1 U103 ( .A1(a[14]), .A2(b[14]), .ZN(y[238]) );
  OR2_X1 U103bar ( .A1(abar[14]), .A2(bbar[14]), .ZN(ybar[238]);
  AND2_X1 U104 ( .A1(a[14]), .A2(b[13]), .ZN(y[237]) );
  OR2_X1 U104bar ( .A1(abar[14]), .A2(bbar[13]), .ZN(ybar[237]);
  AND2_X1 U105 ( .A1(a[14]), .A2(b[12]), .ZN(y[236]) );
  OR2_X1 U105bar ( .A1(abar[14]), .A2(bbar[12]), .ZN(ybar[236]);
  AND2_X1 U106 ( .A1(a[14]), .A2(b[11]), .ZN(y[235]) );
  OR2_X1 U106bar ( .A1(abar[14]), .A2(bbar[11]), .ZN(ybar[235]);
  AND2_X1 U107 ( .A1(a[14]), .A2(b[10]), .ZN(y[234]) );
  OR2_X1 U107bar ( .A1(abar[14]), .A2(bbar[10]), .ZN(ybar[234]);
  AND2_X1 U108 ( .A1(a[14]), .A2(b[9]), .ZN(y[233]) );
  OR2_X1 U108bar ( .A1(abar[14]), .A2(bbar[9]), .ZN(ybar[233]);
  AND2_X1 U109 ( .A1(a[14]), .A2(b[8]), .ZN(y[232]) );
  OR2_X1 U109bar ( .A1(abar[14]), .A2(bbar[8]), .ZN(ybar[232]);
  AND2_X1 U110 ( .A1(a[14]), .A2(b[7]), .ZN(y[231]) );
  OR2_X1 U110bar ( .A1(abar[14]), .A2(bbar[7]), .ZN(ybar[231]);
  AND2_X1 U111 ( .A1(a[14]), .A2(b[6]), .ZN(y[230]) );
  OR2_X1 U111bar ( .A1(abar[14]), .A2(bbar[6]), .ZN(ybar[230]);
  AND2_X1 U112 ( .A1(a[1]), .A2(b[6]), .ZN(y[22]) );
  OR2_X1 U112bar ( .A1(abar[1]), .A2(bbar[6]), .ZN(ybar[22]);
  AND2_X1 U113 ( .A1(a[14]), .A2(b[5]), .ZN(y[229]) );
  OR2_X1 U113bar ( .A1(abar[14]), .A2(bbar[5]), .ZN(ybar[229]);
  AND2_X1 U114 ( .A1(a[14]), .A2(b[4]), .ZN(y[228]) );
  OR2_X1 U114bar ( .A1(abar[14]), .A2(bbar[4]), .ZN(ybar[228]);
  AND2_X1 U115 ( .A1(a[14]), .A2(b[3]), .ZN(y[227]) );
  OR2_X1 U115bar ( .A1(abar[14]), .A2(bbar[3]), .ZN(ybar[227]);
  AND2_X1 U116 ( .A1(a[14]), .A2(b[2]), .ZN(y[226]) );
  OR2_X1 U116bar ( .A1(abar[14]), .A2(bbar[2]), .ZN(ybar[226]);
  AND2_X1 U117 ( .A1(a[14]), .A2(b[1]), .ZN(y[225]) );
  OR2_X1 U117bar ( .A1(abar[14]), .A2(bbar[1]), .ZN(ybar[225]);
  AND2_X1 U118 ( .A1(a[14]), .A2(b[0]), .ZN(y[224]) );
  OR2_X1 U118bar ( .A1(abar[14]), .A2(bbar[0]), .ZN(ybar[224]);
  AND2_X1 U119 ( .A1(a[13]), .A2(b[15]), .ZN(y[223]) );
  OR2_X1 U119bar ( .A1(abar[13]), .A2(bbar[15]), .ZN(ybar[223]);
  AND2_X1 U120 ( .A1(a[13]), .A2(b[14]), .ZN(y[222]) );
  OR2_X1 U120bar ( .A1(abar[13]), .A2(bbar[14]), .ZN(ybar[222]);
  AND2_X1 U121 ( .A1(a[13]), .A2(b[13]), .ZN(y[221]) );
  OR2_X1 U121bar ( .A1(abar[13]), .A2(bbar[13]), .ZN(ybar[221]);
  AND2_X1 U122 ( .A1(a[13]), .A2(b[12]), .ZN(y[220]) );
  OR2_X1 U122bar ( .A1(abar[13]), .A2(bbar[12]), .ZN(ybar[220]);
  AND2_X1 U123 ( .A1(a[1]), .A2(b[5]), .ZN(y[21]) );
  OR2_X1 U123bar ( .A1(abar[1]), .A2(bbar[5]), .ZN(ybar[21]);
  AND2_X1 U124 ( .A1(a[13]), .A2(b[11]), .ZN(y[219]) );
  OR2_X1 U124bar ( .A1(abar[13]), .A2(bbar[11]), .ZN(ybar[219]);
  AND2_X1 U125 ( .A1(a[13]), .A2(b[10]), .ZN(y[218]) );
  OR2_X1 U125bar ( .A1(abar[13]), .A2(bbar[10]), .ZN(ybar[218]);
  AND2_X1 U126 ( .A1(a[13]), .A2(b[9]), .ZN(y[217]) );
  OR2_X1 U126bar ( .A1(abar[13]), .A2(bbar[9]), .ZN(ybar[217]);
  AND2_X1 U127 ( .A1(a[13]), .A2(b[8]), .ZN(y[216]) );
  OR2_X1 U127bar ( .A1(abar[13]), .A2(bbar[8]), .ZN(ybar[216]);
  AND2_X1 U128 ( .A1(a[13]), .A2(b[7]), .ZN(y[215]) );
  OR2_X1 U128bar ( .A1(abar[13]), .A2(bbar[7]), .ZN(ybar[215]);
  AND2_X1 U129 ( .A1(a[13]), .A2(b[6]), .ZN(y[214]) );
  OR2_X1 U129bar ( .A1(abar[13]), .A2(bbar[6]), .ZN(ybar[214]);
  AND2_X1 U130 ( .A1(a[13]), .A2(b[5]), .ZN(y[213]) );
  OR2_X1 U130bar ( .A1(abar[13]), .A2(bbar[5]), .ZN(ybar[213]);
  AND2_X1 U131 ( .A1(a[13]), .A2(b[4]), .ZN(y[212]) );
  OR2_X1 U131bar ( .A1(abar[13]), .A2(bbar[4]), .ZN(ybar[212]);
  AND2_X1 U132 ( .A1(a[13]), .A2(b[3]), .ZN(y[211]) );
  OR2_X1 U132bar ( .A1(abar[13]), .A2(bbar[3]), .ZN(ybar[211]);
  AND2_X1 U133 ( .A1(a[13]), .A2(b[2]), .ZN(y[210]) );
  OR2_X1 U133bar ( .A1(abar[13]), .A2(bbar[2]), .ZN(ybar[210]);
  AND2_X1 U134 ( .A1(a[1]), .A2(b[4]), .ZN(y[20]) );
  OR2_X1 U134bar ( .A1(abar[1]), .A2(bbar[4]), .ZN(ybar[20]);
  AND2_X1 U135 ( .A1(a[13]), .A2(b[1]), .ZN(y[209]) );
  OR2_X1 U135bar ( .A1(abar[13]), .A2(bbar[1]), .ZN(ybar[209]);
  AND2_X1 U136 ( .A1(a[13]), .A2(b[0]), .ZN(y[208]) );
  OR2_X1 U136bar ( .A1(abar[13]), .A2(bbar[0]), .ZN(ybar[208]);
  AND2_X1 U137 ( .A1(a[12]), .A2(b[15]), .ZN(y[207]) );
  OR2_X1 U137bar ( .A1(abar[12]), .A2(bbar[15]), .ZN(ybar[207]);
  AND2_X1 U138 ( .A1(a[12]), .A2(b[14]), .ZN(y[206]) );
  OR2_X1 U138bar ( .A1(abar[12]), .A2(bbar[14]), .ZN(ybar[206]);
  AND2_X1 U139 ( .A1(a[12]), .A2(b[13]), .ZN(y[205]) );
  OR2_X1 U139bar ( .A1(abar[12]), .A2(bbar[13]), .ZN(ybar[205]);
  AND2_X1 U140 ( .A1(a[12]), .A2(b[12]), .ZN(y[204]) );
  OR2_X1 U140bar ( .A1(abar[12]), .A2(bbar[12]), .ZN(ybar[204]);
  AND2_X1 U141 ( .A1(a[12]), .A2(b[11]), .ZN(y[203]) );
  OR2_X1 U141bar ( .A1(abar[12]), .A2(bbar[11]), .ZN(ybar[203]);
  AND2_X1 U142 ( .A1(a[12]), .A2(b[10]), .ZN(y[202]) );
  OR2_X1 U142bar ( .A1(abar[12]), .A2(bbar[10]), .ZN(ybar[202]);
  AND2_X1 U143 ( .A1(a[12]), .A2(b[9]), .ZN(y[201]) );
  OR2_X1 U143bar ( .A1(abar[12]), .A2(bbar[9]), .ZN(ybar[201]);
  AND2_X1 U144 ( .A1(a[12]), .A2(b[8]), .ZN(y[200]) );
  OR2_X1 U144bar ( .A1(abar[12]), .A2(bbar[8]), .ZN(ybar[200]);
  AND2_X1 U145 ( .A1(b[1]), .A2(a[0]), .ZN(y[1]) );
  OR2_X1 U145bar ( .A1(bbar[1]), .A2(abar[0]), .ZN(ybar[1]);
  AND2_X1 U146 ( .A1(a[1]), .A2(b[3]), .ZN(y[19]) );
  OR2_X1 U146bar ( .A1(abar[1]), .A2(bbar[3]), .ZN(ybar[19]);
  AND2_X1 U147 ( .A1(a[12]), .A2(b[7]), .ZN(y[199]) );
  OR2_X1 U147bar ( .A1(abar[12]), .A2(bbar[7]), .ZN(ybar[199]);
  AND2_X1 U148 ( .A1(a[12]), .A2(b[6]), .ZN(y[198]) );
  OR2_X1 U148bar ( .A1(abar[12]), .A2(bbar[6]), .ZN(ybar[198]);
  AND2_X1 U149 ( .A1(a[12]), .A2(b[5]), .ZN(y[197]) );
  OR2_X1 U149bar ( .A1(abar[12]), .A2(bbar[5]), .ZN(ybar[197]);
  AND2_X1 U150 ( .A1(a[12]), .A2(b[4]), .ZN(y[196]) );
  OR2_X1 U150bar ( .A1(abar[12]), .A2(bbar[4]), .ZN(ybar[196]);
  AND2_X1 U151 ( .A1(a[12]), .A2(b[3]), .ZN(y[195]) );
  OR2_X1 U151bar ( .A1(abar[12]), .A2(bbar[3]), .ZN(ybar[195]);
  AND2_X1 U152 ( .A1(a[12]), .A2(b[2]), .ZN(y[194]) );
  OR2_X1 U152bar ( .A1(abar[12]), .A2(bbar[2]), .ZN(ybar[194]);
  AND2_X1 U153 ( .A1(a[12]), .A2(b[1]), .ZN(y[193]) );
  OR2_X1 U153bar ( .A1(abar[12]), .A2(bbar[1]), .ZN(ybar[193]);
  AND2_X1 U154 ( .A1(a[12]), .A2(b[0]), .ZN(y[192]) );
  OR2_X1 U154bar ( .A1(abar[12]), .A2(bbar[0]), .ZN(ybar[192]);
  AND2_X1 U155 ( .A1(a[11]), .A2(b[15]), .ZN(y[191]) );
  OR2_X1 U155bar ( .A1(abar[11]), .A2(bbar[15]), .ZN(ybar[191]);
  AND2_X1 U156 ( .A1(a[11]), .A2(b[14]), .ZN(y[190]) );
  OR2_X1 U156bar ( .A1(abar[11]), .A2(bbar[14]), .ZN(ybar[190]);
  AND2_X1 U157 ( .A1(a[1]), .A2(b[2]), .ZN(y[18]) );
  OR2_X1 U157bar ( .A1(abar[1]), .A2(bbar[2]), .ZN(ybar[18]);
  AND2_X1 U158 ( .A1(a[11]), .A2(b[13]), .ZN(y[189]) );
  OR2_X1 U158bar ( .A1(abar[11]), .A2(bbar[13]), .ZN(ybar[189]);
  AND2_X1 U159 ( .A1(a[11]), .A2(b[12]), .ZN(y[188]) );
  OR2_X1 U159bar ( .A1(abar[11]), .A2(bbar[12]), .ZN(ybar[188]);
  AND2_X1 U160 ( .A1(a[11]), .A2(b[11]), .ZN(y[187]) );
  OR2_X1 U160bar ( .A1(abar[11]), .A2(bbar[11]), .ZN(ybar[187]);
  AND2_X1 U161 ( .A1(a[11]), .A2(b[10]), .ZN(y[186]) );
  OR2_X1 U161bar ( .A1(abar[11]), .A2(bbar[10]), .ZN(ybar[186]);
  AND2_X1 U162 ( .A1(a[11]), .A2(b[9]), .ZN(y[185]) );
  OR2_X1 U162bar ( .A1(abar[11]), .A2(bbar[9]), .ZN(ybar[185]);
  AND2_X1 U163 ( .A1(a[11]), .A2(b[8]), .ZN(y[184]) );
  OR2_X1 U163bar ( .A1(abar[11]), .A2(bbar[8]), .ZN(ybar[184]);
  AND2_X1 U164 ( .A1(a[11]), .A2(b[7]), .ZN(y[183]) );
  OR2_X1 U164bar ( .A1(abar[11]), .A2(bbar[7]), .ZN(ybar[183]);
  AND2_X1 U165 ( .A1(a[11]), .A2(b[6]), .ZN(y[182]) );
  OR2_X1 U165bar ( .A1(abar[11]), .A2(bbar[6]), .ZN(ybar[182]);
  AND2_X1 U166 ( .A1(a[11]), .A2(b[5]), .ZN(y[181]) );
  OR2_X1 U166bar ( .A1(abar[11]), .A2(bbar[5]), .ZN(ybar[181]);
  AND2_X1 U167 ( .A1(a[11]), .A2(b[4]), .ZN(y[180]) );
  OR2_X1 U167bar ( .A1(abar[11]), .A2(bbar[4]), .ZN(ybar[180]);
  AND2_X1 U168 ( .A1(a[1]), .A2(b[1]), .ZN(y[17]) );
  OR2_X1 U168bar ( .A1(abar[1]), .A2(bbar[1]), .ZN(ybar[17]);
  AND2_X1 U169 ( .A1(a[11]), .A2(b[3]), .ZN(y[179]) );
  OR2_X1 U169bar ( .A1(abar[11]), .A2(bbar[3]), .ZN(ybar[179]);
  AND2_X1 U170 ( .A1(a[11]), .A2(b[2]), .ZN(y[178]) );
  OR2_X1 U170bar ( .A1(abar[11]), .A2(bbar[2]), .ZN(ybar[178]);
  AND2_X1 U171 ( .A1(a[11]), .A2(b[1]), .ZN(y[177]) );
  OR2_X1 U171bar ( .A1(abar[11]), .A2(bbar[1]), .ZN(ybar[177]);
  AND2_X1 U172 ( .A1(a[11]), .A2(b[0]), .ZN(y[176]) );
  OR2_X1 U172bar ( .A1(abar[11]), .A2(bbar[0]), .ZN(ybar[176]);
  AND2_X1 U173 ( .A1(a[10]), .A2(b[15]), .ZN(y[175]) );
  OR2_X1 U173bar ( .A1(abar[10]), .A2(bbar[15]), .ZN(ybar[175]);
  AND2_X1 U174 ( .A1(a[10]), .A2(b[14]), .ZN(y[174]) );
  OR2_X1 U174bar ( .A1(abar[10]), .A2(bbar[14]), .ZN(ybar[174]);
  AND2_X1 U175 ( .A1(a[10]), .A2(b[13]), .ZN(y[173]) );
  OR2_X1 U175bar ( .A1(abar[10]), .A2(bbar[13]), .ZN(ybar[173]);
  AND2_X1 U176 ( .A1(a[10]), .A2(b[12]), .ZN(y[172]) );
  OR2_X1 U176bar ( .A1(abar[10]), .A2(bbar[12]), .ZN(ybar[172]);
  AND2_X1 U177 ( .A1(a[10]), .A2(b[11]), .ZN(y[171]) );
  OR2_X1 U177bar ( .A1(abar[10]), .A2(bbar[11]), .ZN(ybar[171]);
  AND2_X1 U178 ( .A1(a[10]), .A2(b[10]), .ZN(y[170]) );
  OR2_X1 U178bar ( .A1(abar[10]), .A2(bbar[10]), .ZN(ybar[170]);
  AND2_X1 U179 ( .A1(a[1]), .A2(b[0]), .ZN(y[16]) );
  OR2_X1 U179bar ( .A1(abar[1]), .A2(bbar[0]), .ZN(ybar[16]);
  AND2_X1 U180 ( .A1(a[10]), .A2(b[9]), .ZN(y[169]) );
  OR2_X1 U180bar ( .A1(abar[10]), .A2(bbar[9]), .ZN(ybar[169]);
  AND2_X1 U181 ( .A1(a[10]), .A2(b[8]), .ZN(y[168]) );
  OR2_X1 U181bar ( .A1(abar[10]), .A2(bbar[8]), .ZN(ybar[168]);
  AND2_X1 U182 ( .A1(a[10]), .A2(b[7]), .ZN(y[167]) );
  OR2_X1 U182bar ( .A1(abar[10]), .A2(bbar[7]), .ZN(ybar[167]);
  AND2_X1 U183 ( .A1(a[10]), .A2(b[6]), .ZN(y[166]) );
  OR2_X1 U183bar ( .A1(abar[10]), .A2(bbar[6]), .ZN(ybar[166]);
  AND2_X1 U184 ( .A1(a[10]), .A2(b[5]), .ZN(y[165]) );
  OR2_X1 U184bar ( .A1(abar[10]), .A2(bbar[5]), .ZN(ybar[165]);
  AND2_X1 U185 ( .A1(a[10]), .A2(b[4]), .ZN(y[164]) );
  OR2_X1 U185bar ( .A1(abar[10]), .A2(bbar[4]), .ZN(ybar[164]);
  AND2_X1 U186 ( .A1(a[10]), .A2(b[3]), .ZN(y[163]) );
  OR2_X1 U186bar ( .A1(abar[10]), .A2(bbar[3]), .ZN(ybar[163]);
  AND2_X1 U187 ( .A1(a[10]), .A2(b[2]), .ZN(y[162]) );
  OR2_X1 U187bar ( .A1(abar[10]), .A2(bbar[2]), .ZN(ybar[162]);
  AND2_X1 U188 ( .A1(a[10]), .A2(b[1]), .ZN(y[161]) );
  OR2_X1 U188bar ( .A1(abar[10]), .A2(bbar[1]), .ZN(ybar[161]);
  AND2_X1 U189 ( .A1(a[10]), .A2(b[0]), .ZN(y[160]) );
  OR2_X1 U189bar ( .A1(abar[10]), .A2(bbar[0]), .ZN(ybar[160]);
  AND2_X1 U190 ( .A1(b[15]), .A2(a[0]), .ZN(y[15]) );
  OR2_X1 U190bar ( .A1(bbar[15]), .A2(abar[0]), .ZN(ybar[15]);
  AND2_X1 U191 ( .A1(a[9]), .A2(b[15]), .ZN(y[159]) );
  OR2_X1 U191bar ( .A1(abar[9]), .A2(bbar[15]), .ZN(ybar[159]);
  AND2_X1 U192 ( .A1(a[9]), .A2(b[14]), .ZN(y[158]) );
  OR2_X1 U192bar ( .A1(abar[9]), .A2(bbar[14]), .ZN(ybar[158]);
  AND2_X1 U193 ( .A1(a[9]), .A2(b[13]), .ZN(y[157]) );
  OR2_X1 U193bar ( .A1(abar[9]), .A2(bbar[13]), .ZN(ybar[157]);
  AND2_X1 U194 ( .A1(a[9]), .A2(b[12]), .ZN(y[156]) );
  OR2_X1 U194bar ( .A1(abar[9]), .A2(bbar[12]), .ZN(ybar[156]);
  AND2_X1 U195 ( .A1(a[9]), .A2(b[11]), .ZN(y[155]) );
  OR2_X1 U195bar ( .A1(abar[9]), .A2(bbar[11]), .ZN(ybar[155]);
  AND2_X1 U196 ( .A1(a[9]), .A2(b[10]), .ZN(y[154]) );
  OR2_X1 U196bar ( .A1(abar[9]), .A2(bbar[10]), .ZN(ybar[154]);
  AND2_X1 U197 ( .A1(a[9]), .A2(b[9]), .ZN(y[153]) );
  OR2_X1 U197bar ( .A1(abar[9]), .A2(bbar[9]), .ZN(ybar[153]);
  AND2_X1 U198 ( .A1(a[9]), .A2(b[8]), .ZN(y[152]) );
  OR2_X1 U198bar ( .A1(abar[9]), .A2(bbar[8]), .ZN(ybar[152]);
  AND2_X1 U199 ( .A1(a[9]), .A2(b[7]), .ZN(y[151]) );
  OR2_X1 U199bar ( .A1(abar[9]), .A2(bbar[7]), .ZN(ybar[151]);
  AND2_X1 U200 ( .A1(a[9]), .A2(b[6]), .ZN(y[150]) );
  OR2_X1 U200bar ( .A1(abar[9]), .A2(bbar[6]), .ZN(ybar[150]);
  AND2_X1 U201 ( .A1(b[14]), .A2(a[0]), .ZN(y[14]) );
  OR2_X1 U201bar ( .A1(bbar[14]), .A2(abar[0]), .ZN(ybar[14]);
  AND2_X1 U202 ( .A1(a[9]), .A2(b[5]), .ZN(y[149]) );
  OR2_X1 U202bar ( .A1(abar[9]), .A2(bbar[5]), .ZN(ybar[149]);
  AND2_X1 U203 ( .A1(a[9]), .A2(b[4]), .ZN(y[148]) );
  OR2_X1 U203bar ( .A1(abar[9]), .A2(bbar[4]), .ZN(ybar[148]);
  AND2_X1 U204 ( .A1(a[9]), .A2(b[3]), .ZN(y[147]) );
  OR2_X1 U204bar ( .A1(abar[9]), .A2(bbar[3]), .ZN(ybar[147]);
  AND2_X1 U205 ( .A1(a[9]), .A2(b[2]), .ZN(y[146]) );
  OR2_X1 U205bar ( .A1(abar[9]), .A2(bbar[2]), .ZN(ybar[146]);
  AND2_X1 U206 ( .A1(a[9]), .A2(b[1]), .ZN(y[145]) );
  OR2_X1 U206bar ( .A1(abar[9]), .A2(bbar[1]), .ZN(ybar[145]);
  AND2_X1 U207 ( .A1(a[9]), .A2(b[0]), .ZN(y[144]) );
  OR2_X1 U207bar ( .A1(abar[9]), .A2(bbar[0]), .ZN(ybar[144]);
  AND2_X1 U208 ( .A1(a[8]), .A2(b[15]), .ZN(y[143]) );
  OR2_X1 U208bar ( .A1(abar[8]), .A2(bbar[15]), .ZN(ybar[143]);
  AND2_X1 U209 ( .A1(a[8]), .A2(b[14]), .ZN(y[142]) );
  OR2_X1 U209bar ( .A1(abar[8]), .A2(bbar[14]), .ZN(ybar[142]);
  AND2_X1 U210 ( .A1(a[8]), .A2(b[13]), .ZN(y[141]) );
  OR2_X1 U210bar ( .A1(abar[8]), .A2(bbar[13]), .ZN(ybar[141]);
  AND2_X1 U211 ( .A1(a[8]), .A2(b[12]), .ZN(y[140]) );
  OR2_X1 U211bar ( .A1(abar[8]), .A2(bbar[12]), .ZN(ybar[140]);
  AND2_X1 U212 ( .A1(b[13]), .A2(a[0]), .ZN(y[13]) );
  OR2_X1 U212bar ( .A1(bbar[13]), .A2(abar[0]), .ZN(ybar[13]);
  AND2_X1 U213 ( .A1(a[8]), .A2(b[11]), .ZN(y[139]) );
  OR2_X1 U213bar ( .A1(abar[8]), .A2(bbar[11]), .ZN(ybar[139]);
  AND2_X1 U214 ( .A1(a[8]), .A2(b[10]), .ZN(y[138]) );
  OR2_X1 U214bar ( .A1(abar[8]), .A2(bbar[10]), .ZN(ybar[138]);
  AND2_X1 U215 ( .A1(a[8]), .A2(b[9]), .ZN(y[137]) );
  OR2_X1 U215bar ( .A1(abar[8]), .A2(bbar[9]), .ZN(ybar[137]);
  AND2_X1 U216 ( .A1(a[8]), .A2(b[8]), .ZN(y[136]) );
  OR2_X1 U216bar ( .A1(abar[8]), .A2(bbar[8]), .ZN(ybar[136]);
  AND2_X1 U217 ( .A1(a[8]), .A2(b[7]), .ZN(y[135]) );
  OR2_X1 U217bar ( .A1(abar[8]), .A2(bbar[7]), .ZN(ybar[135]);
  AND2_X1 U218 ( .A1(a[8]), .A2(b[6]), .ZN(y[134]) );
  OR2_X1 U218bar ( .A1(abar[8]), .A2(bbar[6]), .ZN(ybar[134]);
  AND2_X1 U219 ( .A1(a[8]), .A2(b[5]), .ZN(y[133]) );
  OR2_X1 U219bar ( .A1(abar[8]), .A2(bbar[5]), .ZN(ybar[133]);
  AND2_X1 U220 ( .A1(a[8]), .A2(b[4]), .ZN(y[132]) );
  OR2_X1 U220bar ( .A1(abar[8]), .A2(bbar[4]), .ZN(ybar[132]);
  AND2_X1 U221 ( .A1(a[8]), .A2(b[3]), .ZN(y[131]) );
  OR2_X1 U221bar ( .A1(abar[8]), .A2(bbar[3]), .ZN(ybar[131]);
  AND2_X1 U222 ( .A1(a[8]), .A2(b[2]), .ZN(y[130]) );
  OR2_X1 U222bar ( .A1(abar[8]), .A2(bbar[2]), .ZN(ybar[130]);
  AND2_X1 U223 ( .A1(b[12]), .A2(a[0]), .ZN(y[12]) );
  OR2_X1 U223bar ( .A1(bbar[12]), .A2(abar[0]), .ZN(ybar[12]);
  AND2_X1 U224 ( .A1(a[8]), .A2(b[1]), .ZN(y[129]) );
  OR2_X1 U224bar ( .A1(abar[8]), .A2(bbar[1]), .ZN(ybar[129]);
  AND2_X1 U225 ( .A1(a[8]), .A2(b[0]), .ZN(y[128]) );
  OR2_X1 U225bar ( .A1(abar[8]), .A2(bbar[0]), .ZN(ybar[128]);
  AND2_X1 U226 ( .A1(a[7]), .A2(b[15]), .ZN(y[127]) );
  OR2_X1 U226bar ( .A1(abar[7]), .A2(bbar[15]), .ZN(ybar[127]);
  AND2_X1 U227 ( .A1(a[7]), .A2(b[14]), .ZN(y[126]) );
  OR2_X1 U227bar ( .A1(abar[7]), .A2(bbar[14]), .ZN(ybar[126]);
  AND2_X1 U228 ( .A1(a[7]), .A2(b[13]), .ZN(y[125]) );
  OR2_X1 U228bar ( .A1(abar[7]), .A2(bbar[13]), .ZN(ybar[125]);
  AND2_X1 U229 ( .A1(a[7]), .A2(b[12]), .ZN(y[124]) );
  OR2_X1 U229bar ( .A1(abar[7]), .A2(bbar[12]), .ZN(ybar[124]);
  AND2_X1 U230 ( .A1(a[7]), .A2(b[11]), .ZN(y[123]) );
  OR2_X1 U230bar ( .A1(abar[7]), .A2(bbar[11]), .ZN(ybar[123]);
  AND2_X1 U231 ( .A1(a[7]), .A2(b[10]), .ZN(y[122]) );
  OR2_X1 U231bar ( .A1(abar[7]), .A2(bbar[10]), .ZN(ybar[122]);
  AND2_X1 U232 ( .A1(a[7]), .A2(b[9]), .ZN(y[121]) );
  OR2_X1 U232bar ( .A1(abar[7]), .A2(bbar[9]), .ZN(ybar[121]);
  AND2_X1 U233 ( .A1(a[7]), .A2(b[8]), .ZN(y[120]) );
  OR2_X1 U233bar ( .A1(abar[7]), .A2(bbar[8]), .ZN(ybar[120]);
  AND2_X1 U234 ( .A1(b[11]), .A2(a[0]), .ZN(y[11]) );
  OR2_X1 U234bar ( .A1(bbar[11]), .A2(abar[0]), .ZN(ybar[11]);
  AND2_X1 U235 ( .A1(a[7]), .A2(b[7]), .ZN(y[119]) );
  OR2_X1 U235bar ( .A1(abar[7]), .A2(bbar[7]), .ZN(ybar[119]);
  AND2_X1 U236 ( .A1(a[7]), .A2(b[6]), .ZN(y[118]) );
  OR2_X1 U236bar ( .A1(abar[7]), .A2(bbar[6]), .ZN(ybar[118]);
  AND2_X1 U237 ( .A1(a[7]), .A2(b[5]), .ZN(y[117]) );
  OR2_X1 U237bar ( .A1(abar[7]), .A2(bbar[5]), .ZN(ybar[117]);
  AND2_X1 U238 ( .A1(a[7]), .A2(b[4]), .ZN(y[116]) );
  OR2_X1 U238bar ( .A1(abar[7]), .A2(bbar[4]), .ZN(ybar[116]);
  AND2_X1 U239 ( .A1(a[7]), .A2(b[3]), .ZN(y[115]) );
  OR2_X1 U239bar ( .A1(abar[7]), .A2(bbar[3]), .ZN(ybar[115]);
  AND2_X1 U240 ( .A1(a[7]), .A2(b[2]), .ZN(y[114]) );
  OR2_X1 U240bar ( .A1(abar[7]), .A2(bbar[2]), .ZN(ybar[114]);
  AND2_X1 U241 ( .A1(a[7]), .A2(b[1]), .ZN(y[113]) );
  OR2_X1 U241bar ( .A1(abar[7]), .A2(bbar[1]), .ZN(ybar[113]);
  AND2_X1 U242 ( .A1(a[7]), .A2(b[0]), .ZN(y[112]) );
  OR2_X1 U242bar ( .A1(abar[7]), .A2(bbar[0]), .ZN(ybar[112]);
  AND2_X1 U243 ( .A1(b[15]), .A2(a[6]), .ZN(y[111]) );
  OR2_X1 U243bar ( .A1(bbar[15]), .A2(abar[6]), .ZN(ybar[111]);
  AND2_X1 U244 ( .A1(b[14]), .A2(a[6]), .ZN(y[110]) );
  OR2_X1 U244bar ( .A1(bbar[14]), .A2(abar[6]), .ZN(ybar[110]);
  AND2_X1 U245 ( .A1(b[10]), .A2(a[0]), .ZN(y[10]) );
  OR2_X1 U245bar ( .A1(bbar[10]), .A2(abar[0]), .ZN(ybar[10]);
  AND2_X1 U246 ( .A1(b[13]), .A2(a[6]), .ZN(y[109]) );
  OR2_X1 U246bar ( .A1(bbar[13]), .A2(abar[6]), .ZN(ybar[109]);
  AND2_X1 U247 ( .A1(b[12]), .A2(a[6]), .ZN(y[108]) );
  OR2_X1 U247bar ( .A1(bbar[12]), .A2(abar[6]), .ZN(ybar[108]);
  AND2_X1 U248 ( .A1(b[11]), .A2(a[6]), .ZN(y[107]) );
  OR2_X1 U248bar ( .A1(bbar[11]), .A2(abar[6]), .ZN(ybar[107]);
  AND2_X1 U249 ( .A1(b[10]), .A2(a[6]), .ZN(y[106]) );
  OR2_X1 U249bar ( .A1(bbar[10]), .A2(abar[6]), .ZN(ybar[106]);
  AND2_X1 U250 ( .A1(a[6]), .A2(b[9]), .ZN(y[105]) );
  OR2_X1 U250bar ( .A1(abar[6]), .A2(bbar[9]), .ZN(ybar[105]);
  AND2_X1 U251 ( .A1(b[8]), .A2(a[6]), .ZN(y[104]) );
  OR2_X1 U251bar ( .A1(bbar[8]), .A2(abar[6]), .ZN(ybar[104]);
  AND2_X1 U252 ( .A1(b[7]), .A2(a[6]), .ZN(y[103]) );
  OR2_X1 U252bar ( .A1(bbar[7]), .A2(abar[6]), .ZN(ybar[103]);
  AND2_X1 U253 ( .A1(b[6]), .A2(a[6]), .ZN(y[102]) );
  OR2_X1 U253bar ( .A1(bbar[6]), .A2(abar[6]), .ZN(ybar[102]);
  AND2_X1 U254 ( .A1(b[5]), .A2(a[6]), .ZN(y[101]) );
  OR2_X1 U254bar ( .A1(bbar[5]), .A2(abar[6]), .ZN(ybar[101]);
  AND2_X1 U255 ( .A1(b[4]), .A2(a[6]), .ZN(y[100]) );
  OR2_X1 U255bar ( .A1(bbar[4]), .A2(abar[6]), .ZN(ybar[100]);
  AND2_X1 U256 ( .A1(b[0]), .A2(a[0]), .ZN(y[0]) );
  OR2_X1 U256bar ( .A1(bbar[0]), .A2(abar[0]), .ZN(ybar[0]);
endmodule




module decode_19 ( in, out );
  input [7:0] in;
  //input_done

  output [255:0] out;
  //output_done

  wire   [15:0] level1;
  wire   [31:0] level2;
  //wire_done

  CD2_76 cd_l1_1 ( .a(in[1]), .b(in[0]), .y(level1[3:0]) );
  CD2_75 cd_l1_2 ( .a(in[3]), .b(in[2]), .y(level1[7:4]) );
  CD2_74 cd_l1_3 ( .a(in[5]), .b(in[4]), .y(level1[11:8]) );
  CD2_73 cd_l1_4 ( .a(in[7]), .b(in[6]), .y(level1[15:12]) );
  CD4_38 cd_l2_1 ( .a(level1[7:4]), .b(level1[3:0]), .y(level2[15:0]) );
  CD4_37 cd_l2_2 ( .a(level1[15:12]), .b(level1[11:8]), .y(level2[31:16]) );
  CD16_19 cd_l3 ( .a(level2[31:16]), .b(level2[15:0]), .y(out) );
endmodule


module encode_19 ( in, out );
  input [255:0] in;
  assign inbar[0] = ~in[0];
  assign inbar[1] = ~in[1];
  assign inbar[2] = ~in[2];
  assign inbar[3] = ~in[3];
  assign inbar[4] = ~in[4];
  assign inbar[5] = ~in[5];
  assign inbar[6] = ~in[6];
  assign inbar[7] = ~in[7];
  assign inbar[8] = ~in[8];
  assign inbar[9] = ~in[9];
  assign inbar[10] = ~in[10];
  assign inbar[11] = ~in[11];
  assign inbar[12] = ~in[12];
  assign inbar[13] = ~in[13];
  assign inbar[14] = ~in[14];
  assign inbar[15] = ~in[15];
  assign inbar[16] = ~in[16];
  assign inbar[17] = ~in[17];
  assign inbar[18] = ~in[18];
  assign inbar[19] = ~in[19];
  assign inbar[20] = ~in[20];
  assign inbar[21] = ~in[21];
  assign inbar[22] = ~in[22];
  assign inbar[23] = ~in[23];
  assign inbar[24] = ~in[24];
  assign inbar[25] = ~in[25];
  assign inbar[26] = ~in[26];
  assign inbar[27] = ~in[27];
  assign inbar[28] = ~in[28];
  assign inbar[29] = ~in[29];
  assign inbar[30] = ~in[30];
  assign inbar[31] = ~in[31];
  assign inbar[32] = ~in[32];
  assign inbar[33] = ~in[33];
  assign inbar[34] = ~in[34];
  assign inbar[35] = ~in[35];
  assign inbar[36] = ~in[36];
  assign inbar[37] = ~in[37];
  assign inbar[38] = ~in[38];
  assign inbar[39] = ~in[39];
  assign inbar[40] = ~in[40];
  assign inbar[41] = ~in[41];
  assign inbar[42] = ~in[42];
  assign inbar[43] = ~in[43];
  assign inbar[44] = ~in[44];
  assign inbar[45] = ~in[45];
  assign inbar[46] = ~in[46];
  assign inbar[47] = ~in[47];
  assign inbar[48] = ~in[48];
  assign inbar[49] = ~in[49];
  assign inbar[50] = ~in[50];
  assign inbar[51] = ~in[51];
  assign inbar[52] = ~in[52];
  assign inbar[53] = ~in[53];
  assign inbar[54] = ~in[54];
  assign inbar[55] = ~in[55];
  assign inbar[56] = ~in[56];
  assign inbar[57] = ~in[57];
  assign inbar[58] = ~in[58];
  assign inbar[59] = ~in[59];
  assign inbar[60] = ~in[60];
  assign inbar[61] = ~in[61];
  assign inbar[62] = ~in[62];
  assign inbar[63] = ~in[63];
  assign inbar[64] = ~in[64];
  assign inbar[65] = ~in[65];
  assign inbar[66] = ~in[66];
  assign inbar[67] = ~in[67];
  assign inbar[68] = ~in[68];
  assign inbar[69] = ~in[69];
  assign inbar[70] = ~in[70];
  assign inbar[71] = ~in[71];
  assign inbar[72] = ~in[72];
  assign inbar[73] = ~in[73];
  assign inbar[74] = ~in[74];
  assign inbar[75] = ~in[75];
  assign inbar[76] = ~in[76];
  assign inbar[77] = ~in[77];
  assign inbar[78] = ~in[78];
  assign inbar[79] = ~in[79];
  assign inbar[80] = ~in[80];
  assign inbar[81] = ~in[81];
  assign inbar[82] = ~in[82];
  assign inbar[83] = ~in[83];
  assign inbar[84] = ~in[84];
  assign inbar[85] = ~in[85];
  assign inbar[86] = ~in[86];
  assign inbar[87] = ~in[87];
  assign inbar[88] = ~in[88];
  assign inbar[89] = ~in[89];
  assign inbar[90] = ~in[90];
  assign inbar[91] = ~in[91];
  assign inbar[92] = ~in[92];
  assign inbar[93] = ~in[93];
  assign inbar[94] = ~in[94];
  assign inbar[95] = ~in[95];
  assign inbar[96] = ~in[96];
  assign inbar[97] = ~in[97];
  assign inbar[98] = ~in[98];
  assign inbar[99] = ~in[99];
  assign inbar[100] = ~in[100];
  assign inbar[101] = ~in[101];
  assign inbar[102] = ~in[102];
  assign inbar[103] = ~in[103];
  assign inbar[104] = ~in[104];
  assign inbar[105] = ~in[105];
  assign inbar[106] = ~in[106];
  assign inbar[107] = ~in[107];
  assign inbar[108] = ~in[108];
  assign inbar[109] = ~in[109];
  assign inbar[110] = ~in[110];
  assign inbar[111] = ~in[111];
  assign inbar[112] = ~in[112];
  assign inbar[113] = ~in[113];
  assign inbar[114] = ~in[114];
  assign inbar[115] = ~in[115];
  assign inbar[116] = ~in[116];
  assign inbar[117] = ~in[117];
  assign inbar[118] = ~in[118];
  assign inbar[119] = ~in[119];
  assign inbar[120] = ~in[120];
  assign inbar[121] = ~in[121];
  assign inbar[122] = ~in[122];
  assign inbar[123] = ~in[123];
  assign inbar[124] = ~in[124];
  assign inbar[125] = ~in[125];
  assign inbar[126] = ~in[126];
  assign inbar[127] = ~in[127];
  assign inbar[128] = ~in[128];
  assign inbar[129] = ~in[129];
  assign inbar[130] = ~in[130];
  assign inbar[131] = ~in[131];
  assign inbar[132] = ~in[132];
  assign inbar[133] = ~in[133];
  assign inbar[134] = ~in[134];
  assign inbar[135] = ~in[135];
  assign inbar[136] = ~in[136];
  assign inbar[137] = ~in[137];
  assign inbar[138] = ~in[138];
  assign inbar[139] = ~in[139];
  assign inbar[140] = ~in[140];
  assign inbar[141] = ~in[141];
  assign inbar[142] = ~in[142];
  assign inbar[143] = ~in[143];
  assign inbar[144] = ~in[144];
  assign inbar[145] = ~in[145];
  assign inbar[146] = ~in[146];
  assign inbar[147] = ~in[147];
  assign inbar[148] = ~in[148];
  assign inbar[149] = ~in[149];
  assign inbar[150] = ~in[150];
  assign inbar[151] = ~in[151];
  assign inbar[152] = ~in[152];
  assign inbar[153] = ~in[153];
  assign inbar[154] = ~in[154];
  assign inbar[155] = ~in[155];
  assign inbar[156] = ~in[156];
  assign inbar[157] = ~in[157];
  assign inbar[158] = ~in[158];
  assign inbar[159] = ~in[159];
  assign inbar[160] = ~in[160];
  assign inbar[161] = ~in[161];
  assign inbar[162] = ~in[162];
  assign inbar[163] = ~in[163];
  assign inbar[164] = ~in[164];
  assign inbar[165] = ~in[165];
  assign inbar[166] = ~in[166];
  assign inbar[167] = ~in[167];
  assign inbar[168] = ~in[168];
  assign inbar[169] = ~in[169];
  assign inbar[170] = ~in[170];
  assign inbar[171] = ~in[171];
  assign inbar[172] = ~in[172];
  assign inbar[173] = ~in[173];
  assign inbar[174] = ~in[174];
  assign inbar[175] = ~in[175];
  assign inbar[176] = ~in[176];
  assign inbar[177] = ~in[177];
  assign inbar[178] = ~in[178];
  assign inbar[179] = ~in[179];
  assign inbar[180] = ~in[180];
  assign inbar[181] = ~in[181];
  assign inbar[182] = ~in[182];
  assign inbar[183] = ~in[183];
  assign inbar[184] = ~in[184];
  assign inbar[185] = ~in[185];
  assign inbar[186] = ~in[186];
  assign inbar[187] = ~in[187];
  assign inbar[188] = ~in[188];
  assign inbar[189] = ~in[189];
  assign inbar[190] = ~in[190];
  assign inbar[191] = ~in[191];
  assign inbar[192] = ~in[192];
  assign inbar[193] = ~in[193];
  assign inbar[194] = ~in[194];
  assign inbar[195] = ~in[195];
  assign inbar[196] = ~in[196];
  assign inbar[197] = ~in[197];
  assign inbar[198] = ~in[198];
  assign inbar[199] = ~in[199];
  assign inbar[200] = ~in[200];
  assign inbar[201] = ~in[201];
  assign inbar[202] = ~in[202];
  assign inbar[203] = ~in[203];
  assign inbar[204] = ~in[204];
  assign inbar[205] = ~in[205];
  assign inbar[206] = ~in[206];
  assign inbar[207] = ~in[207];
  assign inbar[208] = ~in[208];
  assign inbar[209] = ~in[209];
  assign inbar[210] = ~in[210];
  assign inbar[211] = ~in[211];
  assign inbar[212] = ~in[212];
  assign inbar[213] = ~in[213];
  assign inbar[214] = ~in[214];
  assign inbar[215] = ~in[215];
  assign inbar[216] = ~in[216];
  assign inbar[217] = ~in[217];
  assign inbar[218] = ~in[218];
  assign inbar[219] = ~in[219];
  assign inbar[220] = ~in[220];
  assign inbar[221] = ~in[221];
  assign inbar[222] = ~in[222];
  assign inbar[223] = ~in[223];
  assign inbar[224] = ~in[224];
  assign inbar[225] = ~in[225];
  assign inbar[226] = ~in[226];
  assign inbar[227] = ~in[227];
  assign inbar[228] = ~in[228];
  assign inbar[229] = ~in[229];
  assign inbar[230] = ~in[230];
  assign inbar[231] = ~in[231];
  assign inbar[232] = ~in[232];
  assign inbar[233] = ~in[233];
  assign inbar[234] = ~in[234];
  assign inbar[235] = ~in[235];
  assign inbar[236] = ~in[236];
  assign inbar[237] = ~in[237];
  assign inbar[238] = ~in[238];
  assign inbar[239] = ~in[239];
  assign inbar[240] = ~in[240];
  assign inbar[241] = ~in[241];
  assign inbar[242] = ~in[242];
  assign inbar[243] = ~in[243];
  assign inbar[244] = ~in[244];
  assign inbar[245] = ~in[245];
  assign inbar[246] = ~in[246];
  assign inbar[247] = ~in[247];
  assign inbar[248] = ~in[248];
  assign inbar[249] = ~in[249];
  assign inbar[250] = ~in[250];
  assign inbar[251] = ~in[251];
  assign inbar[252] = ~in[252];
  assign inbar[253] = ~in[253];
  assign inbar[254] = ~in[254];
  assign inbar[255] = ~in[255];
  //input_done

  output [7:0] out;
  reg [7:0] outbar;
  //output_done

  wire   in_81, in_80, in_79, in_78, in_77, in_76, in_75, in_74, in_73, in_72,
         in_71, in_70, in_69, in_68, in_67, in_66, in_65, in_64, in_63, in_62,
         in_61, in_60, in_59, in_58, in_57, in_56, in_55, in_54, in_53, in_52,
         in_51, in_50, in_49, in_48, in_47, in_46, in_45, in_44, in_43, in_42,
         in_41, in_40, in_39, in_38, in_37, in_36, in_35, in_34, in_33, in_32,
         in_31, in_30, in_29, in_28, in_27, in_26, in_25, in_24, in_23, in_22,
         in_21, in_20, in_19, in_18, in_17, in_16, in_15, in_14, in_13, in_12,
         in_11, in_10, in_9, in_8, in_7, in_6, in_5, in_4, in_3, in_2, in_1,
         in_0, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972;
  wire in_81bar, in_80bar, in_79bar, in_78bar, in_77bar, in_76bar, in_75bar, in_74bar, in_73bar, in_72bar, in_71bar, in_70bar, in_69bar, in_68bar, in_67bar, in_66bar, in_65bar, in_64bar, in_63bar, in_62bar, in_61bar, in_60bar, in_59bar, in_58bar, in_57bar, in_56bar, in_55bar, in_54bar, in_53bar, in_52bar, in_51bar, in_50bar, in_49bar, in_48bar, in_47bar, in_46bar, in_45bar, in_44bar, in_43bar, in_42bar, in_41bar, in_40bar, in_39bar, in_38bar, in_37bar, in_36bar, in_35bar, in_34bar, in_33bar, in_32bar, in_31bar, in_30bar, in_29bar, in_28bar, in_27bar, in_26bar, in_25bar, in_24bar, in_23bar, in_22bar, in_21bar, in_20bar, in_19bar, in_18bar, in_17bar, in_16bar, in_15bar, in_14bar, in_13bar, in_12bar, in_11bar, in_10bar, in_9bar, in_8bar, in_7bar, in_6bar, in_5bar, in_4bar, in_3bar, in_2bar, in_1bar, in_0bar, n487bar, n488bar, n489bar, n490bar, n491bar, n492bar, n493bar, n494bar, n495bar, n496bar, n497bar, n498bar, n499bar, n500bar, n501bar, n502bar, n503bar, n504bar, n505bar, n506bar, n507bar, n508bar, n509bar, n510bar, n511bar, n512bar, n513bar, n514bar, n515bar, n516bar, n517bar, n518bar, n519bar, n520bar, n521bar, n522bar, n523bar, n524bar, n525bar, n526bar, n527bar, n528bar, n529bar, n530bar, n531bar, n532bar, n533bar, n534bar, n535bar, n536bar, n537bar, n538bar, n539bar, n540bar, n541bar, n542bar, n543bar, n544bar, n545bar, n546bar, n547bar, n548bar, n549bar, n550bar, n551bar, n552bar, n553bar, n554bar, n555bar, n556bar, n557bar, n558bar, n559bar, n560bar, n561bar, n562bar, n563bar, n564bar, n565bar, n566bar, n567bar, n568bar, n569bar, n570bar, n571bar, n572bar, n573bar, n574bar, n575bar, n576bar, n577bar, n578bar, n579bar, n580bar, n581bar, n582bar, n583bar, n584bar, n585bar, n586bar, n587bar, n588bar, n589bar, n590bar, n591bar, n592bar, n593bar, n594bar, n595bar, n596bar, n597bar, n598bar, n599bar, n600bar, n601bar, n602bar, n603bar, n604bar, n605bar, n606bar, n607bar, n608bar, n609bar, n610bar, n611bar, n612bar, n613bar, n614bar, n615bar, n616bar, n617bar, n618bar, n619bar, n620bar, n621bar, n622bar, n623bar, n624bar, n625bar, n626bar, n627bar, n628bar, n629bar, n630bar, n631bar, n632bar, n633bar, n634bar, n635bar, n636bar, n637bar, n638bar, n639bar, n640bar, n641bar, n642bar, n643bar, n644bar, n645bar, n646bar, n647bar, n648bar, n649bar, n650bar, n651bar, n652bar, n653bar, n654bar, n655bar, n656bar, n657bar, n658bar, n659bar, n660bar, n661bar, n662bar, n663bar, n664bar, n665bar, n666bar, n667bar, n668bar, n669bar, n670bar, n671bar, n672bar, n673bar, n674bar, n675bar, n676bar, n677bar, n678bar, n679bar, n680bar, n681bar, n682bar, n683bar, n684bar, n685bar, n686bar, n687bar, n688bar, n689bar, n690bar, n691bar, n692bar, n693bar, n694bar, n695bar, n696bar, n697bar, n698bar, n699bar, n700bar, n701bar, n702bar, n703bar, n704bar, n705bar, n706bar, n707bar, n708bar, n709bar, n710bar, n711bar, n712bar, n713bar, n714bar, n715bar, n716bar, n717bar, n718bar, n719bar, n720bar, n721bar, n722bar, n723bar, n724bar, n725bar, n726bar, n727bar, n728bar, n729bar, n730bar, n731bar, n732bar, n733bar, n734bar, n735bar, n736bar, n737bar, n738bar, n739bar, n740bar, n741bar, n742bar, n743bar, n744bar, n745bar, n746bar, n747bar, n748bar, n749bar, n750bar, n751bar, n752bar, n753bar, n754bar, n755bar, n756bar, n757bar, n758bar, n759bar, n760bar, n761bar, n762bar, n763bar, n764bar, n765bar, n766bar, n767bar, n768bar, n769bar, n770bar, n771bar, n772bar, n773bar, n774bar, n775bar, n776bar, n777bar, n778bar, n779bar, n780bar, n781bar, n782bar, n783bar, n784bar, n785bar, n786bar, n787bar, n788bar, n789bar, n790bar, n791bar, n792bar, n793bar, n794bar, n795bar, n796bar, n797bar, n798bar, n799bar, n800bar, n801bar, n802bar, n803bar, n804bar, n805bar, n806bar, n807bar, n808bar, n809bar, n810bar, n811bar, n812bar, n813bar, n814bar, n815bar, n816bar, n817bar, n818bar, n819bar, n820bar, n821bar, n822bar, n823bar, n824bar, n825bar, n826bar, n827bar, n828bar, n829bar, n830bar, n831bar, n832bar, n833bar, n834bar, n835bar, n836bar, n837bar, n838bar, n839bar, n840bar, n841bar, n842bar, n843bar, n844bar, n845bar, n846bar, n847bar, n848bar, n849bar, n850bar, n851bar, n852bar, n853bar, n854bar, n855bar, n856bar, n857bar, n858bar, n859bar, n860bar, n861bar, n862bar, n863bar, n864bar, n865bar, n866bar, n867bar, n868bar, n869bar, n870bar, n871bar, n872bar, n873bar, n874bar, n875bar, n876bar, n877bar, n878bar, n879bar, n880bar, n881bar, n882bar, n883bar, n884bar, n885bar, n886bar, n887bar, n888bar, n889bar, n890bar, n891bar, n892bar, n893bar, n894bar, n895bar, n896bar, n897bar, n898bar, n899bar, n900bar, n901bar, n902bar, n903bar, n904bar, n905bar, n906bar, n907bar, n908bar, n909bar, n910bar, n911bar, n912bar, n913bar, n914bar, n915bar, n916bar, n917bar, n918bar, n919bar, n920bar, n921bar, n922bar, n923bar, n924bar, n925bar, n926bar, n927bar, n928bar, n929bar, n930bar, n931bar, n932bar, n933bar, n934bar, n935bar, n936bar, n937bar, n938bar, n939bar, n940bar, n941bar, n942bar, n943bar, n944bar, n945bar, n946bar, n947bar, n948bar, n949bar, n950bar, n951bar, n952bar, n953bar, n954bar, n955bar, n956bar, n957bar, n958bar, n959bar, n960bar, n961bar, n962bar, n963bar, n964bar, n965bar, n966bar, n967bar, n968bar, n969bar, n970bar, n971bar, n972bar;
  //wire_done

  assign in_81 = in[81];
  assign in_80 = in[80];
  assign in_79 = in[79];
  assign in_78 = in[78];
  assign in_77 = in[77];
  assign in_76 = in[76];
  assign in_75 = in[75];
  assign in_74 = in[74];
  assign in_73 = in[73];
  assign in_72 = in[72];
  assign in_71 = in[71];
  assign in_70 = in[70];
  assign in_69 = in[69];
  assign in_68 = in[68];
  assign in_67 = in[67];
  assign in_66 = in[66];
  assign in_65 = in[65];
  assign in_64 = in[64];
  assign in_63 = in[63];
  assign in_62 = in[62];
  assign in_61 = in[61];
  assign in_60 = in[60];
  assign in_59 = in[59];
  assign in_58 = in[58];
  assign in_57 = in[57];
  assign in_56 = in[56];
  assign in_55 = in[55];
  assign in_54 = in[54];
  assign in_53 = in[53];
  assign in_52 = in[52];
  assign in_51 = in[51];
  assign in_50 = in[50];
  assign in_49 = in[49];
  assign in_48 = in[48];
  assign in_47 = in[47];
  assign in_46 = in[46];
  assign in_45 = in[45];
  assign in_44 = in[44];
  assign in_43 = in[43];
  assign in_42 = in[42];
  assign in_41 = in[41];
  assign in_40 = in[40];
  assign in_39 = in[39];
  assign in_38 = in[38];
  assign in_37 = in[37];
  assign in_36 = in[36];
  assign in_35 = in[35];
  assign in_34 = in[34];
  assign in_33 = in[33];
  assign in_32 = in[32];
  assign in_31 = in[31];
  assign in_30 = in[30];
  assign in_29 = in[29];
  assign in_28 = in[28];
  assign in_27 = in[27];
  assign in_26 = in[26];
  assign in_25 = in[25];
  assign in_24 = in[24];
  assign in_23 = in[23];
  assign in_22 = in[22];
  assign in_21 = in[21];
  assign in_20 = in[20];
  assign in_19 = in[19];
  assign in_18 = in[18];
  assign in_17 = in[17];
  assign in_16 = in[16];
  assign in_15 = in[15];
  assign in_14 = in[14];
  assign in_13 = in[13];
  assign in_12 = in[12];
  assign in_11 = in[11];
  assign in_10 = in[10];
  assign in_9 = in[9];
  assign in_8 = in[8];
  assign in_7 = in[7];
  assign in_6 = in[6];
  assign in_5 = in[5];
  assign in_4 = in[4];
  assign in_3 = in[3];
  assign in_2 = in[2];
  assign in_1 = in[1];
  assign in_0 = in[0];

  OR2_X1 U1 ( .A1(n972), .A2(n971), .ZN(out[7]) );
  AND2_X1 U1bar ( .A1(n972bar), .A2(n971bar), .ZN(outbar[7]);
  OR2_X1 U2 ( .A1(n970), .A2(n969), .ZN(n971) );
  AND2_X1 U2bar ( .A1(n970bar), .A2(n969bar), .ZN(n971bar);
  OR2_X1 U3 ( .A1(n968), .A2(n967), .ZN(n969) );
  AND2_X1 U3bar ( .A1(n968bar), .A2(n967bar), .ZN(n969bar);
  OR2_X1 U4 ( .A1(n966), .A2(n965), .ZN(n967) );
  AND2_X1 U4bar ( .A1(n966bar), .A2(n965bar), .ZN(n967bar);
  OR2_X1 U5 ( .A1(n964), .A2(n963), .ZN(n968) );
  AND2_X1 U5bar ( .A1(n964bar), .A2(n963bar), .ZN(n968bar);
  OR2_X1 U6 ( .A1(in[116]), .A2(n962), .ZN(n963) );
  AND2_X1 U6bar ( .A1(inbar[116]), .A2(n962bar), .ZN(n963bar);
  OR2_X1 U7 ( .A1(n961), .A2(n960), .ZN(n970) );
  AND2_X1 U7bar ( .A1(n961bar), .A2(n960bar), .ZN(n970bar);
  OR2_X1 U8 ( .A1(in[150]), .A2(in[127]), .ZN(n960) );
  AND2_X1 U8bar ( .A1(inbar[150]), .A2(inbar[127]), .ZN(n960bar);
  OR2_X1 U9 ( .A1(in[160]), .A2(n959), .ZN(n961) );
  AND2_X1 U9bar ( .A1(inbar[160]), .A2(n959bar), .ZN(n961bar);
  OR2_X1 U10 ( .A1(in[252]), .A2(in[168]), .ZN(n959) );
  AND2_X1 U10bar ( .A1(inbar[252]), .A2(inbar[168]), .ZN(n959bar);
  OR2_X1 U11 ( .A1(n958), .A2(n957), .ZN(n972) );
  AND2_X1 U11bar ( .A1(n958bar), .A2(n957bar), .ZN(n972bar);
  OR2_X1 U12 ( .A1(n956), .A2(n955), .ZN(n957) );
  AND2_X1 U12bar ( .A1(n956bar), .A2(n955bar), .ZN(n957bar);
  OR2_X1 U13 ( .A1(in_17), .A2(in[96]), .ZN(n955) );
  AND2_X1 U13bar ( .A1(in_17bar), .A2(inbar[96]), .ZN(n955bar);
  OR2_X1 U14 ( .A1(in_23), .A2(n954), .ZN(n956) );
  AND2_X1 U14bar ( .A1(in_23bar), .A2(n954bar), .ZN(n956bar);
  OR2_X1 U15 ( .A1(in_31), .A2(in_26), .ZN(n954) );
  AND2_X1 U15bar ( .A1(in_31bar), .A2(in_26bar), .ZN(n954bar);
  OR2_X1 U16 ( .A1(n953), .A2(n952), .ZN(n958) );
  AND2_X1 U16bar ( .A1(n953bar), .A2(n952bar), .ZN(n958bar);
  OR2_X1 U17 ( .A1(in_58), .A2(in_4), .ZN(n952) );
  AND2_X1 U17bar ( .A1(in_58bar), .A2(in_4bar), .ZN(n952bar);
  OR2_X1 U18 ( .A1(in_59), .A2(n951), .ZN(n953) );
  AND2_X1 U18bar ( .A1(in_59bar), .A2(n951bar), .ZN(n953bar);
  OR2_X1 U19 ( .A1(in_71), .A2(in_62), .ZN(n951) );
  AND2_X1 U19bar ( .A1(in_71bar), .A2(in_62bar), .ZN(n951bar);
  OR2_X1 U20 ( .A1(n950), .A2(n949), .ZN(out[6]) );
  AND2_X1 U20bar ( .A1(n950bar), .A2(n949bar), .ZN(outbar[6]);
  OR2_X1 U21 ( .A1(n948), .A2(n947), .ZN(n949) );
  AND2_X1 U21bar ( .A1(n948bar), .A2(n947bar), .ZN(n949bar);
  OR2_X1 U22 ( .A1(n946), .A2(n945), .ZN(n947) );
  AND2_X1 U22bar ( .A1(n946bar), .A2(n945bar), .ZN(n947bar);
  OR2_X1 U23 ( .A1(n944), .A2(n943), .ZN(n945) );
  AND2_X1 U23bar ( .A1(n944bar), .A2(n943bar), .ZN(n945bar);
  OR2_X1 U24 ( .A1(n942), .A2(n941), .ZN(n946) );
  AND2_X1 U24bar ( .A1(n942bar), .A2(n941bar), .ZN(n946bar);
  OR2_X1 U25 ( .A1(in[101]), .A2(n940), .ZN(n941) );
  AND2_X1 U25bar ( .A1(inbar[101]), .A2(n940bar), .ZN(n941bar);
  OR2_X1 U26 ( .A1(n939), .A2(n938), .ZN(n948) );
  AND2_X1 U26bar ( .A1(n939bar), .A2(n938bar), .ZN(n948bar);
  OR2_X1 U27 ( .A1(in[114]), .A2(in[104]), .ZN(n938) );
  AND2_X1 U27bar ( .A1(inbar[114]), .A2(inbar[104]), .ZN(n938bar);
  OR2_X1 U28 ( .A1(in[128]), .A2(n937), .ZN(n939) );
  AND2_X1 U28bar ( .A1(inbar[128]), .A2(n937bar), .ZN(n939bar);
  OR2_X1 U29 ( .A1(in[136]), .A2(in[134]), .ZN(n937) );
  AND2_X1 U29bar ( .A1(inbar[136]), .A2(inbar[134]), .ZN(n937bar);
  OR2_X1 U30 ( .A1(n936), .A2(n935), .ZN(n950) );
  AND2_X1 U30bar ( .A1(n936bar), .A2(n935bar), .ZN(n950bar);
  OR2_X1 U31 ( .A1(n934), .A2(n933), .ZN(n935) );
  AND2_X1 U31bar ( .A1(n934bar), .A2(n933bar), .ZN(n935bar);
  OR2_X1 U32 ( .A1(in[177]), .A2(in[164]), .ZN(n933) );
  AND2_X1 U32bar ( .A1(inbar[177]), .A2(inbar[164]), .ZN(n933bar);
  OR2_X1 U33 ( .A1(in[212]), .A2(n932), .ZN(n934) );
  AND2_X1 U33bar ( .A1(inbar[212]), .A2(n932bar), .ZN(n934bar);
  OR2_X1 U34 ( .A1(in[248]), .A2(in[221]), .ZN(n932) );
  AND2_X1 U34bar ( .A1(inbar[248]), .A2(inbar[221]), .ZN(n932bar);
  OR2_X1 U35 ( .A1(n931), .A2(n930), .ZN(n936) );
  AND2_X1 U35bar ( .A1(n931bar), .A2(n930bar), .ZN(n936bar);
  OR2_X1 U36 ( .A1(in_18), .A2(in[93]), .ZN(n930) );
  AND2_X1 U36bar ( .A1(in_18bar), .A2(inbar[93]), .ZN(n930bar);
  OR2_X1 U37 ( .A1(in_31), .A2(n929), .ZN(n931) );
  AND2_X1 U37bar ( .A1(in_31bar), .A2(n929bar), .ZN(n931bar);
  OR2_X1 U38 ( .A1(in_7), .A2(in_39), .ZN(n929) );
  AND2_X1 U38bar ( .A1(in_7bar), .A2(in_39bar), .ZN(n929bar);
  OR2_X1 U39 ( .A1(n928), .A2(n927), .ZN(out[5]) );
  AND2_X1 U39bar ( .A1(n928bar), .A2(n927bar), .ZN(outbar[5]);
  OR2_X1 U40 ( .A1(n926), .A2(n925), .ZN(n927) );
  AND2_X1 U40bar ( .A1(n926bar), .A2(n925bar), .ZN(n927bar);
  OR2_X1 U41 ( .A1(n924), .A2(n923), .ZN(n925) );
  AND2_X1 U41bar ( .A1(n924bar), .A2(n923bar), .ZN(n925bar);
  OR2_X1 U42 ( .A1(n922), .A2(n921), .ZN(n923) );
  AND2_X1 U42bar ( .A1(n922bar), .A2(n921bar), .ZN(n923bar);
  OR2_X1 U43 ( .A1(n940), .A2(n920), .ZN(n924) );
  AND2_X1 U43bar ( .A1(n940bar), .A2(n920bar), .ZN(n924bar);
  OR2_X1 U44 ( .A1(in[111]), .A2(n919), .ZN(n920) );
  AND2_X1 U44bar ( .A1(inbar[111]), .A2(n919bar), .ZN(n920bar);
  OR2_X1 U45 ( .A1(n918), .A2(n917), .ZN(n940) );
  AND2_X1 U45bar ( .A1(n918bar), .A2(n917bar), .ZN(n940bar);
  OR2_X1 U46 ( .A1(n916), .A2(n915), .ZN(n917) );
  AND2_X1 U46bar ( .A1(n916bar), .A2(n915bar), .ZN(n917bar);
  OR2_X1 U47 ( .A1(n914), .A2(n913), .ZN(n915) );
  AND2_X1 U47bar ( .A1(n914bar), .A2(n913bar), .ZN(n915bar);
  OR2_X1 U48 ( .A1(in[140]), .A2(in[131]), .ZN(n913) );
  AND2_X1 U48bar ( .A1(inbar[140]), .A2(inbar[131]), .ZN(n913bar);
  OR2_X1 U49 ( .A1(in[160]), .A2(in[144]), .ZN(n914) );
  AND2_X1 U49bar ( .A1(inbar[160]), .A2(inbar[144]), .ZN(n914bar);
  OR2_X1 U50 ( .A1(n912), .A2(n911), .ZN(n916) );
  AND2_X1 U50bar ( .A1(n912bar), .A2(n911bar), .ZN(n916bar);
  OR2_X1 U51 ( .A1(in[179]), .A2(in[174]), .ZN(n911) );
  AND2_X1 U51bar ( .A1(inbar[179]), .A2(inbar[174]), .ZN(n911bar);
  OR2_X1 U52 ( .A1(in[188]), .A2(in[184]), .ZN(n912) );
  AND2_X1 U52bar ( .A1(inbar[188]), .A2(inbar[184]), .ZN(n912bar);
  OR2_X1 U53 ( .A1(n910), .A2(n909), .ZN(n918) );
  AND2_X1 U53bar ( .A1(n910bar), .A2(n909bar), .ZN(n918bar);
  OR2_X1 U54 ( .A1(n908), .A2(n907), .ZN(n909) );
  AND2_X1 U54bar ( .A1(n908bar), .A2(n907bar), .ZN(n909bar);
  OR2_X1 U55 ( .A1(in[216]), .A2(in[200]), .ZN(n907) );
  AND2_X1 U55bar ( .A1(inbar[216]), .A2(inbar[200]), .ZN(n907bar);
  OR2_X1 U56 ( .A1(in[228]), .A2(in[224]), .ZN(n908) );
  AND2_X1 U56bar ( .A1(inbar[228]), .A2(inbar[224]), .ZN(n908bar);
  OR2_X1 U57 ( .A1(n906), .A2(n905), .ZN(n910) );
  AND2_X1 U57bar ( .A1(n906bar), .A2(n905bar), .ZN(n910bar);
  OR2_X1 U58 ( .A1(in[247]), .A2(in[235]), .ZN(n905) );
  AND2_X1 U58bar ( .A1(inbar[247]), .A2(inbar[235]), .ZN(n905bar);
  OR2_X1 U59 ( .A1(in_42), .A2(in[83]), .ZN(n906) );
  AND2_X1 U59bar ( .A1(in_42bar), .A2(inbar[83]), .ZN(n906bar);
  OR2_X1 U60 ( .A1(n904), .A2(n903), .ZN(n926) );
  AND2_X1 U60bar ( .A1(n904bar), .A2(n903bar), .ZN(n926bar);
  OR2_X1 U61 ( .A1(in[166]), .A2(in[123]), .ZN(n903) );
  AND2_X1 U61bar ( .A1(inbar[166]), .A2(inbar[123]), .ZN(n903bar);
  OR2_X1 U62 ( .A1(in[170]), .A2(n902), .ZN(n904) );
  AND2_X1 U62bar ( .A1(inbar[170]), .A2(n902bar), .ZN(n904bar);
  OR2_X1 U63 ( .A1(in[194]), .A2(in[183]), .ZN(n902) );
  AND2_X1 U63bar ( .A1(inbar[194]), .A2(inbar[183]), .ZN(n902bar);
  OR2_X1 U64 ( .A1(n901), .A2(n900), .ZN(n928) );
  AND2_X1 U64bar ( .A1(n901bar), .A2(n900bar), .ZN(n928bar);
  OR2_X1 U65 ( .A1(n899), .A2(n898), .ZN(n900) );
  AND2_X1 U65bar ( .A1(n899bar), .A2(n898bar), .ZN(n900bar);
  OR2_X1 U66 ( .A1(in[241]), .A2(in[238]), .ZN(n898) );
  AND2_X1 U66bar ( .A1(inbar[241]), .A2(inbar[238]), .ZN(n898bar);
  OR2_X1 U67 ( .A1(in[250]), .A2(n897), .ZN(n899) );
  AND2_X1 U67bar ( .A1(inbar[250]), .A2(n897bar), .ZN(n899bar);
  OR2_X1 U68 ( .A1(in_24), .A2(in[84]), .ZN(n897) );
  AND2_X1 U68bar ( .A1(in_24bar), .A2(inbar[84]), .ZN(n897bar);
  OR2_X1 U69 ( .A1(n896), .A2(n895), .ZN(n901) );
  AND2_X1 U69bar ( .A1(n896bar), .A2(n895bar), .ZN(n901bar);
  OR2_X1 U70 ( .A1(in_41), .A2(in_29), .ZN(n895) );
  AND2_X1 U70bar ( .A1(in_41bar), .A2(in_29bar), .ZN(n895bar);
  OR2_X1 U71 ( .A1(in_66), .A2(n894), .ZN(n896) );
  AND2_X1 U71bar ( .A1(in_66bar), .A2(n894bar), .ZN(n896bar);
  OR2_X1 U72 ( .A1(in_76), .A2(in_71), .ZN(n894) );
  AND2_X1 U72bar ( .A1(in_76bar), .A2(in_71bar), .ZN(n894bar);
  OR2_X1 U73 ( .A1(n893), .A2(n892), .ZN(out[4]) );
  AND2_X1 U73bar ( .A1(n893bar), .A2(n892bar), .ZN(outbar[4]);
  OR2_X1 U74 ( .A1(n891), .A2(n890), .ZN(n892) );
  AND2_X1 U74bar ( .A1(n891bar), .A2(n890bar), .ZN(n892bar);
  OR2_X1 U75 ( .A1(n889), .A2(n888), .ZN(n890) );
  AND2_X1 U75bar ( .A1(n889bar), .A2(n888bar), .ZN(n890bar);
  OR2_X1 U76 ( .A1(n922), .A2(n887), .ZN(n888) );
  AND2_X1 U76bar ( .A1(n922bar), .A2(n887bar), .ZN(n888bar);
  OR2_X1 U77 ( .A1(n886), .A2(n885), .ZN(n922) );
  AND2_X1 U77bar ( .A1(n886bar), .A2(n885bar), .ZN(n922bar);
  OR2_X1 U78 ( .A1(n884), .A2(n883), .ZN(n885) );
  AND2_X1 U78bar ( .A1(n884bar), .A2(n883bar), .ZN(n885bar);
  OR2_X1 U79 ( .A1(n882), .A2(n881), .ZN(n883) );
  AND2_X1 U79bar ( .A1(n882bar), .A2(n881bar), .ZN(n883bar);
  OR2_X1 U80 ( .A1(in[118]), .A2(in[109]), .ZN(n881) );
  AND2_X1 U80bar ( .A1(inbar[118]), .A2(inbar[109]), .ZN(n881bar);
  OR2_X1 U81 ( .A1(in[139]), .A2(in[120]), .ZN(n882) );
  AND2_X1 U81bar ( .A1(inbar[139]), .A2(inbar[120]), .ZN(n882bar);
  OR2_X1 U82 ( .A1(n880), .A2(n879), .ZN(n884) );
  AND2_X1 U82bar ( .A1(n880bar), .A2(n879bar), .ZN(n884bar);
  OR2_X1 U83 ( .A1(in[198]), .A2(in[154]), .ZN(n879) );
  AND2_X1 U83bar ( .A1(inbar[198]), .A2(inbar[154]), .ZN(n879bar);
  OR2_X1 U84 ( .A1(in[210]), .A2(in[205]), .ZN(n880) );
  AND2_X1 U84bar ( .A1(inbar[210]), .A2(inbar[205]), .ZN(n880bar);
  OR2_X1 U85 ( .A1(n878), .A2(n877), .ZN(n886) );
  AND2_X1 U85bar ( .A1(n878bar), .A2(n877bar), .ZN(n886bar);
  OR2_X1 U86 ( .A1(n876), .A2(n875), .ZN(n877) );
  AND2_X1 U86bar ( .A1(n876bar), .A2(n875bar), .ZN(n877bar);
  OR2_X1 U87 ( .A1(in[219]), .A2(in[217]), .ZN(n875) );
  AND2_X1 U87bar ( .A1(inbar[219]), .A2(inbar[217]), .ZN(n875bar);
  OR2_X1 U88 ( .A1(in[86]), .A2(in[252]), .ZN(n876) );
  AND2_X1 U88bar ( .A1(inbar[86]), .A2(inbar[252]), .ZN(n876bar);
  OR2_X1 U89 ( .A1(n874), .A2(n873), .ZN(n878) );
  AND2_X1 U89bar ( .A1(n874bar), .A2(n873bar), .ZN(n878bar);
  OR2_X1 U90 ( .A1(in_40), .A2(in[91]), .ZN(n873) );
  AND2_X1 U90bar ( .A1(in_40bar), .A2(inbar[91]), .ZN(n873bar);
  OR2_X1 U91 ( .A1(in_8), .A2(in_46), .ZN(n874) );
  AND2_X1 U91bar ( .A1(in_8bar), .A2(in_46bar), .ZN(n874bar);
  OR2_X1 U92 ( .A1(n872), .A2(n871), .ZN(n889) );
  AND2_X1 U92bar ( .A1(n872bar), .A2(n871bar), .ZN(n889bar);
  OR2_X1 U93 ( .A1(in[117]), .A2(n943), .ZN(n871) );
  AND2_X1 U93bar ( .A1(inbar[117]), .A2(n943bar), .ZN(n871bar);
  OR2_X1 U94 ( .A1(n870), .A2(n869), .ZN(n943) );
  AND2_X1 U94bar ( .A1(n870bar), .A2(n869bar), .ZN(n943bar);
  OR2_X1 U95 ( .A1(n868), .A2(n867), .ZN(n869) );
  AND2_X1 U95bar ( .A1(n868bar), .A2(n867bar), .ZN(n869bar);
  OR2_X1 U96 ( .A1(n866), .A2(n865), .ZN(n867) );
  AND2_X1 U96bar ( .A1(n866bar), .A2(n865bar), .ZN(n867bar);
  OR2_X1 U97 ( .A1(n864), .A2(n863), .ZN(n865) );
  AND2_X1 U97bar ( .A1(n864bar), .A2(n863bar), .ZN(n865bar);
  OR2_X1 U98 ( .A1(in[108]), .A2(n919), .ZN(n866) );
  AND2_X1 U98bar ( .A1(inbar[108]), .A2(n919bar), .ZN(n866bar);
  OR2_X1 U99 ( .A1(n862), .A2(n861), .ZN(n919) );
  AND2_X1 U99bar ( .A1(n862bar), .A2(n861bar), .ZN(n919bar);
  OR2_X1 U100 ( .A1(n860), .A2(n859), .ZN(n861) );
  AND2_X1 U100bar ( .A1(n860bar), .A2(n859bar), .ZN(n861bar);
  OR2_X1 U101 ( .A1(n858), .A2(n857), .ZN(n859) );
  AND2_X1 U101bar ( .A1(n858bar), .A2(n857bar), .ZN(n859bar);
  OR2_X1 U102 ( .A1(in[119]), .A2(in[105]), .ZN(n857) );
  AND2_X1 U102bar ( .A1(inbar[119]), .A2(inbar[105]), .ZN(n857bar);
  OR2_X1 U103 ( .A1(in[186]), .A2(in[175]), .ZN(n858) );
  AND2_X1 U103bar ( .A1(inbar[186]), .A2(inbar[175]), .ZN(n858bar);
  OR2_X1 U104 ( .A1(n856), .A2(n855), .ZN(n860) );
  AND2_X1 U104bar ( .A1(n856bar), .A2(n855bar), .ZN(n860bar);
  OR2_X1 U105 ( .A1(in[202]), .A2(in[193]), .ZN(n855) );
  AND2_X1 U105bar ( .A1(inbar[202]), .A2(inbar[193]), .ZN(n855bar);
  OR2_X1 U106 ( .A1(in[225]), .A2(in[208]), .ZN(n856) );
  AND2_X1 U106bar ( .A1(inbar[225]), .A2(inbar[208]), .ZN(n856bar);
  OR2_X1 U107 ( .A1(n854), .A2(n853), .ZN(n862) );
  AND2_X1 U107bar ( .A1(n854bar), .A2(n853bar), .ZN(n862bar);
  OR2_X1 U108 ( .A1(n852), .A2(n851), .ZN(n853) );
  AND2_X1 U108bar ( .A1(n852bar), .A2(n851bar), .ZN(n853bar);
  OR2_X1 U109 ( .A1(in_1), .A2(in[85]), .ZN(n851) );
  AND2_X1 U109bar ( .A1(in_1bar), .A2(inbar[85]), .ZN(n851bar);
  OR2_X1 U110 ( .A1(in_23), .A2(in_19), .ZN(n852) );
  AND2_X1 U110bar ( .A1(in_23bar), .A2(in_19bar), .ZN(n852bar);
  OR2_X1 U111 ( .A1(n850), .A2(n849), .ZN(n854) );
  AND2_X1 U111bar ( .A1(n850bar), .A2(n849bar), .ZN(n854bar);
  OR2_X1 U112 ( .A1(in_43), .A2(in_33), .ZN(n849) );
  AND2_X1 U112bar ( .A1(in_43bar), .A2(in_33bar), .ZN(n849bar);
  OR2_X1 U113 ( .A1(in_63), .A2(in_44), .ZN(n850) );
  AND2_X1 U113bar ( .A1(in_63bar), .A2(in_44bar), .ZN(n850bar);
  OR2_X1 U114 ( .A1(n848), .A2(n847), .ZN(n868) );
  AND2_X1 U114bar ( .A1(n848bar), .A2(n847bar), .ZN(n868bar);
  OR2_X1 U115 ( .A1(in[141]), .A2(in[112]), .ZN(n847) );
  AND2_X1 U115bar ( .A1(inbar[141]), .A2(inbar[112]), .ZN(n847bar);
  OR2_X1 U116 ( .A1(in[147]), .A2(n846), .ZN(n848) );
  AND2_X1 U116bar ( .A1(inbar[147]), .A2(n846bar), .ZN(n848bar);
  OR2_X1 U117 ( .A1(in[181]), .A2(in[167]), .ZN(n846) );
  AND2_X1 U117bar ( .A1(inbar[181]), .A2(inbar[167]), .ZN(n846bar);
  OR2_X1 U118 ( .A1(n845), .A2(n844), .ZN(n870) );
  AND2_X1 U118bar ( .A1(n845bar), .A2(n844bar), .ZN(n870bar);
  OR2_X1 U119 ( .A1(n843), .A2(n842), .ZN(n844) );
  AND2_X1 U119bar ( .A1(n843bar), .A2(n842bar), .ZN(n844bar);
  OR2_X1 U120 ( .A1(in[229]), .A2(in[201]), .ZN(n842) );
  AND2_X1 U120bar ( .A1(inbar[229]), .A2(inbar[201]), .ZN(n842bar);
  OR2_X1 U121 ( .A1(in[237]), .A2(n841), .ZN(n843) );
  AND2_X1 U121bar ( .A1(inbar[237]), .A2(n841bar), .ZN(n843bar);
  OR2_X1 U122 ( .A1(in[94]), .A2(in[253]), .ZN(n841) );
  AND2_X1 U122bar ( .A1(inbar[94]), .A2(inbar[253]), .ZN(n841bar);
  OR2_X1 U123 ( .A1(n840), .A2(n839), .ZN(n845) );
  AND2_X1 U123bar ( .A1(n840bar), .A2(n839bar), .ZN(n845bar);
  OR2_X1 U124 ( .A1(in_21), .A2(in[96]), .ZN(n839) );
  AND2_X1 U124bar ( .A1(in_21bar), .A2(inbar[96]), .ZN(n839bar);
  OR2_X1 U125 ( .A1(in_25), .A2(n838), .ZN(n840) );
  AND2_X1 U125bar ( .A1(in_25bar), .A2(n838bar), .ZN(n840bar);
  OR2_X1 U126 ( .A1(in_81), .A2(in_45), .ZN(n838) );
  AND2_X1 U126bar ( .A1(in_81bar), .A2(in_45bar), .ZN(n838bar);
  OR2_X1 U127 ( .A1(n837), .A2(n836), .ZN(n891) );
  AND2_X1 U127bar ( .A1(n837bar), .A2(n836bar), .ZN(n891bar);
  OR2_X1 U128 ( .A1(in[142]), .A2(in[124]), .ZN(n836) );
  AND2_X1 U128bar ( .A1(inbar[142]), .A2(inbar[124]), .ZN(n836bar);
  OR2_X1 U129 ( .A1(in[150]), .A2(n835), .ZN(n837) );
  AND2_X1 U129bar ( .A1(inbar[150]), .A2(n835bar), .ZN(n837bar);
  OR2_X1 U130 ( .A1(in[172]), .A2(in[155]), .ZN(n835) );
  AND2_X1 U130bar ( .A1(inbar[172]), .A2(inbar[155]), .ZN(n835bar);
  OR2_X1 U131 ( .A1(n834), .A2(n833), .ZN(n893) );
  AND2_X1 U131bar ( .A1(n834bar), .A2(n833bar), .ZN(n893bar);
  OR2_X1 U132 ( .A1(n832), .A2(n831), .ZN(n833) );
  AND2_X1 U132bar ( .A1(n832bar), .A2(n831bar), .ZN(n833bar);
  OR2_X1 U133 ( .A1(in[196]), .A2(in[173]), .ZN(n831) );
  AND2_X1 U133bar ( .A1(inbar[196]), .A2(inbar[173]), .ZN(n831bar);
  OR2_X1 U134 ( .A1(in[222]), .A2(n830), .ZN(n832) );
  AND2_X1 U134bar ( .A1(inbar[222]), .A2(n830bar), .ZN(n832bar);
  OR2_X1 U135 ( .A1(in[227]), .A2(in[226]), .ZN(n830) );
  AND2_X1 U135bar ( .A1(inbar[227]), .A2(inbar[226]), .ZN(n830bar);
  OR2_X1 U136 ( .A1(n829), .A2(n828), .ZN(n834) );
  AND2_X1 U136bar ( .A1(n829bar), .A2(n828bar), .ZN(n834bar);
  OR2_X1 U137 ( .A1(in[249]), .A2(in[231]), .ZN(n828) );
  AND2_X1 U137bar ( .A1(inbar[249]), .A2(inbar[231]), .ZN(n828bar);
  OR2_X1 U138 ( .A1(in_28), .A2(n827), .ZN(n829) );
  AND2_X1 U138bar ( .A1(in_28bar), .A2(n827bar), .ZN(n829bar);
  OR2_X1 U139 ( .A1(in_52), .A2(in_47), .ZN(n827) );
  AND2_X1 U139bar ( .A1(in_52bar), .A2(in_47bar), .ZN(n827bar);
  OR2_X1 U140 ( .A1(n826), .A2(n825), .ZN(out[3]) );
  AND2_X1 U140bar ( .A1(n826bar), .A2(n825bar), .ZN(outbar[3]);
  OR2_X1 U141 ( .A1(n824), .A2(n823), .ZN(n825) );
  AND2_X1 U141bar ( .A1(n824bar), .A2(n823bar), .ZN(n825bar);
  OR2_X1 U142 ( .A1(n822), .A2(n821), .ZN(n823) );
  AND2_X1 U142bar ( .A1(n822bar), .A2(n821bar), .ZN(n823bar);
  OR2_X1 U143 ( .A1(n820), .A2(n819), .ZN(n821) );
  AND2_X1 U143bar ( .A1(n820bar), .A2(n819bar), .ZN(n821bar);
  OR2_X1 U144 ( .A1(n964), .A2(n818), .ZN(n822) );
  AND2_X1 U144bar ( .A1(n964bar), .A2(n818bar), .ZN(n822bar);
  OR2_X1 U145 ( .A1(in[118]), .A2(n817), .ZN(n818) );
  AND2_X1 U145bar ( .A1(inbar[118]), .A2(n817bar), .ZN(n818bar);
  OR2_X1 U146 ( .A1(n816), .A2(n815), .ZN(n964) );
  AND2_X1 U146bar ( .A1(n816bar), .A2(n815bar), .ZN(n964bar);
  OR2_X1 U147 ( .A1(n814), .A2(n813), .ZN(n815) );
  AND2_X1 U147bar ( .A1(n814bar), .A2(n813bar), .ZN(n815bar);
  OR2_X1 U148 ( .A1(n812), .A2(n811), .ZN(n813) );
  AND2_X1 U148bar ( .A1(n812bar), .A2(n811bar), .ZN(n813bar);
  OR2_X1 U149 ( .A1(in[122]), .A2(in[111]), .ZN(n811) );
  AND2_X1 U149bar ( .A1(inbar[122]), .A2(inbar[111]), .ZN(n811bar);
  OR2_X1 U150 ( .A1(in[154]), .A2(in[151]), .ZN(n812) );
  AND2_X1 U150bar ( .A1(inbar[154]), .A2(inbar[151]), .ZN(n812bar);
  OR2_X1 U151 ( .A1(n810), .A2(n809), .ZN(n814) );
  AND2_X1 U151bar ( .A1(n810bar), .A2(n809bar), .ZN(n814bar);
  OR2_X1 U152 ( .A1(in[187]), .A2(in[177]), .ZN(n809) );
  AND2_X1 U152bar ( .A1(inbar[187]), .A2(inbar[177]), .ZN(n809bar);
  OR2_X1 U153 ( .A1(in[200]), .A2(in[192]), .ZN(n810) );
  AND2_X1 U153bar ( .A1(inbar[200]), .A2(inbar[192]), .ZN(n810bar);
  OR2_X1 U154 ( .A1(n808), .A2(n807), .ZN(n816) );
  AND2_X1 U154bar ( .A1(n808bar), .A2(n807bar), .ZN(n816bar);
  OR2_X1 U155 ( .A1(n806), .A2(n805), .ZN(n807) );
  AND2_X1 U155bar ( .A1(n806bar), .A2(n805bar), .ZN(n807bar);
  OR2_X1 U156 ( .A1(in[225]), .A2(in[207]), .ZN(n805) );
  AND2_X1 U156bar ( .A1(inbar[225]), .A2(inbar[207]), .ZN(n805bar);
  OR2_X1 U157 ( .A1(in[98]), .A2(in[226]), .ZN(n806) );
  AND2_X1 U157bar ( .A1(inbar[98]), .A2(inbar[226]), .ZN(n806bar);
  OR2_X1 U158 ( .A1(n804), .A2(n803), .ZN(n808) );
  AND2_X1 U158bar ( .A1(n804bar), .A2(n803bar), .ZN(n808bar);
  OR2_X1 U159 ( .A1(in_20), .A2(in_16), .ZN(n803) );
  AND2_X1 U159bar ( .A1(in_20bar), .A2(in_16bar), .ZN(n803bar);
  OR2_X1 U160 ( .A1(in_55), .A2(in_45), .ZN(n804) );
  AND2_X1 U160bar ( .A1(in_55bar), .A2(in_45bar), .ZN(n804bar);
  OR2_X1 U161 ( .A1(n802), .A2(n801), .ZN(n824) );
  AND2_X1 U161bar ( .A1(n802bar), .A2(n801bar), .ZN(n824bar);
  OR2_X1 U162 ( .A1(in[162]), .A2(in[149]), .ZN(n801) );
  AND2_X1 U162bar ( .A1(inbar[162]), .A2(inbar[149]), .ZN(n801bar);
  OR2_X1 U163 ( .A1(in[163]), .A2(n800), .ZN(n802) );
  AND2_X1 U163bar ( .A1(inbar[163]), .A2(n800bar), .ZN(n802bar);
  OR2_X1 U164 ( .A1(in[191]), .A2(in[189]), .ZN(n800) );
  AND2_X1 U164bar ( .A1(inbar[191]), .A2(inbar[189]), .ZN(n800bar);
  OR2_X1 U165 ( .A1(n799), .A2(n798), .ZN(n826) );
  AND2_X1 U165bar ( .A1(n799bar), .A2(n798bar), .ZN(n826bar);
  OR2_X1 U166 ( .A1(n797), .A2(n796), .ZN(n798) );
  AND2_X1 U166bar ( .A1(n797bar), .A2(n796bar), .ZN(n798bar);
  OR2_X1 U167 ( .A1(in[212]), .A2(in[193]), .ZN(n796) );
  AND2_X1 U167bar ( .A1(inbar[212]), .A2(inbar[193]), .ZN(n796bar);
  OR2_X1 U168 ( .A1(in[238]), .A2(n795), .ZN(n797) );
  AND2_X1 U168bar ( .A1(inbar[238]), .A2(n795bar), .ZN(n797bar);
  OR2_X1 U169 ( .A1(in[88]), .A2(in[247]), .ZN(n795) );
  AND2_X1 U169bar ( .A1(inbar[88]), .A2(inbar[247]), .ZN(n795bar);
  OR2_X1 U170 ( .A1(n794), .A2(n793), .ZN(n799) );
  AND2_X1 U170bar ( .A1(n794bar), .A2(n793bar), .ZN(n799bar);
  OR2_X1 U171 ( .A1(in[94]), .A2(in[92]), .ZN(n793) );
  AND2_X1 U171bar ( .A1(inbar[94]), .A2(inbar[92]), .ZN(n793bar);
  OR2_X1 U172 ( .A1(in_52), .A2(n792), .ZN(n794) );
  AND2_X1 U172bar ( .A1(in_52bar), .A2(n792bar), .ZN(n794bar);
  OR2_X1 U173 ( .A1(in_70), .A2(in_67), .ZN(n792) );
  AND2_X1 U173bar ( .A1(in_70bar), .A2(in_67bar), .ZN(n792bar);
  OR2_X1 U174 ( .A1(n791), .A2(n790), .ZN(out[2]) );
  AND2_X1 U174bar ( .A1(n791bar), .A2(n790bar), .ZN(outbar[2]);
  OR2_X1 U175 ( .A1(n789), .A2(n788), .ZN(n790) );
  AND2_X1 U175bar ( .A1(n789bar), .A2(n788bar), .ZN(n790bar);
  OR2_X1 U176 ( .A1(n787), .A2(n786), .ZN(n788) );
  AND2_X1 U176bar ( .A1(n787bar), .A2(n786bar), .ZN(n788bar);
  OR2_X1 U177 ( .A1(n819), .A2(n785), .ZN(n786) );
  AND2_X1 U177bar ( .A1(n819bar), .A2(n785bar), .ZN(n786bar);
  OR2_X1 U178 ( .A1(n784), .A2(n783), .ZN(n819) );
  AND2_X1 U178bar ( .A1(n784bar), .A2(n783bar), .ZN(n819bar);
  OR2_X1 U179 ( .A1(n782), .A2(n781), .ZN(n783) );
  AND2_X1 U179bar ( .A1(n782bar), .A2(n781bar), .ZN(n783bar);
  OR2_X1 U180 ( .A1(n780), .A2(n779), .ZN(n781) );
  AND2_X1 U180bar ( .A1(n780bar), .A2(n779bar), .ZN(n781bar);
  OR2_X1 U181 ( .A1(n962), .A2(n778), .ZN(n779) );
  AND2_X1 U181bar ( .A1(n962bar), .A2(n778bar), .ZN(n779bar);
  OR2_X1 U182 ( .A1(n777), .A2(n776), .ZN(n962) );
  AND2_X1 U182bar ( .A1(n777bar), .A2(n776bar), .ZN(n962bar);
  OR2_X1 U183 ( .A1(n775), .A2(n774), .ZN(n776) );
  AND2_X1 U183bar ( .A1(n775bar), .A2(n774bar), .ZN(n776bar);
  OR2_X1 U184 ( .A1(n773), .A2(n772), .ZN(n774) );
  AND2_X1 U184bar ( .A1(n773bar), .A2(n772bar), .ZN(n774bar);
  OR2_X1 U185 ( .A1(in[131]), .A2(in[120]), .ZN(n772) );
  AND2_X1 U185bar ( .A1(inbar[131]), .A2(inbar[120]), .ZN(n772bar);
  OR2_X1 U186 ( .A1(in[153]), .A2(in[147]), .ZN(n773) );
  AND2_X1 U186bar ( .A1(inbar[153]), .A2(inbar[147]), .ZN(n773bar);
  OR2_X1 U187 ( .A1(n771), .A2(n770), .ZN(n775) );
  AND2_X1 U187bar ( .A1(n771bar), .A2(n770bar), .ZN(n775bar);
  OR2_X1 U188 ( .A1(in[170]), .A2(in[156]), .ZN(n770) );
  AND2_X1 U188bar ( .A1(inbar[170]), .A2(inbar[156]), .ZN(n770bar);
  OR2_X1 U189 ( .A1(in[223]), .A2(in[190]), .ZN(n771) );
  AND2_X1 U189bar ( .A1(inbar[223]), .A2(inbar[190]), .ZN(n771bar);
  OR2_X1 U190 ( .A1(n769), .A2(n768), .ZN(n777) );
  AND2_X1 U190bar ( .A1(n769bar), .A2(n768bar), .ZN(n777bar);
  OR2_X1 U191 ( .A1(n767), .A2(n766), .ZN(n768) );
  AND2_X1 U191bar ( .A1(n767bar), .A2(n766bar), .ZN(n768bar);
  OR2_X1 U192 ( .A1(in[236]), .A2(in[230]), .ZN(n766) );
  AND2_X1 U192bar ( .A1(inbar[236]), .A2(inbar[230]), .ZN(n766bar);
  OR2_X1 U193 ( .A1(in[85]), .A2(in[240]), .ZN(n767) );
  AND2_X1 U193bar ( .A1(inbar[85]), .A2(inbar[240]), .ZN(n767bar);
  OR2_X1 U194 ( .A1(n765), .A2(n764), .ZN(n769) );
  AND2_X1 U194bar ( .A1(n765bar), .A2(n764bar), .ZN(n769bar);
  OR2_X1 U195 ( .A1(in_12), .A2(in[90]), .ZN(n764) );
  AND2_X1 U195bar ( .A1(in_12bar), .A2(inbar[90]), .ZN(n764bar);
  OR2_X1 U196 ( .A1(in_39), .A2(in_28), .ZN(n765) );
  AND2_X1 U196bar ( .A1(in_39bar), .A2(in_28bar), .ZN(n765bar);
  OR2_X1 U197 ( .A1(in[109]), .A2(n763), .ZN(n780) );
  AND2_X1 U197bar ( .A1(inbar[109]), .A2(n763bar), .ZN(n780bar);
  OR2_X1 U198 ( .A1(n762), .A2(n761), .ZN(n782) );
  AND2_X1 U198bar ( .A1(n762bar), .A2(n761bar), .ZN(n782bar);
  OR2_X1 U199 ( .A1(in[138]), .A2(in[129]), .ZN(n761) );
  AND2_X1 U199bar ( .A1(inbar[138]), .A2(inbar[129]), .ZN(n761bar);
  OR2_X1 U200 ( .A1(in[157]), .A2(n760), .ZN(n762) );
  AND2_X1 U200bar ( .A1(inbar[157]), .A2(n760bar), .ZN(n762bar);
  OR2_X1 U201 ( .A1(in[182]), .A2(in[167]), .ZN(n760) );
  AND2_X1 U201bar ( .A1(inbar[182]), .A2(inbar[167]), .ZN(n760bar);
  OR2_X1 U202 ( .A1(n759), .A2(n758), .ZN(n784) );
  AND2_X1 U202bar ( .A1(n759bar), .A2(n758bar), .ZN(n784bar);
  OR2_X1 U203 ( .A1(n757), .A2(n756), .ZN(n758) );
  AND2_X1 U203bar ( .A1(n757bar), .A2(n756bar), .ZN(n758bar);
  OR2_X1 U204 ( .A1(in[195]), .A2(in[184]), .ZN(n756) );
  AND2_X1 U204bar ( .A1(inbar[195]), .A2(inbar[184]), .ZN(n756bar);
  OR2_X1 U205 ( .A1(in[196]), .A2(n755), .ZN(n757) );
  AND2_X1 U205bar ( .A1(inbar[196]), .A2(n755bar), .ZN(n757bar);
  OR2_X1 U206 ( .A1(in[215]), .A2(in[209]), .ZN(n755) );
  AND2_X1 U206bar ( .A1(inbar[215]), .A2(inbar[209]), .ZN(n755bar);
  OR2_X1 U207 ( .A1(n754), .A2(n753), .ZN(n759) );
  AND2_X1 U207bar ( .A1(n754bar), .A2(n753bar), .ZN(n759bar);
  OR2_X1 U208 ( .A1(in[93]), .A2(in[233]), .ZN(n753) );
  AND2_X1 U208bar ( .A1(inbar[93]), .A2(inbar[233]), .ZN(n753bar);
  OR2_X1 U209 ( .A1(in_1), .A2(n752), .ZN(n754) );
  AND2_X1 U209bar ( .A1(in_1bar), .A2(n752bar), .ZN(n754bar);
  OR2_X1 U210 ( .A1(in_69), .A2(in_66), .ZN(n752) );
  AND2_X1 U210bar ( .A1(in_69bar), .A2(in_66bar), .ZN(n752bar);
  OR2_X1 U211 ( .A1(n966), .A2(n751), .ZN(n787) );
  AND2_X1 U211bar ( .A1(n966bar), .A2(n751bar), .ZN(n787bar);
  OR2_X1 U212 ( .A1(in[134]), .A2(n750), .ZN(n751) );
  AND2_X1 U212bar ( .A1(inbar[134]), .A2(n750bar), .ZN(n751bar);
  OR2_X1 U213 ( .A1(n749), .A2(n748), .ZN(n966) );
  AND2_X1 U213bar ( .A1(n749bar), .A2(n748bar), .ZN(n966bar);
  OR2_X1 U214 ( .A1(n747), .A2(n746), .ZN(n748) );
  AND2_X1 U214bar ( .A1(n747bar), .A2(n746bar), .ZN(n748bar);
  OR2_X1 U215 ( .A1(n745), .A2(n744), .ZN(n746) );
  AND2_X1 U215bar ( .A1(n745bar), .A2(n744bar), .ZN(n746bar);
  OR2_X1 U216 ( .A1(in[136]), .A2(in[121]), .ZN(n744) );
  AND2_X1 U216bar ( .A1(inbar[136]), .A2(inbar[121]), .ZN(n744bar);
  OR2_X1 U217 ( .A1(in[186]), .A2(in[174]), .ZN(n745) );
  AND2_X1 U217bar ( .A1(inbar[186]), .A2(inbar[174]), .ZN(n745bar);
  OR2_X1 U218 ( .A1(n743), .A2(n742), .ZN(n747) );
  AND2_X1 U218bar ( .A1(n743bar), .A2(n742bar), .ZN(n747bar);
  OR2_X1 U219 ( .A1(in[198]), .A2(in[197]), .ZN(n742) );
  AND2_X1 U219bar ( .A1(inbar[198]), .A2(inbar[197]), .ZN(n742bar);
  OR2_X1 U220 ( .A1(in[214]), .A2(in[199]), .ZN(n743) );
  AND2_X1 U220bar ( .A1(inbar[214]), .A2(inbar[199]), .ZN(n743bar);
  OR2_X1 U221 ( .A1(n741), .A2(n740), .ZN(n749) );
  AND2_X1 U221bar ( .A1(n741bar), .A2(n740bar), .ZN(n749bar);
  OR2_X1 U222 ( .A1(n739), .A2(n738), .ZN(n740) );
  AND2_X1 U222bar ( .A1(n739bar), .A2(n738bar), .ZN(n740bar);
  OR2_X1 U223 ( .A1(in[231]), .A2(in[220]), .ZN(n738) );
  AND2_X1 U223bar ( .A1(inbar[231]), .A2(inbar[220]), .ZN(n738bar);
  OR2_X1 U224 ( .A1(in_25), .A2(in[245]), .ZN(n739) );
  AND2_X1 U224bar ( .A1(in_25bar), .A2(inbar[245]), .ZN(n739bar);
  OR2_X1 U225 ( .A1(n737), .A2(n736), .ZN(n741) );
  AND2_X1 U225bar ( .A1(n737bar), .A2(n736bar), .ZN(n741bar);
  OR2_X1 U226 ( .A1(in_53), .A2(in_29), .ZN(n736) );
  AND2_X1 U226bar ( .A1(in_53bar), .A2(in_29bar), .ZN(n736bar);
  OR2_X1 U227 ( .A1(in_79), .A2(in_74), .ZN(n737) );
  AND2_X1 U227bar ( .A1(in_79bar), .A2(in_74bar), .ZN(n737bar);
  OR2_X1 U228 ( .A1(n735), .A2(n734), .ZN(n789) );
  AND2_X1 U228bar ( .A1(n735bar), .A2(n734bar), .ZN(n789bar);
  OR2_X1 U229 ( .A1(in[152]), .A2(in[140]), .ZN(n734) );
  AND2_X1 U229bar ( .A1(inbar[152]), .A2(inbar[140]), .ZN(n734bar);
  OR2_X1 U230 ( .A1(in[155]), .A2(n733), .ZN(n735) );
  AND2_X1 U230bar ( .A1(inbar[155]), .A2(n733bar), .ZN(n735bar);
  OR2_X1 U231 ( .A1(in[166]), .A2(in[165]), .ZN(n733) );
  AND2_X1 U231bar ( .A1(inbar[166]), .A2(inbar[165]), .ZN(n733bar);
  OR2_X1 U232 ( .A1(n732), .A2(n731), .ZN(n791) );
  AND2_X1 U232bar ( .A1(n732bar), .A2(n731bar), .ZN(n791bar);
  OR2_X1 U233 ( .A1(n730), .A2(n729), .ZN(n731) );
  AND2_X1 U233bar ( .A1(n730bar), .A2(n729bar), .ZN(n731bar);
  OR2_X1 U234 ( .A1(in[202]), .A2(in[185]), .ZN(n729) );
  AND2_X1 U234bar ( .A1(inbar[202]), .A2(inbar[185]), .ZN(n729bar);
  OR2_X1 U235 ( .A1(in[211]), .A2(n728), .ZN(n730) );
  AND2_X1 U235bar ( .A1(inbar[211]), .A2(n728bar), .ZN(n730bar);
  OR2_X1 U236 ( .A1(in[255]), .A2(in[253]), .ZN(n728) );
  AND2_X1 U236bar ( .A1(inbar[255]), .A2(inbar[253]), .ZN(n728bar);
  OR2_X1 U237 ( .A1(n727), .A2(n726), .ZN(n732) );
  AND2_X1 U237bar ( .A1(n727bar), .A2(n726bar), .ZN(n732bar);
  OR2_X1 U238 ( .A1(in_35), .A2(in_15), .ZN(n726) );
  AND2_X1 U238bar ( .A1(in_35bar), .A2(in_15bar), .ZN(n726bar);
  OR2_X1 U239 ( .A1(in_36), .A2(n725), .ZN(n727) );
  AND2_X1 U239bar ( .A1(in_36bar), .A2(n725bar), .ZN(n727bar);
  OR2_X1 U240 ( .A1(in_48), .A2(in_40), .ZN(n725) );
  AND2_X1 U240bar ( .A1(in_48bar), .A2(in_40bar), .ZN(n725bar);
  OR2_X1 U241 ( .A1(n724), .A2(n723), .ZN(out[1]) );
  AND2_X1 U241bar ( .A1(n724bar), .A2(n723bar), .ZN(outbar[1]);
  OR2_X1 U242 ( .A1(n722), .A2(n721), .ZN(n723) );
  AND2_X1 U242bar ( .A1(n722bar), .A2(n721bar), .ZN(n723bar);
  OR2_X1 U243 ( .A1(n720), .A2(n719), .ZN(n721) );
  AND2_X1 U243bar ( .A1(n720bar), .A2(n719bar), .ZN(n721bar);
  OR2_X1 U244 ( .A1(n921), .A2(n887), .ZN(n719) );
  AND2_X1 U244bar ( .A1(n921bar), .A2(n887bar), .ZN(n719bar);
  OR2_X1 U245 ( .A1(n718), .A2(n717), .ZN(n887) );
  AND2_X1 U245bar ( .A1(n718bar), .A2(n717bar), .ZN(n887bar);
  OR2_X1 U246 ( .A1(n716), .A2(n715), .ZN(n717) );
  AND2_X1 U246bar ( .A1(n716bar), .A2(n715bar), .ZN(n717bar);
  OR2_X1 U247 ( .A1(n714), .A2(n713), .ZN(n715) );
  AND2_X1 U247bar ( .A1(n714bar), .A2(n713bar), .ZN(n715bar);
  OR2_X1 U248 ( .A1(in[116]), .A2(in[110]), .ZN(n713) );
  AND2_X1 U248bar ( .A1(inbar[116]), .A2(inbar[110]), .ZN(n713bar);
  OR2_X1 U249 ( .A1(in[133]), .A2(in[130]), .ZN(n714) );
  AND2_X1 U249bar ( .A1(inbar[133]), .A2(inbar[130]), .ZN(n714bar);
  OR2_X1 U250 ( .A1(n712), .A2(n711), .ZN(n716) );
  AND2_X1 U250bar ( .A1(n712bar), .A2(n711bar), .ZN(n716bar);
  OR2_X1 U251 ( .A1(in[203]), .A2(in[135]), .ZN(n711) );
  AND2_X1 U251bar ( .A1(inbar[203]), .A2(inbar[135]), .ZN(n711bar);
  OR2_X1 U252 ( .A1(in[232]), .A2(in[223]), .ZN(n712) );
  AND2_X1 U252bar ( .A1(inbar[232]), .A2(inbar[223]), .ZN(n712bar);
  OR2_X1 U253 ( .A1(n710), .A2(n709), .ZN(n718) );
  AND2_X1 U253bar ( .A1(n710bar), .A2(n709bar), .ZN(n718bar);
  OR2_X1 U254 ( .A1(n708), .A2(n707), .ZN(n709) );
  AND2_X1 U254bar ( .A1(n708bar), .A2(n707bar), .ZN(n709bar);
  OR2_X1 U255 ( .A1(in[255]), .A2(in[233]), .ZN(n707) );
  AND2_X1 U255bar ( .A1(inbar[255]), .A2(inbar[233]), .ZN(n707bar);
  OR2_X1 U256 ( .A1(in_53), .A2(in_34), .ZN(n708) );
  AND2_X1 U256bar ( .A1(in_53bar), .A2(in_34bar), .ZN(n708bar);
  OR2_X1 U257 ( .A1(n706), .A2(n705), .ZN(n710) );
  AND2_X1 U257bar ( .A1(n706bar), .A2(n705bar), .ZN(n710bar);
  OR2_X1 U258 ( .A1(in_57), .A2(in_55), .ZN(n705) );
  AND2_X1 U258bar ( .A1(in_57bar), .A2(in_55bar), .ZN(n705bar);
  OR2_X1 U259 ( .A1(in_68), .A2(in_67), .ZN(n706) );
  AND2_X1 U259bar ( .A1(in_68bar), .A2(in_67bar), .ZN(n706bar);
  OR2_X1 U260 ( .A1(n704), .A2(n703), .ZN(n921) );
  AND2_X1 U260bar ( .A1(n704bar), .A2(n703bar), .ZN(n921bar);
  OR2_X1 U261 ( .A1(n702), .A2(n701), .ZN(n703) );
  AND2_X1 U261bar ( .A1(n702bar), .A2(n701bar), .ZN(n703bar);
  OR2_X1 U262 ( .A1(n700), .A2(n699), .ZN(n701) );
  AND2_X1 U262bar ( .A1(n700bar), .A2(n699bar), .ZN(n701bar);
  OR2_X1 U263 ( .A1(n944), .A2(n872), .ZN(n699) );
  AND2_X1 U263bar ( .A1(n944bar), .A2(n872bar), .ZN(n699bar);
  OR2_X1 U264 ( .A1(n698), .A2(n697), .ZN(n872) );
  AND2_X1 U264bar ( .A1(n698bar), .A2(n697bar), .ZN(n872bar);
  OR2_X1 U265 ( .A1(n696), .A2(n695), .ZN(n697) );
  AND2_X1 U265bar ( .A1(n696bar), .A2(n695bar), .ZN(n697bar);
  OR2_X1 U266 ( .A1(n694), .A2(n693), .ZN(n695) );
  AND2_X1 U266bar ( .A1(n694bar), .A2(n693bar), .ZN(n695bar);
  OR2_X1 U267 ( .A1(in[121]), .A2(in[102]), .ZN(n693) );
  AND2_X1 U267bar ( .A1(inbar[121]), .A2(inbar[102]), .ZN(n693bar);
  OR2_X1 U268 ( .A1(in[162]), .A2(in[161]), .ZN(n694) );
  AND2_X1 U268bar ( .A1(inbar[162]), .A2(inbar[161]), .ZN(n694bar);
  OR2_X1 U269 ( .A1(n692), .A2(n691), .ZN(n696) );
  AND2_X1 U269bar ( .A1(n692bar), .A2(n691bar), .ZN(n696bar);
  OR2_X1 U270 ( .A1(in[192]), .A2(in[178]), .ZN(n691) );
  AND2_X1 U270bar ( .A1(inbar[192]), .A2(inbar[178]), .ZN(n691bar);
  OR2_X1 U271 ( .A1(in[244]), .A2(in[209]), .ZN(n692) );
  AND2_X1 U271bar ( .A1(inbar[244]), .A2(inbar[209]), .ZN(n692bar);
  OR2_X1 U272 ( .A1(n690), .A2(n689), .ZN(n698) );
  AND2_X1 U272bar ( .A1(n690bar), .A2(n689bar), .ZN(n698bar);
  OR2_X1 U273 ( .A1(n688), .A2(n687), .ZN(n689) );
  AND2_X1 U273bar ( .A1(n688bar), .A2(n687bar), .ZN(n689bar);
  OR2_X1 U274 ( .A1(in[90]), .A2(in[254]), .ZN(n687) );
  AND2_X1 U274bar ( .A1(inbar[90]), .A2(inbar[254]), .ZN(n687bar);
  OR2_X1 U275 ( .A1(in_36), .A2(in_32), .ZN(n688) );
  AND2_X1 U275bar ( .A1(in_36bar), .A2(in_32bar), .ZN(n688bar);
  OR2_X1 U276 ( .A1(n686), .A2(n685), .ZN(n690) );
  AND2_X1 U276bar ( .A1(n686bar), .A2(n685bar), .ZN(n690bar);
  OR2_X1 U277 ( .A1(in_62), .A2(in_37), .ZN(n685) );
  AND2_X1 U277bar ( .A1(in_62bar), .A2(in_37bar), .ZN(n685bar);
  OR2_X1 U278 ( .A1(in_75), .A2(in_73), .ZN(n686) );
  AND2_X1 U278bar ( .A1(in_75bar), .A2(in_73bar), .ZN(n686bar);
  OR2_X1 U279 ( .A1(n684), .A2(n683), .ZN(n944) );
  AND2_X1 U279bar ( .A1(n684bar), .A2(n683bar), .ZN(n944bar);
  OR2_X1 U280 ( .A1(n682), .A2(n681), .ZN(n683) );
  AND2_X1 U280bar ( .A1(n682bar), .A2(n681bar), .ZN(n683bar);
  OR2_X1 U281 ( .A1(n680), .A2(n679), .ZN(n681) );
  AND2_X1 U281bar ( .A1(n680bar), .A2(n679bar), .ZN(n681bar);
  OR2_X1 U282 ( .A1(in[171]), .A2(in[153]), .ZN(n679) );
  AND2_X1 U282bar ( .A1(inbar[171]), .A2(inbar[153]), .ZN(n679bar);
  OR2_X1 U283 ( .A1(in[187]), .A2(in[176]), .ZN(n680) );
  AND2_X1 U283bar ( .A1(inbar[187]), .A2(inbar[176]), .ZN(n680bar);
  OR2_X1 U284 ( .A1(n678), .A2(n677), .ZN(n682) );
  AND2_X1 U284bar ( .A1(n678bar), .A2(n677bar), .ZN(n682bar);
  OR2_X1 U285 ( .A1(in[245]), .A2(in[211]), .ZN(n677) );
  AND2_X1 U285bar ( .A1(inbar[245]), .A2(inbar[211]), .ZN(n677bar);
  OR2_X1 U286 ( .A1(in[97]), .A2(in[88]), .ZN(n678) );
  AND2_X1 U286bar ( .A1(inbar[97]), .A2(inbar[88]), .ZN(n678bar);
  OR2_X1 U287 ( .A1(n676), .A2(n675), .ZN(n684) );
  AND2_X1 U287bar ( .A1(n676bar), .A2(n675bar), .ZN(n684bar);
  OR2_X1 U288 ( .A1(n674), .A2(n673), .ZN(n675) );
  AND2_X1 U288bar ( .A1(n674bar), .A2(n673bar), .ZN(n675bar);
  OR2_X1 U289 ( .A1(in_10), .A2(in_0), .ZN(n673) );
  AND2_X1 U289bar ( .A1(in_10bar), .A2(in_0bar), .ZN(n673bar);
  OR2_X1 U290 ( .A1(in_59), .A2(in_5), .ZN(n674) );
  AND2_X1 U290bar ( .A1(in_59bar), .A2(in_5bar), .ZN(n674bar);
  OR2_X1 U291 ( .A1(n672), .A2(n671), .ZN(n676) );
  AND2_X1 U291bar ( .A1(n672bar), .A2(n671bar), .ZN(n676bar);
  OR2_X1 U292 ( .A1(in_60), .A2(in_6), .ZN(n671) );
  AND2_X1 U292bar ( .A1(in_60bar), .A2(in_6bar), .ZN(n671bar);
  OR2_X1 U293 ( .A1(in_77), .A2(in_69), .ZN(n672) );
  AND2_X1 U293bar ( .A1(in_77bar), .A2(in_69bar), .ZN(n672bar);
  OR2_X1 U294 ( .A1(in[113]), .A2(n864), .ZN(n700) );
  AND2_X1 U294bar ( .A1(inbar[113]), .A2(n864bar), .ZN(n700bar);
  OR2_X1 U295 ( .A1(n670), .A2(n669), .ZN(n864) );
  AND2_X1 U295bar ( .A1(n670bar), .A2(n669bar), .ZN(n864bar);
  OR2_X1 U296 ( .A1(n668), .A2(n667), .ZN(n669) );
  AND2_X1 U296bar ( .A1(n668bar), .A2(n667bar), .ZN(n669bar);
  OR2_X1 U297 ( .A1(n666), .A2(n665), .ZN(n667) );
  AND2_X1 U297bar ( .A1(n666bar), .A2(n665bar), .ZN(n667bar);
  OR2_X1 U298 ( .A1(in[125]), .A2(in[107]), .ZN(n665) );
  AND2_X1 U298bar ( .A1(inbar[125]), .A2(inbar[107]), .ZN(n665bar);
  OR2_X1 U299 ( .A1(in[138]), .A2(in[126]), .ZN(n666) );
  AND2_X1 U299bar ( .A1(inbar[138]), .A2(inbar[126]), .ZN(n666bar);
  OR2_X1 U300 ( .A1(n664), .A2(n663), .ZN(n668) );
  AND2_X1 U300bar ( .A1(n664bar), .A2(n663bar), .ZN(n668bar);
  OR2_X1 U301 ( .A1(in[189]), .A2(in[143]), .ZN(n663) );
  AND2_X1 U301bar ( .A1(inbar[189]), .A2(inbar[143]), .ZN(n663bar);
  OR2_X1 U302 ( .A1(in[99]), .A2(in[214]), .ZN(n664) );
  AND2_X1 U302bar ( .A1(inbar[99]), .A2(inbar[214]), .ZN(n664bar);
  OR2_X1 U303 ( .A1(n662), .A2(n661), .ZN(n670) );
  AND2_X1 U303bar ( .A1(n662bar), .A2(n661bar), .ZN(n670bar);
  OR2_X1 U304 ( .A1(n660), .A2(n659), .ZN(n661) );
  AND2_X1 U304bar ( .A1(n660bar), .A2(n659bar), .ZN(n661bar);
  OR2_X1 U305 ( .A1(in_15), .A2(in_12), .ZN(n659) );
  AND2_X1 U305bar ( .A1(in_15bar), .A2(in_12bar), .ZN(n659bar);
  OR2_X1 U306 ( .A1(in_20), .A2(in_2), .ZN(n660) );
  AND2_X1 U306bar ( .A1(in_20bar), .A2(in_2bar), .ZN(n660bar);
  OR2_X1 U307 ( .A1(n658), .A2(n657), .ZN(n662) );
  AND2_X1 U307bar ( .A1(n658bar), .A2(n657bar), .ZN(n662bar);
  OR2_X1 U308 ( .A1(in_30), .A2(in_3), .ZN(n657) );
  AND2_X1 U308bar ( .A1(in_30bar), .A2(in_3bar), .ZN(n657bar);
  OR2_X1 U309 ( .A1(in_4), .A2(in_38), .ZN(n658) );
  AND2_X1 U309bar ( .A1(in_4bar), .A2(in_38bar), .ZN(n658bar);
  OR2_X1 U310 ( .A1(n656), .A2(n655), .ZN(n702) );
  AND2_X1 U310bar ( .A1(n656bar), .A2(n655bar), .ZN(n702bar);
  OR2_X1 U311 ( .A1(in[148]), .A2(in[137]), .ZN(n655) );
  AND2_X1 U311bar ( .A1(inbar[148]), .A2(inbar[137]), .ZN(n655bar);
  OR2_X1 U312 ( .A1(in[149]), .A2(n654), .ZN(n656) );
  AND2_X1 U312bar ( .A1(inbar[149]), .A2(n654bar), .ZN(n656bar);
  OR2_X1 U313 ( .A1(in[195]), .A2(in[190]), .ZN(n654) );
  AND2_X1 U313bar ( .A1(inbar[195]), .A2(inbar[190]), .ZN(n654bar);
  OR2_X1 U314 ( .A1(n653), .A2(n652), .ZN(n704) );
  AND2_X1 U314bar ( .A1(n653bar), .A2(n652bar), .ZN(n704bar);
  OR2_X1 U315 ( .A1(n651), .A2(n650), .ZN(n652) );
  AND2_X1 U315bar ( .A1(n651bar), .A2(n650bar), .ZN(n652bar);
  OR2_X1 U316 ( .A1(in[98]), .A2(in[197]), .ZN(n650) );
  AND2_X1 U316bar ( .A1(inbar[98]), .A2(inbar[197]), .ZN(n650bar);
  OR2_X1 U317 ( .A1(in_11), .A2(n649), .ZN(n651) );
  AND2_X1 U317bar ( .A1(in_11bar), .A2(n649bar), .ZN(n651bar);
  OR2_X1 U318 ( .A1(in_26), .A2(in_14), .ZN(n649) );
  AND2_X1 U318bar ( .A1(in_26bar), .A2(in_14bar), .ZN(n649bar);
  OR2_X1 U319 ( .A1(n648), .A2(n647), .ZN(n653) );
  AND2_X1 U319bar ( .A1(n648bar), .A2(n647bar), .ZN(n653bar);
  OR2_X1 U320 ( .A1(in_35), .A2(in_27), .ZN(n647) );
  AND2_X1 U320bar ( .A1(in_35bar), .A2(in_27bar), .ZN(n647bar);
  OR2_X1 U321 ( .A1(in_50), .A2(n646), .ZN(n648) );
  AND2_X1 U321bar ( .A1(in_50bar), .A2(n646bar), .ZN(n648bar);
  OR2_X1 U322 ( .A1(in_78), .A2(in_61), .ZN(n646) );
  AND2_X1 U322bar ( .A1(in_78bar), .A2(in_61bar), .ZN(n646bar);
  OR2_X1 U323 ( .A1(n942), .A2(n645), .ZN(n720) );
  AND2_X1 U323bar ( .A1(n942bar), .A2(n645bar), .ZN(n720bar);
  OR2_X1 U324 ( .A1(in[106]), .A2(n863), .ZN(n645) );
  AND2_X1 U324bar ( .A1(inbar[106]), .A2(n863bar), .ZN(n645bar);
  OR2_X1 U325 ( .A1(n644), .A2(n643), .ZN(n863) );
  AND2_X1 U325bar ( .A1(n644bar), .A2(n643bar), .ZN(n863bar);
  OR2_X1 U326 ( .A1(n642), .A2(n641), .ZN(n643) );
  AND2_X1 U326bar ( .A1(n642bar), .A2(n641bar), .ZN(n643bar);
  OR2_X1 U327 ( .A1(n640), .A2(n639), .ZN(n641) );
  AND2_X1 U327bar ( .A1(n640bar), .A2(n639bar), .ZN(n641bar);
  OR2_X1 U328 ( .A1(in[127]), .A2(in[122]), .ZN(n639) );
  AND2_X1 U328bar ( .A1(inbar[127]), .A2(inbar[122]), .ZN(n639bar);
  OR2_X1 U329 ( .A1(in[156]), .A2(in[132]), .ZN(n640) );
  AND2_X1 U329bar ( .A1(inbar[156]), .A2(inbar[132]), .ZN(n640bar);
  OR2_X1 U330 ( .A1(n638), .A2(n637), .ZN(n642) );
  AND2_X1 U330bar ( .A1(n638bar), .A2(n637bar), .ZN(n642bar);
  OR2_X1 U331 ( .A1(in[159]), .A2(in[157]), .ZN(n637) );
  AND2_X1 U331bar ( .A1(inbar[159]), .A2(inbar[157]), .ZN(n637bar);
  OR2_X1 U332 ( .A1(in[185]), .A2(in[169]), .ZN(n638) );
  AND2_X1 U332bar ( .A1(inbar[185]), .A2(inbar[169]), .ZN(n638bar);
  OR2_X1 U333 ( .A1(n636), .A2(n635), .ZN(n644) );
  AND2_X1 U333bar ( .A1(n636bar), .A2(n635bar), .ZN(n644bar);
  OR2_X1 U334 ( .A1(n634), .A2(n633), .ZN(n635) );
  AND2_X1 U334bar ( .A1(n634bar), .A2(n633bar), .ZN(n635bar);
  OR2_X1 U335 ( .A1(in[239]), .A2(in[218]), .ZN(n633) );
  AND2_X1 U335bar ( .A1(inbar[239]), .A2(inbar[218]), .ZN(n633bar);
  OR2_X1 U336 ( .A1(in_13), .A2(in[87]), .ZN(n634) );
  AND2_X1 U336bar ( .A1(in_13bar), .A2(inbar[87]), .ZN(n634bar);
  OR2_X1 U337 ( .A1(n632), .A2(n631), .ZN(n636) );
  AND2_X1 U337bar ( .A1(n632bar), .A2(n631bar), .ZN(n636bar);
  OR2_X1 U338 ( .A1(in_72), .A2(in_70), .ZN(n631) );
  AND2_X1 U338bar ( .A1(in_72bar), .A2(in_70bar), .ZN(n631bar);
  OR2_X1 U339 ( .A1(in_80), .A2(in_74), .ZN(n632) );
  AND2_X1 U339bar ( .A1(in_80bar), .A2(in_74bar), .ZN(n632bar);
  OR2_X1 U340 ( .A1(n630), .A2(n629), .ZN(n942) );
  AND2_X1 U340bar ( .A1(n630bar), .A2(n629bar), .ZN(n942bar);
  OR2_X1 U341 ( .A1(n628), .A2(n627), .ZN(n629) );
  AND2_X1 U341bar ( .A1(n628bar), .A2(n627bar), .ZN(n629bar);
  OR2_X1 U342 ( .A1(n626), .A2(n625), .ZN(n627) );
  AND2_X1 U342bar ( .A1(n626bar), .A2(n625bar), .ZN(n627bar);
  OR2_X1 U343 ( .A1(in[146]), .A2(in[100]), .ZN(n625) );
  AND2_X1 U343bar ( .A1(inbar[146]), .A2(inbar[100]), .ZN(n625bar);
  OR2_X1 U344 ( .A1(in[168]), .A2(in[152]), .ZN(n626) );
  AND2_X1 U344bar ( .A1(inbar[168]), .A2(inbar[152]), .ZN(n626bar);
  OR2_X1 U345 ( .A1(n624), .A2(n623), .ZN(n628) );
  AND2_X1 U345bar ( .A1(n624bar), .A2(n623bar), .ZN(n628bar);
  OR2_X1 U346 ( .A1(in[199]), .A2(in[182]), .ZN(n623) );
  AND2_X1 U346bar ( .A1(inbar[199]), .A2(inbar[182]), .ZN(n623bar);
  OR2_X1 U347 ( .A1(in[236]), .A2(in[204]), .ZN(n624) );
  AND2_X1 U347bar ( .A1(inbar[236]), .A2(inbar[204]), .ZN(n624bar);
  OR2_X1 U348 ( .A1(n622), .A2(n621), .ZN(n630) );
  AND2_X1 U348bar ( .A1(n622bar), .A2(n621bar), .ZN(n630bar);
  OR2_X1 U349 ( .A1(n620), .A2(n619), .ZN(n621) );
  AND2_X1 U349bar ( .A1(n620bar), .A2(n619bar), .ZN(n621bar);
  OR2_X1 U350 ( .A1(in[89]), .A2(in[246]), .ZN(n619) );
  AND2_X1 U350bar ( .A1(inbar[89]), .A2(inbar[246]), .ZN(n619bar);
  OR2_X1 U351 ( .A1(in[95]), .A2(in[92]), .ZN(n620) );
  AND2_X1 U351bar ( .A1(inbar[95]), .A2(inbar[92]), .ZN(n620bar);
  OR2_X1 U352 ( .A1(n618), .A2(n617), .ZN(n622) );
  AND2_X1 U352bar ( .A1(n618bar), .A2(n617bar), .ZN(n622bar);
  OR2_X1 U353 ( .A1(in_22), .A2(in_16), .ZN(n617) );
  AND2_X1 U353bar ( .A1(in_22bar), .A2(in_16bar), .ZN(n617bar);
  OR2_X1 U354 ( .A1(in_51), .A2(in_49), .ZN(n618) );
  AND2_X1 U354bar ( .A1(in_51bar), .A2(in_49bar), .ZN(n618bar);
  OR2_X1 U355 ( .A1(n616), .A2(n615), .ZN(n722) );
  AND2_X1 U355bar ( .A1(n616bar), .A2(n615bar), .ZN(n722bar);
  OR2_X1 U356 ( .A1(in[158]), .A2(in[115]), .ZN(n615) );
  AND2_X1 U356bar ( .A1(inbar[158]), .A2(inbar[115]), .ZN(n615bar);
  OR2_X1 U357 ( .A1(in[163]), .A2(n614), .ZN(n616) );
  AND2_X1 U357bar ( .A1(inbar[163]), .A2(n614bar), .ZN(n616bar);
  OR2_X1 U358 ( .A1(in[206]), .A2(in[165]), .ZN(n614) );
  AND2_X1 U358bar ( .A1(inbar[206]), .A2(inbar[165]), .ZN(n614bar);
  OR2_X1 U359 ( .A1(n613), .A2(n612), .ZN(n724) );
  AND2_X1 U359bar ( .A1(n613bar), .A2(n612bar), .ZN(n724bar);
  OR2_X1 U360 ( .A1(n611), .A2(n610), .ZN(n612) );
  AND2_X1 U360bar ( .A1(n611bar), .A2(n610bar), .ZN(n612bar);
  OR2_X1 U361 ( .A1(in[213]), .A2(in[207]), .ZN(n610) );
  AND2_X1 U361bar ( .A1(inbar[213]), .A2(inbar[207]), .ZN(n610bar);
  OR2_X1 U362 ( .A1(in[215]), .A2(n609), .ZN(n611) );
  AND2_X1 U362bar ( .A1(inbar[215]), .A2(n609bar), .ZN(n611bar);
  OR2_X1 U363 ( .A1(in[230]), .A2(in[220]), .ZN(n609) );
  AND2_X1 U363bar ( .A1(inbar[230]), .A2(inbar[220]), .ZN(n609bar);
  OR2_X1 U364 ( .A1(n608), .A2(n607), .ZN(n613) );
  AND2_X1 U364bar ( .A1(n608bar), .A2(n607bar), .ZN(n613bar);
  OR2_X1 U365 ( .A1(in[251]), .A2(in[234]), .ZN(n607) );
  AND2_X1 U365bar ( .A1(inbar[251]), .A2(inbar[234]), .ZN(n607bar);
  OR2_X1 U366 ( .A1(in_17), .A2(n606), .ZN(n608) );
  AND2_X1 U366bar ( .A1(in_17bar), .A2(n606bar), .ZN(n608bar);
  OR2_X1 U367 ( .A1(in_65), .A2(in_56), .ZN(n606) );
  AND2_X1 U367bar ( .A1(in_65bar), .A2(in_56bar), .ZN(n606bar);
  OR2_X1 U368 ( .A1(n605), .A2(n604), .ZN(out[0]) );
  AND2_X1 U368bar ( .A1(n605bar), .A2(n604bar), .ZN(outbar[0]);
  OR2_X1 U369 ( .A1(n603), .A2(n602), .ZN(n604) );
  AND2_X1 U369bar ( .A1(n603bar), .A2(n602bar), .ZN(n604bar);
  OR2_X1 U370 ( .A1(n601), .A2(n600), .ZN(n602) );
  AND2_X1 U370bar ( .A1(n601bar), .A2(n600bar), .ZN(n602bar);
  OR2_X1 U371 ( .A1(n820), .A2(n785), .ZN(n600) );
  AND2_X1 U371bar ( .A1(n820bar), .A2(n785bar), .ZN(n600bar);
  OR2_X1 U372 ( .A1(n599), .A2(n598), .ZN(n785) );
  AND2_X1 U372bar ( .A1(n599bar), .A2(n598bar), .ZN(n785bar);
  OR2_X1 U373 ( .A1(n597), .A2(n596), .ZN(n598) );
  AND2_X1 U373bar ( .A1(n597bar), .A2(n596bar), .ZN(n598bar);
  OR2_X1 U374 ( .A1(n595), .A2(n594), .ZN(n596) );
  AND2_X1 U374bar ( .A1(n595bar), .A2(n594bar), .ZN(n596bar);
  OR2_X1 U375 ( .A1(in[135]), .A2(in[104]), .ZN(n594) );
  AND2_X1 U375bar ( .A1(inbar[135]), .A2(inbar[104]), .ZN(n594bar);
  OR2_X1 U376 ( .A1(in[188]), .A2(in[178]), .ZN(n595) );
  AND2_X1 U376bar ( .A1(inbar[188]), .A2(inbar[178]), .ZN(n595bar);
  OR2_X1 U377 ( .A1(n593), .A2(n592), .ZN(n597) );
  AND2_X1 U377bar ( .A1(n593bar), .A2(n592bar), .ZN(n597bar);
  OR2_X1 U378 ( .A1(in[217]), .A2(in[194]), .ZN(n592) );
  AND2_X1 U378bar ( .A1(inbar[217]), .A2(inbar[194]), .ZN(n592bar);
  OR2_X1 U379 ( .A1(in[237]), .A2(in[218]), .ZN(n593) );
  AND2_X1 U379bar ( .A1(inbar[237]), .A2(inbar[218]), .ZN(n593bar);
  OR2_X1 U380 ( .A1(n591), .A2(n590), .ZN(n599) );
  AND2_X1 U380bar ( .A1(n591bar), .A2(n590bar), .ZN(n599bar);
  OR2_X1 U381 ( .A1(n589), .A2(n588), .ZN(n590) );
  AND2_X1 U381bar ( .A1(n589bar), .A2(n588bar), .ZN(n590bar);
  OR2_X1 U382 ( .A1(in_2), .A2(in_10), .ZN(n588) );
  AND2_X1 U382bar ( .A1(in_2bar), .A2(in_10bar), .ZN(n588bar);
  OR2_X1 U383 ( .A1(in_47), .A2(in_22), .ZN(n589) );
  AND2_X1 U383bar ( .A1(in_47bar), .A2(in_22bar), .ZN(n589bar);
  OR2_X1 U384 ( .A1(n587), .A2(n586), .ZN(n591) );
  AND2_X1 U384bar ( .A1(n587bar), .A2(n586bar), .ZN(n591bar);
  OR2_X1 U385 ( .A1(in_56), .A2(in_54), .ZN(n586) );
  AND2_X1 U385bar ( .A1(in_56bar), .A2(in_54bar), .ZN(n586bar);
  OR2_X1 U386 ( .A1(in_63), .A2(in_61), .ZN(n587) );
  AND2_X1 U386bar ( .A1(in_63bar), .A2(in_61bar), .ZN(n587bar);
  OR2_X1 U387 ( .A1(n585), .A2(n584), .ZN(n820) );
  AND2_X1 U387bar ( .A1(n585bar), .A2(n584bar), .ZN(n820bar);
  OR2_X1 U388 ( .A1(n583), .A2(n582), .ZN(n584) );
  AND2_X1 U388bar ( .A1(n583bar), .A2(n582bar), .ZN(n584bar);
  OR2_X1 U389 ( .A1(n581), .A2(n580), .ZN(n582) );
  AND2_X1 U389bar ( .A1(n581bar), .A2(n580bar), .ZN(n582bar);
  OR2_X1 U390 ( .A1(in[158]), .A2(in[142]), .ZN(n580) );
  AND2_X1 U390bar ( .A1(inbar[158]), .A2(inbar[142]), .ZN(n580bar);
  OR2_X1 U391 ( .A1(in[175]), .A2(in[164]), .ZN(n581) );
  AND2_X1 U391bar ( .A1(inbar[175]), .A2(inbar[164]), .ZN(n581bar);
  OR2_X1 U392 ( .A1(n579), .A2(n578), .ZN(n583) );
  AND2_X1 U392bar ( .A1(n579bar), .A2(n578bar), .ZN(n583bar);
  OR2_X1 U393 ( .A1(in[228]), .A2(in[204]), .ZN(n578) );
  AND2_X1 U393bar ( .A1(inbar[228]), .A2(inbar[204]), .ZN(n578bar);
  OR2_X1 U394 ( .A1(in[91]), .A2(in[87]), .ZN(n579) );
  AND2_X1 U394bar ( .A1(inbar[91]), .A2(inbar[87]), .ZN(n579bar);
  OR2_X1 U395 ( .A1(n577), .A2(n576), .ZN(n585) );
  AND2_X1 U395bar ( .A1(n577bar), .A2(n576bar), .ZN(n585bar);
  OR2_X1 U396 ( .A1(n575), .A2(n574), .ZN(n576) );
  AND2_X1 U396bar ( .A1(n575bar), .A2(n574bar), .ZN(n576bar);
  OR2_X1 U397 ( .A1(in_21), .A2(in_11), .ZN(n574) );
  AND2_X1 U397bar ( .A1(in_21bar), .A2(in_11bar), .ZN(n574bar);
  OR2_X1 U398 ( .A1(in_5), .A2(in_3), .ZN(n575) );
  AND2_X1 U398bar ( .A1(in_5bar), .A2(in_3bar), .ZN(n575bar);
  OR2_X1 U399 ( .A1(n573), .A2(n572), .ZN(n577) );
  AND2_X1 U399bar ( .A1(n573bar), .A2(n572bar), .ZN(n577bar);
  OR2_X1 U400 ( .A1(in_68), .A2(in_64), .ZN(n572) );
  AND2_X1 U400bar ( .A1(in_68bar), .A2(in_64bar), .ZN(n572bar);
  OR2_X1 U401 ( .A1(in_76), .A2(in_73), .ZN(n573) );
  AND2_X1 U401bar ( .A1(in_76bar), .A2(in_73bar), .ZN(n573bar);
  OR2_X1 U402 ( .A1(n778), .A2(n571), .ZN(n601) );
  AND2_X1 U402bar ( .A1(n778bar), .A2(n571bar), .ZN(n601bar);
  OR2_X1 U403 ( .A1(in[100]), .A2(n965), .ZN(n571) );
  AND2_X1 U403bar ( .A1(inbar[100]), .A2(n965bar), .ZN(n571bar);
  OR2_X1 U404 ( .A1(n570), .A2(n569), .ZN(n965) );
  AND2_X1 U404bar ( .A1(n570bar), .A2(n569bar), .ZN(n965bar);
  OR2_X1 U405 ( .A1(n568), .A2(n567), .ZN(n569) );
  AND2_X1 U405bar ( .A1(n568bar), .A2(n567bar), .ZN(n569bar);
  OR2_X1 U406 ( .A1(n566), .A2(n565), .ZN(n567) );
  AND2_X1 U406bar ( .A1(n566bar), .A2(n565bar), .ZN(n567bar);
  OR2_X1 U407 ( .A1(n817), .A2(n750), .ZN(n565) );
  AND2_X1 U407bar ( .A1(n817bar), .A2(n750bar), .ZN(n565bar);
  OR2_X1 U408 ( .A1(n564), .A2(n563), .ZN(n750) );
  AND2_X1 U408bar ( .A1(n564bar), .A2(n563bar), .ZN(n750bar);
  OR2_X1 U409 ( .A1(n562), .A2(n561), .ZN(n563) );
  AND2_X1 U409bar ( .A1(n562bar), .A2(n561bar), .ZN(n563bar);
  OR2_X1 U410 ( .A1(n560), .A2(n559), .ZN(n561) );
  AND2_X1 U410bar ( .A1(n560bar), .A2(n559bar), .ZN(n561bar);
  OR2_X1 U411 ( .A1(in[119]), .A2(in[103]), .ZN(n559) );
  AND2_X1 U411bar ( .A1(inbar[119]), .A2(inbar[103]), .ZN(n559bar);
  OR2_X1 U412 ( .A1(in[137]), .A2(in[133]), .ZN(n560) );
  AND2_X1 U412bar ( .A1(inbar[137]), .A2(inbar[133]), .ZN(n560bar);
  OR2_X1 U413 ( .A1(n558), .A2(n557), .ZN(n562) );
  AND2_X1 U413bar ( .A1(n558bar), .A2(n557bar), .ZN(n562bar);
  OR2_X1 U414 ( .A1(in[176]), .A2(in[173]), .ZN(n557) );
  AND2_X1 U414bar ( .A1(inbar[176]), .A2(inbar[173]), .ZN(n557bar);
  OR2_X1 U415 ( .A1(in[210]), .A2(in[181]), .ZN(n558) );
  AND2_X1 U415bar ( .A1(inbar[210]), .A2(inbar[181]), .ZN(n558bar);
  OR2_X1 U416 ( .A1(n556), .A2(n555), .ZN(n564) );
  AND2_X1 U416bar ( .A1(n556bar), .A2(n555bar), .ZN(n564bar);
  OR2_X1 U417 ( .A1(n554), .A2(n553), .ZN(n555) );
  AND2_X1 U417bar ( .A1(n554bar), .A2(n553bar), .ZN(n555bar);
  OR2_X1 U418 ( .A1(in_13), .A2(in[234]), .ZN(n553) );
  AND2_X1 U418bar ( .A1(in_13bar), .A2(inbar[234]), .ZN(n553bar);
  OR2_X1 U419 ( .A1(in_38), .A2(in_32), .ZN(n554) );
  AND2_X1 U419bar ( .A1(in_38bar), .A2(in_32bar), .ZN(n554bar);
  OR2_X1 U420 ( .A1(n552), .A2(n551), .ZN(n556) );
  AND2_X1 U420bar ( .A1(n552bar), .A2(n551bar), .ZN(n556bar);
  OR2_X1 U421 ( .A1(in_42), .A2(in_41), .ZN(n551) );
  AND2_X1 U421bar ( .A1(in_42bar), .A2(in_41bar), .ZN(n551bar);
  OR2_X1 U422 ( .A1(in_7), .A2(in_49), .ZN(n552) );
  AND2_X1 U422bar ( .A1(in_7bar), .A2(in_49bar), .ZN(n552bar);
  OR2_X1 U423 ( .A1(n550), .A2(n549), .ZN(n817) );
  AND2_X1 U423bar ( .A1(n550bar), .A2(n549bar), .ZN(n817bar);
  OR2_X1 U424 ( .A1(n548), .A2(n547), .ZN(n549) );
  AND2_X1 U424bar ( .A1(n548bar), .A2(n547bar), .ZN(n549bar);
  OR2_X1 U425 ( .A1(n546), .A2(n545), .ZN(n547) );
  AND2_X1 U425bar ( .A1(n546bar), .A2(n545bar), .ZN(n547bar);
  OR2_X1 U426 ( .A1(in[159]), .A2(in[105]), .ZN(n545) );
  AND2_X1 U426bar ( .A1(inbar[159]), .A2(inbar[105]), .ZN(n545bar);
  OR2_X1 U427 ( .A1(in[206]), .A2(in[183]), .ZN(n546) );
  AND2_X1 U427bar ( .A1(inbar[206]), .A2(inbar[183]), .ZN(n546bar);
  OR2_X1 U428 ( .A1(n544), .A2(n543), .ZN(n548) );
  AND2_X1 U428bar ( .A1(n544bar), .A2(n543bar), .ZN(n548bar);
  OR2_X1 U429 ( .A1(in[229]), .A2(in[219]), .ZN(n543) );
  AND2_X1 U429bar ( .A1(inbar[229]), .A2(inbar[219]), .ZN(n543bar);
  OR2_X1 U430 ( .A1(in[235]), .A2(in[232]), .ZN(n544) );
  AND2_X1 U430bar ( .A1(inbar[235]), .A2(inbar[232]), .ZN(n544bar);
  OR2_X1 U431 ( .A1(n542), .A2(n541), .ZN(n550) );
  AND2_X1 U431bar ( .A1(n542bar), .A2(n541bar), .ZN(n550bar);
  OR2_X1 U432 ( .A1(n540), .A2(n539), .ZN(n541) );
  AND2_X1 U432bar ( .A1(n540bar), .A2(n539bar), .ZN(n541bar);
  OR2_X1 U433 ( .A1(in[249]), .A2(in[242]), .ZN(n539) );
  AND2_X1 U433bar ( .A1(inbar[249]), .A2(inbar[242]), .ZN(n539bar);
  OR2_X1 U434 ( .A1(in[89]), .A2(in[254]), .ZN(n540) );
  AND2_X1 U434bar ( .A1(inbar[89]), .A2(inbar[254]), .ZN(n540bar);
  OR2_X1 U435 ( .A1(n538), .A2(n537), .ZN(n542) );
  AND2_X1 U435bar ( .A1(n538bar), .A2(n537bar), .ZN(n542bar);
  OR2_X1 U436 ( .A1(in_14), .A2(in[99]), .ZN(n537) );
  AND2_X1 U436bar ( .A1(in_14bar), .A2(inbar[99]), .ZN(n537bar);
  OR2_X1 U437 ( .A1(in_60), .A2(in_18), .ZN(n538) );
  AND2_X1 U437bar ( .A1(in_60bar), .A2(in_18bar), .ZN(n538bar);
  OR2_X1 U438 ( .A1(in[113]), .A2(n763), .ZN(n566) );
  AND2_X1 U438bar ( .A1(inbar[113]), .A2(n763bar), .ZN(n566bar);
  OR2_X1 U439 ( .A1(n536), .A2(n535), .ZN(n763) );
  AND2_X1 U439bar ( .A1(n536bar), .A2(n535bar), .ZN(n763bar);
  OR2_X1 U440 ( .A1(n534), .A2(n533), .ZN(n535) );
  AND2_X1 U440bar ( .A1(n534bar), .A2(n533bar), .ZN(n535bar);
  OR2_X1 U441 ( .A1(n532), .A2(n531), .ZN(n533) );
  AND2_X1 U441bar ( .A1(n532bar), .A2(n531bar), .ZN(n533bar);
  OR2_X1 U442 ( .A1(in[115]), .A2(in[110]), .ZN(n531) );
  AND2_X1 U442bar ( .A1(inbar[115]), .A2(inbar[110]), .ZN(n531bar);
  OR2_X1 U443 ( .A1(in[125]), .A2(in[117]), .ZN(n532) );
  AND2_X1 U443bar ( .A1(inbar[125]), .A2(inbar[117]), .ZN(n532bar);
  OR2_X1 U444 ( .A1(n530), .A2(n529), .ZN(n534) );
  AND2_X1 U444bar ( .A1(n530bar), .A2(n529bar), .ZN(n534bar);
  OR2_X1 U445 ( .A1(in[180]), .A2(in[128]), .ZN(n529) );
  AND2_X1 U445bar ( .A1(inbar[180]), .A2(inbar[128]), .ZN(n529bar);
  OR2_X1 U446 ( .A1(in[205]), .A2(in[201]), .ZN(n530) );
  AND2_X1 U446bar ( .A1(inbar[205]), .A2(inbar[201]), .ZN(n530bar);
  OR2_X1 U447 ( .A1(n528), .A2(n527), .ZN(n536) );
  AND2_X1 U447bar ( .A1(n528bar), .A2(n527bar), .ZN(n536bar);
  OR2_X1 U448 ( .A1(n526), .A2(n525), .ZN(n527) );
  AND2_X1 U448bar ( .A1(n526bar), .A2(n525bar), .ZN(n527bar);
  OR2_X1 U449 ( .A1(in[244]), .A2(in[239]), .ZN(n525) );
  AND2_X1 U449bar ( .A1(inbar[244]), .A2(inbar[239]), .ZN(n525bar);
  OR2_X1 U450 ( .A1(in[95]), .A2(in[83]), .ZN(n526) );
  AND2_X1 U450bar ( .A1(inbar[95]), .A2(inbar[83]), .ZN(n526bar);
  OR2_X1 U451 ( .A1(n524), .A2(n523), .ZN(n528) );
  AND2_X1 U451bar ( .A1(n524bar), .A2(n523bar), .ZN(n528bar);
  OR2_X1 U452 ( .A1(in_24), .A2(in[97]), .ZN(n523) );
  AND2_X1 U452bar ( .A1(in_24bar), .A2(inbar[97]), .ZN(n523bar);
  OR2_X1 U453 ( .A1(in_33), .A2(in_27), .ZN(n524) );
  AND2_X1 U453bar ( .A1(in_33bar), .A2(in_27bar), .ZN(n524bar);
  OR2_X1 U454 ( .A1(n522), .A2(n521), .ZN(n568) );
  AND2_X1 U454bar ( .A1(n522bar), .A2(n521bar), .ZN(n568bar);
  OR2_X1 U455 ( .A1(in[145]), .A2(in[126]), .ZN(n521) );
  AND2_X1 U455bar ( .A1(inbar[145]), .A2(inbar[126]), .ZN(n521bar);
  OR2_X1 U456 ( .A1(in[169]), .A2(n520), .ZN(n522) );
  AND2_X1 U456bar ( .A1(inbar[169]), .A2(n520bar), .ZN(n522bar);
  OR2_X1 U457 ( .A1(in[221]), .A2(in[172]), .ZN(n520) );
  AND2_X1 U457bar ( .A1(inbar[221]), .A2(inbar[172]), .ZN(n520bar);
  OR2_X1 U458 ( .A1(n519), .A2(n518), .ZN(n570) );
  AND2_X1 U458bar ( .A1(n519bar), .A2(n518bar), .ZN(n570bar);
  OR2_X1 U459 ( .A1(n517), .A2(n516), .ZN(n518) );
  AND2_X1 U459bar ( .A1(n517bar), .A2(n516bar), .ZN(n518bar);
  OR2_X1 U460 ( .A1(in[241]), .A2(in[224]), .ZN(n516) );
  AND2_X1 U460bar ( .A1(inbar[241]), .A2(inbar[224]), .ZN(n516bar);
  OR2_X1 U461 ( .A1(in[86]), .A2(n515), .ZN(n517) );
  AND2_X1 U461bar ( .A1(inbar[86]), .A2(n515bar), .ZN(n517bar);
  OR2_X1 U462 ( .A1(in_43), .A2(in_34), .ZN(n515) );
  AND2_X1 U462bar ( .A1(in_43bar), .A2(in_34bar), .ZN(n515bar);
  OR2_X1 U463 ( .A1(n514), .A2(n513), .ZN(n519) );
  AND2_X1 U463bar ( .A1(n514bar), .A2(n513bar), .ZN(n519bar);
  OR2_X1 U464 ( .A1(in_65), .A2(in_51), .ZN(n513) );
  AND2_X1 U464bar ( .A1(in_65bar), .A2(in_51bar), .ZN(n513bar);
  OR2_X1 U465 ( .A1(in_75), .A2(n512), .ZN(n514) );
  AND2_X1 U465bar ( .A1(in_75bar), .A2(n512bar), .ZN(n514bar);
  OR2_X1 U466 ( .A1(in_81), .A2(in_77), .ZN(n512) );
  AND2_X1 U466bar ( .A1(in_81bar), .A2(in_77bar), .ZN(n512bar);
  OR2_X1 U467 ( .A1(n511), .A2(n510), .ZN(n778) );
  AND2_X1 U467bar ( .A1(n511bar), .A2(n510bar), .ZN(n778bar);
  OR2_X1 U468 ( .A1(n509), .A2(n508), .ZN(n510) );
  AND2_X1 U468bar ( .A1(n509bar), .A2(n508bar), .ZN(n510bar);
  OR2_X1 U469 ( .A1(n507), .A2(n506), .ZN(n508) );
  AND2_X1 U469bar ( .A1(n507bar), .A2(n506bar), .ZN(n508bar);
  OR2_X1 U470 ( .A1(in[107]), .A2(in[101]), .ZN(n506) );
  AND2_X1 U470bar ( .A1(inbar[107]), .A2(inbar[101]), .ZN(n506bar);
  OR2_X1 U471 ( .A1(in[139]), .A2(in[132]), .ZN(n507) );
  AND2_X1 U471bar ( .A1(inbar[139]), .A2(inbar[132]), .ZN(n507bar);
  OR2_X1 U472 ( .A1(n505), .A2(n504), .ZN(n509) );
  AND2_X1 U472bar ( .A1(n505bar), .A2(n504bar), .ZN(n509bar);
  OR2_X1 U473 ( .A1(in[146]), .A2(in[141]), .ZN(n504) );
  AND2_X1 U473bar ( .A1(inbar[146]), .A2(inbar[141]), .ZN(n504bar);
  OR2_X1 U474 ( .A1(in[203]), .A2(in[179]), .ZN(n505) );
  AND2_X1 U474bar ( .A1(inbar[203]), .A2(inbar[179]), .ZN(n505bar);
  OR2_X1 U475 ( .A1(n503), .A2(n502), .ZN(n511) );
  AND2_X1 U475bar ( .A1(n503bar), .A2(n502bar), .ZN(n511bar);
  OR2_X1 U476 ( .A1(n501), .A2(n500), .ZN(n502) );
  AND2_X1 U476bar ( .A1(n501bar), .A2(n500bar), .ZN(n502bar);
  OR2_X1 U477 ( .A1(in[243]), .A2(in[222]), .ZN(n500) );
  AND2_X1 U477bar ( .A1(inbar[243]), .A2(inbar[222]), .ZN(n500bar);
  OR2_X1 U478 ( .A1(in[251]), .A2(in[250]), .ZN(n501) );
  AND2_X1 U478bar ( .A1(inbar[251]), .A2(inbar[250]), .ZN(n501bar);
  OR2_X1 U479 ( .A1(n499), .A2(n498), .ZN(n503) );
  AND2_X1 U479bar ( .A1(n499bar), .A2(n498bar), .ZN(n503bar);
  OR2_X1 U480 ( .A1(in_37), .A2(in_19), .ZN(n498) );
  AND2_X1 U480bar ( .A1(in_37bar), .A2(in_19bar), .ZN(n498bar);
  OR2_X1 U481 ( .A1(in_78), .A2(in_6), .ZN(n499) );
  AND2_X1 U481bar ( .A1(in_78bar), .A2(in_6bar), .ZN(n499bar);
  OR2_X1 U482 ( .A1(n497), .A2(n496), .ZN(n603) );
  AND2_X1 U482bar ( .A1(n497bar), .A2(n496bar), .ZN(n603bar);
  OR2_X1 U483 ( .A1(in[112]), .A2(in[102]), .ZN(n496) );
  AND2_X1 U483bar ( .A1(inbar[112]), .A2(inbar[102]), .ZN(n496bar);
  OR2_X1 U484 ( .A1(in[123]), .A2(n495), .ZN(n497) );
  AND2_X1 U484bar ( .A1(inbar[123]), .A2(n495bar), .ZN(n497bar);
  OR2_X1 U485 ( .A1(in[143]), .A2(in[130]), .ZN(n495) );
  AND2_X1 U485bar ( .A1(inbar[143]), .A2(inbar[130]), .ZN(n495bar);
  OR2_X1 U486 ( .A1(n494), .A2(n493), .ZN(n605) );
  AND2_X1 U486bar ( .A1(n494bar), .A2(n493bar), .ZN(n605bar);
  OR2_X1 U487 ( .A1(n492), .A2(n491), .ZN(n493) );
  AND2_X1 U487bar ( .A1(n492bar), .A2(n491bar), .ZN(n493bar);
  OR2_X1 U488 ( .A1(in[216]), .A2(in[213]), .ZN(n491) );
  AND2_X1 U488bar ( .A1(inbar[216]), .A2(inbar[213]), .ZN(n491bar);
  OR2_X1 U489 ( .A1(in[227]), .A2(n490), .ZN(n492) );
  AND2_X1 U489bar ( .A1(inbar[227]), .A2(n490bar), .ZN(n492bar);
  OR2_X1 U490 ( .A1(in_0), .A2(in[248]), .ZN(n490) );
  AND2_X1 U490bar ( .A1(in_0bar), .A2(inbar[248]), .ZN(n490bar);
  OR2_X1 U491 ( .A1(n489), .A2(n488), .ZN(n494) );
  AND2_X1 U491bar ( .A1(n489bar), .A2(n488bar), .ZN(n494bar);
  OR2_X1 U492 ( .A1(in_46), .A2(in_44), .ZN(n488) );
  AND2_X1 U492bar ( .A1(in_46bar), .A2(in_44bar), .ZN(n488bar);
  OR2_X1 U493 ( .A1(in_50), .A2(n487), .ZN(n489) );
  AND2_X1 U493bar ( .A1(in_50bar), .A2(n487bar), .ZN(n489bar);
  OR2_X1 U494 ( .A1(in_9), .A2(in_80), .ZN(n487) );
  AND2_X1 U494bar ( .A1(in_9bar), .A2(in_80bar), .ZN(n487bar);
endmodule




module sBox_19 ( in, out );
  input [7:0] in;
  //input_done

  output [7:0] out;
  //output_done

  wire   [255:0] decodeOut;
  //wire_done

  decode_19 dec ( .in(in), .out(decodeOut) );
  encode_19 enc ( .in(decodeOut), .out(out) );
endmodule


module scale2_1 ( in, out );
  input [7:0] in;
  //input_done

  output [7:0] out;
  //output_done

  wire   in_0, \in[6] , \in[5] , \in[4] , \in[1] , \in[7] , n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20;
  //wire_done

  assign in_0 = in[0];
  assign out[7] = \in[6] ;
  assign \in[6]  = in[6];
  assign out[6] = \in[5] ;
  assign \in[5]  = in[5];
  assign out[5] = \in[4] ;
  assign \in[4]  = in[4];
  assign out[2] = \in[1] ;
  assign \in[1]  = in[1];
  assign out[0] = \in[7] ;
  assign \in[7]  = in[7];

  INV_X1 U1 ( .A(\in[7]), .ZN(n20) );
  INV_X1 U2 ( .A(in[3]), .ZN(n19) );
  INV_X1 U3 ( .A(in[2]), .ZN(n18) );
  INV_X1 U4 ( .A(in_0), .ZN(n17) );
  OR2_X1 U5 ( .A1(n16), .A2(n15), .ZN(out[4]) );
  AND2_X1 U6 ( .A1(in[3]), .A2(n20), .ZN(n15) );
  AND2_X1 U7 ( .A1(\in[7]), .A2(n19), .ZN(n16) );
  OR2_X1 U8 ( .A1(n14), .A2(n13), .ZN(out[3]) );
  AND2_X1 U9 ( .A1(in[2]), .A2(n20), .ZN(n13) );
  AND2_X1 U10 ( .A1(\in[7]), .A2(n18), .ZN(n14) );
  OR2_X1 U11 ( .A1(n12), .A2(n11), .ZN(out[1]) );
  AND2_X1 U12 ( .A1(in_0), .A2(n20), .ZN(n11) );
  AND2_X1 U13 ( .A1(\in[7]), .A2(n17), .ZN(n12) );
endmodule


module scale2_2 ( in, out );
  input [7:0] in;
  //input_done

  output [7:0] out;
  //output_done

  wire   in_0, \in[6] , \in[5] , \in[4] , \in[1] , \in[7] , n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20;
  //wire_done

  assign in_0 = in[0];
  assign out[7] = \in[6] ;
  assign \in[6]  = in[6];
  assign out[6] = \in[5] ;
  assign \in[5]  = in[5];
  assign out[5] = \in[4] ;
  assign \in[4]  = in[4];
  assign out[2] = \in[1] ;
  assign \in[1]  = in[1];
  assign out[0] = \in[7] ;
  assign \in[7]  = in[7];

  INV_X1 U1 ( .A(\in[7]), .ZN(n20) );
  INV_X1 U2 ( .A(in[3]), .ZN(n19) );
  INV_X1 U3 ( .A(in[2]), .ZN(n18) );
  INV_X1 U4 ( .A(in_0), .ZN(n17) );
  OR2_X1 U5 ( .A1(n16), .A2(n15), .ZN(out[4]) );
  AND2_X1 U6 ( .A1(in[3]), .A2(n20), .ZN(n15) );
  AND2_X1 U7 ( .A1(\in[7]), .A2(n19), .ZN(n16) );
  OR2_X1 U8 ( .A1(n14), .A2(n13), .ZN(out[3]) );
  AND2_X1 U9 ( .A1(in[2]), .A2(n20), .ZN(n13) );
  AND2_X1 U10 ( .A1(\in[7]), .A2(n18), .ZN(n14) );
  OR2_X1 U11 ( .A1(n12), .A2(n11), .ZN(out[1]) );
  AND2_X1 U12 ( .A1(in_0), .A2(n20), .ZN(n11) );
  AND2_X1 U13 ( .A1(\in[7]), .A2(n17), .ZN(n12) );
endmodule


module scale2_3 ( in, out );
  input [7:0] in;
  //input_done

  output [7:0] out;
  //output_done

  wire   in_0, \in[6] , \in[5] , \in[4] , \in[1] , \in[7] , n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20;
  //wire_done
  assign in_0 = in[0];
  assign out[7] = \in[6] ;
  assign \in[6]  = in[6];
  assign out[6] = \in[5] ;
  assign \in[5]  = in[5];
  assign out[5] = \in[4] ;
  assign \in[4]  = in[4];
  assign out[2] = \in[1] ;
  assign \in[1]  = in[1];
  assign out[0] = \in[7] ;
  assign \in[7]  = in[7];

  INV_X1 U1 ( .A(\in[7]), .ZN(n20) );
  INV_X1 U2 ( .A(in[3]), .ZN(n19) );
  INV_X1 U3 ( .A(in[2]), .ZN(n18) );
  INV_X1 U4 ( .A(in_0), .ZN(n17) );
  OR2_X1 U5 ( .A1(n16), .A2(n15), .ZN(out[4]) );
  AND2_X1 U6 ( .A1(in[3]), .A2(n20), .ZN(n15) );
  AND2_X1 U7 ( .A1(\in[7]), .A2(n19), .ZN(n16) );
  OR2_X1 U8 ( .A1(n14), .A2(n13), .ZN(out[3]) );
  AND2_X1 U9 ( .A1(in[2]), .A2(n20), .ZN(n13) );
  AND2_X1 U10 ( .A1(\in[7]), .A2(n18), .ZN(n14) );
  OR2_X1 U11 ( .A1(n12), .A2(n11), .ZN(out[1]) );
  AND2_X1 U12 ( .A1(in_0), .A2(n20), .ZN(n11) );
  AND2_X1 U13 ( .A1(\in[7]), .A2(n17), .ZN(n12) );
endmodule


module scale2_4 ( in, out );
  input [7:0] in;
  //input_done

  output [7:0] out;
  //output_done

  wire   in_0, \in[6] , \in[5] , \in[4] , \in[1] , \in[7] , n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20;
  //wire_done
  assign in_0 = in[0];
  assign out[7] = \in[6] ;
  assign \in[6]  = in[6];
  assign out[6] = \in[5] ;
  assign \in[5]  = in[5];
  assign out[5] = \in[4] ;
  assign \in[4]  = in[4];
  assign out[2] = \in[1] ;
  assign \in[1]  = in[1];
  assign out[0] = \in[7] ;
  assign \in[7]  = in[7];

  INV_X1 U1 ( .A(\in[7]), .ZN(n20) );
  INV_X1 U2 ( .A(in[3]), .ZN(n19) );
  INV_X1 U3 ( .A(in[2]), .ZN(n18) );
  INV_X1 U4 ( .A(in_0), .ZN(n17) );
  OR2_X1 U5 ( .A1(n16), .A2(n15), .ZN(out[4]) );
  AND2_X1 U6 ( .A1(in[3]), .A2(n20), .ZN(n15) );
  AND2_X1 U7 ( .A1(\in[7]), .A2(n19), .ZN(n16) );
  OR2_X1 U8 ( .A1(n14), .A2(n13), .ZN(out[3]) );
  AND2_X1 U9 ( .A1(in[2]), .A2(n20), .ZN(n13) );
  AND2_X1 U10 ( .A1(\in[7]), .A2(n18), .ZN(n14) );
  OR2_X1 U11 ( .A1(n12), .A2(n11), .ZN(out[1]) );
  AND2_X1 U12 ( .A1(in_0), .A2(n20), .ZN(n11) );
  AND2_X1 U13 ( .A1(\in[7]), .A2(n17), .ZN(n12) );
endmodule


module byteXor_2 ( a, b, y );
  input [7:0] a;
  input [7:0] b;
  //input_done

  output [7:0] y;
  //output_done

  wire   n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64;
  //wire_done

  INV_X1 U1 ( .A(n47), .ZN(n64) );
  INV_X1 U2 ( .A(a[7]), .ZN(n63) );
  INV_X1 U3 ( .A(n45), .ZN(n62) );
  INV_X1 U4 ( .A(a[6]), .ZN(n61) );
  INV_X1 U5 ( .A(n43), .ZN(n60) );
  INV_X1 U6 ( .A(a[5]), .ZN(n59) );
  INV_X1 U7 ( .A(n41), .ZN(n58) );
  INV_X1 U8 ( .A(a[4]), .ZN(n57) );
  INV_X1 U9 ( .A(n39), .ZN(n56) );
  INV_X1 U10 ( .A(a[3]), .ZN(n55) );
  INV_X1 U11 ( .A(n37), .ZN(n54) );
  INV_X1 U12 ( .A(a[2]), .ZN(n53) );
  INV_X1 U13 ( .A(n35), .ZN(n52) );
  INV_X1 U14 ( .A(a[1]), .ZN(n51) );
  INV_X1 U15 ( .A(n33), .ZN(n50) );
  INV_X1 U16 ( .A(a[0]), .ZN(n49) );
  OR2_X1 U17 ( .A1(n48), .A2(n64), .ZN(y[7]) );
  OR2_X1 U18 ( .A1(n63), .A2(b[7]), .ZN(n47) );
  AND2_X1 U19 ( .A1(b[7]), .A2(n63), .ZN(n48) );
  OR2_X1 U20 ( .A1(n46), .A2(n62), .ZN(y[6]) );
  OR2_X1 U21 ( .A1(n61), .A2(b[6]), .ZN(n45) );
  AND2_X1 U22 ( .A1(b[6]), .A2(n61), .ZN(n46) );
  OR2_X1 U23 ( .A1(n44), .A2(n60), .ZN(y[5]) );
  OR2_X1 U24 ( .A1(n59), .A2(b[5]), .ZN(n43) );
  AND2_X1 U25 ( .A1(b[5]), .A2(n59), .ZN(n44) );
  OR2_X1 U26 ( .A1(n42), .A2(n58), .ZN(y[4]) );
  OR2_X1 U27 ( .A1(n57), .A2(b[4]), .ZN(n41) );
  AND2_X1 U28 ( .A1(b[4]), .A2(n57), .ZN(n42) );
  OR2_X1 U29 ( .A1(n40), .A2(n56), .ZN(y[3]) );
  OR2_X1 U30 ( .A1(n55), .A2(b[3]), .ZN(n39) );
  AND2_X1 U31 ( .A1(b[3]), .A2(n55), .ZN(n40) );
  OR2_X1 U32 ( .A1(n38), .A2(n54), .ZN(y[2]) );
  OR2_X1 U33 ( .A1(n53), .A2(b[2]), .ZN(n37) );
  AND2_X1 U34 ( .A1(b[2]), .A2(n53), .ZN(n38) );
  OR2_X1 U35 ( .A1(n36), .A2(n52), .ZN(y[1]) );
  OR2_X1 U36 ( .A1(n51), .A2(b[1]), .ZN(n35) );
  AND2_X1 U37 ( .A1(b[1]), .A2(n51), .ZN(n36) );
  OR2_X1 U38 ( .A1(n34), .A2(n50), .ZN(y[0]) );
  OR2_X1 U39 ( .A1(n49), .A2(b[0]), .ZN(n33) );
  AND2_X1 U40 ( .A1(b[0]), .A2(n49), .ZN(n34) );
endmodule


module byteXor_3 ( a, b, y );
  input [7:0] a;
  input [7:0] b;
  //input_done

  output [7:0] y;
  //output_done

  wire   n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64;
  //wire_done

  INV_X1 U1 ( .A(n47), .ZN(n64) );
  INV_X1 U2 ( .A(a[7]), .ZN(n63) );
  INV_X1 U3 ( .A(n45), .ZN(n62) );
  INV_X1 U4 ( .A(a[6]), .ZN(n61) );
  INV_X1 U5 ( .A(n43), .ZN(n60) );
  INV_X1 U6 ( .A(a[5]), .ZN(n59) );
  INV_X1 U7 ( .A(n41), .ZN(n58) );
  INV_X1 U8 ( .A(a[4]), .ZN(n57) );
  INV_X1 U9 ( .A(n39), .ZN(n56) );
  INV_X1 U10 ( .A(a[3]), .ZN(n55) );
  INV_X1 U11 ( .A(n37), .ZN(n54) );
  INV_X1 U12 ( .A(a[2]), .ZN(n53) );
  INV_X1 U13 ( .A(n35), .ZN(n52) );
  INV_X1 U14 ( .A(a[1]), .ZN(n51) );
  INV_X1 U15 ( .A(n33), .ZN(n50) );
  INV_X1 U16 ( .A(a[0]), .ZN(n49) );
  OR2_X1 U17 ( .A1(n48), .A2(n64), .ZN(y[7]) );
  OR2_X1 U18 ( .A1(n63), .A2(b[7]), .ZN(n47) );
  AND2_X1 U19 ( .A1(b[7]), .A2(n63), .ZN(n48) );
  OR2_X1 U20 ( .A1(n46), .A2(n62), .ZN(y[6]) );
  OR2_X1 U21 ( .A1(n61), .A2(b[6]), .ZN(n45) );
  AND2_X1 U22 ( .A1(b[6]), .A2(n61), .ZN(n46) );
  OR2_X1 U23 ( .A1(n44), .A2(n60), .ZN(y[5]) );
  OR2_X1 U24 ( .A1(n59), .A2(b[5]), .ZN(n43) );
  AND2_X1 U25 ( .A1(b[5]), .A2(n59), .ZN(n44) );
  OR2_X1 U26 ( .A1(n42), .A2(n58), .ZN(y[4]) );
  OR2_X1 U27 ( .A1(n57), .A2(b[4]), .ZN(n41) );
  AND2_X1 U28 ( .A1(b[4]), .A2(n57), .ZN(n42) );
  OR2_X1 U29 ( .A1(n40), .A2(n56), .ZN(y[3]) );
  OR2_X1 U30 ( .A1(n55), .A2(b[3]), .ZN(n39) );
  AND2_X1 U31 ( .A1(b[3]), .A2(n55), .ZN(n40) );
  OR2_X1 U32 ( .A1(n38), .A2(n54), .ZN(y[2]) );
  OR2_X1 U33 ( .A1(n53), .A2(b[2]), .ZN(n37) );
  AND2_X1 U34 ( .A1(b[2]), .A2(n53), .ZN(n38) );
  OR2_X1 U35 ( .A1(n36), .A2(n52), .ZN(y[1]) );
  OR2_X1 U36 ( .A1(n51), .A2(b[1]), .ZN(n35) );
  AND2_X1 U37 ( .A1(b[1]), .A2(n51), .ZN(n36) );
  OR2_X1 U38 ( .A1(n34), .A2(n50), .ZN(y[0]) );
  OR2_X1 U39 ( .A1(n49), .A2(b[0]), .ZN(n33) );
  AND2_X1 U40 ( .A1(b[0]), .A2(n49), .ZN(n34) );
endmodule


module byteXor_4 ( a, b, y );
  input [7:0] a;
  input [7:0] b;
  //input_done

  output [7:0] y;
  //output_done

  wire   n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64;
  //wire_done

  INV_X1 U1 ( .A(n47), .ZN(n64) );
  INV_X1 U2 ( .A(a[7]), .ZN(n63) );
  INV_X1 U3 ( .A(n45), .ZN(n62) );
  INV_X1 U4 ( .A(a[6]), .ZN(n61) );
  INV_X1 U5 ( .A(n43), .ZN(n60) );
  INV_X1 U6 ( .A(a[5]), .ZN(n59) );
  INV_X1 U7 ( .A(n41), .ZN(n58) );
  INV_X1 U8 ( .A(a[4]), .ZN(n57) );
  INV_X1 U9 ( .A(n39), .ZN(n56) );
  INV_X1 U10 ( .A(a[3]), .ZN(n55) );
  INV_X1 U11 ( .A(n37), .ZN(n54) );
  INV_X1 U12 ( .A(a[2]), .ZN(n53) );
  INV_X1 U13 ( .A(n35), .ZN(n52) );
  INV_X1 U14 ( .A(a[1]), .ZN(n51) );
  INV_X1 U15 ( .A(n33), .ZN(n50) );
  INV_X1 U16 ( .A(a[0]), .ZN(n49) );
  OR2_X1 U17 ( .A1(n48), .A2(n64), .ZN(y[7]) );
  OR2_X1 U18 ( .A1(n63), .A2(b[7]), .ZN(n47) );
  AND2_X1 U19 ( .A1(b[7]), .A2(n63), .ZN(n48) );
  OR2_X1 U20 ( .A1(n46), .A2(n62), .ZN(y[6]) );
  OR2_X1 U21 ( .A1(n61), .A2(b[6]), .ZN(n45) );
  AND2_X1 U22 ( .A1(b[6]), .A2(n61), .ZN(n46) );
  OR2_X1 U23 ( .A1(n44), .A2(n60), .ZN(y[5]) );
  OR2_X1 U24 ( .A1(n59), .A2(b[5]), .ZN(n43) );
  AND2_X1 U25 ( .A1(b[5]), .A2(n59), .ZN(n44) );
  OR2_X1 U26 ( .A1(n42), .A2(n58), .ZN(y[4]) );
  OR2_X1 U27 ( .A1(n57), .A2(b[4]), .ZN(n41) );
  AND2_X1 U28 ( .A1(b[4]), .A2(n57), .ZN(n42) );
  OR2_X1 U29 ( .A1(n40), .A2(n56), .ZN(y[3]) );
  OR2_X1 U30 ( .A1(n55), .A2(b[3]), .ZN(n39) );
  AND2_X1 U31 ( .A1(b[3]), .A2(n55), .ZN(n40) );
  OR2_X1 U32 ( .A1(n38), .A2(n54), .ZN(y[2]) );
  OR2_X1 U33 ( .A1(n53), .A2(b[2]), .ZN(n37) );
  AND2_X1 U34 ( .A1(b[2]), .A2(n53), .ZN(n38) );
  OR2_X1 U35 ( .A1(n36), .A2(n52), .ZN(y[1]) );
  OR2_X1 U36 ( .A1(n51), .A2(b[1]), .ZN(n35) );
  AND2_X1 U37 ( .A1(b[1]), .A2(n51), .ZN(n36) );
  OR2_X1 U38 ( .A1(n34), .A2(n50), .ZN(y[0]) );
  OR2_X1 U39 ( .A1(n49), .A2(b[0]), .ZN(n33) );
  AND2_X1 U40 ( .A1(b[0]), .A2(n49), .ZN(n34) );
endmodule


module byteXor_5 ( a, b, y );
  input [7:0] a;
  input [7:0] b;
  //input_done

  output [7:0] y;
  //output_done

  wire   n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64;
  //wire_done

  INV_X1 U1 ( .A(n47), .ZN(n64) );
  INV_X1 U2 ( .A(a[7]), .ZN(n63) );
  INV_X1 U3 ( .A(n45), .ZN(n62) );
  INV_X1 U4 ( .A(a[6]), .ZN(n61) );
  INV_X1 U5 ( .A(n43), .ZN(n60) );
  INV_X1 U6 ( .A(a[5]), .ZN(n59) );
  INV_X1 U7 ( .A(n41), .ZN(n58) );
  INV_X1 U8 ( .A(a[4]), .ZN(n57) );
  INV_X1 U9 ( .A(n39), .ZN(n56) );
  INV_X1 U10 ( .A(a[3]), .ZN(n55) );
  INV_X1 U11 ( .A(n37), .ZN(n54) );
  INV_X1 U12 ( .A(a[2]), .ZN(n53) );
  INV_X1 U13 ( .A(n35), .ZN(n52) );
  INV_X1 U14 ( .A(a[1]), .ZN(n51) );
  INV_X1 U15 ( .A(n33), .ZN(n50) );
  INV_X1 U16 ( .A(a[0]), .ZN(n49) );
  OR2_X1 U17 ( .A1(n48), .A2(n64), .ZN(y[7]) );
  OR2_X1 U18 ( .A1(n63), .A2(b[7]), .ZN(n47) );
  AND2_X1 U19 ( .A1(b[7]), .A2(n63), .ZN(n48) );
  OR2_X1 U20 ( .A1(n46), .A2(n62), .ZN(y[6]) );
  OR2_X1 U21 ( .A1(n61), .A2(b[6]), .ZN(n45) );
  AND2_X1 U22 ( .A1(b[6]), .A2(n61), .ZN(n46) );
  OR2_X1 U23 ( .A1(n44), .A2(n60), .ZN(y[5]) );
  OR2_X1 U24 ( .A1(n59), .A2(b[5]), .ZN(n43) );
  AND2_X1 U25 ( .A1(b[5]), .A2(n59), .ZN(n44) );
  OR2_X1 U26 ( .A1(n42), .A2(n58), .ZN(y[4]) );
  OR2_X1 U27 ( .A1(n57), .A2(b[4]), .ZN(n41) );
  AND2_X1 U28 ( .A1(b[4]), .A2(n57), .ZN(n42) );
  OR2_X1 U29 ( .A1(n40), .A2(n56), .ZN(y[3]) );
  OR2_X1 U30 ( .A1(n55), .A2(b[3]), .ZN(n39) );
  AND2_X1 U31 ( .A1(b[3]), .A2(n55), .ZN(n40) );
  OR2_X1 U32 ( .A1(n38), .A2(n54), .ZN(y[2]) );
  OR2_X1 U33 ( .A1(n53), .A2(b[2]), .ZN(n37) );
  AND2_X1 U34 ( .A1(b[2]), .A2(n53), .ZN(n38) );
  OR2_X1 U35 ( .A1(n36), .A2(n52), .ZN(y[1]) );
  OR2_X1 U36 ( .A1(n51), .A2(b[1]), .ZN(n35) );
  AND2_X1 U37 ( .A1(b[1]), .A2(n51), .ZN(n36) );
  OR2_X1 U38 ( .A1(n34), .A2(n50), .ZN(y[0]) );
  OR2_X1 U39 ( .A1(n49), .A2(b[0]), .ZN(n33) );
  AND2_X1 U40 ( .A1(b[0]), .A2(n49), .ZN(n34) );
endmodule


module byteXor4_1 ( a, b, c, d, y );
  input [7:0] a;
  input [7:0] b;
  input [7:0] c;
  input [7:0] d;
  //input_done

  output [7:0] y;
  //output_done

  wire   n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224;
  //wire_done

  INV_X1 U1 ( .A(n175), .ZN(n224) );
  INV_X1 U2 ( .A(a[7]), .ZN(n223) );
  INV_X1 U3 ( .A(n167), .ZN(n222) );
  INV_X1 U4 ( .A(a[6]), .ZN(n221) );
  INV_X1 U5 ( .A(n159), .ZN(n220) );
  INV_X1 U6 ( .A(a[5]), .ZN(n219) );
  INV_X1 U7 ( .A(n151), .ZN(n218) );
  INV_X1 U8 ( .A(a[4]), .ZN(n217) );
  INV_X1 U9 ( .A(n143), .ZN(n216) );
  INV_X1 U10 ( .A(a[3]), .ZN(n215) );
  INV_X1 U11 ( .A(n135), .ZN(n214) );
  INV_X1 U12 ( .A(a[2]), .ZN(n213) );
  INV_X1 U13 ( .A(n127), .ZN(n212) );
  INV_X1 U14 ( .A(a[1]), .ZN(n211) );
  INV_X1 U15 ( .A(n119), .ZN(n210) );
  INV_X1 U16 ( .A(a[0]), .ZN(n209) );
  INV_X1 U17 ( .A(b[7]), .ZN(n208) );
  INV_X1 U18 ( .A(b[6]), .ZN(n207) );
  INV_X1 U19 ( .A(b[5]), .ZN(n206) );
  INV_X1 U20 ( .A(b[4]), .ZN(n205) );
  INV_X1 U21 ( .A(b[3]), .ZN(n204) );
  INV_X1 U22 ( .A(b[2]), .ZN(n203) );
  INV_X1 U23 ( .A(b[1]), .ZN(n202) );
  INV_X1 U24 ( .A(b[0]), .ZN(n201) );
  INV_X1 U25 ( .A(n171), .ZN(n200) );
  INV_X1 U26 ( .A(c[7]), .ZN(n199) );
  INV_X1 U27 ( .A(n163), .ZN(n198) );
  INV_X1 U28 ( .A(c[6]), .ZN(n197) );
  INV_X1 U29 ( .A(n155), .ZN(n196) );
  INV_X1 U30 ( .A(c[5]), .ZN(n195) );
  INV_X1 U31 ( .A(n147), .ZN(n194) );
  INV_X1 U32 ( .A(c[4]), .ZN(n193) );
  INV_X1 U33 ( .A(n139), .ZN(n192) );
  INV_X1 U34 ( .A(c[3]), .ZN(n191) );
  INV_X1 U35 ( .A(n131), .ZN(n190) );
  INV_X1 U36 ( .A(c[2]), .ZN(n189) );
  INV_X1 U37 ( .A(n123), .ZN(n188) );
  INV_X1 U38 ( .A(c[1]), .ZN(n187) );
  INV_X1 U39 ( .A(n115), .ZN(n186) );
  INV_X1 U40 ( .A(c[0]), .ZN(n185) );
  INV_X1 U41 ( .A(d[7]), .ZN(n184) );
  INV_X1 U42 ( .A(d[6]), .ZN(n183) );
  INV_X1 U43 ( .A(d[5]), .ZN(n182) );
  INV_X1 U44 ( .A(d[4]), .ZN(n181) );
  INV_X1 U45 ( .A(d[3]), .ZN(n180) );
  INV_X1 U46 ( .A(d[2]), .ZN(n179) );
  INV_X1 U47 ( .A(d[1]), .ZN(n178) );
  INV_X1 U48 ( .A(d[0]), .ZN(n177) );
  OR2_X1 U49 ( .A1(n176), .A2(n224), .ZN(y[7]) );
  OR2_X1 U50 ( .A1(n174), .A2(n200), .ZN(n175) );
  AND2_X1 U51 ( .A1(n200), .A2(n174), .ZN(n176) );
  AND2_X1 U52 ( .A1(n173), .A2(n172), .ZN(n174) );
  OR2_X1 U53 ( .A1(n223), .A2(b[7]), .ZN(n172) );
  OR2_X1 U54 ( .A1(n208), .A2(a[7]), .ZN(n173) );
  AND2_X1 U55 ( .A1(n170), .A2(n169), .ZN(n171) );
  OR2_X1 U56 ( .A1(n199), .A2(d[7]), .ZN(n169) );
  OR2_X1 U57 ( .A1(n184), .A2(c[7]), .ZN(n170) );
  OR2_X1 U58 ( .A1(n168), .A2(n222), .ZN(y[6]) );
  OR2_X1 U59 ( .A1(n166), .A2(n198), .ZN(n167) );
  AND2_X1 U60 ( .A1(n198), .A2(n166), .ZN(n168) );
  AND2_X1 U61 ( .A1(n165), .A2(n164), .ZN(n166) );
  OR2_X1 U62 ( .A1(n221), .A2(b[6]), .ZN(n164) );
  OR2_X1 U63 ( .A1(n207), .A2(a[6]), .ZN(n165) );
  AND2_X1 U64 ( .A1(n162), .A2(n161), .ZN(n163) );
  OR2_X1 U65 ( .A1(n197), .A2(d[6]), .ZN(n161) );
  OR2_X1 U66 ( .A1(n183), .A2(c[6]), .ZN(n162) );
  OR2_X1 U67 ( .A1(n160), .A2(n220), .ZN(y[5]) );
  OR2_X1 U68 ( .A1(n158), .A2(n196), .ZN(n159) );
  AND2_X1 U69 ( .A1(n196), .A2(n158), .ZN(n160) );
  AND2_X1 U70 ( .A1(n157), .A2(n156), .ZN(n158) );
  OR2_X1 U71 ( .A1(n219), .A2(b[5]), .ZN(n156) );
  OR2_X1 U72 ( .A1(n206), .A2(a[5]), .ZN(n157) );
  AND2_X1 U73 ( .A1(n154), .A2(n153), .ZN(n155) );
  OR2_X1 U74 ( .A1(n195), .A2(d[5]), .ZN(n153) );
  OR2_X1 U75 ( .A1(n182), .A2(c[5]), .ZN(n154) );
  OR2_X1 U76 ( .A1(n152), .A2(n218), .ZN(y[4]) );
  OR2_X1 U77 ( .A1(n150), .A2(n194), .ZN(n151) );
  AND2_X1 U78 ( .A1(n194), .A2(n150), .ZN(n152) );
  AND2_X1 U79 ( .A1(n149), .A2(n148), .ZN(n150) );
  OR2_X1 U80 ( .A1(n217), .A2(b[4]), .ZN(n148) );
  OR2_X1 U81 ( .A1(n205), .A2(a[4]), .ZN(n149) );
  AND2_X1 U82 ( .A1(n146), .A2(n145), .ZN(n147) );
  OR2_X1 U83 ( .A1(n193), .A2(d[4]), .ZN(n145) );
  OR2_X1 U84 ( .A1(n181), .A2(c[4]), .ZN(n146) );
  OR2_X1 U85 ( .A1(n144), .A2(n216), .ZN(y[3]) );
  OR2_X1 U86 ( .A1(n142), .A2(n192), .ZN(n143) );
  AND2_X1 U87 ( .A1(n192), .A2(n142), .ZN(n144) );
  AND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(n142) );
  OR2_X1 U89 ( .A1(n215), .A2(b[3]), .ZN(n140) );
  OR2_X1 U90 ( .A1(n204), .A2(a[3]), .ZN(n141) );
  AND2_X1 U91 ( .A1(n138), .A2(n137), .ZN(n139) );
  OR2_X1 U92 ( .A1(n191), .A2(d[3]), .ZN(n137) );
  OR2_X1 U93 ( .A1(n180), .A2(c[3]), .ZN(n138) );
  OR2_X1 U94 ( .A1(n136), .A2(n214), .ZN(y[2]) );
  OR2_X1 U95 ( .A1(n134), .A2(n190), .ZN(n135) );
  AND2_X1 U96 ( .A1(n190), .A2(n134), .ZN(n136) );
  AND2_X1 U97 ( .A1(n133), .A2(n132), .ZN(n134) );
  OR2_X1 U98 ( .A1(n213), .A2(b[2]), .ZN(n132) );
  OR2_X1 U99 ( .A1(n203), .A2(a[2]), .ZN(n133) );
  AND2_X1 U100 ( .A1(n130), .A2(n129), .ZN(n131) );
  OR2_X1 U101 ( .A1(n189), .A2(d[2]), .ZN(n129) );
  OR2_X1 U102 ( .A1(n179), .A2(c[2]), .ZN(n130) );
  OR2_X1 U103 ( .A1(n128), .A2(n212), .ZN(y[1]) );
  OR2_X1 U104 ( .A1(n126), .A2(n188), .ZN(n127) );
  AND2_X1 U105 ( .A1(n188), .A2(n126), .ZN(n128) );
  AND2_X1 U106 ( .A1(n125), .A2(n124), .ZN(n126) );
  OR2_X1 U107 ( .A1(n211), .A2(b[1]), .ZN(n124) );
  OR2_X1 U108 ( .A1(n202), .A2(a[1]), .ZN(n125) );
  AND2_X1 U109 ( .A1(n122), .A2(n121), .ZN(n123) );
  OR2_X1 U110 ( .A1(n187), .A2(d[1]), .ZN(n121) );
  OR2_X1 U111 ( .A1(n178), .A2(c[1]), .ZN(n122) );
  OR2_X1 U112 ( .A1(n120), .A2(n210), .ZN(y[0]) );
  OR2_X1 U113 ( .A1(n118), .A2(n186), .ZN(n119) );
  AND2_X1 U114 ( .A1(n186), .A2(n118), .ZN(n120) );
  AND2_X1 U115 ( .A1(n117), .A2(n116), .ZN(n118) );
  OR2_X1 U116 ( .A1(n209), .A2(b[0]), .ZN(n116) );
  OR2_X1 U117 ( .A1(n201), .A2(a[0]), .ZN(n117) );
  AND2_X1 U118 ( .A1(n114), .A2(n113), .ZN(n115) );
  OR2_X1 U119 ( .A1(n185), .A2(d[0]), .ZN(n113) );
  OR2_X1 U120 ( .A1(n177), .A2(c[0]), .ZN(n114) );
endmodule


module byteXor4_2 ( a, b, c, d, y );
  input [7:0] a;
  input [7:0] b;
  input [7:0] c;
  input [7:0] d;
  //input_done

  output [7:0] y;
  //output_done

  wire   n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224;
  //wire_done

  INV_X1 U1 ( .A(n175), .ZN(n224) );
  INV_X1 U2 ( .A(a[7]), .ZN(n223) );
  INV_X1 U3 ( .A(n167), .ZN(n222) );
  INV_X1 U4 ( .A(a[6]), .ZN(n221) );
  INV_X1 U5 ( .A(n159), .ZN(n220) );
  INV_X1 U6 ( .A(a[5]), .ZN(n219) );
  INV_X1 U7 ( .A(n151), .ZN(n218) );
  INV_X1 U8 ( .A(a[4]), .ZN(n217) );
  INV_X1 U9 ( .A(n143), .ZN(n216) );
  INV_X1 U10 ( .A(a[3]), .ZN(n215) );
  INV_X1 U11 ( .A(n135), .ZN(n214) );
  INV_X1 U12 ( .A(a[2]), .ZN(n213) );
  INV_X1 U13 ( .A(n127), .ZN(n212) );
  INV_X1 U14 ( .A(a[1]), .ZN(n211) );
  INV_X1 U15 ( .A(n119), .ZN(n210) );
  INV_X1 U16 ( .A(a[0]), .ZN(n209) );
  INV_X1 U17 ( .A(b[7]), .ZN(n208) );
  INV_X1 U18 ( .A(b[6]), .ZN(n207) );
  INV_X1 U19 ( .A(b[5]), .ZN(n206) );
  INV_X1 U20 ( .A(b[4]), .ZN(n205) );
  INV_X1 U21 ( .A(b[3]), .ZN(n204) );
  INV_X1 U22 ( .A(b[2]), .ZN(n203) );
  INV_X1 U23 ( .A(b[1]), .ZN(n202) );
  INV_X1 U24 ( .A(b[0]), .ZN(n201) );
  INV_X1 U25 ( .A(n171), .ZN(n200) );
  INV_X1 U26 ( .A(c[7]), .ZN(n199) );
  INV_X1 U27 ( .A(n163), .ZN(n198) );
  INV_X1 U28 ( .A(c[6]), .ZN(n197) );
  INV_X1 U29 ( .A(n155), .ZN(n196) );
  INV_X1 U30 ( .A(c[5]), .ZN(n195) );
  INV_X1 U31 ( .A(n147), .ZN(n194) );
  INV_X1 U32 ( .A(c[4]), .ZN(n193) );
  INV_X1 U33 ( .A(n139), .ZN(n192) );
  INV_X1 U34 ( .A(c[3]), .ZN(n191) );
  INV_X1 U35 ( .A(n131), .ZN(n190) );
  INV_X1 U36 ( .A(c[2]), .ZN(n189) );
  INV_X1 U37 ( .A(n123), .ZN(n188) );
  INV_X1 U38 ( .A(c[1]), .ZN(n187) );
  INV_X1 U39 ( .A(n115), .ZN(n186) );
  INV_X1 U40 ( .A(c[0]), .ZN(n185) );
  INV_X1 U41 ( .A(d[7]), .ZN(n184) );
  INV_X1 U42 ( .A(d[6]), .ZN(n183) );
  INV_X1 U43 ( .A(d[5]), .ZN(n182) );
  INV_X1 U44 ( .A(d[4]), .ZN(n181) );
  INV_X1 U45 ( .A(d[3]), .ZN(n180) );
  INV_X1 U46 ( .A(d[2]), .ZN(n179) );
  INV_X1 U47 ( .A(d[1]), .ZN(n178) );
  INV_X1 U48 ( .A(d[0]), .ZN(n177) );
  OR2_X1 U49 ( .A1(n176), .A2(n224), .ZN(y[7]) );
  OR2_X1 U50 ( .A1(n174), .A2(n200), .ZN(n175) );
  AND2_X1 U51 ( .A1(n200), .A2(n174), .ZN(n176) );
  AND2_X1 U52 ( .A1(n173), .A2(n172), .ZN(n174) );
  OR2_X1 U53 ( .A1(n223), .A2(b[7]), .ZN(n172) );
  OR2_X1 U54 ( .A1(n208), .A2(a[7]), .ZN(n173) );
  AND2_X1 U55 ( .A1(n170), .A2(n169), .ZN(n171) );
  OR2_X1 U56 ( .A1(n199), .A2(d[7]), .ZN(n169) );
  OR2_X1 U57 ( .A1(n184), .A2(c[7]), .ZN(n170) );
  OR2_X1 U58 ( .A1(n168), .A2(n222), .ZN(y[6]) );
  OR2_X1 U59 ( .A1(n166), .A2(n198), .ZN(n167) );
  AND2_X1 U60 ( .A1(n198), .A2(n166), .ZN(n168) );
  AND2_X1 U61 ( .A1(n165), .A2(n164), .ZN(n166) );
  OR2_X1 U62 ( .A1(n221), .A2(b[6]), .ZN(n164) );
  OR2_X1 U63 ( .A1(n207), .A2(a[6]), .ZN(n165) );
  AND2_X1 U64 ( .A1(n162), .A2(n161), .ZN(n163) );
  OR2_X1 U65 ( .A1(n197), .A2(d[6]), .ZN(n161) );
  OR2_X1 U66 ( .A1(n183), .A2(c[6]), .ZN(n162) );
  OR2_X1 U67 ( .A1(n160), .A2(n220), .ZN(y[5]) );
  OR2_X1 U68 ( .A1(n158), .A2(n196), .ZN(n159) );
  AND2_X1 U69 ( .A1(n196), .A2(n158), .ZN(n160) );
  AND2_X1 U70 ( .A1(n157), .A2(n156), .ZN(n158) );
  OR2_X1 U71 ( .A1(n219), .A2(b[5]), .ZN(n156) );
  OR2_X1 U72 ( .A1(n206), .A2(a[5]), .ZN(n157) );
  AND2_X1 U73 ( .A1(n154), .A2(n153), .ZN(n155) );
  OR2_X1 U74 ( .A1(n195), .A2(d[5]), .ZN(n153) );
  OR2_X1 U75 ( .A1(n182), .A2(c[5]), .ZN(n154) );
  OR2_X1 U76 ( .A1(n152), .A2(n218), .ZN(y[4]) );
  OR2_X1 U77 ( .A1(n150), .A2(n194), .ZN(n151) );
  AND2_X1 U78 ( .A1(n194), .A2(n150), .ZN(n152) );
  AND2_X1 U79 ( .A1(n149), .A2(n148), .ZN(n150) );
  OR2_X1 U80 ( .A1(n217), .A2(b[4]), .ZN(n148) );
  OR2_X1 U81 ( .A1(n205), .A2(a[4]), .ZN(n149) );
  AND2_X1 U82 ( .A1(n146), .A2(n145), .ZN(n147) );
  OR2_X1 U83 ( .A1(n193), .A2(d[4]), .ZN(n145) );
  OR2_X1 U84 ( .A1(n181), .A2(c[4]), .ZN(n146) );
  OR2_X1 U85 ( .A1(n144), .A2(n216), .ZN(y[3]) );
  OR2_X1 U86 ( .A1(n142), .A2(n192), .ZN(n143) );
  AND2_X1 U87 ( .A1(n192), .A2(n142), .ZN(n144) );
  AND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(n142) );
  OR2_X1 U89 ( .A1(n215), .A2(b[3]), .ZN(n140) );
  OR2_X1 U90 ( .A1(n204), .A2(a[3]), .ZN(n141) );
  AND2_X1 U91 ( .A1(n138), .A2(n137), .ZN(n139) );
  OR2_X1 U92 ( .A1(n191), .A2(d[3]), .ZN(n137) );
  OR2_X1 U93 ( .A1(n180), .A2(c[3]), .ZN(n138) );
  OR2_X1 U94 ( .A1(n136), .A2(n214), .ZN(y[2]) );
  OR2_X1 U95 ( .A1(n134), .A2(n190), .ZN(n135) );
  AND2_X1 U96 ( .A1(n190), .A2(n134), .ZN(n136) );
  AND2_X1 U97 ( .A1(n133), .A2(n132), .ZN(n134) );
  OR2_X1 U98 ( .A1(n213), .A2(b[2]), .ZN(n132) );
  OR2_X1 U99 ( .A1(n203), .A2(a[2]), .ZN(n133) );
  AND2_X1 U100 ( .A1(n130), .A2(n129), .ZN(n131) );
  OR2_X1 U101 ( .A1(n189), .A2(d[2]), .ZN(n129) );
  OR2_X1 U102 ( .A1(n179), .A2(c[2]), .ZN(n130) );
  OR2_X1 U103 ( .A1(n128), .A2(n212), .ZN(y[1]) );
  OR2_X1 U104 ( .A1(n126), .A2(n188), .ZN(n127) );
  AND2_X1 U105 ( .A1(n188), .A2(n126), .ZN(n128) );
  AND2_X1 U106 ( .A1(n125), .A2(n124), .ZN(n126) );
  OR2_X1 U107 ( .A1(n211), .A2(b[1]), .ZN(n124) );
  OR2_X1 U108 ( .A1(n202), .A2(a[1]), .ZN(n125) );
  AND2_X1 U109 ( .A1(n122), .A2(n121), .ZN(n123) );
  OR2_X1 U110 ( .A1(n187), .A2(d[1]), .ZN(n121) );
  OR2_X1 U111 ( .A1(n178), .A2(c[1]), .ZN(n122) );
  OR2_X1 U112 ( .A1(n120), .A2(n210), .ZN(y[0]) );
  OR2_X1 U113 ( .A1(n118), .A2(n186), .ZN(n119) );
  AND2_X1 U114 ( .A1(n186), .A2(n118), .ZN(n120) );
  AND2_X1 U115 ( .A1(n117), .A2(n116), .ZN(n118) );
  OR2_X1 U116 ( .A1(n209), .A2(b[0]), .ZN(n116) );
  OR2_X1 U117 ( .A1(n201), .A2(a[0]), .ZN(n117) );
  AND2_X1 U118 ( .A1(n114), .A2(n113), .ZN(n115) );
  OR2_X1 U119 ( .A1(n185), .A2(d[0]), .ZN(n113) );
  OR2_X1 U120 ( .A1(n177), .A2(c[0]), .ZN(n114) );
endmodule


module byteXor4_3 ( a, b, c, d, y );
  input [7:0] a;
  input [7:0] b;
  input [7:0] c;
  input [7:0] d;
  //input_done

  output [7:0] y;
  //output_done

  wire   n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224;
  //wire_done

  INV_X1 U1 ( .A(n175), .ZN(n224) );
  INV_X1 U2 ( .A(a[7]), .ZN(n223) );
  INV_X1 U3 ( .A(n167), .ZN(n222) );
  INV_X1 U4 ( .A(a[6]), .ZN(n221) );
  INV_X1 U5 ( .A(n159), .ZN(n220) );
  INV_X1 U6 ( .A(a[5]), .ZN(n219) );
  INV_X1 U7 ( .A(n151), .ZN(n218) );
  INV_X1 U8 ( .A(a[4]), .ZN(n217) );
  INV_X1 U9 ( .A(n143), .ZN(n216) );
  INV_X1 U10 ( .A(a[3]), .ZN(n215) );
  INV_X1 U11 ( .A(n135), .ZN(n214) );
  INV_X1 U12 ( .A(a[2]), .ZN(n213) );
  INV_X1 U13 ( .A(n127), .ZN(n212) );
  INV_X1 U14 ( .A(a[1]), .ZN(n211) );
  INV_X1 U15 ( .A(n119), .ZN(n210) );
  INV_X1 U16 ( .A(a[0]), .ZN(n209) );
  INV_X1 U17 ( .A(b[7]), .ZN(n208) );
  INV_X1 U18 ( .A(b[6]), .ZN(n207) );
  INV_X1 U19 ( .A(b[5]), .ZN(n206) );
  INV_X1 U20 ( .A(b[4]), .ZN(n205) );
  INV_X1 U21 ( .A(b[3]), .ZN(n204) );
  INV_X1 U22 ( .A(b[2]), .ZN(n203) );
  INV_X1 U23 ( .A(b[1]), .ZN(n202) );
  INV_X1 U24 ( .A(b[0]), .ZN(n201) );
  INV_X1 U25 ( .A(n171), .ZN(n200) );
  INV_X1 U26 ( .A(c[7]), .ZN(n199) );
  INV_X1 U27 ( .A(n163), .ZN(n198) );
  INV_X1 U28 ( .A(c[6]), .ZN(n197) );
  INV_X1 U29 ( .A(n155), .ZN(n196) );
  INV_X1 U30 ( .A(c[5]), .ZN(n195) );
  INV_X1 U31 ( .A(n147), .ZN(n194) );
  INV_X1 U32 ( .A(c[4]), .ZN(n193) );
  INV_X1 U33 ( .A(n139), .ZN(n192) );
  INV_X1 U34 ( .A(c[3]), .ZN(n191) );
  INV_X1 U35 ( .A(n131), .ZN(n190) );
  INV_X1 U36 ( .A(c[2]), .ZN(n189) );
  INV_X1 U37 ( .A(n123), .ZN(n188) );
  INV_X1 U38 ( .A(c[1]), .ZN(n187) );
  INV_X1 U39 ( .A(n115), .ZN(n186) );
  INV_X1 U40 ( .A(c[0]), .ZN(n185) );
  INV_X1 U41 ( .A(d[7]), .ZN(n184) );
  INV_X1 U42 ( .A(d[6]), .ZN(n183) );
  INV_X1 U43 ( .A(d[5]), .ZN(n182) );
  INV_X1 U44 ( .A(d[4]), .ZN(n181) );
  INV_X1 U45 ( .A(d[3]), .ZN(n180) );
  INV_X1 U46 ( .A(d[2]), .ZN(n179) );
  INV_X1 U47 ( .A(d[1]), .ZN(n178) );
  INV_X1 U48 ( .A(d[0]), .ZN(n177) );
  OR2_X1 U49 ( .A1(n176), .A2(n224), .ZN(y[7]) );
  OR2_X1 U50 ( .A1(n174), .A2(n200), .ZN(n175) );
  AND2_X1 U51 ( .A1(n200), .A2(n174), .ZN(n176) );
  AND2_X1 U52 ( .A1(n173), .A2(n172), .ZN(n174) );
  OR2_X1 U53 ( .A1(n223), .A2(b[7]), .ZN(n172) );
  OR2_X1 U54 ( .A1(n208), .A2(a[7]), .ZN(n173) );
  AND2_X1 U55 ( .A1(n170), .A2(n169), .ZN(n171) );
  OR2_X1 U56 ( .A1(n199), .A2(d[7]), .ZN(n169) );
  OR2_X1 U57 ( .A1(n184), .A2(c[7]), .ZN(n170) );
  OR2_X1 U58 ( .A1(n168), .A2(n222), .ZN(y[6]) );
  OR2_X1 U59 ( .A1(n166), .A2(n198), .ZN(n167) );
  AND2_X1 U60 ( .A1(n198), .A2(n166), .ZN(n168) );
  AND2_X1 U61 ( .A1(n165), .A2(n164), .ZN(n166) );
  OR2_X1 U62 ( .A1(n221), .A2(b[6]), .ZN(n164) );
  OR2_X1 U63 ( .A1(n207), .A2(a[6]), .ZN(n165) );
  AND2_X1 U64 ( .A1(n162), .A2(n161), .ZN(n163) );
  OR2_X1 U65 ( .A1(n197), .A2(d[6]), .ZN(n161) );
  OR2_X1 U66 ( .A1(n183), .A2(c[6]), .ZN(n162) );
  OR2_X1 U67 ( .A1(n160), .A2(n220), .ZN(y[5]) );
  OR2_X1 U68 ( .A1(n158), .A2(n196), .ZN(n159) );
  AND2_X1 U69 ( .A1(n196), .A2(n158), .ZN(n160) );
  AND2_X1 U70 ( .A1(n157), .A2(n156), .ZN(n158) );
  OR2_X1 U71 ( .A1(n219), .A2(b[5]), .ZN(n156) );
  OR2_X1 U72 ( .A1(n206), .A2(a[5]), .ZN(n157) );
  AND2_X1 U73 ( .A1(n154), .A2(n153), .ZN(n155) );
  OR2_X1 U74 ( .A1(n195), .A2(d[5]), .ZN(n153) );
  OR2_X1 U75 ( .A1(n182), .A2(c[5]), .ZN(n154) );
  OR2_X1 U76 ( .A1(n152), .A2(n218), .ZN(y[4]) );
  OR2_X1 U77 ( .A1(n150), .A2(n194), .ZN(n151) );
  AND2_X1 U78 ( .A1(n194), .A2(n150), .ZN(n152) );
  AND2_X1 U79 ( .A1(n149), .A2(n148), .ZN(n150) );
  OR2_X1 U80 ( .A1(n217), .A2(b[4]), .ZN(n148) );
  OR2_X1 U81 ( .A1(n205), .A2(a[4]), .ZN(n149) );
  AND2_X1 U82 ( .A1(n146), .A2(n145), .ZN(n147) );
  OR2_X1 U83 ( .A1(n193), .A2(d[4]), .ZN(n145) );
  OR2_X1 U84 ( .A1(n181), .A2(c[4]), .ZN(n146) );
  OR2_X1 U85 ( .A1(n144), .A2(n216), .ZN(y[3]) );
  OR2_X1 U86 ( .A1(n142), .A2(n192), .ZN(n143) );
  AND2_X1 U87 ( .A1(n192), .A2(n142), .ZN(n144) );
  AND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(n142) );
  OR2_X1 U89 ( .A1(n215), .A2(b[3]), .ZN(n140) );
  OR2_X1 U90 ( .A1(n204), .A2(a[3]), .ZN(n141) );
  AND2_X1 U91 ( .A1(n138), .A2(n137), .ZN(n139) );
  OR2_X1 U92 ( .A1(n191), .A2(d[3]), .ZN(n137) );
  OR2_X1 U93 ( .A1(n180), .A2(c[3]), .ZN(n138) );
  OR2_X1 U94 ( .A1(n136), .A2(n214), .ZN(y[2]) );
  OR2_X1 U95 ( .A1(n134), .A2(n190), .ZN(n135) );
  AND2_X1 U96 ( .A1(n190), .A2(n134), .ZN(n136) );
  AND2_X1 U97 ( .A1(n133), .A2(n132), .ZN(n134) );
  OR2_X1 U98 ( .A1(n213), .A2(b[2]), .ZN(n132) );
  OR2_X1 U99 ( .A1(n203), .A2(a[2]), .ZN(n133) );
  AND2_X1 U100 ( .A1(n130), .A2(n129), .ZN(n131) );
  OR2_X1 U101 ( .A1(n189), .A2(d[2]), .ZN(n129) );
  OR2_X1 U102 ( .A1(n179), .A2(c[2]), .ZN(n130) );
  OR2_X1 U103 ( .A1(n128), .A2(n212), .ZN(y[1]) );
  OR2_X1 U104 ( .A1(n126), .A2(n188), .ZN(n127) );
  AND2_X1 U105 ( .A1(n188), .A2(n126), .ZN(n128) );
  AND2_X1 U106 ( .A1(n125), .A2(n124), .ZN(n126) );
  OR2_X1 U107 ( .A1(n211), .A2(b[1]), .ZN(n124) );
  OR2_X1 U108 ( .A1(n202), .A2(a[1]), .ZN(n125) );
  AND2_X1 U109 ( .A1(n122), .A2(n121), .ZN(n123) );
  OR2_X1 U110 ( .A1(n187), .A2(d[1]), .ZN(n121) );
  OR2_X1 U111 ( .A1(n178), .A2(c[1]), .ZN(n122) );
  OR2_X1 U112 ( .A1(n120), .A2(n210), .ZN(y[0]) );
  OR2_X1 U113 ( .A1(n118), .A2(n186), .ZN(n119) );
  AND2_X1 U114 ( .A1(n186), .A2(n118), .ZN(n120) );
  AND2_X1 U115 ( .A1(n117), .A2(n116), .ZN(n118) );
  OR2_X1 U116 ( .A1(n209), .A2(b[0]), .ZN(n116) );
  OR2_X1 U117 ( .A1(n201), .A2(a[0]), .ZN(n117) );
  AND2_X1 U118 ( .A1(n114), .A2(n113), .ZN(n115) );
  OR2_X1 U119 ( .A1(n185), .A2(d[0]), .ZN(n113) );
  OR2_X1 U120 ( .A1(n177), .A2(c[0]), .ZN(n114) );
endmodule


module byteXor4_4 ( a, b, c, d, y );
  input [7:0] a;
  input [7:0] b;
  input [7:0] c;
  input [7:0] d;
  //input_done

  output [7:0] y;
  //output_done

  wire   n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224;
  //wire_done

  INV_X1 U1 ( .A(n175), .ZN(n224) );
  INV_X1 U2 ( .A(a[7]), .ZN(n223) );
  INV_X1 U3 ( .A(n167), .ZN(n222) );
  INV_X1 U4 ( .A(a[6]), .ZN(n221) );
  INV_X1 U5 ( .A(n159), .ZN(n220) );
  INV_X1 U6 ( .A(a[5]), .ZN(n219) );
  INV_X1 U7 ( .A(n151), .ZN(n218) );
  INV_X1 U8 ( .A(a[4]), .ZN(n217) );
  INV_X1 U9 ( .A(n143), .ZN(n216) );
  INV_X1 U10 ( .A(a[3]), .ZN(n215) );
  INV_X1 U11 ( .A(n135), .ZN(n214) );
  INV_X1 U12 ( .A(a[2]), .ZN(n213) );
  INV_X1 U13 ( .A(n127), .ZN(n212) );
  INV_X1 U14 ( .A(a[1]), .ZN(n211) );
  INV_X1 U15 ( .A(n119), .ZN(n210) );
  INV_X1 U16 ( .A(a[0]), .ZN(n209) );
  INV_X1 U17 ( .A(b[7]), .ZN(n208) );
  INV_X1 U18 ( .A(b[6]), .ZN(n207) );
  INV_X1 U19 ( .A(b[5]), .ZN(n206) );
  INV_X1 U20 ( .A(b[4]), .ZN(n205) );
  INV_X1 U21 ( .A(b[3]), .ZN(n204) );
  INV_X1 U22 ( .A(b[2]), .ZN(n203) );
  INV_X1 U23 ( .A(b[1]), .ZN(n202) );
  INV_X1 U24 ( .A(b[0]), .ZN(n201) );
  INV_X1 U25 ( .A(n171), .ZN(n200) );
  INV_X1 U26 ( .A(c[7]), .ZN(n199) );
  INV_X1 U27 ( .A(n163), .ZN(n198) );
  INV_X1 U28 ( .A(c[6]), .ZN(n197) );
  INV_X1 U29 ( .A(n155), .ZN(n196) );
  INV_X1 U30 ( .A(c[5]), .ZN(n195) );
  INV_X1 U31 ( .A(n147), .ZN(n194) );
  INV_X1 U32 ( .A(c[4]), .ZN(n193) );
  INV_X1 U33 ( .A(n139), .ZN(n192) );
  INV_X1 U34 ( .A(c[3]), .ZN(n191) );
  INV_X1 U35 ( .A(n131), .ZN(n190) );
  INV_X1 U36 ( .A(c[2]), .ZN(n189) );
  INV_X1 U37 ( .A(n123), .ZN(n188) );
  INV_X1 U38 ( .A(c[1]), .ZN(n187) );
  INV_X1 U39 ( .A(n115), .ZN(n186) );
  INV_X1 U40 ( .A(c[0]), .ZN(n185) );
  INV_X1 U41 ( .A(d[7]), .ZN(n184) );
  INV_X1 U42 ( .A(d[6]), .ZN(n183) );
  INV_X1 U43 ( .A(d[5]), .ZN(n182) );
  INV_X1 U44 ( .A(d[4]), .ZN(n181) );
  INV_X1 U45 ( .A(d[3]), .ZN(n180) );
  INV_X1 U46 ( .A(d[2]), .ZN(n179) );
  INV_X1 U47 ( .A(d[1]), .ZN(n178) );
  INV_X1 U48 ( .A(d[0]), .ZN(n177) );
  OR2_X1 U49 ( .A1(n176), .A2(n224), .ZN(y[7]) );
  OR2_X1 U50 ( .A1(n174), .A2(n200), .ZN(n175) );
  AND2_X1 U51 ( .A1(n200), .A2(n174), .ZN(n176) );
  AND2_X1 U52 ( .A1(n173), .A2(n172), .ZN(n174) );
  OR2_X1 U53 ( .A1(n223), .A2(b[7]), .ZN(n172) );
  OR2_X1 U54 ( .A1(n208), .A2(a[7]), .ZN(n173) );
  AND2_X1 U55 ( .A1(n170), .A2(n169), .ZN(n171) );
  OR2_X1 U56 ( .A1(n199), .A2(d[7]), .ZN(n169) );
  OR2_X1 U57 ( .A1(n184), .A2(c[7]), .ZN(n170) );
  OR2_X1 U58 ( .A1(n168), .A2(n222), .ZN(y[6]) );
  OR2_X1 U59 ( .A1(n166), .A2(n198), .ZN(n167) );
  AND2_X1 U60 ( .A1(n198), .A2(n166), .ZN(n168) );
  AND2_X1 U61 ( .A1(n165), .A2(n164), .ZN(n166) );
  OR2_X1 U62 ( .A1(n221), .A2(b[6]), .ZN(n164) );
  OR2_X1 U63 ( .A1(n207), .A2(a[6]), .ZN(n165) );
  AND2_X1 U64 ( .A1(n162), .A2(n161), .ZN(n163) );
  OR2_X1 U65 ( .A1(n197), .A2(d[6]), .ZN(n161) );
  OR2_X1 U66 ( .A1(n183), .A2(c[6]), .ZN(n162) );
  OR2_X1 U67 ( .A1(n160), .A2(n220), .ZN(y[5]) );
  OR2_X1 U68 ( .A1(n158), .A2(n196), .ZN(n159) );
  AND2_X1 U69 ( .A1(n196), .A2(n158), .ZN(n160) );
  AND2_X1 U70 ( .A1(n157), .A2(n156), .ZN(n158) );
  OR2_X1 U71 ( .A1(n219), .A2(b[5]), .ZN(n156) );
  OR2_X1 U72 ( .A1(n206), .A2(a[5]), .ZN(n157) );
  AND2_X1 U73 ( .A1(n154), .A2(n153), .ZN(n155) );
  OR2_X1 U74 ( .A1(n195), .A2(d[5]), .ZN(n153) );
  OR2_X1 U75 ( .A1(n182), .A2(c[5]), .ZN(n154) );
  OR2_X1 U76 ( .A1(n152), .A2(n218), .ZN(y[4]) );
  OR2_X1 U77 ( .A1(n150), .A2(n194), .ZN(n151) );
  AND2_X1 U78 ( .A1(n194), .A2(n150), .ZN(n152) );
  AND2_X1 U79 ( .A1(n149), .A2(n148), .ZN(n150) );
  OR2_X1 U80 ( .A1(n217), .A2(b[4]), .ZN(n148) );
  OR2_X1 U81 ( .A1(n205), .A2(a[4]), .ZN(n149) );
  AND2_X1 U82 ( .A1(n146), .A2(n145), .ZN(n147) );
  OR2_X1 U83 ( .A1(n193), .A2(d[4]), .ZN(n145) );
  OR2_X1 U84 ( .A1(n181), .A2(c[4]), .ZN(n146) );
  OR2_X1 U85 ( .A1(n144), .A2(n216), .ZN(y[3]) );
  OR2_X1 U86 ( .A1(n142), .A2(n192), .ZN(n143) );
  AND2_X1 U87 ( .A1(n192), .A2(n142), .ZN(n144) );
  AND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(n142) );
  OR2_X1 U89 ( .A1(n215), .A2(b[3]), .ZN(n140) );
  OR2_X1 U90 ( .A1(n204), .A2(a[3]), .ZN(n141) );
  AND2_X1 U91 ( .A1(n138), .A2(n137), .ZN(n139) );
  OR2_X1 U92 ( .A1(n191), .A2(d[3]), .ZN(n137) );
  OR2_X1 U93 ( .A1(n180), .A2(c[3]), .ZN(n138) );
  OR2_X1 U94 ( .A1(n136), .A2(n214), .ZN(y[2]) );
  OR2_X1 U95 ( .A1(n134), .A2(n190), .ZN(n135) );
  AND2_X1 U96 ( .A1(n190), .A2(n134), .ZN(n136) );
  AND2_X1 U97 ( .A1(n133), .A2(n132), .ZN(n134) );
  OR2_X1 U98 ( .A1(n213), .A2(b[2]), .ZN(n132) );
  OR2_X1 U99 ( .A1(n203), .A2(a[2]), .ZN(n133) );
  AND2_X1 U100 ( .A1(n130), .A2(n129), .ZN(n131) );
  OR2_X1 U101 ( .A1(n189), .A2(d[2]), .ZN(n129) );
  OR2_X1 U102 ( .A1(n179), .A2(c[2]), .ZN(n130) );
  OR2_X1 U103 ( .A1(n128), .A2(n212), .ZN(y[1]) );
  OR2_X1 U104 ( .A1(n126), .A2(n188), .ZN(n127) );
  AND2_X1 U105 ( .A1(n188), .A2(n126), .ZN(n128) );
  AND2_X1 U106 ( .A1(n125), .A2(n124), .ZN(n126) );
  OR2_X1 U107 ( .A1(n211), .A2(b[1]), .ZN(n124) );
  OR2_X1 U108 ( .A1(n202), .A2(a[1]), .ZN(n125) );
  AND2_X1 U109 ( .A1(n122), .A2(n121), .ZN(n123) );
  OR2_X1 U110 ( .A1(n187), .A2(d[1]), .ZN(n121) );
  OR2_X1 U111 ( .A1(n178), .A2(c[1]), .ZN(n122) );
  OR2_X1 U112 ( .A1(n120), .A2(n210), .ZN(y[0]) );
  OR2_X1 U113 ( .A1(n118), .A2(n186), .ZN(n119) );
  AND2_X1 U114 ( .A1(n186), .A2(n118), .ZN(n120) );
  AND2_X1 U115 ( .A1(n117), .A2(n116), .ZN(n118) );
  OR2_X1 U116 ( .A1(n209), .A2(b[0]), .ZN(n116) );
  OR2_X1 U117 ( .A1(n201), .A2(a[0]), .ZN(n117) );
  AND2_X1 U118 ( .A1(n114), .A2(n113), .ZN(n115) );
  OR2_X1 U119 ( .A1(n185), .A2(d[0]), .ZN(n113) );
  OR2_X1 U120 ( .A1(n177), .A2(c[0]), .ZN(n114) );
endmodule


module mixCol_1 ( in, out );
  input [31:0] in;
  //input_done

  output [31:0] out;
  //output_done

  wire   [7:0] b0_s2;
  wire   [7:0] b1_s2;
  wire   [7:0] b2_s2;
  wire   [7:0] b3_s2;
  wire   [7:0] b0_s3;
  wire   [7:0] b1_s3;
  wire   [7:0] b2_s3;
  wire   [7:0] b3_s3;
  //wire_done

  scale2_4 b0_scale2 ( .in(in[31:24]), .out(b0_s2) );
  scale2_3 b1_scale2 ( .in(in[23:16]), .out(b1_s2) );
  scale2_2 b2_scale2 ( .in(in[15:8]), .out(b2_s2) );
  scale2_1 b3_scale2 ( .in(in[7:0]), .out(b3_s2) );
  byteXor_5 b0_scale3 ( .a(in[31:24]), .b(b0_s2), .y(b0_s3) );
  byteXor_4 b1_scale3 ( .a(in[23:16]), .b(b1_s2), .y(b1_s3) );
  byteXor_3 b2_scale3 ( .a(in[15:8]), .b(b2_s2), .y(b2_s3) );
  byteXor_2 b3_scale3 ( .a(in[7:0]), .b(b3_s2), .y(b3_s3) );
  byteXor4_4 out0 ( .a(b0_s2), .b(b1_s3), .c(in[15:8]), .d(in[7:0]), .y(
        out[31:24]) );
  byteXor4_3 out1 ( .a(in[31:24]), .b(b1_s2), .c(b2_s3), .d(in[7:0]), .y(
        out[23:16]) );
  byteXor4_2 out2 ( .a(in[31:24]), .b(in[23:16]), .c(b2_s2), .d(b3_s3), .y(
        out[15:8]) );
  byteXor4_1 out3 ( .a(b0_s3), .b(in[23:16]), .c(in[15:8]), .d(b3_s2), .y(
        out[7:0]) );
endmodule


module scale2_5 ( in, out );
  input [7:0] in;
  //input_done

  output [7:0] out;
  //output_done

  wire   in_0, \in[6] , \in[5] , \in[4] , \in[1] , \in[7] , n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20;
  //wire_done

  assign in_0 = in[0];
  assign out[7] = \in[6] ;
  assign \in[6]  = in[6];
  assign out[6] = \in[5] ;
  assign \in[5]  = in[5];
  assign out[5] = \in[4] ;
  assign \in[4]  = in[4];
  assign out[2] = \in[1] ;
  assign \in[1]  = in[1];
  assign out[0] = \in[7] ;
  assign \in[7]  = in[7];

  INV_X1 U1 ( .A(\in[7]), .ZN(n20) );
  INV_X1 U2 ( .A(in[3]), .ZN(n19) );
  INV_X1 U3 ( .A(in[2]), .ZN(n18) );
  INV_X1 U4 ( .A(in_0), .ZN(n17) );
  OR2_X1 U5 ( .A1(n16), .A2(n15), .ZN(out[4]) );
  AND2_X1 U6 ( .A1(in[3]), .A2(n20), .ZN(n15) );
  AND2_X1 U7 ( .A1(\in[7]), .A2(n19), .ZN(n16) );
  OR2_X1 U8 ( .A1(n14), .A2(n13), .ZN(out[3]) );
  AND2_X1 U9 ( .A1(in[2]), .A2(n20), .ZN(n13) );
  AND2_X1 U10 ( .A1(\in[7]), .A2(n18), .ZN(n14) );
  OR2_X1 U11 ( .A1(n12), .A2(n11), .ZN(out[1]) );
  AND2_X1 U12 ( .A1(in_0), .A2(n20), .ZN(n11) );
  AND2_X1 U13 ( .A1(\in[7]), .A2(n17), .ZN(n12) );
endmodule


module scale2_6 ( in, out );
  input [7:0] in;
  //input_done

  output [7:0] out;
  //output_done

  wire   in_0, \in[6] , \in[5] , \in[4] , \in[1] , \in[7] , n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20;
  //wire_done

  assign in_0 = in[0];
  assign out[7] = \in[6] ;
  assign \in[6]  = in[6];
  assign out[6] = \in[5] ;
  assign \in[5]  = in[5];
  assign out[5] = \in[4] ;
  assign \in[4]  = in[4];
  assign out[2] = \in[1] ;
  assign \in[1]  = in[1];
  assign out[0] = \in[7] ;
  assign \in[7]  = in[7];

  INV_X1 U1 ( .A(\in[7]), .ZN(n20) );
  INV_X1 U2 ( .A(in[3]), .ZN(n19) );
  INV_X1 U3 ( .A(in[2]), .ZN(n18) );
  INV_X1 U4 ( .A(in_0), .ZN(n17) );
  OR2_X1 U5 ( .A1(n16), .A2(n15), .ZN(out[4]) );
  AND2_X1 U6 ( .A1(in[3]), .A2(n20), .ZN(n15) );
  AND2_X1 U7 ( .A1(\in[7]), .A2(n19), .ZN(n16) );
  OR2_X1 U8 ( .A1(n14), .A2(n13), .ZN(out[3]) );
  AND2_X1 U9 ( .A1(in[2]), .A2(n20), .ZN(n13) );
  AND2_X1 U10 ( .A1(\in[7]), .A2(n18), .ZN(n14) );
  OR2_X1 U11 ( .A1(n12), .A2(n11), .ZN(out[1]) );
  AND2_X1 U12 ( .A1(in_0), .A2(n20), .ZN(n11) );
  AND2_X1 U13 ( .A1(\in[7]), .A2(n17), .ZN(n12) );
endmodule


module scale2_7 ( in, out );
  input [7:0] in;
  //input_done

  output [7:0] out;
  //output_done

  wire   in_0, \in[6] , \in[5] , \in[4] , \in[1] , \in[7] , n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20;
  //wire_done

  assign in_0 = in[0];
  assign out[7] = \in[6] ;
  assign \in[6]  = in[6];
  assign out[6] = \in[5] ;
  assign \in[5]  = in[5];
  assign out[5] = \in[4] ;
  assign \in[4]  = in[4];
  assign out[2] = \in[1] ;
  assign \in[1]  = in[1];
  assign out[0] = \in[7] ;
  assign \in[7]  = in[7];

  INV_X1 U1 ( .A(\in[7]), .ZN(n20) );
  INV_X1 U2 ( .A(in[3]), .ZN(n19) );
  INV_X1 U3 ( .A(in[2]), .ZN(n18) );
  INV_X1 U4 ( .A(in_0), .ZN(n17) );
  OR2_X1 U5 ( .A1(n16), .A2(n15), .ZN(out[4]) );
  AND2_X1 U6 ( .A1(in[3]), .A2(n20), .ZN(n15) );
  AND2_X1 U7 ( .A1(\in[7]), .A2(n19), .ZN(n16) );
  OR2_X1 U8 ( .A1(n14), .A2(n13), .ZN(out[3]) );
  AND2_X1 U9 ( .A1(in[2]), .A2(n20), .ZN(n13) );
  AND2_X1 U10 ( .A1(\in[7]), .A2(n18), .ZN(n14) );
  OR2_X1 U11 ( .A1(n12), .A2(n11), .ZN(out[1]) );
  AND2_X1 U12 ( .A1(in_0), .A2(n20), .ZN(n11) );
  AND2_X1 U13 ( .A1(\in[7]), .A2(n17), .ZN(n12) );
endmodule


module scale2_8 ( in, out );
  input [7:0] in;
  //input_done

  output [7:0] out;
  //output_done

  wire   in_0, \in[6] , \in[5] , \in[4] , \in[1] , \in[7] , n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20;
  //wire_done

  assign in_0 = in[0];
  assign out[7] = \in[6] ;
  assign \in[6]  = in[6];
  assign out[6] = \in[5] ;
  assign \in[5]  = in[5];
  assign out[5] = \in[4] ;
  assign \in[4]  = in[4];
  assign out[2] = \in[1] ;
  assign \in[1]  = in[1];
  assign out[0] = \in[7] ;
  assign \in[7]  = in[7];

  INV_X1 U1 ( .A(\in[7]), .ZN(n20) );
  INV_X1 U2 ( .A(in[3]), .ZN(n19) );
  INV_X1 U3 ( .A(in[2]), .ZN(n18) );
  INV_X1 U4 ( .A(in_0), .ZN(n17) );
  OR2_X1 U5 ( .A1(n16), .A2(n15), .ZN(out[4]) );
  AND2_X1 U6 ( .A1(in[3]), .A2(n20), .ZN(n15) );
  AND2_X1 U7 ( .A1(\in[7]), .A2(n19), .ZN(n16) );
  OR2_X1 U8 ( .A1(n14), .A2(n13), .ZN(out[3]) );
  AND2_X1 U9 ( .A1(in[2]), .A2(n20), .ZN(n13) );
  AND2_X1 U10 ( .A1(\in[7]), .A2(n18), .ZN(n14) );
  OR2_X1 U11 ( .A1(n12), .A2(n11), .ZN(out[1]) );
  AND2_X1 U12 ( .A1(in_0), .A2(n20), .ZN(n11) );
  AND2_X1 U13 ( .A1(\in[7]), .A2(n17), .ZN(n12) );
endmodule


module byteXor_6 ( a, b, y );
  input [7:0] a;
  input [7:0] b;
  //input_done

  output [7:0] y;
  //output_done

  wire   n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64;
  //wire_done

  INV_X1 U1 ( .A(n47), .ZN(n64) );
  INV_X1 U2 ( .A(a[7]), .ZN(n63) );
  INV_X1 U3 ( .A(n45), .ZN(n62) );
  INV_X1 U4 ( .A(a[6]), .ZN(n61) );
  INV_X1 U5 ( .A(n43), .ZN(n60) );
  INV_X1 U6 ( .A(a[5]), .ZN(n59) );
  INV_X1 U7 ( .A(n41), .ZN(n58) );
  INV_X1 U8 ( .A(a[4]), .ZN(n57) );
  INV_X1 U9 ( .A(n39), .ZN(n56) );
  INV_X1 U10 ( .A(a[3]), .ZN(n55) );
  INV_X1 U11 ( .A(n37), .ZN(n54) );
  INV_X1 U12 ( .A(a[2]), .ZN(n53) );
  INV_X1 U13 ( .A(n35), .ZN(n52) );
  INV_X1 U14 ( .A(a[1]), .ZN(n51) );
  INV_X1 U15 ( .A(n33), .ZN(n50) );
  INV_X1 U16 ( .A(a[0]), .ZN(n49) );
  OR2_X1 U17 ( .A1(n48), .A2(n64), .ZN(y[7]) );
  OR2_X1 U18 ( .A1(n63), .A2(b[7]), .ZN(n47) );
  AND2_X1 U19 ( .A1(b[7]), .A2(n63), .ZN(n48) );
  OR2_X1 U20 ( .A1(n46), .A2(n62), .ZN(y[6]) );
  OR2_X1 U21 ( .A1(n61), .A2(b[6]), .ZN(n45) );
  AND2_X1 U22 ( .A1(b[6]), .A2(n61), .ZN(n46) );
  OR2_X1 U23 ( .A1(n44), .A2(n60), .ZN(y[5]) );
  OR2_X1 U24 ( .A1(n59), .A2(b[5]), .ZN(n43) );
  AND2_X1 U25 ( .A1(b[5]), .A2(n59), .ZN(n44) );
  OR2_X1 U26 ( .A1(n42), .A2(n58), .ZN(y[4]) );
  OR2_X1 U27 ( .A1(n57), .A2(b[4]), .ZN(n41) );
  AND2_X1 U28 ( .A1(b[4]), .A2(n57), .ZN(n42) );
  OR2_X1 U29 ( .A1(n40), .A2(n56), .ZN(y[3]) );
  OR2_X1 U30 ( .A1(n55), .A2(b[3]), .ZN(n39) );
  AND2_X1 U31 ( .A1(b[3]), .A2(n55), .ZN(n40) );
  OR2_X1 U32 ( .A1(n38), .A2(n54), .ZN(y[2]) );
  OR2_X1 U33 ( .A1(n53), .A2(b[2]), .ZN(n37) );
  AND2_X1 U34 ( .A1(b[2]), .A2(n53), .ZN(n38) );
  OR2_X1 U35 ( .A1(n36), .A2(n52), .ZN(y[1]) );
  OR2_X1 U36 ( .A1(n51), .A2(b[1]), .ZN(n35) );
  AND2_X1 U37 ( .A1(b[1]), .A2(n51), .ZN(n36) );
  OR2_X1 U38 ( .A1(n34), .A2(n50), .ZN(y[0]) );
  OR2_X1 U39 ( .A1(n49), .A2(b[0]), .ZN(n33) );
  AND2_X1 U40 ( .A1(b[0]), .A2(n49), .ZN(n34) );
endmodule


module byteXor_7 ( a, b, y );
  input [7:0] a;
  input [7:0] b;
  //input_done

  output [7:0] y;
  //output_done

  wire   n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64;
  //wire_done

  INV_X1 U1 ( .A(n47), .ZN(n64) );
  INV_X1 U2 ( .A(a[7]), .ZN(n63) );
  INV_X1 U3 ( .A(n45), .ZN(n62) );
  INV_X1 U4 ( .A(a[6]), .ZN(n61) );
  INV_X1 U5 ( .A(n43), .ZN(n60) );
  INV_X1 U6 ( .A(a[5]), .ZN(n59) );
  INV_X1 U7 ( .A(n41), .ZN(n58) );
  INV_X1 U8 ( .A(a[4]), .ZN(n57) );
  INV_X1 U9 ( .A(n39), .ZN(n56) );
  INV_X1 U10 ( .A(a[3]), .ZN(n55) );
  INV_X1 U11 ( .A(n37), .ZN(n54) );
  INV_X1 U12 ( .A(a[2]), .ZN(n53) );
  INV_X1 U13 ( .A(n35), .ZN(n52) );
  INV_X1 U14 ( .A(a[1]), .ZN(n51) );
  INV_X1 U15 ( .A(n33), .ZN(n50) );
  INV_X1 U16 ( .A(a[0]), .ZN(n49) );
  OR2_X1 U17 ( .A1(n48), .A2(n64), .ZN(y[7]) );
  OR2_X1 U18 ( .A1(n63), .A2(b[7]), .ZN(n47) );
  AND2_X1 U19 ( .A1(b[7]), .A2(n63), .ZN(n48) );
  OR2_X1 U20 ( .A1(n46), .A2(n62), .ZN(y[6]) );
  OR2_X1 U21 ( .A1(n61), .A2(b[6]), .ZN(n45) );
  AND2_X1 U22 ( .A1(b[6]), .A2(n61), .ZN(n46) );
  OR2_X1 U23 ( .A1(n44), .A2(n60), .ZN(y[5]) );
  OR2_X1 U24 ( .A1(n59), .A2(b[5]), .ZN(n43) );
  AND2_X1 U25 ( .A1(b[5]), .A2(n59), .ZN(n44) );
  OR2_X1 U26 ( .A1(n42), .A2(n58), .ZN(y[4]) );
  OR2_X1 U27 ( .A1(n57), .A2(b[4]), .ZN(n41) );
  AND2_X1 U28 ( .A1(b[4]), .A2(n57), .ZN(n42) );
  OR2_X1 U29 ( .A1(n40), .A2(n56), .ZN(y[3]) );
  OR2_X1 U30 ( .A1(n55), .A2(b[3]), .ZN(n39) );
  AND2_X1 U31 ( .A1(b[3]), .A2(n55), .ZN(n40) );
  OR2_X1 U32 ( .A1(n38), .A2(n54), .ZN(y[2]) );
  OR2_X1 U33 ( .A1(n53), .A2(b[2]), .ZN(n37) );
  AND2_X1 U34 ( .A1(b[2]), .A2(n53), .ZN(n38) );
  OR2_X1 U35 ( .A1(n36), .A2(n52), .ZN(y[1]) );
  OR2_X1 U36 ( .A1(n51), .A2(b[1]), .ZN(n35) );
  AND2_X1 U37 ( .A1(b[1]), .A2(n51), .ZN(n36) );
  OR2_X1 U38 ( .A1(n34), .A2(n50), .ZN(y[0]) );
  OR2_X1 U39 ( .A1(n49), .A2(b[0]), .ZN(n33) );
  AND2_X1 U40 ( .A1(b[0]), .A2(n49), .ZN(n34) );
endmodule


module byteXor_8 ( a, b, y );
  input [7:0] a;
  input [7:0] b;
  //input_done

  output [7:0] y;
  //output_done

  wire   n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64;
  //wire_done

  INV_X1 U1 ( .A(n47), .ZN(n64) );
  INV_X1 U2 ( .A(a[7]), .ZN(n63) );
  INV_X1 U3 ( .A(n45), .ZN(n62) );
  INV_X1 U4 ( .A(a[6]), .ZN(n61) );
  INV_X1 U5 ( .A(n43), .ZN(n60) );
  INV_X1 U6 ( .A(a[5]), .ZN(n59) );
  INV_X1 U7 ( .A(n41), .ZN(n58) );
  INV_X1 U8 ( .A(a[4]), .ZN(n57) );
  INV_X1 U9 ( .A(n39), .ZN(n56) );
  INV_X1 U10 ( .A(a[3]), .ZN(n55) );
  INV_X1 U11 ( .A(n37), .ZN(n54) );
  INV_X1 U12 ( .A(a[2]), .ZN(n53) );
  INV_X1 U13 ( .A(n35), .ZN(n52) );
  INV_X1 U14 ( .A(a[1]), .ZN(n51) );
  INV_X1 U15 ( .A(n33), .ZN(n50) );
  INV_X1 U16 ( .A(a[0]), .ZN(n49) );
  OR2_X1 U17 ( .A1(n48), .A2(n64), .ZN(y[7]) );
  OR2_X1 U18 ( .A1(n63), .A2(b[7]), .ZN(n47) );
  AND2_X1 U19 ( .A1(b[7]), .A2(n63), .ZN(n48) );
  OR2_X1 U20 ( .A1(n46), .A2(n62), .ZN(y[6]) );
  OR2_X1 U21 ( .A1(n61), .A2(b[6]), .ZN(n45) );
  AND2_X1 U22 ( .A1(b[6]), .A2(n61), .ZN(n46) );
  OR2_X1 U23 ( .A1(n44), .A2(n60), .ZN(y[5]) );
  OR2_X1 U24 ( .A1(n59), .A2(b[5]), .ZN(n43) );
  AND2_X1 U25 ( .A1(b[5]), .A2(n59), .ZN(n44) );
  OR2_X1 U26 ( .A1(n42), .A2(n58), .ZN(y[4]) );
  OR2_X1 U27 ( .A1(n57), .A2(b[4]), .ZN(n41) );
  AND2_X1 U28 ( .A1(b[4]), .A2(n57), .ZN(n42) );
  OR2_X1 U29 ( .A1(n40), .A2(n56), .ZN(y[3]) );
  OR2_X1 U30 ( .A1(n55), .A2(b[3]), .ZN(n39) );
  AND2_X1 U31 ( .A1(b[3]), .A2(n55), .ZN(n40) );
  OR2_X1 U32 ( .A1(n38), .A2(n54), .ZN(y[2]) );
  OR2_X1 U33 ( .A1(n53), .A2(b[2]), .ZN(n37) );
  AND2_X1 U34 ( .A1(b[2]), .A2(n53), .ZN(n38) );
  OR2_X1 U35 ( .A1(n36), .A2(n52), .ZN(y[1]) );
  OR2_X1 U36 ( .A1(n51), .A2(b[1]), .ZN(n35) );
  AND2_X1 U37 ( .A1(b[1]), .A2(n51), .ZN(n36) );
  OR2_X1 U38 ( .A1(n34), .A2(n50), .ZN(y[0]) );
  OR2_X1 U39 ( .A1(n49), .A2(b[0]), .ZN(n33) );
  AND2_X1 U40 ( .A1(b[0]), .A2(n49), .ZN(n34) );
endmodule


module byteXor_9 ( a, b, y );
  input [7:0] a;
  input [7:0] b;
  //input_done

  output [7:0] y;
  //output_done

  wire   n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64;
  //wire_done

  INV_X1 U1 ( .A(n47), .ZN(n64) );
  INV_X1 U2 ( .A(a[7]), .ZN(n63) );
  INV_X1 U3 ( .A(n45), .ZN(n62) );
  INV_X1 U4 ( .A(a[6]), .ZN(n61) );
  INV_X1 U5 ( .A(n43), .ZN(n60) );
  INV_X1 U6 ( .A(a[5]), .ZN(n59) );
  INV_X1 U7 ( .A(n41), .ZN(n58) );
  INV_X1 U8 ( .A(a[4]), .ZN(n57) );
  INV_X1 U9 ( .A(n39), .ZN(n56) );
  INV_X1 U10 ( .A(a[3]), .ZN(n55) );
  INV_X1 U11 ( .A(n37), .ZN(n54) );
  INV_X1 U12 ( .A(a[2]), .ZN(n53) );
  INV_X1 U13 ( .A(n35), .ZN(n52) );
  INV_X1 U14 ( .A(a[1]), .ZN(n51) );
  INV_X1 U15 ( .A(n33), .ZN(n50) );
  INV_X1 U16 ( .A(a[0]), .ZN(n49) );
  OR2_X1 U17 ( .A1(n48), .A2(n64), .ZN(y[7]) );
  OR2_X1 U18 ( .A1(n63), .A2(b[7]), .ZN(n47) );
  AND2_X1 U19 ( .A1(b[7]), .A2(n63), .ZN(n48) );
  OR2_X1 U20 ( .A1(n46), .A2(n62), .ZN(y[6]) );
  OR2_X1 U21 ( .A1(n61), .A2(b[6]), .ZN(n45) );
  AND2_X1 U22 ( .A1(b[6]), .A2(n61), .ZN(n46) );
  OR2_X1 U23 ( .A1(n44), .A2(n60), .ZN(y[5]) );
  OR2_X1 U24 ( .A1(n59), .A2(b[5]), .ZN(n43) );
  AND2_X1 U25 ( .A1(b[5]), .A2(n59), .ZN(n44) );
  OR2_X1 U26 ( .A1(n42), .A2(n58), .ZN(y[4]) );
  OR2_X1 U27 ( .A1(n57), .A2(b[4]), .ZN(n41) );
  AND2_X1 U28 ( .A1(b[4]), .A2(n57), .ZN(n42) );
  OR2_X1 U29 ( .A1(n40), .A2(n56), .ZN(y[3]) );
  OR2_X1 U30 ( .A1(n55), .A2(b[3]), .ZN(n39) );
  AND2_X1 U31 ( .A1(b[3]), .A2(n55), .ZN(n40) );
  OR2_X1 U32 ( .A1(n38), .A2(n54), .ZN(y[2]) );
  OR2_X1 U33 ( .A1(n53), .A2(b[2]), .ZN(n37) );
  AND2_X1 U34 ( .A1(b[2]), .A2(n53), .ZN(n38) );
  OR2_X1 U35 ( .A1(n36), .A2(n52), .ZN(y[1]) );
  OR2_X1 U36 ( .A1(n51), .A2(b[1]), .ZN(n35) );
  AND2_X1 U37 ( .A1(b[1]), .A2(n51), .ZN(n36) );
  OR2_X1 U38 ( .A1(n34), .A2(n50), .ZN(y[0]) );
  OR2_X1 U39 ( .A1(n49), .A2(b[0]), .ZN(n33) );
  AND2_X1 U40 ( .A1(b[0]), .A2(n49), .ZN(n34) );
endmodule


module byteXor4_5 ( a, b, c, d, y );
  input [7:0] a;
  input [7:0] b;
  input [7:0] c;
  input [7:0] d;
  //input_done

  output [7:0] y;
  //output_done

  wire   n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224;
  //wire_done

  INV_X1 U1 ( .A(n175), .ZN(n224) );
  INV_X1 U2 ( .A(a[7]), .ZN(n223) );
  INV_X1 U3 ( .A(n167), .ZN(n222) );
  INV_X1 U4 ( .A(a[6]), .ZN(n221) );
  INV_X1 U5 ( .A(n159), .ZN(n220) );
  INV_X1 U6 ( .A(a[5]), .ZN(n219) );
  INV_X1 U7 ( .A(n151), .ZN(n218) );
  INV_X1 U8 ( .A(a[4]), .ZN(n217) );
  INV_X1 U9 ( .A(n143), .ZN(n216) );
  INV_X1 U10 ( .A(a[3]), .ZN(n215) );
  INV_X1 U11 ( .A(n135), .ZN(n214) );
  INV_X1 U12 ( .A(a[2]), .ZN(n213) );
  INV_X1 U13 ( .A(n127), .ZN(n212) );
  INV_X1 U14 ( .A(a[1]), .ZN(n211) );
  INV_X1 U15 ( .A(n119), .ZN(n210) );
  INV_X1 U16 ( .A(a[0]), .ZN(n209) );
  INV_X1 U17 ( .A(b[7]), .ZN(n208) );
  INV_X1 U18 ( .A(b[6]), .ZN(n207) );
  INV_X1 U19 ( .A(b[5]), .ZN(n206) );
  INV_X1 U20 ( .A(b[4]), .ZN(n205) );
  INV_X1 U21 ( .A(b[3]), .ZN(n204) );
  INV_X1 U22 ( .A(b[2]), .ZN(n203) );
  INV_X1 U23 ( .A(b[1]), .ZN(n202) );
  INV_X1 U24 ( .A(b[0]), .ZN(n201) );
  INV_X1 U25 ( .A(n171), .ZN(n200) );
  INV_X1 U26 ( .A(c[7]), .ZN(n199) );
  INV_X1 U27 ( .A(n163), .ZN(n198) );
  INV_X1 U28 ( .A(c[6]), .ZN(n197) );
  INV_X1 U29 ( .A(n155), .ZN(n196) );
  INV_X1 U30 ( .A(c[5]), .ZN(n195) );
  INV_X1 U31 ( .A(n147), .ZN(n194) );
  INV_X1 U32 ( .A(c[4]), .ZN(n193) );
  INV_X1 U33 ( .A(n139), .ZN(n192) );
  INV_X1 U34 ( .A(c[3]), .ZN(n191) );
  INV_X1 U35 ( .A(n131), .ZN(n190) );
  INV_X1 U36 ( .A(c[2]), .ZN(n189) );
  INV_X1 U37 ( .A(n123), .ZN(n188) );
  INV_X1 U38 ( .A(c[1]), .ZN(n187) );
  INV_X1 U39 ( .A(n115), .ZN(n186) );
  INV_X1 U40 ( .A(c[0]), .ZN(n185) );
  INV_X1 U41 ( .A(d[7]), .ZN(n184) );
  INV_X1 U42 ( .A(d[6]), .ZN(n183) );
  INV_X1 U43 ( .A(d[5]), .ZN(n182) );
  INV_X1 U44 ( .A(d[4]), .ZN(n181) );
  INV_X1 U45 ( .A(d[3]), .ZN(n180) );
  INV_X1 U46 ( .A(d[2]), .ZN(n179) );
  INV_X1 U47 ( .A(d[1]), .ZN(n178) );
  INV_X1 U48 ( .A(d[0]), .ZN(n177) );
  OR2_X1 U49 ( .A1(n176), .A2(n224), .ZN(y[7]) );
  OR2_X1 U50 ( .A1(n174), .A2(n200), .ZN(n175) );
  AND2_X1 U51 ( .A1(n200), .A2(n174), .ZN(n176) );
  AND2_X1 U52 ( .A1(n173), .A2(n172), .ZN(n174) );
  OR2_X1 U53 ( .A1(n223), .A2(b[7]), .ZN(n172) );
  OR2_X1 U54 ( .A1(n208), .A2(a[7]), .ZN(n173) );
  AND2_X1 U55 ( .A1(n170), .A2(n169), .ZN(n171) );
  OR2_X1 U56 ( .A1(n199), .A2(d[7]), .ZN(n169) );
  OR2_X1 U57 ( .A1(n184), .A2(c[7]), .ZN(n170) );
  OR2_X1 U58 ( .A1(n168), .A2(n222), .ZN(y[6]) );
  OR2_X1 U59 ( .A1(n166), .A2(n198), .ZN(n167) );
  AND2_X1 U60 ( .A1(n198), .A2(n166), .ZN(n168) );
  AND2_X1 U61 ( .A1(n165), .A2(n164), .ZN(n166) );
  OR2_X1 U62 ( .A1(n221), .A2(b[6]), .ZN(n164) );
  OR2_X1 U63 ( .A1(n207), .A2(a[6]), .ZN(n165) );
  AND2_X1 U64 ( .A1(n162), .A2(n161), .ZN(n163) );
  OR2_X1 U65 ( .A1(n197), .A2(d[6]), .ZN(n161) );
  OR2_X1 U66 ( .A1(n183), .A2(c[6]), .ZN(n162) );
  OR2_X1 U67 ( .A1(n160), .A2(n220), .ZN(y[5]) );
  OR2_X1 U68 ( .A1(n158), .A2(n196), .ZN(n159) );
  AND2_X1 U69 ( .A1(n196), .A2(n158), .ZN(n160) );
  AND2_X1 U70 ( .A1(n157), .A2(n156), .ZN(n158) );
  OR2_X1 U71 ( .A1(n219), .A2(b[5]), .ZN(n156) );
  OR2_X1 U72 ( .A1(n206), .A2(a[5]), .ZN(n157) );
  AND2_X1 U73 ( .A1(n154), .A2(n153), .ZN(n155) );
  OR2_X1 U74 ( .A1(n195), .A2(d[5]), .ZN(n153) );
  OR2_X1 U75 ( .A1(n182), .A2(c[5]), .ZN(n154) );
  OR2_X1 U76 ( .A1(n152), .A2(n218), .ZN(y[4]) );
  OR2_X1 U77 ( .A1(n150), .A2(n194), .ZN(n151) );
  AND2_X1 U78 ( .A1(n194), .A2(n150), .ZN(n152) );
  AND2_X1 U79 ( .A1(n149), .A2(n148), .ZN(n150) );
  OR2_X1 U80 ( .A1(n217), .A2(b[4]), .ZN(n148) );
  OR2_X1 U81 ( .A1(n205), .A2(a[4]), .ZN(n149) );
  AND2_X1 U82 ( .A1(n146), .A2(n145), .ZN(n147) );
  OR2_X1 U83 ( .A1(n193), .A2(d[4]), .ZN(n145) );
  OR2_X1 U84 ( .A1(n181), .A2(c[4]), .ZN(n146) );
  OR2_X1 U85 ( .A1(n144), .A2(n216), .ZN(y[3]) );
  OR2_X1 U86 ( .A1(n142), .A2(n192), .ZN(n143) );
  AND2_X1 U87 ( .A1(n192), .A2(n142), .ZN(n144) );
  AND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(n142) );
  OR2_X1 U89 ( .A1(n215), .A2(b[3]), .ZN(n140) );
  OR2_X1 U90 ( .A1(n204), .A2(a[3]), .ZN(n141) );
  AND2_X1 U91 ( .A1(n138), .A2(n137), .ZN(n139) );
  OR2_X1 U92 ( .A1(n191), .A2(d[3]), .ZN(n137) );
  OR2_X1 U93 ( .A1(n180), .A2(c[3]), .ZN(n138) );
  OR2_X1 U94 ( .A1(n136), .A2(n214), .ZN(y[2]) );
  OR2_X1 U95 ( .A1(n134), .A2(n190), .ZN(n135) );
  AND2_X1 U96 ( .A1(n190), .A2(n134), .ZN(n136) );
  AND2_X1 U97 ( .A1(n133), .A2(n132), .ZN(n134) );
  OR2_X1 U98 ( .A1(n213), .A2(b[2]), .ZN(n132) );
  OR2_X1 U99 ( .A1(n203), .A2(a[2]), .ZN(n133) );
  AND2_X1 U100 ( .A1(n130), .A2(n129), .ZN(n131) );
  OR2_X1 U101 ( .A1(n189), .A2(d[2]), .ZN(n129) );
  OR2_X1 U102 ( .A1(n179), .A2(c[2]), .ZN(n130) );
  OR2_X1 U103 ( .A1(n128), .A2(n212), .ZN(y[1]) );
  OR2_X1 U104 ( .A1(n126), .A2(n188), .ZN(n127) );
  AND2_X1 U105 ( .A1(n188), .A2(n126), .ZN(n128) );
  AND2_X1 U106 ( .A1(n125), .A2(n124), .ZN(n126) );
  OR2_X1 U107 ( .A1(n211), .A2(b[1]), .ZN(n124) );
  OR2_X1 U108 ( .A1(n202), .A2(a[1]), .ZN(n125) );
  AND2_X1 U109 ( .A1(n122), .A2(n121), .ZN(n123) );
  OR2_X1 U110 ( .A1(n187), .A2(d[1]), .ZN(n121) );
  OR2_X1 U111 ( .A1(n178), .A2(c[1]), .ZN(n122) );
  OR2_X1 U112 ( .A1(n120), .A2(n210), .ZN(y[0]) );
  OR2_X1 U113 ( .A1(n118), .A2(n186), .ZN(n119) );
  AND2_X1 U114 ( .A1(n186), .A2(n118), .ZN(n120) );
  AND2_X1 U115 ( .A1(n117), .A2(n116), .ZN(n118) );
  OR2_X1 U116 ( .A1(n209), .A2(b[0]), .ZN(n116) );
  OR2_X1 U117 ( .A1(n201), .A2(a[0]), .ZN(n117) );
  AND2_X1 U118 ( .A1(n114), .A2(n113), .ZN(n115) );
  OR2_X1 U119 ( .A1(n185), .A2(d[0]), .ZN(n113) );
  OR2_X1 U120 ( .A1(n177), .A2(c[0]), .ZN(n114) );
endmodule


module byteXor4_6 ( a, b, c, d, y );
  input [7:0] a;
  input [7:0] b;
  input [7:0] c;
  input [7:0] d;
  //input_done

  output [7:0] y;
  //output_done

  wire   n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224;
  //wire_done

  INV_X1 U1 ( .A(n175), .ZN(n224) );
  INV_X1 U2 ( .A(a[7]), .ZN(n223) );
  INV_X1 U3 ( .A(n167), .ZN(n222) );
  INV_X1 U4 ( .A(a[6]), .ZN(n221) );
  INV_X1 U5 ( .A(n159), .ZN(n220) );
  INV_X1 U6 ( .A(a[5]), .ZN(n219) );
  INV_X1 U7 ( .A(n151), .ZN(n218) );
  INV_X1 U8 ( .A(a[4]), .ZN(n217) );
  INV_X1 U9 ( .A(n143), .ZN(n216) );
  INV_X1 U10 ( .A(a[3]), .ZN(n215) );
  INV_X1 U11 ( .A(n135), .ZN(n214) );
  INV_X1 U12 ( .A(a[2]), .ZN(n213) );
  INV_X1 U13 ( .A(n127), .ZN(n212) );
  INV_X1 U14 ( .A(a[1]), .ZN(n211) );
  INV_X1 U15 ( .A(n119), .ZN(n210) );
  INV_X1 U16 ( .A(a[0]), .ZN(n209) );
  INV_X1 U17 ( .A(b[7]), .ZN(n208) );
  INV_X1 U18 ( .A(b[6]), .ZN(n207) );
  INV_X1 U19 ( .A(b[5]), .ZN(n206) );
  INV_X1 U20 ( .A(b[4]), .ZN(n205) );
  INV_X1 U21 ( .A(b[3]), .ZN(n204) );
  INV_X1 U22 ( .A(b[2]), .ZN(n203) );
  INV_X1 U23 ( .A(b[1]), .ZN(n202) );
  INV_X1 U24 ( .A(b[0]), .ZN(n201) );
  INV_X1 U25 ( .A(n171), .ZN(n200) );
  INV_X1 U26 ( .A(c[7]), .ZN(n199) );
  INV_X1 U27 ( .A(n163), .ZN(n198) );
  INV_X1 U28 ( .A(c[6]), .ZN(n197) );
  INV_X1 U29 ( .A(n155), .ZN(n196) );
  INV_X1 U30 ( .A(c[5]), .ZN(n195) );
  INV_X1 U31 ( .A(n147), .ZN(n194) );
  INV_X1 U32 ( .A(c[4]), .ZN(n193) );
  INV_X1 U33 ( .A(n139), .ZN(n192) );
  INV_X1 U34 ( .A(c[3]), .ZN(n191) );
  INV_X1 U35 ( .A(n131), .ZN(n190) );
  INV_X1 U36 ( .A(c[2]), .ZN(n189) );
  INV_X1 U37 ( .A(n123), .ZN(n188) );
  INV_X1 U38 ( .A(c[1]), .ZN(n187) );
  INV_X1 U39 ( .A(n115), .ZN(n186) );
  INV_X1 U40 ( .A(c[0]), .ZN(n185) );
  INV_X1 U41 ( .A(d[7]), .ZN(n184) );
  INV_X1 U42 ( .A(d[6]), .ZN(n183) );
  INV_X1 U43 ( .A(d[5]), .ZN(n182) );
  INV_X1 U44 ( .A(d[4]), .ZN(n181) );
  INV_X1 U45 ( .A(d[3]), .ZN(n180) );
  INV_X1 U46 ( .A(d[2]), .ZN(n179) );
  INV_X1 U47 ( .A(d[1]), .ZN(n178) );
  INV_X1 U48 ( .A(d[0]), .ZN(n177) );
  OR2_X1 U49 ( .A1(n176), .A2(n224), .ZN(y[7]) );
  OR2_X1 U50 ( .A1(n174), .A2(n200), .ZN(n175) );
  AND2_X1 U51 ( .A1(n200), .A2(n174), .ZN(n176) );
  AND2_X1 U52 ( .A1(n173), .A2(n172), .ZN(n174) );
  OR2_X1 U53 ( .A1(n223), .A2(b[7]), .ZN(n172) );
  OR2_X1 U54 ( .A1(n208), .A2(a[7]), .ZN(n173) );
  AND2_X1 U55 ( .A1(n170), .A2(n169), .ZN(n171) );
  OR2_X1 U56 ( .A1(n199), .A2(d[7]), .ZN(n169) );
  OR2_X1 U57 ( .A1(n184), .A2(c[7]), .ZN(n170) );
  OR2_X1 U58 ( .A1(n168), .A2(n222), .ZN(y[6]) );
  OR2_X1 U59 ( .A1(n166), .A2(n198), .ZN(n167) );
  AND2_X1 U60 ( .A1(n198), .A2(n166), .ZN(n168) );
  AND2_X1 U61 ( .A1(n165), .A2(n164), .ZN(n166) );
  OR2_X1 U62 ( .A1(n221), .A2(b[6]), .ZN(n164) );
  OR2_X1 U63 ( .A1(n207), .A2(a[6]), .ZN(n165) );
  AND2_X1 U64 ( .A1(n162), .A2(n161), .ZN(n163) );
  OR2_X1 U65 ( .A1(n197), .A2(d[6]), .ZN(n161) );
  OR2_X1 U66 ( .A1(n183), .A2(c[6]), .ZN(n162) );
  OR2_X1 U67 ( .A1(n160), .A2(n220), .ZN(y[5]) );
  OR2_X1 U68 ( .A1(n158), .A2(n196), .ZN(n159) );
  AND2_X1 U69 ( .A1(n196), .A2(n158), .ZN(n160) );
  AND2_X1 U70 ( .A1(n157), .A2(n156), .ZN(n158) );
  OR2_X1 U71 ( .A1(n219), .A2(b[5]), .ZN(n156) );
  OR2_X1 U72 ( .A1(n206), .A2(a[5]), .ZN(n157) );
  AND2_X1 U73 ( .A1(n154), .A2(n153), .ZN(n155) );
  OR2_X1 U74 ( .A1(n195), .A2(d[5]), .ZN(n153) );
  OR2_X1 U75 ( .A1(n182), .A2(c[5]), .ZN(n154) );
  OR2_X1 U76 ( .A1(n152), .A2(n218), .ZN(y[4]) );
  OR2_X1 U77 ( .A1(n150), .A2(n194), .ZN(n151) );
  AND2_X1 U78 ( .A1(n194), .A2(n150), .ZN(n152) );
  AND2_X1 U79 ( .A1(n149), .A2(n148), .ZN(n150) );
  OR2_X1 U80 ( .A1(n217), .A2(b[4]), .ZN(n148) );
  OR2_X1 U81 ( .A1(n205), .A2(a[4]), .ZN(n149) );
  AND2_X1 U82 ( .A1(n146), .A2(n145), .ZN(n147) );
  OR2_X1 U83 ( .A1(n193), .A2(d[4]), .ZN(n145) );
  OR2_X1 U84 ( .A1(n181), .A2(c[4]), .ZN(n146) );
  OR2_X1 U85 ( .A1(n144), .A2(n216), .ZN(y[3]) );
  OR2_X1 U86 ( .A1(n142), .A2(n192), .ZN(n143) );
  AND2_X1 U87 ( .A1(n192), .A2(n142), .ZN(n144) );
  AND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(n142) );
  OR2_X1 U89 ( .A1(n215), .A2(b[3]), .ZN(n140) );
  OR2_X1 U90 ( .A1(n204), .A2(a[3]), .ZN(n141) );
  AND2_X1 U91 ( .A1(n138), .A2(n137), .ZN(n139) );
  OR2_X1 U92 ( .A1(n191), .A2(d[3]), .ZN(n137) );
  OR2_X1 U93 ( .A1(n180), .A2(c[3]), .ZN(n138) );
  OR2_X1 U94 ( .A1(n136), .A2(n214), .ZN(y[2]) );
  OR2_X1 U95 ( .A1(n134), .A2(n190), .ZN(n135) );
  AND2_X1 U96 ( .A1(n190), .A2(n134), .ZN(n136) );
  AND2_X1 U97 ( .A1(n133), .A2(n132), .ZN(n134) );
  OR2_X1 U98 ( .A1(n213), .A2(b[2]), .ZN(n132) );
  OR2_X1 U99 ( .A1(n203), .A2(a[2]), .ZN(n133) );
  AND2_X1 U100 ( .A1(n130), .A2(n129), .ZN(n131) );
  OR2_X1 U101 ( .A1(n189), .A2(d[2]), .ZN(n129) );
  OR2_X1 U102 ( .A1(n179), .A2(c[2]), .ZN(n130) );
  OR2_X1 U103 ( .A1(n128), .A2(n212), .ZN(y[1]) );
  OR2_X1 U104 ( .A1(n126), .A2(n188), .ZN(n127) );
  AND2_X1 U105 ( .A1(n188), .A2(n126), .ZN(n128) );
  AND2_X1 U106 ( .A1(n125), .A2(n124), .ZN(n126) );
  OR2_X1 U107 ( .A1(n211), .A2(b[1]), .ZN(n124) );
  OR2_X1 U108 ( .A1(n202), .A2(a[1]), .ZN(n125) );
  AND2_X1 U109 ( .A1(n122), .A2(n121), .ZN(n123) );
  OR2_X1 U110 ( .A1(n187), .A2(d[1]), .ZN(n121) );
  OR2_X1 U111 ( .A1(n178), .A2(c[1]), .ZN(n122) );
  OR2_X1 U112 ( .A1(n120), .A2(n210), .ZN(y[0]) );
  OR2_X1 U113 ( .A1(n118), .A2(n186), .ZN(n119) );
  AND2_X1 U114 ( .A1(n186), .A2(n118), .ZN(n120) );
  AND2_X1 U115 ( .A1(n117), .A2(n116), .ZN(n118) );
  OR2_X1 U116 ( .A1(n209), .A2(b[0]), .ZN(n116) );
  OR2_X1 U117 ( .A1(n201), .A2(a[0]), .ZN(n117) );
  AND2_X1 U118 ( .A1(n114), .A2(n113), .ZN(n115) );
  OR2_X1 U119 ( .A1(n185), .A2(d[0]), .ZN(n113) );
  OR2_X1 U120 ( .A1(n177), .A2(c[0]), .ZN(n114) );
endmodule


module byteXor4_7 ( a, b, c, d, y );
  input [7:0] a;
  input [7:0] b;
  input [7:0] c;
  input [7:0] d;
  //input_done

  output [7:0] y;
  //output_done

  wire   n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224;
  //wire_done

  INV_X1 U1 ( .A(n175), .ZN(n224) );
  INV_X1 U2 ( .A(a[7]), .ZN(n223) );
  INV_X1 U3 ( .A(n167), .ZN(n222) );
  INV_X1 U4 ( .A(a[6]), .ZN(n221) );
  INV_X1 U5 ( .A(n159), .ZN(n220) );
  INV_X1 U6 ( .A(a[5]), .ZN(n219) );
  INV_X1 U7 ( .A(n151), .ZN(n218) );
  INV_X1 U8 ( .A(a[4]), .ZN(n217) );
  INV_X1 U9 ( .A(n143), .ZN(n216) );
  INV_X1 U10 ( .A(a[3]), .ZN(n215) );
  INV_X1 U11 ( .A(n135), .ZN(n214) );
  INV_X1 U12 ( .A(a[2]), .ZN(n213) );
  INV_X1 U13 ( .A(n127), .ZN(n212) );
  INV_X1 U14 ( .A(a[1]), .ZN(n211) );
  INV_X1 U15 ( .A(n119), .ZN(n210) );
  INV_X1 U16 ( .A(a[0]), .ZN(n209) );
  INV_X1 U17 ( .A(b[7]), .ZN(n208) );
  INV_X1 U18 ( .A(b[6]), .ZN(n207) );
  INV_X1 U19 ( .A(b[5]), .ZN(n206) );
  INV_X1 U20 ( .A(b[4]), .ZN(n205) );
  INV_X1 U21 ( .A(b[3]), .ZN(n204) );
  INV_X1 U22 ( .A(b[2]), .ZN(n203) );
  INV_X1 U23 ( .A(b[1]), .ZN(n202) );
  INV_X1 U24 ( .A(b[0]), .ZN(n201) );
  INV_X1 U25 ( .A(n171), .ZN(n200) );
  INV_X1 U26 ( .A(c[7]), .ZN(n199) );
  INV_X1 U27 ( .A(n163), .ZN(n198) );
  INV_X1 U28 ( .A(c[6]), .ZN(n197) );
  INV_X1 U29 ( .A(n155), .ZN(n196) );
  INV_X1 U30 ( .A(c[5]), .ZN(n195) );
  INV_X1 U31 ( .A(n147), .ZN(n194) );
  INV_X1 U32 ( .A(c[4]), .ZN(n193) );
  INV_X1 U33 ( .A(n139), .ZN(n192) );
  INV_X1 U34 ( .A(c[3]), .ZN(n191) );
  INV_X1 U35 ( .A(n131), .ZN(n190) );
  INV_X1 U36 ( .A(c[2]), .ZN(n189) );
  INV_X1 U37 ( .A(n123), .ZN(n188) );
  INV_X1 U38 ( .A(c[1]), .ZN(n187) );
  INV_X1 U39 ( .A(n115), .ZN(n186) );
  INV_X1 U40 ( .A(c[0]), .ZN(n185) );
  INV_X1 U41 ( .A(d[7]), .ZN(n184) );
  INV_X1 U42 ( .A(d[6]), .ZN(n183) );
  INV_X1 U43 ( .A(d[5]), .ZN(n182) );
  INV_X1 U44 ( .A(d[4]), .ZN(n181) );
  INV_X1 U45 ( .A(d[3]), .ZN(n180) );
  INV_X1 U46 ( .A(d[2]), .ZN(n179) );
  INV_X1 U47 ( .A(d[1]), .ZN(n178) );
  INV_X1 U48 ( .A(d[0]), .ZN(n177) );
  OR2_X1 U49 ( .A1(n176), .A2(n224), .ZN(y[7]) );
  OR2_X1 U50 ( .A1(n174), .A2(n200), .ZN(n175) );
  AND2_X1 U51 ( .A1(n200), .A2(n174), .ZN(n176) );
  AND2_X1 U52 ( .A1(n173), .A2(n172), .ZN(n174) );
  OR2_X1 U53 ( .A1(n223), .A2(b[7]), .ZN(n172) );
  OR2_X1 U54 ( .A1(n208), .A2(a[7]), .ZN(n173) );
  AND2_X1 U55 ( .A1(n170), .A2(n169), .ZN(n171) );
  OR2_X1 U56 ( .A1(n199), .A2(d[7]), .ZN(n169) );
  OR2_X1 U57 ( .A1(n184), .A2(c[7]), .ZN(n170) );
  OR2_X1 U58 ( .A1(n168), .A2(n222), .ZN(y[6]) );
  OR2_X1 U59 ( .A1(n166), .A2(n198), .ZN(n167) );
  AND2_X1 U60 ( .A1(n198), .A2(n166), .ZN(n168) );
  AND2_X1 U61 ( .A1(n165), .A2(n164), .ZN(n166) );
  OR2_X1 U62 ( .A1(n221), .A2(b[6]), .ZN(n164) );
  OR2_X1 U63 ( .A1(n207), .A2(a[6]), .ZN(n165) );
  AND2_X1 U64 ( .A1(n162), .A2(n161), .ZN(n163) );
  OR2_X1 U65 ( .A1(n197), .A2(d[6]), .ZN(n161) );
  OR2_X1 U66 ( .A1(n183), .A2(c[6]), .ZN(n162) );
  OR2_X1 U67 ( .A1(n160), .A2(n220), .ZN(y[5]) );
  OR2_X1 U68 ( .A1(n158), .A2(n196), .ZN(n159) );
  AND2_X1 U69 ( .A1(n196), .A2(n158), .ZN(n160) );
  AND2_X1 U70 ( .A1(n157), .A2(n156), .ZN(n158) );
  OR2_X1 U71 ( .A1(n219), .A2(b[5]), .ZN(n156) );
  OR2_X1 U72 ( .A1(n206), .A2(a[5]), .ZN(n157) );
  AND2_X1 U73 ( .A1(n154), .A2(n153), .ZN(n155) );
  OR2_X1 U74 ( .A1(n195), .A2(d[5]), .ZN(n153) );
  OR2_X1 U75 ( .A1(n182), .A2(c[5]), .ZN(n154) );
  OR2_X1 U76 ( .A1(n152), .A2(n218), .ZN(y[4]) );
  OR2_X1 U77 ( .A1(n150), .A2(n194), .ZN(n151) );
  AND2_X1 U78 ( .A1(n194), .A2(n150), .ZN(n152) );
  AND2_X1 U79 ( .A1(n149), .A2(n148), .ZN(n150) );
  OR2_X1 U80 ( .A1(n217), .A2(b[4]), .ZN(n148) );
  OR2_X1 U81 ( .A1(n205), .A2(a[4]), .ZN(n149) );
  AND2_X1 U82 ( .A1(n146), .A2(n145), .ZN(n147) );
  OR2_X1 U83 ( .A1(n193), .A2(d[4]), .ZN(n145) );
  OR2_X1 U84 ( .A1(n181), .A2(c[4]), .ZN(n146) );
  OR2_X1 U85 ( .A1(n144), .A2(n216), .ZN(y[3]) );
  OR2_X1 U86 ( .A1(n142), .A2(n192), .ZN(n143) );
  AND2_X1 U87 ( .A1(n192), .A2(n142), .ZN(n144) );
  AND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(n142) );
  OR2_X1 U89 ( .A1(n215), .A2(b[3]), .ZN(n140) );
  OR2_X1 U90 ( .A1(n204), .A2(a[3]), .ZN(n141) );
  AND2_X1 U91 ( .A1(n138), .A2(n137), .ZN(n139) );
  OR2_X1 U92 ( .A1(n191), .A2(d[3]), .ZN(n137) );
  OR2_X1 U93 ( .A1(n180), .A2(c[3]), .ZN(n138) );
  OR2_X1 U94 ( .A1(n136), .A2(n214), .ZN(y[2]) );
  OR2_X1 U95 ( .A1(n134), .A2(n190), .ZN(n135) );
  AND2_X1 U96 ( .A1(n190), .A2(n134), .ZN(n136) );
  AND2_X1 U97 ( .A1(n133), .A2(n132), .ZN(n134) );
  OR2_X1 U98 ( .A1(n213), .A2(b[2]), .ZN(n132) );
  OR2_X1 U99 ( .A1(n203), .A2(a[2]), .ZN(n133) );
  AND2_X1 U100 ( .A1(n130), .A2(n129), .ZN(n131) );
  OR2_X1 U101 ( .A1(n189), .A2(d[2]), .ZN(n129) );
  OR2_X1 U102 ( .A1(n179), .A2(c[2]), .ZN(n130) );
  OR2_X1 U103 ( .A1(n128), .A2(n212), .ZN(y[1]) );
  OR2_X1 U104 ( .A1(n126), .A2(n188), .ZN(n127) );
  AND2_X1 U105 ( .A1(n188), .A2(n126), .ZN(n128) );
  AND2_X1 U106 ( .A1(n125), .A2(n124), .ZN(n126) );
  OR2_X1 U107 ( .A1(n211), .A2(b[1]), .ZN(n124) );
  OR2_X1 U108 ( .A1(n202), .A2(a[1]), .ZN(n125) );
  AND2_X1 U109 ( .A1(n122), .A2(n121), .ZN(n123) );
  OR2_X1 U110 ( .A1(n187), .A2(d[1]), .ZN(n121) );
  OR2_X1 U111 ( .A1(n178), .A2(c[1]), .ZN(n122) );
  OR2_X1 U112 ( .A1(n120), .A2(n210), .ZN(y[0]) );
  OR2_X1 U113 ( .A1(n118), .A2(n186), .ZN(n119) );
  AND2_X1 U114 ( .A1(n186), .A2(n118), .ZN(n120) );
  AND2_X1 U115 ( .A1(n117), .A2(n116), .ZN(n118) );
  OR2_X1 U116 ( .A1(n209), .A2(b[0]), .ZN(n116) );
  OR2_X1 U117 ( .A1(n201), .A2(a[0]), .ZN(n117) );
  AND2_X1 U118 ( .A1(n114), .A2(n113), .ZN(n115) );
  OR2_X1 U119 ( .A1(n185), .A2(d[0]), .ZN(n113) );
  OR2_X1 U120 ( .A1(n177), .A2(c[0]), .ZN(n114) );
endmodule


module byteXor4_8 ( a, b, c, d, y );
  input [7:0] a;
  input [7:0] b;
  input [7:0] c;
  input [7:0] d;
  //input_done

  output [7:0] y;
  //output_done

  wire   n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224;
  //wire_done

  INV_X1 U1 ( .A(n175), .ZN(n224) );
  INV_X1 U2 ( .A(a[7]), .ZN(n223) );
  INV_X1 U3 ( .A(n167), .ZN(n222) );
  INV_X1 U4 ( .A(a[6]), .ZN(n221) );
  INV_X1 U5 ( .A(n159), .ZN(n220) );
  INV_X1 U6 ( .A(a[5]), .ZN(n219) );
  INV_X1 U7 ( .A(n151), .ZN(n218) );
  INV_X1 U8 ( .A(a[4]), .ZN(n217) );
  INV_X1 U9 ( .A(n143), .ZN(n216) );
  INV_X1 U10 ( .A(a[3]), .ZN(n215) );
  INV_X1 U11 ( .A(n135), .ZN(n214) );
  INV_X1 U12 ( .A(a[2]), .ZN(n213) );
  INV_X1 U13 ( .A(n127), .ZN(n212) );
  INV_X1 U14 ( .A(a[1]), .ZN(n211) );
  INV_X1 U15 ( .A(n119), .ZN(n210) );
  INV_X1 U16 ( .A(a[0]), .ZN(n209) );
  INV_X1 U17 ( .A(b[7]), .ZN(n208) );
  INV_X1 U18 ( .A(b[6]), .ZN(n207) );
  INV_X1 U19 ( .A(b[5]), .ZN(n206) );
  INV_X1 U20 ( .A(b[4]), .ZN(n205) );
  INV_X1 U21 ( .A(b[3]), .ZN(n204) );
  INV_X1 U22 ( .A(b[2]), .ZN(n203) );
  INV_X1 U23 ( .A(b[1]), .ZN(n202) );
  INV_X1 U24 ( .A(b[0]), .ZN(n201) );
  INV_X1 U25 ( .A(n171), .ZN(n200) );
  INV_X1 U26 ( .A(c[7]), .ZN(n199) );
  INV_X1 U27 ( .A(n163), .ZN(n198) );
  INV_X1 U28 ( .A(c[6]), .ZN(n197) );
  INV_X1 U29 ( .A(n155), .ZN(n196) );
  INV_X1 U30 ( .A(c[5]), .ZN(n195) );
  INV_X1 U31 ( .A(n147), .ZN(n194) );
  INV_X1 U32 ( .A(c[4]), .ZN(n193) );
  INV_X1 U33 ( .A(n139), .ZN(n192) );
  INV_X1 U34 ( .A(c[3]), .ZN(n191) );
  INV_X1 U35 ( .A(n131), .ZN(n190) );
  INV_X1 U36 ( .A(c[2]), .ZN(n189) );
  INV_X1 U37 ( .A(n123), .ZN(n188) );
  INV_X1 U38 ( .A(c[1]), .ZN(n187) );
  INV_X1 U39 ( .A(n115), .ZN(n186) );
  INV_X1 U40 ( .A(c[0]), .ZN(n185) );
  INV_X1 U41 ( .A(d[7]), .ZN(n184) );
  INV_X1 U42 ( .A(d[6]), .ZN(n183) );
  INV_X1 U43 ( .A(d[5]), .ZN(n182) );
  INV_X1 U44 ( .A(d[4]), .ZN(n181) );
  INV_X1 U45 ( .A(d[3]), .ZN(n180) );
  INV_X1 U46 ( .A(d[2]), .ZN(n179) );
  INV_X1 U47 ( .A(d[1]), .ZN(n178) );
  INV_X1 U48 ( .A(d[0]), .ZN(n177) );
  OR2_X1 U49 ( .A1(n176), .A2(n224), .ZN(y[7]) );
  OR2_X1 U50 ( .A1(n174), .A2(n200), .ZN(n175) );
  AND2_X1 U51 ( .A1(n200), .A2(n174), .ZN(n176) );
  AND2_X1 U52 ( .A1(n173), .A2(n172), .ZN(n174) );
  OR2_X1 U53 ( .A1(n223), .A2(b[7]), .ZN(n172) );
  OR2_X1 U54 ( .A1(n208), .A2(a[7]), .ZN(n173) );
  AND2_X1 U55 ( .A1(n170), .A2(n169), .ZN(n171) );
  OR2_X1 U56 ( .A1(n199), .A2(d[7]), .ZN(n169) );
  OR2_X1 U57 ( .A1(n184), .A2(c[7]), .ZN(n170) );
  OR2_X1 U58 ( .A1(n168), .A2(n222), .ZN(y[6]) );
  OR2_X1 U59 ( .A1(n166), .A2(n198), .ZN(n167) );
  AND2_X1 U60 ( .A1(n198), .A2(n166), .ZN(n168) );
  AND2_X1 U61 ( .A1(n165), .A2(n164), .ZN(n166) );
  OR2_X1 U62 ( .A1(n221), .A2(b[6]), .ZN(n164) );
  OR2_X1 U63 ( .A1(n207), .A2(a[6]), .ZN(n165) );
  AND2_X1 U64 ( .A1(n162), .A2(n161), .ZN(n163) );
  OR2_X1 U65 ( .A1(n197), .A2(d[6]), .ZN(n161) );
  OR2_X1 U66 ( .A1(n183), .A2(c[6]), .ZN(n162) );
  OR2_X1 U67 ( .A1(n160), .A2(n220), .ZN(y[5]) );
  OR2_X1 U68 ( .A1(n158), .A2(n196), .ZN(n159) );
  AND2_X1 U69 ( .A1(n196), .A2(n158), .ZN(n160) );
  AND2_X1 U70 ( .A1(n157), .A2(n156), .ZN(n158) );
  OR2_X1 U71 ( .A1(n219), .A2(b[5]), .ZN(n156) );
  OR2_X1 U72 ( .A1(n206), .A2(a[5]), .ZN(n157) );
  AND2_X1 U73 ( .A1(n154), .A2(n153), .ZN(n155) );
  OR2_X1 U74 ( .A1(n195), .A2(d[5]), .ZN(n153) );
  OR2_X1 U75 ( .A1(n182), .A2(c[5]), .ZN(n154) );
  OR2_X1 U76 ( .A1(n152), .A2(n218), .ZN(y[4]) );
  OR2_X1 U77 ( .A1(n150), .A2(n194), .ZN(n151) );
  AND2_X1 U78 ( .A1(n194), .A2(n150), .ZN(n152) );
  AND2_X1 U79 ( .A1(n149), .A2(n148), .ZN(n150) );
  OR2_X1 U80 ( .A1(n217), .A2(b[4]), .ZN(n148) );
  OR2_X1 U81 ( .A1(n205), .A2(a[4]), .ZN(n149) );
  AND2_X1 U82 ( .A1(n146), .A2(n145), .ZN(n147) );
  OR2_X1 U83 ( .A1(n193), .A2(d[4]), .ZN(n145) );
  OR2_X1 U84 ( .A1(n181), .A2(c[4]), .ZN(n146) );
  OR2_X1 U85 ( .A1(n144), .A2(n216), .ZN(y[3]) );
  OR2_X1 U86 ( .A1(n142), .A2(n192), .ZN(n143) );
  AND2_X1 U87 ( .A1(n192), .A2(n142), .ZN(n144) );
  AND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(n142) );
  OR2_X1 U89 ( .A1(n215), .A2(b[3]), .ZN(n140) );
  OR2_X1 U90 ( .A1(n204), .A2(a[3]), .ZN(n141) );
  AND2_X1 U91 ( .A1(n138), .A2(n137), .ZN(n139) );
  OR2_X1 U92 ( .A1(n191), .A2(d[3]), .ZN(n137) );
  OR2_X1 U93 ( .A1(n180), .A2(c[3]), .ZN(n138) );
  OR2_X1 U94 ( .A1(n136), .A2(n214), .ZN(y[2]) );
  OR2_X1 U95 ( .A1(n134), .A2(n190), .ZN(n135) );
  AND2_X1 U96 ( .A1(n190), .A2(n134), .ZN(n136) );
  AND2_X1 U97 ( .A1(n133), .A2(n132), .ZN(n134) );
  OR2_X1 U98 ( .A1(n213), .A2(b[2]), .ZN(n132) );
  OR2_X1 U99 ( .A1(n203), .A2(a[2]), .ZN(n133) );
  AND2_X1 U100 ( .A1(n130), .A2(n129), .ZN(n131) );
  OR2_X1 U101 ( .A1(n189), .A2(d[2]), .ZN(n129) );
  OR2_X1 U102 ( .A1(n179), .A2(c[2]), .ZN(n130) );
  OR2_X1 U103 ( .A1(n128), .A2(n212), .ZN(y[1]) );
  OR2_X1 U104 ( .A1(n126), .A2(n188), .ZN(n127) );
  AND2_X1 U105 ( .A1(n188), .A2(n126), .ZN(n128) );
  AND2_X1 U106 ( .A1(n125), .A2(n124), .ZN(n126) );
  OR2_X1 U107 ( .A1(n211), .A2(b[1]), .ZN(n124) );
  OR2_X1 U108 ( .A1(n202), .A2(a[1]), .ZN(n125) );
  AND2_X1 U109 ( .A1(n122), .A2(n121), .ZN(n123) );
  OR2_X1 U110 ( .A1(n187), .A2(d[1]), .ZN(n121) );
  OR2_X1 U111 ( .A1(n178), .A2(c[1]), .ZN(n122) );
  OR2_X1 U112 ( .A1(n120), .A2(n210), .ZN(y[0]) );
  OR2_X1 U113 ( .A1(n118), .A2(n186), .ZN(n119) );
  AND2_X1 U114 ( .A1(n186), .A2(n118), .ZN(n120) );
  AND2_X1 U115 ( .A1(n117), .A2(n116), .ZN(n118) );
  OR2_X1 U116 ( .A1(n209), .A2(b[0]), .ZN(n116) );
  OR2_X1 U117 ( .A1(n201), .A2(a[0]), .ZN(n117) );
  AND2_X1 U118 ( .A1(n114), .A2(n113), .ZN(n115) );
  OR2_X1 U119 ( .A1(n185), .A2(d[0]), .ZN(n113) );
  OR2_X1 U120 ( .A1(n177), .A2(c[0]), .ZN(n114) );
endmodule


module mixCol_2 ( in, out );
  input [31:0] in;
  //input_done

  output [31:0] out;
  //output_done

  wire   [7:0] b0_s2;
  wire   [7:0] b1_s2;
  wire   [7:0] b2_s2;
  wire   [7:0] b3_s2;
  wire   [7:0] b0_s3;
  wire   [7:0] b1_s3;
  wire   [7:0] b2_s3;
  wire   [7:0] b3_s3;
  //wire_done

  scale2_8 b0_scale2 ( .in(in[31:24]), .out(b0_s2) );
  scale2_7 b1_scale2 ( .in(in[23:16]), .out(b1_s2) );
  scale2_6 b2_scale2 ( .in(in[15:8]), .out(b2_s2) );
  scale2_5 b3_scale2 ( .in(in[7:0]), .out(b3_s2) );
  byteXor_9 b0_scale3 ( .a(in[31:24]), .b(b0_s2), .y(b0_s3) );
  byteXor_8 b1_scale3 ( .a(in[23:16]), .b(b1_s2), .y(b1_s3) );
  byteXor_7 b2_scale3 ( .a(in[15:8]), .b(b2_s2), .y(b2_s3) );
  byteXor_6 b3_scale3 ( .a(in[7:0]), .b(b3_s2), .y(b3_s3) );
  byteXor4_8 out0 ( .a(b0_s2), .b(b1_s3), .c(in[15:8]), .d(in[7:0]), .y(
        out[31:24]) );
  byteXor4_7 out1 ( .a(in[31:24]), .b(b1_s2), .c(b2_s3), .d(in[7:0]), .y(
        out[23:16]) );
  byteXor4_6 out2 ( .a(in[31:24]), .b(in[23:16]), .c(b2_s2), .d(b3_s3), .y(
        out[15:8]) );
  byteXor4_5 out3 ( .a(b0_s3), .b(in[23:16]), .c(in[15:8]), .d(b3_s2), .y(
        out[7:0]) );
endmodule


module scale2_9 ( in, out );
  input [7:0] in;
  //input_done

  output [7:0] out;
  //output_done

  wire   in_0, \in[6] , \in[5] , \in[4] , \in[1] , \in[7] , n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20;
  //wire_done

  assign in_0 = in[0];
  assign out[7] = \in[6] ;
  assign \in[6]  = in[6];
  assign out[6] = \in[5] ;
  assign \in[5]  = in[5];
  assign out[5] = \in[4] ;
  assign \in[4]  = in[4];
  assign out[2] = \in[1] ;
  assign \in[1]  = in[1];
  assign out[0] = \in[7] ;
  assign \in[7]  = in[7];

  INV_X1 U1 ( .A(\in[7]), .ZN(n20) );
  INV_X1 U2 ( .A(in[3]), .ZN(n19) );
  INV_X1 U3 ( .A(in[2]), .ZN(n18) );
  INV_X1 U4 ( .A(in_0), .ZN(n17) );
  OR2_X1 U5 ( .A1(n16), .A2(n15), .ZN(out[4]) );
  AND2_X1 U6 ( .A1(in[3]), .A2(n20), .ZN(n15) );
  AND2_X1 U7 ( .A1(\in[7]), .A2(n19), .ZN(n16) );
  OR2_X1 U8 ( .A1(n14), .A2(n13), .ZN(out[3]) );
  AND2_X1 U9 ( .A1(in[2]), .A2(n20), .ZN(n13) );
  AND2_X1 U10 ( .A1(\in[7]), .A2(n18), .ZN(n14) );
  OR2_X1 U11 ( .A1(n12), .A2(n11), .ZN(out[1]) );
  AND2_X1 U12 ( .A1(in_0), .A2(n20), .ZN(n11) );
  AND2_X1 U13 ( .A1(\in[7]), .A2(n17), .ZN(n12) );
endmodule


module scale2_10 ( in, out );
  input [7:0] in;
  //input_done

  output [7:0] out;
  //output_done

  wire   in_0, \in[6] , \in[5] , \in[4] , \in[1] , \in[7] , n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20;
  //wire_done

  assign in_0 = in[0];
  assign out[7] = \in[6] ;
  assign \in[6]  = in[6];
  assign out[6] = \in[5] ;
  assign \in[5]  = in[5];
  assign out[5] = \in[4] ;
  assign \in[4]  = in[4];
  assign out[2] = \in[1] ;
  assign \in[1]  = in[1];
  assign out[0] = \in[7] ;
  assign \in[7]  = in[7];

  INV_X1 U1 ( .A(\in[7]), .ZN(n20) );
  INV_X1 U2 ( .A(in[3]), .ZN(n19) );
  INV_X1 U3 ( .A(in[2]), .ZN(n18) );
  INV_X1 U4 ( .A(in_0), .ZN(n17) );
  OR2_X1 U5 ( .A1(n16), .A2(n15), .ZN(out[4]) );
  AND2_X1 U6 ( .A1(in[3]), .A2(n20), .ZN(n15) );
  AND2_X1 U7 ( .A1(\in[7]), .A2(n19), .ZN(n16) );
  OR2_X1 U8 ( .A1(n14), .A2(n13), .ZN(out[3]) );
  AND2_X1 U9 ( .A1(in[2]), .A2(n20), .ZN(n13) );
  AND2_X1 U10 ( .A1(\in[7]), .A2(n18), .ZN(n14) );
  OR2_X1 U11 ( .A1(n12), .A2(n11), .ZN(out[1]) );
  AND2_X1 U12 ( .A1(in_0), .A2(n20), .ZN(n11) );
  AND2_X1 U13 ( .A1(\in[7]), .A2(n17), .ZN(n12) );
endmodule


module scale2_11 ( in, out );
  input [7:0] in;
  //input_done

  output [7:0] out;
  //output_done

  wire   in_0, \in[6] , \in[5] , \in[4] , \in[1] , \in[7] , n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20;
  //wire_done

  assign in_0 = in[0];
  assign out[7] = \in[6] ;
  assign \in[6]  = in[6];
  assign out[6] = \in[5] ;
  assign \in[5]  = in[5];
  assign out[5] = \in[4] ;
  assign \in[4]  = in[4];
  assign out[2] = \in[1] ;
  assign \in[1]  = in[1];
  assign out[0] = \in[7] ;
  assign \in[7]  = in[7];

  INV_X1 U1 ( .A(\in[7]), .ZN(n20) );
  INV_X1 U2 ( .A(in[3]), .ZN(n19) );
  INV_X1 U3 ( .A(in[2]), .ZN(n18) );
  INV_X1 U4 ( .A(in_0), .ZN(n17) );
  OR2_X1 U5 ( .A1(n16), .A2(n15), .ZN(out[4]) );
  AND2_X1 U6 ( .A1(in[3]), .A2(n20), .ZN(n15) );
  AND2_X1 U7 ( .A1(\in[7]), .A2(n19), .ZN(n16) );
  OR2_X1 U8 ( .A1(n14), .A2(n13), .ZN(out[3]) );
  AND2_X1 U9 ( .A1(in[2]), .A2(n20), .ZN(n13) );
  AND2_X1 U10 ( .A1(\in[7]), .A2(n18), .ZN(n14) );
  OR2_X1 U11 ( .A1(n12), .A2(n11), .ZN(out[1]) );
  AND2_X1 U12 ( .A1(in_0), .A2(n20), .ZN(n11) );
  AND2_X1 U13 ( .A1(\in[7]), .A2(n17), .ZN(n12) );
endmodule


module scale2_12 ( in, out );
  input [7:0] in;
  //input_done

  output [7:0] out;
  //output_done

  wire   in_0, \in[6] , \in[5] , \in[4] , \in[1] , \in[7] , n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20;
  //wire_done

  assign in_0 = in[0];
  assign out[7] = \in[6] ;
  assign \in[6]  = in[6];
  assign out[6] = \in[5] ;
  assign \in[5]  = in[5];
  assign out[5] = \in[4] ;
  assign \in[4]  = in[4];
  assign out[2] = \in[1] ;
  assign \in[1]  = in[1];
  assign out[0] = \in[7] ;
  assign \in[7]  = in[7];

  INV_X1 U1 ( .A(\in[7]), .ZN(n20) );
  INV_X1 U2 ( .A(in[3]), .ZN(n19) );
  INV_X1 U3 ( .A(in[2]), .ZN(n18) );
  INV_X1 U4 ( .A(in_0), .ZN(n17) );
  OR2_X1 U5 ( .A1(n16), .A2(n15), .ZN(out[4]) );
  AND2_X1 U6 ( .A1(in[3]), .A2(n20), .ZN(n15) );
  AND2_X1 U7 ( .A1(\in[7]), .A2(n19), .ZN(n16) );
  OR2_X1 U8 ( .A1(n14), .A2(n13), .ZN(out[3]) );
  AND2_X1 U9 ( .A1(in[2]), .A2(n20), .ZN(n13) );
  AND2_X1 U10 ( .A1(\in[7]), .A2(n18), .ZN(n14) );
  OR2_X1 U11 ( .A1(n12), .A2(n11), .ZN(out[1]) );
  AND2_X1 U12 ( .A1(in_0), .A2(n20), .ZN(n11) );
  AND2_X1 U13 ( .A1(\in[7]), .A2(n17), .ZN(n12) );
endmodule


module byteXor_10 ( a, b, y );
  input [7:0] a;
  input [7:0] b;
  //input_done

  output [7:0] y;
  //output_done

  wire   n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64;
  //wire_done

  INV_X1 U1 ( .A(n47), .ZN(n64) );
  INV_X1 U2 ( .A(a[7]), .ZN(n63) );
  INV_X1 U3 ( .A(n45), .ZN(n62) );
  INV_X1 U4 ( .A(a[6]), .ZN(n61) );
  INV_X1 U5 ( .A(n43), .ZN(n60) );
  INV_X1 U6 ( .A(a[5]), .ZN(n59) );
  INV_X1 U7 ( .A(n41), .ZN(n58) );
  INV_X1 U8 ( .A(a[4]), .ZN(n57) );
  INV_X1 U9 ( .A(n39), .ZN(n56) );
  INV_X1 U10 ( .A(a[3]), .ZN(n55) );
  INV_X1 U11 ( .A(n37), .ZN(n54) );
  INV_X1 U12 ( .A(a[2]), .ZN(n53) );
  INV_X1 U13 ( .A(n35), .ZN(n52) );
  INV_X1 U14 ( .A(a[1]), .ZN(n51) );
  INV_X1 U15 ( .A(n33), .ZN(n50) );
  INV_X1 U16 ( .A(a[0]), .ZN(n49) );
  OR2_X1 U17 ( .A1(n48), .A2(n64), .ZN(y[7]) );
  OR2_X1 U18 ( .A1(n63), .A2(b[7]), .ZN(n47) );
  AND2_X1 U19 ( .A1(b[7]), .A2(n63), .ZN(n48) );
  OR2_X1 U20 ( .A1(n46), .A2(n62), .ZN(y[6]) );
  OR2_X1 U21 ( .A1(n61), .A2(b[6]), .ZN(n45) );
  AND2_X1 U22 ( .A1(b[6]), .A2(n61), .ZN(n46) );
  OR2_X1 U23 ( .A1(n44), .A2(n60), .ZN(y[5]) );
  OR2_X1 U24 ( .A1(n59), .A2(b[5]), .ZN(n43) );
  AND2_X1 U25 ( .A1(b[5]), .A2(n59), .ZN(n44) );
  OR2_X1 U26 ( .A1(n42), .A2(n58), .ZN(y[4]) );
  OR2_X1 U27 ( .A1(n57), .A2(b[4]), .ZN(n41) );
  AND2_X1 U28 ( .A1(b[4]), .A2(n57), .ZN(n42) );
  OR2_X1 U29 ( .A1(n40), .A2(n56), .ZN(y[3]) );
  OR2_X1 U30 ( .A1(n55), .A2(b[3]), .ZN(n39) );
  AND2_X1 U31 ( .A1(b[3]), .A2(n55), .ZN(n40) );
  OR2_X1 U32 ( .A1(n38), .A2(n54), .ZN(y[2]) );
  OR2_X1 U33 ( .A1(n53), .A2(b[2]), .ZN(n37) );
  AND2_X1 U34 ( .A1(b[2]), .A2(n53), .ZN(n38) );
  OR2_X1 U35 ( .A1(n36), .A2(n52), .ZN(y[1]) );
  OR2_X1 U36 ( .A1(n51), .A2(b[1]), .ZN(n35) );
  AND2_X1 U37 ( .A1(b[1]), .A2(n51), .ZN(n36) );
  OR2_X1 U38 ( .A1(n34), .A2(n50), .ZN(y[0]) );
  OR2_X1 U39 ( .A1(n49), .A2(b[0]), .ZN(n33) );
  AND2_X1 U40 ( .A1(b[0]), .A2(n49), .ZN(n34) );
endmodule


module byteXor_11 ( a, b, y );
  input [7:0] a;
  input [7:0] b;
  //input_done

  output [7:0] y;
  //output_done

  wire   n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64;
  //wire_done

  INV_X1 U1 ( .A(n47), .ZN(n64) );
  INV_X1 U2 ( .A(a[7]), .ZN(n63) );
  INV_X1 U3 ( .A(n45), .ZN(n62) );
  INV_X1 U4 ( .A(a[6]), .ZN(n61) );
  INV_X1 U5 ( .A(n43), .ZN(n60) );
  INV_X1 U6 ( .A(a[5]), .ZN(n59) );
  INV_X1 U7 ( .A(n41), .ZN(n58) );
  INV_X1 U8 ( .A(a[4]), .ZN(n57) );
  INV_X1 U9 ( .A(n39), .ZN(n56) );
  INV_X1 U10 ( .A(a[3]), .ZN(n55) );
  INV_X1 U11 ( .A(n37), .ZN(n54) );
  INV_X1 U12 ( .A(a[2]), .ZN(n53) );
  INV_X1 U13 ( .A(n35), .ZN(n52) );
  INV_X1 U14 ( .A(a[1]), .ZN(n51) );
  INV_X1 U15 ( .A(n33), .ZN(n50) );
  INV_X1 U16 ( .A(a[0]), .ZN(n49) );
  OR2_X1 U17 ( .A1(n48), .A2(n64), .ZN(y[7]) );
  OR2_X1 U18 ( .A1(n63), .A2(b[7]), .ZN(n47) );
  AND2_X1 U19 ( .A1(b[7]), .A2(n63), .ZN(n48) );
  OR2_X1 U20 ( .A1(n46), .A2(n62), .ZN(y[6]) );
  OR2_X1 U21 ( .A1(n61), .A2(b[6]), .ZN(n45) );
  AND2_X1 U22 ( .A1(b[6]), .A2(n61), .ZN(n46) );
  OR2_X1 U23 ( .A1(n44), .A2(n60), .ZN(y[5]) );
  OR2_X1 U24 ( .A1(n59), .A2(b[5]), .ZN(n43) );
  AND2_X1 U25 ( .A1(b[5]), .A2(n59), .ZN(n44) );
  OR2_X1 U26 ( .A1(n42), .A2(n58), .ZN(y[4]) );
  OR2_X1 U27 ( .A1(n57), .A2(b[4]), .ZN(n41) );
  AND2_X1 U28 ( .A1(b[4]), .A2(n57), .ZN(n42) );
  OR2_X1 U29 ( .A1(n40), .A2(n56), .ZN(y[3]) );
  OR2_X1 U30 ( .A1(n55), .A2(b[3]), .ZN(n39) );
  AND2_X1 U31 ( .A1(b[3]), .A2(n55), .ZN(n40) );
  OR2_X1 U32 ( .A1(n38), .A2(n54), .ZN(y[2]) );
  OR2_X1 U33 ( .A1(n53), .A2(b[2]), .ZN(n37) );
  AND2_X1 U34 ( .A1(b[2]), .A2(n53), .ZN(n38) );
  OR2_X1 U35 ( .A1(n36), .A2(n52), .ZN(y[1]) );
  OR2_X1 U36 ( .A1(n51), .A2(b[1]), .ZN(n35) );
  AND2_X1 U37 ( .A1(b[1]), .A2(n51), .ZN(n36) );
  OR2_X1 U38 ( .A1(n34), .A2(n50), .ZN(y[0]) );
  OR2_X1 U39 ( .A1(n49), .A2(b[0]), .ZN(n33) );
  AND2_X1 U40 ( .A1(b[0]), .A2(n49), .ZN(n34) );
endmodule


module byteXor_12 ( a, b, y );
  input [7:0] a;
  input [7:0] b;
  //input_done

  output [7:0] y;
  //output_done

  wire   n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64;
  //wire_done

  INV_X1 U1 ( .A(n47), .ZN(n64) );
  INV_X1 U2 ( .A(a[7]), .ZN(n63) );
  INV_X1 U3 ( .A(n45), .ZN(n62) );
  INV_X1 U4 ( .A(a[6]), .ZN(n61) );
  INV_X1 U5 ( .A(n43), .ZN(n60) );
  INV_X1 U6 ( .A(a[5]), .ZN(n59) );
  INV_X1 U7 ( .A(n41), .ZN(n58) );
  INV_X1 U8 ( .A(a[4]), .ZN(n57) );
  INV_X1 U9 ( .A(n39), .ZN(n56) );
  INV_X1 U10 ( .A(a[3]), .ZN(n55) );
  INV_X1 U11 ( .A(n37), .ZN(n54) );
  INV_X1 U12 ( .A(a[2]), .ZN(n53) );
  INV_X1 U13 ( .A(n35), .ZN(n52) );
  INV_X1 U14 ( .A(a[1]), .ZN(n51) );
  INV_X1 U15 ( .A(n33), .ZN(n50) );
  INV_X1 U16 ( .A(a[0]), .ZN(n49) );
  OR2_X1 U17 ( .A1(n48), .A2(n64), .ZN(y[7]) );
  OR2_X1 U18 ( .A1(n63), .A2(b[7]), .ZN(n47) );
  AND2_X1 U19 ( .A1(b[7]), .A2(n63), .ZN(n48) );
  OR2_X1 U20 ( .A1(n46), .A2(n62), .ZN(y[6]) );
  OR2_X1 U21 ( .A1(n61), .A2(b[6]), .ZN(n45) );
  AND2_X1 U22 ( .A1(b[6]), .A2(n61), .ZN(n46) );
  OR2_X1 U23 ( .A1(n44), .A2(n60), .ZN(y[5]) );
  OR2_X1 U24 ( .A1(n59), .A2(b[5]), .ZN(n43) );
  AND2_X1 U25 ( .A1(b[5]), .A2(n59), .ZN(n44) );
  OR2_X1 U26 ( .A1(n42), .A2(n58), .ZN(y[4]) );
  OR2_X1 U27 ( .A1(n57), .A2(b[4]), .ZN(n41) );
  AND2_X1 U28 ( .A1(b[4]), .A2(n57), .ZN(n42) );
  OR2_X1 U29 ( .A1(n40), .A2(n56), .ZN(y[3]) );
  OR2_X1 U30 ( .A1(n55), .A2(b[3]), .ZN(n39) );
  AND2_X1 U31 ( .A1(b[3]), .A2(n55), .ZN(n40) );
  OR2_X1 U32 ( .A1(n38), .A2(n54), .ZN(y[2]) );
  OR2_X1 U33 ( .A1(n53), .A2(b[2]), .ZN(n37) );
  AND2_X1 U34 ( .A1(b[2]), .A2(n53), .ZN(n38) );
  OR2_X1 U35 ( .A1(n36), .A2(n52), .ZN(y[1]) );
  OR2_X1 U36 ( .A1(n51), .A2(b[1]), .ZN(n35) );
  AND2_X1 U37 ( .A1(b[1]), .A2(n51), .ZN(n36) );
  OR2_X1 U38 ( .A1(n34), .A2(n50), .ZN(y[0]) );
  OR2_X1 U39 ( .A1(n49), .A2(b[0]), .ZN(n33) );
  AND2_X1 U40 ( .A1(b[0]), .A2(n49), .ZN(n34) );
endmodule


module byteXor_13 ( a, b, y );
  input [7:0] a;
  input [7:0] b;
  //input_done

  output [7:0] y;
  //output_done

  wire   n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64;
  //wire_done

  INV_X1 U1 ( .A(n47), .ZN(n64) );
  INV_X1 U2 ( .A(a[7]), .ZN(n63) );
  INV_X1 U3 ( .A(n45), .ZN(n62) );
  INV_X1 U4 ( .A(a[6]), .ZN(n61) );
  INV_X1 U5 ( .A(n43), .ZN(n60) );
  INV_X1 U6 ( .A(a[5]), .ZN(n59) );
  INV_X1 U7 ( .A(n41), .ZN(n58) );
  INV_X1 U8 ( .A(a[4]), .ZN(n57) );
  INV_X1 U9 ( .A(n39), .ZN(n56) );
  INV_X1 U10 ( .A(a[3]), .ZN(n55) );
  INV_X1 U11 ( .A(n37), .ZN(n54) );
  INV_X1 U12 ( .A(a[2]), .ZN(n53) );
  INV_X1 U13 ( .A(n35), .ZN(n52) );
  INV_X1 U14 ( .A(a[1]), .ZN(n51) );
  INV_X1 U15 ( .A(n33), .ZN(n50) );
  INV_X1 U16 ( .A(a[0]), .ZN(n49) );
  OR2_X1 U17 ( .A1(n48), .A2(n64), .ZN(y[7]) );
  OR2_X1 U18 ( .A1(n63), .A2(b[7]), .ZN(n47) );
  AND2_X1 U19 ( .A1(b[7]), .A2(n63), .ZN(n48) );
  OR2_X1 U20 ( .A1(n46), .A2(n62), .ZN(y[6]) );
  OR2_X1 U21 ( .A1(n61), .A2(b[6]), .ZN(n45) );
  AND2_X1 U22 ( .A1(b[6]), .A2(n61), .ZN(n46) );
  OR2_X1 U23 ( .A1(n44), .A2(n60), .ZN(y[5]) );
  OR2_X1 U24 ( .A1(n59), .A2(b[5]), .ZN(n43) );
  AND2_X1 U25 ( .A1(b[5]), .A2(n59), .ZN(n44) );
  OR2_X1 U26 ( .A1(n42), .A2(n58), .ZN(y[4]) );
  OR2_X1 U27 ( .A1(n57), .A2(b[4]), .ZN(n41) );
  AND2_X1 U28 ( .A1(b[4]), .A2(n57), .ZN(n42) );
  OR2_X1 U29 ( .A1(n40), .A2(n56), .ZN(y[3]) );
  OR2_X1 U30 ( .A1(n55), .A2(b[3]), .ZN(n39) );
  AND2_X1 U31 ( .A1(b[3]), .A2(n55), .ZN(n40) );
  OR2_X1 U32 ( .A1(n38), .A2(n54), .ZN(y[2]) );
  OR2_X1 U33 ( .A1(n53), .A2(b[2]), .ZN(n37) );
  AND2_X1 U34 ( .A1(b[2]), .A2(n53), .ZN(n38) );
  OR2_X1 U35 ( .A1(n36), .A2(n52), .ZN(y[1]) );
  OR2_X1 U36 ( .A1(n51), .A2(b[1]), .ZN(n35) );
  AND2_X1 U37 ( .A1(b[1]), .A2(n51), .ZN(n36) );
  OR2_X1 U38 ( .A1(n34), .A2(n50), .ZN(y[0]) );
  OR2_X1 U39 ( .A1(n49), .A2(b[0]), .ZN(n33) );
  AND2_X1 U40 ( .A1(b[0]), .A2(n49), .ZN(n34) );
endmodule


module byteXor4_9 ( a, b, c, d, y );
  input [7:0] a;
  input [7:0] b;
  input [7:0] c;
  input [7:0] d;
  //input_done

  output [7:0] y;
  //output_done

  wire   n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224;
  //wire_done

  INV_X1 U1 ( .A(n175), .ZN(n224) );
  INV_X1 U2 ( .A(a[7]), .ZN(n223) );
  INV_X1 U3 ( .A(n167), .ZN(n222) );
  INV_X1 U4 ( .A(a[6]), .ZN(n221) );
  INV_X1 U5 ( .A(n159), .ZN(n220) );
  INV_X1 U6 ( .A(a[5]), .ZN(n219) );
  INV_X1 U7 ( .A(n151), .ZN(n218) );
  INV_X1 U8 ( .A(a[4]), .ZN(n217) );
  INV_X1 U9 ( .A(n143), .ZN(n216) );
  INV_X1 U10 ( .A(a[3]), .ZN(n215) );
  INV_X1 U11 ( .A(n135), .ZN(n214) );
  INV_X1 U12 ( .A(a[2]), .ZN(n213) );
  INV_X1 U13 ( .A(n127), .ZN(n212) );
  INV_X1 U14 ( .A(a[1]), .ZN(n211) );
  INV_X1 U15 ( .A(n119), .ZN(n210) );
  INV_X1 U16 ( .A(a[0]), .ZN(n209) );
  INV_X1 U17 ( .A(b[7]), .ZN(n208) );
  INV_X1 U18 ( .A(b[6]), .ZN(n207) );
  INV_X1 U19 ( .A(b[5]), .ZN(n206) );
  INV_X1 U20 ( .A(b[4]), .ZN(n205) );
  INV_X1 U21 ( .A(b[3]), .ZN(n204) );
  INV_X1 U22 ( .A(b[2]), .ZN(n203) );
  INV_X1 U23 ( .A(b[1]), .ZN(n202) );
  INV_X1 U24 ( .A(b[0]), .ZN(n201) );
  INV_X1 U25 ( .A(n171), .ZN(n200) );
  INV_X1 U26 ( .A(c[7]), .ZN(n199) );
  INV_X1 U27 ( .A(n163), .ZN(n198) );
  INV_X1 U28 ( .A(c[6]), .ZN(n197) );
  INV_X1 U29 ( .A(n155), .ZN(n196) );
  INV_X1 U30 ( .A(c[5]), .ZN(n195) );
  INV_X1 U31 ( .A(n147), .ZN(n194) );
  INV_X1 U32 ( .A(c[4]), .ZN(n193) );
  INV_X1 U33 ( .A(n139), .ZN(n192) );
  INV_X1 U34 ( .A(c[3]), .ZN(n191) );
  INV_X1 U35 ( .A(n131), .ZN(n190) );
  INV_X1 U36 ( .A(c[2]), .ZN(n189) );
  INV_X1 U37 ( .A(n123), .ZN(n188) );
  INV_X1 U38 ( .A(c[1]), .ZN(n187) );
  INV_X1 U39 ( .A(n115), .ZN(n186) );
  INV_X1 U40 ( .A(c[0]), .ZN(n185) );
  INV_X1 U41 ( .A(d[7]), .ZN(n184) );
  INV_X1 U42 ( .A(d[6]), .ZN(n183) );
  INV_X1 U43 ( .A(d[5]), .ZN(n182) );
  INV_X1 U44 ( .A(d[4]), .ZN(n181) );
  INV_X1 U45 ( .A(d[3]), .ZN(n180) );
  INV_X1 U46 ( .A(d[2]), .ZN(n179) );
  INV_X1 U47 ( .A(d[1]), .ZN(n178) );
  INV_X1 U48 ( .A(d[0]), .ZN(n177) );
  OR2_X1 U49 ( .A1(n176), .A2(n224), .ZN(y[7]) );
  OR2_X1 U50 ( .A1(n174), .A2(n200), .ZN(n175) );
  AND2_X1 U51 ( .A1(n200), .A2(n174), .ZN(n176) );
  AND2_X1 U52 ( .A1(n173), .A2(n172), .ZN(n174) );
  OR2_X1 U53 ( .A1(n223), .A2(b[7]), .ZN(n172) );
  OR2_X1 U54 ( .A1(n208), .A2(a[7]), .ZN(n173) );
  AND2_X1 U55 ( .A1(n170), .A2(n169), .ZN(n171) );
  OR2_X1 U56 ( .A1(n199), .A2(d[7]), .ZN(n169) );
  OR2_X1 U57 ( .A1(n184), .A2(c[7]), .ZN(n170) );
  OR2_X1 U58 ( .A1(n168), .A2(n222), .ZN(y[6]) );
  OR2_X1 U59 ( .A1(n166), .A2(n198), .ZN(n167) );
  AND2_X1 U60 ( .A1(n198), .A2(n166), .ZN(n168) );
  AND2_X1 U61 ( .A1(n165), .A2(n164), .ZN(n166) );
  OR2_X1 U62 ( .A1(n221), .A2(b[6]), .ZN(n164) );
  OR2_X1 U63 ( .A1(n207), .A2(a[6]), .ZN(n165) );
  AND2_X1 U64 ( .A1(n162), .A2(n161), .ZN(n163) );
  OR2_X1 U65 ( .A1(n197), .A2(d[6]), .ZN(n161) );
  OR2_X1 U66 ( .A1(n183), .A2(c[6]), .ZN(n162) );
  OR2_X1 U67 ( .A1(n160), .A2(n220), .ZN(y[5]) );
  OR2_X1 U68 ( .A1(n158), .A2(n196), .ZN(n159) );
  AND2_X1 U69 ( .A1(n196), .A2(n158), .ZN(n160) );
  AND2_X1 U70 ( .A1(n157), .A2(n156), .ZN(n158) );
  OR2_X1 U71 ( .A1(n219), .A2(b[5]), .ZN(n156) );
  OR2_X1 U72 ( .A1(n206), .A2(a[5]), .ZN(n157) );
  AND2_X1 U73 ( .A1(n154), .A2(n153), .ZN(n155) );
  OR2_X1 U74 ( .A1(n195), .A2(d[5]), .ZN(n153) );
  OR2_X1 U75 ( .A1(n182), .A2(c[5]), .ZN(n154) );
  OR2_X1 U76 ( .A1(n152), .A2(n218), .ZN(y[4]) );
  OR2_X1 U77 ( .A1(n150), .A2(n194), .ZN(n151) );
  AND2_X1 U78 ( .A1(n194), .A2(n150), .ZN(n152) );
  AND2_X1 U79 ( .A1(n149), .A2(n148), .ZN(n150) );
  OR2_X1 U80 ( .A1(n217), .A2(b[4]), .ZN(n148) );
  OR2_X1 U81 ( .A1(n205), .A2(a[4]), .ZN(n149) );
  AND2_X1 U82 ( .A1(n146), .A2(n145), .ZN(n147) );
  OR2_X1 U83 ( .A1(n193), .A2(d[4]), .ZN(n145) );
  OR2_X1 U84 ( .A1(n181), .A2(c[4]), .ZN(n146) );
  OR2_X1 U85 ( .A1(n144), .A2(n216), .ZN(y[3]) );
  OR2_X1 U86 ( .A1(n142), .A2(n192), .ZN(n143) );
  AND2_X1 U87 ( .A1(n192), .A2(n142), .ZN(n144) );
  AND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(n142) );
  OR2_X1 U89 ( .A1(n215), .A2(b[3]), .ZN(n140) );
  OR2_X1 U90 ( .A1(n204), .A2(a[3]), .ZN(n141) );
  AND2_X1 U91 ( .A1(n138), .A2(n137), .ZN(n139) );
  OR2_X1 U92 ( .A1(n191), .A2(d[3]), .ZN(n137) );
  OR2_X1 U93 ( .A1(n180), .A2(c[3]), .ZN(n138) );
  OR2_X1 U94 ( .A1(n136), .A2(n214), .ZN(y[2]) );
  OR2_X1 U95 ( .A1(n134), .A2(n190), .ZN(n135) );
  AND2_X1 U96 ( .A1(n190), .A2(n134), .ZN(n136) );
  AND2_X1 U97 ( .A1(n133), .A2(n132), .ZN(n134) );
  OR2_X1 U98 ( .A1(n213), .A2(b[2]), .ZN(n132) );
  OR2_X1 U99 ( .A1(n203), .A2(a[2]), .ZN(n133) );
  AND2_X1 U100 ( .A1(n130), .A2(n129), .ZN(n131) );
  OR2_X1 U101 ( .A1(n189), .A2(d[2]), .ZN(n129) );
  OR2_X1 U102 ( .A1(n179), .A2(c[2]), .ZN(n130) );
  OR2_X1 U103 ( .A1(n128), .A2(n212), .ZN(y[1]) );
  OR2_X1 U104 ( .A1(n126), .A2(n188), .ZN(n127) );
  AND2_X1 U105 ( .A1(n188), .A2(n126), .ZN(n128) );
  AND2_X1 U106 ( .A1(n125), .A2(n124), .ZN(n126) );
  OR2_X1 U107 ( .A1(n211), .A2(b[1]), .ZN(n124) );
  OR2_X1 U108 ( .A1(n202), .A2(a[1]), .ZN(n125) );
  AND2_X1 U109 ( .A1(n122), .A2(n121), .ZN(n123) );
  OR2_X1 U110 ( .A1(n187), .A2(d[1]), .ZN(n121) );
  OR2_X1 U111 ( .A1(n178), .A2(c[1]), .ZN(n122) );
  OR2_X1 U112 ( .A1(n120), .A2(n210), .ZN(y[0]) );
  OR2_X1 U113 ( .A1(n118), .A2(n186), .ZN(n119) );
  AND2_X1 U114 ( .A1(n186), .A2(n118), .ZN(n120) );
  AND2_X1 U115 ( .A1(n117), .A2(n116), .ZN(n118) );
  OR2_X1 U116 ( .A1(n209), .A2(b[0]), .ZN(n116) );
  OR2_X1 U117 ( .A1(n201), .A2(a[0]), .ZN(n117) );
  AND2_X1 U118 ( .A1(n114), .A2(n113), .ZN(n115) );
  OR2_X1 U119 ( .A1(n185), .A2(d[0]), .ZN(n113) );
  OR2_X1 U120 ( .A1(n177), .A2(c[0]), .ZN(n114) );
endmodule


module byteXor4_10 ( a, b, c, d, y );
  input [7:0] a;
  input [7:0] b;
  input [7:0] c;
  input [7:0] d;
  //input_done

  output [7:0] y;
  //output_done

  wire   n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224;
  //wire_done

  INV_X1 U1 ( .A(n175), .ZN(n224) );
  INV_X1 U2 ( .A(a[7]), .ZN(n223) );
  INV_X1 U3 ( .A(n167), .ZN(n222) );
  INV_X1 U4 ( .A(a[6]), .ZN(n221) );
  INV_X1 U5 ( .A(n159), .ZN(n220) );
  INV_X1 U6 ( .A(a[5]), .ZN(n219) );
  INV_X1 U7 ( .A(n151), .ZN(n218) );
  INV_X1 U8 ( .A(a[4]), .ZN(n217) );
  INV_X1 U9 ( .A(n143), .ZN(n216) );
  INV_X1 U10 ( .A(a[3]), .ZN(n215) );
  INV_X1 U11 ( .A(n135), .ZN(n214) );
  INV_X1 U12 ( .A(a[2]), .ZN(n213) );
  INV_X1 U13 ( .A(n127), .ZN(n212) );
  INV_X1 U14 ( .A(a[1]), .ZN(n211) );
  INV_X1 U15 ( .A(n119), .ZN(n210) );
  INV_X1 U16 ( .A(a[0]), .ZN(n209) );
  INV_X1 U17 ( .A(b[7]), .ZN(n208) );
  INV_X1 U18 ( .A(b[6]), .ZN(n207) );
  INV_X1 U19 ( .A(b[5]), .ZN(n206) );
  INV_X1 U20 ( .A(b[4]), .ZN(n205) );
  INV_X1 U21 ( .A(b[3]), .ZN(n204) );
  INV_X1 U22 ( .A(b[2]), .ZN(n203) );
  INV_X1 U23 ( .A(b[1]), .ZN(n202) );
  INV_X1 U24 ( .A(b[0]), .ZN(n201) );
  INV_X1 U25 ( .A(n171), .ZN(n200) );
  INV_X1 U26 ( .A(c[7]), .ZN(n199) );
  INV_X1 U27 ( .A(n163), .ZN(n198) );
  INV_X1 U28 ( .A(c[6]), .ZN(n197) );
  INV_X1 U29 ( .A(n155), .ZN(n196) );
  INV_X1 U30 ( .A(c[5]), .ZN(n195) );
  INV_X1 U31 ( .A(n147), .ZN(n194) );
  INV_X1 U32 ( .A(c[4]), .ZN(n193) );
  INV_X1 U33 ( .A(n139), .ZN(n192) );
  INV_X1 U34 ( .A(c[3]), .ZN(n191) );
  INV_X1 U35 ( .A(n131), .ZN(n190) );
  INV_X1 U36 ( .A(c[2]), .ZN(n189) );
  INV_X1 U37 ( .A(n123), .ZN(n188) );
  INV_X1 U38 ( .A(c[1]), .ZN(n187) );
  INV_X1 U39 ( .A(n115), .ZN(n186) );
  INV_X1 U40 ( .A(c[0]), .ZN(n185) );
  INV_X1 U41 ( .A(d[7]), .ZN(n184) );
  INV_X1 U42 ( .A(d[6]), .ZN(n183) );
  INV_X1 U43 ( .A(d[5]), .ZN(n182) );
  INV_X1 U44 ( .A(d[4]), .ZN(n181) );
  INV_X1 U45 ( .A(d[3]), .ZN(n180) );
  INV_X1 U46 ( .A(d[2]), .ZN(n179) );
  INV_X1 U47 ( .A(d[1]), .ZN(n178) );
  INV_X1 U48 ( .A(d[0]), .ZN(n177) );
  OR2_X1 U49 ( .A1(n176), .A2(n224), .ZN(y[7]) );
  OR2_X1 U50 ( .A1(n174), .A2(n200), .ZN(n175) );
  AND2_X1 U51 ( .A1(n200), .A2(n174), .ZN(n176) );
  AND2_X1 U52 ( .A1(n173), .A2(n172), .ZN(n174) );
  OR2_X1 U53 ( .A1(n223), .A2(b[7]), .ZN(n172) );
  OR2_X1 U54 ( .A1(n208), .A2(a[7]), .ZN(n173) );
  AND2_X1 U55 ( .A1(n170), .A2(n169), .ZN(n171) );
  OR2_X1 U56 ( .A1(n199), .A2(d[7]), .ZN(n169) );
  OR2_X1 U57 ( .A1(n184), .A2(c[7]), .ZN(n170) );
  OR2_X1 U58 ( .A1(n168), .A2(n222), .ZN(y[6]) );
  OR2_X1 U59 ( .A1(n166), .A2(n198), .ZN(n167) );
  AND2_X1 U60 ( .A1(n198), .A2(n166), .ZN(n168) );
  AND2_X1 U61 ( .A1(n165), .A2(n164), .ZN(n166) );
  OR2_X1 U62 ( .A1(n221), .A2(b[6]), .ZN(n164) );
  OR2_X1 U63 ( .A1(n207), .A2(a[6]), .ZN(n165) );
  AND2_X1 U64 ( .A1(n162), .A2(n161), .ZN(n163) );
  OR2_X1 U65 ( .A1(n197), .A2(d[6]), .ZN(n161) );
  OR2_X1 U66 ( .A1(n183), .A2(c[6]), .ZN(n162) );
  OR2_X1 U67 ( .A1(n160), .A2(n220), .ZN(y[5]) );
  OR2_X1 U68 ( .A1(n158), .A2(n196), .ZN(n159) );
  AND2_X1 U69 ( .A1(n196), .A2(n158), .ZN(n160) );
  AND2_X1 U70 ( .A1(n157), .A2(n156), .ZN(n158) );
  OR2_X1 U71 ( .A1(n219), .A2(b[5]), .ZN(n156) );
  OR2_X1 U72 ( .A1(n206), .A2(a[5]), .ZN(n157) );
  AND2_X1 U73 ( .A1(n154), .A2(n153), .ZN(n155) );
  OR2_X1 U74 ( .A1(n195), .A2(d[5]), .ZN(n153) );
  OR2_X1 U75 ( .A1(n182), .A2(c[5]), .ZN(n154) );
  OR2_X1 U76 ( .A1(n152), .A2(n218), .ZN(y[4]) );
  OR2_X1 U77 ( .A1(n150), .A2(n194), .ZN(n151) );
  AND2_X1 U78 ( .A1(n194), .A2(n150), .ZN(n152) );
  AND2_X1 U79 ( .A1(n149), .A2(n148), .ZN(n150) );
  OR2_X1 U80 ( .A1(n217), .A2(b[4]), .ZN(n148) );
  OR2_X1 U81 ( .A1(n205), .A2(a[4]), .ZN(n149) );
  AND2_X1 U82 ( .A1(n146), .A2(n145), .ZN(n147) );
  OR2_X1 U83 ( .A1(n193), .A2(d[4]), .ZN(n145) );
  OR2_X1 U84 ( .A1(n181), .A2(c[4]), .ZN(n146) );
  OR2_X1 U85 ( .A1(n144), .A2(n216), .ZN(y[3]) );
  OR2_X1 U86 ( .A1(n142), .A2(n192), .ZN(n143) );
  AND2_X1 U87 ( .A1(n192), .A2(n142), .ZN(n144) );
  AND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(n142) );
  OR2_X1 U89 ( .A1(n215), .A2(b[3]), .ZN(n140) );
  OR2_X1 U90 ( .A1(n204), .A2(a[3]), .ZN(n141) );
  AND2_X1 U91 ( .A1(n138), .A2(n137), .ZN(n139) );
  OR2_X1 U92 ( .A1(n191), .A2(d[3]), .ZN(n137) );
  OR2_X1 U93 ( .A1(n180), .A2(c[3]), .ZN(n138) );
  OR2_X1 U94 ( .A1(n136), .A2(n214), .ZN(y[2]) );
  OR2_X1 U95 ( .A1(n134), .A2(n190), .ZN(n135) );
  AND2_X1 U96 ( .A1(n190), .A2(n134), .ZN(n136) );
  AND2_X1 U97 ( .A1(n133), .A2(n132), .ZN(n134) );
  OR2_X1 U98 ( .A1(n213), .A2(b[2]), .ZN(n132) );
  OR2_X1 U99 ( .A1(n203), .A2(a[2]), .ZN(n133) );
  AND2_X1 U100 ( .A1(n130), .A2(n129), .ZN(n131) );
  OR2_X1 U101 ( .A1(n189), .A2(d[2]), .ZN(n129) );
  OR2_X1 U102 ( .A1(n179), .A2(c[2]), .ZN(n130) );
  OR2_X1 U103 ( .A1(n128), .A2(n212), .ZN(y[1]) );
  OR2_X1 U104 ( .A1(n126), .A2(n188), .ZN(n127) );
  AND2_X1 U105 ( .A1(n188), .A2(n126), .ZN(n128) );
  AND2_X1 U106 ( .A1(n125), .A2(n124), .ZN(n126) );
  OR2_X1 U107 ( .A1(n211), .A2(b[1]), .ZN(n124) );
  OR2_X1 U108 ( .A1(n202), .A2(a[1]), .ZN(n125) );
  AND2_X1 U109 ( .A1(n122), .A2(n121), .ZN(n123) );
  OR2_X1 U110 ( .A1(n187), .A2(d[1]), .ZN(n121) );
  OR2_X1 U111 ( .A1(n178), .A2(c[1]), .ZN(n122) );
  OR2_X1 U112 ( .A1(n120), .A2(n210), .ZN(y[0]) );
  OR2_X1 U113 ( .A1(n118), .A2(n186), .ZN(n119) );
  AND2_X1 U114 ( .A1(n186), .A2(n118), .ZN(n120) );
  AND2_X1 U115 ( .A1(n117), .A2(n116), .ZN(n118) );
  OR2_X1 U116 ( .A1(n209), .A2(b[0]), .ZN(n116) );
  OR2_X1 U117 ( .A1(n201), .A2(a[0]), .ZN(n117) );
  AND2_X1 U118 ( .A1(n114), .A2(n113), .ZN(n115) );
  OR2_X1 U119 ( .A1(n185), .A2(d[0]), .ZN(n113) );
  OR2_X1 U120 ( .A1(n177), .A2(c[0]), .ZN(n114) );
endmodule


module byteXor4_11 ( a, b, c, d, y );
  input [7:0] a;
  input [7:0] b;
  input [7:0] c;
  input [7:0] d;
  //input_done

  output [7:0] y;
  //output_done

  wire   n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224;
  //wire_done

  INV_X1 U1 ( .A(n175), .ZN(n224) );
  INV_X1 U2 ( .A(a[7]), .ZN(n223) );
  INV_X1 U3 ( .A(n167), .ZN(n222) );
  INV_X1 U4 ( .A(a[6]), .ZN(n221) );
  INV_X1 U5 ( .A(n159), .ZN(n220) );
  INV_X1 U6 ( .A(a[5]), .ZN(n219) );
  INV_X1 U7 ( .A(n151), .ZN(n218) );
  INV_X1 U8 ( .A(a[4]), .ZN(n217) );
  INV_X1 U9 ( .A(n143), .ZN(n216) );
  INV_X1 U10 ( .A(a[3]), .ZN(n215) );
  INV_X1 U11 ( .A(n135), .ZN(n214) );
  INV_X1 U12 ( .A(a[2]), .ZN(n213) );
  INV_X1 U13 ( .A(n127), .ZN(n212) );
  INV_X1 U14 ( .A(a[1]), .ZN(n211) );
  INV_X1 U15 ( .A(n119), .ZN(n210) );
  INV_X1 U16 ( .A(a[0]), .ZN(n209) );
  INV_X1 U17 ( .A(b[7]), .ZN(n208) );
  INV_X1 U18 ( .A(b[6]), .ZN(n207) );
  INV_X1 U19 ( .A(b[5]), .ZN(n206) );
  INV_X1 U20 ( .A(b[4]), .ZN(n205) );
  INV_X1 U21 ( .A(b[3]), .ZN(n204) );
  INV_X1 U22 ( .A(b[2]), .ZN(n203) );
  INV_X1 U23 ( .A(b[1]), .ZN(n202) );
  INV_X1 U24 ( .A(b[0]), .ZN(n201) );
  INV_X1 U25 ( .A(n171), .ZN(n200) );
  INV_X1 U26 ( .A(c[7]), .ZN(n199) );
  INV_X1 U27 ( .A(n163), .ZN(n198) );
  INV_X1 U28 ( .A(c[6]), .ZN(n197) );
  INV_X1 U29 ( .A(n155), .ZN(n196) );
  INV_X1 U30 ( .A(c[5]), .ZN(n195) );
  INV_X1 U31 ( .A(n147), .ZN(n194) );
  INV_X1 U32 ( .A(c[4]), .ZN(n193) );
  INV_X1 U33 ( .A(n139), .ZN(n192) );
  INV_X1 U34 ( .A(c[3]), .ZN(n191) );
  INV_X1 U35 ( .A(n131), .ZN(n190) );
  INV_X1 U36 ( .A(c[2]), .ZN(n189) );
  INV_X1 U37 ( .A(n123), .ZN(n188) );
  INV_X1 U38 ( .A(c[1]), .ZN(n187) );
  INV_X1 U39 ( .A(n115), .ZN(n186) );
  INV_X1 U40 ( .A(c[0]), .ZN(n185) );
  INV_X1 U41 ( .A(d[7]), .ZN(n184) );
  INV_X1 U42 ( .A(d[6]), .ZN(n183) );
  INV_X1 U43 ( .A(d[5]), .ZN(n182) );
  INV_X1 U44 ( .A(d[4]), .ZN(n181) );
  INV_X1 U45 ( .A(d[3]), .ZN(n180) );
  INV_X1 U46 ( .A(d[2]), .ZN(n179) );
  INV_X1 U47 ( .A(d[1]), .ZN(n178) );
  INV_X1 U48 ( .A(d[0]), .ZN(n177) );
  OR2_X1 U49 ( .A1(n176), .A2(n224), .ZN(y[7]) );
  OR2_X1 U50 ( .A1(n174), .A2(n200), .ZN(n175) );
  AND2_X1 U51 ( .A1(n200), .A2(n174), .ZN(n176) );
  AND2_X1 U52 ( .A1(n173), .A2(n172), .ZN(n174) );
  OR2_X1 U53 ( .A1(n223), .A2(b[7]), .ZN(n172) );
  OR2_X1 U54 ( .A1(n208), .A2(a[7]), .ZN(n173) );
  AND2_X1 U55 ( .A1(n170), .A2(n169), .ZN(n171) );
  OR2_X1 U56 ( .A1(n199), .A2(d[7]), .ZN(n169) );
  OR2_X1 U57 ( .A1(n184), .A2(c[7]), .ZN(n170) );
  OR2_X1 U58 ( .A1(n168), .A2(n222), .ZN(y[6]) );
  OR2_X1 U59 ( .A1(n166), .A2(n198), .ZN(n167) );
  AND2_X1 U60 ( .A1(n198), .A2(n166), .ZN(n168) );
  AND2_X1 U61 ( .A1(n165), .A2(n164), .ZN(n166) );
  OR2_X1 U62 ( .A1(n221), .A2(b[6]), .ZN(n164) );
  OR2_X1 U63 ( .A1(n207), .A2(a[6]), .ZN(n165) );
  AND2_X1 U64 ( .A1(n162), .A2(n161), .ZN(n163) );
  OR2_X1 U65 ( .A1(n197), .A2(d[6]), .ZN(n161) );
  OR2_X1 U66 ( .A1(n183), .A2(c[6]), .ZN(n162) );
  OR2_X1 U67 ( .A1(n160), .A2(n220), .ZN(y[5]) );
  OR2_X1 U68 ( .A1(n158), .A2(n196), .ZN(n159) );
  AND2_X1 U69 ( .A1(n196), .A2(n158), .ZN(n160) );
  AND2_X1 U70 ( .A1(n157), .A2(n156), .ZN(n158) );
  OR2_X1 U71 ( .A1(n219), .A2(b[5]), .ZN(n156) );
  OR2_X1 U72 ( .A1(n206), .A2(a[5]), .ZN(n157) );
  AND2_X1 U73 ( .A1(n154), .A2(n153), .ZN(n155) );
  OR2_X1 U74 ( .A1(n195), .A2(d[5]), .ZN(n153) );
  OR2_X1 U75 ( .A1(n182), .A2(c[5]), .ZN(n154) );
  OR2_X1 U76 ( .A1(n152), .A2(n218), .ZN(y[4]) );
  OR2_X1 U77 ( .A1(n150), .A2(n194), .ZN(n151) );
  AND2_X1 U78 ( .A1(n194), .A2(n150), .ZN(n152) );
  AND2_X1 U79 ( .A1(n149), .A2(n148), .ZN(n150) );
  OR2_X1 U80 ( .A1(n217), .A2(b[4]), .ZN(n148) );
  OR2_X1 U81 ( .A1(n205), .A2(a[4]), .ZN(n149) );
  AND2_X1 U82 ( .A1(n146), .A2(n145), .ZN(n147) );
  OR2_X1 U83 ( .A1(n193), .A2(d[4]), .ZN(n145) );
  OR2_X1 U84 ( .A1(n181), .A2(c[4]), .ZN(n146) );
  OR2_X1 U85 ( .A1(n144), .A2(n216), .ZN(y[3]) );
  OR2_X1 U86 ( .A1(n142), .A2(n192), .ZN(n143) );
  AND2_X1 U87 ( .A1(n192), .A2(n142), .ZN(n144) );
  AND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(n142) );
  OR2_X1 U89 ( .A1(n215), .A2(b[3]), .ZN(n140) );
  OR2_X1 U90 ( .A1(n204), .A2(a[3]), .ZN(n141) );
  AND2_X1 U91 ( .A1(n138), .A2(n137), .ZN(n139) );
  OR2_X1 U92 ( .A1(n191), .A2(d[3]), .ZN(n137) );
  OR2_X1 U93 ( .A1(n180), .A2(c[3]), .ZN(n138) );
  OR2_X1 U94 ( .A1(n136), .A2(n214), .ZN(y[2]) );
  OR2_X1 U95 ( .A1(n134), .A2(n190), .ZN(n135) );
  AND2_X1 U96 ( .A1(n190), .A2(n134), .ZN(n136) );
  AND2_X1 U97 ( .A1(n133), .A2(n132), .ZN(n134) );
  OR2_X1 U98 ( .A1(n213), .A2(b[2]), .ZN(n132) );
  OR2_X1 U99 ( .A1(n203), .A2(a[2]), .ZN(n133) );
  AND2_X1 U100 ( .A1(n130), .A2(n129), .ZN(n131) );
  OR2_X1 U101 ( .A1(n189), .A2(d[2]), .ZN(n129) );
  OR2_X1 U102 ( .A1(n179), .A2(c[2]), .ZN(n130) );
  OR2_X1 U103 ( .A1(n128), .A2(n212), .ZN(y[1]) );
  OR2_X1 U104 ( .A1(n126), .A2(n188), .ZN(n127) );
  AND2_X1 U105 ( .A1(n188), .A2(n126), .ZN(n128) );
  AND2_X1 U106 ( .A1(n125), .A2(n124), .ZN(n126) );
  OR2_X1 U107 ( .A1(n211), .A2(b[1]), .ZN(n124) );
  OR2_X1 U108 ( .A1(n202), .A2(a[1]), .ZN(n125) );
  AND2_X1 U109 ( .A1(n122), .A2(n121), .ZN(n123) );
  OR2_X1 U110 ( .A1(n187), .A2(d[1]), .ZN(n121) );
  OR2_X1 U111 ( .A1(n178), .A2(c[1]), .ZN(n122) );
  OR2_X1 U112 ( .A1(n120), .A2(n210), .ZN(y[0]) );
  OR2_X1 U113 ( .A1(n118), .A2(n186), .ZN(n119) );
  AND2_X1 U114 ( .A1(n186), .A2(n118), .ZN(n120) );
  AND2_X1 U115 ( .A1(n117), .A2(n116), .ZN(n118) );
  OR2_X1 U116 ( .A1(n209), .A2(b[0]), .ZN(n116) );
  OR2_X1 U117 ( .A1(n201), .A2(a[0]), .ZN(n117) );
  AND2_X1 U118 ( .A1(n114), .A2(n113), .ZN(n115) );
  OR2_X1 U119 ( .A1(n185), .A2(d[0]), .ZN(n113) );
  OR2_X1 U120 ( .A1(n177), .A2(c[0]), .ZN(n114) );
endmodule


module byteXor4_12 ( a, b, c, d, y );
  input [7:0] a;
  input [7:0] b;
  input [7:0] c;
  input [7:0] d;
  //input_done

  output [7:0] y;
  //output_done

  wire   n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224;
  //wire_done

  INV_X1 U1 ( .A(n175), .ZN(n224) );
  INV_X1 U2 ( .A(a[7]), .ZN(n223) );
  INV_X1 U3 ( .A(n167), .ZN(n222) );
  INV_X1 U4 ( .A(a[6]), .ZN(n221) );
  INV_X1 U5 ( .A(n159), .ZN(n220) );
  INV_X1 U6 ( .A(a[5]), .ZN(n219) );
  INV_X1 U7 ( .A(n151), .ZN(n218) );
  INV_X1 U8 ( .A(a[4]), .ZN(n217) );
  INV_X1 U9 ( .A(n143), .ZN(n216) );
  INV_X1 U10 ( .A(a[3]), .ZN(n215) );
  INV_X1 U11 ( .A(n135), .ZN(n214) );
  INV_X1 U12 ( .A(a[2]), .ZN(n213) );
  INV_X1 U13 ( .A(n127), .ZN(n212) );
  INV_X1 U14 ( .A(a[1]), .ZN(n211) );
  INV_X1 U15 ( .A(n119), .ZN(n210) );
  INV_X1 U16 ( .A(a[0]), .ZN(n209) );
  INV_X1 U17 ( .A(b[7]), .ZN(n208) );
  INV_X1 U18 ( .A(b[6]), .ZN(n207) );
  INV_X1 U19 ( .A(b[5]), .ZN(n206) );
  INV_X1 U20 ( .A(b[4]), .ZN(n205) );
  INV_X1 U21 ( .A(b[3]), .ZN(n204) );
  INV_X1 U22 ( .A(b[2]), .ZN(n203) );
  INV_X1 U23 ( .A(b[1]), .ZN(n202) );
  INV_X1 U24 ( .A(b[0]), .ZN(n201) );
  INV_X1 U25 ( .A(n171), .ZN(n200) );
  INV_X1 U26 ( .A(c[7]), .ZN(n199) );
  INV_X1 U27 ( .A(n163), .ZN(n198) );
  INV_X1 U28 ( .A(c[6]), .ZN(n197) );
  INV_X1 U29 ( .A(n155), .ZN(n196) );
  INV_X1 U30 ( .A(c[5]), .ZN(n195) );
  INV_X1 U31 ( .A(n147), .ZN(n194) );
  INV_X1 U32 ( .A(c[4]), .ZN(n193) );
  INV_X1 U33 ( .A(n139), .ZN(n192) );
  INV_X1 U34 ( .A(c[3]), .ZN(n191) );
  INV_X1 U35 ( .A(n131), .ZN(n190) );
  INV_X1 U36 ( .A(c[2]), .ZN(n189) );
  INV_X1 U37 ( .A(n123), .ZN(n188) );
  INV_X1 U38 ( .A(c[1]), .ZN(n187) );
  INV_X1 U39 ( .A(n115), .ZN(n186) );
  INV_X1 U40 ( .A(c[0]), .ZN(n185) );
  INV_X1 U41 ( .A(d[7]), .ZN(n184) );
  INV_X1 U42 ( .A(d[6]), .ZN(n183) );
  INV_X1 U43 ( .A(d[5]), .ZN(n182) );
  INV_X1 U44 ( .A(d[4]), .ZN(n181) );
  INV_X1 U45 ( .A(d[3]), .ZN(n180) );
  INV_X1 U46 ( .A(d[2]), .ZN(n179) );
  INV_X1 U47 ( .A(d[1]), .ZN(n178) );
  INV_X1 U48 ( .A(d[0]), .ZN(n177) );
  OR2_X1 U49 ( .A1(n176), .A2(n224), .ZN(y[7]) );
  OR2_X1 U50 ( .A1(n174), .A2(n200), .ZN(n175) );
  AND2_X1 U51 ( .A1(n200), .A2(n174), .ZN(n176) );
  AND2_X1 U52 ( .A1(n173), .A2(n172), .ZN(n174) );
  OR2_X1 U53 ( .A1(n223), .A2(b[7]), .ZN(n172) );
  OR2_X1 U54 ( .A1(n208), .A2(a[7]), .ZN(n173) );
  AND2_X1 U55 ( .A1(n170), .A2(n169), .ZN(n171) );
  OR2_X1 U56 ( .A1(n199), .A2(d[7]), .ZN(n169) );
  OR2_X1 U57 ( .A1(n184), .A2(c[7]), .ZN(n170) );
  OR2_X1 U58 ( .A1(n168), .A2(n222), .ZN(y[6]) );
  OR2_X1 U59 ( .A1(n166), .A2(n198), .ZN(n167) );
  AND2_X1 U60 ( .A1(n198), .A2(n166), .ZN(n168) );
  AND2_X1 U61 ( .A1(n165), .A2(n164), .ZN(n166) );
  OR2_X1 U62 ( .A1(n221), .A2(b[6]), .ZN(n164) );
  OR2_X1 U63 ( .A1(n207), .A2(a[6]), .ZN(n165) );
  AND2_X1 U64 ( .A1(n162), .A2(n161), .ZN(n163) );
  OR2_X1 U65 ( .A1(n197), .A2(d[6]), .ZN(n161) );
  OR2_X1 U66 ( .A1(n183), .A2(c[6]), .ZN(n162) );
  OR2_X1 U67 ( .A1(n160), .A2(n220), .ZN(y[5]) );
  OR2_X1 U68 ( .A1(n158), .A2(n196), .ZN(n159) );
  AND2_X1 U69 ( .A1(n196), .A2(n158), .ZN(n160) );
  AND2_X1 U70 ( .A1(n157), .A2(n156), .ZN(n158) );
  OR2_X1 U71 ( .A1(n219), .A2(b[5]), .ZN(n156) );
  OR2_X1 U72 ( .A1(n206), .A2(a[5]), .ZN(n157) );
  AND2_X1 U73 ( .A1(n154), .A2(n153), .ZN(n155) );
  OR2_X1 U74 ( .A1(n195), .A2(d[5]), .ZN(n153) );
  OR2_X1 U75 ( .A1(n182), .A2(c[5]), .ZN(n154) );
  OR2_X1 U76 ( .A1(n152), .A2(n218), .ZN(y[4]) );
  OR2_X1 U77 ( .A1(n150), .A2(n194), .ZN(n151) );
  AND2_X1 U78 ( .A1(n194), .A2(n150), .ZN(n152) );
  AND2_X1 U79 ( .A1(n149), .A2(n148), .ZN(n150) );
  OR2_X1 U80 ( .A1(n217), .A2(b[4]), .ZN(n148) );
  OR2_X1 U81 ( .A1(n205), .A2(a[4]), .ZN(n149) );
  AND2_X1 U82 ( .A1(n146), .A2(n145), .ZN(n147) );
  OR2_X1 U83 ( .A1(n193), .A2(d[4]), .ZN(n145) );
  OR2_X1 U84 ( .A1(n181), .A2(c[4]), .ZN(n146) );
  OR2_X1 U85 ( .A1(n144), .A2(n216), .ZN(y[3]) );
  OR2_X1 U86 ( .A1(n142), .A2(n192), .ZN(n143) );
  AND2_X1 U87 ( .A1(n192), .A2(n142), .ZN(n144) );
  AND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(n142) );
  OR2_X1 U89 ( .A1(n215), .A2(b[3]), .ZN(n140) );
  OR2_X1 U90 ( .A1(n204), .A2(a[3]), .ZN(n141) );
  AND2_X1 U91 ( .A1(n138), .A2(n137), .ZN(n139) );
  OR2_X1 U92 ( .A1(n191), .A2(d[3]), .ZN(n137) );
  OR2_X1 U93 ( .A1(n180), .A2(c[3]), .ZN(n138) );
  OR2_X1 U94 ( .A1(n136), .A2(n214), .ZN(y[2]) );
  OR2_X1 U95 ( .A1(n134), .A2(n190), .ZN(n135) );
  AND2_X1 U96 ( .A1(n190), .A2(n134), .ZN(n136) );
  AND2_X1 U97 ( .A1(n133), .A2(n132), .ZN(n134) );
  OR2_X1 U98 ( .A1(n213), .A2(b[2]), .ZN(n132) );
  OR2_X1 U99 ( .A1(n203), .A2(a[2]), .ZN(n133) );
  AND2_X1 U100 ( .A1(n130), .A2(n129), .ZN(n131) );
  OR2_X1 U101 ( .A1(n189), .A2(d[2]), .ZN(n129) );
  OR2_X1 U102 ( .A1(n179), .A2(c[2]), .ZN(n130) );
  OR2_X1 U103 ( .A1(n128), .A2(n212), .ZN(y[1]) );
  OR2_X1 U104 ( .A1(n126), .A2(n188), .ZN(n127) );
  AND2_X1 U105 ( .A1(n188), .A2(n126), .ZN(n128) );
  AND2_X1 U106 ( .A1(n125), .A2(n124), .ZN(n126) );
  OR2_X1 U107 ( .A1(n211), .A2(b[1]), .ZN(n124) );
  OR2_X1 U108 ( .A1(n202), .A2(a[1]), .ZN(n125) );
  AND2_X1 U109 ( .A1(n122), .A2(n121), .ZN(n123) );
  OR2_X1 U110 ( .A1(n187), .A2(d[1]), .ZN(n121) );
  OR2_X1 U111 ( .A1(n178), .A2(c[1]), .ZN(n122) );
  OR2_X1 U112 ( .A1(n120), .A2(n210), .ZN(y[0]) );
  OR2_X1 U113 ( .A1(n118), .A2(n186), .ZN(n119) );
  AND2_X1 U114 ( .A1(n186), .A2(n118), .ZN(n120) );
  AND2_X1 U115 ( .A1(n117), .A2(n116), .ZN(n118) );
  OR2_X1 U116 ( .A1(n209), .A2(b[0]), .ZN(n116) );
  OR2_X1 U117 ( .A1(n201), .A2(a[0]), .ZN(n117) );
  AND2_X1 U118 ( .A1(n114), .A2(n113), .ZN(n115) );
  OR2_X1 U119 ( .A1(n185), .A2(d[0]), .ZN(n113) );
  OR2_X1 U120 ( .A1(n177), .A2(c[0]), .ZN(n114) );
endmodule


module mixCol_3 ( in, out );
  input [31:0] in;
  //input_done

  output [31:0] out;
  //output_done

  wire   [7:0] b0_s2;
  wire   [7:0] b1_s2;
  wire   [7:0] b2_s2;
  wire   [7:0] b3_s2;
  wire   [7:0] b0_s3;
  wire   [7:0] b1_s3;
  wire   [7:0] b2_s3;
  wire   [7:0] b3_s3;
  //wire_done

  scale2_12 b0_scale2 ( .in(in[31:24]), .out(b0_s2) );
  scale2_11 b1_scale2 ( .in(in[23:16]), .out(b1_s2) );
  scale2_10 b2_scale2 ( .in(in[15:8]), .out(b2_s2) );
  scale2_9 b3_scale2 ( .in(in[7:0]), .out(b3_s2) );
  byteXor_13 b0_scale3 ( .a(in[31:24]), .b(b0_s2), .y(b0_s3) );
  byteXor_12 b1_scale3 ( .a(in[23:16]), .b(b1_s2), .y(b1_s3) );
  byteXor_11 b2_scale3 ( .a(in[15:8]), .b(b2_s2), .y(b2_s3) );
  byteXor_10 b3_scale3 ( .a(in[7:0]), .b(b3_s2), .y(b3_s3) );
  byteXor4_12 out0 ( .a(b0_s2), .b(b1_s3), .c(in[15:8]), .d(in[7:0]), .y(
        out[31:24]) );
  byteXor4_11 out1 ( .a(in[31:24]), .b(b1_s2), .c(b2_s3), .d(in[7:0]), .y(
        out[23:16]) );
  byteXor4_10 out2 ( .a(in[31:24]), .b(in[23:16]), .c(b2_s2), .d(b3_s3), .y(
        out[15:8]) );
  byteXor4_9 out3 ( .a(b0_s3), .b(in[23:16]), .c(in[15:8]), .d(b3_s2), .y(
        out[7:0]) );
endmodule


module aes_128 ( clk, data, key, firstRound, final_round, round_const, out );
  input [127:0] data;
  input [127:0] key;
  input [7:0] round_const;
  input clk, firstRound, final_round;
  //input_done

  output [127:0] out;
  //output_done
  
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773;
  wire   [127:0] state;
  wire   [127:0] data_in;
  wire   [127:0] addKey_out;
  wire   [127:0] sr_out;
  wire   [127:0] sBox_out;
  wire   [127:0] mixCol_out_temp;
  wire   [127:0] mixCol_out;
  wire   [127:0] key_out;
  //wire_done

  mux128_0 dataMux ( .a(out), .b(state), .sel(firstRound), .y(data_in) );
  shiftRows sr ( .in(data_in), .out(sr_out) );
  sBox_0 s0 ( .in(sr_out[127:120]), .out(sBox_out[127:120]) );
  sBox_19 s1 ( .in(sr_out[119:112]), .out(sBox_out[119:112]) );
  sBox_18 s2 ( .in(sr_out[111:104]), .out(sBox_out[111:104]) );
  sBox_17 s3 ( .in(sr_out[103:96]), .out(sBox_out[103:96]) );
  sBox_16 s4 ( .in(sr_out[95:88]), .out(sBox_out[95:88]) );
  sBox_15 s5 ( .in(sr_out[87:80]), .out(sBox_out[87:80]) );
  sBox_14 s6 ( .in(sr_out[79:72]), .out(sBox_out[79:72]) );
  sBox_13 s7 ( .in(sr_out[71:64]), .out(sBox_out[71:64]) );
  sBox_12 s8 ( .in(sr_out[63:56]), .out(sBox_out[63:56]) );
  sBox_11 s9 ( .in(sr_out[55:48]), .out(sBox_out[55:48]) );
  sBox_10 s10 ( .in(sr_out[47:40]), .out(sBox_out[47:40]) );
  sBox_9 s11 ( .in(sr_out[39:32]), .out(sBox_out[39:32]) );
  sBox_8 s12 ( .in(sr_out[31:24]), .out(sBox_out[31:24]) );
  sBox_7 s13 ( .in(sr_out[23:16]), .out(sBox_out[23:16]) );
  sBox_6 s14 ( .in(sr_out[15:8]), .out(sBox_out[15:8]) );
  sBox_5 s15 ( .in(sr_out[7:0]), .out(sBox_out[7:0]) );
  mixCol_0 mc0 ( .in(sBox_out[127:96]), .out(mixCol_out_temp[127:96]) );
  mixCol_3 mc1 ( .in(sBox_out[95:64]), .out(mixCol_out_temp[95:64]) );
  mixCol_2 mc2 ( .in(sBox_out[63:32]), .out(mixCol_out_temp[63:32]) );
  mixCol_1 mc3 ( .in(sBox_out[31:0]), .out(mixCol_out_temp[31:0]) );
  keyExpansion ke ( .key_in(key), .clk(clk), .firstRound(firstRound), 
        .round_const(round_const), .key_out(key_out) );
  addKey ak0 ( .data(mixCol_out), .key(key_out), .out(addKey_out) );
  DFF_X1 \out_reg[0]  ( .D(addKey_out[0]), .CK(clk), .Q(out[0]) );
  DFF_X1 \out_reg[1]  ( .D(addKey_out[1]), .CK(clk), .Q(out[1]) );
  DFF_X1 \out_reg[2]  ( .D(addKey_out[2]), .CK(clk), .Q(out[2]) );
  DFF_X1 \out_reg[3]  ( .D(addKey_out[3]), .CK(clk), .Q(out[3]) );
  DFF_X1 \out_reg[4]  ( .D(addKey_out[4]), .CK(clk), .Q(out[4]) );
  DFF_X1 \out_reg[5]  ( .D(addKey_out[5]), .CK(clk), .Q(out[5]) );
  DFF_X1 \out_reg[6]  ( .D(addKey_out[6]), .CK(clk), .Q(out[6]) );
  DFF_X1 \out_reg[7]  ( .D(addKey_out[7]), .CK(clk), .Q(out[7]) );
  DFF_X1 \out_reg[8]  ( .D(addKey_out[8]), .CK(clk), .Q(out[8]) );
  DFF_X1 \out_reg[9]  ( .D(addKey_out[9]), .CK(clk), .Q(out[9]) );
  DFF_X1 \out_reg[10]  ( .D(addKey_out[10]), .CK(clk), .Q(out[10]) );
  DFF_X1 \out_reg[11]  ( .D(addKey_out[11]), .CK(clk), .Q(out[11]) );
  DFF_X1 \out_reg[12]  ( .D(addKey_out[12]), .CK(clk), .Q(out[12]) );
  DFF_X1 \out_reg[13]  ( .D(addKey_out[13]), .CK(clk), .Q(out[13]) );
  DFF_X1 \out_reg[14]  ( .D(addKey_out[14]), .CK(clk), .Q(out[14]) );
  DFF_X1 \out_reg[15]  ( .D(addKey_out[15]), .CK(clk), .Q(out[15]) );
  DFF_X1 \out_reg[16]  ( .D(addKey_out[16]), .CK(clk), .Q(out[16]) );
  DFF_X1 \out_reg[17]  ( .D(addKey_out[17]), .CK(clk), .Q(out[17]) );
  DFF_X1 \out_reg[18]  ( .D(addKey_out[18]), .CK(clk), .Q(out[18]) );
  DFF_X1 \out_reg[19]  ( .D(addKey_out[19]), .CK(clk), .Q(out[19]) );
  DFF_X1 \out_reg[20]  ( .D(addKey_out[20]), .CK(clk), .Q(out[20]) );
  DFF_X1 \out_reg[21]  ( .D(addKey_out[21]), .CK(clk), .Q(out[21]) );
  DFF_X1 \out_reg[22]  ( .D(addKey_out[22]), .CK(clk), .Q(out[22]) );
  DFF_X1 \out_reg[23]  ( .D(addKey_out[23]), .CK(clk), .Q(out[23]) );
  DFF_X1 \out_reg[24]  ( .D(addKey_out[24]), .CK(clk), .Q(out[24]) );
  DFF_X1 \out_reg[25]  ( .D(addKey_out[25]), .CK(clk), .Q(out[25]) );
  DFF_X1 \out_reg[26]  ( .D(addKey_out[26]), .CK(clk), .Q(out[26]) );
  DFF_X1 \out_reg[27]  ( .D(addKey_out[27]), .CK(clk), .Q(out[27]) );
  DFF_X1 \out_reg[28]  ( .D(addKey_out[28]), .CK(clk), .Q(out[28]) );
  DFF_X1 \out_reg[29]  ( .D(addKey_out[29]), .CK(clk), .Q(out[29]) );
  DFF_X1 \out_reg[30]  ( .D(addKey_out[30]), .CK(clk), .Q(out[30]) );
  DFF_X1 \out_reg[31]  ( .D(addKey_out[31]), .CK(clk), .Q(out[31]) );
  DFF_X1 \out_reg[32]  ( .D(addKey_out[32]), .CK(clk), .Q(out[32]) );
  DFF_X1 \out_reg[33]  ( .D(addKey_out[33]), .CK(clk), .Q(out[33]) );
  DFF_X1 \out_reg[34]  ( .D(addKey_out[34]), .CK(clk), .Q(out[34]) );
  DFF_X1 \out_reg[35]  ( .D(addKey_out[35]), .CK(clk), .Q(out[35]) );
  DFF_X1 \out_reg[36]  ( .D(addKey_out[36]), .CK(clk), .Q(out[36]) );
  DFF_X1 \out_reg[37]  ( .D(addKey_out[37]), .CK(clk), .Q(out[37]) );
  DFF_X1 \out_reg[38]  ( .D(addKey_out[38]), .CK(clk), .Q(out[38]) );
  DFF_X1 \out_reg[39]  ( .D(addKey_out[39]), .CK(clk), .Q(out[39]) );
  DFF_X1 \out_reg[40]  ( .D(addKey_out[40]), .CK(clk), .Q(out[40]) );
  DFF_X1 \out_reg[41]  ( .D(addKey_out[41]), .CK(clk), .Q(out[41]) );
  DFF_X1 \out_reg[42]  ( .D(addKey_out[42]), .CK(clk), .Q(out[42]) );
  DFF_X1 \out_reg[43]  ( .D(addKey_out[43]), .CK(clk), .Q(out[43]) );
  DFF_X1 \out_reg[44]  ( .D(addKey_out[44]), .CK(clk), .Q(out[44]) );
  DFF_X1 \out_reg[45]  ( .D(addKey_out[45]), .CK(clk), .Q(out[45]) );
  DFF_X1 \out_reg[46]  ( .D(addKey_out[46]), .CK(clk), .Q(out[46]) );
  DFF_X1 \out_reg[47]  ( .D(addKey_out[47]), .CK(clk), .Q(out[47]) );
  DFF_X1 \out_reg[48]  ( .D(addKey_out[48]), .CK(clk), .Q(out[48]) );
  DFF_X1 \out_reg[49]  ( .D(addKey_out[49]), .CK(clk), .Q(out[49]) );
  DFF_X1 \out_reg[50]  ( .D(addKey_out[50]), .CK(clk), .Q(out[50]) );
  DFF_X1 \out_reg[51]  ( .D(addKey_out[51]), .CK(clk), .Q(out[51]) );
  DFF_X1 \out_reg[52]  ( .D(addKey_out[52]), .CK(clk), .Q(out[52]) );
  DFF_X1 \out_reg[53]  ( .D(addKey_out[53]), .CK(clk), .Q(out[53]) );
  DFF_X1 \out_reg[54]  ( .D(addKey_out[54]), .CK(clk), .Q(out[54]) );
  DFF_X1 \out_reg[55]  ( .D(addKey_out[55]), .CK(clk), .Q(out[55]) );
  DFF_X1 \out_reg[56]  ( .D(addKey_out[56]), .CK(clk), .Q(out[56]) );
  DFF_X1 \out_reg[57]  ( .D(addKey_out[57]), .CK(clk), .Q(out[57]) );
  DFF_X1 \out_reg[58]  ( .D(addKey_out[58]), .CK(clk), .Q(out[58]) );
  DFF_X1 \out_reg[59]  ( .D(addKey_out[59]), .CK(clk), .Q(out[59]) );
  DFF_X1 \out_reg[60]  ( .D(addKey_out[60]), .CK(clk), .Q(out[60]) );
  DFF_X1 \out_reg[61]  ( .D(addKey_out[61]), .CK(clk), .Q(out[61]) );
  DFF_X1 \out_reg[62]  ( .D(addKey_out[62]), .CK(clk), .Q(out[62]) );
  DFF_X1 \out_reg[63]  ( .D(addKey_out[63]), .CK(clk), .Q(out[63]) );
  DFF_X1 \out_reg[64]  ( .D(addKey_out[64]), .CK(clk), .Q(out[64]) );
  DFF_X1 \out_reg[65]  ( .D(addKey_out[65]), .CK(clk), .Q(out[65]) );
  DFF_X1 \out_reg[66]  ( .D(addKey_out[66]), .CK(clk), .Q(out[66]) );
  DFF_X1 \out_reg[67]  ( .D(addKey_out[67]), .CK(clk), .Q(out[67]) );
  DFF_X1 \out_reg[68]  ( .D(addKey_out[68]), .CK(clk), .Q(out[68]) );
  DFF_X1 \out_reg[69]  ( .D(addKey_out[69]), .CK(clk), .Q(out[69]) );
  DFF_X1 \out_reg[70]  ( .D(addKey_out[70]), .CK(clk), .Q(out[70]) );
  DFF_X1 \out_reg[71]  ( .D(addKey_out[71]), .CK(clk), .Q(out[71]) );
  DFF_X1 \out_reg[72]  ( .D(addKey_out[72]), .CK(clk), .Q(out[72]) );
  DFF_X1 \out_reg[73]  ( .D(addKey_out[73]), .CK(clk), .Q(out[73]) );
  DFF_X1 \out_reg[74]  ( .D(addKey_out[74]), .CK(clk), .Q(out[74]) );
  DFF_X1 \out_reg[75]  ( .D(addKey_out[75]), .CK(clk), .Q(out[75]) );
  DFF_X1 \out_reg[76]  ( .D(addKey_out[76]), .CK(clk), .Q(out[76]) );
  DFF_X1 \out_reg[77]  ( .D(addKey_out[77]), .CK(clk), .Q(out[77]) );
  DFF_X1 \out_reg[78]  ( .D(addKey_out[78]), .CK(clk), .Q(out[78]) );
  DFF_X1 \out_reg[79]  ( .D(addKey_out[79]), .CK(clk), .Q(out[79]) );
  DFF_X1 \out_reg[80]  ( .D(addKey_out[80]), .CK(clk), .Q(out[80]) );
  DFF_X1 \out_reg[81]  ( .D(addKey_out[81]), .CK(clk), .Q(out[81]) );
  DFF_X1 \out_reg[82]  ( .D(addKey_out[82]), .CK(clk), .Q(out[82]) );
  DFF_X1 \out_reg[83]  ( .D(addKey_out[83]), .CK(clk), .Q(out[83]) );
  DFF_X1 \out_reg[84]  ( .D(addKey_out[84]), .CK(clk), .Q(out[84]) );
  DFF_X1 \out_reg[85]  ( .D(addKey_out[85]), .CK(clk), .Q(out[85]) );
  DFF_X1 \out_reg[86]  ( .D(addKey_out[86]), .CK(clk), .Q(out[86]) );
  DFF_X1 \out_reg[87]  ( .D(addKey_out[87]), .CK(clk), .Q(out[87]) );
  DFF_X1 \out_reg[88]  ( .D(addKey_out[88]), .CK(clk), .Q(out[88]) );
  DFF_X1 \out_reg[89]  ( .D(addKey_out[89]), .CK(clk), .Q(out[89]) );
  DFF_X1 \out_reg[90]  ( .D(addKey_out[90]), .CK(clk), .Q(out[90]) );
  DFF_X1 \out_reg[91]  ( .D(addKey_out[91]), .CK(clk), .Q(out[91]) );
  DFF_X1 \out_reg[92]  ( .D(addKey_out[92]), .CK(clk), .Q(out[92]) );
  DFF_X1 \out_reg[93]  ( .D(addKey_out[93]), .CK(clk), .Q(out[93]) );
  DFF_X1 \out_reg[94]  ( .D(addKey_out[94]), .CK(clk), .Q(out[94]) );
  DFF_X1 \out_reg[95]  ( .D(addKey_out[95]), .CK(clk), .Q(out[95]) );
  DFF_X1 \out_reg[96]  ( .D(addKey_out[96]), .CK(clk), .Q(out[96]) );
  DFF_X1 \out_reg[97]  ( .D(addKey_out[97]), .CK(clk), .Q(out[97]) );
  DFF_X1 \out_reg[98]  ( .D(addKey_out[98]), .CK(clk), .Q(out[98]) );
  DFF_X1 \out_reg[99]  ( .D(addKey_out[99]), .CK(clk), .Q(out[99]) );
  DFF_X1 \out_reg[100]  ( .D(addKey_out[100]), .CK(clk), .Q(out[100]) );
  DFF_X1 \out_reg[101]  ( .D(addKey_out[101]), .CK(clk), .Q(out[101]) );
  DFF_X1 \out_reg[102]  ( .D(addKey_out[102]), .CK(clk), .Q(out[102]) );
  DFF_X1 \out_reg[103]  ( .D(addKey_out[103]), .CK(clk), .Q(out[103]) );
  DFF_X1 \out_reg[104]  ( .D(addKey_out[104]), .CK(clk), .Q(out[104]) );
  DFF_X1 \out_reg[105]  ( .D(addKey_out[105]), .CK(clk), .Q(out[105]) );
  DFF_X1 \out_reg[106]  ( .D(addKey_out[106]), .CK(clk), .Q(out[106]) );
  DFF_X1 \out_reg[107]  ( .D(addKey_out[107]), .CK(clk), .Q(out[107]) );
  DFF_X1 \out_reg[108]  ( .D(addKey_out[108]), .CK(clk), .Q(out[108]) );
  DFF_X1 \out_reg[109]  ( .D(addKey_out[109]), .CK(clk), .Q(out[109]) );
  DFF_X1 \out_reg[110]  ( .D(addKey_out[110]), .CK(clk), .Q(out[110]) );
  DFF_X1 \out_reg[111]  ( .D(addKey_out[111]), .CK(clk), .Q(out[111]) );
  DFF_X1 \out_reg[112]  ( .D(addKey_out[112]), .CK(clk), .Q(out[112]) );
  DFF_X1 \out_reg[113]  ( .D(addKey_out[113]), .CK(clk), .Q(out[113]) );
  DFF_X1 \out_reg[114]  ( .D(addKey_out[114]), .CK(clk), .Q(out[114]) );
  DFF_X1 \out_reg[115]  ( .D(addKey_out[115]), .CK(clk), .Q(out[115]) );
  DFF_X1 \out_reg[116]  ( .D(addKey_out[116]), .CK(clk), .Q(out[116]) );
  DFF_X1 \out_reg[117]  ( .D(addKey_out[117]), .CK(clk), .Q(out[117]) );
  DFF_X1 \out_reg[118]  ( .D(addKey_out[118]), .CK(clk), .Q(out[118]) );
  DFF_X1 \out_reg[119]  ( .D(addKey_out[119]), .CK(clk), .Q(out[119]) );
  DFF_X1 \out_reg[120]  ( .D(addKey_out[120]), .CK(clk), .Q(out[120]) );
  DFF_X1 \out_reg[121]  ( .D(addKey_out[121]), .CK(clk), .Q(out[121]) );
  DFF_X1 \out_reg[122]  ( .D(addKey_out[122]), .CK(clk), .Q(out[122]) );
  DFF_X1 \out_reg[123]  ( .D(addKey_out[123]), .CK(clk), .Q(out[123]) );
  DFF_X1 \out_reg[124]  ( .D(addKey_out[124]), .CK(clk), .Q(out[124]) );
  DFF_X1 \out_reg[125]  ( .D(addKey_out[125]), .CK(clk), .Q(out[125]) );
  DFF_X1 \out_reg[126]  ( .D(addKey_out[126]), .CK(clk), .Q(out[126]) );
  DFF_X1 \out_reg[127]  ( .D(addKey_out[127]), .CK(clk), .Q(out[127]) );
  INV_X1 U3 ( .A(n453), .ZN(n1) );
  INV_X1 U4 ( .A(data[127]), .ZN(n2) );
  INV_X1 U5 ( .A(n455), .ZN(n3) );
  INV_X1 U6 ( .A(data[126]), .ZN(n4) );
  INV_X1 U7 ( .A(n457), .ZN(n5) );
  INV_X1 U8 ( .A(data[125]), .ZN(n6) );
  INV_X1 U9 ( .A(n459), .ZN(n7) );
  INV_X1 U10 ( .A(data[124]), .ZN(n8) );
  INV_X1 U11 ( .A(n461), .ZN(n9) );
  INV_X1 U12 ( .A(data[123]), .ZN(n10) );
  INV_X1 U13 ( .A(n463), .ZN(n11) );
  INV_X1 U14 ( .A(data[122]), .ZN(n12) );
  INV_X1 U15 ( .A(n465), .ZN(n13) );
  INV_X1 U16 ( .A(data[121]), .ZN(n14) );
  INV_X1 U17 ( .A(n467), .ZN(n15) );
  INV_X1 U18 ( .A(data[120]), .ZN(n16) );
  INV_X1 U19 ( .A(n471), .ZN(n17) );
  INV_X1 U20 ( .A(data[119]), .ZN(n18) );
  INV_X1 U21 ( .A(n473), .ZN(n19) );
  INV_X1 U22 ( .A(data[118]), .ZN(n20) );
  INV_X1 U23 ( .A(n475), .ZN(n21) );
  INV_X1 U24 ( .A(data[117]), .ZN(n22) );
  INV_X1 U25 ( .A(n477), .ZN(n23) );
  INV_X1 U26 ( .A(data[116]), .ZN(n24) );
  INV_X1 U27 ( .A(n479), .ZN(n25) );
  INV_X1 U28 ( .A(data[115]), .ZN(n26) );
  INV_X1 U29 ( .A(n481), .ZN(n27) );
  INV_X1 U30 ( .A(data[114]), .ZN(n28) );
  INV_X1 U31 ( .A(n483), .ZN(n29) );
  INV_X1 U32 ( .A(data[113]), .ZN(n30) );
  INV_X1 U33 ( .A(n485), .ZN(n31) );
  INV_X1 U34 ( .A(data[112]), .ZN(n32) );
  INV_X1 U35 ( .A(n487), .ZN(n33) );
  INV_X1 U36 ( .A(data[111]), .ZN(n34) );
  INV_X1 U37 ( .A(n489), .ZN(n35) );
  INV_X1 U38 ( .A(data[110]), .ZN(n36) );
  INV_X1 U39 ( .A(n493), .ZN(n37) );
  INV_X1 U40 ( .A(data[109]), .ZN(n38) );
  INV_X1 U41 ( .A(n495), .ZN(n39) );
  INV_X1 U42 ( .A(data[108]), .ZN(n40) );
  INV_X1 U43 ( .A(n497), .ZN(n41) );
  INV_X1 U44 ( .A(data[107]), .ZN(n42) );
  INV_X1 U45 ( .A(n499), .ZN(n43) );
  INV_X1 U46 ( .A(data[106]), .ZN(n44) );
  INV_X1 U47 ( .A(n501), .ZN(n45) );
  INV_X1 U48 ( .A(data[105]), .ZN(n46) );
  INV_X1 U49 ( .A(n503), .ZN(n47) );
  INV_X1 U50 ( .A(data[104]), .ZN(n48) );
  INV_X1 U51 ( .A(n505), .ZN(n49) );
  INV_X1 U52 ( .A(data[103]), .ZN(n50) );
  INV_X1 U53 ( .A(n507), .ZN(n51) );
  INV_X1 U54 ( .A(data[102]), .ZN(n52) );
  INV_X1 U55 ( .A(n509), .ZN(n53) );
  INV_X1 U56 ( .A(data[101]), .ZN(n54) );
  INV_X1 U57 ( .A(n511), .ZN(n55) );
  INV_X1 U58 ( .A(data[100]), .ZN(n56) );
  INV_X1 U59 ( .A(n261), .ZN(n57) );
  INV_X1 U60 ( .A(data[99]), .ZN(n58) );
  INV_X1 U61 ( .A(n263), .ZN(n59) );
  INV_X1 U62 ( .A(data[98]), .ZN(n60) );
  INV_X1 U63 ( .A(n265), .ZN(n61) );
  INV_X1 U64 ( .A(data[97]), .ZN(n62) );
  INV_X1 U65 ( .A(n267), .ZN(n63) );
  INV_X1 U66 ( .A(data[96]), .ZN(n64) );
  INV_X1 U67 ( .A(n269), .ZN(n65) );
  INV_X1 U68 ( .A(data[95]), .ZN(n66) );
  INV_X1 U69 ( .A(n271), .ZN(n67) );
  INV_X1 U70 ( .A(data[94]), .ZN(n68) );
  INV_X1 U71 ( .A(n273), .ZN(n69) );
  INV_X1 U72 ( .A(data[93]), .ZN(n70) );
  INV_X1 U73 ( .A(n275), .ZN(n71) );
  INV_X1 U74 ( .A(data[92]), .ZN(n72) );
  INV_X1 U75 ( .A(n277), .ZN(n73) );
  INV_X1 U76 ( .A(data[91]), .ZN(n74) );
  INV_X1 U77 ( .A(n279), .ZN(n75) );
  INV_X1 U78 ( .A(data[90]), .ZN(n76) );
  INV_X1 U79 ( .A(n283), .ZN(n77) );
  INV_X1 U80 ( .A(data[89]), .ZN(n78) );
  INV_X1 U81 ( .A(n285), .ZN(n79) );
  INV_X1 U82 ( .A(data[88]), .ZN(n80) );
  INV_X1 U83 ( .A(n287), .ZN(n81) );
  INV_X1 U84 ( .A(data[87]), .ZN(n82) );
  INV_X1 U85 ( .A(n289), .ZN(n83) );
  INV_X1 U86 ( .A(data[86]), .ZN(n84) );
  INV_X1 U87 ( .A(n291), .ZN(n85) );
  INV_X1 U88 ( .A(data[85]), .ZN(n86) );
  INV_X1 U89 ( .A(n293), .ZN(n87) );
  INV_X1 U90 ( .A(data[84]), .ZN(n88) );
  INV_X1 U91 ( .A(n295), .ZN(n89) );
  INV_X1 U92 ( .A(data[83]), .ZN(n90) );
  INV_X1 U93 ( .A(n297), .ZN(n91) );
  INV_X1 U94 ( .A(data[82]), .ZN(n92) );
  INV_X1 U95 ( .A(n299), .ZN(n93) );
  INV_X1 U96 ( .A(data[81]), .ZN(n94) );
  INV_X1 U97 ( .A(n301), .ZN(n95) );
  INV_X1 U98 ( .A(data[80]), .ZN(n96) );
  INV_X1 U99 ( .A(n305), .ZN(n97) );
  INV_X1 U100 ( .A(data[79]), .ZN(n98) );
  INV_X1 U101 ( .A(n307), .ZN(n99) );
  INV_X1 U102 ( .A(data[78]), .ZN(n100) );
  INV_X1 U103 ( .A(n309), .ZN(n101) );
  INV_X1 U104 ( .A(data[77]), .ZN(n102) );
  INV_X1 U105 ( .A(n311), .ZN(n103) );
  INV_X1 U106 ( .A(data[76]), .ZN(n104) );
  INV_X1 U107 ( .A(n313), .ZN(n105) );
  INV_X1 U108 ( .A(data[75]), .ZN(n106) );
  INV_X1 U109 ( .A(n315), .ZN(n107) );
  INV_X1 U110 ( .A(data[74]), .ZN(n108) );
  INV_X1 U111 ( .A(n317), .ZN(n109) );
  INV_X1 U112 ( .A(data[73]), .ZN(n110) );
  INV_X1 U113 ( .A(n319), .ZN(n111) );
  INV_X1 U114 ( .A(data[72]), .ZN(n112) );
  INV_X1 U115 ( .A(n321), .ZN(n113) );
  INV_X1 U116 ( .A(data[71]), .ZN(n114) );
  INV_X1 U117 ( .A(n323), .ZN(n115) );
  INV_X1 U118 ( .A(data[70]), .ZN(n116) );
  INV_X1 U119 ( .A(n327), .ZN(n117) );
  INV_X1 U120 ( .A(data[69]), .ZN(n118) );
  INV_X1 U121 ( .A(n329), .ZN(n119) );
  INV_X1 U122 ( .A(data[68]), .ZN(n120) );
  INV_X1 U123 ( .A(n331), .ZN(n121) );
  INV_X1 U124 ( .A(data[67]), .ZN(n122) );
  INV_X1 U125 ( .A(n333), .ZN(n123) );
  INV_X1 U126 ( .A(data[66]), .ZN(n124) );
  INV_X1 U127 ( .A(n335), .ZN(n125) );
  INV_X1 U128 ( .A(data[65]), .ZN(n126) );
  INV_X1 U129 ( .A(n337), .ZN(n127) );
  INV_X1 U130 ( .A(data[64]), .ZN(n128) );
  INV_X1 U131 ( .A(n339), .ZN(n129) );
  INV_X1 U132 ( .A(data[63]), .ZN(n130) );
  INV_X1 U133 ( .A(n341), .ZN(n131) );
  INV_X1 U134 ( .A(data[62]), .ZN(n132) );
  INV_X1 U135 ( .A(n343), .ZN(n133) );
  INV_X1 U136 ( .A(data[61]), .ZN(n134) );
  INV_X1 U137 ( .A(n345), .ZN(n135) );
  INV_X1 U138 ( .A(data[60]), .ZN(n136) );
  INV_X1 U139 ( .A(n349), .ZN(n137) );
  INV_X1 U140 ( .A(data[59]), .ZN(n138) );
  INV_X1 U141 ( .A(n351), .ZN(n139) );
  INV_X1 U142 ( .A(data[58]), .ZN(n140) );
  INV_X1 U143 ( .A(n353), .ZN(n141) );
  INV_X1 U144 ( .A(data[57]), .ZN(n142) );
  INV_X1 U145 ( .A(n355), .ZN(n143) );
  INV_X1 U146 ( .A(data[56]), .ZN(n144) );
  INV_X1 U147 ( .A(n357), .ZN(n145) );
  INV_X1 U148 ( .A(data[55]), .ZN(n146) );
  INV_X1 U149 ( .A(n359), .ZN(n147) );
  INV_X1 U150 ( .A(data[54]), .ZN(n148) );
  INV_X1 U151 ( .A(n361), .ZN(n149) );
  INV_X1 U152 ( .A(data[53]), .ZN(n150) );
  INV_X1 U153 ( .A(n363), .ZN(n151) );
  INV_X1 U154 ( .A(data[52]), .ZN(n152) );
  INV_X1 U155 ( .A(n365), .ZN(n153) );
  INV_X1 U156 ( .A(data[51]), .ZN(n154) );
  INV_X1 U157 ( .A(n367), .ZN(n155) );
  INV_X1 U158 ( .A(data[50]), .ZN(n156) );
  INV_X1 U159 ( .A(n371), .ZN(n157) );
  INV_X1 U160 ( .A(data[49]), .ZN(n158) );
  INV_X1 U161 ( .A(n373), .ZN(n159) );
  INV_X1 U162 ( .A(data[48]), .ZN(n160) );
  INV_X1 U163 ( .A(n375), .ZN(n161) );
  INV_X1 U164 ( .A(data[47]), .ZN(n162) );
  INV_X1 U165 ( .A(n377), .ZN(n163) );
  INV_X1 U166 ( .A(data[46]), .ZN(n164) );
  INV_X1 U167 ( .A(n379), .ZN(n165) );
  INV_X1 U168 ( .A(data[45]), .ZN(n166) );
  INV_X1 U169 ( .A(n381), .ZN(n167) );
  INV_X1 U170 ( .A(data[44]), .ZN(n168) );
  INV_X1 U171 ( .A(n383), .ZN(n169) );
  INV_X1 U172 ( .A(data[43]), .ZN(n170) );
  INV_X1 U173 ( .A(n385), .ZN(n171) );
  INV_X1 U174 ( .A(data[42]), .ZN(n172) );
  INV_X1 U175 ( .A(n387), .ZN(n173) );
  INV_X1 U176 ( .A(data[41]), .ZN(n174) );
  INV_X1 U177 ( .A(n389), .ZN(n175) );
  INV_X1 U178 ( .A(data[40]), .ZN(n176) );
  INV_X1 U179 ( .A(n393), .ZN(n177) );
  INV_X1 U180 ( .A(data[39]), .ZN(n178) );
  INV_X1 U181 ( .A(n395), .ZN(n179) );
  INV_X1 U182 ( .A(data[38]), .ZN(n180) );
  INV_X1 U183 ( .A(n397), .ZN(n181) );
  INV_X1 U184 ( .A(data[37]), .ZN(n182) );
  INV_X1 U185 ( .A(n399), .ZN(n183) );
  INV_X1 U186 ( .A(data[36]), .ZN(n184) );
  INV_X1 U187 ( .A(n401), .ZN(n185) );
  INV_X1 U188 ( .A(data[35]), .ZN(n186) );
  INV_X1 U189 ( .A(n403), .ZN(n187) );
  INV_X1 U190 ( .A(data[34]), .ZN(n188) );
  INV_X1 U191 ( .A(n405), .ZN(n189) );
  INV_X1 U192 ( .A(data[33]), .ZN(n190) );
  INV_X1 U193 ( .A(n407), .ZN(n191) );
  INV_X1 U194 ( .A(data[32]), .ZN(n192) );
  INV_X1 U195 ( .A(n409), .ZN(n193) );
  INV_X1 U196 ( .A(data[31]), .ZN(n194) );
  INV_X1 U197 ( .A(n411), .ZN(n195) );
  INV_X1 U198 ( .A(data[30]), .ZN(n196) );
  INV_X1 U199 ( .A(n415), .ZN(n197) );
  INV_X1 U200 ( .A(data[29]), .ZN(n198) );
  INV_X1 U201 ( .A(n417), .ZN(n199) );
  INV_X1 U202 ( .A(data[28]), .ZN(n200) );
  INV_X1 U203 ( .A(n419), .ZN(n201) );
  INV_X1 U204 ( .A(data[27]), .ZN(n202) );
  INV_X1 U205 ( .A(n421), .ZN(n203) );
  INV_X1 U206 ( .A(data[26]), .ZN(n204) );
  INV_X1 U207 ( .A(n423), .ZN(n205) );
  INV_X1 U208 ( .A(data[25]), .ZN(n206) );
  INV_X1 U209 ( .A(n425), .ZN(n207) );
  INV_X1 U210 ( .A(data[24]), .ZN(n208) );
  INV_X1 U211 ( .A(n427), .ZN(n209) );
  INV_X1 U212 ( .A(data[23]), .ZN(n210) );
  INV_X1 U213 ( .A(n429), .ZN(n211) );
  INV_X1 U214 ( .A(data[22]), .ZN(n212) );
  INV_X1 U215 ( .A(n431), .ZN(n213) );
  INV_X1 U216 ( .A(data[21]), .ZN(n214) );
  INV_X1 U217 ( .A(n433), .ZN(n215) );
  INV_X1 U218 ( .A(data[20]), .ZN(n216) );
  INV_X1 U219 ( .A(n437), .ZN(n217) );
  INV_X1 U220 ( .A(data[19]), .ZN(n218) );
  INV_X1 U221 ( .A(n439), .ZN(n219) );
  INV_X1 U222 ( .A(data[18]), .ZN(n220) );
  INV_X1 U223 ( .A(n441), .ZN(n221) );
  INV_X1 U224 ( .A(data[17]), .ZN(n222) );
  INV_X1 U225 ( .A(n443), .ZN(n223) );
  INV_X1 U226 ( .A(data[16]), .ZN(n224) );
  INV_X1 U227 ( .A(n445), .ZN(n225) );
  INV_X1 U228 ( .A(data[15]), .ZN(n226) );
  INV_X1 U229 ( .A(n447), .ZN(n227) );
  INV_X1 U230 ( .A(data[14]), .ZN(n228) );
  INV_X1 U231 ( .A(n449), .ZN(n229) );
  INV_X1 U232 ( .A(data[13]), .ZN(n230) );
  INV_X1 U233 ( .A(n451), .ZN(n231) );
  INV_X1 U234 ( .A(data[12]), .ZN(n232) );
  INV_X1 U235 ( .A(n469), .ZN(n233) );
  INV_X1 U236 ( .A(data[11]), .ZN(n234) );
  INV_X1 U237 ( .A(n491), .ZN(n235) );
  INV_X1 U238 ( .A(data[10]), .ZN(n236) );
  INV_X1 U239 ( .A(n259), .ZN(n237) );
  INV_X1 U240 ( .A(data[9]), .ZN(n238) );
  INV_X1 U241 ( .A(n281), .ZN(n239) );
  INV_X1 U242 ( .A(data[8]), .ZN(n240) );
  INV_X1 U243 ( .A(n303), .ZN(n241) );
  INV_X1 U244 ( .A(data[7]), .ZN(n242) );
  INV_X1 U245 ( .A(n325), .ZN(n243) );
  INV_X1 U246 ( .A(data[6]), .ZN(n244) );
  INV_X1 U247 ( .A(n347), .ZN(n245) );
  INV_X1 U248 ( .A(data[5]), .ZN(n246) );
  INV_X1 U249 ( .A(n369), .ZN(n247) );
  INV_X1 U250 ( .A(data[4]), .ZN(n248) );
  INV_X1 U251 ( .A(n391), .ZN(n249) );
  INV_X1 U252 ( .A(data[3]), .ZN(n250) );
  INV_X1 U253 ( .A(n413), .ZN(n251) );
  INV_X1 U254 ( .A(data[2]), .ZN(n252) );
  INV_X1 U255 ( .A(n435), .ZN(n253) );
  INV_X1 U256 ( .A(data[1]), .ZN(n254) );
  INV_X1 U257 ( .A(n513), .ZN(n255) );
  INV_X1 U258 ( .A(data[0]), .ZN(n256) );
  OR2_X1 U260 ( .A1(n258), .A2(n237), .ZN(state[9]) );
  OR2_X1 U261 ( .A1(n238), .A2(key[9]), .ZN(n259) );
  AND2_X1 U262 ( .A1(key[9]), .A2(n238), .ZN(n258) );
  OR2_X1 U263 ( .A1(n260), .A2(n57), .ZN(state[99]) );
  OR2_X1 U264 ( .A1(n58), .A2(key[99]), .ZN(n261) );
  AND2_X1 U265 ( .A1(key[99]), .A2(n58), .ZN(n260) );
  OR2_X1 U266 ( .A1(n262), .A2(n59), .ZN(state[98]) );
  OR2_X1 U267 ( .A1(n60), .A2(key[98]), .ZN(n263) );
  AND2_X1 U268 ( .A1(key[98]), .A2(n60), .ZN(n262) );
  OR2_X1 U269 ( .A1(n264), .A2(n61), .ZN(state[97]) );
  OR2_X1 U270 ( .A1(n62), .A2(key[97]), .ZN(n265) );
  AND2_X1 U271 ( .A1(key[97]), .A2(n62), .ZN(n264) );
  OR2_X1 U272 ( .A1(n266), .A2(n63), .ZN(state[96]) );
  OR2_X1 U273 ( .A1(n64), .A2(key[96]), .ZN(n267) );
  AND2_X1 U274 ( .A1(key[96]), .A2(n64), .ZN(n266) );
  OR2_X1 U275 ( .A1(n268), .A2(n65), .ZN(state[95]) );
  OR2_X1 U276 ( .A1(n66), .A2(key[95]), .ZN(n269) );
  AND2_X1 U277 ( .A1(key[95]), .A2(n66), .ZN(n268) );
  OR2_X1 U278 ( .A1(n270), .A2(n67), .ZN(state[94]) );
  OR2_X1 U279 ( .A1(n68), .A2(key[94]), .ZN(n271) );
  AND2_X1 U280 ( .A1(key[94]), .A2(n68), .ZN(n270) );
  OR2_X1 U281 ( .A1(n272), .A2(n69), .ZN(state[93]) );
  OR2_X1 U282 ( .A1(n70), .A2(key[93]), .ZN(n273) );
  AND2_X1 U283 ( .A1(key[93]), .A2(n70), .ZN(n272) );
  OR2_X1 U284 ( .A1(n274), .A2(n71), .ZN(state[92]) );
  OR2_X1 U285 ( .A1(n72), .A2(key[92]), .ZN(n275) );
  AND2_X1 U286 ( .A1(key[92]), .A2(n72), .ZN(n274) );
  OR2_X1 U287 ( .A1(n276), .A2(n73), .ZN(state[91]) );
  OR2_X1 U288 ( .A1(n74), .A2(key[91]), .ZN(n277) );
  AND2_X1 U289 ( .A1(key[91]), .A2(n74), .ZN(n276) );
  OR2_X1 U290 ( .A1(n278), .A2(n75), .ZN(state[90]) );
  OR2_X1 U291 ( .A1(n76), .A2(key[90]), .ZN(n279) );
  AND2_X1 U292 ( .A1(key[90]), .A2(n76), .ZN(n278) );
  OR2_X1 U293 ( .A1(n280), .A2(n239), .ZN(state[8]) );
  OR2_X1 U294 ( .A1(n240), .A2(key[8]), .ZN(n281) );
  AND2_X1 U295 ( .A1(key[8]), .A2(n240), .ZN(n280) );
  OR2_X1 U296 ( .A1(n282), .A2(n77), .ZN(state[89]) );
  OR2_X1 U297 ( .A1(n78), .A2(key[89]), .ZN(n283) );
  AND2_X1 U298 ( .A1(key[89]), .A2(n78), .ZN(n282) );
  OR2_X1 U299 ( .A1(n284), .A2(n79), .ZN(state[88]) );
  OR2_X1 U300 ( .A1(n80), .A2(key[88]), .ZN(n285) );
  AND2_X1 U301 ( .A1(key[88]), .A2(n80), .ZN(n284) );
  OR2_X1 U302 ( .A1(n286), .A2(n81), .ZN(state[87]) );
  OR2_X1 U303 ( .A1(n82), .A2(key[87]), .ZN(n287) );
  AND2_X1 U304 ( .A1(key[87]), .A2(n82), .ZN(n286) );
  OR2_X1 U305 ( .A1(n288), .A2(n83), .ZN(state[86]) );
  OR2_X1 U306 ( .A1(n84), .A2(key[86]), .ZN(n289) );
  AND2_X1 U307 ( .A1(key[86]), .A2(n84), .ZN(n288) );
  OR2_X1 U308 ( .A1(n290), .A2(n85), .ZN(state[85]) );
  OR2_X1 U309 ( .A1(n86), .A2(key[85]), .ZN(n291) );
  AND2_X1 U310 ( .A1(key[85]), .A2(n86), .ZN(n290) );
  OR2_X1 U311 ( .A1(n292), .A2(n87), .ZN(state[84]) );
  OR2_X1 U312 ( .A1(n88), .A2(key[84]), .ZN(n293) );
  AND2_X1 U313 ( .A1(key[84]), .A2(n88), .ZN(n292) );
  OR2_X1 U314 ( .A1(n294), .A2(n89), .ZN(state[83]) );
  OR2_X1 U315 ( .A1(n90), .A2(key[83]), .ZN(n295) );
  AND2_X1 U316 ( .A1(key[83]), .A2(n90), .ZN(n294) );
  OR2_X1 U317 ( .A1(n296), .A2(n91), .ZN(state[82]) );
  OR2_X1 U318 ( .A1(n92), .A2(key[82]), .ZN(n297) );
  AND2_X1 U319 ( .A1(key[82]), .A2(n92), .ZN(n296) );
  OR2_X1 U320 ( .A1(n298), .A2(n93), .ZN(state[81]) );
  OR2_X1 U321 ( .A1(n94), .A2(key[81]), .ZN(n299) );
  AND2_X1 U322 ( .A1(key[81]), .A2(n94), .ZN(n298) );
  OR2_X1 U323 ( .A1(n300), .A2(n95), .ZN(state[80]) );
  OR2_X1 U324 ( .A1(n96), .A2(key[80]), .ZN(n301) );
  AND2_X1 U325 ( .A1(key[80]), .A2(n96), .ZN(n300) );
  OR2_X1 U326 ( .A1(n302), .A2(n241), .ZN(state[7]) );
  OR2_X1 U327 ( .A1(n242), .A2(key[7]), .ZN(n303) );
  AND2_X1 U328 ( .A1(key[7]), .A2(n242), .ZN(n302) );
  OR2_X1 U329 ( .A1(n304), .A2(n97), .ZN(state[79]) );
  OR2_X1 U330 ( .A1(n98), .A2(key[79]), .ZN(n305) );
  AND2_X1 U331 ( .A1(key[79]), .A2(n98), .ZN(n304) );
  OR2_X1 U332 ( .A1(n306), .A2(n99), .ZN(state[78]) );
  OR2_X1 U333 ( .A1(n100), .A2(key[78]), .ZN(n307) );
  AND2_X1 U334 ( .A1(key[78]), .A2(n100), .ZN(n306) );
  OR2_X1 U335 ( .A1(n308), .A2(n101), .ZN(state[77]) );
  OR2_X1 U336 ( .A1(n102), .A2(key[77]), .ZN(n309) );
  AND2_X1 U337 ( .A1(key[77]), .A2(n102), .ZN(n308) );
  OR2_X1 U338 ( .A1(n310), .A2(n103), .ZN(state[76]) );
  OR2_X1 U339 ( .A1(n104), .A2(key[76]), .ZN(n311) );
  AND2_X1 U340 ( .A1(key[76]), .A2(n104), .ZN(n310) );
  OR2_X1 U341 ( .A1(n312), .A2(n105), .ZN(state[75]) );
  OR2_X1 U342 ( .A1(n106), .A2(key[75]), .ZN(n313) );
  AND2_X1 U343 ( .A1(key[75]), .A2(n106), .ZN(n312) );
  OR2_X1 U344 ( .A1(n314), .A2(n107), .ZN(state[74]) );
  OR2_X1 U345 ( .A1(n108), .A2(key[74]), .ZN(n315) );
  AND2_X1 U346 ( .A1(key[74]), .A2(n108), .ZN(n314) );
  OR2_X1 U347 ( .A1(n316), .A2(n109), .ZN(state[73]) );
  OR2_X1 U348 ( .A1(n110), .A2(key[73]), .ZN(n317) );
  AND2_X1 U349 ( .A1(key[73]), .A2(n110), .ZN(n316) );
  OR2_X1 U350 ( .A1(n318), .A2(n111), .ZN(state[72]) );
  OR2_X1 U351 ( .A1(n112), .A2(key[72]), .ZN(n319) );
  AND2_X1 U352 ( .A1(key[72]), .A2(n112), .ZN(n318) );
  OR2_X1 U353 ( .A1(n320), .A2(n113), .ZN(state[71]) );
  OR2_X1 U354 ( .A1(n114), .A2(key[71]), .ZN(n321) );
  AND2_X1 U355 ( .A1(key[71]), .A2(n114), .ZN(n320) );
  OR2_X1 U356 ( .A1(n322), .A2(n115), .ZN(state[70]) );
  OR2_X1 U357 ( .A1(n116), .A2(key[70]), .ZN(n323) );
  AND2_X1 U358 ( .A1(key[70]), .A2(n116), .ZN(n322) );
  OR2_X1 U359 ( .A1(n324), .A2(n243), .ZN(state[6]) );
  OR2_X1 U360 ( .A1(n244), .A2(key[6]), .ZN(n325) );
  AND2_X1 U361 ( .A1(key[6]), .A2(n244), .ZN(n324) );
  OR2_X1 U362 ( .A1(n326), .A2(n117), .ZN(state[69]) );
  OR2_X1 U363 ( .A1(n118), .A2(key[69]), .ZN(n327) );
  AND2_X1 U364 ( .A1(key[69]), .A2(n118), .ZN(n326) );
  OR2_X1 U365 ( .A1(n328), .A2(n119), .ZN(state[68]) );
  OR2_X1 U366 ( .A1(n120), .A2(key[68]), .ZN(n329) );
  AND2_X1 U367 ( .A1(key[68]), .A2(n120), .ZN(n328) );
  OR2_X1 U368 ( .A1(n330), .A2(n121), .ZN(state[67]) );
  OR2_X1 U369 ( .A1(n122), .A2(key[67]), .ZN(n331) );
  AND2_X1 U370 ( .A1(key[67]), .A2(n122), .ZN(n330) );
  OR2_X1 U371 ( .A1(n332), .A2(n123), .ZN(state[66]) );
  OR2_X1 U372 ( .A1(n124), .A2(key[66]), .ZN(n333) );
  AND2_X1 U373 ( .A1(key[66]), .A2(n124), .ZN(n332) );
  OR2_X1 U374 ( .A1(n334), .A2(n125), .ZN(state[65]) );
  OR2_X1 U375 ( .A1(n126), .A2(key[65]), .ZN(n335) );
  AND2_X1 U376 ( .A1(key[65]), .A2(n126), .ZN(n334) );
  OR2_X1 U377 ( .A1(n336), .A2(n127), .ZN(state[64]) );
  OR2_X1 U378 ( .A1(n128), .A2(key[64]), .ZN(n337) );
  AND2_X1 U379 ( .A1(key[64]), .A2(n128), .ZN(n336) );
  OR2_X1 U380 ( .A1(n338), .A2(n129), .ZN(state[63]) );
  OR2_X1 U381 ( .A1(n130), .A2(key[63]), .ZN(n339) );
  AND2_X1 U382 ( .A1(key[63]), .A2(n130), .ZN(n338) );
  OR2_X1 U383 ( .A1(n340), .A2(n131), .ZN(state[62]) );
  OR2_X1 U384 ( .A1(n132), .A2(key[62]), .ZN(n341) );
  AND2_X1 U385 ( .A1(key[62]), .A2(n132), .ZN(n340) );
  OR2_X1 U386 ( .A1(n342), .A2(n133), .ZN(state[61]) );
  OR2_X1 U387 ( .A1(n134), .A2(key[61]), .ZN(n343) );
  AND2_X1 U388 ( .A1(key[61]), .A2(n134), .ZN(n342) );
  OR2_X1 U389 ( .A1(n344), .A2(n135), .ZN(state[60]) );
  OR2_X1 U390 ( .A1(n136), .A2(key[60]), .ZN(n345) );
  AND2_X1 U391 ( .A1(key[60]), .A2(n136), .ZN(n344) );
  OR2_X1 U392 ( .A1(n346), .A2(n245), .ZN(state[5]) );
  OR2_X1 U393 ( .A1(n246), .A2(key[5]), .ZN(n347) );
  AND2_X1 U394 ( .A1(key[5]), .A2(n246), .ZN(n346) );
  OR2_X1 U395 ( .A1(n348), .A2(n137), .ZN(state[59]) );
  OR2_X1 U396 ( .A1(n138), .A2(key[59]), .ZN(n349) );
  AND2_X1 U397 ( .A1(key[59]), .A2(n138), .ZN(n348) );
  OR2_X1 U398 ( .A1(n350), .A2(n139), .ZN(state[58]) );
  OR2_X1 U399 ( .A1(n140), .A2(key[58]), .ZN(n351) );
  AND2_X1 U400 ( .A1(key[58]), .A2(n140), .ZN(n350) );
  OR2_X1 U401 ( .A1(n352), .A2(n141), .ZN(state[57]) );
  OR2_X1 U402 ( .A1(n142), .A2(key[57]), .ZN(n353) );
  AND2_X1 U403 ( .A1(key[57]), .A2(n142), .ZN(n352) );
  OR2_X1 U404 ( .A1(n354), .A2(n143), .ZN(state[56]) );
  OR2_X1 U405 ( .A1(n144), .A2(key[56]), .ZN(n355) );
  AND2_X1 U406 ( .A1(key[56]), .A2(n144), .ZN(n354) );
  OR2_X1 U407 ( .A1(n356), .A2(n145), .ZN(state[55]) );
  OR2_X1 U408 ( .A1(n146), .A2(key[55]), .ZN(n357) );
  AND2_X1 U409 ( .A1(key[55]), .A2(n146), .ZN(n356) );
  OR2_X1 U410 ( .A1(n358), .A2(n147), .ZN(state[54]) );
  OR2_X1 U411 ( .A1(n148), .A2(key[54]), .ZN(n359) );
  AND2_X1 U412 ( .A1(key[54]), .A2(n148), .ZN(n358) );
  OR2_X1 U413 ( .A1(n360), .A2(n149), .ZN(state[53]) );
  OR2_X1 U414 ( .A1(n150), .A2(key[53]), .ZN(n361) );
  AND2_X1 U415 ( .A1(key[53]), .A2(n150), .ZN(n360) );
  OR2_X1 U416 ( .A1(n362), .A2(n151), .ZN(state[52]) );
  OR2_X1 U417 ( .A1(n152), .A2(key[52]), .ZN(n363) );
  AND2_X1 U418 ( .A1(key[52]), .A2(n152), .ZN(n362) );
  OR2_X1 U419 ( .A1(n364), .A2(n153), .ZN(state[51]) );
  OR2_X1 U420 ( .A1(n154), .A2(key[51]), .ZN(n365) );
  AND2_X1 U421 ( .A1(key[51]), .A2(n154), .ZN(n364) );
  OR2_X1 U422 ( .A1(n366), .A2(n155), .ZN(state[50]) );
  OR2_X1 U423 ( .A1(n156), .A2(key[50]), .ZN(n367) );
  AND2_X1 U424 ( .A1(key[50]), .A2(n156), .ZN(n366) );
  OR2_X1 U425 ( .A1(n368), .A2(n247), .ZN(state[4]) );
  OR2_X1 U426 ( .A1(n248), .A2(key[4]), .ZN(n369) );
  AND2_X1 U427 ( .A1(key[4]), .A2(n248), .ZN(n368) );
  OR2_X1 U428 ( .A1(n370), .A2(n157), .ZN(state[49]) );
  OR2_X1 U429 ( .A1(n158), .A2(key[49]), .ZN(n371) );
  AND2_X1 U430 ( .A1(key[49]), .A2(n158), .ZN(n370) );
  OR2_X1 U431 ( .A1(n372), .A2(n159), .ZN(state[48]) );
  OR2_X1 U432 ( .A1(n160), .A2(key[48]), .ZN(n373) );
  AND2_X1 U433 ( .A1(key[48]), .A2(n160), .ZN(n372) );
  OR2_X1 U434 ( .A1(n374), .A2(n161), .ZN(state[47]) );
  OR2_X1 U435 ( .A1(n162), .A2(key[47]), .ZN(n375) );
  AND2_X1 U436 ( .A1(key[47]), .A2(n162), .ZN(n374) );
  OR2_X1 U437 ( .A1(n376), .A2(n163), .ZN(state[46]) );
  OR2_X1 U438 ( .A1(n164), .A2(key[46]), .ZN(n377) );
  AND2_X1 U439 ( .A1(key[46]), .A2(n164), .ZN(n376) );
  OR2_X1 U440 ( .A1(n378), .A2(n165), .ZN(state[45]) );
  OR2_X1 U441 ( .A1(n166), .A2(key[45]), .ZN(n379) );
  AND2_X1 U442 ( .A1(key[45]), .A2(n166), .ZN(n378) );
  OR2_X1 U443 ( .A1(n380), .A2(n167), .ZN(state[44]) );
  OR2_X1 U444 ( .A1(n168), .A2(key[44]), .ZN(n381) );
  AND2_X1 U445 ( .A1(key[44]), .A2(n168), .ZN(n380) );
  OR2_X1 U446 ( .A1(n382), .A2(n169), .ZN(state[43]) );
  OR2_X1 U447 ( .A1(n170), .A2(key[43]), .ZN(n383) );
  AND2_X1 U448 ( .A1(key[43]), .A2(n170), .ZN(n382) );
  OR2_X1 U449 ( .A1(n384), .A2(n171), .ZN(state[42]) );
  OR2_X1 U450 ( .A1(n172), .A2(key[42]), .ZN(n385) );
  AND2_X1 U451 ( .A1(key[42]), .A2(n172), .ZN(n384) );
  OR2_X1 U452 ( .A1(n386), .A2(n173), .ZN(state[41]) );
  OR2_X1 U453 ( .A1(n174), .A2(key[41]), .ZN(n387) );
  AND2_X1 U454 ( .A1(key[41]), .A2(n174), .ZN(n386) );
  OR2_X1 U455 ( .A1(n388), .A2(n175), .ZN(state[40]) );
  OR2_X1 U456 ( .A1(n176), .A2(key[40]), .ZN(n389) );
  AND2_X1 U457 ( .A1(key[40]), .A2(n176), .ZN(n388) );
  OR2_X1 U458 ( .A1(n390), .A2(n249), .ZN(state[3]) );
  OR2_X1 U459 ( .A1(n250), .A2(key[3]), .ZN(n391) );
  AND2_X1 U460 ( .A1(key[3]), .A2(n250), .ZN(n390) );
  OR2_X1 U461 ( .A1(n392), .A2(n177), .ZN(state[39]) );
  OR2_X1 U462 ( .A1(n178), .A2(key[39]), .ZN(n393) );
  AND2_X1 U463 ( .A1(key[39]), .A2(n178), .ZN(n392) );
  OR2_X1 U464 ( .A1(n394), .A2(n179), .ZN(state[38]) );
  OR2_X1 U465 ( .A1(n180), .A2(key[38]), .ZN(n395) );
  AND2_X1 U466 ( .A1(key[38]), .A2(n180), .ZN(n394) );
  OR2_X1 U467 ( .A1(n396), .A2(n181), .ZN(state[37]) );
  OR2_X1 U468 ( .A1(n182), .A2(key[37]), .ZN(n397) );
  AND2_X1 U469 ( .A1(key[37]), .A2(n182), .ZN(n396) );
  OR2_X1 U470 ( .A1(n398), .A2(n183), .ZN(state[36]) );
  OR2_X1 U471 ( .A1(n184), .A2(key[36]), .ZN(n399) );
  AND2_X1 U472 ( .A1(key[36]), .A2(n184), .ZN(n398) );
  OR2_X1 U473 ( .A1(n400), .A2(n185), .ZN(state[35]) );
  OR2_X1 U474 ( .A1(n186), .A2(key[35]), .ZN(n401) );
  AND2_X1 U475 ( .A1(key[35]), .A2(n186), .ZN(n400) );
  OR2_X1 U476 ( .A1(n402), .A2(n187), .ZN(state[34]) );
  OR2_X1 U477 ( .A1(n188), .A2(key[34]), .ZN(n403) );
  AND2_X1 U478 ( .A1(key[34]), .A2(n188), .ZN(n402) );
  OR2_X1 U479 ( .A1(n404), .A2(n189), .ZN(state[33]) );
  OR2_X1 U480 ( .A1(n190), .A2(key[33]), .ZN(n405) );
  AND2_X1 U481 ( .A1(key[33]), .A2(n190), .ZN(n404) );
  OR2_X1 U482 ( .A1(n406), .A2(n191), .ZN(state[32]) );
  OR2_X1 U483 ( .A1(n192), .A2(key[32]), .ZN(n407) );
  AND2_X1 U484 ( .A1(key[32]), .A2(n192), .ZN(n406) );
  OR2_X1 U485 ( .A1(n408), .A2(n193), .ZN(state[31]) );
  OR2_X1 U486 ( .A1(n194), .A2(key[31]), .ZN(n409) );
  AND2_X1 U487 ( .A1(key[31]), .A2(n194), .ZN(n408) );
  OR2_X1 U488 ( .A1(n410), .A2(n195), .ZN(state[30]) );
  OR2_X1 U489 ( .A1(n196), .A2(key[30]), .ZN(n411) );
  AND2_X1 U490 ( .A1(key[30]), .A2(n196), .ZN(n410) );
  OR2_X1 U491 ( .A1(n412), .A2(n251), .ZN(state[2]) );
  OR2_X1 U492 ( .A1(n252), .A2(key[2]), .ZN(n413) );
  AND2_X1 U493 ( .A1(key[2]), .A2(n252), .ZN(n412) );
  OR2_X1 U494 ( .A1(n414), .A2(n197), .ZN(state[29]) );
  OR2_X1 U495 ( .A1(n198), .A2(key[29]), .ZN(n415) );
  AND2_X1 U496 ( .A1(key[29]), .A2(n198), .ZN(n414) );
  OR2_X1 U497 ( .A1(n416), .A2(n199), .ZN(state[28]) );
  OR2_X1 U498 ( .A1(n200), .A2(key[28]), .ZN(n417) );
  AND2_X1 U499 ( .A1(key[28]), .A2(n200), .ZN(n416) );
  OR2_X1 U500 ( .A1(n418), .A2(n201), .ZN(state[27]) );
  OR2_X1 U501 ( .A1(n202), .A2(key[27]), .ZN(n419) );
  AND2_X1 U502 ( .A1(key[27]), .A2(n202), .ZN(n418) );
  OR2_X1 U503 ( .A1(n420), .A2(n203), .ZN(state[26]) );
  OR2_X1 U504 ( .A1(n204), .A2(key[26]), .ZN(n421) );
  AND2_X1 U505 ( .A1(key[26]), .A2(n204), .ZN(n420) );
  OR2_X1 U506 ( .A1(n422), .A2(n205), .ZN(state[25]) );
  OR2_X1 U507 ( .A1(n206), .A2(key[25]), .ZN(n423) );
  AND2_X1 U508 ( .A1(key[25]), .A2(n206), .ZN(n422) );
  OR2_X1 U509 ( .A1(n424), .A2(n207), .ZN(state[24]) );
  OR2_X1 U510 ( .A1(n208), .A2(key[24]), .ZN(n425) );
  AND2_X1 U511 ( .A1(key[24]), .A2(n208), .ZN(n424) );
  OR2_X1 U512 ( .A1(n426), .A2(n209), .ZN(state[23]) );
  OR2_X1 U513 ( .A1(n210), .A2(key[23]), .ZN(n427) );
  AND2_X1 U514 ( .A1(key[23]), .A2(n210), .ZN(n426) );
  OR2_X1 U515 ( .A1(n428), .A2(n211), .ZN(state[22]) );
  OR2_X1 U516 ( .A1(n212), .A2(key[22]), .ZN(n429) );
  AND2_X1 U517 ( .A1(key[22]), .A2(n212), .ZN(n428) );
  OR2_X1 U518 ( .A1(n430), .A2(n213), .ZN(state[21]) );
  OR2_X1 U519 ( .A1(n214), .A2(key[21]), .ZN(n431) );
  AND2_X1 U520 ( .A1(key[21]), .A2(n214), .ZN(n430) );
  OR2_X1 U521 ( .A1(n432), .A2(n215), .ZN(state[20]) );
  OR2_X1 U522 ( .A1(n216), .A2(key[20]), .ZN(n433) );
  AND2_X1 U523 ( .A1(key[20]), .A2(n216), .ZN(n432) );
  OR2_X1 U524 ( .A1(n434), .A2(n253), .ZN(state[1]) );
  OR2_X1 U525 ( .A1(n254), .A2(key[1]), .ZN(n435) );
  AND2_X1 U526 ( .A1(key[1]), .A2(n254), .ZN(n434) );
  OR2_X1 U527 ( .A1(n436), .A2(n217), .ZN(state[19]) );
  OR2_X1 U528 ( .A1(n218), .A2(key[19]), .ZN(n437) );
  AND2_X1 U529 ( .A1(key[19]), .A2(n218), .ZN(n436) );
  OR2_X1 U530 ( .A1(n438), .A2(n219), .ZN(state[18]) );
  OR2_X1 U531 ( .A1(n220), .A2(key[18]), .ZN(n439) );
  AND2_X1 U532 ( .A1(key[18]), .A2(n220), .ZN(n438) );
  OR2_X1 U533 ( .A1(n440), .A2(n221), .ZN(state[17]) );
  OR2_X1 U534 ( .A1(n222), .A2(key[17]), .ZN(n441) );
  AND2_X1 U535 ( .A1(key[17]), .A2(n222), .ZN(n440) );
  OR2_X1 U536 ( .A1(n442), .A2(n223), .ZN(state[16]) );
  OR2_X1 U537 ( .A1(n224), .A2(key[16]), .ZN(n443) );
  AND2_X1 U538 ( .A1(key[16]), .A2(n224), .ZN(n442) );
  OR2_X1 U539 ( .A1(n444), .A2(n225), .ZN(state[15]) );
  OR2_X1 U540 ( .A1(n226), .A2(key[15]), .ZN(n445) );
  AND2_X1 U541 ( .A1(key[15]), .A2(n226), .ZN(n444) );
  OR2_X1 U542 ( .A1(n446), .A2(n227), .ZN(state[14]) );
  OR2_X1 U543 ( .A1(n228), .A2(key[14]), .ZN(n447) );
  AND2_X1 U544 ( .A1(key[14]), .A2(n228), .ZN(n446) );
  OR2_X1 U545 ( .A1(n448), .A2(n229), .ZN(state[13]) );
  OR2_X1 U546 ( .A1(n230), .A2(key[13]), .ZN(n449) );
  AND2_X1 U547 ( .A1(key[13]), .A2(n230), .ZN(n448) );
  OR2_X1 U548 ( .A1(n450), .A2(n231), .ZN(state[12]) );
  OR2_X1 U549 ( .A1(n232), .A2(key[12]), .ZN(n451) );
  AND2_X1 U550 ( .A1(key[12]), .A2(n232), .ZN(n450) );
  OR2_X1 U551 ( .A1(n452), .A2(n1), .ZN(state[127]) );
  OR2_X1 U552 ( .A1(n2), .A2(key[127]), .ZN(n453) );
  AND2_X1 U553 ( .A1(key[127]), .A2(n2), .ZN(n452) );
  OR2_X1 U554 ( .A1(n454), .A2(n3), .ZN(state[126]) );
  OR2_X1 U555 ( .A1(n4), .A2(key[126]), .ZN(n455) );
  AND2_X1 U556 ( .A1(key[126]), .A2(n4), .ZN(n454) );
  OR2_X1 U557 ( .A1(n456), .A2(n5), .ZN(state[125]) );
  OR2_X1 U558 ( .A1(n6), .A2(key[125]), .ZN(n457) );
  AND2_X1 U559 ( .A1(key[125]), .A2(n6), .ZN(n456) );
  OR2_X1 U560 ( .A1(n458), .A2(n7), .ZN(state[124]) );
  OR2_X1 U561 ( .A1(n8), .A2(key[124]), .ZN(n459) );
  AND2_X1 U562 ( .A1(key[124]), .A2(n8), .ZN(n458) );
  OR2_X1 U563 ( .A1(n460), .A2(n9), .ZN(state[123]) );
  OR2_X1 U564 ( .A1(n10), .A2(key[123]), .ZN(n461) );
  AND2_X1 U565 ( .A1(key[123]), .A2(n10), .ZN(n460) );
  OR2_X1 U566 ( .A1(n462), .A2(n11), .ZN(state[122]) );
  OR2_X1 U567 ( .A1(n12), .A2(key[122]), .ZN(n463) );
  AND2_X1 U568 ( .A1(key[122]), .A2(n12), .ZN(n462) );
  OR2_X1 U569 ( .A1(n464), .A2(n13), .ZN(state[121]) );
  OR2_X1 U570 ( .A1(n14), .A2(key[121]), .ZN(n465) );
  AND2_X1 U571 ( .A1(key[121]), .A2(n14), .ZN(n464) );
  OR2_X1 U572 ( .A1(n466), .A2(n15), .ZN(state[120]) );
  OR2_X1 U573 ( .A1(n16), .A2(key[120]), .ZN(n467) );
  AND2_X1 U574 ( .A1(key[120]), .A2(n16), .ZN(n466) );
  OR2_X1 U575 ( .A1(n468), .A2(n233), .ZN(state[11]) );
  OR2_X1 U576 ( .A1(n234), .A2(key[11]), .ZN(n469) );
  AND2_X1 U577 ( .A1(key[11]), .A2(n234), .ZN(n468) );
  OR2_X1 U578 ( .A1(n470), .A2(n17), .ZN(state[119]) );
  OR2_X1 U579 ( .A1(n18), .A2(key[119]), .ZN(n471) );
  AND2_X1 U580 ( .A1(key[119]), .A2(n18), .ZN(n470) );
  OR2_X1 U581 ( .A1(n472), .A2(n19), .ZN(state[118]) );
  OR2_X1 U582 ( .A1(n20), .A2(key[118]), .ZN(n473) );
  AND2_X1 U583 ( .A1(key[118]), .A2(n20), .ZN(n472) );
  OR2_X1 U584 ( .A1(n474), .A2(n21), .ZN(state[117]) );
  OR2_X1 U585 ( .A1(n22), .A2(key[117]), .ZN(n475) );
  AND2_X1 U586 ( .A1(key[117]), .A2(n22), .ZN(n474) );
  OR2_X1 U587 ( .A1(n476), .A2(n23), .ZN(state[116]) );
  OR2_X1 U588 ( .A1(n24), .A2(key[116]), .ZN(n477) );
  AND2_X1 U589 ( .A1(key[116]), .A2(n24), .ZN(n476) );
  OR2_X1 U590 ( .A1(n478), .A2(n25), .ZN(state[115]) );
  OR2_X1 U591 ( .A1(n26), .A2(key[115]), .ZN(n479) );
  AND2_X1 U592 ( .A1(key[115]), .A2(n26), .ZN(n478) );
  OR2_X1 U593 ( .A1(n480), .A2(n27), .ZN(state[114]) );
  OR2_X1 U594 ( .A1(n28), .A2(key[114]), .ZN(n481) );
  AND2_X1 U595 ( .A1(key[114]), .A2(n28), .ZN(n480) );
  OR2_X1 U596 ( .A1(n482), .A2(n29), .ZN(state[113]) );
  OR2_X1 U597 ( .A1(n30), .A2(key[113]), .ZN(n483) );
  AND2_X1 U598 ( .A1(key[113]), .A2(n30), .ZN(n482) );
  OR2_X1 U599 ( .A1(n484), .A2(n31), .ZN(state[112]) );
  OR2_X1 U600 ( .A1(n32), .A2(key[112]), .ZN(n485) );
  AND2_X1 U601 ( .A1(key[112]), .A2(n32), .ZN(n484) );
  OR2_X1 U602 ( .A1(n486), .A2(n33), .ZN(state[111]) );
  OR2_X1 U603 ( .A1(n34), .A2(key[111]), .ZN(n487) );
  AND2_X1 U604 ( .A1(key[111]), .A2(n34), .ZN(n486) );
  OR2_X1 U605 ( .A1(n488), .A2(n35), .ZN(state[110]) );
  OR2_X1 U606 ( .A1(n36), .A2(key[110]), .ZN(n489) );
  AND2_X1 U607 ( .A1(key[110]), .A2(n36), .ZN(n488) );
  OR2_X1 U608 ( .A1(n490), .A2(n235), .ZN(state[10]) );
  OR2_X1 U609 ( .A1(n236), .A2(key[10]), .ZN(n491) );
  AND2_X1 U610 ( .A1(key[10]), .A2(n236), .ZN(n490) );
  OR2_X1 U611 ( .A1(n492), .A2(n37), .ZN(state[109]) );
  OR2_X1 U612 ( .A1(n38), .A2(key[109]), .ZN(n493) );
  AND2_X1 U613 ( .A1(key[109]), .A2(n38), .ZN(n492) );
  OR2_X1 U614 ( .A1(n494), .A2(n39), .ZN(state[108]) );
  OR2_X1 U615 ( .A1(n40), .A2(key[108]), .ZN(n495) );
  AND2_X1 U616 ( .A1(key[108]), .A2(n40), .ZN(n494) );
  OR2_X1 U617 ( .A1(n496), .A2(n41), .ZN(state[107]) );
  OR2_X1 U618 ( .A1(n42), .A2(key[107]), .ZN(n497) );
  AND2_X1 U619 ( .A1(key[107]), .A2(n42), .ZN(n496) );
  OR2_X1 U620 ( .A1(n498), .A2(n43), .ZN(state[106]) );
  OR2_X1 U621 ( .A1(n44), .A2(key[106]), .ZN(n499) );
  AND2_X1 U622 ( .A1(key[106]), .A2(n44), .ZN(n498) );
  OR2_X1 U623 ( .A1(n500), .A2(n45), .ZN(state[105]) );
  OR2_X1 U624 ( .A1(n46), .A2(key[105]), .ZN(n501) );
  AND2_X1 U625 ( .A1(key[105]), .A2(n46), .ZN(n500) );
  OR2_X1 U626 ( .A1(n502), .A2(n47), .ZN(state[104]) );
  OR2_X1 U627 ( .A1(n48), .A2(key[104]), .ZN(n503) );
  AND2_X1 U628 ( .A1(key[104]), .A2(n48), .ZN(n502) );
  OR2_X1 U629 ( .A1(n504), .A2(n49), .ZN(state[103]) );
  OR2_X1 U630 ( .A1(n50), .A2(key[103]), .ZN(n505) );
  AND2_X1 U631 ( .A1(key[103]), .A2(n50), .ZN(n504) );
  OR2_X1 U632 ( .A1(n506), .A2(n51), .ZN(state[102]) );
  OR2_X1 U633 ( .A1(n52), .A2(key[102]), .ZN(n507) );
  AND2_X1 U634 ( .A1(key[102]), .A2(n52), .ZN(n506) );
  OR2_X1 U635 ( .A1(n508), .A2(n53), .ZN(state[101]) );
  OR2_X1 U636 ( .A1(n54), .A2(key[101]), .ZN(n509) );
  AND2_X1 U637 ( .A1(key[101]), .A2(n54), .ZN(n508) );
  OR2_X1 U638 ( .A1(n510), .A2(n55), .ZN(state[100]) );
  OR2_X1 U639 ( .A1(n56), .A2(key[100]), .ZN(n511) );
  AND2_X1 U640 ( .A1(key[100]), .A2(n56), .ZN(n510) );
  OR2_X1 U641 ( .A1(n512), .A2(n255), .ZN(state[0]) );
  OR2_X1 U642 ( .A1(n256), .A2(key[0]), .ZN(n513) );
  AND2_X1 U643 ( .A1(key[0]), .A2(n256), .ZN(n512) );
  OR2_X1 U644 ( .A1(n514), .A2(n515), .ZN(mixCol_out[9]) );
  AND2_X1 U645 ( .A1(sBox_out[9]), .A2(final_round), .ZN(n515) );
  AND2_X1 U646 ( .A1(mixCol_out_temp[9]), .A2(n772), .ZN(n514) );
  OR2_X1 U647 ( .A1(n516), .A2(n517), .ZN(mixCol_out[99]) );
  AND2_X1 U648 ( .A1(sBox_out[99]), .A2(final_round), .ZN(n517) );
  AND2_X1 U649 ( .A1(mixCol_out_temp[99]), .A2(n771), .ZN(n516) );
  OR2_X1 U650 ( .A1(n518), .A2(n519), .ZN(mixCol_out[98]) );
  AND2_X1 U651 ( .A1(sBox_out[98]), .A2(final_round), .ZN(n519) );
  AND2_X1 U652 ( .A1(mixCol_out_temp[98]), .A2(n770), .ZN(n518) );
  OR2_X1 U653 ( .A1(n520), .A2(n521), .ZN(mixCol_out[97]) );
  AND2_X1 U654 ( .A1(sBox_out[97]), .A2(final_round), .ZN(n521) );
  AND2_X1 U655 ( .A1(mixCol_out_temp[97]), .A2(n771), .ZN(n520) );
  OR2_X1 U656 ( .A1(n522), .A2(n523), .ZN(mixCol_out[96]) );
  AND2_X1 U657 ( .A1(sBox_out[96]), .A2(final_round), .ZN(n523) );
  AND2_X1 U658 ( .A1(mixCol_out_temp[96]), .A2(n770), .ZN(n522) );
  OR2_X1 U659 ( .A1(n524), .A2(n525), .ZN(mixCol_out[95]) );
  AND2_X1 U660 ( .A1(sBox_out[95]), .A2(final_round), .ZN(n525) );
  AND2_X1 U661 ( .A1(mixCol_out_temp[95]), .A2(n771), .ZN(n524) );
  OR2_X1 U662 ( .A1(n526), .A2(n527), .ZN(mixCol_out[94]) );
  AND2_X1 U663 ( .A1(sBox_out[94]), .A2(final_round), .ZN(n527) );
  AND2_X1 U664 ( .A1(mixCol_out_temp[94]), .A2(n773), .ZN(n526) );
  OR2_X1 U665 ( .A1(n528), .A2(n529), .ZN(mixCol_out[93]) );
  AND2_X1 U666 ( .A1(sBox_out[93]), .A2(final_round), .ZN(n529) );
  AND2_X1 U667 ( .A1(mixCol_out_temp[93]), .A2(n772), .ZN(n528) );
  OR2_X1 U668 ( .A1(n530), .A2(n531), .ZN(mixCol_out[92]) );
  AND2_X1 U669 ( .A1(sBox_out[92]), .A2(final_round), .ZN(n531) );
  AND2_X1 U670 ( .A1(mixCol_out_temp[92]), .A2(n770), .ZN(n530) );
  OR2_X1 U671 ( .A1(n532), .A2(n533), .ZN(mixCol_out[91]) );
  AND2_X1 U672 ( .A1(sBox_out[91]), .A2(final_round), .ZN(n533) );
  AND2_X1 U673 ( .A1(mixCol_out_temp[91]), .A2(n772), .ZN(n532) );
  OR2_X1 U674 ( .A1(n534), .A2(n535), .ZN(mixCol_out[90]) );
  AND2_X1 U675 ( .A1(sBox_out[90]), .A2(final_round), .ZN(n535) );
  AND2_X1 U676 ( .A1(mixCol_out_temp[90]), .A2(n770), .ZN(n534) );
  OR2_X1 U677 ( .A1(n536), .A2(n537), .ZN(mixCol_out[8]) );
  AND2_X1 U678 ( .A1(sBox_out[8]), .A2(final_round), .ZN(n537) );
  AND2_X1 U679 ( .A1(mixCol_out_temp[8]), .A2(n771), .ZN(n536) );
  OR2_X1 U680 ( .A1(n538), .A2(n539), .ZN(mixCol_out[89]) );
  AND2_X1 U681 ( .A1(sBox_out[89]), .A2(final_round), .ZN(n539) );
  AND2_X1 U682 ( .A1(mixCol_out_temp[89]), .A2(n771), .ZN(n538) );
  OR2_X1 U683 ( .A1(n540), .A2(n541), .ZN(mixCol_out[88]) );
  AND2_X1 U684 ( .A1(sBox_out[88]), .A2(final_round), .ZN(n541) );
  AND2_X1 U685 ( .A1(mixCol_out_temp[88]), .A2(n771), .ZN(n540) );
  OR2_X1 U686 ( .A1(n542), .A2(n543), .ZN(mixCol_out[87]) );
  AND2_X1 U687 ( .A1(sBox_out[87]), .A2(final_round), .ZN(n543) );
  AND2_X1 U688 ( .A1(mixCol_out_temp[87]), .A2(n770), .ZN(n542) );
  OR2_X1 U689 ( .A1(n544), .A2(n545), .ZN(mixCol_out[86]) );
  AND2_X1 U690 ( .A1(sBox_out[86]), .A2(final_round), .ZN(n545) );
  AND2_X1 U691 ( .A1(mixCol_out_temp[86]), .A2(n773), .ZN(n544) );
  OR2_X1 U692 ( .A1(n546), .A2(n547), .ZN(mixCol_out[85]) );
  AND2_X1 U693 ( .A1(sBox_out[85]), .A2(final_round), .ZN(n547) );
  AND2_X1 U694 ( .A1(mixCol_out_temp[85]), .A2(n772), .ZN(n546) );
  OR2_X1 U695 ( .A1(n548), .A2(n549), .ZN(mixCol_out[84]) );
  AND2_X1 U696 ( .A1(sBox_out[84]), .A2(final_round), .ZN(n549) );
  AND2_X1 U697 ( .A1(mixCol_out_temp[84]), .A2(n772), .ZN(n548) );
  OR2_X1 U698 ( .A1(n550), .A2(n551), .ZN(mixCol_out[83]) );
  AND2_X1 U699 ( .A1(sBox_out[83]), .A2(final_round), .ZN(n551) );
  AND2_X1 U700 ( .A1(mixCol_out_temp[83]), .A2(n773), .ZN(n550) );
  OR2_X1 U701 ( .A1(n552), .A2(n553), .ZN(mixCol_out[82]) );
  AND2_X1 U702 ( .A1(sBox_out[82]), .A2(final_round), .ZN(n553) );
  AND2_X1 U703 ( .A1(mixCol_out_temp[82]), .A2(n773), .ZN(n552) );
  OR2_X1 U704 ( .A1(n554), .A2(n555), .ZN(mixCol_out[81]) );
  AND2_X1 U705 ( .A1(sBox_out[81]), .A2(final_round), .ZN(n555) );
  AND2_X1 U706 ( .A1(mixCol_out_temp[81]), .A2(n771), .ZN(n554) );
  OR2_X1 U707 ( .A1(n556), .A2(n557), .ZN(mixCol_out[80]) );
  AND2_X1 U708 ( .A1(sBox_out[80]), .A2(final_round), .ZN(n557) );
  AND2_X1 U709 ( .A1(mixCol_out_temp[80]), .A2(n772), .ZN(n556) );
  OR2_X1 U710 ( .A1(n558), .A2(n559), .ZN(mixCol_out[7]) );
  AND2_X1 U711 ( .A1(sBox_out[7]), .A2(final_round), .ZN(n559) );
  AND2_X1 U712 ( .A1(mixCol_out_temp[7]), .A2(n772), .ZN(n558) );
  OR2_X1 U713 ( .A1(n560), .A2(n561), .ZN(mixCol_out[79]) );
  AND2_X1 U714 ( .A1(sBox_out[79]), .A2(final_round), .ZN(n561) );
  AND2_X1 U715 ( .A1(mixCol_out_temp[79]), .A2(n771), .ZN(n560) );
  OR2_X1 U716 ( .A1(n562), .A2(n563), .ZN(mixCol_out[78]) );
  AND2_X1 U717 ( .A1(sBox_out[78]), .A2(final_round), .ZN(n563) );
  AND2_X1 U718 ( .A1(mixCol_out_temp[78]), .A2(n773), .ZN(n562) );
  OR2_X1 U719 ( .A1(n564), .A2(n565), .ZN(mixCol_out[77]) );
  AND2_X1 U720 ( .A1(sBox_out[77]), .A2(final_round), .ZN(n565) );
  AND2_X1 U721 ( .A1(mixCol_out_temp[77]), .A2(n772), .ZN(n564) );
  OR2_X1 U722 ( .A1(n566), .A2(n567), .ZN(mixCol_out[76]) );
  AND2_X1 U723 ( .A1(sBox_out[76]), .A2(final_round), .ZN(n567) );
  AND2_X1 U724 ( .A1(mixCol_out_temp[76]), .A2(n773), .ZN(n566) );
  OR2_X1 U725 ( .A1(n568), .A2(n569), .ZN(mixCol_out[75]) );
  AND2_X1 U726 ( .A1(sBox_out[75]), .A2(final_round), .ZN(n569) );
  AND2_X1 U727 ( .A1(mixCol_out_temp[75]), .A2(n772), .ZN(n568) );
  OR2_X1 U728 ( .A1(n570), .A2(n571), .ZN(mixCol_out[74]) );
  AND2_X1 U729 ( .A1(sBox_out[74]), .A2(final_round), .ZN(n571) );
  AND2_X1 U730 ( .A1(mixCol_out_temp[74]), .A2(n771), .ZN(n570) );
  OR2_X1 U731 ( .A1(n572), .A2(n573), .ZN(mixCol_out[73]) );
  AND2_X1 U732 ( .A1(sBox_out[73]), .A2(final_round), .ZN(n573) );
  AND2_X1 U733 ( .A1(mixCol_out_temp[73]), .A2(n771), .ZN(n572) );
  OR2_X1 U734 ( .A1(n574), .A2(n575), .ZN(mixCol_out[72]) );
  AND2_X1 U735 ( .A1(sBox_out[72]), .A2(final_round), .ZN(n575) );
  AND2_X1 U736 ( .A1(mixCol_out_temp[72]), .A2(n771), .ZN(n574) );
  OR2_X1 U737 ( .A1(n576), .A2(n577), .ZN(mixCol_out[71]) );
  AND2_X1 U738 ( .A1(sBox_out[71]), .A2(final_round), .ZN(n577) );
  AND2_X1 U739 ( .A1(mixCol_out_temp[71]), .A2(n771), .ZN(n576) );
  OR2_X1 U740 ( .A1(n578), .A2(n579), .ZN(mixCol_out[70]) );
  AND2_X1 U741 ( .A1(sBox_out[70]), .A2(final_round), .ZN(n579) );
  AND2_X1 U742 ( .A1(mixCol_out_temp[70]), .A2(n771), .ZN(n578) );
  OR2_X1 U743 ( .A1(n580), .A2(n581), .ZN(mixCol_out[6]) );
  AND2_X1 U744 ( .A1(sBox_out[6]), .A2(final_round), .ZN(n581) );
  AND2_X1 U745 ( .A1(mixCol_out_temp[6]), .A2(n770), .ZN(n580) );
  OR2_X1 U746 ( .A1(n582), .A2(n583), .ZN(mixCol_out[69]) );
  AND2_X1 U747 ( .A1(sBox_out[69]), .A2(final_round), .ZN(n583) );
  AND2_X1 U748 ( .A1(mixCol_out_temp[69]), .A2(n770), .ZN(n582) );
  OR2_X1 U749 ( .A1(n584), .A2(n585), .ZN(mixCol_out[68]) );
  AND2_X1 U750 ( .A1(sBox_out[68]), .A2(final_round), .ZN(n585) );
  AND2_X1 U751 ( .A1(mixCol_out_temp[68]), .A2(n771), .ZN(n584) );
  OR2_X1 U752 ( .A1(n586), .A2(n587), .ZN(mixCol_out[67]) );
  AND2_X1 U753 ( .A1(sBox_out[67]), .A2(final_round), .ZN(n587) );
  AND2_X1 U754 ( .A1(mixCol_out_temp[67]), .A2(n771), .ZN(n586) );
  OR2_X1 U755 ( .A1(n588), .A2(n589), .ZN(mixCol_out[66]) );
  AND2_X1 U756 ( .A1(sBox_out[66]), .A2(final_round), .ZN(n589) );
  AND2_X1 U757 ( .A1(mixCol_out_temp[66]), .A2(n773), .ZN(n588) );
  OR2_X1 U758 ( .A1(n590), .A2(n591), .ZN(mixCol_out[65]) );
  AND2_X1 U759 ( .A1(sBox_out[65]), .A2(final_round), .ZN(n591) );
  AND2_X1 U760 ( .A1(mixCol_out_temp[65]), .A2(n771), .ZN(n590) );
  OR2_X1 U761 ( .A1(n592), .A2(n593), .ZN(mixCol_out[64]) );
  AND2_X1 U762 ( .A1(sBox_out[64]), .A2(final_round), .ZN(n593) );
  AND2_X1 U763 ( .A1(mixCol_out_temp[64]), .A2(n772), .ZN(n592) );
  OR2_X1 U764 ( .A1(n594), .A2(n595), .ZN(mixCol_out[63]) );
  AND2_X1 U765 ( .A1(sBox_out[63]), .A2(final_round), .ZN(n595) );
  AND2_X1 U766 ( .A1(mixCol_out_temp[63]), .A2(n771), .ZN(n594) );
  OR2_X1 U767 ( .A1(n596), .A2(n597), .ZN(mixCol_out[62]) );
  AND2_X1 U768 ( .A1(sBox_out[62]), .A2(final_round), .ZN(n597) );
  AND2_X1 U769 ( .A1(mixCol_out_temp[62]), .A2(n770), .ZN(n596) );
  OR2_X1 U770 ( .A1(n598), .A2(n599), .ZN(mixCol_out[61]) );
  AND2_X1 U771 ( .A1(sBox_out[61]), .A2(final_round), .ZN(n599) );
  AND2_X1 U772 ( .A1(mixCol_out_temp[61]), .A2(n770), .ZN(n598) );
  OR2_X1 U773 ( .A1(n600), .A2(n601), .ZN(mixCol_out[60]) );
  AND2_X1 U774 ( .A1(sBox_out[60]), .A2(final_round), .ZN(n601) );
  AND2_X1 U775 ( .A1(mixCol_out_temp[60]), .A2(n771), .ZN(n600) );
  OR2_X1 U776 ( .A1(n602), .A2(n603), .ZN(mixCol_out[5]) );
  AND2_X1 U777 ( .A1(sBox_out[5]), .A2(final_round), .ZN(n603) );
  AND2_X1 U778 ( .A1(mixCol_out_temp[5]), .A2(n770), .ZN(n602) );
  OR2_X1 U779 ( .A1(n604), .A2(n605), .ZN(mixCol_out[59]) );
  AND2_X1 U780 ( .A1(sBox_out[59]), .A2(final_round), .ZN(n605) );
  AND2_X1 U781 ( .A1(mixCol_out_temp[59]), .A2(n770), .ZN(n604) );
  OR2_X1 U782 ( .A1(n606), .A2(n607), .ZN(mixCol_out[58]) );
  AND2_X1 U783 ( .A1(sBox_out[58]), .A2(final_round), .ZN(n607) );
  AND2_X1 U784 ( .A1(mixCol_out_temp[58]), .A2(n771), .ZN(n606) );
  OR2_X1 U785 ( .A1(n608), .A2(n609), .ZN(mixCol_out[57]) );
  AND2_X1 U786 ( .A1(sBox_out[57]), .A2(final_round), .ZN(n609) );
  AND2_X1 U787 ( .A1(mixCol_out_temp[57]), .A2(n773), .ZN(n608) );
  OR2_X1 U788 ( .A1(n610), .A2(n611), .ZN(mixCol_out[56]) );
  AND2_X1 U789 ( .A1(sBox_out[56]), .A2(final_round), .ZN(n611) );
  AND2_X1 U790 ( .A1(mixCol_out_temp[56]), .A2(n771), .ZN(n610) );
  OR2_X1 U791 ( .A1(n612), .A2(n613), .ZN(mixCol_out[55]) );
  AND2_X1 U792 ( .A1(sBox_out[55]), .A2(final_round), .ZN(n613) );
  AND2_X1 U793 ( .A1(mixCol_out_temp[55]), .A2(n770), .ZN(n612) );
  OR2_X1 U794 ( .A1(n614), .A2(n615), .ZN(mixCol_out[54]) );
  AND2_X1 U795 ( .A1(sBox_out[54]), .A2(final_round), .ZN(n615) );
  AND2_X1 U796 ( .A1(mixCol_out_temp[54]), .A2(n770), .ZN(n614) );
  OR2_X1 U797 ( .A1(n616), .A2(n617), .ZN(mixCol_out[53]) );
  AND2_X1 U798 ( .A1(sBox_out[53]), .A2(final_round), .ZN(n617) );
  AND2_X1 U799 ( .A1(mixCol_out_temp[53]), .A2(n771), .ZN(n616) );
  OR2_X1 U800 ( .A1(n618), .A2(n619), .ZN(mixCol_out[52]) );
  AND2_X1 U801 ( .A1(sBox_out[52]), .A2(final_round), .ZN(n619) );
  AND2_X1 U802 ( .A1(mixCol_out_temp[52]), .A2(n770), .ZN(n618) );
  OR2_X1 U803 ( .A1(n620), .A2(n621), .ZN(mixCol_out[51]) );
  AND2_X1 U804 ( .A1(sBox_out[51]), .A2(final_round), .ZN(n621) );
  AND2_X1 U805 ( .A1(mixCol_out_temp[51]), .A2(n772), .ZN(n620) );
  OR2_X1 U806 ( .A1(n622), .A2(n623), .ZN(mixCol_out[50]) );
  AND2_X1 U807 ( .A1(sBox_out[50]), .A2(final_round), .ZN(n623) );
  AND2_X1 U808 ( .A1(mixCol_out_temp[50]), .A2(n771), .ZN(n622) );
  OR2_X1 U809 ( .A1(n624), .A2(n625), .ZN(mixCol_out[4]) );
  AND2_X1 U810 ( .A1(sBox_out[4]), .A2(final_round), .ZN(n625) );
  AND2_X1 U811 ( .A1(mixCol_out_temp[4]), .A2(n772), .ZN(n624) );
  OR2_X1 U812 ( .A1(n626), .A2(n627), .ZN(mixCol_out[49]) );
  AND2_X1 U813 ( .A1(sBox_out[49]), .A2(final_round), .ZN(n627) );
  AND2_X1 U814 ( .A1(mixCol_out_temp[49]), .A2(n770), .ZN(n626) );
  OR2_X1 U815 ( .A1(n628), .A2(n629), .ZN(mixCol_out[48]) );
  AND2_X1 U816 ( .A1(sBox_out[48]), .A2(final_round), .ZN(n629) );
  AND2_X1 U817 ( .A1(mixCol_out_temp[48]), .A2(n770), .ZN(n628) );
  OR2_X1 U818 ( .A1(n630), .A2(n631), .ZN(mixCol_out[47]) );
  AND2_X1 U819 ( .A1(sBox_out[47]), .A2(final_round), .ZN(n631) );
  AND2_X1 U820 ( .A1(mixCol_out_temp[47]), .A2(n771), .ZN(n630) );
  OR2_X1 U821 ( .A1(n632), .A2(n633), .ZN(mixCol_out[46]) );
  AND2_X1 U822 ( .A1(sBox_out[46]), .A2(final_round), .ZN(n633) );
  AND2_X1 U823 ( .A1(mixCol_out_temp[46]), .A2(n771), .ZN(n632) );
  OR2_X1 U824 ( .A1(n634), .A2(n635), .ZN(mixCol_out[45]) );
  AND2_X1 U825 ( .A1(sBox_out[45]), .A2(final_round), .ZN(n635) );
  AND2_X1 U826 ( .A1(mixCol_out_temp[45]), .A2(n770), .ZN(n634) );
  OR2_X1 U827 ( .A1(n636), .A2(n637), .ZN(mixCol_out[44]) );
  AND2_X1 U828 ( .A1(sBox_out[44]), .A2(final_round), .ZN(n637) );
  AND2_X1 U829 ( .A1(mixCol_out_temp[44]), .A2(n770), .ZN(n636) );
  OR2_X1 U830 ( .A1(n638), .A2(n639), .ZN(mixCol_out[43]) );
  AND2_X1 U831 ( .A1(sBox_out[43]), .A2(final_round), .ZN(n639) );
  AND2_X1 U832 ( .A1(mixCol_out_temp[43]), .A2(n773), .ZN(n638) );
  OR2_X1 U833 ( .A1(n640), .A2(n641), .ZN(mixCol_out[42]) );
  AND2_X1 U834 ( .A1(sBox_out[42]), .A2(final_round), .ZN(n641) );
  AND2_X1 U835 ( .A1(mixCol_out_temp[42]), .A2(n771), .ZN(n640) );
  OR2_X1 U836 ( .A1(n642), .A2(n643), .ZN(mixCol_out[41]) );
  AND2_X1 U837 ( .A1(sBox_out[41]), .A2(final_round), .ZN(n643) );
  AND2_X1 U838 ( .A1(mixCol_out_temp[41]), .A2(n771), .ZN(n642) );
  OR2_X1 U839 ( .A1(n644), .A2(n645), .ZN(mixCol_out[40]) );
  AND2_X1 U840 ( .A1(sBox_out[40]), .A2(final_round), .ZN(n645) );
  AND2_X1 U841 ( .A1(mixCol_out_temp[40]), .A2(n773), .ZN(n644) );
  OR2_X1 U842 ( .A1(n646), .A2(n647), .ZN(mixCol_out[3]) );
  AND2_X1 U843 ( .A1(sBox_out[3]), .A2(final_round), .ZN(n647) );
  AND2_X1 U844 ( .A1(mixCol_out_temp[3]), .A2(n770), .ZN(n646) );
  OR2_X1 U845 ( .A1(n648), .A2(n649), .ZN(mixCol_out[39]) );
  AND2_X1 U846 ( .A1(sBox_out[39]), .A2(final_round), .ZN(n649) );
  AND2_X1 U847 ( .A1(mixCol_out_temp[39]), .A2(n771), .ZN(n648) );
  OR2_X1 U848 ( .A1(n650), .A2(n651), .ZN(mixCol_out[38]) );
  AND2_X1 U849 ( .A1(sBox_out[38]), .A2(final_round), .ZN(n651) );
  AND2_X1 U850 ( .A1(mixCol_out_temp[38]), .A2(n770), .ZN(n650) );
  OR2_X1 U851 ( .A1(n652), .A2(n653), .ZN(mixCol_out[37]) );
  AND2_X1 U852 ( .A1(sBox_out[37]), .A2(final_round), .ZN(n653) );
  AND2_X1 U853 ( .A1(mixCol_out_temp[37]), .A2(n773), .ZN(n652) );
  OR2_X1 U854 ( .A1(n654), .A2(n655), .ZN(mixCol_out[36]) );
  AND2_X1 U855 ( .A1(sBox_out[36]), .A2(final_round), .ZN(n655) );
  AND2_X1 U856 ( .A1(mixCol_out_temp[36]), .A2(n772), .ZN(n654) );
  OR2_X1 U857 ( .A1(n656), .A2(n657), .ZN(mixCol_out[35]) );
  AND2_X1 U858 ( .A1(sBox_out[35]), .A2(final_round), .ZN(n657) );
  AND2_X1 U859 ( .A1(mixCol_out_temp[35]), .A2(n770), .ZN(n656) );
  OR2_X1 U860 ( .A1(n658), .A2(n659), .ZN(mixCol_out[34]) );
  AND2_X1 U861 ( .A1(sBox_out[34]), .A2(final_round), .ZN(n659) );
  AND2_X1 U862 ( .A1(mixCol_out_temp[34]), .A2(n771), .ZN(n658) );
  OR2_X1 U863 ( .A1(n660), .A2(n661), .ZN(mixCol_out[33]) );
  AND2_X1 U864 ( .A1(sBox_out[33]), .A2(final_round), .ZN(n661) );
  AND2_X1 U865 ( .A1(mixCol_out_temp[33]), .A2(n773), .ZN(n660) );
  OR2_X1 U866 ( .A1(n662), .A2(n663), .ZN(mixCol_out[32]) );
  AND2_X1 U867 ( .A1(sBox_out[32]), .A2(final_round), .ZN(n663) );
  AND2_X1 U868 ( .A1(mixCol_out_temp[32]), .A2(n772), .ZN(n662) );
  OR2_X1 U869 ( .A1(n664), .A2(n665), .ZN(mixCol_out[31]) );
  AND2_X1 U870 ( .A1(sBox_out[31]), .A2(final_round), .ZN(n665) );
  AND2_X1 U871 ( .A1(mixCol_out_temp[31]), .A2(n771), .ZN(n664) );
  OR2_X1 U872 ( .A1(n666), .A2(n667), .ZN(mixCol_out[30]) );
  AND2_X1 U873 ( .A1(sBox_out[30]), .A2(final_round), .ZN(n667) );
  AND2_X1 U874 ( .A1(mixCol_out_temp[30]), .A2(n770), .ZN(n666) );
  OR2_X1 U875 ( .A1(n668), .A2(n669), .ZN(mixCol_out[2]) );
  AND2_X1 U876 ( .A1(sBox_out[2]), .A2(final_round), .ZN(n669) );
  AND2_X1 U877 ( .A1(mixCol_out_temp[2]), .A2(n770), .ZN(n668) );
  OR2_X1 U878 ( .A1(n670), .A2(n671), .ZN(mixCol_out[29]) );
  AND2_X1 U879 ( .A1(sBox_out[29]), .A2(final_round), .ZN(n671) );
  AND2_X1 U880 ( .A1(mixCol_out_temp[29]), .A2(n770), .ZN(n670) );
  OR2_X1 U881 ( .A1(n672), .A2(n673), .ZN(mixCol_out[28]) );
  AND2_X1 U882 ( .A1(sBox_out[28]), .A2(final_round), .ZN(n673) );
  AND2_X1 U883 ( .A1(mixCol_out_temp[28]), .A2(n773), .ZN(n672) );
  OR2_X1 U884 ( .A1(n674), .A2(n675), .ZN(mixCol_out[27]) );
  AND2_X1 U885 ( .A1(sBox_out[27]), .A2(final_round), .ZN(n675) );
  AND2_X1 U886 ( .A1(mixCol_out_temp[27]), .A2(n773), .ZN(n674) );
  OR2_X1 U887 ( .A1(n676), .A2(n677), .ZN(mixCol_out[26]) );
  AND2_X1 U888 ( .A1(sBox_out[26]), .A2(final_round), .ZN(n677) );
  AND2_X1 U889 ( .A1(mixCol_out_temp[26]), .A2(n772), .ZN(n676) );
  OR2_X1 U890 ( .A1(n678), .A2(n679), .ZN(mixCol_out[25]) );
  AND2_X1 U891 ( .A1(sBox_out[25]), .A2(final_round), .ZN(n679) );
  AND2_X1 U892 ( .A1(mixCol_out_temp[25]), .A2(n770), .ZN(n678) );
  OR2_X1 U893 ( .A1(n680), .A2(n681), .ZN(mixCol_out[24]) );
  AND2_X1 U894 ( .A1(sBox_out[24]), .A2(final_round), .ZN(n681) );
  AND2_X1 U895 ( .A1(mixCol_out_temp[24]), .A2(n773), .ZN(n680) );
  OR2_X1 U896 ( .A1(n682), .A2(n683), .ZN(mixCol_out[23]) );
  AND2_X1 U897 ( .A1(sBox_out[23]), .A2(final_round), .ZN(n683) );
  AND2_X1 U898 ( .A1(mixCol_out_temp[23]), .A2(n772), .ZN(n682) );
  OR2_X1 U899 ( .A1(n684), .A2(n685), .ZN(mixCol_out[22]) );
  AND2_X1 U900 ( .A1(sBox_out[22]), .A2(final_round), .ZN(n685) );
  AND2_X1 U901 ( .A1(mixCol_out_temp[22]), .A2(n773), .ZN(n684) );
  OR2_X1 U902 ( .A1(n686), .A2(n687), .ZN(mixCol_out[21]) );
  AND2_X1 U903 ( .A1(sBox_out[21]), .A2(final_round), .ZN(n687) );
  AND2_X1 U904 ( .A1(mixCol_out_temp[21]), .A2(n772), .ZN(n686) );
  OR2_X1 U905 ( .A1(n688), .A2(n689), .ZN(mixCol_out[20]) );
  AND2_X1 U906 ( .A1(sBox_out[20]), .A2(final_round), .ZN(n689) );
  AND2_X1 U907 ( .A1(mixCol_out_temp[20]), .A2(n770), .ZN(n688) );
  OR2_X1 U908 ( .A1(n690), .A2(n691), .ZN(mixCol_out[1]) );
  AND2_X1 U909 ( .A1(sBox_out[1]), .A2(final_round), .ZN(n691) );
  AND2_X1 U910 ( .A1(mixCol_out_temp[1]), .A2(n773), .ZN(n690) );
  OR2_X1 U911 ( .A1(n692), .A2(n693), .ZN(mixCol_out[19]) );
  AND2_X1 U912 ( .A1(sBox_out[19]), .A2(final_round), .ZN(n693) );
  AND2_X1 U913 ( .A1(mixCol_out_temp[19]), .A2(n770), .ZN(n692) );
  OR2_X1 U914 ( .A1(n694), .A2(n695), .ZN(mixCol_out[18]) );
  AND2_X1 U915 ( .A1(sBox_out[18]), .A2(final_round), .ZN(n695) );
  AND2_X1 U916 ( .A1(mixCol_out_temp[18]), .A2(n773), .ZN(n694) );
  OR2_X1 U917 ( .A1(n696), .A2(n697), .ZN(mixCol_out[17]) );
  AND2_X1 U918 ( .A1(sBox_out[17]), .A2(final_round), .ZN(n697) );
  AND2_X1 U919 ( .A1(mixCol_out_temp[17]), .A2(n773), .ZN(n696) );
  OR2_X1 U920 ( .A1(n698), .A2(n699), .ZN(mixCol_out[16]) );
  AND2_X1 U921 ( .A1(sBox_out[16]), .A2(final_round), .ZN(n699) );
  AND2_X1 U922 ( .A1(mixCol_out_temp[16]), .A2(n772), .ZN(n698) );
  OR2_X1 U923 ( .A1(n700), .A2(n701), .ZN(mixCol_out[15]) );
  AND2_X1 U924 ( .A1(sBox_out[15]), .A2(final_round), .ZN(n701) );
  AND2_X1 U925 ( .A1(mixCol_out_temp[15]), .A2(n770), .ZN(n700) );
  OR2_X1 U926 ( .A1(n702), .A2(n703), .ZN(mixCol_out[14]) );
  AND2_X1 U927 ( .A1(sBox_out[14]), .A2(final_round), .ZN(n703) );
  AND2_X1 U928 ( .A1(mixCol_out_temp[14]), .A2(n772), .ZN(n702) );
  OR2_X1 U929 ( .A1(n704), .A2(n705), .ZN(mixCol_out[13]) );
  AND2_X1 U930 ( .A1(sBox_out[13]), .A2(final_round), .ZN(n705) );
  AND2_X1 U931 ( .A1(mixCol_out_temp[13]), .A2(n771), .ZN(n704) );
  OR2_X1 U932 ( .A1(n706), .A2(n707), .ZN(mixCol_out[12]) );
  AND2_X1 U933 ( .A1(sBox_out[12]), .A2(final_round), .ZN(n707) );
  AND2_X1 U934 ( .A1(mixCol_out_temp[12]), .A2(n772), .ZN(n706) );
  OR2_X1 U935 ( .A1(n708), .A2(n709), .ZN(mixCol_out[127]) );
  AND2_X1 U936 ( .A1(sBox_out[127]), .A2(final_round), .ZN(n709) );
  AND2_X1 U937 ( .A1(mixCol_out_temp[127]), .A2(n773), .ZN(n708) );
  OR2_X1 U938 ( .A1(n710), .A2(n711), .ZN(mixCol_out[126]) );
  AND2_X1 U939 ( .A1(sBox_out[126]), .A2(final_round), .ZN(n711) );
  AND2_X1 U940 ( .A1(mixCol_out_temp[126]), .A2(n772), .ZN(n710) );
  OR2_X1 U941 ( .A1(n712), .A2(n713), .ZN(mixCol_out[125]) );
  AND2_X1 U942 ( .A1(sBox_out[125]), .A2(final_round), .ZN(n713) );
  AND2_X1 U943 ( .A1(mixCol_out_temp[125]), .A2(n772), .ZN(n712) );
  OR2_X1 U944 ( .A1(n714), .A2(n715), .ZN(mixCol_out[124]) );
  AND2_X1 U945 ( .A1(sBox_out[124]), .A2(final_round), .ZN(n715) );
  AND2_X1 U946 ( .A1(mixCol_out_temp[124]), .A2(n772), .ZN(n714) );
  OR2_X1 U947 ( .A1(n716), .A2(n717), .ZN(mixCol_out[123]) );
  AND2_X1 U948 ( .A1(sBox_out[123]), .A2(final_round), .ZN(n717) );
  AND2_X1 U949 ( .A1(mixCol_out_temp[123]), .A2(n772), .ZN(n716) );
  OR2_X1 U950 ( .A1(n718), .A2(n719), .ZN(mixCol_out[122]) );
  AND2_X1 U951 ( .A1(sBox_out[122]), .A2(final_round), .ZN(n719) );
  AND2_X1 U952 ( .A1(mixCol_out_temp[122]), .A2(n772), .ZN(n718) );
  OR2_X1 U953 ( .A1(n720), .A2(n721), .ZN(mixCol_out[121]) );
  AND2_X1 U954 ( .A1(sBox_out[121]), .A2(final_round), .ZN(n721) );
  AND2_X1 U955 ( .A1(mixCol_out_temp[121]), .A2(n772), .ZN(n720) );
  OR2_X1 U956 ( .A1(n722), .A2(n723), .ZN(mixCol_out[120]) );
  AND2_X1 U957 ( .A1(sBox_out[120]), .A2(final_round), .ZN(n723) );
  AND2_X1 U958 ( .A1(mixCol_out_temp[120]), .A2(n772), .ZN(n722) );
  OR2_X1 U959 ( .A1(n724), .A2(n725), .ZN(mixCol_out[11]) );
  AND2_X1 U960 ( .A1(sBox_out[11]), .A2(final_round), .ZN(n725) );
  AND2_X1 U961 ( .A1(mixCol_out_temp[11]), .A2(n772), .ZN(n724) );
  OR2_X1 U962 ( .A1(n726), .A2(n727), .ZN(mixCol_out[119]) );
  AND2_X1 U963 ( .A1(sBox_out[119]), .A2(final_round), .ZN(n727) );
  AND2_X1 U964 ( .A1(mixCol_out_temp[119]), .A2(n772), .ZN(n726) );
  OR2_X1 U965 ( .A1(n728), .A2(n729), .ZN(mixCol_out[118]) );
  AND2_X1 U966 ( .A1(sBox_out[118]), .A2(final_round), .ZN(n729) );
  AND2_X1 U967 ( .A1(mixCol_out_temp[118]), .A2(n772), .ZN(n728) );
  OR2_X1 U968 ( .A1(n730), .A2(n731), .ZN(mixCol_out[117]) );
  AND2_X1 U969 ( .A1(sBox_out[117]), .A2(final_round), .ZN(n731) );
  AND2_X1 U970 ( .A1(mixCol_out_temp[117]), .A2(n772), .ZN(n730) );
  OR2_X1 U971 ( .A1(n732), .A2(n733), .ZN(mixCol_out[116]) );
  AND2_X1 U972 ( .A1(sBox_out[116]), .A2(final_round), .ZN(n733) );
  AND2_X1 U973 ( .A1(mixCol_out_temp[116]), .A2(n772), .ZN(n732) );
  OR2_X1 U974 ( .A1(n734), .A2(n735), .ZN(mixCol_out[115]) );
  AND2_X1 U975 ( .A1(sBox_out[115]), .A2(final_round), .ZN(n735) );
  AND2_X1 U976 ( .A1(mixCol_out_temp[115]), .A2(n773), .ZN(n734) );
  OR2_X1 U977 ( .A1(n736), .A2(n737), .ZN(mixCol_out[114]) );
  AND2_X1 U978 ( .A1(sBox_out[114]), .A2(final_round), .ZN(n737) );
  AND2_X1 U979 ( .A1(mixCol_out_temp[114]), .A2(n773), .ZN(n736) );
  OR2_X1 U980 ( .A1(n738), .A2(n739), .ZN(mixCol_out[113]) );
  AND2_X1 U981 ( .A1(sBox_out[113]), .A2(final_round), .ZN(n739) );
  AND2_X1 U982 ( .A1(mixCol_out_temp[113]), .A2(n773), .ZN(n738) );
  OR2_X1 U983 ( .A1(n740), .A2(n741), .ZN(mixCol_out[112]) );
  AND2_X1 U984 ( .A1(sBox_out[112]), .A2(final_round), .ZN(n741) );
  AND2_X1 U985 ( .A1(mixCol_out_temp[112]), .A2(n773), .ZN(n740) );
  OR2_X1 U986 ( .A1(n742), .A2(n743), .ZN(mixCol_out[111]) );
  AND2_X1 U987 ( .A1(sBox_out[111]), .A2(final_round), .ZN(n743) );
  AND2_X1 U988 ( .A1(mixCol_out_temp[111]), .A2(n773), .ZN(n742) );
  OR2_X1 U989 ( .A1(n744), .A2(n745), .ZN(mixCol_out[110]) );
  AND2_X1 U990 ( .A1(sBox_out[110]), .A2(final_round), .ZN(n745) );
  AND2_X1 U991 ( .A1(mixCol_out_temp[110]), .A2(n773), .ZN(n744) );
  OR2_X1 U992 ( .A1(n746), .A2(n747), .ZN(mixCol_out[10]) );
  AND2_X1 U993 ( .A1(sBox_out[10]), .A2(final_round), .ZN(n747) );
  AND2_X1 U994 ( .A1(mixCol_out_temp[10]), .A2(n773), .ZN(n746) );
  OR2_X1 U995 ( .A1(n748), .A2(n749), .ZN(mixCol_out[109]) );
  AND2_X1 U996 ( .A1(sBox_out[109]), .A2(final_round), .ZN(n749) );
  AND2_X1 U997 ( .A1(mixCol_out_temp[109]), .A2(n773), .ZN(n748) );
  OR2_X1 U998 ( .A1(n750), .A2(n751), .ZN(mixCol_out[108]) );
  AND2_X1 U999 ( .A1(sBox_out[108]), .A2(final_round), .ZN(n751) );
  AND2_X1 U1000 ( .A1(mixCol_out_temp[108]), .A2(n773), .ZN(n750) );
  OR2_X1 U1001 ( .A1(n752), .A2(n753), .ZN(mixCol_out[107]) );
  AND2_X1 U1002 ( .A1(sBox_out[107]), .A2(final_round), .ZN(n753) );
  AND2_X1 U1003 ( .A1(mixCol_out_temp[107]), .A2(n773), .ZN(n752) );
  OR2_X1 U1004 ( .A1(n754), .A2(n755), .ZN(mixCol_out[106]) );
  AND2_X1 U1005 ( .A1(sBox_out[106]), .A2(final_round), .ZN(n755) );
  AND2_X1 U1006 ( .A1(mixCol_out_temp[106]), .A2(n773), .ZN(n754) );
  OR2_X1 U1007 ( .A1(n756), .A2(n757), .ZN(mixCol_out[105]) );
  AND2_X1 U1008 ( .A1(sBox_out[105]), .A2(final_round), .ZN(n757) );
  AND2_X1 U1009 ( .A1(mixCol_out_temp[105]), .A2(n770), .ZN(n756) );
  OR2_X1 U1010 ( .A1(n758), .A2(n759), .ZN(mixCol_out[104]) );
  AND2_X1 U1011 ( .A1(sBox_out[104]), .A2(final_round), .ZN(n759) );
  AND2_X1 U1012 ( .A1(mixCol_out_temp[104]), .A2(n771), .ZN(n758) );
  OR2_X1 U1013 ( .A1(n760), .A2(n761), .ZN(mixCol_out[103]) );
  AND2_X1 U1014 ( .A1(sBox_out[103]), .A2(final_round), .ZN(n761) );
  AND2_X1 U1015 ( .A1(mixCol_out_temp[103]), .A2(n773), .ZN(n760) );
  OR2_X1 U1016 ( .A1(n762), .A2(n763), .ZN(mixCol_out[102]) );
  AND2_X1 U1017 ( .A1(sBox_out[102]), .A2(final_round), .ZN(n763) );
  AND2_X1 U1018 ( .A1(mixCol_out_temp[102]), .A2(n772), .ZN(n762) );
  OR2_X1 U1019 ( .A1(n764), .A2(n765), .ZN(mixCol_out[101]) );
  AND2_X1 U1020 ( .A1(sBox_out[101]), .A2(final_round), .ZN(n765) );
  AND2_X1 U1021 ( .A1(mixCol_out_temp[101]), .A2(n770), .ZN(n764) );
  OR2_X1 U1022 ( .A1(n766), .A2(n767), .ZN(mixCol_out[100]) );
  AND2_X1 U1023 ( .A1(sBox_out[100]), .A2(final_round), .ZN(n767) );
  AND2_X1 U1024 ( .A1(mixCol_out_temp[100]), .A2(n771), .ZN(n766) );
  OR2_X1 U1025 ( .A1(n768), .A2(n769), .ZN(mixCol_out[0]) );
  AND2_X1 U1026 ( .A1(sBox_out[0]), .A2(final_round), .ZN(n769) );
  AND2_X1 U1027 ( .A1(mixCol_out_temp[0]), .A2(n773), .ZN(n768) );
  INV_X1 U1028 ( .A(final_round), .ZN(n770) );
  INV_X1 U1029 ( .A(final_round), .ZN(n771) );
  INV_X1 U1030 ( .A(final_round), .ZN(n772) );
  INV_X1 U1031 ( .A(final_round), .ZN(n773) );
endmodule

//done
