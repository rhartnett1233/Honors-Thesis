module addRoundKey ( data, key, out );
  input [127:0] data;
  input [127:0] key;
  //input_done

  output [127:0] out;
  //output_done

  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512;
  //wire_done

  INV_X1 U1 ( .A(n452), .ZN(n1) );
  INV_X1 U2 ( .A(data[127]), .ZN(n2) );
  INV_X1 U3 ( .A(n454), .ZN(n3) );
  INV_X1 U4 ( .A(data[126]), .ZN(n4) );
  INV_X1 U5 ( .A(n456), .ZN(n5) );
  INV_X1 U6 ( .A(data[125]), .ZN(n6) );
  INV_X1 U7 ( .A(n458), .ZN(n7) );
  INV_X1 U8 ( .A(data[124]), .ZN(n8) );
  INV_X1 U9 ( .A(n460), .ZN(n9) );
  INV_X1 U10 ( .A(data[123]), .ZN(n10) );
  INV_X1 U11 ( .A(n462), .ZN(n11) );
  INV_X1 U12 ( .A(data[122]), .ZN(n12) );
  INV_X1 U13 ( .A(n464), .ZN(n13) );
  INV_X1 U14 ( .A(data[121]), .ZN(n14) );
  INV_X1 U15 ( .A(n466), .ZN(n15) );
  INV_X1 U16 ( .A(data[120]), .ZN(n16) );
  INV_X1 U17 ( .A(n470), .ZN(n17) );
  INV_X1 U18 ( .A(data[119]), .ZN(n18) );
  INV_X1 U19 ( .A(n472), .ZN(n19) );
  INV_X1 U20 ( .A(data[118]), .ZN(n20) );
  INV_X1 U21 ( .A(n474), .ZN(n21) );
  INV_X1 U22 ( .A(data[117]), .ZN(n22) );
  INV_X1 U23 ( .A(n476), .ZN(n23) );
  INV_X1 U24 ( .A(data[116]), .ZN(n24) );
  INV_X1 U25 ( .A(n478), .ZN(n25) );
  INV_X1 U26 ( .A(data[115]), .ZN(n26) );
  INV_X1 U27 ( .A(n480), .ZN(n27) );
  INV_X1 U28 ( .A(data[114]), .ZN(n28) );
  INV_X1 U29 ( .A(n482), .ZN(n29) );
  INV_X1 U30 ( .A(data[113]), .ZN(n30) );
  INV_X1 U31 ( .A(n484), .ZN(n31) );
  INV_X1 U32 ( .A(data[112]), .ZN(n32) );
  INV_X1 U33 ( .A(n486), .ZN(n33) );
  INV_X1 U34 ( .A(data[111]), .ZN(n34) );
  INV_X1 U35 ( .A(n488), .ZN(n35) );
  INV_X1 U36 ( .A(data[110]), .ZN(n36) );
  INV_X1 U37 ( .A(n492), .ZN(n37) );
  INV_X1 U38 ( .A(data[109]), .ZN(n38) );
  INV_X1 U39 ( .A(n494), .ZN(n39) );
  INV_X1 U40 ( .A(data[108]), .ZN(n40) );
  INV_X1 U41 ( .A(n496), .ZN(n41) );
  INV_X1 U42 ( .A(data[107]), .ZN(n42) );
  INV_X1 U43 ( .A(n498), .ZN(n43) );
  INV_X1 U44 ( .A(data[106]), .ZN(n44) );
  INV_X1 U45 ( .A(n500), .ZN(n45) );
  INV_X1 U46 ( .A(data[105]), .ZN(n46) );
  INV_X1 U47 ( .A(n502), .ZN(n47) );
  INV_X1 U48 ( .A(data[104]), .ZN(n48) );
  INV_X1 U49 ( .A(n504), .ZN(n49) );
  INV_X1 U50 ( .A(data[103]), .ZN(n50) );
  INV_X1 U51 ( .A(n506), .ZN(n51) );
  INV_X1 U52 ( .A(data[102]), .ZN(n52) );
  INV_X1 U53 ( .A(n508), .ZN(n53) );
  INV_X1 U54 ( .A(data[101]), .ZN(n54) );
  INV_X1 U55 ( .A(n510), .ZN(n55) );
  INV_X1 U56 ( .A(data[100]), .ZN(n56) );
  INV_X1 U57 ( .A(n260), .ZN(n57) );
  INV_X1 U58 ( .A(data[99]), .ZN(n58) );
  INV_X1 U59 ( .A(n262), .ZN(n59) );
  INV_X1 U60 ( .A(data[98]), .ZN(n60) );
  INV_X1 U61 ( .A(n264), .ZN(n61) );
  INV_X1 U62 ( .A(data[97]), .ZN(n62) );
  INV_X1 U63 ( .A(n266), .ZN(n63) );
  INV_X1 U64 ( .A(data[96]), .ZN(n64) );
  INV_X1 U65 ( .A(n268), .ZN(n65) );
  INV_X1 U66 ( .A(data[95]), .ZN(n66) );
  INV_X1 U67 ( .A(n270), .ZN(n67) );
  INV_X1 U68 ( .A(data[94]), .ZN(n68) );
  INV_X1 U69 ( .A(n272), .ZN(n69) );
  INV_X1 U70 ( .A(data[93]), .ZN(n70) );
  INV_X1 U71 ( .A(n274), .ZN(n71) );
  INV_X1 U72 ( .A(data[92]), .ZN(n72) );
  INV_X1 U73 ( .A(n276), .ZN(n73) );
  INV_X1 U74 ( .A(data[91]), .ZN(n74) );
  INV_X1 U75 ( .A(n278), .ZN(n75) );
  INV_X1 U76 ( .A(data[90]), .ZN(n76) );
  INV_X1 U77 ( .A(n282), .ZN(n77) );
  INV_X1 U78 ( .A(data[89]), .ZN(n78) );
  INV_X1 U79 ( .A(n284), .ZN(n79) );
  INV_X1 U80 ( .A(data[88]), .ZN(n80) );
  INV_X1 U81 ( .A(n286), .ZN(n81) );
  INV_X1 U82 ( .A(data[87]), .ZN(n82) );
  INV_X1 U83 ( .A(n288), .ZN(n83) );
  INV_X1 U84 ( .A(data[86]), .ZN(n84) );
  INV_X1 U85 ( .A(n290), .ZN(n85) );
  INV_X1 U86 ( .A(data[85]), .ZN(n86) );
  INV_X1 U87 ( .A(n292), .ZN(n87) );
  INV_X1 U88 ( .A(data[84]), .ZN(n88) );
  INV_X1 U89 ( .A(n294), .ZN(n89) );
  INV_X1 U90 ( .A(data[83]), .ZN(n90) );
  INV_X1 U91 ( .A(n296), .ZN(n91) );
  INV_X1 U92 ( .A(data[82]), .ZN(n92) );
  INV_X1 U93 ( .A(n298), .ZN(n93) );
  INV_X1 U94 ( .A(data[81]), .ZN(n94) );
  INV_X1 U95 ( .A(n300), .ZN(n95) );
  INV_X1 U96 ( .A(data[80]), .ZN(n96) );
  INV_X1 U97 ( .A(n304), .ZN(n97) );
  INV_X1 U98 ( .A(data[79]), .ZN(n98) );
  INV_X1 U99 ( .A(n306), .ZN(n99) );
  INV_X1 U100 ( .A(data[78]), .ZN(n100) );
  INV_X1 U101 ( .A(n308), .ZN(n101) );
  INV_X1 U102 ( .A(data[77]), .ZN(n102) );
  INV_X1 U103 ( .A(n310), .ZN(n103) );
  INV_X1 U104 ( .A(data[76]), .ZN(n104) );
  INV_X1 U105 ( .A(n312), .ZN(n105) );
  INV_X1 U106 ( .A(data[75]), .ZN(n106) );
  INV_X1 U107 ( .A(n314), .ZN(n107) );
  INV_X1 U108 ( .A(data[74]), .ZN(n108) );
  INV_X1 U109 ( .A(n316), .ZN(n109) );
  INV_X1 U110 ( .A(data[73]), .ZN(n110) );
  INV_X1 U111 ( .A(n318), .ZN(n111) );
  INV_X1 U112 ( .A(data[72]), .ZN(n112) );
  INV_X1 U113 ( .A(n320), .ZN(n113) );
  INV_X1 U114 ( .A(data[71]), .ZN(n114) );
  INV_X1 U115 ( .A(n322), .ZN(n115) );
  INV_X1 U116 ( .A(data[70]), .ZN(n116) );
  INV_X1 U117 ( .A(n326), .ZN(n117) );
  INV_X1 U118 ( .A(data[69]), .ZN(n118) );
  INV_X1 U119 ( .A(n328), .ZN(n119) );
  INV_X1 U120 ( .A(data[68]), .ZN(n120) );
  INV_X1 U121 ( .A(n330), .ZN(n121) );
  INV_X1 U122 ( .A(data[67]), .ZN(n122) );
  INV_X1 U123 ( .A(n332), .ZN(n123) );
  INV_X1 U124 ( .A(data[66]), .ZN(n124) );
  INV_X1 U125 ( .A(n334), .ZN(n125) );
  INV_X1 U126 ( .A(data[65]), .ZN(n126) );
  INV_X1 U127 ( .A(n336), .ZN(n127) );
  INV_X1 U128 ( .A(data[64]), .ZN(n128) );
  INV_X1 U129 ( .A(n338), .ZN(n129) );
  INV_X1 U130 ( .A(data[63]), .ZN(n130) );
  INV_X1 U131 ( .A(n340), .ZN(n131) );
  INV_X1 U132 ( .A(data[62]), .ZN(n132) );
  INV_X1 U133 ( .A(n342), .ZN(n133) );
  INV_X1 U134 ( .A(data[61]), .ZN(n134) );
  INV_X1 U135 ( .A(n344), .ZN(n135) );
  INV_X1 U136 ( .A(data[60]), .ZN(n136) );
  INV_X1 U137 ( .A(n348), .ZN(n137) );
  INV_X1 U138 ( .A(data[59]), .ZN(n138) );
  INV_X1 U139 ( .A(n350), .ZN(n139) );
  INV_X1 U140 ( .A(data[58]), .ZN(n140) );
  INV_X1 U141 ( .A(n352), .ZN(n141) );
  INV_X1 U142 ( .A(data[57]), .ZN(n142) );
  INV_X1 U143 ( .A(n354), .ZN(n143) );
  INV_X1 U144 ( .A(data[56]), .ZN(n144) );
  INV_X1 U145 ( .A(n356), .ZN(n145) );
  INV_X1 U146 ( .A(data[55]), .ZN(n146) );
  INV_X1 U147 ( .A(n358), .ZN(n147) );
  INV_X1 U148 ( .A(data[54]), .ZN(n148) );
  INV_X1 U149 ( .A(n360), .ZN(n149) );
  INV_X1 U150 ( .A(data[53]), .ZN(n150) );
  INV_X1 U151 ( .A(n362), .ZN(n151) );
  INV_X1 U152 ( .A(data[52]), .ZN(n152) );
  INV_X1 U153 ( .A(n364), .ZN(n153) );
  INV_X1 U154 ( .A(data[51]), .ZN(n154) );
  INV_X1 U155 ( .A(n366), .ZN(n155) );
  INV_X1 U156 ( .A(data[50]), .ZN(n156) );
  INV_X1 U157 ( .A(n370), .ZN(n157) );
  INV_X1 U158 ( .A(data[49]), .ZN(n158) );
  INV_X1 U159 ( .A(n372), .ZN(n159) );
  INV_X1 U160 ( .A(data[48]), .ZN(n160) );
  INV_X1 U161 ( .A(n374), .ZN(n161) );
  INV_X1 U162 ( .A(data[47]), .ZN(n162) );
  INV_X1 U163 ( .A(n376), .ZN(n163) );
  INV_X1 U164 ( .A(data[46]), .ZN(n164) );
  INV_X1 U165 ( .A(n378), .ZN(n165) );
  INV_X1 U166 ( .A(data[45]), .ZN(n166) );
  INV_X1 U167 ( .A(n380), .ZN(n167) );
  INV_X1 U168 ( .A(data[44]), .ZN(n168) );
  INV_X1 U169 ( .A(n382), .ZN(n169) );
  INV_X1 U170 ( .A(data[43]), .ZN(n170) );
  INV_X1 U171 ( .A(n384), .ZN(n171) );
  INV_X1 U172 ( .A(data[42]), .ZN(n172) );
  INV_X1 U173 ( .A(n386), .ZN(n173) );
  INV_X1 U174 ( .A(data[41]), .ZN(n174) );
  INV_X1 U175 ( .A(n388), .ZN(n175) );
  INV_X1 U176 ( .A(data[40]), .ZN(n176) );
  INV_X1 U177 ( .A(n392), .ZN(n177) );
  INV_X1 U178 ( .A(data[39]), .ZN(n178) );
  INV_X1 U179 ( .A(n394), .ZN(n179) );
  INV_X1 U180 ( .A(data[38]), .ZN(n180) );
  INV_X1 U181 ( .A(n396), .ZN(n181) );
  INV_X1 U182 ( .A(data[37]), .ZN(n182) );
  INV_X1 U183 ( .A(n398), .ZN(n183) );
  INV_X1 U184 ( .A(data[36]), .ZN(n184) );
  INV_X1 U185 ( .A(n400), .ZN(n185) );
  INV_X1 U186 ( .A(data[35]), .ZN(n186) );
  INV_X1 U187 ( .A(n402), .ZN(n187) );
  INV_X1 U188 ( .A(data[34]), .ZN(n188) );
  INV_X1 U189 ( .A(n404), .ZN(n189) );
  INV_X1 U190 ( .A(data[33]), .ZN(n190) );
  INV_X1 U191 ( .A(n406), .ZN(n191) );
  INV_X1 U192 ( .A(data[32]), .ZN(n192) );
  INV_X1 U193 ( .A(n408), .ZN(n193) );
  INV_X1 U194 ( .A(data[31]), .ZN(n194) );
  INV_X1 U195 ( .A(n410), .ZN(n195) );
  INV_X1 U196 ( .A(data[30]), .ZN(n196) );
  INV_X1 U197 ( .A(n414), .ZN(n197) );
  INV_X1 U198 ( .A(data[29]), .ZN(n198) );
  INV_X1 U199 ( .A(n416), .ZN(n199) );
  INV_X1 U200 ( .A(data[28]), .ZN(n200) );
  INV_X1 U201 ( .A(n418), .ZN(n201) );
  INV_X1 U202 ( .A(data[27]), .ZN(n202) );
  INV_X1 U203 ( .A(n420), .ZN(n203) );
  INV_X1 U204 ( .A(data[26]), .ZN(n204) );
  INV_X1 U205 ( .A(n422), .ZN(n205) );
  INV_X1 U206 ( .A(data[25]), .ZN(n206) );
  INV_X1 U207 ( .A(n424), .ZN(n207) );
  INV_X1 U208 ( .A(data[24]), .ZN(n208) );
  INV_X1 U209 ( .A(n426), .ZN(n209) );
  INV_X1 U210 ( .A(data[23]), .ZN(n210) );
  INV_X1 U211 ( .A(n428), .ZN(n211) );
  INV_X1 U212 ( .A(data[22]), .ZN(n212) );
  INV_X1 U213 ( .A(n430), .ZN(n213) );
  INV_X1 U214 ( .A(data[21]), .ZN(n214) );
  INV_X1 U215 ( .A(n432), .ZN(n215) );
  INV_X1 U216 ( .A(data[20]), .ZN(n216) );
  INV_X1 U217 ( .A(n436), .ZN(n217) );
  INV_X1 U218 ( .A(data[19]), .ZN(n218) );
  INV_X1 U219 ( .A(n438), .ZN(n219) );
  INV_X1 U220 ( .A(data[18]), .ZN(n220) );
  INV_X1 U221 ( .A(n440), .ZN(n221) );
  INV_X1 U222 ( .A(data[17]), .ZN(n222) );
  INV_X1 U223 ( .A(n442), .ZN(n223) );
  INV_X1 U224 ( .A(data[16]), .ZN(n224) );
  INV_X1 U225 ( .A(n444), .ZN(n225) );
  INV_X1 U226 ( .A(data[15]), .ZN(n226) );
  INV_X1 U227 ( .A(n446), .ZN(n227) );
  INV_X1 U228 ( .A(data[14]), .ZN(n228) );
  INV_X1 U229 ( .A(n448), .ZN(n229) );
  INV_X1 U230 ( .A(data[13]), .ZN(n230) );
  INV_X1 U231 ( .A(n450), .ZN(n231) );
  INV_X1 U232 ( .A(data[12]), .ZN(n232) );
  INV_X1 U233 ( .A(n468), .ZN(n233) );
  INV_X1 U234 ( .A(data[11]), .ZN(n234) );
  INV_X1 U235 ( .A(n490), .ZN(n235) );
  INV_X1 U236 ( .A(data[10]), .ZN(n236) );
  INV_X1 U237 ( .A(n258), .ZN(n237) );
  INV_X1 U238 ( .A(data[9]), .ZN(n238) );
  INV_X1 U239 ( .A(n280), .ZN(n239) );
  INV_X1 U240 ( .A(data[8]), .ZN(n240) );
  INV_X1 U241 ( .A(n302), .ZN(n241) );
  INV_X1 U242 ( .A(data[7]), .ZN(n242) );
  INV_X1 U243 ( .A(n324), .ZN(n243) );
  INV_X1 U244 ( .A(data[6]), .ZN(n244) );
  INV_X1 U245 ( .A(n346), .ZN(n245) );
  INV_X1 U246 ( .A(data[5]), .ZN(n246) );
  INV_X1 U247 ( .A(n368), .ZN(n247) );
  INV_X1 U248 ( .A(data[4]), .ZN(n248) );
  INV_X1 U249 ( .A(n390), .ZN(n249) );
  INV_X1 U250 ( .A(data[3]), .ZN(n250) );
  INV_X1 U251 ( .A(n412), .ZN(n251) );
  INV_X1 U252 ( .A(data[2]), .ZN(n252) );
  INV_X1 U253 ( .A(n434), .ZN(n253) );
  INV_X1 U254 ( .A(data[1]), .ZN(n254) );
  INV_X1 U255 ( .A(n512), .ZN(n255) );
  INV_X1 U256 ( .A(data[0]), .ZN(n256) );
  OR2_X1 U257 ( .A1(n257), .A2(n237), .ZN(out[9]) );
  OR2_X1 U258 ( .A1(n238), .A2(key[9]), .ZN(n258) );
  AND2_X1 U259 ( .A1(key[9]), .A2(n238), .ZN(n257) );
  OR2_X1 U260 ( .A1(n259), .A2(n57), .ZN(out[99]) );
  OR2_X1 U261 ( .A1(n58), .A2(key[99]), .ZN(n260) );
  AND2_X1 U262 ( .A1(key[99]), .A2(n58), .ZN(n259) );
  OR2_X1 U263 ( .A1(n261), .A2(n59), .ZN(out[98]) );
  OR2_X1 U264 ( .A1(n60), .A2(key[98]), .ZN(n262) );
  AND2_X1 U265 ( .A1(key[98]), .A2(n60), .ZN(n261) );
  OR2_X1 U266 ( .A1(n263), .A2(n61), .ZN(out[97]) );
  OR2_X1 U267 ( .A1(n62), .A2(key[97]), .ZN(n264) );
  AND2_X1 U268 ( .A1(key[97]), .A2(n62), .ZN(n263) );
  OR2_X1 U269 ( .A1(n265), .A2(n63), .ZN(out[96]) );
  OR2_X1 U270 ( .A1(n64), .A2(key[96]), .ZN(n266) );
  AND2_X1 U271 ( .A1(key[96]), .A2(n64), .ZN(n265) );
  OR2_X1 U272 ( .A1(n267), .A2(n65), .ZN(out[95]) );
  OR2_X1 U273 ( .A1(n66), .A2(key[95]), .ZN(n268) );
  AND2_X1 U274 ( .A1(key[95]), .A2(n66), .ZN(n267) );
  OR2_X1 U275 ( .A1(n269), .A2(n67), .ZN(out[94]) );
  OR2_X1 U276 ( .A1(n68), .A2(key[94]), .ZN(n270) );
  AND2_X1 U277 ( .A1(key[94]), .A2(n68), .ZN(n269) );
  OR2_X1 U278 ( .A1(n271), .A2(n69), .ZN(out[93]) );
  OR2_X1 U279 ( .A1(n70), .A2(key[93]), .ZN(n272) );
  AND2_X1 U280 ( .A1(key[93]), .A2(n70), .ZN(n271) );
  OR2_X1 U281 ( .A1(n273), .A2(n71), .ZN(out[92]) );
  OR2_X1 U282 ( .A1(n72), .A2(key[92]), .ZN(n274) );
  AND2_X1 U283 ( .A1(key[92]), .A2(n72), .ZN(n273) );
  OR2_X1 U284 ( .A1(n275), .A2(n73), .ZN(out[91]) );
  OR2_X1 U285 ( .A1(n74), .A2(key[91]), .ZN(n276) );
  AND2_X1 U286 ( .A1(key[91]), .A2(n74), .ZN(n275) );
  OR2_X1 U287 ( .A1(n277), .A2(n75), .ZN(out[90]) );
  OR2_X1 U288 ( .A1(n76), .A2(key[90]), .ZN(n278) );
  AND2_X1 U289 ( .A1(key[90]), .A2(n76), .ZN(n277) );
  OR2_X1 U290 ( .A1(n279), .A2(n239), .ZN(out[8]) );
  OR2_X1 U291 ( .A1(n240), .A2(key[8]), .ZN(n280) );
  AND2_X1 U292 ( .A1(key[8]), .A2(n240), .ZN(n279) );
  OR2_X1 U293 ( .A1(n281), .A2(n77), .ZN(out[89]) );
  OR2_X1 U294 ( .A1(n78), .A2(key[89]), .ZN(n282) );
  AND2_X1 U295 ( .A1(key[89]), .A2(n78), .ZN(n281) );
  OR2_X1 U296 ( .A1(n283), .A2(n79), .ZN(out[88]) );
  OR2_X1 U297 ( .A1(n80), .A2(key[88]), .ZN(n284) );
  AND2_X1 U298 ( .A1(key[88]), .A2(n80), .ZN(n283) );
  OR2_X1 U299 ( .A1(n285), .A2(n81), .ZN(out[87]) );
  OR2_X1 U300 ( .A1(n82), .A2(key[87]), .ZN(n286) );
  AND2_X1 U301 ( .A1(key[87]), .A2(n82), .ZN(n285) );
  OR2_X1 U302 ( .A1(n287), .A2(n83), .ZN(out[86]) );
  OR2_X1 U303 ( .A1(n84), .A2(key[86]), .ZN(n288) );
  AND2_X1 U304 ( .A1(key[86]), .A2(n84), .ZN(n287) );
  OR2_X1 U305 ( .A1(n289), .A2(n85), .ZN(out[85]) );
  OR2_X1 U306 ( .A1(n86), .A2(key[85]), .ZN(n290) );
  AND2_X1 U307 ( .A1(key[85]), .A2(n86), .ZN(n289) );
  OR2_X1 U308 ( .A1(n291), .A2(n87), .ZN(out[84]) );
  OR2_X1 U309 ( .A1(n88), .A2(key[84]), .ZN(n292) );
  AND2_X1 U310 ( .A1(key[84]), .A2(n88), .ZN(n291) );
  OR2_X1 U311 ( .A1(n293), .A2(n89), .ZN(out[83]) );
  OR2_X1 U312 ( .A1(n90), .A2(key[83]), .ZN(n294) );
  AND2_X1 U313 ( .A1(key[83]), .A2(n90), .ZN(n293) );
  OR2_X1 U314 ( .A1(n295), .A2(n91), .ZN(out[82]) );
  OR2_X1 U315 ( .A1(n92), .A2(key[82]), .ZN(n296) );
  AND2_X1 U316 ( .A1(key[82]), .A2(n92), .ZN(n295) );
  OR2_X1 U317 ( .A1(n297), .A2(n93), .ZN(out[81]) );
  OR2_X1 U318 ( .A1(n94), .A2(key[81]), .ZN(n298) );
  AND2_X1 U319 ( .A1(key[81]), .A2(n94), .ZN(n297) );
  OR2_X1 U320 ( .A1(n299), .A2(n95), .ZN(out[80]) );
  OR2_X1 U321 ( .A1(n96), .A2(key[80]), .ZN(n300) );
  AND2_X1 U322 ( .A1(key[80]), .A2(n96), .ZN(n299) );
  OR2_X1 U323 ( .A1(n301), .A2(n241), .ZN(out[7]) );
  OR2_X1 U324 ( .A1(n242), .A2(key[7]), .ZN(n302) );
  AND2_X1 U325 ( .A1(key[7]), .A2(n242), .ZN(n301) );
  OR2_X1 U326 ( .A1(n303), .A2(n97), .ZN(out[79]) );
  OR2_X1 U327 ( .A1(n98), .A2(key[79]), .ZN(n304) );
  AND2_X1 U328 ( .A1(key[79]), .A2(n98), .ZN(n303) );
  OR2_X1 U329 ( .A1(n305), .A2(n99), .ZN(out[78]) );
  OR2_X1 U330 ( .A1(n100), .A2(key[78]), .ZN(n306) );
  AND2_X1 U331 ( .A1(key[78]), .A2(n100), .ZN(n305) );
  OR2_X1 U332 ( .A1(n307), .A2(n101), .ZN(out[77]) );
  OR2_X1 U333 ( .A1(n102), .A2(key[77]), .ZN(n308) );
  AND2_X1 U334 ( .A1(key[77]), .A2(n102), .ZN(n307) );
  OR2_X1 U335 ( .A1(n309), .A2(n103), .ZN(out[76]) );
  OR2_X1 U336 ( .A1(n104), .A2(key[76]), .ZN(n310) );
  AND2_X1 U337 ( .A1(key[76]), .A2(n104), .ZN(n309) );
  OR2_X1 U338 ( .A1(n311), .A2(n105), .ZN(out[75]) );
  OR2_X1 U339 ( .A1(n106), .A2(key[75]), .ZN(n312) );
  AND2_X1 U340 ( .A1(key[75]), .A2(n106), .ZN(n311) );
  OR2_X1 U341 ( .A1(n313), .A2(n107), .ZN(out[74]) );
  OR2_X1 U342 ( .A1(n108), .A2(key[74]), .ZN(n314) );
  AND2_X1 U343 ( .A1(key[74]), .A2(n108), .ZN(n313) );
  OR2_X1 U344 ( .A1(n315), .A2(n109), .ZN(out[73]) );
  OR2_X1 U345 ( .A1(n110), .A2(key[73]), .ZN(n316) );
  AND2_X1 U346 ( .A1(key[73]), .A2(n110), .ZN(n315) );
  OR2_X1 U347 ( .A1(n317), .A2(n111), .ZN(out[72]) );
  OR2_X1 U348 ( .A1(n112), .A2(key[72]), .ZN(n318) );
  AND2_X1 U349 ( .A1(key[72]), .A2(n112), .ZN(n317) );
  OR2_X1 U350 ( .A1(n319), .A2(n113), .ZN(out[71]) );
  OR2_X1 U351 ( .A1(n114), .A2(key[71]), .ZN(n320) );
  AND2_X1 U352 ( .A1(key[71]), .A2(n114), .ZN(n319) );
  OR2_X1 U353 ( .A1(n321), .A2(n115), .ZN(out[70]) );
  OR2_X1 U354 ( .A1(n116), .A2(key[70]), .ZN(n322) );
  AND2_X1 U355 ( .A1(key[70]), .A2(n116), .ZN(n321) );
  OR2_X1 U356 ( .A1(n323), .A2(n243), .ZN(out[6]) );
  OR2_X1 U357 ( .A1(n244), .A2(key[6]), .ZN(n324) );
  AND2_X1 U358 ( .A1(key[6]), .A2(n244), .ZN(n323) );
  OR2_X1 U359 ( .A1(n325), .A2(n117), .ZN(out[69]) );
  OR2_X1 U360 ( .A1(n118), .A2(key[69]), .ZN(n326) );
  AND2_X1 U361 ( .A1(key[69]), .A2(n118), .ZN(n325) );
  OR2_X1 U362 ( .A1(n327), .A2(n119), .ZN(out[68]) );
  OR2_X1 U363 ( .A1(n120), .A2(key[68]), .ZN(n328) );
  AND2_X1 U364 ( .A1(key[68]), .A2(n120), .ZN(n327) );
  OR2_X1 U365 ( .A1(n329), .A2(n121), .ZN(out[67]) );
  OR2_X1 U366 ( .A1(n122), .A2(key[67]), .ZN(n330) );
  AND2_X1 U367 ( .A1(key[67]), .A2(n122), .ZN(n329) );
  OR2_X1 U368 ( .A1(n331), .A2(n123), .ZN(out[66]) );
  OR2_X1 U369 ( .A1(n124), .A2(key[66]), .ZN(n332) );
  AND2_X1 U370 ( .A1(key[66]), .A2(n124), .ZN(n331) );
  OR2_X1 U371 ( .A1(n333), .A2(n125), .ZN(out[65]) );
  OR2_X1 U372 ( .A1(n126), .A2(key[65]), .ZN(n334) );
  AND2_X1 U373 ( .A1(key[65]), .A2(n126), .ZN(n333) );
  OR2_X1 U374 ( .A1(n335), .A2(n127), .ZN(out[64]) );
  OR2_X1 U375 ( .A1(n128), .A2(key[64]), .ZN(n336) );
  AND2_X1 U376 ( .A1(key[64]), .A2(n128), .ZN(n335) );
  OR2_X1 U377 ( .A1(n337), .A2(n129), .ZN(out[63]) );
  OR2_X1 U378 ( .A1(n130), .A2(key[63]), .ZN(n338) );
  AND2_X1 U379 ( .A1(key[63]), .A2(n130), .ZN(n337) );
  OR2_X1 U380 ( .A1(n339), .A2(n131), .ZN(out[62]) );
  OR2_X1 U381 ( .A1(n132), .A2(key[62]), .ZN(n340) );
  AND2_X1 U382 ( .A1(key[62]), .A2(n132), .ZN(n339) );
  OR2_X1 U383 ( .A1(n341), .A2(n133), .ZN(out[61]) );
  OR2_X1 U384 ( .A1(n134), .A2(key[61]), .ZN(n342) );
  AND2_X1 U385 ( .A1(key[61]), .A2(n134), .ZN(n341) );
  OR2_X1 U386 ( .A1(n343), .A2(n135), .ZN(out[60]) );
  OR2_X1 U387 ( .A1(n136), .A2(key[60]), .ZN(n344) );
  AND2_X1 U388 ( .A1(key[60]), .A2(n136), .ZN(n343) );
  OR2_X1 U389 ( .A1(n345), .A2(n245), .ZN(out[5]) );
  OR2_X1 U390 ( .A1(n246), .A2(key[5]), .ZN(n346) );
  AND2_X1 U391 ( .A1(key[5]), .A2(n246), .ZN(n345) );
  OR2_X1 U392 ( .A1(n347), .A2(n137), .ZN(out[59]) );
  OR2_X1 U393 ( .A1(n138), .A2(key[59]), .ZN(n348) );
  AND2_X1 U394 ( .A1(key[59]), .A2(n138), .ZN(n347) );
  OR2_X1 U395 ( .A1(n349), .A2(n139), .ZN(out[58]) );
  OR2_X1 U396 ( .A1(n140), .A2(key[58]), .ZN(n350) );
  AND2_X1 U397 ( .A1(key[58]), .A2(n140), .ZN(n349) );
  OR2_X1 U398 ( .A1(n351), .A2(n141), .ZN(out[57]) );
  OR2_X1 U399 ( .A1(n142), .A2(key[57]), .ZN(n352) );
  AND2_X1 U400 ( .A1(key[57]), .A2(n142), .ZN(n351) );
  OR2_X1 U401 ( .A1(n353), .A2(n143), .ZN(out[56]) );
  OR2_X1 U402 ( .A1(n144), .A2(key[56]), .ZN(n354) );
  AND2_X1 U403 ( .A1(key[56]), .A2(n144), .ZN(n353) );
  OR2_X1 U404 ( .A1(n355), .A2(n145), .ZN(out[55]) );
  OR2_X1 U405 ( .A1(n146), .A2(key[55]), .ZN(n356) );
  AND2_X1 U406 ( .A1(key[55]), .A2(n146), .ZN(n355) );
  OR2_X1 U407 ( .A1(n357), .A2(n147), .ZN(out[54]) );
  OR2_X1 U408 ( .A1(n148), .A2(key[54]), .ZN(n358) );
  AND2_X1 U409 ( .A1(key[54]), .A2(n148), .ZN(n357) );
  OR2_X1 U410 ( .A1(n359), .A2(n149), .ZN(out[53]) );
  OR2_X1 U411 ( .A1(n150), .A2(key[53]), .ZN(n360) );
  AND2_X1 U412 ( .A1(key[53]), .A2(n150), .ZN(n359) );
  OR2_X1 U413 ( .A1(n361), .A2(n151), .ZN(out[52]) );
  OR2_X1 U414 ( .A1(n152), .A2(key[52]), .ZN(n362) );
  AND2_X1 U415 ( .A1(key[52]), .A2(n152), .ZN(n361) );
  OR2_X1 U416 ( .A1(n363), .A2(n153), .ZN(out[51]) );
  OR2_X1 U417 ( .A1(n154), .A2(key[51]), .ZN(n364) );
  AND2_X1 U418 ( .A1(key[51]), .A2(n154), .ZN(n363) );
  OR2_X1 U419 ( .A1(n365), .A2(n155), .ZN(out[50]) );
  OR2_X1 U420 ( .A1(n156), .A2(key[50]), .ZN(n366) );
  AND2_X1 U421 ( .A1(key[50]), .A2(n156), .ZN(n365) );
  OR2_X1 U422 ( .A1(n367), .A2(n247), .ZN(out[4]) );
  OR2_X1 U423 ( .A1(n248), .A2(key[4]), .ZN(n368) );
  AND2_X1 U424 ( .A1(key[4]), .A2(n248), .ZN(n367) );
  OR2_X1 U425 ( .A1(n369), .A2(n157), .ZN(out[49]) );
  OR2_X1 U426 ( .A1(n158), .A2(key[49]), .ZN(n370) );
  AND2_X1 U427 ( .A1(key[49]), .A2(n158), .ZN(n369) );
  OR2_X1 U428 ( .A1(n371), .A2(n159), .ZN(out[48]) );
  OR2_X1 U429 ( .A1(n160), .A2(key[48]), .ZN(n372) );
  AND2_X1 U430 ( .A1(key[48]), .A2(n160), .ZN(n371) );
  OR2_X1 U431 ( .A1(n373), .A2(n161), .ZN(out[47]) );
  OR2_X1 U432 ( .A1(n162), .A2(key[47]), .ZN(n374) );
  AND2_X1 U433 ( .A1(key[47]), .A2(n162), .ZN(n373) );
  OR2_X1 U434 ( .A1(n375), .A2(n163), .ZN(out[46]) );
  OR2_X1 U435 ( .A1(n164), .A2(key[46]), .ZN(n376) );
  AND2_X1 U436 ( .A1(key[46]), .A2(n164), .ZN(n375) );
  OR2_X1 U437 ( .A1(n377), .A2(n165), .ZN(out[45]) );
  OR2_X1 U438 ( .A1(n166), .A2(key[45]), .ZN(n378) );
  AND2_X1 U439 ( .A1(key[45]), .A2(n166), .ZN(n377) );
  OR2_X1 U440 ( .A1(n379), .A2(n167), .ZN(out[44]) );
  OR2_X1 U441 ( .A1(n168), .A2(key[44]), .ZN(n380) );
  AND2_X1 U442 ( .A1(key[44]), .A2(n168), .ZN(n379) );
  OR2_X1 U443 ( .A1(n381), .A2(n169), .ZN(out[43]) );
  OR2_X1 U444 ( .A1(n170), .A2(key[43]), .ZN(n382) );
  AND2_X1 U445 ( .A1(key[43]), .A2(n170), .ZN(n381) );
  OR2_X1 U446 ( .A1(n383), .A2(n171), .ZN(out[42]) );
  OR2_X1 U447 ( .A1(n172), .A2(key[42]), .ZN(n384) );
  AND2_X1 U448 ( .A1(key[42]), .A2(n172), .ZN(n383) );
  OR2_X1 U449 ( .A1(n385), .A2(n173), .ZN(out[41]) );
  OR2_X1 U450 ( .A1(n174), .A2(key[41]), .ZN(n386) );
  AND2_X1 U451 ( .A1(key[41]), .A2(n174), .ZN(n385) );
  OR2_X1 U452 ( .A1(n387), .A2(n175), .ZN(out[40]) );
  OR2_X1 U453 ( .A1(n176), .A2(key[40]), .ZN(n388) );
  AND2_X1 U454 ( .A1(key[40]), .A2(n176), .ZN(n387) );
  OR2_X1 U455 ( .A1(n389), .A2(n249), .ZN(out[3]) );
  OR2_X1 U456 ( .A1(n250), .A2(key[3]), .ZN(n390) );
  AND2_X1 U457 ( .A1(key[3]), .A2(n250), .ZN(n389) );
  OR2_X1 U458 ( .A1(n391), .A2(n177), .ZN(out[39]) );
  OR2_X1 U459 ( .A1(n178), .A2(key[39]), .ZN(n392) );
  AND2_X1 U460 ( .A1(key[39]), .A2(n178), .ZN(n391) );
  OR2_X1 U461 ( .A1(n393), .A2(n179), .ZN(out[38]) );
  OR2_X1 U462 ( .A1(n180), .A2(key[38]), .ZN(n394) );
  AND2_X1 U463 ( .A1(key[38]), .A2(n180), .ZN(n393) );
  OR2_X1 U464 ( .A1(n395), .A2(n181), .ZN(out[37]) );
  OR2_X1 U465 ( .A1(n182), .A2(key[37]), .ZN(n396) );
  AND2_X1 U466 ( .A1(key[37]), .A2(n182), .ZN(n395) );
  OR2_X1 U467 ( .A1(n397), .A2(n183), .ZN(out[36]) );
  OR2_X1 U468 ( .A1(n184), .A2(key[36]), .ZN(n398) );
  AND2_X1 U469 ( .A1(key[36]), .A2(n184), .ZN(n397) );
  OR2_X1 U470 ( .A1(n399), .A2(n185), .ZN(out[35]) );
  OR2_X1 U471 ( .A1(n186), .A2(key[35]), .ZN(n400) );
  AND2_X1 U472 ( .A1(key[35]), .A2(n186), .ZN(n399) );
  OR2_X1 U473 ( .A1(n401), .A2(n187), .ZN(out[34]) );
  OR2_X1 U474 ( .A1(n188), .A2(key[34]), .ZN(n402) );
  AND2_X1 U475 ( .A1(key[34]), .A2(n188), .ZN(n401) );
  OR2_X1 U476 ( .A1(n403), .A2(n189), .ZN(out[33]) );
  OR2_X1 U477 ( .A1(n190), .A2(key[33]), .ZN(n404) );
  AND2_X1 U478 ( .A1(key[33]), .A2(n190), .ZN(n403) );
  OR2_X1 U479 ( .A1(n405), .A2(n191), .ZN(out[32]) );
  OR2_X1 U480 ( .A1(n192), .A2(key[32]), .ZN(n406) );
  AND2_X1 U481 ( .A1(key[32]), .A2(n192), .ZN(n405) );
  OR2_X1 U482 ( .A1(n407), .A2(n193), .ZN(out[31]) );
  OR2_X1 U483 ( .A1(n194), .A2(key[31]), .ZN(n408) );
  AND2_X1 U484 ( .A1(key[31]), .A2(n194), .ZN(n407) );
  OR2_X1 U485 ( .A1(n409), .A2(n195), .ZN(out[30]) );
  OR2_X1 U486 ( .A1(n196), .A2(key[30]), .ZN(n410) );
  AND2_X1 U487 ( .A1(key[30]), .A2(n196), .ZN(n409) );
  OR2_X1 U488 ( .A1(n411), .A2(n251), .ZN(out[2]) );
  OR2_X1 U489 ( .A1(n252), .A2(key[2]), .ZN(n412) );
  AND2_X1 U490 ( .A1(key[2]), .A2(n252), .ZN(n411) );
  OR2_X1 U491 ( .A1(n413), .A2(n197), .ZN(out[29]) );
  OR2_X1 U492 ( .A1(n198), .A2(key[29]), .ZN(n414) );
  AND2_X1 U493 ( .A1(key[29]), .A2(n198), .ZN(n413) );
  OR2_X1 U494 ( .A1(n415), .A2(n199), .ZN(out[28]) );
  OR2_X1 U495 ( .A1(n200), .A2(key[28]), .ZN(n416) );
  AND2_X1 U496 ( .A1(key[28]), .A2(n200), .ZN(n415) );
  OR2_X1 U497 ( .A1(n417), .A2(n201), .ZN(out[27]) );
  OR2_X1 U498 ( .A1(n202), .A2(key[27]), .ZN(n418) );
  AND2_X1 U499 ( .A1(key[27]), .A2(n202), .ZN(n417) );
  OR2_X1 U500 ( .A1(n419), .A2(n203), .ZN(out[26]) );
  OR2_X1 U501 ( .A1(n204), .A2(key[26]), .ZN(n420) );
  AND2_X1 U502 ( .A1(key[26]), .A2(n204), .ZN(n419) );
  OR2_X1 U503 ( .A1(n421), .A2(n205), .ZN(out[25]) );
  OR2_X1 U504 ( .A1(n206), .A2(key[25]), .ZN(n422) );
  AND2_X1 U505 ( .A1(key[25]), .A2(n206), .ZN(n421) );
  OR2_X1 U506 ( .A1(n423), .A2(n207), .ZN(out[24]) );
  OR2_X1 U507 ( .A1(n208), .A2(key[24]), .ZN(n424) );
  AND2_X1 U508 ( .A1(key[24]), .A2(n208), .ZN(n423) );
  OR2_X1 U509 ( .A1(n425), .A2(n209), .ZN(out[23]) );
  OR2_X1 U510 ( .A1(n210), .A2(key[23]), .ZN(n426) );
  AND2_X1 U511 ( .A1(key[23]), .A2(n210), .ZN(n425) );
  OR2_X1 U512 ( .A1(n427), .A2(n211), .ZN(out[22]) );
  OR2_X1 U513 ( .A1(n212), .A2(key[22]), .ZN(n428) );
  AND2_X1 U514 ( .A1(key[22]), .A2(n212), .ZN(n427) );
  OR2_X1 U515 ( .A1(n429), .A2(n213), .ZN(out[21]) );
  OR2_X1 U516 ( .A1(n214), .A2(key[21]), .ZN(n430) );
  AND2_X1 U517 ( .A1(key[21]), .A2(n214), .ZN(n429) );
  OR2_X1 U518 ( .A1(n431), .A2(n215), .ZN(out[20]) );
  OR2_X1 U519 ( .A1(n216), .A2(key[20]), .ZN(n432) );
  AND2_X1 U520 ( .A1(key[20]), .A2(n216), .ZN(n431) );
  OR2_X1 U521 ( .A1(n433), .A2(n253), .ZN(out[1]) );
  OR2_X1 U522 ( .A1(n254), .A2(key[1]), .ZN(n434) );
  AND2_X1 U523 ( .A1(key[1]), .A2(n254), .ZN(n433) );
  OR2_X1 U524 ( .A1(n435), .A2(n217), .ZN(out[19]) );
  OR2_X1 U525 ( .A1(n218), .A2(key[19]), .ZN(n436) );
  AND2_X1 U526 ( .A1(key[19]), .A2(n218), .ZN(n435) );
  OR2_X1 U527 ( .A1(n437), .A2(n219), .ZN(out[18]) );
  OR2_X1 U528 ( .A1(n220), .A2(key[18]), .ZN(n438) );
  AND2_X1 U529 ( .A1(key[18]), .A2(n220), .ZN(n437) );
  OR2_X1 U530 ( .A1(n439), .A2(n221), .ZN(out[17]) );
  OR2_X1 U531 ( .A1(n222), .A2(key[17]), .ZN(n440) );
  AND2_X1 U532 ( .A1(key[17]), .A2(n222), .ZN(n439) );
  OR2_X1 U533 ( .A1(n441), .A2(n223), .ZN(out[16]) );
  OR2_X1 U534 ( .A1(n224), .A2(key[16]), .ZN(n442) );
  AND2_X1 U535 ( .A1(key[16]), .A2(n224), .ZN(n441) );
  OR2_X1 U536 ( .A1(n443), .A2(n225), .ZN(out[15]) );
  OR2_X1 U537 ( .A1(n226), .A2(key[15]), .ZN(n444) );
  AND2_X1 U538 ( .A1(key[15]), .A2(n226), .ZN(n443) );
  OR2_X1 U539 ( .A1(n445), .A2(n227), .ZN(out[14]) );
  OR2_X1 U540 ( .A1(n228), .A2(key[14]), .ZN(n446) );
  AND2_X1 U541 ( .A1(key[14]), .A2(n228), .ZN(n445) );
  OR2_X1 U542 ( .A1(n447), .A2(n229), .ZN(out[13]) );
  OR2_X1 U543 ( .A1(n230), .A2(key[13]), .ZN(n448) );
  AND2_X1 U544 ( .A1(key[13]), .A2(n230), .ZN(n447) );
  OR2_X1 U545 ( .A1(n449), .A2(n231), .ZN(out[12]) );
  OR2_X1 U546 ( .A1(n232), .A2(key[12]), .ZN(n450) );
  AND2_X1 U547 ( .A1(key[12]), .A2(n232), .ZN(n449) );
  OR2_X1 U548 ( .A1(n451), .A2(n1), .ZN(out[127]) );
  OR2_X1 U549 ( .A1(n2), .A2(key[127]), .ZN(n452) );
  AND2_X1 U550 ( .A1(key[127]), .A2(n2), .ZN(n451) );
  OR2_X1 U551 ( .A1(n453), .A2(n3), .ZN(out[126]) );
  OR2_X1 U552 ( .A1(n4), .A2(key[126]), .ZN(n454) );
  AND2_X1 U553 ( .A1(key[126]), .A2(n4), .ZN(n453) );
  OR2_X1 U554 ( .A1(n455), .A2(n5), .ZN(out[125]) );
  OR2_X1 U555 ( .A1(n6), .A2(key[125]), .ZN(n456) );
  AND2_X1 U556 ( .A1(key[125]), .A2(n6), .ZN(n455) );
  OR2_X1 U557 ( .A1(n457), .A2(n7), .ZN(out[124]) );
  OR2_X1 U558 ( .A1(n8), .A2(key[124]), .ZN(n458) );
  AND2_X1 U559 ( .A1(key[124]), .A2(n8), .ZN(n457) );
  OR2_X1 U560 ( .A1(n459), .A2(n9), .ZN(out[123]) );
  OR2_X1 U561 ( .A1(n10), .A2(key[123]), .ZN(n460) );
  AND2_X1 U562 ( .A1(key[123]), .A2(n10), .ZN(n459) );
  OR2_X1 U563 ( .A1(n461), .A2(n11), .ZN(out[122]) );
  OR2_X1 U564 ( .A1(n12), .A2(key[122]), .ZN(n462) );
  AND2_X1 U565 ( .A1(key[122]), .A2(n12), .ZN(n461) );
  OR2_X1 U566 ( .A1(n463), .A2(n13), .ZN(out[121]) );
  OR2_X1 U567 ( .A1(n14), .A2(key[121]), .ZN(n464) );
  AND2_X1 U568 ( .A1(key[121]), .A2(n14), .ZN(n463) );
  OR2_X1 U569 ( .A1(n465), .A2(n15), .ZN(out[120]) );
  OR2_X1 U570 ( .A1(n16), .A2(key[120]), .ZN(n466) );
  AND2_X1 U571 ( .A1(key[120]), .A2(n16), .ZN(n465) );
  OR2_X1 U572 ( .A1(n467), .A2(n233), .ZN(out[11]) );
  OR2_X1 U573 ( .A1(n234), .A2(key[11]), .ZN(n468) );
  AND2_X1 U574 ( .A1(key[11]), .A2(n234), .ZN(n467) );
  OR2_X1 U575 ( .A1(n469), .A2(n17), .ZN(out[119]) );
  OR2_X1 U576 ( .A1(n18), .A2(key[119]), .ZN(n470) );
  AND2_X1 U577 ( .A1(key[119]), .A2(n18), .ZN(n469) );
  OR2_X1 U578 ( .A1(n471), .A2(n19), .ZN(out[118]) );
  OR2_X1 U579 ( .A1(n20), .A2(key[118]), .ZN(n472) );
  AND2_X1 U580 ( .A1(key[118]), .A2(n20), .ZN(n471) );
  OR2_X1 U581 ( .A1(n473), .A2(n21), .ZN(out[117]) );
  OR2_X1 U582 ( .A1(n22), .A2(key[117]), .ZN(n474) );
  AND2_X1 U583 ( .A1(key[117]), .A2(n22), .ZN(n473) );
  OR2_X1 U584 ( .A1(n475), .A2(n23), .ZN(out[116]) );
  OR2_X1 U585 ( .A1(n24), .A2(key[116]), .ZN(n476) );
  AND2_X1 U586 ( .A1(key[116]), .A2(n24), .ZN(n475) );
  OR2_X1 U587 ( .A1(n477), .A2(n25), .ZN(out[115]) );
  OR2_X1 U588 ( .A1(n26), .A2(key[115]), .ZN(n478) );
  AND2_X1 U589 ( .A1(key[115]), .A2(n26), .ZN(n477) );
  OR2_X1 U590 ( .A1(n479), .A2(n27), .ZN(out[114]) );
  OR2_X1 U591 ( .A1(n28), .A2(key[114]), .ZN(n480) );
  AND2_X1 U592 ( .A1(key[114]), .A2(n28), .ZN(n479) );
  OR2_X1 U593 ( .A1(n481), .A2(n29), .ZN(out[113]) );
  OR2_X1 U594 ( .A1(n30), .A2(key[113]), .ZN(n482) );
  AND2_X1 U595 ( .A1(key[113]), .A2(n30), .ZN(n481) );
  OR2_X1 U596 ( .A1(n483), .A2(n31), .ZN(out[112]) );
  OR2_X1 U597 ( .A1(n32), .A2(key[112]), .ZN(n484) );
  AND2_X1 U598 ( .A1(key[112]), .A2(n32), .ZN(n483) );
  OR2_X1 U599 ( .A1(n485), .A2(n33), .ZN(out[111]) );
  OR2_X1 U600 ( .A1(n34), .A2(key[111]), .ZN(n486) );
  AND2_X1 U601 ( .A1(key[111]), .A2(n34), .ZN(n485) );
  OR2_X1 U602 ( .A1(n487), .A2(n35), .ZN(out[110]) );
  OR2_X1 U603 ( .A1(n36), .A2(key[110]), .ZN(n488) );
  AND2_X1 U604 ( .A1(key[110]), .A2(n36), .ZN(n487) );
  OR2_X1 U605 ( .A1(n489), .A2(n235), .ZN(out[10]) );
  OR2_X1 U606 ( .A1(n236), .A2(key[10]), .ZN(n490) );
  AND2_X1 U607 ( .A1(key[10]), .A2(n236), .ZN(n489) );
  OR2_X1 U608 ( .A1(n491), .A2(n37), .ZN(out[109]) );
  OR2_X1 U609 ( .A1(n38), .A2(key[109]), .ZN(n492) );
  AND2_X1 U610 ( .A1(key[109]), .A2(n38), .ZN(n491) );
  OR2_X1 U611 ( .A1(n493), .A2(n39), .ZN(out[108]) );
  OR2_X1 U612 ( .A1(n40), .A2(key[108]), .ZN(n494) );
  AND2_X1 U613 ( .A1(key[108]), .A2(n40), .ZN(n493) );
  OR2_X1 U614 ( .A1(n495), .A2(n41), .ZN(out[107]) );
  OR2_X1 U615 ( .A1(n42), .A2(key[107]), .ZN(n496) );
  AND2_X1 U616 ( .A1(key[107]), .A2(n42), .ZN(n495) );
  OR2_X1 U617 ( .A1(n497), .A2(n43), .ZN(out[106]) );
  OR2_X1 U618 ( .A1(n44), .A2(key[106]), .ZN(n498) );
  AND2_X1 U619 ( .A1(key[106]), .A2(n44), .ZN(n497) );
  OR2_X1 U620 ( .A1(n499), .A2(n45), .ZN(out[105]) );
  OR2_X1 U621 ( .A1(n46), .A2(key[105]), .ZN(n500) );
  AND2_X1 U622 ( .A1(key[105]), .A2(n46), .ZN(n499) );
  OR2_X1 U623 ( .A1(n501), .A2(n47), .ZN(out[104]) );
  OR2_X1 U624 ( .A1(n48), .A2(key[104]), .ZN(n502) );
  AND2_X1 U625 ( .A1(key[104]), .A2(n48), .ZN(n501) );
  OR2_X1 U626 ( .A1(n503), .A2(n49), .ZN(out[103]) );
  OR2_X1 U627 ( .A1(n50), .A2(key[103]), .ZN(n504) );
  AND2_X1 U628 ( .A1(key[103]), .A2(n50), .ZN(n503) );
  OR2_X1 U629 ( .A1(n505), .A2(n51), .ZN(out[102]) );
  OR2_X1 U630 ( .A1(n52), .A2(key[102]), .ZN(n506) );
  AND2_X1 U631 ( .A1(key[102]), .A2(n52), .ZN(n505) );
  OR2_X1 U632 ( .A1(n507), .A2(n53), .ZN(out[101]) );
  OR2_X1 U633 ( .A1(n54), .A2(key[101]), .ZN(n508) );
  AND2_X1 U634 ( .A1(key[101]), .A2(n54), .ZN(n507) );
  OR2_X1 U635 ( .A1(n509), .A2(n55), .ZN(out[100]) );
  OR2_X1 U636 ( .A1(n56), .A2(key[100]), .ZN(n510) );
  AND2_X1 U637 ( .A1(key[100]), .A2(n56), .ZN(n509) );
  OR2_X1 U638 ( .A1(n511), .A2(n255), .ZN(out[0]) );
  OR2_X1 U639 ( .A1(n256), .A2(key[0]), .ZN(n512) );
  AND2_X1 U640 ( .A1(key[0]), .A2(n256), .ZN(n511) );
endmodule

//done